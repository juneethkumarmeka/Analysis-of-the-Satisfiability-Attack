module basic_2000_20000_2500_20_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nor U0 (N_0,In_1512,In_1665);
or U1 (N_1,In_473,In_1187);
nor U2 (N_2,In_1517,In_985);
or U3 (N_3,In_1253,In_971);
or U4 (N_4,In_220,In_329);
nand U5 (N_5,In_1513,In_71);
nand U6 (N_6,In_144,In_1149);
nor U7 (N_7,In_1293,In_64);
nor U8 (N_8,In_76,In_1976);
nor U9 (N_9,In_1762,In_1056);
nand U10 (N_10,In_1717,In_677);
and U11 (N_11,In_631,In_1090);
or U12 (N_12,In_1681,In_552);
nand U13 (N_13,In_791,In_1779);
nor U14 (N_14,In_1939,In_758);
or U15 (N_15,In_1643,In_1788);
nor U16 (N_16,In_1199,In_1395);
nor U17 (N_17,In_1520,In_799);
or U18 (N_18,In_1295,In_182);
nand U19 (N_19,In_1603,In_1749);
nand U20 (N_20,In_618,In_1221);
nand U21 (N_21,In_278,In_1725);
and U22 (N_22,In_448,In_164);
and U23 (N_23,In_514,In_1922);
and U24 (N_24,In_1871,In_613);
or U25 (N_25,In_1731,In_1503);
nand U26 (N_26,In_1605,In_700);
and U27 (N_27,In_731,In_1736);
nand U28 (N_28,In_578,In_795);
xor U29 (N_29,In_774,In_1884);
xnor U30 (N_30,In_1938,In_1078);
nand U31 (N_31,In_272,In_461);
nand U32 (N_32,In_1738,In_1458);
nand U33 (N_33,In_267,In_928);
xor U34 (N_34,In_1310,In_1373);
xor U35 (N_35,In_1836,In_1650);
nand U36 (N_36,In_995,In_1451);
and U37 (N_37,In_1008,In_279);
xor U38 (N_38,In_1421,In_1491);
nand U39 (N_39,In_401,In_1979);
nor U40 (N_40,In_1003,In_128);
or U41 (N_41,In_1761,In_907);
and U42 (N_42,In_1039,In_529);
or U43 (N_43,In_1120,In_1858);
xnor U44 (N_44,In_619,In_416);
or U45 (N_45,In_386,In_1046);
nand U46 (N_46,In_935,In_759);
nand U47 (N_47,In_1740,In_458);
nand U48 (N_48,In_1244,In_1473);
nand U49 (N_49,In_1264,In_185);
nor U50 (N_50,In_351,In_976);
or U51 (N_51,In_451,In_864);
nand U52 (N_52,In_1347,In_1812);
or U53 (N_53,In_992,In_286);
nand U54 (N_54,In_1019,In_150);
or U55 (N_55,In_38,In_270);
and U56 (N_56,In_1743,In_783);
nor U57 (N_57,In_1919,In_979);
or U58 (N_58,In_1125,In_813);
nor U59 (N_59,In_1455,In_1454);
or U60 (N_60,In_92,In_557);
nor U61 (N_61,In_443,In_1435);
nor U62 (N_62,In_1460,In_123);
or U63 (N_63,In_492,In_737);
nand U64 (N_64,In_512,In_1613);
nor U65 (N_65,In_273,In_1035);
nor U66 (N_66,In_404,In_1203);
xnor U67 (N_67,In_1990,In_1186);
nand U68 (N_68,In_1758,In_1929);
xor U69 (N_69,In_866,In_1882);
and U70 (N_70,In_1096,In_1289);
nor U71 (N_71,In_318,In_441);
xor U72 (N_72,In_407,In_491);
or U73 (N_73,In_1196,In_603);
and U74 (N_74,In_1769,In_895);
and U75 (N_75,In_1972,In_1072);
or U76 (N_76,In_1341,In_1070);
xor U77 (N_77,In_103,In_599);
nand U78 (N_78,In_1658,In_434);
nor U79 (N_79,In_753,In_1076);
or U80 (N_80,In_859,In_586);
and U81 (N_81,In_565,In_1278);
nand U82 (N_82,In_1813,In_35);
or U83 (N_83,In_1181,In_1291);
xnor U84 (N_84,In_1870,In_1826);
xnor U85 (N_85,In_1036,In_208);
xor U86 (N_86,In_422,In_236);
nand U87 (N_87,In_176,In_636);
and U88 (N_88,In_348,In_14);
xor U89 (N_89,In_1168,In_1504);
xnor U90 (N_90,In_912,In_1702);
and U91 (N_91,In_1055,In_1638);
nor U92 (N_92,In_913,In_1062);
and U93 (N_93,In_1415,In_1669);
or U94 (N_94,In_710,In_956);
nor U95 (N_95,In_166,In_453);
xor U96 (N_96,In_151,In_1950);
or U97 (N_97,In_777,In_1251);
nor U98 (N_98,In_349,In_1551);
nor U99 (N_99,In_1941,In_1560);
nor U100 (N_100,In_261,In_931);
nand U101 (N_101,In_1479,In_518);
or U102 (N_102,In_1250,In_1607);
nand U103 (N_103,In_1143,In_688);
and U104 (N_104,In_1766,In_477);
or U105 (N_105,In_1686,In_1688);
nand U106 (N_106,In_1350,In_967);
and U107 (N_107,In_1904,In_1084);
nor U108 (N_108,In_548,In_199);
and U109 (N_109,In_104,In_666);
or U110 (N_110,In_516,In_689);
nor U111 (N_111,In_1424,In_732);
xnor U112 (N_112,In_934,In_314);
nand U113 (N_113,In_1441,In_446);
nand U114 (N_114,In_1527,In_232);
xor U115 (N_115,In_852,In_1069);
nand U116 (N_116,In_889,In_1022);
nor U117 (N_117,In_1881,In_583);
nand U118 (N_118,In_1058,In_1034);
xnor U119 (N_119,In_133,In_471);
nand U120 (N_120,In_887,In_553);
or U121 (N_121,In_1127,In_1949);
and U122 (N_122,In_1600,In_1068);
and U123 (N_123,In_1618,In_41);
xnor U124 (N_124,In_1486,In_886);
nor U125 (N_125,In_1173,In_880);
xnor U126 (N_126,In_69,In_1422);
nand U127 (N_127,In_1419,In_1396);
nand U128 (N_128,In_1511,In_1846);
or U129 (N_129,In_1098,In_1863);
xnor U130 (N_130,In_1727,In_85);
and U131 (N_131,In_997,In_1151);
xor U132 (N_132,In_499,In_87);
and U133 (N_133,In_233,In_1053);
and U134 (N_134,In_789,In_1225);
and U135 (N_135,In_1741,In_1585);
and U136 (N_136,In_853,In_1557);
nand U137 (N_137,In_1693,In_1617);
and U138 (N_138,In_277,In_1087);
and U139 (N_139,In_1452,In_1228);
or U140 (N_140,In_860,In_1909);
or U141 (N_141,In_1420,In_307);
nand U142 (N_142,In_322,In_89);
or U143 (N_143,In_345,In_498);
nand U144 (N_144,In_174,In_1796);
and U145 (N_145,In_709,In_1483);
or U146 (N_146,In_544,In_537);
and U147 (N_147,In_1880,In_243);
or U148 (N_148,In_447,In_1208);
and U149 (N_149,In_1166,In_340);
or U150 (N_150,In_496,In_1450);
nor U151 (N_151,In_1664,In_1940);
or U152 (N_152,In_452,In_156);
or U153 (N_153,In_1163,In_36);
or U154 (N_154,In_316,In_896);
nor U155 (N_155,In_1771,In_78);
nand U156 (N_156,In_1633,In_1204);
xnor U157 (N_157,In_23,In_1349);
nor U158 (N_158,In_1367,In_414);
or U159 (N_159,In_1694,In_122);
nand U160 (N_160,In_258,In_531);
nor U161 (N_161,In_1254,In_254);
or U162 (N_162,In_20,In_1885);
nand U163 (N_163,In_1237,In_1108);
nand U164 (N_164,In_1869,In_659);
nor U165 (N_165,In_558,In_1382);
and U166 (N_166,In_1953,In_1780);
or U167 (N_167,In_1328,In_223);
nand U168 (N_168,In_1215,In_1621);
nand U169 (N_169,In_1948,In_765);
nand U170 (N_170,In_1436,In_707);
nand U171 (N_171,In_456,In_1908);
xor U172 (N_172,In_53,In_139);
nor U173 (N_173,In_1141,In_1878);
xnor U174 (N_174,In_1864,In_399);
xnor U175 (N_175,In_1839,In_1002);
xnor U176 (N_176,In_1958,In_1263);
nand U177 (N_177,In_1247,In_1890);
nand U178 (N_178,In_902,In_773);
xor U179 (N_179,In_1509,In_1113);
or U180 (N_180,In_385,In_1932);
nand U181 (N_181,In_1645,In_428);
nor U182 (N_182,In_409,In_1730);
nor U183 (N_183,In_1245,In_980);
nor U184 (N_184,In_336,In_292);
and U185 (N_185,In_1841,In_59);
nand U186 (N_186,In_948,In_61);
nor U187 (N_187,In_382,In_1623);
or U188 (N_188,In_1066,In_478);
xnor U189 (N_189,In_1728,In_682);
nand U190 (N_190,In_1021,In_648);
nand U191 (N_191,In_93,In_1652);
nand U192 (N_192,In_1593,In_1057);
and U193 (N_193,In_1032,In_770);
xnor U194 (N_194,In_1624,In_160);
nor U195 (N_195,In_939,In_1162);
and U196 (N_196,In_925,In_952);
nand U197 (N_197,In_1115,In_1249);
or U198 (N_198,In_1538,In_1029);
xnor U199 (N_199,In_175,In_1789);
xnor U200 (N_200,In_217,In_1256);
nand U201 (N_201,In_1609,In_354);
nand U202 (N_202,In_1447,In_16);
xnor U203 (N_203,In_1272,In_1378);
and U204 (N_204,In_60,In_380);
nor U205 (N_205,In_624,In_660);
nand U206 (N_206,In_1033,In_1260);
nand U207 (N_207,In_1442,In_906);
or U208 (N_208,In_429,In_1357);
or U209 (N_209,In_867,In_405);
and U210 (N_210,In_642,In_417);
nor U211 (N_211,In_127,In_803);
xnor U212 (N_212,In_854,In_432);
or U213 (N_213,In_413,In_847);
nand U214 (N_214,In_1480,In_67);
nand U215 (N_215,In_1594,In_605);
xor U216 (N_216,In_357,In_403);
or U217 (N_217,In_1611,In_1872);
nor U218 (N_218,In_840,In_1676);
and U219 (N_219,In_198,In_1267);
or U220 (N_220,In_324,In_1768);
or U221 (N_221,In_1970,In_1964);
nor U222 (N_222,In_262,In_1161);
xnor U223 (N_223,In_330,In_766);
or U224 (N_224,In_1967,In_724);
or U225 (N_225,In_489,In_844);
nand U226 (N_226,In_309,In_615);
nand U227 (N_227,In_1377,In_595);
or U228 (N_228,In_776,In_226);
nand U229 (N_229,In_589,In_1052);
nor U230 (N_230,In_58,In_520);
and U231 (N_231,In_426,In_398);
xnor U232 (N_232,In_1923,In_579);
or U233 (N_233,In_1490,In_1584);
and U234 (N_234,In_242,In_1816);
nor U235 (N_235,In_505,In_344);
nor U236 (N_236,In_37,In_1038);
xor U237 (N_237,In_1365,In_1227);
xor U238 (N_238,In_374,In_717);
nor U239 (N_239,In_821,In_1670);
and U240 (N_240,In_1041,In_1531);
nand U241 (N_241,In_1942,In_944);
or U242 (N_242,In_989,In_356);
nand U243 (N_243,In_1193,In_362);
or U244 (N_244,In_1859,In_1156);
or U245 (N_245,In_1756,In_8);
and U246 (N_246,In_1580,In_1887);
xor U247 (N_247,In_1380,In_1499);
nor U248 (N_248,In_1317,In_378);
xnor U249 (N_249,In_525,In_1945);
nand U250 (N_250,In_384,In_1918);
or U251 (N_251,In_188,In_1514);
and U252 (N_252,In_805,In_921);
xnor U253 (N_253,In_559,In_360);
xor U254 (N_254,In_305,In_1656);
or U255 (N_255,In_99,In_1361);
or U256 (N_256,In_869,In_1793);
xor U257 (N_257,In_381,In_898);
xnor U258 (N_258,In_650,In_1854);
xor U259 (N_259,In_146,In_706);
xor U260 (N_260,In_1842,In_115);
xor U261 (N_261,In_825,In_159);
and U262 (N_262,In_5,In_1901);
and U263 (N_263,In_1719,In_1674);
xnor U264 (N_264,In_874,In_4);
nor U265 (N_265,In_301,In_410);
nor U266 (N_266,In_1927,In_269);
or U267 (N_267,In_511,In_1372);
nor U268 (N_268,In_500,In_297);
or U269 (N_269,In_1523,In_890);
nand U270 (N_270,In_1238,In_1448);
and U271 (N_271,In_1210,In_1586);
xor U272 (N_272,In_173,In_622);
and U273 (N_273,In_1540,In_1700);
nor U274 (N_274,In_1660,In_810);
nand U275 (N_275,In_756,In_1651);
xor U276 (N_276,In_1860,In_392);
and U277 (N_277,In_457,In_210);
or U278 (N_278,In_1331,In_1018);
nand U279 (N_279,In_24,In_408);
and U280 (N_280,In_1131,In_377);
xor U281 (N_281,In_1539,In_1006);
nor U282 (N_282,In_721,In_321);
and U283 (N_283,In_519,In_1985);
nor U284 (N_284,In_1801,In_1308);
nand U285 (N_285,In_481,In_1152);
and U286 (N_286,In_504,In_730);
and U287 (N_287,In_665,In_515);
xor U288 (N_288,In_1902,In_943);
xnor U289 (N_289,In_207,In_466);
or U290 (N_290,In_1067,In_800);
nor U291 (N_291,In_1074,In_332);
or U292 (N_292,In_1266,In_1031);
nor U293 (N_293,In_1235,In_694);
nand U294 (N_294,In_1246,In_1677);
xnor U295 (N_295,In_1588,In_568);
or U296 (N_296,In_1012,In_1508);
nor U297 (N_297,In_667,In_1489);
or U298 (N_298,In_1843,In_1192);
xor U299 (N_299,In_1202,In_891);
xor U300 (N_300,In_645,In_657);
xor U301 (N_301,In_888,In_1576);
xnor U302 (N_302,In_1099,In_1433);
nand U303 (N_303,In_222,In_849);
nand U304 (N_304,In_170,In_388);
and U305 (N_305,In_1464,In_1834);
nor U306 (N_306,In_1568,In_655);
nand U307 (N_307,In_1616,In_1195);
xnor U308 (N_308,In_1716,In_1696);
nand U309 (N_309,In_1821,In_1574);
and U310 (N_310,In_1386,In_291);
nand U311 (N_311,In_1476,In_1234);
and U312 (N_312,In_1262,In_1122);
or U313 (N_313,In_812,In_1402);
and U314 (N_314,In_397,In_479);
xor U315 (N_315,In_317,In_740);
xor U316 (N_316,In_1144,In_158);
nand U317 (N_317,In_1376,In_627);
xor U318 (N_318,In_1971,In_289);
xnor U319 (N_319,In_1800,In_977);
or U320 (N_320,In_206,In_969);
and U321 (N_321,In_1528,In_1537);
or U322 (N_322,In_1059,In_33);
or U323 (N_323,In_590,In_1370);
nand U324 (N_324,In_135,In_626);
and U325 (N_325,In_1969,In_1627);
xor U326 (N_326,In_1240,In_959);
nand U327 (N_327,In_858,In_244);
and U328 (N_328,In_1086,In_990);
and U329 (N_329,In_112,In_729);
xnor U330 (N_330,In_1760,In_335);
or U331 (N_331,In_364,In_1371);
nor U332 (N_332,In_1129,In_264);
and U333 (N_333,In_1981,In_1270);
nor U334 (N_334,In_1984,In_1430);
xor U335 (N_335,In_1484,In_922);
or U336 (N_336,In_521,In_1468);
xnor U337 (N_337,In_1023,In_1207);
or U338 (N_338,In_1304,In_1493);
xor U339 (N_339,In_179,In_1094);
xor U340 (N_340,In_100,In_543);
nor U341 (N_341,In_1185,In_459);
nor U342 (N_342,In_978,In_83);
or U343 (N_343,In_1720,In_440);
nand U344 (N_344,In_63,In_787);
or U345 (N_345,In_1481,In_882);
nand U346 (N_346,In_247,In_12);
nor U347 (N_347,In_121,In_567);
nor U348 (N_348,In_1427,In_856);
xor U349 (N_349,In_780,In_1340);
or U350 (N_350,In_1721,In_1722);
nand U351 (N_351,In_1437,In_284);
or U352 (N_352,In_1492,In_1963);
xnor U353 (N_353,In_1861,In_1510);
nor U354 (N_354,In_285,In_708);
or U355 (N_355,In_960,In_555);
nor U356 (N_356,In_835,In_562);
or U357 (N_357,In_651,In_1114);
nand U358 (N_358,In_862,In_387);
xnor U359 (N_359,In_1906,In_1502);
xnor U360 (N_360,In_750,In_1577);
xor U361 (N_361,In_157,In_1282);
xor U362 (N_362,In_1302,In_1867);
and U363 (N_363,In_972,In_1243);
and U364 (N_364,In_253,In_1751);
or U365 (N_365,In_124,In_534);
and U366 (N_366,In_302,In_57);
xnor U367 (N_367,In_1232,In_393);
xor U368 (N_368,In_1935,In_926);
nand U369 (N_369,In_577,In_695);
xor U370 (N_370,In_798,In_716);
and U371 (N_371,In_1271,In_1824);
and U372 (N_372,In_355,In_1176);
nand U373 (N_373,In_1578,In_30);
or U374 (N_374,In_1414,In_621);
or U375 (N_375,In_1729,In_1345);
or U376 (N_376,In_674,In_1092);
nand U377 (N_377,In_987,In_342);
nand U378 (N_378,In_1020,In_575);
or U379 (N_379,In_1145,In_1525);
nand U380 (N_380,In_234,In_1024);
nor U381 (N_381,In_1184,In_1288);
and U382 (N_382,In_1432,In_299);
nor U383 (N_383,In_1817,In_1147);
xnor U384 (N_384,In_1679,In_171);
xor U385 (N_385,In_1209,In_1339);
and U386 (N_386,In_480,In_1505);
nand U387 (N_387,In_1191,In_796);
nor U388 (N_388,In_1283,In_701);
nand U389 (N_389,In_450,In_1853);
nor U390 (N_390,In_1966,In_230);
nor U391 (N_391,In_1912,In_1258);
xor U392 (N_392,In_312,In_346);
nand U393 (N_393,In_1487,In_1628);
and U394 (N_394,In_110,In_1672);
nor U395 (N_395,In_193,In_1892);
nand U396 (N_396,In_546,In_1255);
nor U397 (N_397,In_963,In_1978);
or U398 (N_398,In_1564,In_1599);
or U399 (N_399,In_1390,In_506);
xor U400 (N_400,In_493,In_29);
or U401 (N_401,In_1873,In_488);
xor U402 (N_402,In_231,In_871);
nand U403 (N_403,In_975,In_1591);
xor U404 (N_404,In_1274,In_1429);
and U405 (N_405,In_1004,In_804);
nor U406 (N_406,In_116,In_1354);
nor U407 (N_407,In_472,In_1913);
nor U408 (N_408,In_1200,In_319);
and U409 (N_409,In_539,In_1589);
or U410 (N_410,In_1194,In_591);
xor U411 (N_411,In_98,In_161);
or U412 (N_412,In_1412,In_1954);
xor U413 (N_413,In_190,In_154);
and U414 (N_414,In_17,In_957);
nor U415 (N_415,In_955,In_715);
or U416 (N_416,In_837,In_111);
and U417 (N_417,In_581,In_1811);
xor U418 (N_418,In_245,In_215);
nor U419 (N_419,In_201,In_21);
nand U420 (N_420,In_711,In_1037);
xnor U421 (N_421,In_1685,In_746);
nand U422 (N_422,In_930,In_1883);
or U423 (N_423,In_1543,In_415);
nor U424 (N_424,In_1417,In_1797);
and U425 (N_425,In_109,In_771);
or U426 (N_426,In_1825,In_1103);
nor U427 (N_427,In_282,In_361);
xor U428 (N_428,In_663,In_870);
or U429 (N_429,In_80,In_1522);
nand U430 (N_430,In_691,In_1947);
or U431 (N_431,In_1975,In_547);
xnor U432 (N_432,In_108,In_634);
nor U433 (N_433,In_892,In_1351);
nor U434 (N_434,In_596,In_542);
nand U435 (N_435,In_741,In_418);
xnor U436 (N_436,In_431,In_34);
or U437 (N_437,In_917,In_266);
nor U438 (N_438,In_95,In_1818);
xnor U439 (N_439,In_1790,In_1900);
xor U440 (N_440,In_1159,In_830);
nand U441 (N_441,In_1044,In_1307);
or U442 (N_442,In_467,In_1561);
nor U443 (N_443,In_40,In_315);
nor U444 (N_444,In_1991,In_1368);
xor U445 (N_445,In_637,In_1983);
nor U446 (N_446,In_1553,In_827);
nor U447 (N_447,In_617,In_1748);
or U448 (N_448,In_1026,In_1358);
and U449 (N_449,In_439,In_1968);
nor U450 (N_450,In_824,In_1786);
xor U451 (N_451,In_1905,In_368);
nand U452 (N_452,In_72,In_1172);
or U453 (N_453,In_1093,In_949);
or U454 (N_454,In_1635,In_1301);
nand U455 (N_455,In_1726,In_1496);
nand U456 (N_456,In_358,In_683);
or U457 (N_457,In_216,In_1010);
nand U458 (N_458,In_1027,In_742);
or U459 (N_459,In_1851,In_1279);
xnor U460 (N_460,In_927,In_748);
nand U461 (N_461,In_1040,In_1169);
and U462 (N_462,In_1899,In_1408);
and U463 (N_463,In_1257,In_1292);
xnor U464 (N_464,In_712,In_1362);
nand U465 (N_465,In_778,In_1494);
nand U466 (N_466,In_495,In_736);
or U467 (N_467,In_1875,In_1852);
and U468 (N_468,In_52,In_549);
xnor U469 (N_469,In_1164,In_755);
or U470 (N_470,In_962,In_1682);
nor U471 (N_471,In_1545,In_640);
and U472 (N_472,In_788,In_1847);
nand U473 (N_473,In_1774,In_1581);
nor U474 (N_474,In_564,In_1356);
xnor U475 (N_475,In_296,In_1897);
or U476 (N_476,In_685,In_761);
nor U477 (N_477,In_1703,In_81);
and U478 (N_478,In_1868,In_875);
nor U479 (N_479,In_1265,In_936);
xnor U480 (N_480,In_527,In_576);
nand U481 (N_481,In_1737,In_968);
or U482 (N_482,In_1467,In_509);
xnor U483 (N_483,In_1742,In_834);
nand U484 (N_484,In_1575,In_945);
nor U485 (N_485,In_705,In_1724);
or U486 (N_486,In_1081,In_1776);
xor U487 (N_487,In_1907,In_106);
xor U488 (N_488,In_1423,In_1404);
or U489 (N_489,In_240,In_1973);
nor U490 (N_490,In_923,In_1832);
and U491 (N_491,In_363,In_1444);
and U492 (N_492,In_1844,In_460);
xor U493 (N_493,In_1992,In_1625);
nor U494 (N_494,In_768,In_718);
nor U495 (N_495,In_1360,In_684);
nor U496 (N_496,In_1876,In_904);
and U497 (N_497,In_427,In_1587);
xnor U498 (N_498,In_625,In_313);
nor U499 (N_499,In_713,In_359);
xnor U500 (N_500,In_1285,In_47);
nor U501 (N_501,In_1001,In_463);
xor U502 (N_502,In_352,In_1795);
xnor U503 (N_503,In_1445,In_246);
xnor U504 (N_504,In_219,In_1515);
or U505 (N_505,In_785,In_672);
nand U506 (N_506,In_181,In_1562);
xnor U507 (N_507,In_1710,In_900);
nor U508 (N_508,In_396,In_1405);
nor U509 (N_509,In_353,In_592);
and U510 (N_510,In_86,In_1112);
or U511 (N_511,In_74,In_879);
and U512 (N_512,In_79,In_823);
nor U513 (N_513,In_1898,In_1951);
or U514 (N_514,In_1337,In_1640);
nor U515 (N_515,In_1312,In_1190);
nand U516 (N_516,In_423,In_911);
nand U517 (N_517,In_1268,In_999);
xnor U518 (N_518,In_449,In_1309);
nand U519 (N_519,In_196,In_1431);
and U520 (N_520,In_738,In_702);
xor U521 (N_521,In_339,In_1111);
and U522 (N_522,In_268,In_46);
and U523 (N_523,In_1461,In_1217);
xnor U524 (N_524,In_438,In_1140);
xor U525 (N_525,In_503,In_1381);
xnor U526 (N_526,In_1644,In_350);
and U527 (N_527,In_1698,In_1558);
and U528 (N_528,In_1182,In_1222);
nand U529 (N_529,In_195,In_1833);
nand U530 (N_530,In_1383,In_1903);
and U531 (N_531,In_661,In_727);
xnor U532 (N_532,In_692,In_211);
nor U533 (N_533,In_669,In_1687);
nand U534 (N_534,In_1691,In_563);
nand U535 (N_535,In_752,In_229);
nand U536 (N_536,In_251,In_1782);
nand U537 (N_537,In_836,In_1343);
or U538 (N_538,In_1223,In_1178);
nand U539 (N_539,In_981,In_833);
xor U540 (N_540,In_1952,In_25);
xnor U541 (N_541,In_1016,In_885);
nor U542 (N_542,In_723,In_1808);
xnor U543 (N_543,In_275,In_250);
or U544 (N_544,In_1359,In_1128);
nor U545 (N_545,In_1342,In_1709);
xnor U546 (N_546,In_187,In_1596);
nand U547 (N_547,In_1746,In_1226);
and U548 (N_548,In_602,In_1230);
nor U549 (N_549,In_1572,In_806);
nor U550 (N_550,In_391,In_1100);
xnor U551 (N_551,In_545,In_507);
and U552 (N_552,In_125,In_802);
or U553 (N_553,In_9,In_1849);
xnor U554 (N_554,In_1472,In_1158);
xor U555 (N_555,In_1891,In_94);
nor U556 (N_556,In_832,In_1697);
nor U557 (N_557,In_1711,In_628);
or U558 (N_558,In_829,In_126);
xnor U559 (N_559,In_337,In_485);
nand U560 (N_560,In_55,In_1840);
xnor U561 (N_561,In_676,In_1582);
nor U562 (N_562,In_897,In_1048);
and U563 (N_563,In_878,In_1583);
nand U564 (N_564,In_1809,In_1705);
nor U565 (N_565,In_117,In_256);
nand U566 (N_566,In_1798,In_1105);
xnor U567 (N_567,In_508,In_1661);
nand U568 (N_568,In_323,In_1936);
nor U569 (N_569,In_1025,In_1205);
nand U570 (N_570,In_745,In_143);
and U571 (N_571,In_1955,In_113);
and U572 (N_572,In_420,In_1418);
or U573 (N_573,In_697,In_97);
nor U574 (N_574,In_1475,In_826);
nand U575 (N_575,In_366,In_419);
nor U576 (N_576,In_91,In_1773);
or U577 (N_577,In_1219,In_486);
and U578 (N_578,In_1061,In_1626);
xnor U579 (N_579,In_287,In_1180);
nand U580 (N_580,In_865,In_1095);
nor U581 (N_581,In_1662,In_162);
or U582 (N_582,In_1639,In_88);
xor U583 (N_583,In_845,In_749);
and U584 (N_584,In_1119,In_894);
nor U585 (N_585,In_476,In_1313);
and U586 (N_586,In_881,In_526);
nand U587 (N_587,In_1242,In_1287);
nand U588 (N_588,In_15,In_1474);
xor U589 (N_589,In_54,In_877);
nor U590 (N_590,In_1154,In_1831);
xnor U591 (N_591,In_169,In_212);
nor U592 (N_592,In_105,In_1043);
nand U593 (N_593,In_940,In_670);
nor U594 (N_594,In_1957,In_237);
nand U595 (N_595,In_1425,In_1387);
or U596 (N_596,In_908,In_793);
nand U597 (N_597,In_152,In_818);
xor U598 (N_598,In_1252,In_141);
xor U599 (N_599,In_1783,In_373);
or U600 (N_600,In_982,In_996);
nor U601 (N_601,In_1735,In_914);
xor U602 (N_602,In_177,In_1322);
or U603 (N_603,In_1374,In_654);
xnor U604 (N_604,In_1007,In_1236);
xor U605 (N_605,In_214,In_13);
nor U606 (N_606,In_1174,In_1914);
nor U607 (N_607,In_1073,In_389);
or U608 (N_608,In_1428,In_790);
xnor U609 (N_609,In_114,In_375);
and U610 (N_610,In_1280,In_681);
or U611 (N_611,In_772,In_1759);
xnor U612 (N_612,In_1916,In_1498);
xnor U613 (N_613,In_1713,In_1439);
and U614 (N_614,In_1071,In_1284);
xor U615 (N_615,In_1647,In_1353);
or U616 (N_616,In_1530,In_1045);
xnor U617 (N_617,In_11,In_227);
nand U618 (N_618,In_966,In_1352);
nand U619 (N_619,In_300,In_490);
or U620 (N_620,In_280,In_899);
or U621 (N_621,In_1315,In_129);
nor U622 (N_622,In_961,In_1311);
xnor U623 (N_623,In_1324,In_1364);
and U624 (N_624,In_1534,In_1657);
xnor U625 (N_625,In_1675,In_1273);
xor U626 (N_626,In_131,In_1535);
or U627 (N_627,In_1877,In_1465);
nor U628 (N_628,In_1133,In_1126);
or U629 (N_629,In_1079,In_1329);
and U630 (N_630,In_964,In_551);
and U631 (N_631,In_205,In_1463);
and U632 (N_632,In_255,In_238);
or U633 (N_633,In_1920,In_1326);
nand U634 (N_634,In_809,In_998);
nor U635 (N_635,In_142,In_1699);
and U636 (N_636,In_183,In_1519);
nand U637 (N_637,In_1456,In_1388);
nand U638 (N_638,In_462,In_1000);
nor U639 (N_639,In_454,In_1107);
nor U640 (N_640,In_376,In_331);
nor U641 (N_641,In_1830,In_394);
nor U642 (N_642,In_612,In_1893);
nand U643 (N_643,In_580,In_1977);
nor U644 (N_644,In_739,In_271);
nor U645 (N_645,In_1369,In_1690);
nor U646 (N_646,In_1110,In_1139);
xnor U647 (N_647,In_533,In_1556);
and U648 (N_648,In_1471,In_598);
or U649 (N_649,In_1521,In_1518);
nand U650 (N_650,In_1453,In_1765);
xor U651 (N_651,In_638,In_747);
or U652 (N_652,In_538,In_1366);
and U653 (N_653,In_1838,In_569);
or U654 (N_654,In_1438,In_283);
xnor U655 (N_655,In_973,In_1506);
nor U656 (N_656,In_1116,In_1397);
xnor U657 (N_657,In_1874,In_986);
or U658 (N_658,In_1410,In_1684);
or U659 (N_659,In_828,In_1197);
xor U660 (N_660,In_635,In_1379);
nand U661 (N_661,In_425,In_304);
and U662 (N_662,In_876,In_1541);
or U663 (N_663,In_325,In_775);
and U664 (N_664,In_1469,In_633);
and U665 (N_665,In_673,In_1784);
xor U666 (N_666,In_194,In_1548);
xor U667 (N_667,In_1363,In_561);
and U668 (N_668,In_1297,In_1822);
xnor U669 (N_669,In_137,In_1138);
nor U670 (N_670,In_1054,In_556);
and U671 (N_671,In_1188,In_929);
xor U672 (N_672,In_497,In_696);
nand U673 (N_673,In_1298,In_42);
xor U674 (N_674,In_1764,In_1495);
nor U675 (N_675,In_733,In_77);
nor U676 (N_676,In_442,In_958);
and U677 (N_677,In_1346,In_372);
or U678 (N_678,In_1529,In_1987);
nor U679 (N_679,In_1355,In_1015);
xor U680 (N_680,In_167,In_1526);
or U681 (N_681,In_1241,In_1654);
nand U682 (N_682,In_1928,In_764);
nand U683 (N_683,In_412,In_1999);
and U684 (N_684,In_82,In_1049);
nor U685 (N_685,In_1986,In_402);
and U686 (N_686,In_1316,In_184);
or U687 (N_687,In_720,In_690);
or U688 (N_688,In_73,In_1921);
and U689 (N_689,In_1733,In_1142);
nor U690 (N_690,In_1629,In_1201);
xor U691 (N_691,In_1837,In_1524);
and U692 (N_692,In_797,In_1739);
xnor U693 (N_693,In_1106,In_993);
xnor U694 (N_694,In_680,In_1804);
and U695 (N_695,In_464,In_1478);
nor U696 (N_696,In_937,In_298);
and U697 (N_697,In_610,In_18);
and U698 (N_698,In_1167,In_1663);
and U699 (N_699,In_180,In_754);
or U700 (N_700,In_148,In_1013);
or U701 (N_701,In_751,In_550);
nor U702 (N_702,In_1183,In_1763);
or U703 (N_703,In_916,In_1413);
nand U704 (N_704,In_842,In_1745);
and U705 (N_705,In_1075,In_1636);
and U706 (N_706,In_1695,In_991);
nor U707 (N_707,In_646,In_851);
or U708 (N_708,In_45,In_1989);
xor U709 (N_709,In_186,In_1286);
nand U710 (N_710,In_484,In_75);
or U711 (N_711,In_168,In_1641);
and U712 (N_712,In_781,In_1532);
nor U713 (N_713,In_252,In_1715);
nor U714 (N_714,In_469,In_395);
and U715 (N_715,In_483,In_1211);
xnor U716 (N_716,In_1409,In_915);
xnor U717 (N_717,In_792,In_1933);
or U718 (N_718,In_153,In_1101);
nand U719 (N_719,In_406,In_3);
nand U720 (N_720,In_1806,In_763);
xnor U721 (N_721,In_1931,In_1233);
xnor U722 (N_722,In_1384,In_371);
xor U723 (N_723,In_257,In_474);
xnor U724 (N_724,In_1604,In_248);
xor U725 (N_725,In_1823,In_1017);
nand U726 (N_726,In_192,In_138);
and U727 (N_727,In_1065,In_857);
nor U728 (N_728,In_288,In_1886);
or U729 (N_729,In_530,In_1091);
nand U730 (N_730,In_213,In_524);
xnor U731 (N_731,In_1118,In_260);
or U732 (N_732,In_1224,In_988);
xor U733 (N_733,In_873,In_1109);
nor U734 (N_734,In_510,In_1622);
or U735 (N_735,In_259,In_1982);
and U736 (N_736,In_517,In_1894);
xor U737 (N_737,In_1206,In_719);
xnor U738 (N_738,In_611,In_1212);
and U739 (N_739,In_1177,In_1121);
xor U740 (N_740,In_1637,In_411);
xnor U741 (N_741,In_1778,In_1767);
or U742 (N_742,In_686,In_22);
or U743 (N_743,In_1642,In_698);
nor U744 (N_744,In_265,In_1136);
nand U745 (N_745,In_1189,In_652);
or U746 (N_746,In_1117,In_1965);
and U747 (N_747,In_767,In_1426);
and U748 (N_748,In_872,In_585);
or U749 (N_749,In_574,In_1175);
nand U750 (N_750,In_893,In_850);
or U751 (N_751,In_1124,In_241);
and U752 (N_752,In_1393,In_919);
and U753 (N_753,In_1895,In_1544);
nor U754 (N_754,In_1485,In_436);
nand U755 (N_755,In_228,In_1802);
or U756 (N_756,In_1501,In_32);
nor U757 (N_757,In_6,In_1807);
xnor U758 (N_758,In_1239,In_132);
xor U759 (N_759,In_1327,In_1835);
or U760 (N_760,In_1275,In_841);
nor U761 (N_761,In_224,In_1632);
xor U762 (N_762,In_1888,In_347);
or U763 (N_763,In_1259,In_600);
nand U764 (N_764,In_7,In_1500);
nand U765 (N_765,In_1827,In_704);
xnor U766 (N_766,In_1082,In_235);
nand U767 (N_767,In_933,In_263);
and U768 (N_768,In_1411,In_90);
xor U769 (N_769,In_584,In_1792);
nand U770 (N_770,In_468,In_1446);
and U771 (N_771,In_1334,In_725);
and U772 (N_772,In_1457,In_1962);
nand U773 (N_773,In_1290,In_831);
or U774 (N_774,In_572,In_1064);
nor U775 (N_775,In_333,In_941);
nand U776 (N_776,In_31,In_699);
nor U777 (N_777,In_1879,In_808);
nor U778 (N_778,In_1299,In_1335);
xnor U779 (N_779,In_820,In_1009);
nor U780 (N_780,In_814,In_1610);
xnor U781 (N_781,In_1595,In_1862);
xor U782 (N_782,In_341,In_593);
or U783 (N_783,In_1961,In_1546);
nand U784 (N_784,In_1104,In_1130);
nor U785 (N_785,In_221,In_1592);
nand U786 (N_786,In_1406,In_1631);
and U787 (N_787,In_465,In_616);
xnor U788 (N_788,In_1889,In_310);
nand U789 (N_789,In_1567,In_942);
nor U790 (N_790,In_1554,In_365);
nand U791 (N_791,In_1338,In_1323);
and U792 (N_792,In_1753,In_1559);
nand U793 (N_793,In_1943,In_433);
and U794 (N_794,In_369,In_1281);
and U795 (N_795,In_1856,In_421);
or U796 (N_796,In_1750,In_249);
or U797 (N_797,In_664,In_1815);
or U798 (N_798,In_290,In_1718);
or U799 (N_799,In_178,In_1723);
nor U800 (N_800,In_70,In_51);
and U801 (N_801,In_984,In_1294);
and U802 (N_802,In_294,In_643);
nand U803 (N_803,In_430,In_807);
and U804 (N_804,In_536,In_136);
xnor U805 (N_805,In_49,In_1566);
xnor U806 (N_806,In_1988,In_487);
xnor U807 (N_807,In_757,In_1403);
or U808 (N_808,In_1011,In_1590);
or U809 (N_809,In_1330,In_43);
xnor U810 (N_810,In_470,In_101);
and U811 (N_811,In_1319,In_970);
xor U812 (N_812,In_1956,In_145);
or U813 (N_813,In_649,In_1896);
xor U814 (N_814,In_1655,In_1305);
or U815 (N_815,In_1994,In_769);
and U816 (N_816,In_1570,In_1997);
and U817 (N_817,In_909,In_1198);
nor U818 (N_818,In_1602,In_200);
nor U819 (N_819,In_606,In_1137);
nand U820 (N_820,In_1946,In_1787);
xor U821 (N_821,In_1555,In_370);
nor U822 (N_822,In_784,In_535);
nand U823 (N_823,In_1819,In_1276);
nor U824 (N_824,In_320,In_597);
nor U825 (N_825,In_1980,In_1333);
xor U826 (N_826,In_1416,In_1649);
or U827 (N_827,In_96,In_1550);
or U828 (N_828,In_1218,In_1704);
xor U829 (N_829,In_1277,In_27);
and U830 (N_830,In_938,In_1440);
xnor U831 (N_831,In_1348,In_1400);
nand U832 (N_832,In_1634,In_400);
nand U833 (N_833,In_817,In_1959);
or U834 (N_834,In_614,In_1085);
and U835 (N_835,In_1216,In_1375);
xor U836 (N_836,In_1732,In_608);
nand U837 (N_837,In_445,In_1300);
xnor U838 (N_838,In_1088,In_130);
nor U839 (N_839,In_306,In_1320);
nand U840 (N_840,In_1781,In_1855);
or U841 (N_841,In_629,In_522);
nor U842 (N_842,In_1042,In_165);
or U843 (N_843,In_641,In_609);
and U844 (N_844,In_953,In_1332);
xor U845 (N_845,In_779,In_191);
and U846 (N_846,In_839,In_760);
xor U847 (N_847,In_1993,In_140);
or U848 (N_848,In_946,In_647);
or U849 (N_849,In_905,In_1391);
xnor U850 (N_850,In_1213,In_1470);
or U851 (N_851,In_56,In_1805);
and U852 (N_852,In_1434,In_149);
and U853 (N_853,In_1680,In_1296);
or U854 (N_854,In_44,In_1799);
xnor U855 (N_855,In_1569,In_1336);
and U856 (N_856,In_1754,In_119);
nor U857 (N_857,In_1924,In_1398);
or U858 (N_858,In_744,In_1303);
nor U859 (N_859,In_502,In_1030);
and U860 (N_860,In_1747,In_994);
xnor U861 (N_861,In_424,In_855);
and U862 (N_862,In_1814,In_728);
nand U863 (N_863,In_734,In_1394);
or U864 (N_864,In_951,In_1462);
nor U865 (N_865,In_743,In_671);
nor U866 (N_866,In_1407,In_1014);
or U867 (N_867,In_1615,In_1683);
nor U868 (N_868,In_587,In_1060);
nor U869 (N_869,In_163,In_444);
nor U870 (N_870,In_1848,In_155);
nor U871 (N_871,In_1829,In_1714);
nor U872 (N_872,In_1998,In_1925);
and U873 (N_873,In_630,In_172);
nor U874 (N_874,In_1810,In_918);
or U875 (N_875,In_947,In_1678);
nor U876 (N_876,In_1248,In_1960);
xor U877 (N_877,In_924,In_1606);
xnor U878 (N_878,In_1552,In_1153);
xnor U879 (N_879,In_868,In_903);
nand U880 (N_880,In_1220,In_501);
xor U881 (N_881,In_607,In_513);
nand U882 (N_882,In_623,In_134);
or U883 (N_883,In_311,In_1565);
nand U884 (N_884,In_276,In_658);
or U885 (N_885,In_475,In_1389);
xor U886 (N_886,In_1,In_2);
xor U887 (N_887,In_950,In_1449);
and U888 (N_888,In_28,In_1573);
nand U889 (N_889,In_1146,In_1597);
or U890 (N_890,In_848,In_560);
and U891 (N_891,In_0,In_656);
nor U892 (N_892,In_811,In_19);
xnor U893 (N_893,In_203,In_1692);
and U894 (N_894,In_1482,In_48);
or U895 (N_895,In_326,In_1306);
nand U896 (N_896,In_782,In_675);
and U897 (N_897,In_1673,In_1857);
xor U898 (N_898,In_327,In_218);
xnor U899 (N_899,In_189,In_1689);
and U900 (N_900,In_974,In_435);
nand U901 (N_901,In_965,In_1707);
or U902 (N_902,In_1579,In_762);
or U903 (N_903,In_1794,In_1620);
nor U904 (N_904,In_293,In_588);
or U905 (N_905,In_1477,In_1752);
xnor U906 (N_906,In_197,In_714);
and U907 (N_907,In_1542,In_328);
and U908 (N_908,In_1659,In_1653);
nor U909 (N_909,In_1915,In_1612);
and U910 (N_910,In_1671,In_1646);
and U911 (N_911,In_1102,In_679);
or U912 (N_912,In_1443,In_1757);
xnor U913 (N_913,In_1063,In_1160);
or U914 (N_914,In_1974,In_573);
and U915 (N_915,In_1549,In_1850);
and U916 (N_916,In_1123,In_1399);
and U917 (N_917,In_1132,In_1563);
xor U918 (N_918,In_494,In_703);
nor U919 (N_919,In_1734,In_735);
nand U920 (N_920,In_225,In_786);
xor U921 (N_921,In_10,In_1229);
xor U922 (N_922,In_204,In_1668);
and U923 (N_923,In_1944,In_482);
and U924 (N_924,In_1321,In_1231);
xor U925 (N_925,In_639,In_118);
or U926 (N_926,In_303,In_367);
and U927 (N_927,In_1005,In_1150);
and U928 (N_928,In_838,In_1865);
and U929 (N_929,In_1820,In_863);
nand U930 (N_930,In_1755,In_1047);
nand U931 (N_931,In_1261,In_1155);
nand U932 (N_932,In_1157,In_566);
xor U933 (N_933,In_1325,In_65);
and U934 (N_934,In_50,In_1917);
or U935 (N_935,In_1385,In_26);
and U936 (N_936,In_816,In_920);
or U937 (N_937,In_1134,In_668);
nor U938 (N_938,In_1706,In_390);
and U939 (N_939,In_1770,In_620);
or U940 (N_940,In_1828,In_532);
xor U941 (N_941,In_1516,In_843);
nor U942 (N_942,In_794,In_1547);
and U943 (N_943,In_1077,In_1775);
xnor U944 (N_944,In_334,In_102);
xnor U945 (N_945,In_147,In_901);
nor U946 (N_946,In_1269,In_239);
nand U947 (N_947,In_687,In_1866);
and U948 (N_948,In_84,In_678);
or U949 (N_949,In_1608,In_801);
xnor U950 (N_950,In_846,In_541);
xor U951 (N_951,In_1179,In_571);
nor U952 (N_952,In_1080,In_523);
nand U953 (N_953,In_884,In_1934);
or U954 (N_954,In_1148,In_295);
nand U955 (N_955,In_819,In_1097);
xor U956 (N_956,In_343,In_1171);
or U957 (N_957,In_662,In_693);
nand U958 (N_958,In_308,In_68);
xor U959 (N_959,In_1050,In_1488);
or U960 (N_960,In_1165,In_1777);
nand U961 (N_961,In_1910,In_1392);
xnor U962 (N_962,In_1318,In_209);
or U963 (N_963,In_437,In_1401);
and U964 (N_964,In_1083,In_601);
nand U965 (N_965,In_1536,In_954);
nand U966 (N_966,In_1926,In_338);
and U967 (N_967,In_281,In_1785);
xnor U968 (N_968,In_1930,In_910);
nand U969 (N_969,In_632,In_1135);
xor U970 (N_970,In_39,In_62);
xor U971 (N_971,In_653,In_822);
xor U972 (N_972,In_554,In_1937);
or U973 (N_973,In_1466,In_1459);
nand U974 (N_974,In_1744,In_726);
and U975 (N_975,In_1598,In_1028);
or U976 (N_976,In_1344,In_1708);
or U977 (N_977,In_107,In_1803);
xor U978 (N_978,In_274,In_1051);
nor U979 (N_979,In_983,In_528);
or U980 (N_980,In_815,In_379);
or U981 (N_981,In_1533,In_1701);
xor U982 (N_982,In_1648,In_66);
and U983 (N_983,In_582,In_1314);
and U984 (N_984,In_604,In_722);
and U985 (N_985,In_1170,In_202);
and U986 (N_986,In_1712,In_383);
xor U987 (N_987,In_644,In_1630);
nor U988 (N_988,In_932,In_1995);
xnor U989 (N_989,In_1497,In_1772);
nand U990 (N_990,In_1911,In_1619);
or U991 (N_991,In_570,In_120);
xnor U992 (N_992,In_540,In_594);
nand U993 (N_993,In_883,In_455);
and U994 (N_994,In_1214,In_1996);
and U995 (N_995,In_1791,In_861);
and U996 (N_996,In_1667,In_1571);
nand U997 (N_997,In_1845,In_1089);
xor U998 (N_998,In_1507,In_1614);
nand U999 (N_999,In_1666,In_1601);
xnor U1000 (N_1000,N_113,N_820);
and U1001 (N_1001,N_525,N_748);
or U1002 (N_1002,N_838,N_666);
or U1003 (N_1003,N_213,N_429);
xnor U1004 (N_1004,N_544,N_346);
nand U1005 (N_1005,N_32,N_50);
nand U1006 (N_1006,N_702,N_356);
xnor U1007 (N_1007,N_371,N_98);
or U1008 (N_1008,N_347,N_238);
or U1009 (N_1009,N_680,N_788);
xnor U1010 (N_1010,N_104,N_499);
or U1011 (N_1011,N_184,N_248);
nand U1012 (N_1012,N_275,N_16);
xor U1013 (N_1013,N_158,N_786);
nor U1014 (N_1014,N_99,N_504);
nor U1015 (N_1015,N_65,N_168);
or U1016 (N_1016,N_861,N_954);
xnor U1017 (N_1017,N_672,N_412);
or U1018 (N_1018,N_668,N_757);
nor U1019 (N_1019,N_388,N_982);
xnor U1020 (N_1020,N_671,N_214);
and U1021 (N_1021,N_594,N_790);
nor U1022 (N_1022,N_239,N_320);
nand U1023 (N_1023,N_687,N_315);
or U1024 (N_1024,N_586,N_561);
and U1025 (N_1025,N_761,N_90);
xnor U1026 (N_1026,N_628,N_768);
and U1027 (N_1027,N_906,N_457);
nand U1028 (N_1028,N_686,N_23);
nor U1029 (N_1029,N_463,N_829);
xor U1030 (N_1030,N_870,N_636);
nor U1031 (N_1031,N_6,N_278);
and U1032 (N_1032,N_963,N_295);
and U1033 (N_1033,N_314,N_709);
xnor U1034 (N_1034,N_461,N_94);
nor U1035 (N_1035,N_190,N_133);
nor U1036 (N_1036,N_331,N_989);
and U1037 (N_1037,N_580,N_652);
and U1038 (N_1038,N_428,N_690);
nand U1039 (N_1039,N_81,N_382);
xor U1040 (N_1040,N_251,N_336);
nor U1041 (N_1041,N_727,N_9);
nand U1042 (N_1042,N_682,N_816);
nor U1043 (N_1043,N_125,N_302);
xnor U1044 (N_1044,N_489,N_276);
xnor U1045 (N_1045,N_705,N_283);
xnor U1046 (N_1046,N_340,N_827);
or U1047 (N_1047,N_186,N_900);
xor U1048 (N_1048,N_383,N_480);
or U1049 (N_1049,N_610,N_975);
nand U1050 (N_1050,N_500,N_627);
nor U1051 (N_1051,N_294,N_965);
xor U1052 (N_1052,N_44,N_601);
nor U1053 (N_1053,N_940,N_699);
or U1054 (N_1054,N_154,N_341);
or U1055 (N_1055,N_846,N_159);
or U1056 (N_1056,N_365,N_585);
nor U1057 (N_1057,N_25,N_993);
or U1058 (N_1058,N_110,N_150);
or U1059 (N_1059,N_221,N_928);
nor U1060 (N_1060,N_45,N_389);
nor U1061 (N_1061,N_479,N_532);
nor U1062 (N_1062,N_608,N_641);
nor U1063 (N_1063,N_800,N_13);
and U1064 (N_1064,N_811,N_92);
and U1065 (N_1065,N_376,N_316);
nor U1066 (N_1066,N_903,N_157);
or U1067 (N_1067,N_723,N_166);
nor U1068 (N_1068,N_573,N_644);
nor U1069 (N_1069,N_293,N_149);
xnor U1070 (N_1070,N_64,N_357);
or U1071 (N_1071,N_735,N_42);
or U1072 (N_1072,N_679,N_256);
xnor U1073 (N_1073,N_73,N_187);
xnor U1074 (N_1074,N_574,N_889);
and U1075 (N_1075,N_714,N_136);
xor U1076 (N_1076,N_657,N_804);
xnor U1077 (N_1077,N_102,N_191);
or U1078 (N_1078,N_805,N_235);
and U1079 (N_1079,N_775,N_584);
nor U1080 (N_1080,N_950,N_576);
nor U1081 (N_1081,N_393,N_984);
nand U1082 (N_1082,N_462,N_614);
or U1083 (N_1083,N_516,N_62);
nand U1084 (N_1084,N_153,N_442);
nor U1085 (N_1085,N_128,N_173);
nand U1086 (N_1086,N_917,N_247);
nor U1087 (N_1087,N_324,N_893);
nand U1088 (N_1088,N_630,N_338);
nor U1089 (N_1089,N_744,N_834);
and U1090 (N_1090,N_674,N_351);
nor U1091 (N_1091,N_873,N_152);
xor U1092 (N_1092,N_756,N_179);
or U1093 (N_1093,N_66,N_348);
or U1094 (N_1094,N_39,N_103);
and U1095 (N_1095,N_770,N_255);
nand U1096 (N_1096,N_134,N_922);
or U1097 (N_1097,N_857,N_426);
and U1098 (N_1098,N_273,N_28);
and U1099 (N_1099,N_259,N_598);
or U1100 (N_1100,N_175,N_961);
or U1101 (N_1101,N_30,N_223);
and U1102 (N_1102,N_604,N_986);
or U1103 (N_1103,N_664,N_640);
and U1104 (N_1104,N_212,N_261);
or U1105 (N_1105,N_312,N_352);
nor U1106 (N_1106,N_512,N_677);
xor U1107 (N_1107,N_303,N_228);
xor U1108 (N_1108,N_370,N_354);
xor U1109 (N_1109,N_404,N_334);
or U1110 (N_1110,N_427,N_327);
xnor U1111 (N_1111,N_416,N_249);
and U1112 (N_1112,N_34,N_453);
nand U1113 (N_1113,N_531,N_299);
xor U1114 (N_1114,N_911,N_496);
nand U1115 (N_1115,N_291,N_263);
nand U1116 (N_1116,N_758,N_421);
nand U1117 (N_1117,N_855,N_605);
and U1118 (N_1118,N_515,N_0);
xnor U1119 (N_1119,N_321,N_750);
nor U1120 (N_1120,N_880,N_112);
xor U1121 (N_1121,N_969,N_973);
nor U1122 (N_1122,N_445,N_486);
and U1123 (N_1123,N_326,N_519);
nor U1124 (N_1124,N_852,N_527);
and U1125 (N_1125,N_733,N_556);
or U1126 (N_1126,N_147,N_643);
or U1127 (N_1127,N_985,N_550);
nand U1128 (N_1128,N_725,N_131);
and U1129 (N_1129,N_863,N_968);
or U1130 (N_1130,N_737,N_392);
xnor U1131 (N_1131,N_648,N_449);
nand U1132 (N_1132,N_194,N_970);
nor U1133 (N_1133,N_732,N_447);
or U1134 (N_1134,N_625,N_244);
or U1135 (N_1135,N_420,N_58);
nand U1136 (N_1136,N_520,N_237);
and U1137 (N_1137,N_132,N_289);
nand U1138 (N_1138,N_734,N_759);
xor U1139 (N_1139,N_126,N_423);
and U1140 (N_1140,N_407,N_57);
or U1141 (N_1141,N_285,N_116);
nand U1142 (N_1142,N_27,N_994);
nor U1143 (N_1143,N_831,N_465);
nand U1144 (N_1144,N_201,N_367);
or U1145 (N_1145,N_942,N_266);
nor U1146 (N_1146,N_899,N_562);
and U1147 (N_1147,N_4,N_391);
and U1148 (N_1148,N_332,N_858);
xnor U1149 (N_1149,N_74,N_789);
or U1150 (N_1150,N_882,N_595);
nor U1151 (N_1151,N_907,N_205);
xnor U1152 (N_1152,N_162,N_597);
or U1153 (N_1153,N_936,N_559);
xor U1154 (N_1154,N_120,N_773);
or U1155 (N_1155,N_662,N_949);
nand U1156 (N_1156,N_708,N_844);
nor U1157 (N_1157,N_991,N_660);
nand U1158 (N_1158,N_328,N_656);
and U1159 (N_1159,N_538,N_563);
or U1160 (N_1160,N_377,N_529);
nand U1161 (N_1161,N_359,N_91);
or U1162 (N_1162,N_552,N_53);
nand U1163 (N_1163,N_130,N_779);
and U1164 (N_1164,N_912,N_638);
nand U1165 (N_1165,N_943,N_284);
nor U1166 (N_1166,N_141,N_726);
or U1167 (N_1167,N_305,N_864);
or U1168 (N_1168,N_309,N_919);
nor U1169 (N_1169,N_612,N_93);
xnor U1170 (N_1170,N_955,N_84);
nor U1171 (N_1171,N_771,N_891);
and U1172 (N_1172,N_830,N_952);
nand U1173 (N_1173,N_739,N_483);
and U1174 (N_1174,N_452,N_337);
or U1175 (N_1175,N_402,N_358);
xor U1176 (N_1176,N_566,N_31);
xnor U1177 (N_1177,N_491,N_156);
or U1178 (N_1178,N_344,N_583);
and U1179 (N_1179,N_183,N_661);
nand U1180 (N_1180,N_565,N_403);
nor U1181 (N_1181,N_578,N_304);
or U1182 (N_1182,N_799,N_311);
nor U1183 (N_1183,N_883,N_135);
and U1184 (N_1184,N_557,N_956);
xor U1185 (N_1185,N_410,N_808);
or U1186 (N_1186,N_170,N_951);
nand U1187 (N_1187,N_177,N_458);
and U1188 (N_1188,N_242,N_944);
or U1189 (N_1189,N_432,N_897);
nor U1190 (N_1190,N_397,N_859);
and U1191 (N_1191,N_82,N_67);
nand U1192 (N_1192,N_10,N_945);
xor U1193 (N_1193,N_591,N_405);
and U1194 (N_1194,N_105,N_494);
xnor U1195 (N_1195,N_124,N_560);
xor U1196 (N_1196,N_1,N_510);
xnor U1197 (N_1197,N_369,N_22);
nand U1198 (N_1198,N_169,N_929);
xor U1199 (N_1199,N_232,N_570);
and U1200 (N_1200,N_999,N_543);
nor U1201 (N_1201,N_695,N_260);
nor U1202 (N_1202,N_503,N_54);
or U1203 (N_1203,N_617,N_822);
and U1204 (N_1204,N_470,N_33);
nand U1205 (N_1205,N_413,N_697);
nor U1206 (N_1206,N_379,N_509);
xnor U1207 (N_1207,N_785,N_318);
nor U1208 (N_1208,N_689,N_473);
or U1209 (N_1209,N_513,N_987);
nor U1210 (N_1210,N_51,N_654);
xor U1211 (N_1211,N_508,N_751);
xor U1212 (N_1212,N_143,N_366);
xnor U1213 (N_1213,N_724,N_387);
xor U1214 (N_1214,N_363,N_571);
xor U1215 (N_1215,N_862,N_633);
nand U1216 (N_1216,N_224,N_526);
nand U1217 (N_1217,N_868,N_233);
nand U1218 (N_1218,N_207,N_317);
and U1219 (N_1219,N_530,N_47);
xor U1220 (N_1220,N_924,N_720);
nand U1221 (N_1221,N_46,N_460);
nand U1222 (N_1222,N_83,N_69);
nor U1223 (N_1223,N_869,N_579);
or U1224 (N_1224,N_741,N_920);
nor U1225 (N_1225,N_850,N_884);
nor U1226 (N_1226,N_37,N_754);
and U1227 (N_1227,N_776,N_219);
nand U1228 (N_1228,N_921,N_5);
nand U1229 (N_1229,N_52,N_106);
and U1230 (N_1230,N_20,N_781);
nor U1231 (N_1231,N_406,N_189);
nand U1232 (N_1232,N_262,N_916);
xor U1233 (N_1233,N_564,N_990);
xor U1234 (N_1234,N_145,N_441);
or U1235 (N_1235,N_111,N_966);
nor U1236 (N_1236,N_914,N_678);
or U1237 (N_1237,N_373,N_464);
or U1238 (N_1238,N_721,N_218);
and U1239 (N_1239,N_632,N_964);
xor U1240 (N_1240,N_118,N_268);
xor U1241 (N_1241,N_685,N_146);
nor U1242 (N_1242,N_746,N_437);
or U1243 (N_1243,N_319,N_675);
xnor U1244 (N_1244,N_394,N_216);
nand U1245 (N_1245,N_658,N_514);
or U1246 (N_1246,N_645,N_439);
or U1247 (N_1247,N_443,N_254);
nand U1248 (N_1248,N_127,N_88);
xnor U1249 (N_1249,N_901,N_819);
xnor U1250 (N_1250,N_670,N_468);
nor U1251 (N_1251,N_330,N_345);
and U1252 (N_1252,N_611,N_629);
xnor U1253 (N_1253,N_343,N_896);
nor U1254 (N_1254,N_881,N_114);
or U1255 (N_1255,N_307,N_866);
and U1256 (N_1256,N_738,N_182);
nor U1257 (N_1257,N_703,N_817);
nand U1258 (N_1258,N_313,N_151);
nand U1259 (N_1259,N_941,N_204);
xnor U1260 (N_1260,N_15,N_807);
nor U1261 (N_1261,N_706,N_270);
nand U1262 (N_1262,N_109,N_957);
nand U1263 (N_1263,N_841,N_21);
xnor U1264 (N_1264,N_107,N_925);
xnor U1265 (N_1265,N_684,N_414);
nor U1266 (N_1266,N_487,N_581);
and U1267 (N_1267,N_129,N_634);
xor U1268 (N_1268,N_467,N_41);
nor U1269 (N_1269,N_879,N_996);
or U1270 (N_1270,N_743,N_534);
nor U1271 (N_1271,N_430,N_451);
and U1272 (N_1272,N_782,N_108);
xnor U1273 (N_1273,N_333,N_983);
or U1274 (N_1274,N_471,N_24);
nor U1275 (N_1275,N_440,N_481);
and U1276 (N_1276,N_271,N_306);
nor U1277 (N_1277,N_765,N_590);
xnor U1278 (N_1278,N_663,N_878);
nor U1279 (N_1279,N_607,N_995);
or U1280 (N_1280,N_521,N_203);
nand U1281 (N_1281,N_164,N_444);
nand U1282 (N_1282,N_122,N_615);
and U1283 (N_1283,N_596,N_711);
or U1284 (N_1284,N_935,N_475);
and U1285 (N_1285,N_558,N_300);
nor U1286 (N_1286,N_806,N_577);
xnor U1287 (N_1287,N_142,N_138);
xor U1288 (N_1288,N_78,N_613);
and U1289 (N_1289,N_635,N_399);
and U1290 (N_1290,N_553,N_694);
or U1291 (N_1291,N_567,N_849);
nor U1292 (N_1292,N_814,N_745);
xor U1293 (N_1293,N_826,N_419);
nor U1294 (N_1294,N_185,N_325);
nand U1295 (N_1295,N_704,N_226);
nand U1296 (N_1296,N_476,N_502);
nand U1297 (N_1297,N_292,N_227);
nand U1298 (N_1298,N_368,N_140);
xor U1299 (N_1299,N_265,N_192);
or U1300 (N_1300,N_624,N_528);
nor U1301 (N_1301,N_701,N_398);
nand U1302 (N_1302,N_209,N_76);
and U1303 (N_1303,N_243,N_540);
nand U1304 (N_1304,N_2,N_524);
nor U1305 (N_1305,N_812,N_623);
nor U1306 (N_1306,N_839,N_865);
or U1307 (N_1307,N_609,N_976);
xnor U1308 (N_1308,N_715,N_602);
and U1309 (N_1309,N_616,N_930);
nor U1310 (N_1310,N_485,N_698);
xnor U1311 (N_1311,N_281,N_70);
and U1312 (N_1312,N_828,N_448);
nor U1313 (N_1313,N_482,N_395);
and U1314 (N_1314,N_948,N_144);
xnor U1315 (N_1315,N_717,N_823);
xor U1316 (N_1316,N_886,N_848);
nor U1317 (N_1317,N_937,N_980);
nor U1318 (N_1318,N_339,N_653);
and U1319 (N_1319,N_946,N_620);
nor U1320 (N_1320,N_199,N_409);
xnor U1321 (N_1321,N_148,N_301);
and U1322 (N_1322,N_766,N_683);
and U1323 (N_1323,N_161,N_639);
nor U1324 (N_1324,N_760,N_696);
nand U1325 (N_1325,N_72,N_466);
xor U1326 (N_1326,N_77,N_755);
nor U1327 (N_1327,N_163,N_700);
or U1328 (N_1328,N_75,N_18);
xor U1329 (N_1329,N_506,N_763);
xor U1330 (N_1330,N_287,N_234);
nand U1331 (N_1331,N_469,N_49);
or U1332 (N_1332,N_335,N_840);
nor U1333 (N_1333,N_938,N_80);
nand U1334 (N_1334,N_282,N_19);
nand U1335 (N_1335,N_931,N_493);
or U1336 (N_1336,N_752,N_296);
nand U1337 (N_1337,N_240,N_14);
nor U1338 (N_1338,N_913,N_905);
or U1339 (N_1339,N_417,N_362);
or U1340 (N_1340,N_193,N_997);
or U1341 (N_1341,N_48,N_888);
and U1342 (N_1342,N_606,N_290);
nor U1343 (N_1343,N_272,N_511);
and U1344 (N_1344,N_600,N_646);
nand U1345 (N_1345,N_856,N_542);
xnor U1346 (N_1346,N_229,N_424);
and U1347 (N_1347,N_323,N_974);
and U1348 (N_1348,N_8,N_547);
nor U1349 (N_1349,N_908,N_934);
or U1350 (N_1350,N_422,N_716);
nand U1351 (N_1351,N_250,N_972);
or U1352 (N_1352,N_375,N_736);
nand U1353 (N_1353,N_780,N_119);
or U1354 (N_1354,N_978,N_211);
xnor U1355 (N_1355,N_796,N_762);
xnor U1356 (N_1356,N_792,N_548);
or U1357 (N_1357,N_971,N_117);
and U1358 (N_1358,N_435,N_926);
nand U1359 (N_1359,N_286,N_877);
nor U1360 (N_1360,N_722,N_691);
nand U1361 (N_1361,N_433,N_386);
nor U1362 (N_1362,N_208,N_478);
or U1363 (N_1363,N_11,N_507);
or U1364 (N_1364,N_599,N_933);
and U1365 (N_1365,N_274,N_361);
or U1366 (N_1366,N_210,N_3);
nand U1367 (N_1367,N_650,N_349);
or U1368 (N_1368,N_719,N_536);
xor U1369 (N_1369,N_55,N_867);
nor U1370 (N_1370,N_667,N_947);
or U1371 (N_1371,N_876,N_411);
xor U1372 (N_1372,N_582,N_29);
and U1373 (N_1373,N_895,N_139);
xnor U1374 (N_1374,N_195,N_230);
nor U1375 (N_1375,N_35,N_655);
and U1376 (N_1376,N_518,N_533);
xnor U1377 (N_1377,N_554,N_818);
and U1378 (N_1378,N_692,N_206);
or U1379 (N_1379,N_390,N_38);
or U1380 (N_1380,N_434,N_198);
or U1381 (N_1381,N_245,N_631);
nand U1382 (N_1382,N_915,N_225);
nand U1383 (N_1383,N_791,N_767);
nor U1384 (N_1384,N_693,N_798);
xor U1385 (N_1385,N_79,N_787);
and U1386 (N_1386,N_68,N_188);
xnor U1387 (N_1387,N_215,N_847);
and U1388 (N_1388,N_810,N_355);
nand U1389 (N_1389,N_885,N_60);
nor U1390 (N_1390,N_647,N_492);
nor U1391 (N_1391,N_904,N_537);
and U1392 (N_1392,N_196,N_86);
nand U1393 (N_1393,N_269,N_825);
or U1394 (N_1394,N_374,N_833);
nand U1395 (N_1395,N_97,N_96);
nor U1396 (N_1396,N_100,N_505);
nor U1397 (N_1397,N_875,N_436);
nand U1398 (N_1398,N_551,N_87);
and U1399 (N_1399,N_472,N_85);
xnor U1400 (N_1400,N_795,N_575);
nand U1401 (N_1401,N_497,N_438);
or U1402 (N_1402,N_802,N_501);
nand U1403 (N_1403,N_932,N_821);
and U1404 (N_1404,N_592,N_774);
nand U1405 (N_1405,N_56,N_673);
or U1406 (N_1406,N_713,N_960);
nor U1407 (N_1407,N_63,N_953);
xor U1408 (N_1408,N_517,N_431);
and U1409 (N_1409,N_651,N_707);
nor U1410 (N_1410,N_572,N_872);
xnor U1411 (N_1411,N_981,N_626);
xnor U1412 (N_1412,N_353,N_665);
xor U1413 (N_1413,N_258,N_910);
and U1414 (N_1414,N_165,N_381);
or U1415 (N_1415,N_769,N_43);
nand U1416 (N_1416,N_252,N_718);
and U1417 (N_1417,N_7,N_308);
or U1418 (N_1418,N_927,N_962);
xor U1419 (N_1419,N_803,N_740);
and U1420 (N_1420,N_959,N_277);
nor U1421 (N_1421,N_498,N_488);
nand U1422 (N_1422,N_360,N_197);
or U1423 (N_1423,N_396,N_593);
or U1424 (N_1424,N_618,N_415);
xnor U1425 (N_1425,N_523,N_257);
nor U1426 (N_1426,N_778,N_400);
and U1427 (N_1427,N_642,N_589);
nor U1428 (N_1428,N_832,N_621);
and U1429 (N_1429,N_446,N_898);
or U1430 (N_1430,N_992,N_180);
nor U1431 (N_1431,N_851,N_813);
nand U1432 (N_1432,N_710,N_178);
and U1433 (N_1433,N_342,N_793);
nand U1434 (N_1434,N_967,N_742);
xnor U1435 (N_1435,N_115,N_380);
or U1436 (N_1436,N_310,N_772);
nor U1437 (N_1437,N_619,N_918);
nand U1438 (N_1438,N_137,N_425);
xor U1439 (N_1439,N_659,N_874);
and U1440 (N_1440,N_902,N_71);
xor U1441 (N_1441,N_815,N_753);
xor U1442 (N_1442,N_669,N_123);
xor U1443 (N_1443,N_603,N_322);
nand U1444 (N_1444,N_892,N_459);
or U1445 (N_1445,N_329,N_794);
xor U1446 (N_1446,N_174,N_731);
xor U1447 (N_1447,N_854,N_454);
xnor U1448 (N_1448,N_40,N_728);
nor U1449 (N_1449,N_522,N_783);
and U1450 (N_1450,N_181,N_784);
nand U1451 (N_1451,N_890,N_236);
xor U1452 (N_1452,N_555,N_279);
xor U1453 (N_1453,N_729,N_484);
nand U1454 (N_1454,N_241,N_809);
nor U1455 (N_1455,N_246,N_121);
xor U1456 (N_1456,N_569,N_297);
nand U1457 (N_1457,N_998,N_894);
nand U1458 (N_1458,N_280,N_101);
or U1459 (N_1459,N_842,N_988);
xor U1460 (N_1460,N_456,N_546);
or U1461 (N_1461,N_26,N_909);
and U1462 (N_1462,N_887,N_171);
nor U1463 (N_1463,N_549,N_977);
or U1464 (N_1464,N_220,N_845);
xor U1465 (N_1465,N_495,N_939);
xnor U1466 (N_1466,N_36,N_797);
xor U1467 (N_1467,N_622,N_545);
xor U1468 (N_1468,N_17,N_860);
or U1469 (N_1469,N_95,N_12);
xnor U1470 (N_1470,N_167,N_637);
nor U1471 (N_1471,N_764,N_372);
nand U1472 (N_1472,N_455,N_288);
nor U1473 (N_1473,N_539,N_89);
nor U1474 (N_1474,N_253,N_231);
and U1475 (N_1475,N_568,N_408);
xnor U1476 (N_1476,N_837,N_688);
and U1477 (N_1477,N_217,N_474);
xor U1478 (N_1478,N_202,N_824);
nor U1479 (N_1479,N_749,N_384);
xnor U1480 (N_1480,N_801,N_172);
xnor U1481 (N_1481,N_871,N_401);
and U1482 (N_1482,N_364,N_350);
and U1483 (N_1483,N_681,N_843);
or U1484 (N_1484,N_264,N_418);
and U1485 (N_1485,N_853,N_267);
nor U1486 (N_1486,N_835,N_61);
nand U1487 (N_1487,N_59,N_712);
or U1488 (N_1488,N_676,N_155);
nand U1489 (N_1489,N_649,N_298);
and U1490 (N_1490,N_730,N_958);
nor U1491 (N_1491,N_777,N_222);
nand U1492 (N_1492,N_477,N_979);
nand U1493 (N_1493,N_836,N_923);
or U1494 (N_1494,N_176,N_588);
nand U1495 (N_1495,N_200,N_490);
or U1496 (N_1496,N_747,N_450);
xor U1497 (N_1497,N_587,N_541);
nand U1498 (N_1498,N_160,N_535);
nor U1499 (N_1499,N_378,N_385);
or U1500 (N_1500,N_301,N_425);
or U1501 (N_1501,N_121,N_767);
xnor U1502 (N_1502,N_248,N_347);
nor U1503 (N_1503,N_71,N_189);
nand U1504 (N_1504,N_10,N_263);
xnor U1505 (N_1505,N_50,N_493);
nor U1506 (N_1506,N_422,N_744);
xor U1507 (N_1507,N_188,N_916);
nand U1508 (N_1508,N_255,N_175);
and U1509 (N_1509,N_99,N_701);
or U1510 (N_1510,N_118,N_445);
nor U1511 (N_1511,N_694,N_919);
nand U1512 (N_1512,N_930,N_857);
nand U1513 (N_1513,N_727,N_827);
and U1514 (N_1514,N_470,N_62);
nor U1515 (N_1515,N_831,N_171);
nor U1516 (N_1516,N_970,N_349);
nand U1517 (N_1517,N_657,N_907);
xnor U1518 (N_1518,N_709,N_12);
and U1519 (N_1519,N_985,N_264);
nor U1520 (N_1520,N_28,N_433);
nor U1521 (N_1521,N_241,N_639);
nand U1522 (N_1522,N_484,N_28);
nor U1523 (N_1523,N_435,N_292);
nand U1524 (N_1524,N_946,N_270);
xor U1525 (N_1525,N_137,N_34);
or U1526 (N_1526,N_980,N_946);
xor U1527 (N_1527,N_155,N_527);
xnor U1528 (N_1528,N_82,N_421);
nand U1529 (N_1529,N_222,N_312);
or U1530 (N_1530,N_346,N_560);
nand U1531 (N_1531,N_491,N_239);
nand U1532 (N_1532,N_896,N_127);
nand U1533 (N_1533,N_34,N_562);
or U1534 (N_1534,N_67,N_394);
or U1535 (N_1535,N_908,N_368);
nor U1536 (N_1536,N_342,N_143);
or U1537 (N_1537,N_589,N_559);
or U1538 (N_1538,N_912,N_8);
xor U1539 (N_1539,N_435,N_68);
xnor U1540 (N_1540,N_112,N_558);
xnor U1541 (N_1541,N_722,N_438);
nand U1542 (N_1542,N_853,N_249);
nand U1543 (N_1543,N_975,N_250);
and U1544 (N_1544,N_257,N_737);
nand U1545 (N_1545,N_702,N_120);
xnor U1546 (N_1546,N_154,N_357);
xor U1547 (N_1547,N_653,N_5);
xnor U1548 (N_1548,N_377,N_355);
and U1549 (N_1549,N_42,N_461);
nor U1550 (N_1550,N_988,N_501);
nor U1551 (N_1551,N_688,N_609);
xnor U1552 (N_1552,N_175,N_372);
and U1553 (N_1553,N_710,N_498);
nand U1554 (N_1554,N_712,N_937);
xor U1555 (N_1555,N_194,N_125);
or U1556 (N_1556,N_891,N_690);
nor U1557 (N_1557,N_486,N_88);
and U1558 (N_1558,N_568,N_716);
nor U1559 (N_1559,N_17,N_222);
xnor U1560 (N_1560,N_374,N_184);
and U1561 (N_1561,N_413,N_979);
and U1562 (N_1562,N_726,N_657);
and U1563 (N_1563,N_599,N_928);
nor U1564 (N_1564,N_112,N_487);
and U1565 (N_1565,N_400,N_238);
and U1566 (N_1566,N_647,N_905);
nor U1567 (N_1567,N_592,N_15);
nand U1568 (N_1568,N_420,N_429);
or U1569 (N_1569,N_980,N_384);
and U1570 (N_1570,N_781,N_308);
and U1571 (N_1571,N_650,N_284);
nor U1572 (N_1572,N_157,N_236);
nand U1573 (N_1573,N_246,N_73);
or U1574 (N_1574,N_382,N_417);
xnor U1575 (N_1575,N_276,N_512);
nor U1576 (N_1576,N_262,N_841);
nand U1577 (N_1577,N_983,N_252);
nor U1578 (N_1578,N_608,N_540);
nand U1579 (N_1579,N_692,N_315);
nor U1580 (N_1580,N_130,N_800);
or U1581 (N_1581,N_634,N_317);
xnor U1582 (N_1582,N_544,N_56);
xnor U1583 (N_1583,N_663,N_27);
and U1584 (N_1584,N_544,N_111);
nand U1585 (N_1585,N_472,N_809);
nand U1586 (N_1586,N_908,N_199);
xnor U1587 (N_1587,N_792,N_615);
or U1588 (N_1588,N_825,N_450);
or U1589 (N_1589,N_616,N_193);
xor U1590 (N_1590,N_396,N_583);
or U1591 (N_1591,N_952,N_715);
or U1592 (N_1592,N_963,N_348);
and U1593 (N_1593,N_643,N_122);
and U1594 (N_1594,N_959,N_778);
nand U1595 (N_1595,N_549,N_426);
and U1596 (N_1596,N_225,N_311);
nor U1597 (N_1597,N_286,N_939);
or U1598 (N_1598,N_815,N_524);
nand U1599 (N_1599,N_754,N_294);
or U1600 (N_1600,N_561,N_981);
and U1601 (N_1601,N_917,N_565);
nor U1602 (N_1602,N_290,N_733);
xnor U1603 (N_1603,N_218,N_597);
or U1604 (N_1604,N_791,N_128);
xnor U1605 (N_1605,N_406,N_2);
and U1606 (N_1606,N_826,N_671);
nor U1607 (N_1607,N_434,N_714);
and U1608 (N_1608,N_781,N_596);
xor U1609 (N_1609,N_700,N_861);
nand U1610 (N_1610,N_806,N_221);
nand U1611 (N_1611,N_259,N_813);
and U1612 (N_1612,N_178,N_799);
nand U1613 (N_1613,N_368,N_978);
or U1614 (N_1614,N_494,N_833);
nand U1615 (N_1615,N_146,N_364);
nor U1616 (N_1616,N_482,N_398);
nor U1617 (N_1617,N_576,N_361);
nor U1618 (N_1618,N_832,N_234);
xor U1619 (N_1619,N_34,N_350);
nor U1620 (N_1620,N_730,N_935);
nand U1621 (N_1621,N_748,N_254);
nand U1622 (N_1622,N_69,N_286);
and U1623 (N_1623,N_190,N_956);
or U1624 (N_1624,N_296,N_563);
nand U1625 (N_1625,N_752,N_273);
nor U1626 (N_1626,N_607,N_414);
or U1627 (N_1627,N_919,N_337);
nand U1628 (N_1628,N_4,N_395);
and U1629 (N_1629,N_581,N_807);
and U1630 (N_1630,N_918,N_747);
or U1631 (N_1631,N_860,N_453);
xor U1632 (N_1632,N_27,N_431);
xnor U1633 (N_1633,N_576,N_434);
nor U1634 (N_1634,N_528,N_917);
or U1635 (N_1635,N_538,N_237);
and U1636 (N_1636,N_141,N_246);
and U1637 (N_1637,N_837,N_749);
or U1638 (N_1638,N_499,N_372);
and U1639 (N_1639,N_705,N_609);
and U1640 (N_1640,N_812,N_449);
or U1641 (N_1641,N_156,N_279);
and U1642 (N_1642,N_206,N_209);
nor U1643 (N_1643,N_228,N_541);
nor U1644 (N_1644,N_647,N_601);
nand U1645 (N_1645,N_521,N_770);
xnor U1646 (N_1646,N_51,N_469);
nor U1647 (N_1647,N_208,N_299);
and U1648 (N_1648,N_489,N_969);
nor U1649 (N_1649,N_75,N_543);
or U1650 (N_1650,N_478,N_894);
and U1651 (N_1651,N_431,N_800);
nand U1652 (N_1652,N_553,N_793);
nor U1653 (N_1653,N_476,N_175);
nor U1654 (N_1654,N_804,N_938);
and U1655 (N_1655,N_693,N_591);
nor U1656 (N_1656,N_480,N_299);
nor U1657 (N_1657,N_895,N_681);
or U1658 (N_1658,N_978,N_127);
or U1659 (N_1659,N_594,N_528);
nand U1660 (N_1660,N_853,N_516);
xnor U1661 (N_1661,N_164,N_930);
and U1662 (N_1662,N_826,N_546);
xnor U1663 (N_1663,N_458,N_358);
and U1664 (N_1664,N_875,N_17);
xnor U1665 (N_1665,N_824,N_19);
nand U1666 (N_1666,N_25,N_300);
or U1667 (N_1667,N_644,N_921);
nand U1668 (N_1668,N_699,N_899);
nor U1669 (N_1669,N_60,N_721);
or U1670 (N_1670,N_784,N_883);
or U1671 (N_1671,N_304,N_150);
or U1672 (N_1672,N_331,N_533);
or U1673 (N_1673,N_527,N_583);
xnor U1674 (N_1674,N_438,N_738);
and U1675 (N_1675,N_263,N_665);
nor U1676 (N_1676,N_270,N_668);
nand U1677 (N_1677,N_872,N_442);
and U1678 (N_1678,N_279,N_439);
or U1679 (N_1679,N_797,N_183);
nand U1680 (N_1680,N_143,N_13);
and U1681 (N_1681,N_320,N_163);
nor U1682 (N_1682,N_689,N_485);
xor U1683 (N_1683,N_813,N_532);
xor U1684 (N_1684,N_373,N_806);
xnor U1685 (N_1685,N_80,N_409);
or U1686 (N_1686,N_833,N_161);
xnor U1687 (N_1687,N_611,N_125);
nand U1688 (N_1688,N_665,N_750);
nand U1689 (N_1689,N_95,N_974);
or U1690 (N_1690,N_358,N_52);
and U1691 (N_1691,N_183,N_52);
and U1692 (N_1692,N_545,N_6);
or U1693 (N_1693,N_551,N_569);
nand U1694 (N_1694,N_54,N_497);
and U1695 (N_1695,N_352,N_260);
or U1696 (N_1696,N_126,N_221);
or U1697 (N_1697,N_864,N_775);
and U1698 (N_1698,N_753,N_539);
nand U1699 (N_1699,N_795,N_711);
and U1700 (N_1700,N_614,N_495);
nor U1701 (N_1701,N_693,N_836);
nand U1702 (N_1702,N_213,N_682);
nand U1703 (N_1703,N_686,N_218);
and U1704 (N_1704,N_146,N_297);
xnor U1705 (N_1705,N_163,N_809);
xnor U1706 (N_1706,N_811,N_483);
xor U1707 (N_1707,N_281,N_541);
xor U1708 (N_1708,N_692,N_955);
nor U1709 (N_1709,N_439,N_483);
nand U1710 (N_1710,N_578,N_536);
and U1711 (N_1711,N_683,N_123);
nor U1712 (N_1712,N_939,N_911);
and U1713 (N_1713,N_116,N_314);
nor U1714 (N_1714,N_424,N_597);
nor U1715 (N_1715,N_760,N_396);
or U1716 (N_1716,N_258,N_899);
nor U1717 (N_1717,N_810,N_15);
or U1718 (N_1718,N_585,N_605);
and U1719 (N_1719,N_174,N_234);
nor U1720 (N_1720,N_366,N_401);
nand U1721 (N_1721,N_38,N_714);
nand U1722 (N_1722,N_921,N_793);
nor U1723 (N_1723,N_163,N_526);
xnor U1724 (N_1724,N_961,N_534);
nand U1725 (N_1725,N_273,N_632);
or U1726 (N_1726,N_658,N_711);
or U1727 (N_1727,N_358,N_55);
xnor U1728 (N_1728,N_373,N_830);
nand U1729 (N_1729,N_660,N_983);
nor U1730 (N_1730,N_287,N_793);
and U1731 (N_1731,N_417,N_441);
xnor U1732 (N_1732,N_40,N_805);
and U1733 (N_1733,N_666,N_474);
and U1734 (N_1734,N_148,N_831);
and U1735 (N_1735,N_175,N_998);
nor U1736 (N_1736,N_504,N_5);
and U1737 (N_1737,N_929,N_475);
nor U1738 (N_1738,N_275,N_18);
xor U1739 (N_1739,N_198,N_271);
nor U1740 (N_1740,N_320,N_44);
nand U1741 (N_1741,N_892,N_20);
nand U1742 (N_1742,N_173,N_295);
or U1743 (N_1743,N_644,N_17);
and U1744 (N_1744,N_664,N_160);
nor U1745 (N_1745,N_310,N_563);
xnor U1746 (N_1746,N_713,N_256);
xnor U1747 (N_1747,N_404,N_401);
xnor U1748 (N_1748,N_287,N_341);
or U1749 (N_1749,N_506,N_369);
nand U1750 (N_1750,N_220,N_738);
xnor U1751 (N_1751,N_807,N_75);
xor U1752 (N_1752,N_246,N_467);
and U1753 (N_1753,N_685,N_19);
xnor U1754 (N_1754,N_617,N_720);
nand U1755 (N_1755,N_240,N_155);
nand U1756 (N_1756,N_916,N_851);
and U1757 (N_1757,N_218,N_858);
nor U1758 (N_1758,N_418,N_464);
xnor U1759 (N_1759,N_664,N_691);
nand U1760 (N_1760,N_722,N_588);
or U1761 (N_1761,N_232,N_68);
or U1762 (N_1762,N_873,N_14);
xnor U1763 (N_1763,N_486,N_602);
nand U1764 (N_1764,N_105,N_6);
xor U1765 (N_1765,N_471,N_494);
xor U1766 (N_1766,N_818,N_74);
nand U1767 (N_1767,N_439,N_446);
xor U1768 (N_1768,N_416,N_334);
or U1769 (N_1769,N_888,N_45);
and U1770 (N_1770,N_325,N_40);
and U1771 (N_1771,N_973,N_502);
or U1772 (N_1772,N_773,N_696);
xor U1773 (N_1773,N_652,N_559);
xor U1774 (N_1774,N_253,N_96);
nand U1775 (N_1775,N_837,N_803);
nor U1776 (N_1776,N_910,N_792);
xor U1777 (N_1777,N_261,N_173);
nor U1778 (N_1778,N_228,N_784);
or U1779 (N_1779,N_525,N_996);
nand U1780 (N_1780,N_763,N_688);
xnor U1781 (N_1781,N_285,N_897);
nand U1782 (N_1782,N_597,N_335);
nor U1783 (N_1783,N_183,N_492);
nor U1784 (N_1784,N_158,N_640);
nand U1785 (N_1785,N_305,N_467);
or U1786 (N_1786,N_515,N_89);
and U1787 (N_1787,N_873,N_535);
or U1788 (N_1788,N_738,N_509);
xor U1789 (N_1789,N_481,N_246);
nor U1790 (N_1790,N_716,N_695);
and U1791 (N_1791,N_465,N_217);
nand U1792 (N_1792,N_184,N_931);
xnor U1793 (N_1793,N_621,N_26);
xor U1794 (N_1794,N_258,N_810);
xor U1795 (N_1795,N_412,N_341);
xor U1796 (N_1796,N_100,N_750);
nand U1797 (N_1797,N_450,N_417);
nor U1798 (N_1798,N_707,N_73);
or U1799 (N_1799,N_439,N_889);
nor U1800 (N_1800,N_276,N_294);
nor U1801 (N_1801,N_349,N_254);
nand U1802 (N_1802,N_648,N_807);
nand U1803 (N_1803,N_305,N_947);
nor U1804 (N_1804,N_665,N_442);
xor U1805 (N_1805,N_683,N_885);
or U1806 (N_1806,N_849,N_249);
nand U1807 (N_1807,N_767,N_607);
nand U1808 (N_1808,N_974,N_467);
or U1809 (N_1809,N_128,N_492);
or U1810 (N_1810,N_319,N_982);
and U1811 (N_1811,N_550,N_794);
xnor U1812 (N_1812,N_491,N_191);
or U1813 (N_1813,N_857,N_144);
nor U1814 (N_1814,N_736,N_317);
nor U1815 (N_1815,N_490,N_793);
xor U1816 (N_1816,N_594,N_974);
nor U1817 (N_1817,N_168,N_347);
and U1818 (N_1818,N_211,N_320);
and U1819 (N_1819,N_563,N_529);
nor U1820 (N_1820,N_68,N_447);
and U1821 (N_1821,N_453,N_948);
or U1822 (N_1822,N_566,N_645);
xor U1823 (N_1823,N_352,N_104);
nor U1824 (N_1824,N_713,N_115);
and U1825 (N_1825,N_924,N_918);
xor U1826 (N_1826,N_522,N_387);
or U1827 (N_1827,N_140,N_383);
and U1828 (N_1828,N_503,N_552);
nor U1829 (N_1829,N_972,N_227);
nor U1830 (N_1830,N_582,N_839);
or U1831 (N_1831,N_33,N_182);
or U1832 (N_1832,N_557,N_407);
or U1833 (N_1833,N_979,N_607);
xor U1834 (N_1834,N_964,N_142);
and U1835 (N_1835,N_397,N_235);
nand U1836 (N_1836,N_303,N_4);
or U1837 (N_1837,N_320,N_541);
xor U1838 (N_1838,N_381,N_987);
xnor U1839 (N_1839,N_827,N_635);
or U1840 (N_1840,N_27,N_259);
nand U1841 (N_1841,N_589,N_986);
and U1842 (N_1842,N_774,N_214);
nand U1843 (N_1843,N_172,N_30);
or U1844 (N_1844,N_698,N_847);
or U1845 (N_1845,N_517,N_338);
nor U1846 (N_1846,N_423,N_233);
nand U1847 (N_1847,N_729,N_996);
and U1848 (N_1848,N_856,N_757);
or U1849 (N_1849,N_845,N_175);
or U1850 (N_1850,N_245,N_36);
nor U1851 (N_1851,N_761,N_387);
nand U1852 (N_1852,N_9,N_446);
or U1853 (N_1853,N_647,N_163);
xor U1854 (N_1854,N_132,N_852);
nand U1855 (N_1855,N_181,N_114);
or U1856 (N_1856,N_467,N_61);
and U1857 (N_1857,N_364,N_566);
nor U1858 (N_1858,N_676,N_315);
nor U1859 (N_1859,N_571,N_358);
xnor U1860 (N_1860,N_517,N_112);
xnor U1861 (N_1861,N_78,N_824);
and U1862 (N_1862,N_463,N_36);
nand U1863 (N_1863,N_499,N_179);
and U1864 (N_1864,N_430,N_182);
and U1865 (N_1865,N_563,N_785);
nand U1866 (N_1866,N_619,N_491);
or U1867 (N_1867,N_796,N_487);
nand U1868 (N_1868,N_819,N_726);
or U1869 (N_1869,N_78,N_686);
and U1870 (N_1870,N_308,N_628);
nor U1871 (N_1871,N_960,N_252);
and U1872 (N_1872,N_611,N_632);
nand U1873 (N_1873,N_187,N_566);
or U1874 (N_1874,N_967,N_646);
nand U1875 (N_1875,N_318,N_238);
nor U1876 (N_1876,N_160,N_95);
nor U1877 (N_1877,N_308,N_530);
nand U1878 (N_1878,N_399,N_484);
xor U1879 (N_1879,N_170,N_302);
nand U1880 (N_1880,N_348,N_704);
or U1881 (N_1881,N_233,N_226);
or U1882 (N_1882,N_355,N_220);
xor U1883 (N_1883,N_277,N_283);
nor U1884 (N_1884,N_776,N_105);
or U1885 (N_1885,N_935,N_397);
and U1886 (N_1886,N_582,N_919);
nor U1887 (N_1887,N_145,N_464);
or U1888 (N_1888,N_834,N_276);
and U1889 (N_1889,N_567,N_600);
or U1890 (N_1890,N_864,N_356);
xor U1891 (N_1891,N_489,N_639);
nand U1892 (N_1892,N_783,N_868);
xnor U1893 (N_1893,N_457,N_297);
nor U1894 (N_1894,N_95,N_94);
nor U1895 (N_1895,N_128,N_986);
nand U1896 (N_1896,N_571,N_487);
and U1897 (N_1897,N_359,N_714);
and U1898 (N_1898,N_457,N_925);
nor U1899 (N_1899,N_843,N_774);
xor U1900 (N_1900,N_518,N_775);
or U1901 (N_1901,N_800,N_195);
or U1902 (N_1902,N_565,N_332);
nand U1903 (N_1903,N_843,N_928);
nor U1904 (N_1904,N_346,N_827);
or U1905 (N_1905,N_29,N_792);
or U1906 (N_1906,N_51,N_733);
nand U1907 (N_1907,N_946,N_320);
and U1908 (N_1908,N_152,N_911);
and U1909 (N_1909,N_433,N_477);
nand U1910 (N_1910,N_980,N_257);
or U1911 (N_1911,N_915,N_82);
and U1912 (N_1912,N_423,N_68);
nor U1913 (N_1913,N_348,N_167);
nand U1914 (N_1914,N_526,N_858);
and U1915 (N_1915,N_65,N_865);
xor U1916 (N_1916,N_335,N_636);
nor U1917 (N_1917,N_118,N_945);
nor U1918 (N_1918,N_776,N_707);
and U1919 (N_1919,N_157,N_196);
nand U1920 (N_1920,N_489,N_523);
or U1921 (N_1921,N_151,N_222);
xnor U1922 (N_1922,N_216,N_864);
nor U1923 (N_1923,N_332,N_910);
xor U1924 (N_1924,N_55,N_5);
and U1925 (N_1925,N_569,N_152);
or U1926 (N_1926,N_413,N_941);
xor U1927 (N_1927,N_574,N_54);
nor U1928 (N_1928,N_328,N_613);
xnor U1929 (N_1929,N_145,N_747);
or U1930 (N_1930,N_910,N_606);
xor U1931 (N_1931,N_474,N_310);
or U1932 (N_1932,N_783,N_778);
nand U1933 (N_1933,N_959,N_594);
or U1934 (N_1934,N_774,N_444);
or U1935 (N_1935,N_236,N_70);
nor U1936 (N_1936,N_373,N_99);
or U1937 (N_1937,N_94,N_135);
and U1938 (N_1938,N_541,N_829);
or U1939 (N_1939,N_157,N_448);
or U1940 (N_1940,N_79,N_53);
and U1941 (N_1941,N_483,N_883);
nand U1942 (N_1942,N_209,N_829);
xor U1943 (N_1943,N_429,N_788);
or U1944 (N_1944,N_706,N_19);
nor U1945 (N_1945,N_321,N_865);
xnor U1946 (N_1946,N_129,N_811);
xnor U1947 (N_1947,N_757,N_972);
or U1948 (N_1948,N_531,N_944);
xor U1949 (N_1949,N_68,N_663);
nor U1950 (N_1950,N_575,N_227);
nor U1951 (N_1951,N_616,N_911);
or U1952 (N_1952,N_644,N_284);
nor U1953 (N_1953,N_150,N_138);
or U1954 (N_1954,N_972,N_511);
and U1955 (N_1955,N_724,N_158);
nand U1956 (N_1956,N_751,N_697);
xor U1957 (N_1957,N_378,N_149);
nor U1958 (N_1958,N_805,N_777);
and U1959 (N_1959,N_251,N_515);
xnor U1960 (N_1960,N_495,N_418);
and U1961 (N_1961,N_22,N_500);
xnor U1962 (N_1962,N_678,N_765);
and U1963 (N_1963,N_210,N_18);
nor U1964 (N_1964,N_89,N_739);
or U1965 (N_1965,N_308,N_387);
or U1966 (N_1966,N_359,N_111);
nand U1967 (N_1967,N_130,N_670);
nand U1968 (N_1968,N_791,N_549);
nand U1969 (N_1969,N_369,N_158);
nor U1970 (N_1970,N_741,N_852);
and U1971 (N_1971,N_76,N_52);
xnor U1972 (N_1972,N_80,N_285);
nor U1973 (N_1973,N_718,N_79);
xor U1974 (N_1974,N_35,N_828);
nor U1975 (N_1975,N_123,N_728);
xnor U1976 (N_1976,N_567,N_869);
and U1977 (N_1977,N_383,N_699);
xnor U1978 (N_1978,N_88,N_567);
or U1979 (N_1979,N_226,N_322);
or U1980 (N_1980,N_686,N_409);
nor U1981 (N_1981,N_43,N_420);
or U1982 (N_1982,N_414,N_314);
nor U1983 (N_1983,N_223,N_725);
nand U1984 (N_1984,N_708,N_800);
nand U1985 (N_1985,N_847,N_822);
xor U1986 (N_1986,N_2,N_888);
nand U1987 (N_1987,N_248,N_58);
nand U1988 (N_1988,N_257,N_767);
nor U1989 (N_1989,N_9,N_64);
nor U1990 (N_1990,N_767,N_483);
and U1991 (N_1991,N_836,N_114);
nand U1992 (N_1992,N_214,N_803);
or U1993 (N_1993,N_667,N_605);
and U1994 (N_1994,N_407,N_434);
and U1995 (N_1995,N_256,N_617);
or U1996 (N_1996,N_843,N_974);
nor U1997 (N_1997,N_715,N_990);
nand U1998 (N_1998,N_939,N_856);
xnor U1999 (N_1999,N_947,N_465);
nor U2000 (N_2000,N_1885,N_1939);
or U2001 (N_2001,N_1180,N_1892);
or U2002 (N_2002,N_1446,N_1737);
xnor U2003 (N_2003,N_1799,N_1267);
or U2004 (N_2004,N_1889,N_1306);
nor U2005 (N_2005,N_1499,N_1917);
nand U2006 (N_2006,N_1545,N_1578);
nand U2007 (N_2007,N_1583,N_1571);
nor U2008 (N_2008,N_1385,N_1626);
nand U2009 (N_2009,N_1605,N_1593);
or U2010 (N_2010,N_1857,N_1462);
or U2011 (N_2011,N_1068,N_1091);
xnor U2012 (N_2012,N_1404,N_1609);
nor U2013 (N_2013,N_1142,N_1680);
nand U2014 (N_2014,N_1137,N_1188);
nand U2015 (N_2015,N_1454,N_1791);
nand U2016 (N_2016,N_1122,N_1964);
or U2017 (N_2017,N_1480,N_1246);
nor U2018 (N_2018,N_1055,N_1211);
nand U2019 (N_2019,N_1350,N_1401);
and U2020 (N_2020,N_1101,N_1519);
or U2021 (N_2021,N_1093,N_1097);
nor U2022 (N_2022,N_1872,N_1637);
and U2023 (N_2023,N_1636,N_1774);
xor U2024 (N_2024,N_1066,N_1763);
or U2025 (N_2025,N_1397,N_1878);
nor U2026 (N_2026,N_1032,N_1975);
nand U2027 (N_2027,N_1945,N_1342);
xor U2028 (N_2028,N_1380,N_1738);
nor U2029 (N_2029,N_1849,N_1143);
and U2030 (N_2030,N_1445,N_1275);
nand U2031 (N_2031,N_1860,N_1662);
nor U2032 (N_2032,N_1356,N_1094);
nand U2033 (N_2033,N_1811,N_1440);
nand U2034 (N_2034,N_1187,N_1253);
nand U2035 (N_2035,N_1704,N_1428);
and U2036 (N_2036,N_1140,N_1089);
or U2037 (N_2037,N_1853,N_1432);
xor U2038 (N_2038,N_1795,N_1357);
xnor U2039 (N_2039,N_1971,N_1630);
and U2040 (N_2040,N_1219,N_1844);
xnor U2041 (N_2041,N_1335,N_1570);
or U2042 (N_2042,N_1057,N_1284);
nand U2043 (N_2043,N_1222,N_1443);
and U2044 (N_2044,N_1415,N_1381);
or U2045 (N_2045,N_1105,N_1114);
nor U2046 (N_2046,N_1410,N_1161);
nand U2047 (N_2047,N_1809,N_1834);
xnor U2048 (N_2048,N_1937,N_1072);
or U2049 (N_2049,N_1554,N_1002);
nor U2050 (N_2050,N_1374,N_1978);
nor U2051 (N_2051,N_1653,N_1847);
nor U2052 (N_2052,N_1264,N_1320);
nand U2053 (N_2053,N_1254,N_1854);
xnor U2054 (N_2054,N_1539,N_1429);
nand U2055 (N_2055,N_1391,N_1619);
or U2056 (N_2056,N_1363,N_1893);
xnor U2057 (N_2057,N_1150,N_1479);
xor U2058 (N_2058,N_1153,N_1448);
and U2059 (N_2059,N_1595,N_1108);
and U2060 (N_2060,N_1149,N_1011);
xor U2061 (N_2061,N_1651,N_1599);
xor U2062 (N_2062,N_1212,N_1762);
and U2063 (N_2063,N_1262,N_1976);
and U2064 (N_2064,N_1168,N_1044);
or U2065 (N_2065,N_1258,N_1884);
nor U2066 (N_2066,N_1079,N_1934);
nand U2067 (N_2067,N_1483,N_1782);
and U2068 (N_2068,N_1426,N_1814);
or U2069 (N_2069,N_1125,N_1841);
xor U2070 (N_2070,N_1204,N_1887);
nor U2071 (N_2071,N_1989,N_1634);
or U2072 (N_2072,N_1458,N_1229);
nor U2073 (N_2073,N_1899,N_1994);
and U2074 (N_2074,N_1319,N_1327);
or U2075 (N_2075,N_1724,N_1046);
or U2076 (N_2076,N_1160,N_1765);
or U2077 (N_2077,N_1580,N_1243);
xnor U2078 (N_2078,N_1240,N_1829);
nand U2079 (N_2079,N_1713,N_1083);
xor U2080 (N_2080,N_1852,N_1959);
nor U2081 (N_2081,N_1154,N_1777);
nand U2082 (N_2082,N_1620,N_1099);
nand U2083 (N_2083,N_1280,N_1487);
nor U2084 (N_2084,N_1008,N_1496);
and U2085 (N_2085,N_1460,N_1758);
and U2086 (N_2086,N_1076,N_1375);
nand U2087 (N_2087,N_1656,N_1382);
nor U2088 (N_2088,N_1394,N_1276);
or U2089 (N_2089,N_1955,N_1495);
nand U2090 (N_2090,N_1608,N_1957);
nor U2091 (N_2091,N_1654,N_1027);
nor U2092 (N_2092,N_1360,N_1127);
or U2093 (N_2093,N_1497,N_1364);
or U2094 (N_2094,N_1952,N_1058);
nor U2095 (N_2095,N_1017,N_1431);
nand U2096 (N_2096,N_1030,N_1430);
xor U2097 (N_2097,N_1004,N_1753);
and U2098 (N_2098,N_1518,N_1274);
nand U2099 (N_2099,N_1082,N_1312);
and U2100 (N_2100,N_1861,N_1728);
nor U2101 (N_2101,N_1501,N_1128);
nand U2102 (N_2102,N_1242,N_1594);
and U2103 (N_2103,N_1529,N_1929);
xor U2104 (N_2104,N_1468,N_1036);
or U2105 (N_2105,N_1208,N_1616);
and U2106 (N_2106,N_1742,N_1676);
nor U2107 (N_2107,N_1581,N_1308);
nor U2108 (N_2108,N_1493,N_1822);
or U2109 (N_2109,N_1942,N_1711);
xnor U2110 (N_2110,N_1200,N_1326);
nor U2111 (N_2111,N_1456,N_1556);
nor U2112 (N_2112,N_1172,N_1992);
nand U2113 (N_2113,N_1377,N_1831);
nand U2114 (N_2114,N_1792,N_1572);
nor U2115 (N_2115,N_1848,N_1882);
nor U2116 (N_2116,N_1787,N_1673);
nand U2117 (N_2117,N_1494,N_1024);
or U2118 (N_2118,N_1121,N_1198);
and U2119 (N_2119,N_1836,N_1956);
or U2120 (N_2120,N_1489,N_1136);
nand U2121 (N_2121,N_1435,N_1119);
nand U2122 (N_2122,N_1981,N_1686);
nor U2123 (N_2123,N_1111,N_1315);
xor U2124 (N_2124,N_1803,N_1120);
xor U2125 (N_2125,N_1974,N_1131);
nand U2126 (N_2126,N_1896,N_1170);
xnor U2127 (N_2127,N_1486,N_1778);
nand U2128 (N_2128,N_1373,N_1596);
nor U2129 (N_2129,N_1864,N_1370);
nor U2130 (N_2130,N_1592,N_1696);
xor U2131 (N_2131,N_1132,N_1901);
xor U2132 (N_2132,N_1249,N_1801);
nor U2133 (N_2133,N_1721,N_1478);
or U2134 (N_2134,N_1389,N_1573);
or U2135 (N_2135,N_1400,N_1873);
and U2136 (N_2136,N_1190,N_1422);
and U2137 (N_2137,N_1718,N_1839);
or U2138 (N_2138,N_1269,N_1465);
xor U2139 (N_2139,N_1970,N_1145);
or U2140 (N_2140,N_1597,N_1940);
nand U2141 (N_2141,N_1442,N_1338);
or U2142 (N_2142,N_1569,N_1386);
nor U2143 (N_2143,N_1603,N_1492);
or U2144 (N_2144,N_1910,N_1175);
nand U2145 (N_2145,N_1196,N_1085);
or U2146 (N_2146,N_1226,N_1948);
and U2147 (N_2147,N_1271,N_1779);
xnor U2148 (N_2148,N_1176,N_1943);
or U2149 (N_2149,N_1197,N_1255);
nor U2150 (N_2150,N_1126,N_1797);
nor U2151 (N_2151,N_1930,N_1677);
or U2152 (N_2152,N_1071,N_1371);
or U2153 (N_2153,N_1251,N_1946);
nor U2154 (N_2154,N_1833,N_1643);
nand U2155 (N_2155,N_1563,N_1648);
and U2156 (N_2156,N_1202,N_1333);
nor U2157 (N_2157,N_1727,N_1048);
and U2158 (N_2158,N_1328,N_1130);
xor U2159 (N_2159,N_1516,N_1544);
or U2160 (N_2160,N_1709,N_1612);
xnor U2161 (N_2161,N_1039,N_1911);
or U2162 (N_2162,N_1006,N_1966);
nor U2163 (N_2163,N_1895,N_1233);
and U2164 (N_2164,N_1591,N_1512);
nand U2165 (N_2165,N_1850,N_1533);
xnor U2166 (N_2166,N_1977,N_1628);
and U2167 (N_2167,N_1949,N_1793);
nor U2168 (N_2168,N_1352,N_1134);
xor U2169 (N_2169,N_1481,N_1824);
and U2170 (N_2170,N_1313,N_1214);
or U2171 (N_2171,N_1026,N_1666);
nand U2172 (N_2172,N_1546,N_1690);
nor U2173 (N_2173,N_1587,N_1412);
xnor U2174 (N_2174,N_1217,N_1565);
or U2175 (N_2175,N_1610,N_1346);
nor U2176 (N_2176,N_1644,N_1104);
and U2177 (N_2177,N_1972,N_1703);
xor U2178 (N_2178,N_1282,N_1645);
xnor U2179 (N_2179,N_1786,N_1461);
or U2180 (N_2180,N_1498,N_1986);
nor U2181 (N_2181,N_1700,N_1936);
or U2182 (N_2182,N_1606,N_1467);
nand U2183 (N_2183,N_1821,N_1647);
nand U2184 (N_2184,N_1007,N_1220);
and U2185 (N_2185,N_1840,N_1434);
or U2186 (N_2186,N_1103,N_1744);
xnor U2187 (N_2187,N_1726,N_1984);
xor U2188 (N_2188,N_1256,N_1087);
nand U2189 (N_2189,N_1019,N_1421);
and U2190 (N_2190,N_1739,N_1950);
xor U2191 (N_2191,N_1697,N_1025);
nor U2192 (N_2192,N_1543,N_1764);
xnor U2193 (N_2193,N_1416,N_1485);
nor U2194 (N_2194,N_1000,N_1303);
xnor U2195 (N_2195,N_1759,N_1650);
nor U2196 (N_2196,N_1995,N_1668);
and U2197 (N_2197,N_1752,N_1133);
or U2198 (N_2198,N_1655,N_1034);
nand U2199 (N_2199,N_1195,N_1244);
nor U2200 (N_2200,N_1773,N_1148);
nand U2201 (N_2201,N_1828,N_1588);
xor U2202 (N_2202,N_1715,N_1102);
or U2203 (N_2203,N_1684,N_1158);
xor U2204 (N_2204,N_1997,N_1201);
xor U2205 (N_2205,N_1279,N_1216);
nand U2206 (N_2206,N_1252,N_1682);
xnor U2207 (N_2207,N_1527,N_1031);
and U2208 (N_2208,N_1339,N_1155);
or U2209 (N_2209,N_1920,N_1064);
nor U2210 (N_2210,N_1740,N_1403);
or U2211 (N_2211,N_1471,N_1523);
nor U2212 (N_2212,N_1221,N_1392);
nand U2213 (N_2213,N_1323,N_1239);
nor U2214 (N_2214,N_1798,N_1755);
nor U2215 (N_2215,N_1708,N_1598);
nand U2216 (N_2216,N_1367,N_1894);
xnor U2217 (N_2217,N_1151,N_1875);
and U2218 (N_2218,N_1225,N_1913);
xor U2219 (N_2219,N_1053,N_1301);
nor U2220 (N_2220,N_1552,N_1329);
xnor U2221 (N_2221,N_1078,N_1919);
or U2222 (N_2222,N_1542,N_1436);
nand U2223 (N_2223,N_1576,N_1288);
and U2224 (N_2224,N_1473,N_1157);
nand U2225 (N_2225,N_1823,N_1754);
nand U2226 (N_2226,N_1692,N_1819);
nor U2227 (N_2227,N_1685,N_1638);
xor U2228 (N_2228,N_1038,N_1745);
and U2229 (N_2229,N_1362,N_1561);
nor U2230 (N_2230,N_1862,N_1420);
or U2231 (N_2231,N_1877,N_1880);
or U2232 (N_2232,N_1224,N_1156);
nand U2233 (N_2233,N_1474,N_1433);
xnor U2234 (N_2234,N_1866,N_1052);
and U2235 (N_2235,N_1622,N_1402);
nor U2236 (N_2236,N_1012,N_1021);
or U2237 (N_2237,N_1354,N_1450);
xnor U2238 (N_2238,N_1293,N_1163);
nand U2239 (N_2239,N_1999,N_1810);
or U2240 (N_2240,N_1525,N_1750);
nand U2241 (N_2241,N_1614,N_1390);
nand U2242 (N_2242,N_1147,N_1536);
and U2243 (N_2243,N_1250,N_1843);
xnor U2244 (N_2244,N_1664,N_1817);
and U2245 (N_2245,N_1808,N_1453);
nor U2246 (N_2246,N_1705,N_1490);
nor U2247 (N_2247,N_1041,N_1177);
and U2248 (N_2248,N_1965,N_1417);
nor U2249 (N_2249,N_1870,N_1751);
nand U2250 (N_2250,N_1670,N_1567);
nand U2251 (N_2251,N_1186,N_1907);
or U2252 (N_2252,N_1365,N_1729);
nor U2253 (N_2253,N_1618,N_1419);
or U2254 (N_2254,N_1005,N_1503);
nand U2255 (N_2255,N_1235,N_1807);
nor U2256 (N_2256,N_1043,N_1776);
xnor U2257 (N_2257,N_1897,N_1674);
or U2258 (N_2258,N_1347,N_1874);
xor U2259 (N_2259,N_1617,N_1245);
nand U2260 (N_2260,N_1883,N_1660);
nor U2261 (N_2261,N_1259,N_1463);
and U2262 (N_2262,N_1915,N_1590);
and U2263 (N_2263,N_1757,N_1621);
nand U2264 (N_2264,N_1555,N_1028);
nand U2265 (N_2265,N_1452,N_1060);
xnor U2266 (N_2266,N_1733,N_1425);
xnor U2267 (N_2267,N_1183,N_1016);
xor U2268 (N_2268,N_1585,N_1557);
xor U2269 (N_2269,N_1967,N_1234);
xnor U2270 (N_2270,N_1505,N_1800);
or U2271 (N_2271,N_1475,N_1278);
nor U2272 (N_2272,N_1059,N_1921);
nor U2273 (N_2273,N_1806,N_1139);
nand U2274 (N_2274,N_1470,N_1712);
and U2275 (N_2275,N_1291,N_1969);
or U2276 (N_2276,N_1982,N_1173);
nor U2277 (N_2277,N_1586,N_1261);
nand U2278 (N_2278,N_1063,N_1152);
or U2279 (N_2279,N_1337,N_1756);
nand U2280 (N_2280,N_1602,N_1722);
and U2281 (N_2281,N_1918,N_1268);
nor U2282 (N_2282,N_1414,N_1438);
and U2283 (N_2283,N_1054,N_1706);
nand U2284 (N_2284,N_1863,N_1050);
and U2285 (N_2285,N_1820,N_1925);
nand U2286 (N_2286,N_1855,N_1802);
nand U2287 (N_2287,N_1604,N_1772);
or U2288 (N_2288,N_1502,N_1826);
and U2289 (N_2289,N_1169,N_1353);
xnor U2290 (N_2290,N_1182,N_1482);
nor U2291 (N_2291,N_1607,N_1566);
or U2292 (N_2292,N_1075,N_1785);
or U2293 (N_2293,N_1273,N_1096);
xor U2294 (N_2294,N_1858,N_1113);
nand U2295 (N_2295,N_1511,N_1506);
xnor U2296 (N_2296,N_1361,N_1504);
nor U2297 (N_2297,N_1193,N_1926);
and U2298 (N_2298,N_1162,N_1399);
xnor U2299 (N_2299,N_1517,N_1663);
or U2300 (N_2300,N_1725,N_1735);
nor U2301 (N_2301,N_1238,N_1922);
xnor U2302 (N_2302,N_1781,N_1396);
xor U2303 (N_2303,N_1035,N_1968);
nand U2304 (N_2304,N_1209,N_1285);
nand U2305 (N_2305,N_1710,N_1023);
or U2306 (N_2306,N_1691,N_1228);
xor U2307 (N_2307,N_1613,N_1332);
and U2308 (N_2308,N_1961,N_1359);
or U2309 (N_2309,N_1743,N_1014);
nand U2310 (N_2310,N_1299,N_1960);
nand U2311 (N_2311,N_1642,N_1780);
nor U2312 (N_2312,N_1865,N_1931);
xor U2313 (N_2313,N_1941,N_1979);
nor U2314 (N_2314,N_1310,N_1766);
and U2315 (N_2315,N_1439,N_1879);
xor U2316 (N_2316,N_1304,N_1671);
nor U2317 (N_2317,N_1343,N_1372);
xnor U2318 (N_2318,N_1123,N_1215);
nor U2319 (N_2319,N_1090,N_1669);
xor U2320 (N_2320,N_1248,N_1953);
xor U2321 (N_2321,N_1988,N_1784);
and U2322 (N_2322,N_1218,N_1437);
nand U2323 (N_2323,N_1061,N_1286);
nor U2324 (N_2324,N_1300,N_1444);
and U2325 (N_2325,N_1749,N_1171);
and U2326 (N_2326,N_1185,N_1551);
or U2327 (N_2327,N_1292,N_1287);
or U2328 (N_2328,N_1040,N_1307);
and U2329 (N_2329,N_1985,N_1804);
or U2330 (N_2330,N_1524,N_1289);
nand U2331 (N_2331,N_1112,N_1584);
and U2332 (N_2332,N_1927,N_1632);
nor U2333 (N_2333,N_1340,N_1938);
and U2334 (N_2334,N_1575,N_1513);
and U2335 (N_2335,N_1748,N_1615);
or U2336 (N_2336,N_1117,N_1384);
nor U2337 (N_2337,N_1652,N_1484);
nor U2338 (N_2338,N_1827,N_1223);
xnor U2339 (N_2339,N_1906,N_1318);
nand U2340 (N_2340,N_1675,N_1954);
xor U2341 (N_2341,N_1631,N_1813);
or U2342 (N_2342,N_1110,N_1559);
nor U2343 (N_2343,N_1488,N_1734);
nor U2344 (N_2344,N_1933,N_1579);
and U2345 (N_2345,N_1665,N_1203);
xor U2346 (N_2346,N_1167,N_1541);
or U2347 (N_2347,N_1088,N_1747);
or U2348 (N_2348,N_1084,N_1845);
nor U2349 (N_2349,N_1932,N_1891);
nand U2350 (N_2350,N_1876,N_1775);
or U2351 (N_2351,N_1832,N_1816);
nand U2352 (N_2352,N_1368,N_1281);
or U2353 (N_2353,N_1601,N_1194);
nand U2354 (N_2354,N_1409,N_1144);
or U2355 (N_2355,N_1166,N_1769);
or U2356 (N_2356,N_1998,N_1296);
nor U2357 (N_2357,N_1179,N_1683);
nor U2358 (N_2358,N_1741,N_1106);
xnor U2359 (N_2359,N_1900,N_1265);
and U2360 (N_2360,N_1963,N_1851);
nand U2361 (N_2361,N_1657,N_1331);
xnor U2362 (N_2362,N_1407,N_1888);
nand U2363 (N_2363,N_1330,N_1311);
nand U2364 (N_2364,N_1317,N_1681);
nand U2365 (N_2365,N_1695,N_1294);
or U2366 (N_2366,N_1991,N_1914);
or U2367 (N_2367,N_1689,N_1886);
nor U2368 (N_2368,N_1272,N_1640);
nor U2369 (N_2369,N_1393,N_1987);
or U2370 (N_2370,N_1993,N_1589);
and U2371 (N_2371,N_1297,N_1558);
nand U2372 (N_2372,N_1796,N_1164);
xor U2373 (N_2373,N_1476,N_1095);
xnor U2374 (N_2374,N_1716,N_1916);
xnor U2375 (N_2375,N_1424,N_1464);
nor U2376 (N_2376,N_1625,N_1118);
nor U2377 (N_2377,N_1107,N_1207);
nor U2378 (N_2378,N_1547,N_1633);
and U2379 (N_2379,N_1909,N_1334);
nor U2380 (N_2380,N_1564,N_1100);
and U2381 (N_2381,N_1227,N_1124);
xnor U2382 (N_2382,N_1719,N_1577);
and U2383 (N_2383,N_1146,N_1115);
or U2384 (N_2384,N_1098,N_1535);
and U2385 (N_2385,N_1092,N_1947);
nand U2386 (N_2386,N_1013,N_1427);
and U2387 (N_2387,N_1199,N_1345);
nand U2388 (N_2388,N_1070,N_1699);
nor U2389 (N_2389,N_1908,N_1138);
or U2390 (N_2390,N_1534,N_1760);
and U2391 (N_2391,N_1413,N_1509);
xnor U2392 (N_2392,N_1627,N_1835);
xnor U2393 (N_2393,N_1451,N_1646);
or U2394 (N_2394,N_1305,N_1266);
and U2395 (N_2395,N_1344,N_1447);
nand U2396 (N_2396,N_1996,N_1379);
nand U2397 (N_2397,N_1237,N_1010);
nor U2398 (N_2398,N_1029,N_1231);
xnor U2399 (N_2399,N_1550,N_1507);
xor U2400 (N_2400,N_1322,N_1395);
or U2401 (N_2401,N_1341,N_1521);
nor U2402 (N_2402,N_1869,N_1530);
xor U2403 (N_2403,N_1924,N_1962);
nand U2404 (N_2404,N_1459,N_1477);
and U2405 (N_2405,N_1859,N_1898);
xor U2406 (N_2406,N_1159,N_1688);
xnor U2407 (N_2407,N_1109,N_1247);
and U2408 (N_2408,N_1846,N_1260);
and U2409 (N_2409,N_1678,N_1623);
nor U2410 (N_2410,N_1165,N_1672);
xnor U2411 (N_2411,N_1553,N_1045);
nand U2412 (N_2412,N_1522,N_1263);
or U2413 (N_2413,N_1206,N_1635);
nor U2414 (N_2414,N_1073,N_1037);
or U2415 (N_2415,N_1257,N_1351);
xnor U2416 (N_2416,N_1661,N_1520);
xnor U2417 (N_2417,N_1355,N_1951);
nand U2418 (N_2418,N_1531,N_1325);
xor U2419 (N_2419,N_1830,N_1790);
xor U2420 (N_2420,N_1184,N_1624);
and U2421 (N_2421,N_1472,N_1582);
and U2422 (N_2422,N_1174,N_1944);
xor U2423 (N_2423,N_1639,N_1514);
nand U2424 (N_2424,N_1210,N_1549);
xor U2425 (N_2425,N_1761,N_1405);
and U2426 (N_2426,N_1871,N_1720);
or U2427 (N_2427,N_1466,N_1902);
or U2428 (N_2428,N_1074,N_1641);
and U2429 (N_2429,N_1042,N_1129);
xor U2430 (N_2430,N_1069,N_1406);
nor U2431 (N_2431,N_1973,N_1707);
nand U2432 (N_2432,N_1659,N_1904);
and U2433 (N_2433,N_1077,N_1687);
and U2434 (N_2434,N_1805,N_1538);
xnor U2435 (N_2435,N_1812,N_1009);
xnor U2436 (N_2436,N_1736,N_1314);
nand U2437 (N_2437,N_1568,N_1526);
nor U2438 (N_2438,N_1560,N_1051);
and U2439 (N_2439,N_1693,N_1528);
or U2440 (N_2440,N_1056,N_1277);
nor U2441 (N_2441,N_1771,N_1980);
xnor U2442 (N_2442,N_1698,N_1983);
and U2443 (N_2443,N_1469,N_1768);
nand U2444 (N_2444,N_1302,N_1191);
or U2445 (N_2445,N_1213,N_1574);
nor U2446 (N_2446,N_1321,N_1842);
or U2447 (N_2447,N_1881,N_1611);
nand U2448 (N_2448,N_1181,N_1423);
nand U2449 (N_2449,N_1411,N_1730);
or U2450 (N_2450,N_1905,N_1189);
or U2451 (N_2451,N_1062,N_1383);
or U2452 (N_2452,N_1702,N_1418);
nand U2453 (N_2453,N_1717,N_1701);
nor U2454 (N_2454,N_1366,N_1548);
xnor U2455 (N_2455,N_1783,N_1369);
nor U2456 (N_2456,N_1532,N_1455);
and U2457 (N_2457,N_1003,N_1020);
or U2458 (N_2458,N_1408,N_1141);
and U2459 (N_2459,N_1679,N_1270);
xnor U2460 (N_2460,N_1001,N_1500);
and U2461 (N_2461,N_1825,N_1290);
nor U2462 (N_2462,N_1081,N_1388);
or U2463 (N_2463,N_1348,N_1658);
nor U2464 (N_2464,N_1398,N_1241);
and U2465 (N_2465,N_1324,N_1629);
or U2466 (N_2466,N_1856,N_1746);
or U2467 (N_2467,N_1283,N_1018);
nand U2468 (N_2468,N_1890,N_1767);
or U2469 (N_2469,N_1600,N_1232);
nand U2470 (N_2470,N_1537,N_1349);
xor U2471 (N_2471,N_1067,N_1358);
xor U2472 (N_2472,N_1789,N_1694);
nor U2473 (N_2473,N_1794,N_1047);
nand U2474 (N_2474,N_1732,N_1309);
xor U2475 (N_2475,N_1236,N_1192);
xnor U2476 (N_2476,N_1230,N_1295);
and U2477 (N_2477,N_1049,N_1837);
nand U2478 (N_2478,N_1723,N_1376);
or U2479 (N_2479,N_1449,N_1731);
nor U2480 (N_2480,N_1562,N_1457);
and U2481 (N_2481,N_1928,N_1818);
xnor U2482 (N_2482,N_1867,N_1667);
and U2483 (N_2483,N_1788,N_1065);
xnor U2484 (N_2484,N_1205,N_1838);
nand U2485 (N_2485,N_1387,N_1178);
nor U2486 (N_2486,N_1540,N_1958);
xnor U2487 (N_2487,N_1022,N_1714);
nor U2488 (N_2488,N_1033,N_1135);
xnor U2489 (N_2489,N_1116,N_1298);
nand U2490 (N_2490,N_1868,N_1649);
nand U2491 (N_2491,N_1336,N_1086);
nor U2492 (N_2492,N_1510,N_1508);
xnor U2493 (N_2493,N_1903,N_1912);
nand U2494 (N_2494,N_1923,N_1441);
xor U2495 (N_2495,N_1491,N_1990);
xnor U2496 (N_2496,N_1378,N_1515);
or U2497 (N_2497,N_1770,N_1935);
or U2498 (N_2498,N_1080,N_1316);
nor U2499 (N_2499,N_1815,N_1015);
xor U2500 (N_2500,N_1284,N_1935);
or U2501 (N_2501,N_1686,N_1446);
nand U2502 (N_2502,N_1401,N_1708);
nor U2503 (N_2503,N_1162,N_1269);
nand U2504 (N_2504,N_1781,N_1940);
nand U2505 (N_2505,N_1235,N_1852);
nor U2506 (N_2506,N_1252,N_1042);
or U2507 (N_2507,N_1270,N_1135);
nor U2508 (N_2508,N_1099,N_1845);
nand U2509 (N_2509,N_1804,N_1173);
nand U2510 (N_2510,N_1658,N_1272);
or U2511 (N_2511,N_1329,N_1019);
nor U2512 (N_2512,N_1604,N_1554);
nor U2513 (N_2513,N_1801,N_1648);
and U2514 (N_2514,N_1763,N_1159);
nand U2515 (N_2515,N_1920,N_1388);
and U2516 (N_2516,N_1403,N_1321);
or U2517 (N_2517,N_1737,N_1307);
nand U2518 (N_2518,N_1538,N_1125);
nor U2519 (N_2519,N_1169,N_1872);
xor U2520 (N_2520,N_1238,N_1708);
nor U2521 (N_2521,N_1880,N_1052);
or U2522 (N_2522,N_1052,N_1434);
nor U2523 (N_2523,N_1466,N_1007);
xor U2524 (N_2524,N_1453,N_1986);
nand U2525 (N_2525,N_1908,N_1130);
and U2526 (N_2526,N_1140,N_1988);
and U2527 (N_2527,N_1919,N_1043);
and U2528 (N_2528,N_1527,N_1594);
xor U2529 (N_2529,N_1726,N_1927);
and U2530 (N_2530,N_1189,N_1351);
nor U2531 (N_2531,N_1879,N_1798);
nand U2532 (N_2532,N_1968,N_1800);
or U2533 (N_2533,N_1748,N_1473);
nor U2534 (N_2534,N_1055,N_1074);
or U2535 (N_2535,N_1021,N_1936);
and U2536 (N_2536,N_1435,N_1583);
nand U2537 (N_2537,N_1077,N_1886);
xor U2538 (N_2538,N_1882,N_1826);
nor U2539 (N_2539,N_1854,N_1720);
nand U2540 (N_2540,N_1244,N_1302);
or U2541 (N_2541,N_1202,N_1987);
nor U2542 (N_2542,N_1754,N_1971);
nand U2543 (N_2543,N_1090,N_1714);
and U2544 (N_2544,N_1166,N_1517);
nand U2545 (N_2545,N_1599,N_1064);
nand U2546 (N_2546,N_1473,N_1839);
or U2547 (N_2547,N_1668,N_1526);
nand U2548 (N_2548,N_1375,N_1550);
xnor U2549 (N_2549,N_1755,N_1782);
xor U2550 (N_2550,N_1328,N_1433);
nor U2551 (N_2551,N_1820,N_1658);
nand U2552 (N_2552,N_1424,N_1930);
or U2553 (N_2553,N_1892,N_1060);
xnor U2554 (N_2554,N_1716,N_1065);
and U2555 (N_2555,N_1520,N_1580);
nand U2556 (N_2556,N_1568,N_1509);
or U2557 (N_2557,N_1055,N_1007);
nand U2558 (N_2558,N_1983,N_1639);
and U2559 (N_2559,N_1423,N_1035);
xor U2560 (N_2560,N_1640,N_1522);
nand U2561 (N_2561,N_1914,N_1480);
xor U2562 (N_2562,N_1550,N_1702);
xor U2563 (N_2563,N_1422,N_1354);
or U2564 (N_2564,N_1202,N_1353);
nor U2565 (N_2565,N_1509,N_1156);
xor U2566 (N_2566,N_1150,N_1471);
or U2567 (N_2567,N_1267,N_1228);
or U2568 (N_2568,N_1588,N_1048);
nor U2569 (N_2569,N_1021,N_1703);
nor U2570 (N_2570,N_1921,N_1552);
xor U2571 (N_2571,N_1029,N_1947);
and U2572 (N_2572,N_1269,N_1564);
or U2573 (N_2573,N_1366,N_1561);
or U2574 (N_2574,N_1435,N_1266);
nand U2575 (N_2575,N_1429,N_1126);
or U2576 (N_2576,N_1393,N_1834);
or U2577 (N_2577,N_1896,N_1406);
or U2578 (N_2578,N_1889,N_1587);
xor U2579 (N_2579,N_1594,N_1403);
and U2580 (N_2580,N_1584,N_1050);
or U2581 (N_2581,N_1556,N_1596);
or U2582 (N_2582,N_1254,N_1982);
nand U2583 (N_2583,N_1856,N_1394);
nor U2584 (N_2584,N_1605,N_1772);
or U2585 (N_2585,N_1862,N_1181);
nor U2586 (N_2586,N_1216,N_1848);
and U2587 (N_2587,N_1827,N_1813);
xor U2588 (N_2588,N_1122,N_1701);
nand U2589 (N_2589,N_1666,N_1325);
nor U2590 (N_2590,N_1579,N_1201);
nand U2591 (N_2591,N_1615,N_1390);
nor U2592 (N_2592,N_1538,N_1020);
nor U2593 (N_2593,N_1261,N_1836);
xor U2594 (N_2594,N_1861,N_1739);
xor U2595 (N_2595,N_1496,N_1773);
xnor U2596 (N_2596,N_1253,N_1639);
xnor U2597 (N_2597,N_1862,N_1685);
nand U2598 (N_2598,N_1279,N_1669);
and U2599 (N_2599,N_1577,N_1759);
nor U2600 (N_2600,N_1584,N_1257);
and U2601 (N_2601,N_1505,N_1297);
or U2602 (N_2602,N_1912,N_1992);
nand U2603 (N_2603,N_1335,N_1288);
and U2604 (N_2604,N_1286,N_1736);
xor U2605 (N_2605,N_1499,N_1835);
or U2606 (N_2606,N_1186,N_1316);
xor U2607 (N_2607,N_1447,N_1500);
nor U2608 (N_2608,N_1250,N_1564);
and U2609 (N_2609,N_1703,N_1123);
nand U2610 (N_2610,N_1916,N_1359);
nor U2611 (N_2611,N_1575,N_1557);
xor U2612 (N_2612,N_1281,N_1885);
and U2613 (N_2613,N_1391,N_1226);
nor U2614 (N_2614,N_1587,N_1182);
and U2615 (N_2615,N_1420,N_1601);
and U2616 (N_2616,N_1223,N_1872);
nand U2617 (N_2617,N_1653,N_1056);
nor U2618 (N_2618,N_1951,N_1282);
and U2619 (N_2619,N_1562,N_1534);
nor U2620 (N_2620,N_1583,N_1328);
nand U2621 (N_2621,N_1639,N_1930);
nor U2622 (N_2622,N_1939,N_1744);
nor U2623 (N_2623,N_1747,N_1395);
or U2624 (N_2624,N_1692,N_1380);
nand U2625 (N_2625,N_1042,N_1736);
nand U2626 (N_2626,N_1613,N_1066);
xnor U2627 (N_2627,N_1767,N_1776);
and U2628 (N_2628,N_1250,N_1708);
nor U2629 (N_2629,N_1722,N_1811);
nand U2630 (N_2630,N_1462,N_1856);
and U2631 (N_2631,N_1703,N_1285);
nor U2632 (N_2632,N_1616,N_1969);
nor U2633 (N_2633,N_1172,N_1505);
nor U2634 (N_2634,N_1590,N_1472);
nor U2635 (N_2635,N_1720,N_1855);
and U2636 (N_2636,N_1755,N_1756);
nor U2637 (N_2637,N_1098,N_1003);
and U2638 (N_2638,N_1601,N_1313);
and U2639 (N_2639,N_1274,N_1581);
and U2640 (N_2640,N_1949,N_1077);
xor U2641 (N_2641,N_1105,N_1675);
and U2642 (N_2642,N_1599,N_1698);
xnor U2643 (N_2643,N_1698,N_1973);
and U2644 (N_2644,N_1461,N_1057);
nand U2645 (N_2645,N_1372,N_1569);
nor U2646 (N_2646,N_1018,N_1922);
and U2647 (N_2647,N_1348,N_1300);
nor U2648 (N_2648,N_1856,N_1635);
nand U2649 (N_2649,N_1446,N_1203);
and U2650 (N_2650,N_1230,N_1462);
or U2651 (N_2651,N_1603,N_1289);
or U2652 (N_2652,N_1263,N_1257);
or U2653 (N_2653,N_1630,N_1603);
nor U2654 (N_2654,N_1005,N_1211);
nand U2655 (N_2655,N_1238,N_1247);
and U2656 (N_2656,N_1434,N_1412);
or U2657 (N_2657,N_1864,N_1865);
nand U2658 (N_2658,N_1403,N_1129);
nand U2659 (N_2659,N_1110,N_1718);
nor U2660 (N_2660,N_1788,N_1486);
and U2661 (N_2661,N_1392,N_1010);
xor U2662 (N_2662,N_1688,N_1377);
nor U2663 (N_2663,N_1309,N_1288);
or U2664 (N_2664,N_1804,N_1946);
or U2665 (N_2665,N_1758,N_1167);
or U2666 (N_2666,N_1946,N_1919);
xnor U2667 (N_2667,N_1324,N_1102);
and U2668 (N_2668,N_1265,N_1761);
nand U2669 (N_2669,N_1453,N_1595);
nand U2670 (N_2670,N_1004,N_1101);
nor U2671 (N_2671,N_1119,N_1770);
nor U2672 (N_2672,N_1201,N_1807);
or U2673 (N_2673,N_1807,N_1519);
xor U2674 (N_2674,N_1346,N_1622);
nand U2675 (N_2675,N_1984,N_1270);
nor U2676 (N_2676,N_1502,N_1204);
nor U2677 (N_2677,N_1346,N_1307);
nor U2678 (N_2678,N_1568,N_1119);
nor U2679 (N_2679,N_1238,N_1467);
or U2680 (N_2680,N_1752,N_1294);
or U2681 (N_2681,N_1224,N_1227);
and U2682 (N_2682,N_1680,N_1965);
nor U2683 (N_2683,N_1553,N_1535);
or U2684 (N_2684,N_1313,N_1841);
xor U2685 (N_2685,N_1196,N_1949);
and U2686 (N_2686,N_1870,N_1656);
nor U2687 (N_2687,N_1057,N_1638);
xnor U2688 (N_2688,N_1131,N_1829);
nand U2689 (N_2689,N_1031,N_1177);
nand U2690 (N_2690,N_1062,N_1716);
nor U2691 (N_2691,N_1888,N_1420);
xnor U2692 (N_2692,N_1896,N_1953);
xnor U2693 (N_2693,N_1065,N_1833);
xnor U2694 (N_2694,N_1612,N_1007);
or U2695 (N_2695,N_1178,N_1305);
xor U2696 (N_2696,N_1510,N_1816);
nand U2697 (N_2697,N_1930,N_1110);
and U2698 (N_2698,N_1682,N_1751);
nor U2699 (N_2699,N_1378,N_1357);
xnor U2700 (N_2700,N_1453,N_1690);
or U2701 (N_2701,N_1953,N_1324);
and U2702 (N_2702,N_1909,N_1022);
nor U2703 (N_2703,N_1622,N_1103);
xnor U2704 (N_2704,N_1921,N_1240);
xnor U2705 (N_2705,N_1170,N_1685);
and U2706 (N_2706,N_1879,N_1815);
or U2707 (N_2707,N_1055,N_1360);
and U2708 (N_2708,N_1060,N_1969);
or U2709 (N_2709,N_1542,N_1794);
nand U2710 (N_2710,N_1538,N_1890);
nor U2711 (N_2711,N_1890,N_1635);
nand U2712 (N_2712,N_1691,N_1909);
xor U2713 (N_2713,N_1048,N_1745);
and U2714 (N_2714,N_1825,N_1217);
nor U2715 (N_2715,N_1941,N_1384);
nand U2716 (N_2716,N_1265,N_1489);
and U2717 (N_2717,N_1318,N_1248);
and U2718 (N_2718,N_1124,N_1323);
or U2719 (N_2719,N_1673,N_1004);
nor U2720 (N_2720,N_1722,N_1103);
nand U2721 (N_2721,N_1228,N_1422);
nand U2722 (N_2722,N_1755,N_1893);
xor U2723 (N_2723,N_1530,N_1760);
xnor U2724 (N_2724,N_1139,N_1347);
or U2725 (N_2725,N_1759,N_1084);
nor U2726 (N_2726,N_1347,N_1684);
or U2727 (N_2727,N_1543,N_1121);
and U2728 (N_2728,N_1735,N_1210);
xor U2729 (N_2729,N_1423,N_1731);
xnor U2730 (N_2730,N_1045,N_1802);
nand U2731 (N_2731,N_1686,N_1330);
and U2732 (N_2732,N_1355,N_1693);
nand U2733 (N_2733,N_1418,N_1106);
nor U2734 (N_2734,N_1229,N_1988);
and U2735 (N_2735,N_1055,N_1251);
or U2736 (N_2736,N_1535,N_1378);
and U2737 (N_2737,N_1851,N_1995);
nor U2738 (N_2738,N_1257,N_1666);
or U2739 (N_2739,N_1261,N_1192);
nand U2740 (N_2740,N_1077,N_1384);
xnor U2741 (N_2741,N_1649,N_1238);
nand U2742 (N_2742,N_1894,N_1223);
nor U2743 (N_2743,N_1871,N_1927);
and U2744 (N_2744,N_1857,N_1806);
nand U2745 (N_2745,N_1946,N_1247);
nor U2746 (N_2746,N_1851,N_1820);
or U2747 (N_2747,N_1458,N_1461);
xor U2748 (N_2748,N_1476,N_1096);
nor U2749 (N_2749,N_1438,N_1768);
nand U2750 (N_2750,N_1775,N_1895);
and U2751 (N_2751,N_1397,N_1157);
xor U2752 (N_2752,N_1833,N_1300);
nand U2753 (N_2753,N_1114,N_1626);
xnor U2754 (N_2754,N_1773,N_1530);
or U2755 (N_2755,N_1578,N_1275);
nand U2756 (N_2756,N_1393,N_1848);
xnor U2757 (N_2757,N_1526,N_1477);
nor U2758 (N_2758,N_1872,N_1822);
and U2759 (N_2759,N_1727,N_1285);
nand U2760 (N_2760,N_1050,N_1273);
xnor U2761 (N_2761,N_1053,N_1378);
nor U2762 (N_2762,N_1199,N_1475);
or U2763 (N_2763,N_1700,N_1260);
xnor U2764 (N_2764,N_1795,N_1856);
and U2765 (N_2765,N_1326,N_1582);
xor U2766 (N_2766,N_1769,N_1896);
nor U2767 (N_2767,N_1537,N_1601);
and U2768 (N_2768,N_1666,N_1017);
nand U2769 (N_2769,N_1828,N_1165);
nor U2770 (N_2770,N_1280,N_1286);
nand U2771 (N_2771,N_1318,N_1601);
xnor U2772 (N_2772,N_1634,N_1684);
nand U2773 (N_2773,N_1581,N_1802);
xnor U2774 (N_2774,N_1193,N_1149);
or U2775 (N_2775,N_1590,N_1081);
and U2776 (N_2776,N_1399,N_1933);
and U2777 (N_2777,N_1405,N_1677);
nand U2778 (N_2778,N_1149,N_1216);
and U2779 (N_2779,N_1647,N_1361);
nand U2780 (N_2780,N_1367,N_1842);
xnor U2781 (N_2781,N_1730,N_1002);
nand U2782 (N_2782,N_1005,N_1409);
xnor U2783 (N_2783,N_1305,N_1495);
and U2784 (N_2784,N_1280,N_1405);
nor U2785 (N_2785,N_1716,N_1909);
nand U2786 (N_2786,N_1636,N_1886);
nand U2787 (N_2787,N_1412,N_1153);
nand U2788 (N_2788,N_1773,N_1880);
or U2789 (N_2789,N_1460,N_1071);
or U2790 (N_2790,N_1374,N_1260);
and U2791 (N_2791,N_1596,N_1816);
or U2792 (N_2792,N_1930,N_1992);
and U2793 (N_2793,N_1329,N_1781);
and U2794 (N_2794,N_1439,N_1135);
and U2795 (N_2795,N_1969,N_1243);
nor U2796 (N_2796,N_1718,N_1529);
nand U2797 (N_2797,N_1549,N_1527);
or U2798 (N_2798,N_1272,N_1331);
xor U2799 (N_2799,N_1167,N_1366);
nand U2800 (N_2800,N_1399,N_1317);
nor U2801 (N_2801,N_1113,N_1175);
xnor U2802 (N_2802,N_1138,N_1331);
or U2803 (N_2803,N_1647,N_1307);
or U2804 (N_2804,N_1994,N_1336);
or U2805 (N_2805,N_1282,N_1252);
nor U2806 (N_2806,N_1910,N_1326);
or U2807 (N_2807,N_1875,N_1902);
nor U2808 (N_2808,N_1813,N_1799);
and U2809 (N_2809,N_1797,N_1064);
xor U2810 (N_2810,N_1886,N_1440);
xnor U2811 (N_2811,N_1627,N_1706);
xor U2812 (N_2812,N_1357,N_1340);
and U2813 (N_2813,N_1080,N_1923);
xor U2814 (N_2814,N_1369,N_1608);
nand U2815 (N_2815,N_1107,N_1078);
and U2816 (N_2816,N_1663,N_1200);
and U2817 (N_2817,N_1077,N_1309);
or U2818 (N_2818,N_1540,N_1281);
or U2819 (N_2819,N_1933,N_1645);
and U2820 (N_2820,N_1115,N_1149);
or U2821 (N_2821,N_1550,N_1751);
xnor U2822 (N_2822,N_1143,N_1881);
nand U2823 (N_2823,N_1537,N_1788);
nor U2824 (N_2824,N_1601,N_1518);
or U2825 (N_2825,N_1468,N_1703);
and U2826 (N_2826,N_1887,N_1299);
xor U2827 (N_2827,N_1300,N_1023);
or U2828 (N_2828,N_1607,N_1340);
and U2829 (N_2829,N_1496,N_1541);
nor U2830 (N_2830,N_1940,N_1879);
nor U2831 (N_2831,N_1759,N_1730);
nor U2832 (N_2832,N_1839,N_1654);
nand U2833 (N_2833,N_1168,N_1093);
and U2834 (N_2834,N_1167,N_1019);
and U2835 (N_2835,N_1510,N_1260);
and U2836 (N_2836,N_1120,N_1200);
nor U2837 (N_2837,N_1499,N_1990);
or U2838 (N_2838,N_1363,N_1169);
or U2839 (N_2839,N_1424,N_1130);
nor U2840 (N_2840,N_1238,N_1864);
xnor U2841 (N_2841,N_1960,N_1892);
or U2842 (N_2842,N_1914,N_1567);
and U2843 (N_2843,N_1526,N_1607);
nor U2844 (N_2844,N_1995,N_1303);
nor U2845 (N_2845,N_1245,N_1130);
xnor U2846 (N_2846,N_1395,N_1147);
xnor U2847 (N_2847,N_1822,N_1616);
xor U2848 (N_2848,N_1049,N_1119);
xor U2849 (N_2849,N_1505,N_1554);
xnor U2850 (N_2850,N_1585,N_1359);
and U2851 (N_2851,N_1928,N_1943);
or U2852 (N_2852,N_1781,N_1180);
and U2853 (N_2853,N_1944,N_1788);
or U2854 (N_2854,N_1880,N_1268);
and U2855 (N_2855,N_1674,N_1278);
and U2856 (N_2856,N_1319,N_1083);
or U2857 (N_2857,N_1219,N_1000);
xnor U2858 (N_2858,N_1691,N_1479);
nor U2859 (N_2859,N_1542,N_1113);
or U2860 (N_2860,N_1599,N_1748);
or U2861 (N_2861,N_1039,N_1462);
xor U2862 (N_2862,N_1046,N_1658);
nand U2863 (N_2863,N_1987,N_1735);
nor U2864 (N_2864,N_1924,N_1473);
xor U2865 (N_2865,N_1713,N_1172);
nand U2866 (N_2866,N_1624,N_1413);
xnor U2867 (N_2867,N_1342,N_1572);
and U2868 (N_2868,N_1936,N_1629);
or U2869 (N_2869,N_1152,N_1245);
nand U2870 (N_2870,N_1179,N_1699);
and U2871 (N_2871,N_1665,N_1968);
nor U2872 (N_2872,N_1037,N_1735);
and U2873 (N_2873,N_1066,N_1045);
nor U2874 (N_2874,N_1836,N_1066);
or U2875 (N_2875,N_1030,N_1961);
nor U2876 (N_2876,N_1234,N_1982);
nand U2877 (N_2877,N_1129,N_1514);
or U2878 (N_2878,N_1521,N_1559);
and U2879 (N_2879,N_1042,N_1534);
or U2880 (N_2880,N_1081,N_1722);
nand U2881 (N_2881,N_1962,N_1855);
nand U2882 (N_2882,N_1589,N_1601);
or U2883 (N_2883,N_1979,N_1003);
and U2884 (N_2884,N_1621,N_1375);
nor U2885 (N_2885,N_1889,N_1982);
nor U2886 (N_2886,N_1079,N_1303);
and U2887 (N_2887,N_1674,N_1090);
or U2888 (N_2888,N_1345,N_1785);
nand U2889 (N_2889,N_1954,N_1715);
nand U2890 (N_2890,N_1168,N_1457);
nand U2891 (N_2891,N_1568,N_1828);
and U2892 (N_2892,N_1081,N_1750);
xor U2893 (N_2893,N_1191,N_1571);
xor U2894 (N_2894,N_1621,N_1024);
nand U2895 (N_2895,N_1239,N_1825);
or U2896 (N_2896,N_1109,N_1775);
nor U2897 (N_2897,N_1712,N_1509);
or U2898 (N_2898,N_1198,N_1645);
nand U2899 (N_2899,N_1154,N_1740);
or U2900 (N_2900,N_1762,N_1481);
nor U2901 (N_2901,N_1145,N_1573);
nand U2902 (N_2902,N_1245,N_1028);
xnor U2903 (N_2903,N_1282,N_1039);
xnor U2904 (N_2904,N_1637,N_1564);
xor U2905 (N_2905,N_1016,N_1510);
xor U2906 (N_2906,N_1625,N_1377);
nor U2907 (N_2907,N_1125,N_1763);
and U2908 (N_2908,N_1785,N_1357);
nand U2909 (N_2909,N_1610,N_1958);
and U2910 (N_2910,N_1585,N_1208);
or U2911 (N_2911,N_1724,N_1789);
and U2912 (N_2912,N_1586,N_1451);
xnor U2913 (N_2913,N_1739,N_1458);
nor U2914 (N_2914,N_1088,N_1814);
xor U2915 (N_2915,N_1851,N_1098);
xnor U2916 (N_2916,N_1389,N_1715);
and U2917 (N_2917,N_1580,N_1553);
and U2918 (N_2918,N_1820,N_1793);
xor U2919 (N_2919,N_1201,N_1124);
xor U2920 (N_2920,N_1050,N_1748);
xnor U2921 (N_2921,N_1503,N_1721);
or U2922 (N_2922,N_1734,N_1818);
and U2923 (N_2923,N_1698,N_1921);
xnor U2924 (N_2924,N_1442,N_1138);
and U2925 (N_2925,N_1267,N_1176);
xor U2926 (N_2926,N_1313,N_1749);
nor U2927 (N_2927,N_1956,N_1736);
xnor U2928 (N_2928,N_1861,N_1869);
xnor U2929 (N_2929,N_1286,N_1920);
nor U2930 (N_2930,N_1052,N_1817);
nor U2931 (N_2931,N_1599,N_1686);
xor U2932 (N_2932,N_1067,N_1221);
nor U2933 (N_2933,N_1523,N_1516);
nor U2934 (N_2934,N_1603,N_1303);
xnor U2935 (N_2935,N_1766,N_1238);
nand U2936 (N_2936,N_1574,N_1552);
xnor U2937 (N_2937,N_1156,N_1456);
nor U2938 (N_2938,N_1908,N_1673);
xor U2939 (N_2939,N_1649,N_1016);
nand U2940 (N_2940,N_1912,N_1522);
and U2941 (N_2941,N_1056,N_1572);
nor U2942 (N_2942,N_1279,N_1820);
xor U2943 (N_2943,N_1398,N_1836);
nor U2944 (N_2944,N_1444,N_1490);
and U2945 (N_2945,N_1005,N_1776);
or U2946 (N_2946,N_1758,N_1286);
and U2947 (N_2947,N_1089,N_1001);
nor U2948 (N_2948,N_1427,N_1862);
nand U2949 (N_2949,N_1021,N_1268);
and U2950 (N_2950,N_1071,N_1801);
or U2951 (N_2951,N_1573,N_1792);
xnor U2952 (N_2952,N_1330,N_1242);
and U2953 (N_2953,N_1152,N_1273);
nand U2954 (N_2954,N_1522,N_1967);
nand U2955 (N_2955,N_1406,N_1025);
and U2956 (N_2956,N_1053,N_1245);
or U2957 (N_2957,N_1330,N_1732);
nand U2958 (N_2958,N_1812,N_1601);
nor U2959 (N_2959,N_1855,N_1102);
nand U2960 (N_2960,N_1355,N_1039);
nor U2961 (N_2961,N_1355,N_1149);
or U2962 (N_2962,N_1803,N_1604);
xnor U2963 (N_2963,N_1899,N_1392);
and U2964 (N_2964,N_1957,N_1798);
xor U2965 (N_2965,N_1331,N_1690);
and U2966 (N_2966,N_1119,N_1638);
and U2967 (N_2967,N_1871,N_1911);
nand U2968 (N_2968,N_1630,N_1554);
xor U2969 (N_2969,N_1668,N_1438);
nand U2970 (N_2970,N_1838,N_1879);
and U2971 (N_2971,N_1853,N_1290);
nand U2972 (N_2972,N_1303,N_1468);
nand U2973 (N_2973,N_1949,N_1961);
nor U2974 (N_2974,N_1912,N_1897);
and U2975 (N_2975,N_1104,N_1868);
or U2976 (N_2976,N_1380,N_1724);
xnor U2977 (N_2977,N_1479,N_1704);
or U2978 (N_2978,N_1549,N_1845);
and U2979 (N_2979,N_1775,N_1130);
xor U2980 (N_2980,N_1799,N_1646);
nand U2981 (N_2981,N_1660,N_1172);
nor U2982 (N_2982,N_1866,N_1106);
nor U2983 (N_2983,N_1283,N_1809);
nand U2984 (N_2984,N_1955,N_1388);
nor U2985 (N_2985,N_1044,N_1335);
or U2986 (N_2986,N_1322,N_1356);
nand U2987 (N_2987,N_1005,N_1840);
nor U2988 (N_2988,N_1715,N_1713);
xnor U2989 (N_2989,N_1963,N_1955);
and U2990 (N_2990,N_1040,N_1695);
xnor U2991 (N_2991,N_1760,N_1604);
nand U2992 (N_2992,N_1712,N_1893);
or U2993 (N_2993,N_1418,N_1388);
or U2994 (N_2994,N_1243,N_1734);
nor U2995 (N_2995,N_1623,N_1868);
xor U2996 (N_2996,N_1822,N_1199);
and U2997 (N_2997,N_1101,N_1598);
and U2998 (N_2998,N_1223,N_1192);
and U2999 (N_2999,N_1063,N_1325);
nor U3000 (N_3000,N_2041,N_2337);
xor U3001 (N_3001,N_2058,N_2536);
nand U3002 (N_3002,N_2537,N_2001);
nor U3003 (N_3003,N_2121,N_2762);
nand U3004 (N_3004,N_2756,N_2033);
or U3005 (N_3005,N_2675,N_2543);
or U3006 (N_3006,N_2971,N_2046);
or U3007 (N_3007,N_2524,N_2115);
nand U3008 (N_3008,N_2890,N_2530);
or U3009 (N_3009,N_2790,N_2614);
nand U3010 (N_3010,N_2412,N_2110);
xor U3011 (N_3011,N_2229,N_2513);
or U3012 (N_3012,N_2887,N_2789);
xnor U3013 (N_3013,N_2132,N_2137);
xnor U3014 (N_3014,N_2146,N_2753);
and U3015 (N_3015,N_2959,N_2505);
xnor U3016 (N_3016,N_2651,N_2997);
xor U3017 (N_3017,N_2723,N_2181);
nor U3018 (N_3018,N_2244,N_2677);
nand U3019 (N_3019,N_2962,N_2160);
or U3020 (N_3020,N_2552,N_2005);
nor U3021 (N_3021,N_2938,N_2857);
nor U3022 (N_3022,N_2992,N_2426);
or U3023 (N_3023,N_2954,N_2573);
nor U3024 (N_3024,N_2764,N_2534);
nand U3025 (N_3025,N_2777,N_2429);
or U3026 (N_3026,N_2691,N_2193);
xor U3027 (N_3027,N_2101,N_2662);
and U3028 (N_3028,N_2681,N_2714);
xor U3029 (N_3029,N_2161,N_2162);
nand U3030 (N_3030,N_2230,N_2733);
xnor U3031 (N_3031,N_2682,N_2512);
or U3032 (N_3032,N_2563,N_2996);
nor U3033 (N_3033,N_2117,N_2361);
or U3034 (N_3034,N_2377,N_2523);
or U3035 (N_3035,N_2485,N_2297);
nor U3036 (N_3036,N_2170,N_2165);
and U3037 (N_3037,N_2641,N_2300);
nor U3038 (N_3038,N_2087,N_2519);
nand U3039 (N_3039,N_2974,N_2290);
nand U3040 (N_3040,N_2514,N_2478);
nand U3041 (N_3041,N_2815,N_2634);
nor U3042 (N_3042,N_2991,N_2249);
and U3043 (N_3043,N_2284,N_2551);
or U3044 (N_3044,N_2936,N_2602);
nand U3045 (N_3045,N_2555,N_2339);
xor U3046 (N_3046,N_2197,N_2596);
xor U3047 (N_3047,N_2646,N_2059);
xor U3048 (N_3048,N_2250,N_2163);
nand U3049 (N_3049,N_2808,N_2072);
or U3050 (N_3050,N_2898,N_2719);
nand U3051 (N_3051,N_2882,N_2558);
nor U3052 (N_3052,N_2492,N_2801);
and U3053 (N_3053,N_2935,N_2493);
nor U3054 (N_3054,N_2796,N_2124);
nand U3055 (N_3055,N_2647,N_2840);
or U3056 (N_3056,N_2044,N_2703);
or U3057 (N_3057,N_2303,N_2299);
and U3058 (N_3058,N_2574,N_2976);
nand U3059 (N_3059,N_2799,N_2745);
nor U3060 (N_3060,N_2448,N_2358);
and U3061 (N_3061,N_2055,N_2593);
xnor U3062 (N_3062,N_2999,N_2816);
or U3063 (N_3063,N_2051,N_2139);
nor U3064 (N_3064,N_2724,N_2313);
and U3065 (N_3065,N_2771,N_2528);
nor U3066 (N_3066,N_2982,N_2611);
and U3067 (N_3067,N_2482,N_2245);
and U3068 (N_3068,N_2881,N_2052);
xnor U3069 (N_3069,N_2442,N_2374);
or U3070 (N_3070,N_2886,N_2354);
and U3071 (N_3071,N_2952,N_2663);
nor U3072 (N_3072,N_2913,N_2613);
or U3073 (N_3073,N_2000,N_2965);
nand U3074 (N_3074,N_2242,N_2909);
or U3075 (N_3075,N_2867,N_2930);
and U3076 (N_3076,N_2921,N_2670);
nand U3077 (N_3077,N_2093,N_2363);
and U3078 (N_3078,N_2225,N_2054);
nand U3079 (N_3079,N_2252,N_2845);
or U3080 (N_3080,N_2217,N_2415);
xor U3081 (N_3081,N_2606,N_2873);
and U3082 (N_3082,N_2317,N_2770);
nand U3083 (N_3083,N_2399,N_2428);
xor U3084 (N_3084,N_2787,N_2226);
or U3085 (N_3085,N_2362,N_2089);
nor U3086 (N_3086,N_2948,N_2280);
xor U3087 (N_3087,N_2877,N_2879);
or U3088 (N_3088,N_2080,N_2540);
xnor U3089 (N_3089,N_2931,N_2082);
nand U3090 (N_3090,N_2255,N_2383);
xnor U3091 (N_3091,N_2885,N_2452);
and U3092 (N_3092,N_2686,N_2656);
nand U3093 (N_3093,N_2516,N_2731);
nor U3094 (N_3094,N_2016,N_2809);
nand U3095 (N_3095,N_2424,N_2167);
xnor U3096 (N_3096,N_2607,N_2194);
nor U3097 (N_3097,N_2699,N_2640);
and U3098 (N_3098,N_2147,N_2746);
xnor U3099 (N_3099,N_2570,N_2259);
or U3100 (N_3100,N_2783,N_2142);
nand U3101 (N_3101,N_2664,N_2599);
nor U3102 (N_3102,N_2659,N_2324);
nand U3103 (N_3103,N_2715,N_2043);
nand U3104 (N_3104,N_2738,N_2916);
xor U3105 (N_3105,N_2712,N_2618);
xor U3106 (N_3106,N_2073,N_2185);
or U3107 (N_3107,N_2002,N_2907);
nand U3108 (N_3108,N_2705,N_2509);
nor U3109 (N_3109,N_2231,N_2047);
nand U3110 (N_3110,N_2495,N_2995);
nor U3111 (N_3111,N_2768,N_2100);
and U3112 (N_3112,N_2469,N_2347);
xor U3113 (N_3113,N_2458,N_2828);
nand U3114 (N_3114,N_2017,N_2224);
nor U3115 (N_3115,N_2876,N_2944);
or U3116 (N_3116,N_2678,N_2690);
nor U3117 (N_3117,N_2695,N_2106);
nand U3118 (N_3118,N_2108,N_2330);
nand U3119 (N_3119,N_2849,N_2214);
or U3120 (N_3120,N_2189,N_2865);
xor U3121 (N_3121,N_2370,N_2402);
xor U3122 (N_3122,N_2432,N_2583);
xnor U3123 (N_3123,N_2282,N_2569);
nor U3124 (N_3124,N_2869,N_2232);
nor U3125 (N_3125,N_2956,N_2466);
or U3126 (N_3126,N_2933,N_2007);
xor U3127 (N_3127,N_2416,N_2166);
nand U3128 (N_3128,N_2531,N_2425);
and U3129 (N_3129,N_2698,N_2037);
or U3130 (N_3130,N_2134,N_2961);
and U3131 (N_3131,N_2254,N_2474);
and U3132 (N_3132,N_2892,N_2187);
xor U3133 (N_3133,N_2763,N_2639);
nor U3134 (N_3134,N_2554,N_2862);
xor U3135 (N_3135,N_2891,N_2049);
nand U3136 (N_3136,N_2220,N_2465);
xor U3137 (N_3137,N_2628,N_2257);
nor U3138 (N_3138,N_2863,N_2970);
and U3139 (N_3139,N_2261,N_2696);
or U3140 (N_3140,N_2480,N_2152);
xnor U3141 (N_3141,N_2494,N_2623);
or U3142 (N_3142,N_2234,N_2260);
xnor U3143 (N_3143,N_2932,N_2154);
nor U3144 (N_3144,N_2456,N_2518);
nor U3145 (N_3145,N_2526,N_2927);
nand U3146 (N_3146,N_2923,N_2366);
xnor U3147 (N_3147,N_2473,N_2757);
or U3148 (N_3148,N_2446,N_2308);
nor U3149 (N_3149,N_2258,N_2727);
nand U3150 (N_3150,N_2819,N_2972);
and U3151 (N_3151,N_2451,N_2295);
xor U3152 (N_3152,N_2716,N_2195);
or U3153 (N_3153,N_2585,N_2589);
nor U3154 (N_3154,N_2729,N_2042);
nor U3155 (N_3155,N_2463,N_2331);
nor U3156 (N_3156,N_2726,N_2692);
and U3157 (N_3157,N_2550,N_2394);
and U3158 (N_3158,N_2760,N_2011);
nand U3159 (N_3159,N_2521,N_2061);
xnor U3160 (N_3160,N_2103,N_2813);
nor U3161 (N_3161,N_2119,N_2019);
or U3162 (N_3162,N_2924,N_2708);
nor U3163 (N_3163,N_2155,N_2203);
or U3164 (N_3164,N_2437,N_2732);
xor U3165 (N_3165,N_2901,N_2632);
or U3166 (N_3166,N_2311,N_2851);
xnor U3167 (N_3167,N_2918,N_2365);
xor U3168 (N_3168,N_2169,N_2319);
nor U3169 (N_3169,N_2960,N_2198);
nor U3170 (N_3170,N_2159,N_2156);
and U3171 (N_3171,N_2063,N_2409);
or U3172 (N_3172,N_2826,N_2427);
nor U3173 (N_3173,N_2112,N_2630);
and U3174 (N_3174,N_2470,N_2223);
nand U3175 (N_3175,N_2576,N_2070);
nand U3176 (N_3176,N_2275,N_2088);
or U3177 (N_3177,N_2084,N_2627);
nand U3178 (N_3178,N_2202,N_2298);
nor U3179 (N_3179,N_2580,N_2648);
nand U3180 (N_3180,N_2689,N_2859);
xnor U3181 (N_3181,N_2003,N_2071);
nor U3182 (N_3182,N_2751,N_2915);
or U3183 (N_3183,N_2395,N_2401);
or U3184 (N_3184,N_2889,N_2821);
and U3185 (N_3185,N_2592,N_2781);
xnor U3186 (N_3186,N_2942,N_2488);
or U3187 (N_3187,N_2609,N_2802);
xnor U3188 (N_3188,N_2186,N_2140);
nor U3189 (N_3189,N_2793,N_2233);
and U3190 (N_3190,N_2795,N_2545);
and U3191 (N_3191,N_2822,N_2404);
nor U3192 (N_3192,N_2200,N_2767);
nor U3193 (N_3193,N_2460,N_2557);
xor U3194 (N_3194,N_2449,N_2433);
or U3195 (N_3195,N_2179,N_2079);
nand U3196 (N_3196,N_2184,N_2064);
nor U3197 (N_3197,N_2515,N_2905);
or U3198 (N_3198,N_2211,N_2240);
and U3199 (N_3199,N_2814,N_2382);
xnor U3200 (N_3200,N_2341,N_2022);
and U3201 (N_3201,N_2248,N_2844);
and U3202 (N_3202,N_2508,N_2265);
and U3203 (N_3203,N_2653,N_2736);
nand U3204 (N_3204,N_2911,N_2092);
or U3205 (N_3205,N_2018,N_2511);
or U3206 (N_3206,N_2306,N_2704);
xor U3207 (N_3207,N_2925,N_2107);
or U3208 (N_3208,N_2798,N_2755);
and U3209 (N_3209,N_2153,N_2206);
and U3210 (N_3210,N_2342,N_2454);
or U3211 (N_3211,N_2024,N_2173);
and U3212 (N_3212,N_2794,N_2759);
or U3213 (N_3213,N_2786,N_2544);
or U3214 (N_3214,N_2652,N_2839);
xor U3215 (N_3215,N_2669,N_2253);
nand U3216 (N_3216,N_2464,N_2364);
nor U3217 (N_3217,N_2529,N_2920);
nand U3218 (N_3218,N_2285,N_2263);
nor U3219 (N_3219,N_2707,N_2566);
and U3220 (N_3220,N_2713,N_2984);
and U3221 (N_3221,N_2481,N_2950);
xnor U3222 (N_3222,N_2990,N_2392);
or U3223 (N_3223,N_2209,N_2949);
and U3224 (N_3224,N_2279,N_2720);
xor U3225 (N_3225,N_2262,N_2776);
or U3226 (N_3226,N_2345,N_2878);
or U3227 (N_3227,N_2122,N_2274);
xnor U3228 (N_3228,N_2894,N_2467);
and U3229 (N_3229,N_2842,N_2897);
and U3230 (N_3230,N_2722,N_2355);
nand U3231 (N_3231,N_2453,N_2989);
nor U3232 (N_3232,N_2853,N_2434);
xnor U3233 (N_3233,N_2846,N_2009);
xnor U3234 (N_3234,N_2631,N_2038);
nand U3235 (N_3235,N_2617,N_2413);
nor U3236 (N_3236,N_2957,N_2969);
and U3237 (N_3237,N_2532,N_2864);
xnor U3238 (N_3238,N_2711,N_2182);
nor U3239 (N_3239,N_2396,N_2036);
and U3240 (N_3240,N_2098,N_2605);
or U3241 (N_3241,N_2318,N_2053);
or U3242 (N_3242,N_2553,N_2241);
nor U3243 (N_3243,N_2700,N_2329);
nor U3244 (N_3244,N_2291,N_2387);
nor U3245 (N_3245,N_2006,N_2549);
and U3246 (N_3246,N_2993,N_2688);
and U3247 (N_3247,N_2848,N_2572);
nor U3248 (N_3248,N_2951,N_2222);
nand U3249 (N_3249,N_2149,N_2444);
nor U3250 (N_3250,N_2028,N_2183);
and U3251 (N_3251,N_2065,N_2980);
nor U3252 (N_3252,N_2504,N_2158);
nand U3253 (N_3253,N_2739,N_2293);
nand U3254 (N_3254,N_2872,N_2806);
nand U3255 (N_3255,N_2403,N_2490);
xnor U3256 (N_3256,N_2136,N_2774);
and U3257 (N_3257,N_2375,N_2199);
nor U3258 (N_3258,N_2861,N_2013);
or U3259 (N_3259,N_2349,N_2676);
and U3260 (N_3260,N_2097,N_2421);
xor U3261 (N_3261,N_2369,N_2067);
nand U3262 (N_3262,N_2843,N_2479);
xnor U3263 (N_3263,N_2357,N_2955);
xnor U3264 (N_3264,N_2164,N_2272);
or U3265 (N_3265,N_2780,N_2741);
xor U3266 (N_3266,N_2835,N_2568);
or U3267 (N_3267,N_2327,N_2050);
nand U3268 (N_3268,N_2314,N_2650);
or U3269 (N_3269,N_2236,N_2247);
and U3270 (N_3270,N_2393,N_2866);
and U3271 (N_3271,N_2600,N_2977);
and U3272 (N_3272,N_2309,N_2388);
xnor U3273 (N_3273,N_2975,N_2027);
or U3274 (N_3274,N_2679,N_2397);
and U3275 (N_3275,N_2895,N_2517);
and U3276 (N_3276,N_2538,N_2773);
nor U3277 (N_3277,N_2858,N_2129);
nor U3278 (N_3278,N_2709,N_2418);
nor U3279 (N_3279,N_2376,N_2908);
nor U3280 (N_3280,N_2343,N_2384);
or U3281 (N_3281,N_2207,N_2323);
nand U3282 (N_3282,N_2963,N_2477);
nand U3283 (N_3283,N_2212,N_2443);
xnor U3284 (N_3284,N_2694,N_2276);
nand U3285 (N_3285,N_2968,N_2333);
nand U3286 (N_3286,N_2616,N_2350);
nor U3287 (N_3287,N_2032,N_2888);
nand U3288 (N_3288,N_2438,N_2334);
nor U3289 (N_3289,N_2902,N_2304);
nor U3290 (N_3290,N_2829,N_2069);
and U3291 (N_3291,N_2497,N_2943);
or U3292 (N_3292,N_2292,N_2561);
and U3293 (N_3293,N_2348,N_2520);
nor U3294 (N_3294,N_2143,N_2578);
nand U3295 (N_3295,N_2560,N_2312);
and U3296 (N_3296,N_2012,N_2266);
and U3297 (N_3297,N_2579,N_2871);
nand U3298 (N_3298,N_2461,N_2351);
nor U3299 (N_3299,N_2180,N_2827);
and U3300 (N_3300,N_2268,N_2315);
nand U3301 (N_3301,N_2868,N_2527);
or U3302 (N_3302,N_2114,N_2123);
and U3303 (N_3303,N_2803,N_2525);
or U3304 (N_3304,N_2367,N_2946);
xor U3305 (N_3305,N_2496,N_2588);
or U3306 (N_3306,N_2852,N_2487);
and U3307 (N_3307,N_2408,N_2855);
nor U3308 (N_3308,N_2812,N_2359);
and U3309 (N_3309,N_2903,N_2649);
and U3310 (N_3310,N_2216,N_2411);
xor U3311 (N_3311,N_2021,N_2168);
xnor U3312 (N_3312,N_2105,N_2655);
nor U3313 (N_3313,N_2564,N_2747);
xor U3314 (N_3314,N_2235,N_2994);
or U3315 (N_3315,N_2227,N_2800);
or U3316 (N_3316,N_2581,N_2340);
or U3317 (N_3317,N_2023,N_2109);
nor U3318 (N_3318,N_2510,N_2062);
nand U3319 (N_3319,N_2749,N_2144);
and U3320 (N_3320,N_2271,N_2026);
nand U3321 (N_3321,N_2118,N_2015);
xnor U3322 (N_3322,N_2410,N_2056);
nand U3323 (N_3323,N_2127,N_2615);
and U3324 (N_3324,N_2267,N_2457);
nand U3325 (N_3325,N_2575,N_2020);
and U3326 (N_3326,N_2281,N_2310);
or U3327 (N_3327,N_2447,N_2381);
and U3328 (N_3328,N_2440,N_2128);
or U3329 (N_3329,N_2441,N_2503);
nor U3330 (N_3330,N_2338,N_2057);
nand U3331 (N_3331,N_2468,N_2964);
nand U3332 (N_3332,N_2644,N_2133);
nor U3333 (N_3333,N_2620,N_2584);
or U3334 (N_3334,N_2941,N_2398);
or U3335 (N_3335,N_2141,N_2116);
nor U3336 (N_3336,N_2219,N_2660);
nor U3337 (N_3337,N_2256,N_2967);
xnor U3338 (N_3338,N_2718,N_2577);
nand U3339 (N_3339,N_2626,N_2445);
or U3340 (N_3340,N_2937,N_2728);
or U3341 (N_3341,N_2546,N_2847);
nand U3342 (N_3342,N_2326,N_2754);
and U3343 (N_3343,N_2475,N_2177);
and U3344 (N_3344,N_2748,N_2066);
and U3345 (N_3345,N_2597,N_2706);
xor U3346 (N_3346,N_2778,N_2973);
and U3347 (N_3347,N_2998,N_2307);
xor U3348 (N_3348,N_2671,N_2621);
or U3349 (N_3349,N_2603,N_2856);
xnor U3350 (N_3350,N_2204,N_2172);
and U3351 (N_3351,N_2752,N_2353);
nor U3352 (N_3352,N_2215,N_2406);
xor U3353 (N_3353,N_2522,N_2077);
xnor U3354 (N_3354,N_2836,N_2666);
nand U3355 (N_3355,N_2832,N_2148);
nor U3356 (N_3356,N_2818,N_2904);
nor U3357 (N_3357,N_2094,N_2210);
nand U3358 (N_3358,N_2004,N_2880);
xnor U3359 (N_3359,N_2657,N_2784);
nor U3360 (N_3360,N_2201,N_2910);
and U3361 (N_3361,N_2791,N_2817);
nor U3362 (N_3362,N_2294,N_2837);
nand U3363 (N_3363,N_2111,N_2587);
xnor U3364 (N_3364,N_2126,N_2151);
and U3365 (N_3365,N_2668,N_2192);
nor U3366 (N_3366,N_2188,N_2547);
nor U3367 (N_3367,N_2368,N_2068);
and U3368 (N_3368,N_2769,N_2277);
xnor U3369 (N_3369,N_2419,N_2246);
and U3370 (N_3370,N_2654,N_2332);
and U3371 (N_3371,N_2228,N_2860);
nand U3372 (N_3372,N_2811,N_2693);
nand U3373 (N_3373,N_2622,N_2076);
nor U3374 (N_3374,N_2273,N_2883);
nand U3375 (N_3375,N_2758,N_2104);
nor U3376 (N_3376,N_2717,N_2157);
nand U3377 (N_3377,N_2743,N_2571);
or U3378 (N_3378,N_2590,N_2966);
nand U3379 (N_3379,N_2264,N_2237);
nand U3380 (N_3380,N_2251,N_2125);
nand U3381 (N_3381,N_2635,N_2740);
nor U3382 (N_3382,N_2506,N_2336);
nor U3383 (N_3383,N_2988,N_2095);
and U3384 (N_3384,N_2854,N_2765);
xor U3385 (N_3385,N_2096,N_2379);
nand U3386 (N_3386,N_2120,N_2431);
or U3387 (N_3387,N_2344,N_2672);
and U3388 (N_3388,N_2060,N_2029);
nor U3389 (N_3389,N_2629,N_2025);
xnor U3390 (N_3390,N_2078,N_2906);
and U3391 (N_3391,N_2483,N_2685);
and U3392 (N_3392,N_2673,N_2624);
nand U3393 (N_3393,N_2459,N_2591);
xnor U3394 (N_3394,N_2598,N_2083);
and U3395 (N_3395,N_2750,N_2884);
nor U3396 (N_3396,N_2900,N_2288);
nand U3397 (N_3397,N_2684,N_2914);
nor U3398 (N_3398,N_2360,N_2238);
nand U3399 (N_3399,N_2131,N_2178);
and U3400 (N_3400,N_2667,N_2471);
xor U3401 (N_3401,N_2556,N_2283);
xnor U3402 (N_3402,N_2761,N_2825);
or U3403 (N_3403,N_2834,N_2619);
or U3404 (N_3404,N_2734,N_2820);
and U3405 (N_3405,N_2987,N_2661);
xnor U3406 (N_3406,N_2823,N_2643);
or U3407 (N_3407,N_2833,N_2875);
or U3408 (N_3408,N_2562,N_2810);
nor U3409 (N_3409,N_2356,N_2919);
nor U3410 (N_3410,N_2683,N_2958);
or U3411 (N_3411,N_2423,N_2328);
nor U3412 (N_3412,N_2633,N_2174);
or U3413 (N_3413,N_2218,N_2772);
nor U3414 (N_3414,N_2378,N_2542);
nor U3415 (N_3415,N_2371,N_2582);
nand U3416 (N_3416,N_2565,N_2420);
xnor U3417 (N_3417,N_2320,N_2305);
nand U3418 (N_3418,N_2400,N_2874);
and U3419 (N_3419,N_2372,N_2831);
and U3420 (N_3420,N_2113,N_2239);
and U3421 (N_3421,N_2586,N_2680);
xor U3422 (N_3422,N_2014,N_2645);
or U3423 (N_3423,N_2039,N_2986);
xnor U3424 (N_3424,N_2213,N_2928);
and U3425 (N_3425,N_2507,N_2091);
and U3426 (N_3426,N_2335,N_2175);
and U3427 (N_3427,N_2934,N_2735);
and U3428 (N_3428,N_2940,N_2499);
nand U3429 (N_3429,N_2391,N_2830);
nand U3430 (N_3430,N_2476,N_2797);
or U3431 (N_3431,N_2612,N_2595);
nor U3432 (N_3432,N_2548,N_2917);
nand U3433 (N_3433,N_2414,N_2979);
xnor U3434 (N_3434,N_2450,N_2788);
nor U3435 (N_3435,N_2922,N_2702);
or U3436 (N_3436,N_2701,N_2390);
or U3437 (N_3437,N_2559,N_2539);
and U3438 (N_3438,N_2710,N_2725);
or U3439 (N_3439,N_2302,N_2983);
or U3440 (N_3440,N_2804,N_2489);
nor U3441 (N_3441,N_2484,N_2636);
nand U3442 (N_3442,N_2296,N_2455);
xnor U3443 (N_3443,N_2610,N_2608);
and U3444 (N_3444,N_2138,N_2697);
xor U3445 (N_3445,N_2792,N_2805);
nand U3446 (N_3446,N_2737,N_2270);
nand U3447 (N_3447,N_2779,N_2045);
xor U3448 (N_3448,N_2785,N_2491);
or U3449 (N_3449,N_2721,N_2316);
or U3450 (N_3450,N_2034,N_2782);
and U3451 (N_3451,N_2422,N_2150);
nand U3452 (N_3452,N_2638,N_2085);
xnor U3453 (N_3453,N_2130,N_2346);
or U3454 (N_3454,N_2841,N_2658);
xor U3455 (N_3455,N_2221,N_2744);
and U3456 (N_3456,N_2601,N_2775);
or U3457 (N_3457,N_2947,N_2286);
nand U3458 (N_3458,N_2352,N_2981);
nand U3459 (N_3459,N_2462,N_2321);
or U3460 (N_3460,N_2289,N_2048);
nand U3461 (N_3461,N_2325,N_2269);
or U3462 (N_3462,N_2075,N_2373);
and U3463 (N_3463,N_2929,N_2541);
and U3464 (N_3464,N_2322,N_2031);
or U3465 (N_3465,N_2939,N_2176);
nand U3466 (N_3466,N_2191,N_2674);
or U3467 (N_3467,N_2498,N_2896);
nor U3468 (N_3468,N_2893,N_2380);
nand U3469 (N_3469,N_2385,N_2642);
nor U3470 (N_3470,N_2567,N_2135);
xnor U3471 (N_3471,N_2439,N_2500);
nand U3472 (N_3472,N_2625,N_2386);
or U3473 (N_3473,N_2838,N_2190);
xnor U3474 (N_3474,N_2912,N_2807);
xnor U3475 (N_3475,N_2978,N_2985);
and U3476 (N_3476,N_2899,N_2074);
nor U3477 (N_3477,N_2594,N_2417);
and U3478 (N_3478,N_2472,N_2435);
xor U3479 (N_3479,N_2430,N_2533);
and U3480 (N_3480,N_2604,N_2243);
nand U3481 (N_3481,N_2824,N_2389);
or U3482 (N_3482,N_2665,N_2407);
xor U3483 (N_3483,N_2081,N_2086);
xor U3484 (N_3484,N_2278,N_2870);
or U3485 (N_3485,N_2099,N_2008);
and U3486 (N_3486,N_2953,N_2502);
nand U3487 (N_3487,N_2945,N_2030);
or U3488 (N_3488,N_2287,N_2090);
nand U3489 (N_3489,N_2010,N_2637);
nor U3490 (N_3490,N_2405,N_2850);
and U3491 (N_3491,N_2196,N_2040);
nand U3492 (N_3492,N_2742,N_2208);
and U3493 (N_3493,N_2730,N_2687);
xnor U3494 (N_3494,N_2102,N_2766);
and U3495 (N_3495,N_2535,N_2926);
or U3496 (N_3496,N_2145,N_2171);
xnor U3497 (N_3497,N_2501,N_2436);
xnor U3498 (N_3498,N_2205,N_2486);
and U3499 (N_3499,N_2035,N_2301);
nor U3500 (N_3500,N_2874,N_2404);
xor U3501 (N_3501,N_2310,N_2131);
or U3502 (N_3502,N_2345,N_2374);
nand U3503 (N_3503,N_2645,N_2492);
nor U3504 (N_3504,N_2657,N_2330);
xnor U3505 (N_3505,N_2225,N_2897);
nand U3506 (N_3506,N_2026,N_2549);
xor U3507 (N_3507,N_2657,N_2529);
or U3508 (N_3508,N_2996,N_2602);
nor U3509 (N_3509,N_2375,N_2275);
nor U3510 (N_3510,N_2877,N_2687);
nor U3511 (N_3511,N_2608,N_2223);
and U3512 (N_3512,N_2496,N_2481);
nand U3513 (N_3513,N_2079,N_2925);
nor U3514 (N_3514,N_2166,N_2916);
nand U3515 (N_3515,N_2848,N_2282);
nand U3516 (N_3516,N_2781,N_2364);
nand U3517 (N_3517,N_2272,N_2843);
and U3518 (N_3518,N_2300,N_2809);
xnor U3519 (N_3519,N_2956,N_2593);
xor U3520 (N_3520,N_2448,N_2991);
or U3521 (N_3521,N_2864,N_2670);
nand U3522 (N_3522,N_2625,N_2280);
xor U3523 (N_3523,N_2765,N_2617);
or U3524 (N_3524,N_2214,N_2574);
or U3525 (N_3525,N_2359,N_2002);
and U3526 (N_3526,N_2153,N_2745);
and U3527 (N_3527,N_2109,N_2999);
or U3528 (N_3528,N_2838,N_2166);
xor U3529 (N_3529,N_2970,N_2983);
and U3530 (N_3530,N_2225,N_2195);
and U3531 (N_3531,N_2446,N_2361);
nand U3532 (N_3532,N_2266,N_2969);
xnor U3533 (N_3533,N_2128,N_2692);
xor U3534 (N_3534,N_2525,N_2410);
nand U3535 (N_3535,N_2851,N_2569);
nor U3536 (N_3536,N_2872,N_2743);
xor U3537 (N_3537,N_2039,N_2558);
and U3538 (N_3538,N_2619,N_2481);
xor U3539 (N_3539,N_2237,N_2700);
or U3540 (N_3540,N_2865,N_2664);
or U3541 (N_3541,N_2337,N_2380);
nor U3542 (N_3542,N_2356,N_2637);
xnor U3543 (N_3543,N_2676,N_2022);
or U3544 (N_3544,N_2299,N_2106);
or U3545 (N_3545,N_2328,N_2931);
and U3546 (N_3546,N_2899,N_2668);
xor U3547 (N_3547,N_2587,N_2642);
xnor U3548 (N_3548,N_2556,N_2290);
xnor U3549 (N_3549,N_2629,N_2612);
nor U3550 (N_3550,N_2910,N_2378);
nor U3551 (N_3551,N_2026,N_2471);
nand U3552 (N_3552,N_2610,N_2064);
nand U3553 (N_3553,N_2322,N_2773);
nand U3554 (N_3554,N_2727,N_2245);
nand U3555 (N_3555,N_2333,N_2450);
xor U3556 (N_3556,N_2919,N_2585);
nor U3557 (N_3557,N_2369,N_2549);
nor U3558 (N_3558,N_2898,N_2954);
nand U3559 (N_3559,N_2336,N_2848);
nor U3560 (N_3560,N_2335,N_2678);
nand U3561 (N_3561,N_2382,N_2223);
and U3562 (N_3562,N_2376,N_2202);
xor U3563 (N_3563,N_2841,N_2952);
nand U3564 (N_3564,N_2588,N_2525);
or U3565 (N_3565,N_2979,N_2365);
nor U3566 (N_3566,N_2294,N_2193);
or U3567 (N_3567,N_2620,N_2485);
and U3568 (N_3568,N_2599,N_2433);
or U3569 (N_3569,N_2172,N_2438);
nand U3570 (N_3570,N_2346,N_2679);
nor U3571 (N_3571,N_2695,N_2670);
and U3572 (N_3572,N_2527,N_2605);
and U3573 (N_3573,N_2330,N_2696);
or U3574 (N_3574,N_2027,N_2277);
and U3575 (N_3575,N_2083,N_2525);
nor U3576 (N_3576,N_2847,N_2942);
xnor U3577 (N_3577,N_2203,N_2065);
or U3578 (N_3578,N_2652,N_2437);
or U3579 (N_3579,N_2117,N_2550);
and U3580 (N_3580,N_2308,N_2312);
or U3581 (N_3581,N_2834,N_2541);
or U3582 (N_3582,N_2146,N_2125);
or U3583 (N_3583,N_2064,N_2792);
xor U3584 (N_3584,N_2685,N_2111);
and U3585 (N_3585,N_2694,N_2217);
and U3586 (N_3586,N_2204,N_2637);
xnor U3587 (N_3587,N_2889,N_2729);
or U3588 (N_3588,N_2033,N_2988);
nor U3589 (N_3589,N_2813,N_2361);
and U3590 (N_3590,N_2316,N_2455);
or U3591 (N_3591,N_2089,N_2609);
and U3592 (N_3592,N_2548,N_2039);
nor U3593 (N_3593,N_2012,N_2516);
or U3594 (N_3594,N_2798,N_2760);
nand U3595 (N_3595,N_2703,N_2944);
or U3596 (N_3596,N_2241,N_2503);
nand U3597 (N_3597,N_2504,N_2313);
nand U3598 (N_3598,N_2757,N_2414);
nor U3599 (N_3599,N_2005,N_2054);
nor U3600 (N_3600,N_2901,N_2797);
xor U3601 (N_3601,N_2915,N_2753);
xor U3602 (N_3602,N_2629,N_2258);
and U3603 (N_3603,N_2720,N_2073);
nor U3604 (N_3604,N_2291,N_2377);
xnor U3605 (N_3605,N_2756,N_2767);
nor U3606 (N_3606,N_2152,N_2727);
xor U3607 (N_3607,N_2605,N_2266);
xnor U3608 (N_3608,N_2991,N_2014);
or U3609 (N_3609,N_2734,N_2201);
nor U3610 (N_3610,N_2178,N_2924);
or U3611 (N_3611,N_2750,N_2793);
nand U3612 (N_3612,N_2010,N_2162);
nor U3613 (N_3613,N_2173,N_2950);
nand U3614 (N_3614,N_2707,N_2894);
or U3615 (N_3615,N_2567,N_2694);
or U3616 (N_3616,N_2362,N_2779);
and U3617 (N_3617,N_2594,N_2965);
nand U3618 (N_3618,N_2295,N_2299);
nand U3619 (N_3619,N_2906,N_2969);
nand U3620 (N_3620,N_2532,N_2747);
xor U3621 (N_3621,N_2514,N_2289);
or U3622 (N_3622,N_2297,N_2984);
and U3623 (N_3623,N_2959,N_2513);
and U3624 (N_3624,N_2311,N_2588);
or U3625 (N_3625,N_2886,N_2372);
nand U3626 (N_3626,N_2179,N_2823);
or U3627 (N_3627,N_2222,N_2914);
nand U3628 (N_3628,N_2001,N_2758);
nand U3629 (N_3629,N_2767,N_2191);
and U3630 (N_3630,N_2673,N_2060);
nand U3631 (N_3631,N_2139,N_2684);
nor U3632 (N_3632,N_2252,N_2916);
or U3633 (N_3633,N_2733,N_2426);
nand U3634 (N_3634,N_2714,N_2065);
or U3635 (N_3635,N_2127,N_2041);
nand U3636 (N_3636,N_2621,N_2711);
xnor U3637 (N_3637,N_2903,N_2050);
xor U3638 (N_3638,N_2776,N_2117);
nor U3639 (N_3639,N_2517,N_2738);
nor U3640 (N_3640,N_2296,N_2597);
or U3641 (N_3641,N_2887,N_2924);
xor U3642 (N_3642,N_2200,N_2288);
nand U3643 (N_3643,N_2163,N_2838);
or U3644 (N_3644,N_2893,N_2515);
nand U3645 (N_3645,N_2237,N_2318);
and U3646 (N_3646,N_2741,N_2085);
nor U3647 (N_3647,N_2676,N_2443);
or U3648 (N_3648,N_2186,N_2846);
or U3649 (N_3649,N_2075,N_2543);
nand U3650 (N_3650,N_2460,N_2882);
xor U3651 (N_3651,N_2194,N_2722);
nand U3652 (N_3652,N_2434,N_2165);
xnor U3653 (N_3653,N_2790,N_2385);
or U3654 (N_3654,N_2972,N_2853);
xnor U3655 (N_3655,N_2275,N_2877);
and U3656 (N_3656,N_2059,N_2220);
nand U3657 (N_3657,N_2231,N_2227);
xor U3658 (N_3658,N_2084,N_2568);
nor U3659 (N_3659,N_2231,N_2761);
nand U3660 (N_3660,N_2405,N_2699);
xor U3661 (N_3661,N_2576,N_2079);
or U3662 (N_3662,N_2977,N_2720);
or U3663 (N_3663,N_2591,N_2311);
xnor U3664 (N_3664,N_2396,N_2357);
nand U3665 (N_3665,N_2794,N_2508);
and U3666 (N_3666,N_2450,N_2569);
xor U3667 (N_3667,N_2110,N_2712);
xor U3668 (N_3668,N_2156,N_2495);
xor U3669 (N_3669,N_2100,N_2905);
and U3670 (N_3670,N_2932,N_2772);
xnor U3671 (N_3671,N_2462,N_2055);
or U3672 (N_3672,N_2038,N_2211);
nand U3673 (N_3673,N_2089,N_2955);
or U3674 (N_3674,N_2634,N_2594);
xor U3675 (N_3675,N_2545,N_2533);
nand U3676 (N_3676,N_2695,N_2270);
nor U3677 (N_3677,N_2642,N_2927);
and U3678 (N_3678,N_2457,N_2894);
or U3679 (N_3679,N_2610,N_2441);
and U3680 (N_3680,N_2429,N_2764);
xnor U3681 (N_3681,N_2698,N_2182);
or U3682 (N_3682,N_2064,N_2824);
nor U3683 (N_3683,N_2556,N_2903);
nand U3684 (N_3684,N_2209,N_2050);
xor U3685 (N_3685,N_2180,N_2350);
or U3686 (N_3686,N_2421,N_2558);
nand U3687 (N_3687,N_2727,N_2846);
xnor U3688 (N_3688,N_2363,N_2258);
nor U3689 (N_3689,N_2693,N_2915);
and U3690 (N_3690,N_2467,N_2947);
and U3691 (N_3691,N_2513,N_2654);
xnor U3692 (N_3692,N_2338,N_2517);
or U3693 (N_3693,N_2666,N_2351);
xor U3694 (N_3694,N_2003,N_2530);
xnor U3695 (N_3695,N_2258,N_2202);
or U3696 (N_3696,N_2266,N_2022);
nand U3697 (N_3697,N_2199,N_2861);
or U3698 (N_3698,N_2287,N_2222);
nand U3699 (N_3699,N_2299,N_2792);
nor U3700 (N_3700,N_2975,N_2678);
or U3701 (N_3701,N_2645,N_2023);
xor U3702 (N_3702,N_2250,N_2728);
or U3703 (N_3703,N_2952,N_2221);
xor U3704 (N_3704,N_2578,N_2249);
xnor U3705 (N_3705,N_2808,N_2396);
xor U3706 (N_3706,N_2731,N_2701);
xor U3707 (N_3707,N_2233,N_2274);
xor U3708 (N_3708,N_2286,N_2090);
xor U3709 (N_3709,N_2193,N_2878);
nor U3710 (N_3710,N_2299,N_2437);
xor U3711 (N_3711,N_2176,N_2549);
and U3712 (N_3712,N_2008,N_2328);
nand U3713 (N_3713,N_2739,N_2231);
and U3714 (N_3714,N_2417,N_2783);
xnor U3715 (N_3715,N_2151,N_2280);
and U3716 (N_3716,N_2232,N_2123);
nand U3717 (N_3717,N_2924,N_2678);
and U3718 (N_3718,N_2941,N_2900);
xnor U3719 (N_3719,N_2275,N_2741);
nand U3720 (N_3720,N_2341,N_2640);
or U3721 (N_3721,N_2889,N_2027);
nor U3722 (N_3722,N_2479,N_2622);
nor U3723 (N_3723,N_2143,N_2861);
or U3724 (N_3724,N_2979,N_2288);
xnor U3725 (N_3725,N_2483,N_2409);
xor U3726 (N_3726,N_2020,N_2015);
nand U3727 (N_3727,N_2203,N_2834);
xor U3728 (N_3728,N_2640,N_2937);
nor U3729 (N_3729,N_2998,N_2501);
and U3730 (N_3730,N_2735,N_2162);
and U3731 (N_3731,N_2060,N_2645);
and U3732 (N_3732,N_2992,N_2667);
xnor U3733 (N_3733,N_2304,N_2162);
nand U3734 (N_3734,N_2969,N_2102);
nand U3735 (N_3735,N_2993,N_2635);
xor U3736 (N_3736,N_2152,N_2763);
nand U3737 (N_3737,N_2511,N_2644);
xor U3738 (N_3738,N_2640,N_2177);
nand U3739 (N_3739,N_2340,N_2357);
nor U3740 (N_3740,N_2157,N_2078);
and U3741 (N_3741,N_2869,N_2268);
nor U3742 (N_3742,N_2103,N_2078);
or U3743 (N_3743,N_2098,N_2548);
nand U3744 (N_3744,N_2673,N_2236);
or U3745 (N_3745,N_2740,N_2820);
xor U3746 (N_3746,N_2827,N_2828);
or U3747 (N_3747,N_2764,N_2326);
xnor U3748 (N_3748,N_2643,N_2083);
and U3749 (N_3749,N_2242,N_2984);
or U3750 (N_3750,N_2019,N_2577);
or U3751 (N_3751,N_2083,N_2499);
nand U3752 (N_3752,N_2941,N_2685);
or U3753 (N_3753,N_2679,N_2112);
nand U3754 (N_3754,N_2488,N_2504);
or U3755 (N_3755,N_2326,N_2750);
xnor U3756 (N_3756,N_2530,N_2769);
nand U3757 (N_3757,N_2066,N_2623);
and U3758 (N_3758,N_2686,N_2099);
nor U3759 (N_3759,N_2207,N_2257);
nor U3760 (N_3760,N_2597,N_2343);
xor U3761 (N_3761,N_2924,N_2015);
and U3762 (N_3762,N_2179,N_2528);
or U3763 (N_3763,N_2696,N_2258);
nor U3764 (N_3764,N_2981,N_2297);
or U3765 (N_3765,N_2216,N_2705);
and U3766 (N_3766,N_2099,N_2751);
nand U3767 (N_3767,N_2889,N_2575);
nor U3768 (N_3768,N_2033,N_2818);
and U3769 (N_3769,N_2724,N_2872);
and U3770 (N_3770,N_2133,N_2730);
or U3771 (N_3771,N_2982,N_2056);
and U3772 (N_3772,N_2785,N_2081);
xor U3773 (N_3773,N_2386,N_2966);
nor U3774 (N_3774,N_2729,N_2489);
nor U3775 (N_3775,N_2591,N_2738);
and U3776 (N_3776,N_2957,N_2853);
xor U3777 (N_3777,N_2307,N_2526);
xor U3778 (N_3778,N_2189,N_2891);
or U3779 (N_3779,N_2912,N_2355);
and U3780 (N_3780,N_2966,N_2417);
xor U3781 (N_3781,N_2416,N_2834);
and U3782 (N_3782,N_2295,N_2945);
and U3783 (N_3783,N_2791,N_2122);
nor U3784 (N_3784,N_2991,N_2108);
and U3785 (N_3785,N_2803,N_2674);
xnor U3786 (N_3786,N_2421,N_2584);
nand U3787 (N_3787,N_2927,N_2616);
xnor U3788 (N_3788,N_2306,N_2648);
nor U3789 (N_3789,N_2228,N_2837);
nand U3790 (N_3790,N_2303,N_2143);
and U3791 (N_3791,N_2488,N_2429);
nand U3792 (N_3792,N_2749,N_2492);
xor U3793 (N_3793,N_2830,N_2577);
and U3794 (N_3794,N_2857,N_2499);
xor U3795 (N_3795,N_2144,N_2185);
and U3796 (N_3796,N_2421,N_2928);
nand U3797 (N_3797,N_2544,N_2564);
and U3798 (N_3798,N_2194,N_2410);
xor U3799 (N_3799,N_2593,N_2676);
nand U3800 (N_3800,N_2765,N_2129);
xnor U3801 (N_3801,N_2894,N_2061);
and U3802 (N_3802,N_2479,N_2602);
nand U3803 (N_3803,N_2295,N_2139);
xor U3804 (N_3804,N_2285,N_2372);
xor U3805 (N_3805,N_2537,N_2663);
and U3806 (N_3806,N_2805,N_2963);
nand U3807 (N_3807,N_2946,N_2536);
or U3808 (N_3808,N_2531,N_2056);
and U3809 (N_3809,N_2558,N_2048);
or U3810 (N_3810,N_2790,N_2500);
xnor U3811 (N_3811,N_2734,N_2542);
and U3812 (N_3812,N_2176,N_2644);
xor U3813 (N_3813,N_2506,N_2335);
nand U3814 (N_3814,N_2779,N_2533);
and U3815 (N_3815,N_2662,N_2683);
nor U3816 (N_3816,N_2088,N_2204);
nand U3817 (N_3817,N_2798,N_2990);
and U3818 (N_3818,N_2404,N_2397);
or U3819 (N_3819,N_2126,N_2697);
xor U3820 (N_3820,N_2815,N_2169);
nand U3821 (N_3821,N_2217,N_2789);
nor U3822 (N_3822,N_2162,N_2235);
nor U3823 (N_3823,N_2292,N_2151);
or U3824 (N_3824,N_2607,N_2316);
xor U3825 (N_3825,N_2433,N_2542);
xor U3826 (N_3826,N_2243,N_2491);
nor U3827 (N_3827,N_2193,N_2195);
nand U3828 (N_3828,N_2422,N_2426);
nand U3829 (N_3829,N_2560,N_2080);
xnor U3830 (N_3830,N_2602,N_2537);
xnor U3831 (N_3831,N_2458,N_2736);
nand U3832 (N_3832,N_2422,N_2372);
or U3833 (N_3833,N_2524,N_2517);
and U3834 (N_3834,N_2776,N_2964);
nor U3835 (N_3835,N_2934,N_2571);
nor U3836 (N_3836,N_2606,N_2359);
xor U3837 (N_3837,N_2854,N_2789);
xor U3838 (N_3838,N_2546,N_2632);
nor U3839 (N_3839,N_2061,N_2741);
xor U3840 (N_3840,N_2597,N_2377);
or U3841 (N_3841,N_2017,N_2963);
xnor U3842 (N_3842,N_2764,N_2847);
nand U3843 (N_3843,N_2107,N_2418);
nand U3844 (N_3844,N_2587,N_2004);
and U3845 (N_3845,N_2209,N_2607);
and U3846 (N_3846,N_2138,N_2629);
xor U3847 (N_3847,N_2531,N_2215);
nand U3848 (N_3848,N_2002,N_2331);
and U3849 (N_3849,N_2576,N_2141);
xnor U3850 (N_3850,N_2479,N_2024);
nand U3851 (N_3851,N_2316,N_2098);
or U3852 (N_3852,N_2739,N_2540);
nor U3853 (N_3853,N_2440,N_2052);
nor U3854 (N_3854,N_2572,N_2543);
and U3855 (N_3855,N_2480,N_2271);
and U3856 (N_3856,N_2300,N_2162);
and U3857 (N_3857,N_2143,N_2382);
nor U3858 (N_3858,N_2733,N_2623);
and U3859 (N_3859,N_2758,N_2009);
and U3860 (N_3860,N_2997,N_2571);
nand U3861 (N_3861,N_2625,N_2219);
nand U3862 (N_3862,N_2022,N_2739);
nand U3863 (N_3863,N_2422,N_2240);
and U3864 (N_3864,N_2739,N_2294);
nand U3865 (N_3865,N_2540,N_2055);
nor U3866 (N_3866,N_2351,N_2368);
nand U3867 (N_3867,N_2836,N_2572);
nand U3868 (N_3868,N_2938,N_2446);
xnor U3869 (N_3869,N_2896,N_2953);
nor U3870 (N_3870,N_2835,N_2942);
and U3871 (N_3871,N_2496,N_2417);
nand U3872 (N_3872,N_2780,N_2281);
xnor U3873 (N_3873,N_2242,N_2966);
and U3874 (N_3874,N_2025,N_2925);
xor U3875 (N_3875,N_2789,N_2388);
xor U3876 (N_3876,N_2351,N_2981);
xor U3877 (N_3877,N_2872,N_2225);
or U3878 (N_3878,N_2844,N_2204);
nor U3879 (N_3879,N_2424,N_2263);
xnor U3880 (N_3880,N_2528,N_2992);
or U3881 (N_3881,N_2562,N_2077);
nand U3882 (N_3882,N_2469,N_2431);
nor U3883 (N_3883,N_2610,N_2747);
or U3884 (N_3884,N_2567,N_2728);
nand U3885 (N_3885,N_2076,N_2047);
nor U3886 (N_3886,N_2514,N_2883);
and U3887 (N_3887,N_2369,N_2766);
nor U3888 (N_3888,N_2336,N_2603);
nor U3889 (N_3889,N_2173,N_2050);
nor U3890 (N_3890,N_2468,N_2503);
and U3891 (N_3891,N_2058,N_2227);
and U3892 (N_3892,N_2520,N_2390);
nand U3893 (N_3893,N_2621,N_2265);
or U3894 (N_3894,N_2915,N_2118);
nand U3895 (N_3895,N_2775,N_2176);
and U3896 (N_3896,N_2307,N_2514);
or U3897 (N_3897,N_2061,N_2095);
xor U3898 (N_3898,N_2562,N_2972);
nand U3899 (N_3899,N_2269,N_2697);
or U3900 (N_3900,N_2914,N_2717);
nor U3901 (N_3901,N_2204,N_2685);
and U3902 (N_3902,N_2999,N_2241);
or U3903 (N_3903,N_2320,N_2681);
nor U3904 (N_3904,N_2906,N_2563);
nor U3905 (N_3905,N_2577,N_2223);
nand U3906 (N_3906,N_2320,N_2476);
nand U3907 (N_3907,N_2309,N_2910);
nor U3908 (N_3908,N_2947,N_2171);
xnor U3909 (N_3909,N_2461,N_2906);
xor U3910 (N_3910,N_2760,N_2140);
nor U3911 (N_3911,N_2796,N_2651);
xnor U3912 (N_3912,N_2537,N_2146);
nor U3913 (N_3913,N_2125,N_2678);
or U3914 (N_3914,N_2448,N_2610);
nand U3915 (N_3915,N_2517,N_2025);
xnor U3916 (N_3916,N_2586,N_2022);
and U3917 (N_3917,N_2886,N_2498);
xnor U3918 (N_3918,N_2399,N_2041);
nor U3919 (N_3919,N_2790,N_2512);
nand U3920 (N_3920,N_2463,N_2982);
nand U3921 (N_3921,N_2872,N_2359);
and U3922 (N_3922,N_2502,N_2922);
and U3923 (N_3923,N_2792,N_2230);
nand U3924 (N_3924,N_2115,N_2836);
nor U3925 (N_3925,N_2825,N_2065);
and U3926 (N_3926,N_2583,N_2766);
and U3927 (N_3927,N_2732,N_2081);
nor U3928 (N_3928,N_2994,N_2256);
and U3929 (N_3929,N_2739,N_2675);
or U3930 (N_3930,N_2389,N_2270);
or U3931 (N_3931,N_2662,N_2983);
and U3932 (N_3932,N_2138,N_2280);
nand U3933 (N_3933,N_2544,N_2396);
or U3934 (N_3934,N_2480,N_2957);
or U3935 (N_3935,N_2746,N_2732);
nand U3936 (N_3936,N_2094,N_2640);
nor U3937 (N_3937,N_2430,N_2967);
xnor U3938 (N_3938,N_2597,N_2349);
xnor U3939 (N_3939,N_2819,N_2773);
nand U3940 (N_3940,N_2853,N_2598);
nand U3941 (N_3941,N_2487,N_2269);
or U3942 (N_3942,N_2685,N_2906);
and U3943 (N_3943,N_2591,N_2186);
nand U3944 (N_3944,N_2126,N_2247);
xor U3945 (N_3945,N_2504,N_2952);
or U3946 (N_3946,N_2107,N_2871);
nor U3947 (N_3947,N_2364,N_2031);
and U3948 (N_3948,N_2782,N_2095);
xor U3949 (N_3949,N_2056,N_2218);
nand U3950 (N_3950,N_2252,N_2403);
and U3951 (N_3951,N_2091,N_2039);
nand U3952 (N_3952,N_2277,N_2900);
nor U3953 (N_3953,N_2832,N_2871);
nor U3954 (N_3954,N_2211,N_2426);
nor U3955 (N_3955,N_2305,N_2798);
xor U3956 (N_3956,N_2660,N_2947);
xor U3957 (N_3957,N_2032,N_2291);
nand U3958 (N_3958,N_2642,N_2842);
xnor U3959 (N_3959,N_2133,N_2765);
nor U3960 (N_3960,N_2725,N_2824);
nand U3961 (N_3961,N_2896,N_2916);
nand U3962 (N_3962,N_2742,N_2398);
nor U3963 (N_3963,N_2637,N_2378);
xor U3964 (N_3964,N_2047,N_2099);
nand U3965 (N_3965,N_2343,N_2908);
and U3966 (N_3966,N_2370,N_2067);
and U3967 (N_3967,N_2585,N_2438);
xnor U3968 (N_3968,N_2232,N_2956);
and U3969 (N_3969,N_2126,N_2044);
xnor U3970 (N_3970,N_2725,N_2390);
nand U3971 (N_3971,N_2967,N_2540);
nor U3972 (N_3972,N_2294,N_2593);
nor U3973 (N_3973,N_2599,N_2978);
and U3974 (N_3974,N_2374,N_2794);
xnor U3975 (N_3975,N_2935,N_2533);
or U3976 (N_3976,N_2299,N_2128);
nor U3977 (N_3977,N_2167,N_2400);
nor U3978 (N_3978,N_2452,N_2694);
and U3979 (N_3979,N_2928,N_2999);
nand U3980 (N_3980,N_2136,N_2230);
nand U3981 (N_3981,N_2927,N_2039);
and U3982 (N_3982,N_2477,N_2673);
and U3983 (N_3983,N_2465,N_2186);
nor U3984 (N_3984,N_2426,N_2149);
and U3985 (N_3985,N_2218,N_2930);
or U3986 (N_3986,N_2851,N_2003);
nand U3987 (N_3987,N_2099,N_2545);
and U3988 (N_3988,N_2381,N_2023);
nand U3989 (N_3989,N_2284,N_2503);
nand U3990 (N_3990,N_2194,N_2289);
nor U3991 (N_3991,N_2196,N_2954);
xnor U3992 (N_3992,N_2140,N_2384);
nand U3993 (N_3993,N_2218,N_2661);
or U3994 (N_3994,N_2914,N_2084);
nor U3995 (N_3995,N_2298,N_2666);
xor U3996 (N_3996,N_2359,N_2164);
nor U3997 (N_3997,N_2579,N_2828);
xor U3998 (N_3998,N_2351,N_2649);
nor U3999 (N_3999,N_2027,N_2198);
or U4000 (N_4000,N_3688,N_3798);
xor U4001 (N_4001,N_3276,N_3216);
nor U4002 (N_4002,N_3293,N_3926);
and U4003 (N_4003,N_3872,N_3130);
xnor U4004 (N_4004,N_3260,N_3643);
nand U4005 (N_4005,N_3546,N_3939);
nand U4006 (N_4006,N_3889,N_3242);
nand U4007 (N_4007,N_3214,N_3834);
and U4008 (N_4008,N_3149,N_3487);
and U4009 (N_4009,N_3364,N_3739);
or U4010 (N_4010,N_3353,N_3036);
xor U4011 (N_4011,N_3785,N_3005);
nand U4012 (N_4012,N_3104,N_3700);
or U4013 (N_4013,N_3191,N_3317);
xnor U4014 (N_4014,N_3995,N_3135);
and U4015 (N_4015,N_3741,N_3031);
and U4016 (N_4016,N_3103,N_3307);
or U4017 (N_4017,N_3316,N_3596);
or U4018 (N_4018,N_3511,N_3070);
nor U4019 (N_4019,N_3342,N_3318);
or U4020 (N_4020,N_3415,N_3083);
and U4021 (N_4021,N_3057,N_3951);
or U4022 (N_4022,N_3388,N_3246);
nand U4023 (N_4023,N_3780,N_3699);
and U4024 (N_4024,N_3136,N_3393);
nand U4025 (N_4025,N_3618,N_3877);
or U4026 (N_4026,N_3266,N_3380);
and U4027 (N_4027,N_3254,N_3349);
and U4028 (N_4028,N_3114,N_3505);
nand U4029 (N_4029,N_3177,N_3444);
nor U4030 (N_4030,N_3251,N_3760);
and U4031 (N_4031,N_3174,N_3754);
or U4032 (N_4032,N_3331,N_3876);
or U4033 (N_4033,N_3516,N_3059);
nand U4034 (N_4034,N_3740,N_3265);
nand U4035 (N_4035,N_3264,N_3051);
or U4036 (N_4036,N_3115,N_3544);
nor U4037 (N_4037,N_3621,N_3817);
and U4038 (N_4038,N_3608,N_3719);
nand U4039 (N_4039,N_3645,N_3166);
and U4040 (N_4040,N_3284,N_3126);
and U4041 (N_4041,N_3370,N_3923);
nor U4042 (N_4042,N_3198,N_3244);
nor U4043 (N_4043,N_3938,N_3795);
nand U4044 (N_4044,N_3522,N_3549);
and U4045 (N_4045,N_3397,N_3194);
xnor U4046 (N_4046,N_3110,N_3079);
or U4047 (N_4047,N_3997,N_3459);
xnor U4048 (N_4048,N_3150,N_3519);
nor U4049 (N_4049,N_3275,N_3170);
nor U4050 (N_4050,N_3722,N_3774);
nor U4051 (N_4051,N_3196,N_3205);
or U4052 (N_4052,N_3202,N_3704);
or U4053 (N_4053,N_3300,N_3580);
xnor U4054 (N_4054,N_3280,N_3160);
nand U4055 (N_4055,N_3838,N_3658);
or U4056 (N_4056,N_3282,N_3882);
and U4057 (N_4057,N_3241,N_3961);
or U4058 (N_4058,N_3387,N_3382);
nand U4059 (N_4059,N_3861,N_3528);
nand U4060 (N_4060,N_3339,N_3358);
or U4061 (N_4061,N_3678,N_3008);
xor U4062 (N_4062,N_3928,N_3374);
and U4063 (N_4063,N_3237,N_3726);
xnor U4064 (N_4064,N_3659,N_3981);
nor U4065 (N_4065,N_3402,N_3234);
nor U4066 (N_4066,N_3967,N_3586);
or U4067 (N_4067,N_3429,N_3159);
nor U4068 (N_4068,N_3381,N_3482);
xor U4069 (N_4069,N_3035,N_3909);
nor U4070 (N_4070,N_3306,N_3960);
nand U4071 (N_4071,N_3852,N_3014);
nand U4072 (N_4072,N_3994,N_3232);
and U4073 (N_4073,N_3674,N_3099);
xnor U4074 (N_4074,N_3753,N_3844);
or U4075 (N_4075,N_3750,N_3653);
xnor U4076 (N_4076,N_3458,N_3792);
and U4077 (N_4077,N_3779,N_3540);
or U4078 (N_4078,N_3428,N_3343);
nand U4079 (N_4079,N_3421,N_3281);
xnor U4080 (N_4080,N_3527,N_3143);
or U4081 (N_4081,N_3647,N_3408);
nor U4082 (N_4082,N_3466,N_3835);
nor U4083 (N_4083,N_3496,N_3173);
xnor U4084 (N_4084,N_3662,N_3649);
nor U4085 (N_4085,N_3682,N_3425);
or U4086 (N_4086,N_3555,N_3042);
or U4087 (N_4087,N_3144,N_3980);
or U4088 (N_4088,N_3052,N_3147);
xor U4089 (N_4089,N_3705,N_3820);
or U4090 (N_4090,N_3058,N_3289);
and U4091 (N_4091,N_3805,N_3711);
xnor U4092 (N_4092,N_3684,N_3350);
and U4093 (N_4093,N_3533,N_3373);
and U4094 (N_4094,N_3913,N_3475);
and U4095 (N_4095,N_3512,N_3957);
nor U4096 (N_4096,N_3776,N_3292);
nand U4097 (N_4097,N_3590,N_3966);
nand U4098 (N_4098,N_3921,N_3192);
xor U4099 (N_4099,N_3417,N_3568);
xnor U4100 (N_4100,N_3329,N_3165);
nand U4101 (N_4101,N_3901,N_3521);
nor U4102 (N_4102,N_3401,N_3773);
nand U4103 (N_4103,N_3561,N_3255);
and U4104 (N_4104,N_3570,N_3607);
or U4105 (N_4105,N_3133,N_3984);
nand U4106 (N_4106,N_3474,N_3629);
and U4107 (N_4107,N_3573,N_3864);
xnor U4108 (N_4108,N_3377,N_3403);
nor U4109 (N_4109,N_3538,N_3751);
or U4110 (N_4110,N_3341,N_3491);
xor U4111 (N_4111,N_3239,N_3322);
nand U4112 (N_4112,N_3175,N_3526);
xnor U4113 (N_4113,N_3319,N_3932);
nand U4114 (N_4114,N_3167,N_3634);
nand U4115 (N_4115,N_3900,N_3811);
or U4116 (N_4116,N_3182,N_3632);
nor U4117 (N_4117,N_3209,N_3507);
or U4118 (N_4118,N_3438,N_3611);
nand U4119 (N_4119,N_3467,N_3414);
nand U4120 (N_4120,N_3944,N_3652);
xnor U4121 (N_4121,N_3420,N_3825);
xnor U4122 (N_4122,N_3077,N_3724);
or U4123 (N_4123,N_3671,N_3720);
nand U4124 (N_4124,N_3490,N_3016);
and U4125 (N_4125,N_3218,N_3369);
nor U4126 (N_4126,N_3639,N_3023);
xnor U4127 (N_4127,N_3258,N_3504);
or U4128 (N_4128,N_3400,N_3731);
nor U4129 (N_4129,N_3151,N_3513);
nor U4130 (N_4130,N_3821,N_3037);
nor U4131 (N_4131,N_3346,N_3692);
nor U4132 (N_4132,N_3465,N_3934);
nand U4133 (N_4133,N_3423,N_3551);
or U4134 (N_4134,N_3988,N_3911);
xnor U4135 (N_4135,N_3076,N_3125);
xor U4136 (N_4136,N_3840,N_3180);
xor U4137 (N_4137,N_3063,N_3302);
nand U4138 (N_4138,N_3105,N_3195);
nor U4139 (N_4139,N_3587,N_3286);
and U4140 (N_4140,N_3069,N_3577);
and U4141 (N_4141,N_3163,N_3305);
nor U4142 (N_4142,N_3272,N_3560);
or U4143 (N_4143,N_3407,N_3355);
nand U4144 (N_4144,N_3456,N_3865);
nor U4145 (N_4145,N_3563,N_3348);
and U4146 (N_4146,N_3723,N_3368);
and U4147 (N_4147,N_3920,N_3935);
xnor U4148 (N_4148,N_3554,N_3040);
xnor U4149 (N_4149,N_3004,N_3695);
nor U4150 (N_4150,N_3295,N_3553);
nand U4151 (N_4151,N_3033,N_3567);
nor U4152 (N_4152,N_3409,N_3091);
and U4153 (N_4153,N_3015,N_3772);
nor U4154 (N_4154,N_3579,N_3184);
or U4155 (N_4155,N_3333,N_3687);
and U4156 (N_4156,N_3890,N_3313);
or U4157 (N_4157,N_3502,N_3112);
and U4158 (N_4158,N_3169,N_3660);
xor U4159 (N_4159,N_3757,N_3509);
nor U4160 (N_4160,N_3843,N_3460);
or U4161 (N_4161,N_3665,N_3117);
and U4162 (N_4162,N_3116,N_3666);
nor U4163 (N_4163,N_3536,N_3963);
or U4164 (N_4164,N_3481,N_3049);
nor U4165 (N_4165,N_3893,N_3977);
nand U4166 (N_4166,N_3524,N_3702);
nand U4167 (N_4167,N_3569,N_3492);
and U4168 (N_4168,N_3638,N_3734);
nand U4169 (N_4169,N_3298,N_3873);
nand U4170 (N_4170,N_3471,N_3636);
or U4171 (N_4171,N_3948,N_3390);
xor U4172 (N_4172,N_3073,N_3208);
xnor U4173 (N_4173,N_3743,N_3217);
and U4174 (N_4174,N_3245,N_3455);
xnor U4175 (N_4175,N_3120,N_3028);
nor U4176 (N_4176,N_3715,N_3530);
nand U4177 (N_4177,N_3168,N_3261);
xnor U4178 (N_4178,N_3819,N_3712);
nor U4179 (N_4179,N_3219,N_3156);
nand U4180 (N_4180,N_3612,N_3309);
and U4181 (N_4181,N_3867,N_3323);
and U4182 (N_4182,N_3418,N_3493);
nand U4183 (N_4183,N_3367,N_3267);
nor U4184 (N_4184,N_3906,N_3514);
xnor U4185 (N_4185,N_3190,N_3142);
nor U4186 (N_4186,N_3154,N_3845);
or U4187 (N_4187,N_3064,N_3763);
xor U4188 (N_4188,N_3676,N_3379);
and U4189 (N_4189,N_3708,N_3030);
nand U4190 (N_4190,N_3717,N_3398);
or U4191 (N_4191,N_3290,N_3451);
xnor U4192 (N_4192,N_3899,N_3376);
nor U4193 (N_4193,N_3915,N_3791);
xnor U4194 (N_4194,N_3745,N_3206);
or U4195 (N_4195,N_3733,N_3007);
or U4196 (N_4196,N_3849,N_3066);
nor U4197 (N_4197,N_3762,N_3446);
nand U4198 (N_4198,N_3498,N_3878);
or U4199 (N_4199,N_3111,N_3445);
or U4200 (N_4200,N_3314,N_3716);
and U4201 (N_4201,N_3257,N_3140);
nor U4202 (N_4202,N_3998,N_3657);
and U4203 (N_4203,N_3537,N_3097);
or U4204 (N_4204,N_3228,N_3075);
or U4205 (N_4205,N_3161,N_3441);
nor U4206 (N_4206,N_3991,N_3777);
nor U4207 (N_4207,N_3081,N_3404);
nand U4208 (N_4208,N_3749,N_3626);
xnor U4209 (N_4209,N_3324,N_3029);
or U4210 (N_4210,N_3338,N_3085);
nor U4211 (N_4211,N_3363,N_3869);
nand U4212 (N_4212,N_3352,N_3841);
nor U4213 (N_4213,N_3854,N_3972);
nand U4214 (N_4214,N_3227,N_3856);
and U4215 (N_4215,N_3326,N_3970);
or U4216 (N_4216,N_3707,N_3250);
xor U4217 (N_4217,N_3572,N_3898);
nor U4218 (N_4218,N_3017,N_3296);
nand U4219 (N_4219,N_3646,N_3071);
and U4220 (N_4220,N_3449,N_3089);
and U4221 (N_4221,N_3617,N_3478);
nand U4222 (N_4222,N_3788,N_3171);
and U4223 (N_4223,N_3394,N_3846);
xnor U4224 (N_4224,N_3721,N_3279);
and U4225 (N_4225,N_3807,N_3894);
and U4226 (N_4226,N_3690,N_3203);
nand U4227 (N_4227,N_3942,N_3047);
nor U4228 (N_4228,N_3001,N_3936);
nor U4229 (N_4229,N_3210,N_3090);
or U4230 (N_4230,N_3238,N_3584);
and U4231 (N_4231,N_3197,N_3249);
nor U4232 (N_4232,N_3672,N_3480);
or U4233 (N_4233,N_3758,N_3902);
nor U4234 (N_4234,N_3986,N_3386);
nand U4235 (N_4235,N_3709,N_3483);
nand U4236 (N_4236,N_3435,N_3278);
nand U4237 (N_4237,N_3823,N_3153);
or U4238 (N_4238,N_3360,N_3925);
and U4239 (N_4239,N_3106,N_3134);
nor U4240 (N_4240,N_3879,N_3024);
or U4241 (N_4241,N_3630,N_3759);
or U4242 (N_4242,N_3597,N_3912);
nor U4243 (N_4243,N_3439,N_3006);
xor U4244 (N_4244,N_3810,N_3224);
and U4245 (N_4245,N_3178,N_3784);
nand U4246 (N_4246,N_3534,N_3862);
and U4247 (N_4247,N_3914,N_3887);
or U4248 (N_4248,N_3291,N_3800);
nor U4249 (N_4249,N_3486,N_3012);
or U4250 (N_4250,N_3273,N_3189);
xor U4251 (N_4251,N_3510,N_3187);
and U4252 (N_4252,N_3225,N_3801);
and U4253 (N_4253,N_3101,N_3145);
nand U4254 (N_4254,N_3405,N_3330);
nor U4255 (N_4255,N_3742,N_3685);
xnor U4256 (N_4256,N_3571,N_3054);
nor U4257 (N_4257,N_3947,N_3744);
nor U4258 (N_4258,N_3495,N_3892);
nand U4259 (N_4259,N_3804,N_3958);
nor U4260 (N_4260,N_3464,N_3829);
and U4261 (N_4261,N_3904,N_3009);
xor U4262 (N_4262,N_3764,N_3973);
nand U4263 (N_4263,N_3816,N_3631);
nand U4264 (N_4264,N_3728,N_3732);
nand U4265 (N_4265,N_3301,N_3430);
or U4266 (N_4266,N_3769,N_3606);
nor U4267 (N_4267,N_3410,N_3494);
nor U4268 (N_4268,N_3186,N_3088);
nor U4269 (N_4269,N_3508,N_3667);
nand U4270 (N_4270,N_3044,N_3858);
xor U4271 (N_4271,N_3416,N_3351);
nand U4272 (N_4272,N_3883,N_3003);
or U4273 (N_4273,N_3847,N_3055);
or U4274 (N_4274,N_3185,N_3806);
and U4275 (N_4275,N_3974,N_3000);
nor U4276 (N_4276,N_3993,N_3283);
or U4277 (N_4277,N_3499,N_3654);
or U4278 (N_4278,N_3564,N_3484);
nor U4279 (N_4279,N_3321,N_3930);
and U4280 (N_4280,N_3045,N_3679);
or U4281 (N_4281,N_3043,N_3604);
nand U4282 (N_4282,N_3616,N_3886);
or U4283 (N_4283,N_3332,N_3559);
or U4284 (N_4284,N_3593,N_3529);
and U4285 (N_4285,N_3613,N_3327);
and U4286 (N_4286,N_3027,N_3259);
or U4287 (N_4287,N_3814,N_3461);
nor U4288 (N_4288,N_3199,N_3591);
xnor U4289 (N_4289,N_3990,N_3833);
nand U4290 (N_4290,N_3975,N_3830);
nand U4291 (N_4291,N_3062,N_3422);
nor U4292 (N_4292,N_3385,N_3558);
xor U4293 (N_4293,N_3576,N_3213);
xnor U4294 (N_4294,N_3648,N_3952);
nand U4295 (N_4295,N_3022,N_3677);
nor U4296 (N_4296,N_3183,N_3694);
or U4297 (N_4297,N_3675,N_3627);
and U4298 (N_4298,N_3472,N_3927);
nand U4299 (N_4299,N_3770,N_3074);
xnor U4300 (N_4300,N_3176,N_3211);
nor U4301 (N_4301,N_3287,N_3207);
or U4302 (N_4302,N_3485,N_3395);
nand U4303 (N_4303,N_3689,N_3139);
nand U4304 (N_4304,N_3782,N_3406);
nand U4305 (N_4305,N_3794,N_3955);
nand U4306 (N_4306,N_3637,N_3738);
nor U4307 (N_4307,N_3440,N_3065);
nor U4308 (N_4308,N_3710,N_3828);
or U4309 (N_4309,N_3895,N_3378);
nand U4310 (N_4310,N_3940,N_3978);
or U4311 (N_4311,N_3315,N_3262);
nor U4312 (N_4312,N_3413,N_3411);
nor U4313 (N_4313,N_3018,N_3050);
and U4314 (N_4314,N_3714,N_3669);
or U4315 (N_4315,N_3243,N_3971);
and U4316 (N_4316,N_3802,N_3871);
and U4317 (N_4317,N_3761,N_3929);
xnor U4318 (N_4318,N_3989,N_3503);
or U4319 (N_4319,N_3859,N_3875);
xnor U4320 (N_4320,N_3737,N_3515);
or U4321 (N_4321,N_3226,N_3010);
nand U4322 (N_4322,N_3489,N_3918);
xor U4323 (N_4323,N_3556,N_3222);
or U4324 (N_4324,N_3041,N_3727);
nand U4325 (N_4325,N_3910,N_3371);
or U4326 (N_4326,N_3937,N_3651);
nand U4327 (N_4327,N_3565,N_3905);
xnor U4328 (N_4328,N_3897,N_3775);
xnor U4329 (N_4329,N_3954,N_3589);
nor U4330 (N_4330,N_3337,N_3019);
or U4331 (N_4331,N_3545,N_3442);
xnor U4332 (N_4332,N_3223,N_3310);
and U4333 (N_4333,N_3703,N_3344);
nor U4334 (N_4334,N_3020,N_3427);
or U4335 (N_4335,N_3581,N_3119);
xor U4336 (N_4336,N_3131,N_3247);
or U4337 (N_4337,N_3548,N_3949);
nand U4338 (N_4338,N_3221,N_3768);
xor U4339 (N_4339,N_3907,N_3432);
nand U4340 (N_4340,N_3736,N_3888);
xor U4341 (N_4341,N_3582,N_3056);
nand U4342 (N_4342,N_3334,N_3832);
nor U4343 (N_4343,N_3633,N_3599);
nor U4344 (N_4344,N_3320,N_3303);
and U4345 (N_4345,N_3285,N_3434);
nand U4346 (N_4346,N_3547,N_3152);
nor U4347 (N_4347,N_3755,N_3078);
and U4348 (N_4348,N_3746,N_3641);
nor U4349 (N_4349,N_3855,N_3575);
and U4350 (N_4350,N_3706,N_3389);
or U4351 (N_4351,N_3525,N_3375);
nand U4352 (N_4352,N_3297,N_3668);
or U4353 (N_4353,N_3574,N_3808);
nor U4354 (N_4354,N_3725,N_3543);
nand U4355 (N_4355,N_3842,N_3096);
xor U4356 (N_4356,N_3874,N_3697);
and U4357 (N_4357,N_3655,N_3673);
and U4358 (N_4358,N_3236,N_3274);
and U4359 (N_4359,N_3793,N_3122);
and U4360 (N_4360,N_3240,N_3476);
nor U4361 (N_4361,N_3453,N_3870);
and U4362 (N_4362,N_3962,N_3635);
nand U4363 (N_4363,N_3866,N_3470);
and U4364 (N_4364,N_3068,N_3778);
nand U4365 (N_4365,N_3557,N_3229);
nand U4366 (N_4366,N_3092,N_3908);
xnor U4367 (N_4367,N_3796,N_3787);
nand U4368 (N_4368,N_3082,N_3048);
nand U4369 (N_4369,N_3248,N_3881);
or U4370 (N_4370,N_3701,N_3448);
xnor U4371 (N_4371,N_3931,N_3578);
and U4372 (N_4372,N_3462,N_3263);
and U4373 (N_4373,N_3625,N_3797);
nor U4374 (N_4374,N_3128,N_3964);
or U4375 (N_4375,N_3628,N_3138);
xnor U4376 (N_4376,N_3094,N_3396);
or U4377 (N_4377,N_3450,N_3436);
nor U4378 (N_4378,N_3362,N_3880);
or U4379 (N_4379,N_3518,N_3179);
xnor U4380 (N_4380,N_3826,N_3201);
nor U4381 (N_4381,N_3391,N_3468);
nor U4382 (N_4382,N_3691,N_3756);
and U4383 (N_4383,N_3539,N_3809);
or U4384 (N_4384,N_3884,N_3693);
nor U4385 (N_4385,N_3452,N_3137);
nand U4386 (N_4386,N_3968,N_3836);
nand U4387 (N_4387,N_3624,N_3506);
or U4388 (N_4388,N_3956,N_3132);
nor U4389 (N_4389,N_3497,N_3304);
and U4390 (N_4390,N_3299,N_3598);
nand U4391 (N_4391,N_3851,N_3039);
and U4392 (N_4392,N_3002,N_3294);
xor U4393 (N_4393,N_3552,N_3595);
nor U4394 (N_4394,N_3583,N_3277);
and U4395 (N_4395,N_3384,N_3789);
nand U4396 (N_4396,N_3469,N_3288);
nor U4397 (N_4397,N_3399,N_3457);
xor U4398 (N_4398,N_3098,N_3479);
nand U4399 (N_4399,N_3992,N_3347);
or U4400 (N_4400,N_3034,N_3328);
nor U4401 (N_4401,N_3523,N_3193);
or U4402 (N_4402,N_3325,N_3614);
nor U4403 (N_4403,N_3270,N_3146);
nand U4404 (N_4404,N_3520,N_3383);
xnor U4405 (N_4405,N_3609,N_3781);
or U4406 (N_4406,N_3025,N_3500);
nand U4407 (N_4407,N_3412,N_3366);
nand U4408 (N_4408,N_3072,N_3230);
and U4409 (N_4409,N_3477,N_3803);
nor U4410 (N_4410,N_3361,N_3357);
nor U4411 (N_4411,N_3786,N_3959);
and U4412 (N_4412,N_3924,N_3021);
and U4413 (N_4413,N_3437,N_3424);
xnor U4414 (N_4414,N_3747,N_3831);
or U4415 (N_4415,N_3850,N_3681);
xor U4416 (N_4416,N_3969,N_3896);
nand U4417 (N_4417,N_3535,N_3813);
xor U4418 (N_4418,N_3686,N_3670);
nand U4419 (N_4419,N_3100,N_3312);
or U4420 (N_4420,N_3335,N_3982);
and U4421 (N_4421,N_3080,N_3164);
nand U4422 (N_4422,N_3999,N_3155);
nor U4423 (N_4423,N_3650,N_3108);
or U4424 (N_4424,N_3783,N_3550);
nand U4425 (N_4425,N_3588,N_3121);
xnor U4426 (N_4426,N_3188,N_3656);
nand U4427 (N_4427,N_3118,N_3663);
nand U4428 (N_4428,N_3933,N_3824);
or U4429 (N_4429,N_3729,N_3987);
and U4430 (N_4430,N_3696,N_3392);
or U4431 (N_4431,N_3212,N_3113);
nor U4432 (N_4432,N_3356,N_3765);
nand U4433 (N_4433,N_3945,N_3256);
nor U4434 (N_4434,N_3766,N_3231);
and U4435 (N_4435,N_3965,N_3532);
and U4436 (N_4436,N_3235,N_3473);
and U4437 (N_4437,N_3129,N_3046);
nor U4438 (N_4438,N_3107,N_3013);
xor U4439 (N_4439,N_3815,N_3640);
or U4440 (N_4440,N_3853,N_3683);
nand U4441 (N_4441,N_3252,N_3891);
or U4442 (N_4442,N_3067,N_3095);
or U4443 (N_4443,N_3172,N_3433);
and U4444 (N_4444,N_3501,N_3610);
xor U4445 (N_4445,N_3735,N_3308);
or U4446 (N_4446,N_3642,N_3748);
or U4447 (N_4447,N_3517,N_3200);
nor U4448 (N_4448,N_3976,N_3102);
nor U4449 (N_4449,N_3268,N_3790);
nand U4450 (N_4450,N_3087,N_3162);
nand U4451 (N_4451,N_3086,N_3541);
and U4452 (N_4452,N_3032,N_3233);
nand U4453 (N_4453,N_3839,N_3060);
and U4454 (N_4454,N_3916,N_3336);
and U4455 (N_4455,N_3903,N_3799);
xnor U4456 (N_4456,N_3623,N_3127);
nand U4457 (N_4457,N_3426,N_3605);
xor U4458 (N_4458,N_3919,N_3827);
and U4459 (N_4459,N_3141,N_3359);
nor U4460 (N_4460,N_3619,N_3837);
and U4461 (N_4461,N_3592,N_3848);
nand U4462 (N_4462,N_3620,N_3983);
xor U4463 (N_4463,N_3585,N_3953);
nor U4464 (N_4464,N_3941,N_3985);
xor U4465 (N_4465,N_3011,N_3269);
nor U4466 (N_4466,N_3767,N_3488);
nand U4467 (N_4467,N_3812,N_3109);
nor U4468 (N_4468,N_3602,N_3124);
nor U4469 (N_4469,N_3818,N_3615);
nor U4470 (N_4470,N_3311,N_3542);
nand U4471 (N_4471,N_3038,N_3026);
xnor U4472 (N_4472,N_3664,N_3093);
or U4473 (N_4473,N_3372,N_3730);
xnor U4474 (N_4474,N_3061,N_3698);
nor U4475 (N_4475,N_3454,N_3996);
or U4476 (N_4476,N_3603,N_3885);
xor U4477 (N_4477,N_3566,N_3644);
nor U4478 (N_4478,N_3463,N_3345);
xor U4479 (N_4479,N_3443,N_3868);
or U4480 (N_4480,N_3447,N_3123);
nor U4481 (N_4481,N_3340,N_3860);
nor U4482 (N_4482,N_3622,N_3917);
nand U4483 (N_4483,N_3661,N_3220);
xor U4484 (N_4484,N_3562,N_3943);
nand U4485 (N_4485,N_3771,N_3922);
xor U4486 (N_4486,N_3271,N_3946);
nand U4487 (N_4487,N_3601,N_3713);
and U4488 (N_4488,N_3594,N_3215);
nor U4489 (N_4489,N_3822,N_3354);
xnor U4490 (N_4490,N_3718,N_3148);
nand U4491 (N_4491,N_3979,N_3157);
nor U4492 (N_4492,N_3863,N_3680);
nand U4493 (N_4493,N_3084,N_3158);
and U4494 (N_4494,N_3950,N_3857);
nand U4495 (N_4495,N_3600,N_3253);
and U4496 (N_4496,N_3204,N_3431);
nand U4497 (N_4497,N_3752,N_3531);
or U4498 (N_4498,N_3053,N_3419);
or U4499 (N_4499,N_3181,N_3365);
and U4500 (N_4500,N_3711,N_3125);
and U4501 (N_4501,N_3787,N_3710);
nor U4502 (N_4502,N_3246,N_3076);
nand U4503 (N_4503,N_3479,N_3606);
and U4504 (N_4504,N_3712,N_3014);
nor U4505 (N_4505,N_3066,N_3128);
nor U4506 (N_4506,N_3480,N_3565);
nand U4507 (N_4507,N_3883,N_3119);
xor U4508 (N_4508,N_3603,N_3130);
and U4509 (N_4509,N_3154,N_3057);
and U4510 (N_4510,N_3887,N_3573);
nor U4511 (N_4511,N_3831,N_3780);
or U4512 (N_4512,N_3754,N_3059);
or U4513 (N_4513,N_3824,N_3219);
and U4514 (N_4514,N_3127,N_3388);
and U4515 (N_4515,N_3504,N_3719);
nand U4516 (N_4516,N_3990,N_3073);
nor U4517 (N_4517,N_3357,N_3691);
or U4518 (N_4518,N_3079,N_3161);
xor U4519 (N_4519,N_3425,N_3030);
nor U4520 (N_4520,N_3283,N_3998);
xor U4521 (N_4521,N_3588,N_3637);
or U4522 (N_4522,N_3563,N_3557);
nand U4523 (N_4523,N_3590,N_3892);
and U4524 (N_4524,N_3780,N_3966);
nor U4525 (N_4525,N_3858,N_3984);
or U4526 (N_4526,N_3844,N_3237);
or U4527 (N_4527,N_3886,N_3474);
or U4528 (N_4528,N_3798,N_3855);
or U4529 (N_4529,N_3487,N_3444);
nor U4530 (N_4530,N_3041,N_3240);
or U4531 (N_4531,N_3783,N_3530);
nor U4532 (N_4532,N_3617,N_3261);
xnor U4533 (N_4533,N_3664,N_3318);
and U4534 (N_4534,N_3686,N_3585);
xor U4535 (N_4535,N_3247,N_3141);
nand U4536 (N_4536,N_3161,N_3927);
nand U4537 (N_4537,N_3633,N_3772);
and U4538 (N_4538,N_3201,N_3226);
or U4539 (N_4539,N_3606,N_3511);
xor U4540 (N_4540,N_3610,N_3594);
xnor U4541 (N_4541,N_3167,N_3089);
nor U4542 (N_4542,N_3123,N_3601);
xnor U4543 (N_4543,N_3468,N_3001);
nand U4544 (N_4544,N_3999,N_3140);
or U4545 (N_4545,N_3756,N_3709);
nand U4546 (N_4546,N_3273,N_3268);
or U4547 (N_4547,N_3441,N_3711);
or U4548 (N_4548,N_3877,N_3156);
or U4549 (N_4549,N_3006,N_3970);
or U4550 (N_4550,N_3526,N_3938);
nand U4551 (N_4551,N_3473,N_3686);
nand U4552 (N_4552,N_3255,N_3058);
and U4553 (N_4553,N_3752,N_3818);
and U4554 (N_4554,N_3865,N_3611);
nor U4555 (N_4555,N_3226,N_3699);
xnor U4556 (N_4556,N_3341,N_3797);
nand U4557 (N_4557,N_3653,N_3352);
xnor U4558 (N_4558,N_3285,N_3198);
nor U4559 (N_4559,N_3028,N_3248);
nand U4560 (N_4560,N_3166,N_3437);
nor U4561 (N_4561,N_3915,N_3818);
nand U4562 (N_4562,N_3720,N_3240);
nor U4563 (N_4563,N_3940,N_3150);
or U4564 (N_4564,N_3809,N_3632);
xor U4565 (N_4565,N_3701,N_3496);
and U4566 (N_4566,N_3279,N_3239);
and U4567 (N_4567,N_3827,N_3692);
nand U4568 (N_4568,N_3836,N_3879);
xnor U4569 (N_4569,N_3909,N_3648);
xnor U4570 (N_4570,N_3713,N_3475);
xnor U4571 (N_4571,N_3496,N_3131);
or U4572 (N_4572,N_3623,N_3878);
nor U4573 (N_4573,N_3018,N_3468);
or U4574 (N_4574,N_3731,N_3490);
and U4575 (N_4575,N_3812,N_3226);
nand U4576 (N_4576,N_3655,N_3500);
or U4577 (N_4577,N_3605,N_3993);
and U4578 (N_4578,N_3199,N_3175);
and U4579 (N_4579,N_3171,N_3106);
nor U4580 (N_4580,N_3343,N_3910);
xnor U4581 (N_4581,N_3647,N_3306);
nor U4582 (N_4582,N_3376,N_3364);
nor U4583 (N_4583,N_3858,N_3851);
xor U4584 (N_4584,N_3134,N_3478);
xor U4585 (N_4585,N_3095,N_3399);
xnor U4586 (N_4586,N_3575,N_3319);
or U4587 (N_4587,N_3386,N_3330);
nand U4588 (N_4588,N_3039,N_3478);
and U4589 (N_4589,N_3362,N_3942);
nand U4590 (N_4590,N_3742,N_3346);
or U4591 (N_4591,N_3561,N_3874);
or U4592 (N_4592,N_3227,N_3684);
nand U4593 (N_4593,N_3774,N_3328);
and U4594 (N_4594,N_3878,N_3822);
xor U4595 (N_4595,N_3010,N_3372);
xor U4596 (N_4596,N_3567,N_3916);
nand U4597 (N_4597,N_3440,N_3178);
and U4598 (N_4598,N_3087,N_3594);
nand U4599 (N_4599,N_3130,N_3875);
xnor U4600 (N_4600,N_3061,N_3160);
and U4601 (N_4601,N_3744,N_3155);
nand U4602 (N_4602,N_3230,N_3547);
nor U4603 (N_4603,N_3720,N_3168);
or U4604 (N_4604,N_3861,N_3834);
or U4605 (N_4605,N_3552,N_3696);
nand U4606 (N_4606,N_3673,N_3337);
xor U4607 (N_4607,N_3116,N_3962);
nand U4608 (N_4608,N_3439,N_3020);
nor U4609 (N_4609,N_3670,N_3049);
nor U4610 (N_4610,N_3288,N_3227);
nor U4611 (N_4611,N_3999,N_3243);
nor U4612 (N_4612,N_3107,N_3381);
nand U4613 (N_4613,N_3199,N_3643);
and U4614 (N_4614,N_3291,N_3953);
and U4615 (N_4615,N_3238,N_3956);
nor U4616 (N_4616,N_3037,N_3858);
and U4617 (N_4617,N_3846,N_3791);
and U4618 (N_4618,N_3668,N_3885);
or U4619 (N_4619,N_3433,N_3825);
and U4620 (N_4620,N_3926,N_3061);
nand U4621 (N_4621,N_3990,N_3504);
or U4622 (N_4622,N_3747,N_3304);
xor U4623 (N_4623,N_3294,N_3329);
nor U4624 (N_4624,N_3446,N_3966);
xnor U4625 (N_4625,N_3501,N_3297);
nand U4626 (N_4626,N_3407,N_3382);
and U4627 (N_4627,N_3087,N_3587);
nand U4628 (N_4628,N_3367,N_3457);
xnor U4629 (N_4629,N_3667,N_3520);
or U4630 (N_4630,N_3579,N_3633);
and U4631 (N_4631,N_3538,N_3179);
nand U4632 (N_4632,N_3913,N_3432);
and U4633 (N_4633,N_3616,N_3290);
or U4634 (N_4634,N_3838,N_3211);
xor U4635 (N_4635,N_3158,N_3525);
or U4636 (N_4636,N_3654,N_3641);
or U4637 (N_4637,N_3920,N_3980);
or U4638 (N_4638,N_3089,N_3291);
xnor U4639 (N_4639,N_3160,N_3201);
and U4640 (N_4640,N_3391,N_3710);
xor U4641 (N_4641,N_3236,N_3705);
and U4642 (N_4642,N_3978,N_3486);
xnor U4643 (N_4643,N_3805,N_3247);
and U4644 (N_4644,N_3221,N_3153);
or U4645 (N_4645,N_3693,N_3104);
and U4646 (N_4646,N_3439,N_3315);
xnor U4647 (N_4647,N_3921,N_3673);
and U4648 (N_4648,N_3315,N_3539);
xor U4649 (N_4649,N_3601,N_3913);
xnor U4650 (N_4650,N_3775,N_3514);
or U4651 (N_4651,N_3327,N_3268);
xnor U4652 (N_4652,N_3159,N_3475);
or U4653 (N_4653,N_3506,N_3849);
or U4654 (N_4654,N_3991,N_3727);
and U4655 (N_4655,N_3507,N_3865);
nor U4656 (N_4656,N_3880,N_3290);
xnor U4657 (N_4657,N_3988,N_3144);
or U4658 (N_4658,N_3631,N_3515);
nand U4659 (N_4659,N_3401,N_3590);
nand U4660 (N_4660,N_3745,N_3028);
xnor U4661 (N_4661,N_3750,N_3414);
nand U4662 (N_4662,N_3519,N_3528);
and U4663 (N_4663,N_3408,N_3241);
and U4664 (N_4664,N_3876,N_3676);
nor U4665 (N_4665,N_3737,N_3508);
xor U4666 (N_4666,N_3024,N_3495);
and U4667 (N_4667,N_3720,N_3944);
xor U4668 (N_4668,N_3977,N_3872);
nor U4669 (N_4669,N_3748,N_3840);
or U4670 (N_4670,N_3302,N_3628);
or U4671 (N_4671,N_3614,N_3213);
and U4672 (N_4672,N_3694,N_3019);
or U4673 (N_4673,N_3585,N_3036);
xnor U4674 (N_4674,N_3901,N_3279);
xnor U4675 (N_4675,N_3659,N_3060);
and U4676 (N_4676,N_3294,N_3842);
and U4677 (N_4677,N_3839,N_3136);
or U4678 (N_4678,N_3750,N_3789);
xnor U4679 (N_4679,N_3907,N_3972);
or U4680 (N_4680,N_3331,N_3217);
and U4681 (N_4681,N_3773,N_3848);
nor U4682 (N_4682,N_3523,N_3625);
xor U4683 (N_4683,N_3040,N_3873);
xnor U4684 (N_4684,N_3461,N_3026);
nor U4685 (N_4685,N_3689,N_3150);
nand U4686 (N_4686,N_3755,N_3680);
or U4687 (N_4687,N_3134,N_3952);
nor U4688 (N_4688,N_3926,N_3020);
or U4689 (N_4689,N_3784,N_3321);
or U4690 (N_4690,N_3063,N_3689);
nand U4691 (N_4691,N_3571,N_3023);
xnor U4692 (N_4692,N_3345,N_3722);
and U4693 (N_4693,N_3504,N_3433);
xor U4694 (N_4694,N_3326,N_3956);
or U4695 (N_4695,N_3352,N_3833);
or U4696 (N_4696,N_3466,N_3349);
nand U4697 (N_4697,N_3849,N_3234);
xor U4698 (N_4698,N_3516,N_3517);
nand U4699 (N_4699,N_3856,N_3244);
or U4700 (N_4700,N_3866,N_3666);
nand U4701 (N_4701,N_3010,N_3351);
and U4702 (N_4702,N_3577,N_3087);
or U4703 (N_4703,N_3522,N_3177);
nand U4704 (N_4704,N_3529,N_3316);
and U4705 (N_4705,N_3660,N_3381);
or U4706 (N_4706,N_3544,N_3812);
nor U4707 (N_4707,N_3038,N_3081);
or U4708 (N_4708,N_3937,N_3563);
xor U4709 (N_4709,N_3868,N_3686);
and U4710 (N_4710,N_3901,N_3630);
nand U4711 (N_4711,N_3206,N_3756);
nor U4712 (N_4712,N_3110,N_3977);
and U4713 (N_4713,N_3081,N_3658);
nand U4714 (N_4714,N_3652,N_3457);
xor U4715 (N_4715,N_3249,N_3280);
or U4716 (N_4716,N_3406,N_3273);
nor U4717 (N_4717,N_3417,N_3099);
and U4718 (N_4718,N_3885,N_3384);
nor U4719 (N_4719,N_3510,N_3056);
xnor U4720 (N_4720,N_3854,N_3821);
nor U4721 (N_4721,N_3641,N_3607);
xor U4722 (N_4722,N_3167,N_3548);
nand U4723 (N_4723,N_3475,N_3014);
xnor U4724 (N_4724,N_3346,N_3762);
nor U4725 (N_4725,N_3425,N_3695);
nand U4726 (N_4726,N_3291,N_3789);
nor U4727 (N_4727,N_3834,N_3958);
and U4728 (N_4728,N_3410,N_3835);
nor U4729 (N_4729,N_3709,N_3682);
nand U4730 (N_4730,N_3512,N_3193);
xor U4731 (N_4731,N_3108,N_3636);
nand U4732 (N_4732,N_3150,N_3633);
or U4733 (N_4733,N_3398,N_3537);
nand U4734 (N_4734,N_3102,N_3670);
nor U4735 (N_4735,N_3575,N_3712);
nand U4736 (N_4736,N_3724,N_3540);
or U4737 (N_4737,N_3605,N_3213);
nand U4738 (N_4738,N_3588,N_3409);
xor U4739 (N_4739,N_3090,N_3060);
xor U4740 (N_4740,N_3060,N_3000);
nand U4741 (N_4741,N_3250,N_3553);
xor U4742 (N_4742,N_3093,N_3406);
and U4743 (N_4743,N_3664,N_3581);
and U4744 (N_4744,N_3260,N_3407);
xnor U4745 (N_4745,N_3054,N_3798);
or U4746 (N_4746,N_3702,N_3705);
nand U4747 (N_4747,N_3784,N_3761);
nor U4748 (N_4748,N_3761,N_3030);
or U4749 (N_4749,N_3393,N_3097);
nor U4750 (N_4750,N_3086,N_3681);
nand U4751 (N_4751,N_3675,N_3902);
and U4752 (N_4752,N_3403,N_3645);
or U4753 (N_4753,N_3622,N_3815);
nand U4754 (N_4754,N_3910,N_3109);
nand U4755 (N_4755,N_3445,N_3736);
or U4756 (N_4756,N_3400,N_3564);
xor U4757 (N_4757,N_3477,N_3146);
xnor U4758 (N_4758,N_3354,N_3636);
nand U4759 (N_4759,N_3478,N_3079);
and U4760 (N_4760,N_3644,N_3704);
nor U4761 (N_4761,N_3085,N_3951);
nand U4762 (N_4762,N_3019,N_3400);
nor U4763 (N_4763,N_3599,N_3644);
and U4764 (N_4764,N_3991,N_3383);
or U4765 (N_4765,N_3865,N_3470);
or U4766 (N_4766,N_3840,N_3734);
or U4767 (N_4767,N_3644,N_3521);
nor U4768 (N_4768,N_3129,N_3174);
or U4769 (N_4769,N_3406,N_3092);
nand U4770 (N_4770,N_3614,N_3723);
or U4771 (N_4771,N_3160,N_3595);
nand U4772 (N_4772,N_3486,N_3706);
xor U4773 (N_4773,N_3149,N_3596);
xnor U4774 (N_4774,N_3728,N_3695);
or U4775 (N_4775,N_3956,N_3579);
and U4776 (N_4776,N_3710,N_3994);
xnor U4777 (N_4777,N_3841,N_3319);
nand U4778 (N_4778,N_3634,N_3435);
or U4779 (N_4779,N_3733,N_3942);
xor U4780 (N_4780,N_3680,N_3832);
xor U4781 (N_4781,N_3894,N_3330);
nand U4782 (N_4782,N_3967,N_3825);
and U4783 (N_4783,N_3985,N_3946);
and U4784 (N_4784,N_3282,N_3150);
nor U4785 (N_4785,N_3229,N_3763);
nand U4786 (N_4786,N_3013,N_3484);
xnor U4787 (N_4787,N_3391,N_3387);
or U4788 (N_4788,N_3745,N_3562);
nand U4789 (N_4789,N_3117,N_3878);
nand U4790 (N_4790,N_3874,N_3642);
and U4791 (N_4791,N_3132,N_3217);
xnor U4792 (N_4792,N_3753,N_3980);
nor U4793 (N_4793,N_3489,N_3567);
nand U4794 (N_4794,N_3883,N_3071);
or U4795 (N_4795,N_3454,N_3827);
or U4796 (N_4796,N_3034,N_3562);
and U4797 (N_4797,N_3532,N_3579);
xor U4798 (N_4798,N_3110,N_3872);
or U4799 (N_4799,N_3838,N_3177);
or U4800 (N_4800,N_3715,N_3004);
xnor U4801 (N_4801,N_3581,N_3884);
nand U4802 (N_4802,N_3431,N_3901);
nor U4803 (N_4803,N_3650,N_3656);
and U4804 (N_4804,N_3609,N_3811);
nor U4805 (N_4805,N_3281,N_3810);
and U4806 (N_4806,N_3024,N_3393);
nor U4807 (N_4807,N_3145,N_3033);
or U4808 (N_4808,N_3278,N_3788);
and U4809 (N_4809,N_3860,N_3949);
xnor U4810 (N_4810,N_3303,N_3098);
nand U4811 (N_4811,N_3046,N_3956);
and U4812 (N_4812,N_3652,N_3093);
nor U4813 (N_4813,N_3035,N_3818);
nor U4814 (N_4814,N_3610,N_3728);
or U4815 (N_4815,N_3619,N_3145);
xor U4816 (N_4816,N_3155,N_3158);
xor U4817 (N_4817,N_3759,N_3884);
nor U4818 (N_4818,N_3298,N_3311);
nand U4819 (N_4819,N_3453,N_3023);
nor U4820 (N_4820,N_3984,N_3059);
and U4821 (N_4821,N_3897,N_3161);
and U4822 (N_4822,N_3680,N_3861);
xor U4823 (N_4823,N_3067,N_3841);
nand U4824 (N_4824,N_3763,N_3566);
or U4825 (N_4825,N_3222,N_3873);
nor U4826 (N_4826,N_3579,N_3141);
and U4827 (N_4827,N_3442,N_3865);
or U4828 (N_4828,N_3563,N_3497);
or U4829 (N_4829,N_3718,N_3235);
xor U4830 (N_4830,N_3664,N_3390);
nand U4831 (N_4831,N_3691,N_3803);
xnor U4832 (N_4832,N_3343,N_3915);
xnor U4833 (N_4833,N_3224,N_3132);
nand U4834 (N_4834,N_3589,N_3069);
nor U4835 (N_4835,N_3565,N_3647);
xnor U4836 (N_4836,N_3418,N_3274);
and U4837 (N_4837,N_3819,N_3895);
xor U4838 (N_4838,N_3708,N_3128);
nor U4839 (N_4839,N_3767,N_3937);
xnor U4840 (N_4840,N_3098,N_3137);
xnor U4841 (N_4841,N_3554,N_3944);
xor U4842 (N_4842,N_3789,N_3583);
or U4843 (N_4843,N_3399,N_3104);
nor U4844 (N_4844,N_3306,N_3323);
xor U4845 (N_4845,N_3061,N_3683);
or U4846 (N_4846,N_3439,N_3716);
and U4847 (N_4847,N_3175,N_3417);
or U4848 (N_4848,N_3514,N_3867);
nor U4849 (N_4849,N_3647,N_3671);
xnor U4850 (N_4850,N_3973,N_3257);
xor U4851 (N_4851,N_3238,N_3385);
nor U4852 (N_4852,N_3218,N_3926);
nand U4853 (N_4853,N_3619,N_3750);
or U4854 (N_4854,N_3240,N_3954);
or U4855 (N_4855,N_3089,N_3479);
nor U4856 (N_4856,N_3859,N_3125);
nand U4857 (N_4857,N_3077,N_3243);
or U4858 (N_4858,N_3505,N_3752);
and U4859 (N_4859,N_3592,N_3654);
xnor U4860 (N_4860,N_3489,N_3878);
and U4861 (N_4861,N_3955,N_3930);
and U4862 (N_4862,N_3899,N_3161);
nor U4863 (N_4863,N_3312,N_3031);
and U4864 (N_4864,N_3305,N_3022);
and U4865 (N_4865,N_3416,N_3409);
nor U4866 (N_4866,N_3648,N_3435);
and U4867 (N_4867,N_3166,N_3543);
nand U4868 (N_4868,N_3658,N_3111);
or U4869 (N_4869,N_3045,N_3977);
nor U4870 (N_4870,N_3084,N_3879);
nand U4871 (N_4871,N_3184,N_3330);
xor U4872 (N_4872,N_3505,N_3073);
nand U4873 (N_4873,N_3507,N_3720);
xnor U4874 (N_4874,N_3580,N_3190);
and U4875 (N_4875,N_3198,N_3503);
nor U4876 (N_4876,N_3190,N_3309);
xnor U4877 (N_4877,N_3944,N_3283);
or U4878 (N_4878,N_3426,N_3778);
nand U4879 (N_4879,N_3613,N_3597);
and U4880 (N_4880,N_3783,N_3107);
nand U4881 (N_4881,N_3792,N_3026);
xor U4882 (N_4882,N_3920,N_3037);
and U4883 (N_4883,N_3559,N_3683);
nand U4884 (N_4884,N_3517,N_3392);
or U4885 (N_4885,N_3673,N_3305);
xor U4886 (N_4886,N_3730,N_3009);
and U4887 (N_4887,N_3449,N_3853);
and U4888 (N_4888,N_3763,N_3407);
nand U4889 (N_4889,N_3197,N_3487);
nor U4890 (N_4890,N_3176,N_3675);
nor U4891 (N_4891,N_3992,N_3760);
and U4892 (N_4892,N_3416,N_3331);
nor U4893 (N_4893,N_3150,N_3388);
nand U4894 (N_4894,N_3425,N_3450);
xor U4895 (N_4895,N_3646,N_3132);
nor U4896 (N_4896,N_3144,N_3285);
and U4897 (N_4897,N_3812,N_3020);
and U4898 (N_4898,N_3337,N_3996);
and U4899 (N_4899,N_3612,N_3898);
and U4900 (N_4900,N_3049,N_3136);
nand U4901 (N_4901,N_3462,N_3904);
and U4902 (N_4902,N_3181,N_3353);
and U4903 (N_4903,N_3708,N_3267);
or U4904 (N_4904,N_3517,N_3357);
and U4905 (N_4905,N_3938,N_3007);
or U4906 (N_4906,N_3276,N_3864);
nand U4907 (N_4907,N_3661,N_3782);
and U4908 (N_4908,N_3961,N_3681);
or U4909 (N_4909,N_3106,N_3088);
xor U4910 (N_4910,N_3729,N_3033);
nand U4911 (N_4911,N_3325,N_3343);
or U4912 (N_4912,N_3375,N_3321);
xnor U4913 (N_4913,N_3694,N_3006);
nor U4914 (N_4914,N_3895,N_3359);
xor U4915 (N_4915,N_3698,N_3681);
and U4916 (N_4916,N_3818,N_3781);
and U4917 (N_4917,N_3051,N_3098);
xor U4918 (N_4918,N_3725,N_3312);
and U4919 (N_4919,N_3641,N_3492);
and U4920 (N_4920,N_3417,N_3129);
or U4921 (N_4921,N_3847,N_3939);
and U4922 (N_4922,N_3378,N_3853);
and U4923 (N_4923,N_3387,N_3640);
xor U4924 (N_4924,N_3384,N_3902);
nand U4925 (N_4925,N_3359,N_3066);
or U4926 (N_4926,N_3102,N_3653);
and U4927 (N_4927,N_3094,N_3591);
nand U4928 (N_4928,N_3312,N_3166);
nor U4929 (N_4929,N_3618,N_3052);
nor U4930 (N_4930,N_3202,N_3684);
or U4931 (N_4931,N_3081,N_3909);
or U4932 (N_4932,N_3184,N_3194);
xnor U4933 (N_4933,N_3905,N_3780);
nand U4934 (N_4934,N_3043,N_3281);
nor U4935 (N_4935,N_3993,N_3507);
nor U4936 (N_4936,N_3379,N_3860);
or U4937 (N_4937,N_3931,N_3205);
xor U4938 (N_4938,N_3898,N_3968);
nor U4939 (N_4939,N_3678,N_3168);
xnor U4940 (N_4940,N_3559,N_3335);
nor U4941 (N_4941,N_3158,N_3400);
xor U4942 (N_4942,N_3879,N_3077);
or U4943 (N_4943,N_3558,N_3933);
nand U4944 (N_4944,N_3060,N_3448);
nor U4945 (N_4945,N_3322,N_3289);
nor U4946 (N_4946,N_3132,N_3668);
nor U4947 (N_4947,N_3058,N_3187);
and U4948 (N_4948,N_3339,N_3237);
xor U4949 (N_4949,N_3334,N_3085);
or U4950 (N_4950,N_3436,N_3658);
or U4951 (N_4951,N_3324,N_3974);
nand U4952 (N_4952,N_3951,N_3341);
and U4953 (N_4953,N_3144,N_3895);
or U4954 (N_4954,N_3584,N_3068);
and U4955 (N_4955,N_3081,N_3531);
nand U4956 (N_4956,N_3598,N_3008);
xor U4957 (N_4957,N_3596,N_3629);
nand U4958 (N_4958,N_3127,N_3909);
xnor U4959 (N_4959,N_3507,N_3105);
and U4960 (N_4960,N_3343,N_3320);
xor U4961 (N_4961,N_3875,N_3483);
nor U4962 (N_4962,N_3813,N_3020);
xor U4963 (N_4963,N_3047,N_3751);
or U4964 (N_4964,N_3769,N_3708);
xor U4965 (N_4965,N_3628,N_3056);
xnor U4966 (N_4966,N_3465,N_3588);
xor U4967 (N_4967,N_3231,N_3260);
and U4968 (N_4968,N_3817,N_3723);
xnor U4969 (N_4969,N_3617,N_3649);
nor U4970 (N_4970,N_3113,N_3290);
or U4971 (N_4971,N_3614,N_3920);
and U4972 (N_4972,N_3496,N_3737);
nor U4973 (N_4973,N_3595,N_3272);
nand U4974 (N_4974,N_3594,N_3842);
or U4975 (N_4975,N_3179,N_3772);
nor U4976 (N_4976,N_3209,N_3013);
or U4977 (N_4977,N_3614,N_3065);
nor U4978 (N_4978,N_3223,N_3350);
or U4979 (N_4979,N_3813,N_3599);
nand U4980 (N_4980,N_3542,N_3743);
nand U4981 (N_4981,N_3095,N_3009);
xor U4982 (N_4982,N_3869,N_3944);
or U4983 (N_4983,N_3343,N_3224);
nand U4984 (N_4984,N_3024,N_3141);
nor U4985 (N_4985,N_3528,N_3211);
xor U4986 (N_4986,N_3677,N_3018);
nand U4987 (N_4987,N_3104,N_3017);
xnor U4988 (N_4988,N_3065,N_3276);
nand U4989 (N_4989,N_3226,N_3767);
xor U4990 (N_4990,N_3754,N_3994);
and U4991 (N_4991,N_3858,N_3407);
nand U4992 (N_4992,N_3546,N_3149);
nor U4993 (N_4993,N_3801,N_3337);
or U4994 (N_4994,N_3009,N_3388);
nor U4995 (N_4995,N_3317,N_3776);
or U4996 (N_4996,N_3713,N_3814);
or U4997 (N_4997,N_3127,N_3540);
or U4998 (N_4998,N_3479,N_3464);
nand U4999 (N_4999,N_3936,N_3429);
nor U5000 (N_5000,N_4299,N_4414);
and U5001 (N_5001,N_4349,N_4888);
nand U5002 (N_5002,N_4033,N_4461);
nand U5003 (N_5003,N_4228,N_4734);
xnor U5004 (N_5004,N_4927,N_4906);
or U5005 (N_5005,N_4537,N_4398);
or U5006 (N_5006,N_4361,N_4129);
xor U5007 (N_5007,N_4519,N_4433);
nor U5008 (N_5008,N_4000,N_4728);
or U5009 (N_5009,N_4496,N_4588);
xnor U5010 (N_5010,N_4999,N_4152);
nand U5011 (N_5011,N_4786,N_4438);
and U5012 (N_5012,N_4188,N_4360);
nand U5013 (N_5013,N_4612,N_4539);
nand U5014 (N_5014,N_4611,N_4838);
nand U5015 (N_5015,N_4766,N_4536);
or U5016 (N_5016,N_4507,N_4182);
and U5017 (N_5017,N_4825,N_4965);
nor U5018 (N_5018,N_4991,N_4998);
and U5019 (N_5019,N_4269,N_4555);
nor U5020 (N_5020,N_4373,N_4463);
nor U5021 (N_5021,N_4895,N_4111);
xnor U5022 (N_5022,N_4493,N_4038);
nand U5023 (N_5023,N_4098,N_4829);
nand U5024 (N_5024,N_4444,N_4821);
and U5025 (N_5025,N_4562,N_4137);
or U5026 (N_5026,N_4451,N_4558);
xor U5027 (N_5027,N_4871,N_4093);
nand U5028 (N_5028,N_4690,N_4933);
or U5029 (N_5029,N_4079,N_4634);
and U5030 (N_5030,N_4168,N_4792);
nand U5031 (N_5031,N_4559,N_4348);
nor U5032 (N_5032,N_4913,N_4887);
or U5033 (N_5033,N_4099,N_4316);
and U5034 (N_5034,N_4653,N_4532);
xor U5035 (N_5035,N_4787,N_4785);
xor U5036 (N_5036,N_4802,N_4295);
nor U5037 (N_5037,N_4071,N_4541);
xor U5038 (N_5038,N_4637,N_4540);
nor U5039 (N_5039,N_4440,N_4533);
xnor U5040 (N_5040,N_4750,N_4151);
and U5041 (N_5041,N_4312,N_4695);
nor U5042 (N_5042,N_4229,N_4416);
nand U5043 (N_5043,N_4505,N_4307);
nor U5044 (N_5044,N_4359,N_4154);
nor U5045 (N_5045,N_4478,N_4922);
or U5046 (N_5046,N_4718,N_4242);
and U5047 (N_5047,N_4372,N_4121);
or U5048 (N_5048,N_4075,N_4894);
or U5049 (N_5049,N_4022,N_4840);
or U5050 (N_5050,N_4710,N_4934);
nor U5051 (N_5051,N_4325,N_4184);
and U5052 (N_5052,N_4827,N_4595);
nand U5053 (N_5053,N_4816,N_4091);
nor U5054 (N_5054,N_4686,N_4198);
nand U5055 (N_5055,N_4973,N_4962);
nor U5056 (N_5056,N_4388,N_4556);
nor U5057 (N_5057,N_4730,N_4270);
or U5058 (N_5058,N_4082,N_4599);
nor U5059 (N_5059,N_4133,N_4488);
xor U5060 (N_5060,N_4236,N_4631);
nor U5061 (N_5061,N_4849,N_4743);
and U5062 (N_5062,N_4553,N_4338);
or U5063 (N_5063,N_4278,N_4528);
and U5064 (N_5064,N_4592,N_4974);
xor U5065 (N_5065,N_4917,N_4944);
or U5066 (N_5066,N_4890,N_4027);
and U5067 (N_5067,N_4482,N_4935);
nand U5068 (N_5068,N_4243,N_4384);
and U5069 (N_5069,N_4529,N_4609);
nor U5070 (N_5070,N_4551,N_4465);
nand U5071 (N_5071,N_4377,N_4399);
and U5072 (N_5072,N_4097,N_4741);
nand U5073 (N_5073,N_4010,N_4050);
or U5074 (N_5074,N_4657,N_4615);
and U5075 (N_5075,N_4819,N_4445);
nand U5076 (N_5076,N_4323,N_4573);
or U5077 (N_5077,N_4402,N_4200);
xnor U5078 (N_5078,N_4818,N_4251);
nor U5079 (N_5079,N_4112,N_4471);
and U5080 (N_5080,N_4432,N_4409);
and U5081 (N_5081,N_4717,N_4520);
nor U5082 (N_5082,N_4281,N_4502);
and U5083 (N_5083,N_4313,N_4702);
or U5084 (N_5084,N_4645,N_4042);
and U5085 (N_5085,N_4067,N_4515);
xor U5086 (N_5086,N_4512,N_4777);
nor U5087 (N_5087,N_4005,N_4475);
or U5088 (N_5088,N_4382,N_4138);
xnor U5089 (N_5089,N_4814,N_4606);
nand U5090 (N_5090,N_4021,N_4337);
xnor U5091 (N_5091,N_4905,N_4090);
xor U5092 (N_5092,N_4470,N_4310);
or U5093 (N_5093,N_4969,N_4937);
and U5094 (N_5094,N_4193,N_4830);
or U5095 (N_5095,N_4430,N_4566);
or U5096 (N_5096,N_4836,N_4034);
and U5097 (N_5097,N_4638,N_4434);
and U5098 (N_5098,N_4456,N_4145);
and U5099 (N_5099,N_4896,N_4476);
or U5100 (N_5100,N_4736,N_4527);
nor U5101 (N_5101,N_4096,N_4576);
and U5102 (N_5102,N_4923,N_4538);
and U5103 (N_5103,N_4687,N_4087);
or U5104 (N_5104,N_4194,N_4682);
nand U5105 (N_5105,N_4767,N_4492);
xor U5106 (N_5106,N_4760,N_4655);
or U5107 (N_5107,N_4123,N_4288);
nand U5108 (N_5108,N_4253,N_4950);
nor U5109 (N_5109,N_4980,N_4144);
or U5110 (N_5110,N_4237,N_4983);
or U5111 (N_5111,N_4978,N_4778);
or U5112 (N_5112,N_4051,N_4904);
nor U5113 (N_5113,N_4120,N_4513);
xor U5114 (N_5114,N_4779,N_4964);
and U5115 (N_5115,N_4220,N_4635);
and U5116 (N_5116,N_4842,N_4044);
xor U5117 (N_5117,N_4833,N_4380);
nand U5118 (N_5118,N_4248,N_4055);
xor U5119 (N_5119,N_4746,N_4584);
or U5120 (N_5120,N_4720,N_4108);
nor U5121 (N_5121,N_4621,N_4692);
and U5122 (N_5122,N_4117,N_4458);
nand U5123 (N_5123,N_4049,N_4176);
nand U5124 (N_5124,N_4160,N_4632);
nor U5125 (N_5125,N_4343,N_4474);
or U5126 (N_5126,N_4350,N_4642);
xnor U5127 (N_5127,N_4367,N_4627);
nor U5128 (N_5128,N_4996,N_4428);
nand U5129 (N_5129,N_4202,N_4844);
and U5130 (N_5130,N_4158,N_4788);
nand U5131 (N_5131,N_4714,N_4375);
and U5132 (N_5132,N_4058,N_4483);
or U5133 (N_5133,N_4565,N_4708);
xor U5134 (N_5134,N_4912,N_4187);
xor U5135 (N_5135,N_4062,N_4330);
or U5136 (N_5136,N_4397,N_4166);
or U5137 (N_5137,N_4929,N_4826);
or U5138 (N_5138,N_4102,N_4086);
and U5139 (N_5139,N_4776,N_4650);
nor U5140 (N_5140,N_4092,N_4069);
xor U5141 (N_5141,N_4003,N_4164);
nor U5142 (N_5142,N_4285,N_4436);
and U5143 (N_5143,N_4548,N_4578);
xor U5144 (N_5144,N_4329,N_4754);
nor U5145 (N_5145,N_4901,N_4179);
nor U5146 (N_5146,N_4405,N_4169);
nand U5147 (N_5147,N_4389,N_4511);
and U5148 (N_5148,N_4473,N_4334);
and U5149 (N_5149,N_4809,N_4574);
nand U5150 (N_5150,N_4368,N_4413);
and U5151 (N_5151,N_4577,N_4674);
nand U5152 (N_5152,N_4346,N_4012);
or U5153 (N_5153,N_4018,N_4671);
and U5154 (N_5154,N_4489,N_4294);
and U5155 (N_5155,N_4070,N_4823);
or U5156 (N_5156,N_4298,N_4500);
nand U5157 (N_5157,N_4893,N_4870);
nand U5158 (N_5158,N_4932,N_4963);
xor U5159 (N_5159,N_4966,N_4542);
xor U5160 (N_5160,N_4157,N_4805);
or U5161 (N_5161,N_4967,N_4683);
and U5162 (N_5162,N_4410,N_4968);
and U5163 (N_5163,N_4925,N_4335);
nand U5164 (N_5164,N_4271,N_4262);
xnor U5165 (N_5165,N_4457,N_4563);
and U5166 (N_5166,N_4640,N_4585);
nand U5167 (N_5167,N_4586,N_4183);
or U5168 (N_5168,N_4256,N_4684);
or U5169 (N_5169,N_4293,N_4721);
xnor U5170 (N_5170,N_4793,N_4390);
and U5171 (N_5171,N_4404,N_4171);
nor U5172 (N_5172,N_4907,N_4442);
nand U5173 (N_5173,N_4140,N_4411);
or U5174 (N_5174,N_4715,N_4261);
and U5175 (N_5175,N_4172,N_4510);
xor U5176 (N_5176,N_4679,N_4282);
and U5177 (N_5177,N_4688,N_4813);
nor U5178 (N_5178,N_4480,N_4249);
or U5179 (N_5179,N_4088,N_4696);
and U5180 (N_5180,N_4190,N_4425);
and U5181 (N_5181,N_4909,N_4554);
xor U5182 (N_5182,N_4486,N_4061);
nand U5183 (N_5183,N_4740,N_4462);
nor U5184 (N_5184,N_4124,N_4641);
and U5185 (N_5185,N_4569,N_4989);
nand U5186 (N_5186,N_4955,N_4764);
or U5187 (N_5187,N_4835,N_4020);
xnor U5188 (N_5188,N_4834,N_4114);
nand U5189 (N_5189,N_4868,N_4794);
and U5190 (N_5190,N_4352,N_4583);
and U5191 (N_5191,N_4663,N_4659);
nor U5192 (N_5192,N_4046,N_4550);
nand U5193 (N_5193,N_4707,N_4910);
or U5194 (N_5194,N_4723,N_4747);
nand U5195 (N_5195,N_4211,N_4822);
or U5196 (N_5196,N_4644,N_4247);
nor U5197 (N_5197,N_4422,N_4737);
or U5198 (N_5198,N_4617,N_4523);
nand U5199 (N_5199,N_4869,N_4014);
xor U5200 (N_5200,N_4297,N_4233);
or U5201 (N_5201,N_4304,N_4407);
xnor U5202 (N_5202,N_4146,N_4892);
nor U5203 (N_5203,N_4872,N_4607);
and U5204 (N_5204,N_4362,N_4948);
nor U5205 (N_5205,N_4057,N_4284);
or U5206 (N_5206,N_4509,N_4296);
or U5207 (N_5207,N_4712,N_4560);
nor U5208 (N_5208,N_4264,N_4669);
nand U5209 (N_5209,N_4719,N_4775);
nor U5210 (N_5210,N_4567,N_4857);
and U5211 (N_5211,N_4985,N_4147);
nand U5212 (N_5212,N_4326,N_4689);
and U5213 (N_5213,N_4997,N_4387);
and U5214 (N_5214,N_4647,N_4081);
and U5215 (N_5215,N_4127,N_4685);
nor U5216 (N_5216,N_4235,N_4765);
nand U5217 (N_5217,N_4781,N_4455);
or U5218 (N_5218,N_4939,N_4196);
nand U5219 (N_5219,N_4733,N_4421);
xor U5220 (N_5220,N_4711,N_4226);
or U5221 (N_5221,N_4192,N_4238);
xnor U5222 (N_5222,N_4848,N_4315);
nand U5223 (N_5223,N_4303,N_4204);
and U5224 (N_5224,N_4587,N_4756);
xnor U5225 (N_5225,N_4025,N_4751);
nand U5226 (N_5226,N_4029,N_4518);
and U5227 (N_5227,N_4342,N_4678);
nand U5228 (N_5228,N_4861,N_4260);
nor U5229 (N_5229,N_4077,N_4435);
and U5230 (N_5230,N_4280,N_4947);
and U5231 (N_5231,N_4170,N_4516);
and U5232 (N_5232,N_4648,N_4898);
and U5233 (N_5233,N_4993,N_4225);
xor U5234 (N_5234,N_4064,N_4698);
and U5235 (N_5235,N_4920,N_4472);
nand U5236 (N_5236,N_4490,N_4914);
nand U5237 (N_5237,N_4265,N_4415);
nand U5238 (N_5238,N_4782,N_4481);
or U5239 (N_5239,N_4618,N_4804);
nor U5240 (N_5240,N_4068,N_4427);
nand U5241 (N_5241,N_4891,N_4713);
or U5242 (N_5242,N_4203,N_4957);
and U5243 (N_5243,N_4841,N_4995);
nand U5244 (N_5244,N_4530,N_4074);
or U5245 (N_5245,N_4916,N_4218);
or U5246 (N_5246,N_4291,N_4795);
or U5247 (N_5247,N_4662,N_4636);
and U5248 (N_5248,N_4514,N_4122);
xor U5249 (N_5249,N_4812,N_4783);
xnor U5250 (N_5250,N_4552,N_4742);
nor U5251 (N_5251,N_4956,N_4706);
or U5252 (N_5252,N_4596,N_4214);
or U5253 (N_5253,N_4216,N_4953);
and U5254 (N_5254,N_4832,N_4073);
or U5255 (N_5255,N_4448,N_4625);
nand U5256 (N_5256,N_4885,N_4768);
and U5257 (N_5257,N_4201,N_4941);
and U5258 (N_5258,N_4843,N_4860);
or U5259 (N_5259,N_4899,N_4059);
nor U5260 (N_5260,N_4806,N_4649);
or U5261 (N_5261,N_4083,N_4322);
xnor U5262 (N_5262,N_4494,N_4015);
nor U5263 (N_5263,N_4487,N_4403);
and U5264 (N_5264,N_4223,N_4469);
nand U5265 (N_5265,N_4745,N_4704);
or U5266 (N_5266,N_4283,N_4374);
and U5267 (N_5267,N_4495,N_4865);
nand U5268 (N_5268,N_4006,N_4308);
nand U5269 (N_5269,N_4579,N_4633);
and U5270 (N_5270,N_4239,N_4508);
xor U5271 (N_5271,N_4940,N_4942);
nand U5272 (N_5272,N_4884,N_4156);
nand U5273 (N_5273,N_4820,N_4009);
xor U5274 (N_5274,N_4363,N_4109);
xnor U5275 (N_5275,N_4858,N_4694);
or U5276 (N_5276,N_4936,N_4498);
and U5277 (N_5277,N_4651,N_4643);
xor U5278 (N_5278,N_4054,N_4287);
or U5279 (N_5279,N_4545,N_4453);
xnor U5280 (N_5280,N_4420,N_4180);
and U5281 (N_5281,N_4605,N_4013);
or U5282 (N_5282,N_4072,N_4866);
or U5283 (N_5283,N_4732,N_4084);
or U5284 (N_5284,N_4328,N_4406);
or U5285 (N_5285,N_4205,N_4824);
xor U5286 (N_5286,N_4401,N_4085);
and U5287 (N_5287,N_4141,N_4970);
and U5288 (N_5288,N_4060,N_4365);
and U5289 (N_5289,N_4370,N_4594);
nand U5290 (N_5290,N_4106,N_4961);
nand U5291 (N_5291,N_4371,N_4383);
nor U5292 (N_5292,N_4926,N_4676);
or U5293 (N_5293,N_4726,N_4744);
nor U5294 (N_5294,N_4626,N_4784);
or U5295 (N_5295,N_4215,N_4185);
and U5296 (N_5296,N_4811,N_4855);
or U5297 (N_5297,N_4207,N_4629);
nor U5298 (N_5298,N_4452,N_4864);
xor U5299 (N_5299,N_4103,N_4620);
xor U5300 (N_5300,N_4959,N_4725);
nand U5301 (N_5301,N_4881,N_4949);
or U5302 (N_5302,N_4801,N_4976);
xor U5303 (N_5303,N_4052,N_4526);
nor U5304 (N_5304,N_4619,N_4952);
xnor U5305 (N_5305,N_4167,N_4677);
nor U5306 (N_5306,N_4195,N_4001);
xor U5307 (N_5307,N_4104,N_4616);
or U5308 (N_5308,N_4429,N_4602);
and U5309 (N_5309,N_4378,N_4391);
or U5310 (N_5310,N_4116,N_4306);
nor U5311 (N_5311,N_4290,N_4464);
or U5312 (N_5312,N_4672,N_4863);
or U5313 (N_5313,N_4175,N_4244);
or U5314 (N_5314,N_4240,N_4990);
and U5315 (N_5315,N_4447,N_4181);
and U5316 (N_5316,N_4273,N_4155);
and U5317 (N_5317,N_4131,N_4305);
nor U5318 (N_5318,N_4639,N_4041);
nor U5319 (N_5319,N_4673,N_4454);
xor U5320 (N_5320,N_4080,N_4327);
xor U5321 (N_5321,N_4007,N_4771);
nand U5322 (N_5322,N_4219,N_4113);
xor U5323 (N_5323,N_4412,N_4546);
nand U5324 (N_5324,N_4355,N_4986);
and U5325 (N_5325,N_4867,N_4094);
and U5326 (N_5326,N_4418,N_4758);
and U5327 (N_5327,N_4808,N_4597);
and U5328 (N_5328,N_4227,N_4699);
xor U5329 (N_5329,N_4466,N_4030);
or U5330 (N_5330,N_4217,N_4666);
xor U5331 (N_5331,N_4924,N_4268);
nand U5332 (N_5332,N_4255,N_4854);
nor U5333 (N_5333,N_4593,N_4992);
nand U5334 (N_5334,N_4063,N_4501);
nor U5335 (N_5335,N_4267,N_4289);
nand U5336 (N_5336,N_4443,N_4431);
nor U5337 (N_5337,N_4705,N_4697);
and U5338 (N_5338,N_4016,N_4977);
xnor U5339 (N_5339,N_4918,N_4339);
or U5340 (N_5340,N_4210,N_4369);
and U5341 (N_5341,N_4791,N_4873);
xnor U5342 (N_5342,N_4774,N_4570);
xor U5343 (N_5343,N_4119,N_4324);
and U5344 (N_5344,N_4149,N_4224);
or U5345 (N_5345,N_4396,N_4275);
nand U5346 (N_5346,N_4386,N_4408);
nor U5347 (N_5347,N_4807,N_4150);
nor U5348 (N_5348,N_4366,N_4839);
nand U5349 (N_5349,N_4979,N_4943);
nor U5350 (N_5350,N_4749,N_4522);
nor U5351 (N_5351,N_4309,N_4130);
xor U5352 (N_5352,N_4668,N_4880);
nor U5353 (N_5353,N_4700,N_4460);
xnor U5354 (N_5354,N_4045,N_4446);
nor U5355 (N_5355,N_4199,N_4136);
or U5356 (N_5356,N_4797,N_4208);
or U5357 (N_5357,N_4902,N_4789);
or U5358 (N_5358,N_4189,N_4318);
xor U5359 (N_5359,N_4400,N_4798);
or U5360 (N_5360,N_4319,N_4259);
xor U5361 (N_5361,N_4340,N_4089);
or U5362 (N_5362,N_4752,N_4039);
nor U5363 (N_5363,N_4245,N_4173);
nand U5364 (N_5364,N_4748,N_4314);
and U5365 (N_5365,N_4879,N_4345);
or U5366 (N_5366,N_4796,N_4773);
or U5367 (N_5367,N_4601,N_4521);
or U5368 (N_5368,N_4908,N_4568);
nor U5369 (N_5369,N_4279,N_4850);
and U5370 (N_5370,N_4656,N_4915);
xor U5371 (N_5371,N_4665,N_4286);
nor U5372 (N_5372,N_4590,N_4065);
nand U5373 (N_5373,N_4517,N_4759);
or U5374 (N_5374,N_4667,N_4008);
nand U5375 (N_5375,N_4263,N_4497);
xor U5376 (N_5376,N_4604,N_4254);
or U5377 (N_5377,N_4675,N_4467);
nand U5378 (N_5378,N_4139,N_4364);
and U5379 (N_5379,N_4076,N_4722);
nand U5380 (N_5380,N_4477,N_4241);
xor U5381 (N_5381,N_4876,N_4035);
nor U5382 (N_5382,N_4984,N_4028);
and U5383 (N_5383,N_4670,N_4101);
nor U5384 (N_5384,N_4354,N_4479);
nor U5385 (N_5385,N_4351,N_4491);
or U5386 (N_5386,N_4951,N_4800);
nand U5387 (N_5387,N_4132,N_4878);
or U5388 (N_5388,N_4886,N_4394);
or U5389 (N_5389,N_4882,N_4571);
nor U5390 (N_5390,N_4994,N_4105);
and U5391 (N_5391,N_4026,N_4982);
nor U5392 (N_5392,N_4504,N_4928);
nor U5393 (N_5393,N_4439,N_4499);
and U5394 (N_5394,N_4353,N_4037);
and U5395 (N_5395,N_4301,N_4110);
and U5396 (N_5396,N_4379,N_4135);
and U5397 (N_5397,N_4547,N_4234);
nor U5398 (N_5398,N_4300,N_4036);
and U5399 (N_5399,N_4837,N_4534);
xor U5400 (N_5400,N_4831,N_4652);
xnor U5401 (N_5401,N_4209,N_4525);
and U5402 (N_5402,N_4426,N_4213);
nor U5403 (N_5403,N_4610,N_4608);
and U5404 (N_5404,N_4603,N_4790);
xor U5405 (N_5405,N_4877,N_4930);
or U5406 (N_5406,N_4946,N_4727);
and U5407 (N_5407,N_4017,N_4191);
xnor U5408 (N_5408,N_4772,N_4739);
nand U5409 (N_5409,N_4165,N_4142);
and U5410 (N_5410,N_4128,N_4731);
or U5411 (N_5411,N_4333,N_4024);
or U5412 (N_5412,N_4859,N_4958);
nor U5413 (N_5413,N_4660,N_4761);
nor U5414 (N_5414,N_4485,N_4115);
xor U5415 (N_5415,N_4589,N_4531);
or U5416 (N_5416,N_4459,N_4561);
and U5417 (N_5417,N_4661,N_4600);
nor U5418 (N_5418,N_4047,N_4107);
and U5419 (N_5419,N_4628,N_4762);
nor U5420 (N_5420,N_4851,N_4738);
xor U5421 (N_5421,N_4703,N_4691);
nor U5422 (N_5422,N_4078,N_4900);
nor U5423 (N_5423,N_4729,N_4002);
xor U5424 (N_5424,N_4770,N_4311);
or U5425 (N_5425,N_4735,N_4331);
nor U5426 (N_5426,N_4757,N_4381);
or U5427 (N_5427,N_4468,N_4799);
or U5428 (N_5428,N_4975,N_4317);
and U5429 (N_5429,N_4053,N_4357);
nand U5430 (N_5430,N_4344,N_4724);
and U5431 (N_5431,N_4186,N_4023);
nor U5432 (N_5432,N_4437,N_4258);
and U5433 (N_5433,N_4163,N_4828);
and U5434 (N_5434,N_4125,N_4862);
and U5435 (N_5435,N_4056,N_4356);
xnor U5436 (N_5436,N_4613,N_4506);
and U5437 (N_5437,N_4503,N_4709);
nor U5438 (N_5438,N_4230,N_4206);
and U5439 (N_5439,N_4581,N_4161);
nor U5440 (N_5440,N_4681,N_4385);
and U5441 (N_5441,N_4544,N_4250);
or U5442 (N_5442,N_4393,N_4874);
or U5443 (N_5443,N_4630,N_4118);
nor U5444 (N_5444,N_4815,N_4572);
nand U5445 (N_5445,N_4276,N_4153);
xor U5446 (N_5446,N_4852,N_4693);
nor U5447 (N_5447,N_4392,N_4654);
and U5448 (N_5448,N_4763,N_4257);
xnor U5449 (N_5449,N_4043,N_4178);
or U5450 (N_5450,N_4524,N_4277);
xnor U5451 (N_5451,N_4417,N_4535);
and U5452 (N_5452,N_4252,N_4484);
and U5453 (N_5453,N_4845,N_4716);
nand U5454 (N_5454,N_4450,N_4162);
nor U5455 (N_5455,N_4883,N_4031);
nor U5456 (N_5456,N_4395,N_4231);
xor U5457 (N_5457,N_4449,N_4177);
or U5458 (N_5458,N_4302,N_4598);
xor U5459 (N_5459,N_4019,N_4100);
nand U5460 (N_5460,N_4292,N_4358);
nand U5461 (N_5461,N_4174,N_4148);
nand U5462 (N_5462,N_4753,N_4222);
nand U5463 (N_5463,N_4321,N_4332);
xor U5464 (N_5464,N_4680,N_4897);
xnor U5465 (N_5465,N_4622,N_4011);
and U5466 (N_5466,N_4769,N_4575);
nand U5467 (N_5467,N_4274,N_4972);
nor U5468 (N_5468,N_4646,N_4246);
nand U5469 (N_5469,N_4543,N_4272);
and U5470 (N_5470,N_4066,N_4347);
and U5471 (N_5471,N_4376,N_4040);
nor U5472 (N_5472,N_4623,N_4988);
nor U5473 (N_5473,N_4624,N_4320);
nor U5474 (N_5474,N_4853,N_4931);
xor U5475 (N_5475,N_4591,N_4755);
xor U5476 (N_5476,N_4614,N_4846);
or U5477 (N_5477,N_4212,N_4266);
or U5478 (N_5478,N_4875,N_4954);
nor U5479 (N_5479,N_4549,N_4911);
xnor U5480 (N_5480,N_4126,N_4921);
nor U5481 (N_5481,N_4919,N_4048);
nand U5482 (N_5482,N_4903,N_4582);
or U5483 (N_5483,N_4134,N_4441);
nand U5484 (N_5484,N_4564,N_4159);
and U5485 (N_5485,N_4557,N_4981);
and U5486 (N_5486,N_4938,N_4960);
and U5487 (N_5487,N_4856,N_4701);
nor U5488 (N_5488,N_4423,N_4803);
and U5489 (N_5489,N_4664,N_4580);
nor U5490 (N_5490,N_4780,N_4987);
nand U5491 (N_5491,N_4232,N_4419);
or U5492 (N_5492,N_4004,N_4221);
nand U5493 (N_5493,N_4095,N_4032);
and U5494 (N_5494,N_4341,N_4810);
and U5495 (N_5495,N_4336,N_4847);
nand U5496 (N_5496,N_4971,N_4143);
nand U5497 (N_5497,N_4197,N_4945);
nor U5498 (N_5498,N_4658,N_4889);
and U5499 (N_5499,N_4817,N_4424);
and U5500 (N_5500,N_4726,N_4437);
or U5501 (N_5501,N_4428,N_4364);
nor U5502 (N_5502,N_4930,N_4434);
or U5503 (N_5503,N_4007,N_4894);
nor U5504 (N_5504,N_4188,N_4961);
or U5505 (N_5505,N_4170,N_4949);
and U5506 (N_5506,N_4083,N_4329);
xor U5507 (N_5507,N_4519,N_4696);
or U5508 (N_5508,N_4348,N_4671);
or U5509 (N_5509,N_4312,N_4434);
or U5510 (N_5510,N_4750,N_4290);
or U5511 (N_5511,N_4243,N_4610);
and U5512 (N_5512,N_4359,N_4574);
xnor U5513 (N_5513,N_4339,N_4635);
and U5514 (N_5514,N_4665,N_4888);
nor U5515 (N_5515,N_4505,N_4627);
nor U5516 (N_5516,N_4688,N_4276);
nand U5517 (N_5517,N_4904,N_4957);
xor U5518 (N_5518,N_4968,N_4569);
nand U5519 (N_5519,N_4174,N_4252);
or U5520 (N_5520,N_4363,N_4222);
xor U5521 (N_5521,N_4871,N_4576);
or U5522 (N_5522,N_4264,N_4281);
xor U5523 (N_5523,N_4192,N_4389);
nand U5524 (N_5524,N_4096,N_4603);
and U5525 (N_5525,N_4481,N_4389);
nor U5526 (N_5526,N_4696,N_4537);
xnor U5527 (N_5527,N_4945,N_4653);
nand U5528 (N_5528,N_4362,N_4444);
nor U5529 (N_5529,N_4989,N_4004);
xor U5530 (N_5530,N_4609,N_4229);
and U5531 (N_5531,N_4159,N_4186);
nor U5532 (N_5532,N_4292,N_4877);
nor U5533 (N_5533,N_4489,N_4422);
and U5534 (N_5534,N_4860,N_4322);
nor U5535 (N_5535,N_4987,N_4459);
xnor U5536 (N_5536,N_4535,N_4008);
nor U5537 (N_5537,N_4915,N_4737);
nor U5538 (N_5538,N_4689,N_4885);
nand U5539 (N_5539,N_4155,N_4017);
and U5540 (N_5540,N_4291,N_4833);
xnor U5541 (N_5541,N_4911,N_4860);
or U5542 (N_5542,N_4442,N_4124);
nor U5543 (N_5543,N_4926,N_4042);
or U5544 (N_5544,N_4153,N_4795);
nor U5545 (N_5545,N_4959,N_4996);
nand U5546 (N_5546,N_4263,N_4651);
xnor U5547 (N_5547,N_4090,N_4797);
or U5548 (N_5548,N_4523,N_4197);
nor U5549 (N_5549,N_4831,N_4393);
and U5550 (N_5550,N_4953,N_4062);
xnor U5551 (N_5551,N_4226,N_4770);
nor U5552 (N_5552,N_4322,N_4242);
nor U5553 (N_5553,N_4652,N_4835);
or U5554 (N_5554,N_4641,N_4078);
nor U5555 (N_5555,N_4813,N_4307);
or U5556 (N_5556,N_4326,N_4968);
or U5557 (N_5557,N_4146,N_4501);
and U5558 (N_5558,N_4919,N_4702);
or U5559 (N_5559,N_4635,N_4205);
nor U5560 (N_5560,N_4351,N_4232);
or U5561 (N_5561,N_4095,N_4903);
and U5562 (N_5562,N_4422,N_4043);
nand U5563 (N_5563,N_4058,N_4804);
or U5564 (N_5564,N_4980,N_4906);
xor U5565 (N_5565,N_4153,N_4435);
nor U5566 (N_5566,N_4152,N_4884);
nor U5567 (N_5567,N_4668,N_4591);
nor U5568 (N_5568,N_4463,N_4251);
xnor U5569 (N_5569,N_4705,N_4323);
or U5570 (N_5570,N_4651,N_4020);
nand U5571 (N_5571,N_4406,N_4476);
and U5572 (N_5572,N_4936,N_4450);
and U5573 (N_5573,N_4953,N_4494);
and U5574 (N_5574,N_4692,N_4415);
nor U5575 (N_5575,N_4178,N_4524);
nand U5576 (N_5576,N_4001,N_4318);
nor U5577 (N_5577,N_4444,N_4159);
and U5578 (N_5578,N_4469,N_4968);
and U5579 (N_5579,N_4375,N_4622);
nand U5580 (N_5580,N_4934,N_4919);
nand U5581 (N_5581,N_4883,N_4872);
and U5582 (N_5582,N_4379,N_4985);
or U5583 (N_5583,N_4022,N_4842);
and U5584 (N_5584,N_4835,N_4572);
or U5585 (N_5585,N_4532,N_4157);
nand U5586 (N_5586,N_4282,N_4185);
nand U5587 (N_5587,N_4981,N_4735);
nor U5588 (N_5588,N_4341,N_4777);
xnor U5589 (N_5589,N_4100,N_4509);
xor U5590 (N_5590,N_4442,N_4918);
xor U5591 (N_5591,N_4571,N_4654);
nand U5592 (N_5592,N_4541,N_4373);
nor U5593 (N_5593,N_4278,N_4026);
or U5594 (N_5594,N_4797,N_4976);
xnor U5595 (N_5595,N_4599,N_4426);
nand U5596 (N_5596,N_4588,N_4814);
and U5597 (N_5597,N_4996,N_4407);
xnor U5598 (N_5598,N_4862,N_4056);
and U5599 (N_5599,N_4685,N_4307);
xor U5600 (N_5600,N_4682,N_4040);
nor U5601 (N_5601,N_4787,N_4328);
or U5602 (N_5602,N_4578,N_4939);
or U5603 (N_5603,N_4613,N_4333);
xor U5604 (N_5604,N_4941,N_4009);
and U5605 (N_5605,N_4969,N_4487);
xor U5606 (N_5606,N_4152,N_4721);
or U5607 (N_5607,N_4499,N_4303);
nand U5608 (N_5608,N_4411,N_4457);
nand U5609 (N_5609,N_4700,N_4823);
nand U5610 (N_5610,N_4242,N_4272);
nor U5611 (N_5611,N_4903,N_4692);
nand U5612 (N_5612,N_4202,N_4860);
or U5613 (N_5613,N_4518,N_4626);
nand U5614 (N_5614,N_4111,N_4081);
and U5615 (N_5615,N_4618,N_4390);
xor U5616 (N_5616,N_4192,N_4810);
nand U5617 (N_5617,N_4139,N_4677);
nor U5618 (N_5618,N_4637,N_4041);
or U5619 (N_5619,N_4485,N_4514);
nor U5620 (N_5620,N_4619,N_4457);
nand U5621 (N_5621,N_4640,N_4795);
nor U5622 (N_5622,N_4417,N_4856);
or U5623 (N_5623,N_4191,N_4913);
or U5624 (N_5624,N_4783,N_4206);
xnor U5625 (N_5625,N_4788,N_4656);
or U5626 (N_5626,N_4712,N_4858);
and U5627 (N_5627,N_4900,N_4215);
nor U5628 (N_5628,N_4793,N_4585);
xnor U5629 (N_5629,N_4096,N_4502);
nand U5630 (N_5630,N_4170,N_4482);
and U5631 (N_5631,N_4336,N_4004);
nor U5632 (N_5632,N_4268,N_4780);
and U5633 (N_5633,N_4054,N_4258);
and U5634 (N_5634,N_4359,N_4947);
nand U5635 (N_5635,N_4053,N_4240);
xnor U5636 (N_5636,N_4148,N_4318);
nor U5637 (N_5637,N_4913,N_4649);
nand U5638 (N_5638,N_4760,N_4978);
nor U5639 (N_5639,N_4545,N_4205);
and U5640 (N_5640,N_4939,N_4002);
xnor U5641 (N_5641,N_4923,N_4897);
nand U5642 (N_5642,N_4761,N_4273);
nand U5643 (N_5643,N_4012,N_4695);
nor U5644 (N_5644,N_4616,N_4280);
and U5645 (N_5645,N_4224,N_4260);
or U5646 (N_5646,N_4637,N_4267);
and U5647 (N_5647,N_4782,N_4175);
and U5648 (N_5648,N_4342,N_4485);
nand U5649 (N_5649,N_4648,N_4800);
nand U5650 (N_5650,N_4740,N_4666);
nor U5651 (N_5651,N_4067,N_4538);
nor U5652 (N_5652,N_4553,N_4872);
and U5653 (N_5653,N_4633,N_4609);
nor U5654 (N_5654,N_4123,N_4867);
and U5655 (N_5655,N_4571,N_4360);
or U5656 (N_5656,N_4520,N_4476);
or U5657 (N_5657,N_4584,N_4423);
xnor U5658 (N_5658,N_4730,N_4603);
nand U5659 (N_5659,N_4448,N_4529);
xor U5660 (N_5660,N_4435,N_4708);
xor U5661 (N_5661,N_4590,N_4036);
nor U5662 (N_5662,N_4783,N_4976);
nor U5663 (N_5663,N_4111,N_4770);
or U5664 (N_5664,N_4216,N_4440);
or U5665 (N_5665,N_4293,N_4170);
nor U5666 (N_5666,N_4441,N_4462);
nor U5667 (N_5667,N_4604,N_4826);
or U5668 (N_5668,N_4082,N_4951);
nor U5669 (N_5669,N_4670,N_4568);
xnor U5670 (N_5670,N_4832,N_4147);
xor U5671 (N_5671,N_4411,N_4848);
nand U5672 (N_5672,N_4395,N_4155);
xnor U5673 (N_5673,N_4702,N_4145);
nand U5674 (N_5674,N_4789,N_4036);
nand U5675 (N_5675,N_4707,N_4339);
xnor U5676 (N_5676,N_4142,N_4337);
or U5677 (N_5677,N_4556,N_4968);
xnor U5678 (N_5678,N_4103,N_4994);
and U5679 (N_5679,N_4730,N_4302);
nor U5680 (N_5680,N_4526,N_4028);
xnor U5681 (N_5681,N_4375,N_4785);
nor U5682 (N_5682,N_4051,N_4598);
nand U5683 (N_5683,N_4347,N_4767);
or U5684 (N_5684,N_4488,N_4611);
nand U5685 (N_5685,N_4955,N_4264);
or U5686 (N_5686,N_4686,N_4173);
nand U5687 (N_5687,N_4114,N_4187);
nand U5688 (N_5688,N_4637,N_4260);
nand U5689 (N_5689,N_4862,N_4298);
and U5690 (N_5690,N_4553,N_4450);
and U5691 (N_5691,N_4497,N_4719);
nand U5692 (N_5692,N_4488,N_4427);
nand U5693 (N_5693,N_4128,N_4140);
nand U5694 (N_5694,N_4462,N_4001);
nand U5695 (N_5695,N_4903,N_4919);
xor U5696 (N_5696,N_4827,N_4660);
and U5697 (N_5697,N_4478,N_4074);
xnor U5698 (N_5698,N_4694,N_4402);
and U5699 (N_5699,N_4376,N_4440);
xor U5700 (N_5700,N_4573,N_4265);
or U5701 (N_5701,N_4460,N_4278);
or U5702 (N_5702,N_4408,N_4429);
nor U5703 (N_5703,N_4867,N_4138);
and U5704 (N_5704,N_4058,N_4278);
nand U5705 (N_5705,N_4844,N_4257);
nor U5706 (N_5706,N_4223,N_4612);
nand U5707 (N_5707,N_4636,N_4030);
nor U5708 (N_5708,N_4930,N_4542);
nor U5709 (N_5709,N_4818,N_4724);
or U5710 (N_5710,N_4240,N_4667);
or U5711 (N_5711,N_4118,N_4216);
nand U5712 (N_5712,N_4746,N_4485);
xnor U5713 (N_5713,N_4098,N_4503);
and U5714 (N_5714,N_4271,N_4255);
nor U5715 (N_5715,N_4647,N_4295);
or U5716 (N_5716,N_4656,N_4937);
or U5717 (N_5717,N_4428,N_4644);
or U5718 (N_5718,N_4318,N_4443);
or U5719 (N_5719,N_4871,N_4281);
nand U5720 (N_5720,N_4096,N_4014);
and U5721 (N_5721,N_4753,N_4579);
xor U5722 (N_5722,N_4219,N_4593);
or U5723 (N_5723,N_4883,N_4923);
or U5724 (N_5724,N_4674,N_4183);
nor U5725 (N_5725,N_4046,N_4164);
and U5726 (N_5726,N_4231,N_4279);
or U5727 (N_5727,N_4796,N_4511);
and U5728 (N_5728,N_4300,N_4583);
nand U5729 (N_5729,N_4753,N_4575);
nand U5730 (N_5730,N_4305,N_4579);
nor U5731 (N_5731,N_4042,N_4044);
xnor U5732 (N_5732,N_4229,N_4568);
or U5733 (N_5733,N_4441,N_4234);
xor U5734 (N_5734,N_4291,N_4911);
xor U5735 (N_5735,N_4977,N_4231);
nor U5736 (N_5736,N_4936,N_4954);
nor U5737 (N_5737,N_4574,N_4686);
nand U5738 (N_5738,N_4079,N_4350);
and U5739 (N_5739,N_4319,N_4727);
or U5740 (N_5740,N_4071,N_4176);
nor U5741 (N_5741,N_4500,N_4010);
and U5742 (N_5742,N_4131,N_4479);
or U5743 (N_5743,N_4364,N_4691);
nor U5744 (N_5744,N_4778,N_4172);
nor U5745 (N_5745,N_4779,N_4369);
xor U5746 (N_5746,N_4236,N_4898);
nand U5747 (N_5747,N_4490,N_4199);
and U5748 (N_5748,N_4077,N_4836);
or U5749 (N_5749,N_4565,N_4298);
or U5750 (N_5750,N_4925,N_4407);
and U5751 (N_5751,N_4194,N_4345);
and U5752 (N_5752,N_4998,N_4462);
and U5753 (N_5753,N_4053,N_4140);
and U5754 (N_5754,N_4925,N_4376);
or U5755 (N_5755,N_4897,N_4242);
or U5756 (N_5756,N_4394,N_4175);
xnor U5757 (N_5757,N_4140,N_4534);
or U5758 (N_5758,N_4277,N_4981);
and U5759 (N_5759,N_4692,N_4197);
or U5760 (N_5760,N_4097,N_4241);
xnor U5761 (N_5761,N_4988,N_4215);
nand U5762 (N_5762,N_4743,N_4639);
nand U5763 (N_5763,N_4958,N_4197);
or U5764 (N_5764,N_4325,N_4016);
nor U5765 (N_5765,N_4619,N_4085);
or U5766 (N_5766,N_4691,N_4540);
xnor U5767 (N_5767,N_4280,N_4287);
or U5768 (N_5768,N_4617,N_4038);
nor U5769 (N_5769,N_4546,N_4577);
and U5770 (N_5770,N_4903,N_4334);
and U5771 (N_5771,N_4442,N_4749);
and U5772 (N_5772,N_4684,N_4133);
and U5773 (N_5773,N_4350,N_4130);
xnor U5774 (N_5774,N_4787,N_4107);
nor U5775 (N_5775,N_4045,N_4784);
nor U5776 (N_5776,N_4034,N_4412);
or U5777 (N_5777,N_4992,N_4225);
or U5778 (N_5778,N_4186,N_4045);
nor U5779 (N_5779,N_4831,N_4780);
nor U5780 (N_5780,N_4253,N_4354);
and U5781 (N_5781,N_4788,N_4271);
xnor U5782 (N_5782,N_4312,N_4472);
and U5783 (N_5783,N_4310,N_4629);
or U5784 (N_5784,N_4967,N_4812);
nand U5785 (N_5785,N_4590,N_4723);
nand U5786 (N_5786,N_4527,N_4250);
or U5787 (N_5787,N_4955,N_4966);
or U5788 (N_5788,N_4555,N_4539);
or U5789 (N_5789,N_4162,N_4814);
nor U5790 (N_5790,N_4031,N_4334);
nand U5791 (N_5791,N_4391,N_4536);
xnor U5792 (N_5792,N_4663,N_4757);
and U5793 (N_5793,N_4496,N_4820);
nand U5794 (N_5794,N_4786,N_4267);
and U5795 (N_5795,N_4240,N_4387);
xnor U5796 (N_5796,N_4239,N_4846);
nand U5797 (N_5797,N_4222,N_4832);
nor U5798 (N_5798,N_4251,N_4932);
nand U5799 (N_5799,N_4868,N_4841);
xnor U5800 (N_5800,N_4447,N_4023);
xor U5801 (N_5801,N_4176,N_4971);
nand U5802 (N_5802,N_4276,N_4085);
xor U5803 (N_5803,N_4999,N_4308);
or U5804 (N_5804,N_4561,N_4575);
and U5805 (N_5805,N_4434,N_4234);
nor U5806 (N_5806,N_4977,N_4560);
nor U5807 (N_5807,N_4981,N_4081);
or U5808 (N_5808,N_4407,N_4135);
nand U5809 (N_5809,N_4032,N_4565);
or U5810 (N_5810,N_4262,N_4072);
nor U5811 (N_5811,N_4933,N_4938);
nand U5812 (N_5812,N_4130,N_4854);
nand U5813 (N_5813,N_4146,N_4325);
or U5814 (N_5814,N_4597,N_4955);
nand U5815 (N_5815,N_4416,N_4509);
nor U5816 (N_5816,N_4971,N_4679);
nor U5817 (N_5817,N_4777,N_4439);
xnor U5818 (N_5818,N_4435,N_4810);
and U5819 (N_5819,N_4427,N_4872);
or U5820 (N_5820,N_4171,N_4298);
nand U5821 (N_5821,N_4306,N_4676);
nand U5822 (N_5822,N_4549,N_4968);
and U5823 (N_5823,N_4326,N_4451);
nor U5824 (N_5824,N_4098,N_4398);
or U5825 (N_5825,N_4373,N_4811);
nor U5826 (N_5826,N_4879,N_4547);
and U5827 (N_5827,N_4015,N_4505);
nand U5828 (N_5828,N_4346,N_4320);
nand U5829 (N_5829,N_4553,N_4856);
and U5830 (N_5830,N_4989,N_4327);
or U5831 (N_5831,N_4756,N_4681);
nor U5832 (N_5832,N_4923,N_4059);
nand U5833 (N_5833,N_4209,N_4435);
and U5834 (N_5834,N_4881,N_4183);
nand U5835 (N_5835,N_4675,N_4744);
and U5836 (N_5836,N_4109,N_4253);
nor U5837 (N_5837,N_4018,N_4377);
nor U5838 (N_5838,N_4954,N_4683);
nor U5839 (N_5839,N_4311,N_4680);
xor U5840 (N_5840,N_4533,N_4428);
or U5841 (N_5841,N_4485,N_4314);
and U5842 (N_5842,N_4550,N_4495);
or U5843 (N_5843,N_4672,N_4885);
nand U5844 (N_5844,N_4687,N_4537);
nand U5845 (N_5845,N_4214,N_4391);
nor U5846 (N_5846,N_4144,N_4043);
nand U5847 (N_5847,N_4324,N_4552);
nand U5848 (N_5848,N_4119,N_4589);
nor U5849 (N_5849,N_4660,N_4403);
or U5850 (N_5850,N_4303,N_4348);
xnor U5851 (N_5851,N_4004,N_4550);
xor U5852 (N_5852,N_4982,N_4358);
xnor U5853 (N_5853,N_4074,N_4131);
nand U5854 (N_5854,N_4276,N_4997);
or U5855 (N_5855,N_4490,N_4262);
and U5856 (N_5856,N_4685,N_4101);
nor U5857 (N_5857,N_4578,N_4989);
and U5858 (N_5858,N_4854,N_4057);
or U5859 (N_5859,N_4973,N_4009);
or U5860 (N_5860,N_4797,N_4463);
and U5861 (N_5861,N_4002,N_4629);
and U5862 (N_5862,N_4177,N_4674);
xor U5863 (N_5863,N_4399,N_4259);
nor U5864 (N_5864,N_4623,N_4532);
and U5865 (N_5865,N_4287,N_4435);
and U5866 (N_5866,N_4510,N_4141);
and U5867 (N_5867,N_4622,N_4350);
xnor U5868 (N_5868,N_4798,N_4460);
xnor U5869 (N_5869,N_4856,N_4089);
and U5870 (N_5870,N_4960,N_4634);
nor U5871 (N_5871,N_4810,N_4168);
and U5872 (N_5872,N_4889,N_4722);
nor U5873 (N_5873,N_4829,N_4317);
xor U5874 (N_5874,N_4803,N_4712);
or U5875 (N_5875,N_4980,N_4978);
or U5876 (N_5876,N_4109,N_4928);
xnor U5877 (N_5877,N_4145,N_4307);
or U5878 (N_5878,N_4099,N_4217);
and U5879 (N_5879,N_4186,N_4886);
nor U5880 (N_5880,N_4174,N_4661);
and U5881 (N_5881,N_4054,N_4196);
or U5882 (N_5882,N_4266,N_4936);
nor U5883 (N_5883,N_4344,N_4726);
or U5884 (N_5884,N_4577,N_4398);
nor U5885 (N_5885,N_4172,N_4656);
nand U5886 (N_5886,N_4275,N_4126);
and U5887 (N_5887,N_4272,N_4336);
nand U5888 (N_5888,N_4471,N_4886);
xnor U5889 (N_5889,N_4982,N_4661);
and U5890 (N_5890,N_4040,N_4997);
xor U5891 (N_5891,N_4203,N_4081);
nor U5892 (N_5892,N_4263,N_4523);
nand U5893 (N_5893,N_4276,N_4087);
nand U5894 (N_5894,N_4721,N_4677);
nand U5895 (N_5895,N_4458,N_4634);
xnor U5896 (N_5896,N_4957,N_4279);
and U5897 (N_5897,N_4393,N_4108);
xor U5898 (N_5898,N_4416,N_4949);
and U5899 (N_5899,N_4732,N_4604);
and U5900 (N_5900,N_4864,N_4013);
xnor U5901 (N_5901,N_4354,N_4102);
nor U5902 (N_5902,N_4426,N_4061);
nand U5903 (N_5903,N_4589,N_4745);
and U5904 (N_5904,N_4302,N_4915);
nor U5905 (N_5905,N_4864,N_4250);
xor U5906 (N_5906,N_4126,N_4082);
nand U5907 (N_5907,N_4942,N_4820);
xnor U5908 (N_5908,N_4089,N_4065);
xnor U5909 (N_5909,N_4408,N_4622);
xnor U5910 (N_5910,N_4381,N_4278);
nor U5911 (N_5911,N_4978,N_4224);
and U5912 (N_5912,N_4623,N_4599);
or U5913 (N_5913,N_4416,N_4901);
xor U5914 (N_5914,N_4498,N_4982);
and U5915 (N_5915,N_4687,N_4569);
and U5916 (N_5916,N_4321,N_4916);
xor U5917 (N_5917,N_4686,N_4619);
xnor U5918 (N_5918,N_4531,N_4710);
nor U5919 (N_5919,N_4339,N_4721);
or U5920 (N_5920,N_4698,N_4740);
and U5921 (N_5921,N_4096,N_4963);
and U5922 (N_5922,N_4344,N_4682);
nand U5923 (N_5923,N_4383,N_4832);
or U5924 (N_5924,N_4958,N_4573);
xor U5925 (N_5925,N_4574,N_4376);
xor U5926 (N_5926,N_4578,N_4848);
xor U5927 (N_5927,N_4694,N_4720);
xor U5928 (N_5928,N_4466,N_4930);
or U5929 (N_5929,N_4308,N_4650);
and U5930 (N_5930,N_4702,N_4322);
or U5931 (N_5931,N_4789,N_4931);
nand U5932 (N_5932,N_4323,N_4779);
nor U5933 (N_5933,N_4811,N_4049);
nor U5934 (N_5934,N_4348,N_4485);
or U5935 (N_5935,N_4929,N_4272);
nor U5936 (N_5936,N_4865,N_4346);
xnor U5937 (N_5937,N_4550,N_4363);
nor U5938 (N_5938,N_4410,N_4695);
or U5939 (N_5939,N_4642,N_4389);
nand U5940 (N_5940,N_4378,N_4138);
xor U5941 (N_5941,N_4502,N_4284);
and U5942 (N_5942,N_4560,N_4953);
xnor U5943 (N_5943,N_4944,N_4070);
nor U5944 (N_5944,N_4561,N_4581);
and U5945 (N_5945,N_4646,N_4052);
or U5946 (N_5946,N_4922,N_4265);
nand U5947 (N_5947,N_4966,N_4798);
nor U5948 (N_5948,N_4988,N_4336);
nand U5949 (N_5949,N_4833,N_4721);
nor U5950 (N_5950,N_4484,N_4468);
nor U5951 (N_5951,N_4524,N_4570);
xnor U5952 (N_5952,N_4545,N_4808);
xnor U5953 (N_5953,N_4493,N_4242);
nand U5954 (N_5954,N_4218,N_4437);
nor U5955 (N_5955,N_4656,N_4541);
or U5956 (N_5956,N_4202,N_4496);
and U5957 (N_5957,N_4240,N_4047);
xor U5958 (N_5958,N_4174,N_4197);
or U5959 (N_5959,N_4764,N_4954);
nor U5960 (N_5960,N_4713,N_4972);
and U5961 (N_5961,N_4747,N_4946);
or U5962 (N_5962,N_4409,N_4422);
nor U5963 (N_5963,N_4860,N_4997);
and U5964 (N_5964,N_4118,N_4700);
nor U5965 (N_5965,N_4381,N_4627);
xnor U5966 (N_5966,N_4649,N_4872);
nor U5967 (N_5967,N_4556,N_4862);
and U5968 (N_5968,N_4089,N_4611);
nor U5969 (N_5969,N_4286,N_4106);
and U5970 (N_5970,N_4895,N_4327);
nor U5971 (N_5971,N_4632,N_4058);
nand U5972 (N_5972,N_4236,N_4970);
or U5973 (N_5973,N_4663,N_4427);
nor U5974 (N_5974,N_4102,N_4848);
or U5975 (N_5975,N_4406,N_4997);
nor U5976 (N_5976,N_4305,N_4472);
or U5977 (N_5977,N_4367,N_4983);
or U5978 (N_5978,N_4527,N_4489);
or U5979 (N_5979,N_4035,N_4731);
nand U5980 (N_5980,N_4941,N_4763);
nand U5981 (N_5981,N_4463,N_4219);
nor U5982 (N_5982,N_4747,N_4232);
xor U5983 (N_5983,N_4491,N_4800);
nand U5984 (N_5984,N_4182,N_4409);
or U5985 (N_5985,N_4159,N_4920);
nor U5986 (N_5986,N_4277,N_4502);
and U5987 (N_5987,N_4896,N_4685);
nand U5988 (N_5988,N_4896,N_4659);
or U5989 (N_5989,N_4624,N_4755);
or U5990 (N_5990,N_4040,N_4029);
nand U5991 (N_5991,N_4129,N_4119);
and U5992 (N_5992,N_4870,N_4863);
nand U5993 (N_5993,N_4238,N_4132);
and U5994 (N_5994,N_4224,N_4451);
nand U5995 (N_5995,N_4295,N_4974);
or U5996 (N_5996,N_4537,N_4677);
nor U5997 (N_5997,N_4863,N_4577);
and U5998 (N_5998,N_4899,N_4398);
nor U5999 (N_5999,N_4568,N_4967);
and U6000 (N_6000,N_5301,N_5785);
xnor U6001 (N_6001,N_5286,N_5590);
nor U6002 (N_6002,N_5652,N_5223);
nand U6003 (N_6003,N_5791,N_5458);
xnor U6004 (N_6004,N_5868,N_5125);
nand U6005 (N_6005,N_5327,N_5550);
nand U6006 (N_6006,N_5631,N_5807);
nor U6007 (N_6007,N_5692,N_5004);
or U6008 (N_6008,N_5073,N_5849);
xor U6009 (N_6009,N_5872,N_5480);
or U6010 (N_6010,N_5099,N_5437);
or U6011 (N_6011,N_5822,N_5472);
xnor U6012 (N_6012,N_5473,N_5593);
xnor U6013 (N_6013,N_5463,N_5840);
xnor U6014 (N_6014,N_5922,N_5216);
or U6015 (N_6015,N_5426,N_5093);
nand U6016 (N_6016,N_5964,N_5890);
and U6017 (N_6017,N_5324,N_5398);
or U6018 (N_6018,N_5723,N_5674);
or U6019 (N_6019,N_5450,N_5748);
nor U6020 (N_6020,N_5848,N_5756);
nor U6021 (N_6021,N_5635,N_5132);
nor U6022 (N_6022,N_5534,N_5335);
nor U6023 (N_6023,N_5678,N_5016);
nand U6024 (N_6024,N_5133,N_5864);
nor U6025 (N_6025,N_5177,N_5957);
and U6026 (N_6026,N_5955,N_5241);
or U6027 (N_6027,N_5483,N_5516);
xor U6028 (N_6028,N_5414,N_5570);
nor U6029 (N_6029,N_5660,N_5384);
and U6030 (N_6030,N_5992,N_5420);
or U6031 (N_6031,N_5449,N_5110);
nor U6032 (N_6032,N_5743,N_5305);
nand U6033 (N_6033,N_5968,N_5396);
or U6034 (N_6034,N_5428,N_5982);
nor U6035 (N_6035,N_5148,N_5834);
xor U6036 (N_6036,N_5230,N_5271);
nand U6037 (N_6037,N_5724,N_5017);
nor U6038 (N_6038,N_5369,N_5543);
or U6039 (N_6039,N_5841,N_5075);
nand U6040 (N_6040,N_5364,N_5972);
and U6041 (N_6041,N_5595,N_5039);
and U6042 (N_6042,N_5994,N_5047);
and U6043 (N_6043,N_5060,N_5180);
nor U6044 (N_6044,N_5893,N_5446);
xnor U6045 (N_6045,N_5354,N_5197);
and U6046 (N_6046,N_5086,N_5330);
xnor U6047 (N_6047,N_5325,N_5014);
and U6048 (N_6048,N_5510,N_5627);
and U6049 (N_6049,N_5626,N_5676);
nor U6050 (N_6050,N_5439,N_5290);
and U6051 (N_6051,N_5211,N_5936);
or U6052 (N_6052,N_5779,N_5466);
or U6053 (N_6053,N_5235,N_5094);
nor U6054 (N_6054,N_5602,N_5080);
nand U6055 (N_6055,N_5622,N_5255);
xnor U6056 (N_6056,N_5798,N_5797);
nor U6057 (N_6057,N_5373,N_5642);
xor U6058 (N_6058,N_5481,N_5068);
nand U6059 (N_6059,N_5173,N_5682);
or U6060 (N_6060,N_5368,N_5783);
and U6061 (N_6061,N_5708,N_5826);
nor U6062 (N_6062,N_5636,N_5076);
nand U6063 (N_6063,N_5924,N_5781);
and U6064 (N_6064,N_5045,N_5530);
xnor U6065 (N_6065,N_5202,N_5730);
or U6066 (N_6066,N_5453,N_5320);
or U6067 (N_6067,N_5342,N_5009);
or U6068 (N_6068,N_5587,N_5239);
or U6069 (N_6069,N_5338,N_5888);
nor U6070 (N_6070,N_5742,N_5336);
and U6071 (N_6071,N_5619,N_5894);
or U6072 (N_6072,N_5242,N_5511);
nand U6073 (N_6073,N_5668,N_5013);
or U6074 (N_6074,N_5965,N_5171);
nor U6075 (N_6075,N_5529,N_5859);
or U6076 (N_6076,N_5599,N_5489);
nand U6077 (N_6077,N_5140,N_5650);
xnor U6078 (N_6078,N_5119,N_5738);
nand U6079 (N_6079,N_5792,N_5991);
xnor U6080 (N_6080,N_5700,N_5699);
and U6081 (N_6081,N_5467,N_5865);
or U6082 (N_6082,N_5405,N_5808);
or U6083 (N_6083,N_5139,N_5270);
nor U6084 (N_6084,N_5159,N_5763);
nor U6085 (N_6085,N_5664,N_5088);
or U6086 (N_6086,N_5525,N_5617);
nor U6087 (N_6087,N_5918,N_5208);
nor U6088 (N_6088,N_5415,N_5777);
nand U6089 (N_6089,N_5934,N_5735);
xor U6090 (N_6090,N_5395,N_5215);
and U6091 (N_6091,N_5332,N_5609);
and U6092 (N_6092,N_5624,N_5565);
nand U6093 (N_6093,N_5401,N_5112);
or U6094 (N_6094,N_5329,N_5331);
xor U6095 (N_6095,N_5447,N_5015);
xnor U6096 (N_6096,N_5657,N_5632);
nand U6097 (N_6097,N_5572,N_5434);
nor U6098 (N_6098,N_5438,N_5656);
nor U6099 (N_6099,N_5800,N_5000);
xnor U6100 (N_6100,N_5248,N_5302);
nand U6101 (N_6101,N_5231,N_5750);
nor U6102 (N_6102,N_5578,N_5718);
nand U6103 (N_6103,N_5513,N_5031);
or U6104 (N_6104,N_5263,N_5873);
nor U6105 (N_6105,N_5498,N_5705);
nand U6106 (N_6106,N_5028,N_5561);
and U6107 (N_6107,N_5986,N_5853);
and U6108 (N_6108,N_5928,N_5633);
or U6109 (N_6109,N_5034,N_5860);
xnor U6110 (N_6110,N_5704,N_5200);
and U6111 (N_6111,N_5448,N_5930);
and U6112 (N_6112,N_5461,N_5470);
nand U6113 (N_6113,N_5575,N_5973);
or U6114 (N_6114,N_5985,N_5388);
or U6115 (N_6115,N_5341,N_5240);
or U6116 (N_6116,N_5588,N_5762);
nand U6117 (N_6117,N_5616,N_5107);
nand U6118 (N_6118,N_5646,N_5612);
and U6119 (N_6119,N_5983,N_5751);
nor U6120 (N_6120,N_5683,N_5950);
xor U6121 (N_6121,N_5829,N_5024);
nor U6122 (N_6122,N_5558,N_5328);
nor U6123 (N_6123,N_5431,N_5417);
xnor U6124 (N_6124,N_5547,N_5693);
nand U6125 (N_6125,N_5036,N_5711);
xnor U6126 (N_6126,N_5179,N_5085);
or U6127 (N_6127,N_5217,N_5397);
xor U6128 (N_6128,N_5025,N_5352);
xnor U6129 (N_6129,N_5831,N_5541);
and U6130 (N_6130,N_5882,N_5318);
nand U6131 (N_6131,N_5908,N_5677);
or U6132 (N_6132,N_5939,N_5451);
nor U6133 (N_6133,N_5725,N_5518);
or U6134 (N_6134,N_5929,N_5412);
xnor U6135 (N_6135,N_5247,N_5694);
nor U6136 (N_6136,N_5280,N_5746);
nor U6137 (N_6137,N_5687,N_5672);
nand U6138 (N_6138,N_5820,N_5213);
nand U6139 (N_6139,N_5106,N_5596);
nor U6140 (N_6140,N_5760,N_5390);
and U6141 (N_6141,N_5050,N_5297);
nor U6142 (N_6142,N_5287,N_5926);
or U6143 (N_6143,N_5204,N_5351);
nor U6144 (N_6144,N_5744,N_5382);
xor U6145 (N_6145,N_5527,N_5251);
nor U6146 (N_6146,N_5847,N_5193);
xnor U6147 (N_6147,N_5167,N_5460);
xor U6148 (N_6148,N_5150,N_5755);
or U6149 (N_6149,N_5313,N_5101);
nand U6150 (N_6150,N_5224,N_5921);
or U6151 (N_6151,N_5361,N_5374);
xnor U6152 (N_6152,N_5089,N_5257);
nor U6153 (N_6153,N_5192,N_5147);
or U6154 (N_6154,N_5126,N_5933);
nand U6155 (N_6155,N_5274,N_5563);
nor U6156 (N_6156,N_5471,N_5372);
xnor U6157 (N_6157,N_5038,N_5468);
xor U6158 (N_6158,N_5355,N_5772);
nor U6159 (N_6159,N_5589,N_5761);
nand U6160 (N_6160,N_5515,N_5090);
xor U6161 (N_6161,N_5899,N_5878);
and U6162 (N_6162,N_5278,N_5363);
and U6163 (N_6163,N_5954,N_5604);
nor U6164 (N_6164,N_5579,N_5108);
xor U6165 (N_6165,N_5720,N_5375);
nand U6166 (N_6166,N_5914,N_5555);
nor U6167 (N_6167,N_5001,N_5673);
or U6168 (N_6168,N_5520,N_5163);
nand U6169 (N_6169,N_5279,N_5429);
nand U6170 (N_6170,N_5383,N_5662);
nand U6171 (N_6171,N_5281,N_5999);
and U6172 (N_6172,N_5484,N_5862);
xnor U6173 (N_6173,N_5358,N_5131);
xnor U6174 (N_6174,N_5490,N_5680);
and U6175 (N_6175,N_5494,N_5307);
or U6176 (N_6176,N_5802,N_5238);
nand U6177 (N_6177,N_5130,N_5941);
xor U6178 (N_6178,N_5497,N_5365);
xnor U6179 (N_6179,N_5524,N_5519);
nor U6180 (N_6180,N_5441,N_5477);
xor U6181 (N_6181,N_5452,N_5310);
or U6182 (N_6182,N_5979,N_5613);
and U6183 (N_6183,N_5731,N_5292);
nand U6184 (N_6184,N_5900,N_5033);
nand U6185 (N_6185,N_5528,N_5585);
and U6186 (N_6186,N_5823,N_5605);
xnor U6187 (N_6187,N_5237,N_5803);
xor U6188 (N_6188,N_5910,N_5706);
nor U6189 (N_6189,N_5866,N_5962);
nand U6190 (N_6190,N_5095,N_5134);
and U6191 (N_6191,N_5267,N_5026);
or U6192 (N_6192,N_5262,N_5392);
and U6193 (N_6193,N_5898,N_5474);
or U6194 (N_6194,N_5314,N_5158);
or U6195 (N_6195,N_5611,N_5717);
and U6196 (N_6196,N_5421,N_5196);
nor U6197 (N_6197,N_5155,N_5885);
or U6198 (N_6198,N_5114,N_5010);
and U6199 (N_6199,N_5695,N_5951);
xnor U6200 (N_6200,N_5981,N_5078);
or U6201 (N_6201,N_5070,N_5151);
nand U6202 (N_6202,N_5220,N_5185);
or U6203 (N_6203,N_5721,N_5475);
xor U6204 (N_6204,N_5997,N_5686);
nor U6205 (N_6205,N_5011,N_5176);
nor U6206 (N_6206,N_5887,N_5782);
nand U6207 (N_6207,N_5199,N_5172);
and U6208 (N_6208,N_5246,N_5970);
or U6209 (N_6209,N_5006,N_5681);
and U6210 (N_6210,N_5391,N_5117);
xor U6211 (N_6211,N_5495,N_5776);
or U6212 (N_6212,N_5127,N_5618);
xnor U6213 (N_6213,N_5850,N_5881);
or U6214 (N_6214,N_5911,N_5152);
or U6215 (N_6215,N_5040,N_5827);
xnor U6216 (N_6216,N_5178,N_5935);
and U6217 (N_6217,N_5670,N_5067);
and U6218 (N_6218,N_5081,N_5753);
nand U6219 (N_6219,N_5339,N_5165);
nor U6220 (N_6220,N_5049,N_5842);
nand U6221 (N_6221,N_5312,N_5136);
or U6222 (N_6222,N_5225,N_5943);
or U6223 (N_6223,N_5055,N_5294);
or U6224 (N_6224,N_5726,N_5056);
xnor U6225 (N_6225,N_5980,N_5598);
and U6226 (N_6226,N_5580,N_5459);
nand U6227 (N_6227,N_5523,N_5560);
nand U6228 (N_6228,N_5571,N_5256);
and U6229 (N_6229,N_5181,N_5816);
and U6230 (N_6230,N_5586,N_5603);
xor U6231 (N_6231,N_5813,N_5737);
or U6232 (N_6232,N_5115,N_5643);
or U6233 (N_6233,N_5214,N_5858);
or U6234 (N_6234,N_5138,N_5345);
nand U6235 (N_6235,N_5457,N_5259);
nand U6236 (N_6236,N_5424,N_5432);
nor U6237 (N_6237,N_5444,N_5886);
and U6238 (N_6238,N_5282,N_5260);
nor U6239 (N_6239,N_5311,N_5321);
and U6240 (N_6240,N_5562,N_5728);
xor U6241 (N_6241,N_5727,N_5465);
nor U6242 (N_6242,N_5814,N_5061);
and U6243 (N_6243,N_5875,N_5790);
nor U6244 (N_6244,N_5077,N_5566);
nor U6245 (N_6245,N_5897,N_5526);
nor U6246 (N_6246,N_5072,N_5837);
or U6247 (N_6247,N_5844,N_5500);
nand U6248 (N_6248,N_5442,N_5835);
xnor U6249 (N_6249,N_5976,N_5679);
nor U6250 (N_6250,N_5931,N_5404);
nand U6251 (N_6251,N_5573,N_5051);
nand U6252 (N_6252,N_5959,N_5757);
nor U6253 (N_6253,N_5360,N_5714);
and U6254 (N_6254,N_5787,N_5052);
or U6255 (N_6255,N_5109,N_5393);
xor U6256 (N_6256,N_5923,N_5433);
or U6257 (N_6257,N_5896,N_5137);
xnor U6258 (N_6258,N_5833,N_5796);
nand U6259 (N_6259,N_5638,N_5387);
and U6260 (N_6260,N_5852,N_5946);
xnor U6261 (N_6261,N_5810,N_5892);
xor U6262 (N_6262,N_5304,N_5169);
nor U6263 (N_6263,N_5569,N_5296);
nor U6264 (N_6264,N_5639,N_5637);
xnor U6265 (N_6265,N_5344,N_5945);
nor U6266 (N_6266,N_5537,N_5531);
or U6267 (N_6267,N_5476,N_5701);
nand U6268 (N_6268,N_5285,N_5030);
and U6269 (N_6269,N_5268,N_5654);
or U6270 (N_6270,N_5454,N_5594);
and U6271 (N_6271,N_5264,N_5386);
or U6272 (N_6272,N_5340,N_5758);
nor U6273 (N_6273,N_5581,N_5533);
and U6274 (N_6274,N_5492,N_5406);
or U6275 (N_6275,N_5378,N_5851);
nand U6276 (N_6276,N_5408,N_5901);
nor U6277 (N_6277,N_5162,N_5403);
or U6278 (N_6278,N_5799,N_5175);
and U6279 (N_6279,N_5554,N_5356);
xnor U6280 (N_6280,N_5846,N_5653);
xnor U6281 (N_6281,N_5174,N_5741);
xor U6282 (N_6282,N_5659,N_5071);
xor U6283 (N_6283,N_5349,N_5666);
xnor U6284 (N_6284,N_5120,N_5487);
nor U6285 (N_6285,N_5996,N_5161);
nor U6286 (N_6286,N_5749,N_5041);
nand U6287 (N_6287,N_5830,N_5564);
xnor U6288 (N_6288,N_5105,N_5685);
and U6289 (N_6289,N_5303,N_5422);
nand U6290 (N_6290,N_5317,N_5440);
nand U6291 (N_6291,N_5539,N_5658);
and U6292 (N_6292,N_5546,N_5780);
xnor U6293 (N_6293,N_5300,N_5648);
nor U6294 (N_6294,N_5811,N_5867);
nor U6295 (N_6295,N_5445,N_5649);
xnor U6296 (N_6296,N_5407,N_5189);
or U6297 (N_6297,N_5688,N_5545);
nand U6298 (N_6298,N_5733,N_5337);
xor U6299 (N_6299,N_5183,N_5308);
or U6300 (N_6300,N_5517,N_5641);
nor U6301 (N_6301,N_5118,N_5295);
nor U6302 (N_6302,N_5482,N_5628);
nor U6303 (N_6303,N_5855,N_5187);
nand U6304 (N_6304,N_5367,N_5065);
xnor U6305 (N_6305,N_5288,N_5091);
nand U6306 (N_6306,N_5883,N_5399);
xor U6307 (N_6307,N_5043,N_5993);
or U6308 (N_6308,N_5507,N_5008);
xnor U6309 (N_6309,N_5203,N_5032);
nand U6310 (N_6310,N_5505,N_5874);
and U6311 (N_6311,N_5289,N_5007);
nor U6312 (N_6312,N_5098,N_5234);
nand U6313 (N_6313,N_5574,N_5977);
and U6314 (N_6314,N_5958,N_5222);
xnor U6315 (N_6315,N_5111,N_5978);
and U6316 (N_6316,N_5696,N_5116);
nor U6317 (N_6317,N_5804,N_5479);
nor U6318 (N_6318,N_5514,N_5319);
and U6319 (N_6319,N_5128,N_5207);
and U6320 (N_6320,N_5869,N_5647);
nand U6321 (N_6321,N_5828,N_5059);
nor U6322 (N_6322,N_5501,N_5625);
and U6323 (N_6323,N_5503,N_5671);
nand U6324 (N_6324,N_5998,N_5948);
or U6325 (N_6325,N_5509,N_5567);
nand U6326 (N_6326,N_5194,N_5944);
and U6327 (N_6327,N_5917,N_5293);
nand U6328 (N_6328,N_5548,N_5736);
and U6329 (N_6329,N_5801,N_5315);
and U6330 (N_6330,N_5884,N_5502);
nor U6331 (N_6331,N_5266,N_5435);
and U6332 (N_6332,N_5608,N_5496);
nand U6333 (N_6333,N_5362,N_5229);
nor U6334 (N_6334,N_5082,N_5856);
or U6335 (N_6335,N_5722,N_5499);
nor U6336 (N_6336,N_5506,N_5877);
nor U6337 (N_6337,N_5913,N_5766);
or U6338 (N_6338,N_5275,N_5346);
or U6339 (N_6339,N_5254,N_5645);
or U6340 (N_6340,N_5037,N_5226);
xor U6341 (N_6341,N_5283,N_5995);
nand U6342 (N_6342,N_5739,N_5880);
and U6343 (N_6343,N_5644,N_5969);
or U6344 (N_6344,N_5634,N_5663);
nor U6345 (N_6345,N_5987,N_5334);
and U6346 (N_6346,N_5064,N_5048);
xnor U6347 (N_6347,N_5046,N_5153);
xnor U6348 (N_6348,N_5620,N_5916);
and U6349 (N_6349,N_5947,N_5359);
nand U6350 (N_6350,N_5961,N_5952);
and U6351 (N_6351,N_5166,N_5990);
or U6352 (N_6352,N_5054,N_5102);
and U6353 (N_6353,N_5436,N_5023);
or U6354 (N_6354,N_5413,N_5058);
xor U6355 (N_6355,N_5074,N_5291);
or U6356 (N_6356,N_5170,N_5385);
nand U6357 (N_6357,N_5232,N_5538);
or U6358 (N_6358,N_5418,N_5786);
nand U6359 (N_6359,N_5584,N_5577);
or U6360 (N_6360,N_5027,N_5542);
nand U6361 (N_6361,N_5168,N_5876);
and U6362 (N_6362,N_5919,N_5838);
or U6363 (N_6363,N_5553,N_5768);
nand U6364 (N_6364,N_5773,N_5778);
nor U6365 (N_6365,N_5455,N_5097);
nor U6366 (N_6366,N_5411,N_5909);
or U6367 (N_6367,N_5142,N_5597);
nand U6368 (N_6368,N_5521,N_5323);
nor U6369 (N_6369,N_5836,N_5427);
and U6370 (N_6370,N_5568,N_5902);
or U6371 (N_6371,N_5141,N_5784);
and U6372 (N_6372,N_5491,N_5789);
nand U6373 (N_6373,N_5198,N_5824);
and U6374 (N_6374,N_5689,N_5350);
nand U6375 (N_6375,N_5019,N_5100);
xor U6376 (N_6376,N_5160,N_5154);
nor U6377 (N_6377,N_5583,N_5966);
and U6378 (N_6378,N_5253,N_5087);
nor U6379 (N_6379,N_5298,N_5665);
nor U6380 (N_6380,N_5702,N_5767);
and U6381 (N_6381,N_5084,N_5228);
xnor U6382 (N_6382,N_5729,N_5691);
nand U6383 (N_6383,N_5269,N_5188);
nor U6384 (N_6384,N_5854,N_5932);
and U6385 (N_6385,N_5600,N_5029);
nor U6386 (N_6386,N_5079,N_5423);
or U6387 (N_6387,N_5347,N_5124);
and U6388 (N_6388,N_5607,N_5905);
or U6389 (N_6389,N_5066,N_5277);
or U6390 (N_6390,N_5144,N_5103);
and U6391 (N_6391,N_5236,N_5716);
nand U6392 (N_6392,N_5191,N_5249);
nor U6393 (N_6393,N_5348,N_5416);
and U6394 (N_6394,N_5710,N_5443);
xnor U6395 (N_6395,N_5825,N_5333);
or U6396 (N_6396,N_5469,N_5425);
nand U6397 (N_6397,N_5870,N_5640);
xnor U6398 (N_6398,N_5488,N_5552);
xor U6399 (N_6399,N_5817,N_5092);
or U6400 (N_6400,N_5621,N_5551);
xor U6401 (N_6401,N_5149,N_5794);
xnor U6402 (N_6402,N_5839,N_5879);
xnor U6403 (N_6403,N_5532,N_5400);
nor U6404 (N_6404,N_5508,N_5210);
or U6405 (N_6405,N_5614,N_5002);
xnor U6406 (N_6406,N_5903,N_5912);
xnor U6407 (N_6407,N_5927,N_5219);
or U6408 (N_6408,N_5861,N_5486);
nor U6409 (N_6409,N_5669,N_5536);
nand U6410 (N_6410,N_5402,N_5209);
and U6411 (N_6411,N_5366,N_5715);
and U6412 (N_6412,N_5493,N_5156);
or U6413 (N_6413,N_5698,N_5456);
or U6414 (N_6414,N_5719,N_5707);
or U6415 (N_6415,N_5250,N_5629);
xnor U6416 (N_6416,N_5703,N_5667);
or U6417 (N_6417,N_5322,N_5775);
and U6418 (N_6418,N_5769,N_5576);
nor U6419 (N_6419,N_5764,N_5212);
nor U6420 (N_6420,N_5357,N_5745);
and U6421 (N_6421,N_5559,N_5557);
xor U6422 (N_6422,N_5675,N_5272);
or U6423 (N_6423,N_5353,N_5419);
or U6424 (N_6424,N_5069,N_5713);
nor U6425 (N_6425,N_5394,N_5157);
and U6426 (N_6426,N_5857,N_5949);
nand U6427 (N_6427,N_5370,N_5206);
xnor U6428 (N_6428,N_5788,N_5245);
nor U6429 (N_6429,N_5326,N_5907);
and U6430 (N_6430,N_5967,N_5971);
nor U6431 (N_6431,N_5233,N_5218);
xnor U6432 (N_6432,N_5129,N_5227);
nor U6433 (N_6433,N_5409,N_5871);
nor U6434 (N_6434,N_5655,N_5261);
and U6435 (N_6435,N_5690,N_5845);
and U6436 (N_6436,N_5343,N_5774);
nor U6437 (N_6437,N_5410,N_5765);
or U6438 (N_6438,N_5623,N_5747);
and U6439 (N_6439,N_5504,N_5389);
xnor U6440 (N_6440,N_5113,N_5697);
or U6441 (N_6441,N_5035,N_5989);
nor U6442 (N_6442,N_5057,N_5556);
xor U6443 (N_6443,N_5606,N_5740);
xor U6444 (N_6444,N_5610,N_5806);
nand U6445 (N_6445,N_5661,N_5709);
and U6446 (N_6446,N_5812,N_5381);
nor U6447 (N_6447,N_5104,N_5734);
xnor U6448 (N_6448,N_5184,N_5832);
nor U6449 (N_6449,N_5630,N_5430);
and U6450 (N_6450,N_5276,N_5186);
nor U6451 (N_6451,N_5083,N_5135);
nand U6452 (N_6452,N_5793,N_5712);
or U6453 (N_6453,N_5258,N_5754);
or U6454 (N_6454,N_5601,N_5462);
xnor U6455 (N_6455,N_5906,N_5265);
xnor U6456 (N_6456,N_5309,N_5920);
xnor U6457 (N_6457,N_5485,N_5889);
nand U6458 (N_6458,N_5821,N_5937);
and U6459 (N_6459,N_5244,N_5190);
nand U6460 (N_6460,N_5815,N_5164);
xnor U6461 (N_6461,N_5122,N_5752);
xnor U6462 (N_6462,N_5042,N_5284);
and U6463 (N_6463,N_5942,N_5299);
nand U6464 (N_6464,N_5684,N_5022);
xor U6465 (N_6465,N_5145,N_5940);
and U6466 (N_6466,N_5020,N_5809);
nand U6467 (N_6467,N_5956,N_5891);
or U6468 (N_6468,N_5371,N_5925);
xor U6469 (N_6469,N_5953,N_5904);
and U6470 (N_6470,N_5012,N_5535);
nand U6471 (N_6471,N_5121,N_5018);
and U6472 (N_6472,N_5243,N_5096);
nor U6473 (N_6473,N_5053,N_5316);
nand U6474 (N_6474,N_5540,N_5819);
xnor U6475 (N_6475,N_5195,N_5044);
nand U6476 (N_6476,N_5732,N_5549);
and U6477 (N_6477,N_5464,N_5591);
and U6478 (N_6478,N_5379,N_5960);
xnor U6479 (N_6479,N_5143,N_5062);
or U6480 (N_6480,N_5863,N_5770);
and U6481 (N_6481,N_5805,N_5843);
nor U6482 (N_6482,N_5771,N_5582);
xnor U6483 (N_6483,N_5974,N_5063);
and U6484 (N_6484,N_5895,N_5522);
and U6485 (N_6485,N_5201,N_5376);
nor U6486 (N_6486,N_5795,N_5377);
nor U6487 (N_6487,N_5544,N_5759);
and U6488 (N_6488,N_5221,N_5205);
nand U6489 (N_6489,N_5592,N_5651);
or U6490 (N_6490,N_5938,N_5818);
nor U6491 (N_6491,N_5005,N_5306);
nand U6492 (N_6492,N_5615,N_5182);
xnor U6493 (N_6493,N_5984,N_5975);
and U6494 (N_6494,N_5915,N_5478);
nand U6495 (N_6495,N_5273,N_5963);
nor U6496 (N_6496,N_5021,N_5512);
or U6497 (N_6497,N_5252,N_5123);
nor U6498 (N_6498,N_5988,N_5003);
xor U6499 (N_6499,N_5380,N_5146);
and U6500 (N_6500,N_5679,N_5489);
or U6501 (N_6501,N_5944,N_5026);
and U6502 (N_6502,N_5333,N_5676);
or U6503 (N_6503,N_5655,N_5220);
xnor U6504 (N_6504,N_5709,N_5849);
xnor U6505 (N_6505,N_5560,N_5561);
xor U6506 (N_6506,N_5944,N_5640);
xor U6507 (N_6507,N_5984,N_5400);
and U6508 (N_6508,N_5630,N_5004);
and U6509 (N_6509,N_5269,N_5182);
and U6510 (N_6510,N_5741,N_5971);
nand U6511 (N_6511,N_5335,N_5891);
nor U6512 (N_6512,N_5108,N_5888);
xor U6513 (N_6513,N_5290,N_5511);
xor U6514 (N_6514,N_5482,N_5805);
nand U6515 (N_6515,N_5278,N_5773);
and U6516 (N_6516,N_5580,N_5180);
or U6517 (N_6517,N_5573,N_5270);
nor U6518 (N_6518,N_5016,N_5619);
nand U6519 (N_6519,N_5837,N_5719);
nand U6520 (N_6520,N_5782,N_5362);
or U6521 (N_6521,N_5157,N_5061);
xnor U6522 (N_6522,N_5575,N_5609);
xor U6523 (N_6523,N_5985,N_5595);
nand U6524 (N_6524,N_5912,N_5109);
xor U6525 (N_6525,N_5423,N_5189);
and U6526 (N_6526,N_5141,N_5967);
and U6527 (N_6527,N_5055,N_5339);
nor U6528 (N_6528,N_5741,N_5464);
or U6529 (N_6529,N_5000,N_5416);
or U6530 (N_6530,N_5221,N_5641);
nor U6531 (N_6531,N_5479,N_5372);
nand U6532 (N_6532,N_5049,N_5545);
and U6533 (N_6533,N_5043,N_5635);
nor U6534 (N_6534,N_5650,N_5857);
xnor U6535 (N_6535,N_5825,N_5986);
and U6536 (N_6536,N_5702,N_5273);
xnor U6537 (N_6537,N_5652,N_5746);
and U6538 (N_6538,N_5824,N_5240);
or U6539 (N_6539,N_5533,N_5613);
and U6540 (N_6540,N_5202,N_5275);
xor U6541 (N_6541,N_5378,N_5086);
nor U6542 (N_6542,N_5697,N_5002);
nand U6543 (N_6543,N_5069,N_5589);
and U6544 (N_6544,N_5131,N_5572);
xnor U6545 (N_6545,N_5194,N_5523);
nand U6546 (N_6546,N_5544,N_5007);
and U6547 (N_6547,N_5328,N_5616);
nor U6548 (N_6548,N_5246,N_5854);
or U6549 (N_6549,N_5562,N_5559);
or U6550 (N_6550,N_5405,N_5881);
xor U6551 (N_6551,N_5931,N_5294);
and U6552 (N_6552,N_5044,N_5293);
nor U6553 (N_6553,N_5557,N_5265);
nor U6554 (N_6554,N_5139,N_5391);
xor U6555 (N_6555,N_5528,N_5282);
nand U6556 (N_6556,N_5215,N_5911);
or U6557 (N_6557,N_5295,N_5663);
and U6558 (N_6558,N_5750,N_5118);
nor U6559 (N_6559,N_5699,N_5560);
nand U6560 (N_6560,N_5070,N_5342);
or U6561 (N_6561,N_5146,N_5110);
and U6562 (N_6562,N_5583,N_5838);
or U6563 (N_6563,N_5047,N_5198);
or U6564 (N_6564,N_5669,N_5924);
xor U6565 (N_6565,N_5854,N_5137);
nand U6566 (N_6566,N_5021,N_5464);
or U6567 (N_6567,N_5372,N_5189);
nand U6568 (N_6568,N_5566,N_5375);
nor U6569 (N_6569,N_5488,N_5195);
and U6570 (N_6570,N_5631,N_5338);
xor U6571 (N_6571,N_5846,N_5389);
xnor U6572 (N_6572,N_5506,N_5160);
and U6573 (N_6573,N_5471,N_5583);
xor U6574 (N_6574,N_5956,N_5904);
nor U6575 (N_6575,N_5278,N_5090);
nand U6576 (N_6576,N_5070,N_5424);
nand U6577 (N_6577,N_5015,N_5458);
nand U6578 (N_6578,N_5850,N_5606);
or U6579 (N_6579,N_5209,N_5816);
and U6580 (N_6580,N_5724,N_5095);
or U6581 (N_6581,N_5023,N_5116);
nand U6582 (N_6582,N_5559,N_5136);
or U6583 (N_6583,N_5063,N_5607);
and U6584 (N_6584,N_5047,N_5033);
xnor U6585 (N_6585,N_5558,N_5902);
nor U6586 (N_6586,N_5809,N_5863);
xor U6587 (N_6587,N_5876,N_5860);
nand U6588 (N_6588,N_5133,N_5462);
and U6589 (N_6589,N_5464,N_5756);
nand U6590 (N_6590,N_5182,N_5222);
nor U6591 (N_6591,N_5370,N_5486);
xnor U6592 (N_6592,N_5282,N_5790);
or U6593 (N_6593,N_5649,N_5339);
or U6594 (N_6594,N_5465,N_5363);
nand U6595 (N_6595,N_5388,N_5948);
xnor U6596 (N_6596,N_5462,N_5557);
nor U6597 (N_6597,N_5607,N_5526);
or U6598 (N_6598,N_5912,N_5077);
xnor U6599 (N_6599,N_5420,N_5593);
and U6600 (N_6600,N_5941,N_5266);
and U6601 (N_6601,N_5159,N_5239);
nor U6602 (N_6602,N_5046,N_5656);
xor U6603 (N_6603,N_5799,N_5612);
and U6604 (N_6604,N_5024,N_5478);
or U6605 (N_6605,N_5754,N_5467);
nor U6606 (N_6606,N_5055,N_5983);
nand U6607 (N_6607,N_5851,N_5494);
xor U6608 (N_6608,N_5896,N_5971);
and U6609 (N_6609,N_5060,N_5308);
xnor U6610 (N_6610,N_5351,N_5584);
and U6611 (N_6611,N_5624,N_5685);
nand U6612 (N_6612,N_5696,N_5816);
and U6613 (N_6613,N_5971,N_5464);
xnor U6614 (N_6614,N_5523,N_5287);
or U6615 (N_6615,N_5494,N_5083);
and U6616 (N_6616,N_5819,N_5309);
and U6617 (N_6617,N_5506,N_5282);
or U6618 (N_6618,N_5652,N_5881);
xnor U6619 (N_6619,N_5048,N_5472);
nand U6620 (N_6620,N_5510,N_5533);
nor U6621 (N_6621,N_5976,N_5530);
nand U6622 (N_6622,N_5177,N_5529);
xnor U6623 (N_6623,N_5847,N_5881);
nand U6624 (N_6624,N_5910,N_5632);
or U6625 (N_6625,N_5910,N_5626);
xor U6626 (N_6626,N_5464,N_5721);
and U6627 (N_6627,N_5925,N_5289);
xnor U6628 (N_6628,N_5203,N_5293);
xnor U6629 (N_6629,N_5538,N_5898);
nand U6630 (N_6630,N_5396,N_5898);
or U6631 (N_6631,N_5681,N_5038);
nand U6632 (N_6632,N_5477,N_5136);
nand U6633 (N_6633,N_5886,N_5283);
nand U6634 (N_6634,N_5351,N_5626);
xnor U6635 (N_6635,N_5807,N_5790);
xnor U6636 (N_6636,N_5947,N_5869);
and U6637 (N_6637,N_5329,N_5693);
nand U6638 (N_6638,N_5161,N_5341);
and U6639 (N_6639,N_5460,N_5334);
and U6640 (N_6640,N_5071,N_5197);
or U6641 (N_6641,N_5616,N_5087);
nand U6642 (N_6642,N_5968,N_5287);
and U6643 (N_6643,N_5201,N_5609);
nand U6644 (N_6644,N_5082,N_5268);
xnor U6645 (N_6645,N_5048,N_5324);
nand U6646 (N_6646,N_5309,N_5618);
and U6647 (N_6647,N_5359,N_5461);
nor U6648 (N_6648,N_5755,N_5252);
or U6649 (N_6649,N_5073,N_5144);
nor U6650 (N_6650,N_5302,N_5409);
xnor U6651 (N_6651,N_5913,N_5498);
nand U6652 (N_6652,N_5465,N_5623);
nand U6653 (N_6653,N_5145,N_5049);
xnor U6654 (N_6654,N_5763,N_5686);
xor U6655 (N_6655,N_5513,N_5703);
xnor U6656 (N_6656,N_5067,N_5577);
nor U6657 (N_6657,N_5646,N_5533);
xor U6658 (N_6658,N_5774,N_5064);
nand U6659 (N_6659,N_5834,N_5089);
or U6660 (N_6660,N_5091,N_5373);
nand U6661 (N_6661,N_5835,N_5670);
nor U6662 (N_6662,N_5047,N_5042);
nor U6663 (N_6663,N_5926,N_5477);
or U6664 (N_6664,N_5690,N_5008);
or U6665 (N_6665,N_5414,N_5425);
nand U6666 (N_6666,N_5511,N_5520);
or U6667 (N_6667,N_5481,N_5362);
nor U6668 (N_6668,N_5436,N_5320);
nor U6669 (N_6669,N_5895,N_5904);
xnor U6670 (N_6670,N_5138,N_5125);
nand U6671 (N_6671,N_5984,N_5338);
xnor U6672 (N_6672,N_5666,N_5406);
nand U6673 (N_6673,N_5486,N_5992);
or U6674 (N_6674,N_5933,N_5911);
xor U6675 (N_6675,N_5367,N_5232);
nor U6676 (N_6676,N_5767,N_5750);
or U6677 (N_6677,N_5163,N_5877);
and U6678 (N_6678,N_5056,N_5094);
xnor U6679 (N_6679,N_5432,N_5546);
nor U6680 (N_6680,N_5879,N_5299);
and U6681 (N_6681,N_5847,N_5146);
or U6682 (N_6682,N_5293,N_5972);
or U6683 (N_6683,N_5438,N_5967);
nand U6684 (N_6684,N_5399,N_5908);
xor U6685 (N_6685,N_5126,N_5352);
and U6686 (N_6686,N_5493,N_5593);
or U6687 (N_6687,N_5035,N_5319);
nand U6688 (N_6688,N_5357,N_5670);
nand U6689 (N_6689,N_5349,N_5606);
nor U6690 (N_6690,N_5847,N_5950);
xnor U6691 (N_6691,N_5804,N_5688);
nand U6692 (N_6692,N_5959,N_5909);
nand U6693 (N_6693,N_5317,N_5254);
and U6694 (N_6694,N_5212,N_5544);
nand U6695 (N_6695,N_5089,N_5191);
and U6696 (N_6696,N_5846,N_5692);
nand U6697 (N_6697,N_5254,N_5084);
nand U6698 (N_6698,N_5731,N_5063);
nor U6699 (N_6699,N_5622,N_5742);
nor U6700 (N_6700,N_5264,N_5227);
and U6701 (N_6701,N_5977,N_5202);
and U6702 (N_6702,N_5423,N_5350);
xor U6703 (N_6703,N_5116,N_5444);
nand U6704 (N_6704,N_5541,N_5053);
or U6705 (N_6705,N_5686,N_5679);
xor U6706 (N_6706,N_5682,N_5244);
nand U6707 (N_6707,N_5508,N_5673);
nor U6708 (N_6708,N_5592,N_5225);
and U6709 (N_6709,N_5907,N_5993);
or U6710 (N_6710,N_5973,N_5974);
nor U6711 (N_6711,N_5611,N_5762);
and U6712 (N_6712,N_5544,N_5095);
nor U6713 (N_6713,N_5757,N_5539);
or U6714 (N_6714,N_5280,N_5566);
nand U6715 (N_6715,N_5019,N_5081);
nand U6716 (N_6716,N_5038,N_5645);
and U6717 (N_6717,N_5194,N_5961);
and U6718 (N_6718,N_5620,N_5501);
nor U6719 (N_6719,N_5237,N_5996);
xor U6720 (N_6720,N_5547,N_5111);
and U6721 (N_6721,N_5628,N_5821);
and U6722 (N_6722,N_5015,N_5847);
xor U6723 (N_6723,N_5116,N_5375);
xnor U6724 (N_6724,N_5357,N_5454);
and U6725 (N_6725,N_5718,N_5573);
nor U6726 (N_6726,N_5992,N_5304);
and U6727 (N_6727,N_5238,N_5851);
or U6728 (N_6728,N_5431,N_5838);
or U6729 (N_6729,N_5505,N_5171);
xor U6730 (N_6730,N_5611,N_5089);
xnor U6731 (N_6731,N_5409,N_5272);
and U6732 (N_6732,N_5639,N_5624);
xnor U6733 (N_6733,N_5074,N_5808);
or U6734 (N_6734,N_5522,N_5705);
and U6735 (N_6735,N_5728,N_5068);
nor U6736 (N_6736,N_5243,N_5539);
nand U6737 (N_6737,N_5552,N_5041);
and U6738 (N_6738,N_5564,N_5425);
or U6739 (N_6739,N_5078,N_5976);
nand U6740 (N_6740,N_5073,N_5993);
nor U6741 (N_6741,N_5557,N_5838);
nand U6742 (N_6742,N_5271,N_5835);
or U6743 (N_6743,N_5234,N_5691);
nor U6744 (N_6744,N_5028,N_5462);
nand U6745 (N_6745,N_5162,N_5948);
or U6746 (N_6746,N_5451,N_5857);
xnor U6747 (N_6747,N_5725,N_5655);
nand U6748 (N_6748,N_5593,N_5132);
and U6749 (N_6749,N_5948,N_5190);
and U6750 (N_6750,N_5123,N_5239);
xnor U6751 (N_6751,N_5839,N_5837);
and U6752 (N_6752,N_5375,N_5775);
nor U6753 (N_6753,N_5419,N_5373);
nand U6754 (N_6754,N_5870,N_5258);
or U6755 (N_6755,N_5236,N_5784);
xnor U6756 (N_6756,N_5923,N_5910);
nand U6757 (N_6757,N_5795,N_5037);
xor U6758 (N_6758,N_5977,N_5296);
xor U6759 (N_6759,N_5826,N_5127);
xnor U6760 (N_6760,N_5507,N_5393);
or U6761 (N_6761,N_5279,N_5350);
or U6762 (N_6762,N_5865,N_5909);
or U6763 (N_6763,N_5201,N_5318);
nand U6764 (N_6764,N_5978,N_5347);
or U6765 (N_6765,N_5752,N_5599);
and U6766 (N_6766,N_5062,N_5848);
and U6767 (N_6767,N_5449,N_5387);
nand U6768 (N_6768,N_5530,N_5296);
or U6769 (N_6769,N_5694,N_5742);
nor U6770 (N_6770,N_5166,N_5794);
or U6771 (N_6771,N_5833,N_5217);
nor U6772 (N_6772,N_5031,N_5493);
or U6773 (N_6773,N_5853,N_5884);
or U6774 (N_6774,N_5832,N_5308);
or U6775 (N_6775,N_5293,N_5241);
nor U6776 (N_6776,N_5660,N_5442);
nand U6777 (N_6777,N_5236,N_5922);
xor U6778 (N_6778,N_5434,N_5425);
and U6779 (N_6779,N_5838,N_5558);
nand U6780 (N_6780,N_5951,N_5937);
nand U6781 (N_6781,N_5480,N_5392);
or U6782 (N_6782,N_5472,N_5817);
xnor U6783 (N_6783,N_5894,N_5853);
nor U6784 (N_6784,N_5709,N_5482);
and U6785 (N_6785,N_5762,N_5293);
or U6786 (N_6786,N_5024,N_5152);
xnor U6787 (N_6787,N_5609,N_5271);
and U6788 (N_6788,N_5008,N_5622);
or U6789 (N_6789,N_5712,N_5331);
nand U6790 (N_6790,N_5829,N_5259);
and U6791 (N_6791,N_5901,N_5093);
or U6792 (N_6792,N_5318,N_5889);
nand U6793 (N_6793,N_5563,N_5408);
xnor U6794 (N_6794,N_5380,N_5366);
or U6795 (N_6795,N_5915,N_5552);
nand U6796 (N_6796,N_5751,N_5643);
xnor U6797 (N_6797,N_5357,N_5198);
nor U6798 (N_6798,N_5360,N_5373);
nor U6799 (N_6799,N_5344,N_5659);
xnor U6800 (N_6800,N_5302,N_5741);
or U6801 (N_6801,N_5181,N_5090);
nand U6802 (N_6802,N_5032,N_5956);
or U6803 (N_6803,N_5643,N_5282);
nand U6804 (N_6804,N_5897,N_5394);
xor U6805 (N_6805,N_5440,N_5924);
and U6806 (N_6806,N_5853,N_5350);
nor U6807 (N_6807,N_5230,N_5235);
nand U6808 (N_6808,N_5309,N_5541);
or U6809 (N_6809,N_5014,N_5027);
xor U6810 (N_6810,N_5735,N_5021);
nand U6811 (N_6811,N_5634,N_5380);
nand U6812 (N_6812,N_5368,N_5245);
or U6813 (N_6813,N_5232,N_5427);
nand U6814 (N_6814,N_5046,N_5511);
and U6815 (N_6815,N_5582,N_5860);
nand U6816 (N_6816,N_5492,N_5872);
xnor U6817 (N_6817,N_5712,N_5386);
xor U6818 (N_6818,N_5039,N_5916);
or U6819 (N_6819,N_5365,N_5121);
or U6820 (N_6820,N_5275,N_5425);
and U6821 (N_6821,N_5291,N_5749);
xnor U6822 (N_6822,N_5935,N_5680);
and U6823 (N_6823,N_5119,N_5916);
or U6824 (N_6824,N_5056,N_5602);
nand U6825 (N_6825,N_5344,N_5119);
nor U6826 (N_6826,N_5076,N_5834);
or U6827 (N_6827,N_5171,N_5348);
nor U6828 (N_6828,N_5585,N_5736);
xor U6829 (N_6829,N_5264,N_5763);
or U6830 (N_6830,N_5563,N_5887);
nor U6831 (N_6831,N_5489,N_5894);
or U6832 (N_6832,N_5485,N_5223);
nor U6833 (N_6833,N_5948,N_5332);
nand U6834 (N_6834,N_5102,N_5623);
and U6835 (N_6835,N_5361,N_5038);
nor U6836 (N_6836,N_5441,N_5381);
or U6837 (N_6837,N_5793,N_5208);
nand U6838 (N_6838,N_5334,N_5757);
and U6839 (N_6839,N_5489,N_5603);
nor U6840 (N_6840,N_5129,N_5390);
or U6841 (N_6841,N_5582,N_5124);
nand U6842 (N_6842,N_5814,N_5995);
xnor U6843 (N_6843,N_5343,N_5075);
xnor U6844 (N_6844,N_5463,N_5339);
xnor U6845 (N_6845,N_5064,N_5220);
nor U6846 (N_6846,N_5825,N_5490);
nor U6847 (N_6847,N_5246,N_5756);
xor U6848 (N_6848,N_5107,N_5841);
nor U6849 (N_6849,N_5807,N_5502);
or U6850 (N_6850,N_5029,N_5082);
nand U6851 (N_6851,N_5421,N_5815);
nor U6852 (N_6852,N_5219,N_5231);
nand U6853 (N_6853,N_5000,N_5631);
nand U6854 (N_6854,N_5071,N_5600);
nand U6855 (N_6855,N_5506,N_5642);
or U6856 (N_6856,N_5206,N_5484);
or U6857 (N_6857,N_5664,N_5510);
and U6858 (N_6858,N_5415,N_5839);
nand U6859 (N_6859,N_5066,N_5061);
xnor U6860 (N_6860,N_5329,N_5820);
nand U6861 (N_6861,N_5231,N_5923);
and U6862 (N_6862,N_5928,N_5502);
nand U6863 (N_6863,N_5686,N_5943);
or U6864 (N_6864,N_5813,N_5740);
nand U6865 (N_6865,N_5905,N_5086);
nor U6866 (N_6866,N_5028,N_5553);
xnor U6867 (N_6867,N_5375,N_5527);
and U6868 (N_6868,N_5792,N_5544);
nand U6869 (N_6869,N_5636,N_5529);
nor U6870 (N_6870,N_5849,N_5313);
or U6871 (N_6871,N_5367,N_5134);
or U6872 (N_6872,N_5616,N_5646);
or U6873 (N_6873,N_5902,N_5021);
xnor U6874 (N_6874,N_5258,N_5782);
nor U6875 (N_6875,N_5988,N_5622);
or U6876 (N_6876,N_5726,N_5475);
nor U6877 (N_6877,N_5040,N_5912);
or U6878 (N_6878,N_5182,N_5930);
xnor U6879 (N_6879,N_5572,N_5251);
or U6880 (N_6880,N_5505,N_5772);
nor U6881 (N_6881,N_5611,N_5330);
and U6882 (N_6882,N_5053,N_5187);
and U6883 (N_6883,N_5351,N_5156);
xnor U6884 (N_6884,N_5349,N_5858);
xor U6885 (N_6885,N_5737,N_5316);
or U6886 (N_6886,N_5958,N_5678);
xnor U6887 (N_6887,N_5347,N_5193);
or U6888 (N_6888,N_5346,N_5170);
nor U6889 (N_6889,N_5942,N_5880);
or U6890 (N_6890,N_5178,N_5776);
or U6891 (N_6891,N_5254,N_5607);
nand U6892 (N_6892,N_5399,N_5084);
and U6893 (N_6893,N_5744,N_5912);
or U6894 (N_6894,N_5568,N_5291);
nor U6895 (N_6895,N_5754,N_5844);
nor U6896 (N_6896,N_5700,N_5242);
nor U6897 (N_6897,N_5840,N_5845);
xor U6898 (N_6898,N_5429,N_5050);
or U6899 (N_6899,N_5416,N_5849);
nand U6900 (N_6900,N_5063,N_5054);
nor U6901 (N_6901,N_5385,N_5396);
and U6902 (N_6902,N_5243,N_5420);
xor U6903 (N_6903,N_5194,N_5035);
or U6904 (N_6904,N_5884,N_5480);
and U6905 (N_6905,N_5662,N_5095);
nand U6906 (N_6906,N_5035,N_5328);
xnor U6907 (N_6907,N_5467,N_5856);
nand U6908 (N_6908,N_5613,N_5765);
and U6909 (N_6909,N_5167,N_5623);
xnor U6910 (N_6910,N_5806,N_5995);
or U6911 (N_6911,N_5365,N_5065);
or U6912 (N_6912,N_5758,N_5058);
and U6913 (N_6913,N_5828,N_5892);
nand U6914 (N_6914,N_5760,N_5095);
or U6915 (N_6915,N_5099,N_5923);
or U6916 (N_6916,N_5107,N_5691);
or U6917 (N_6917,N_5085,N_5575);
nand U6918 (N_6918,N_5847,N_5218);
xnor U6919 (N_6919,N_5560,N_5106);
or U6920 (N_6920,N_5053,N_5551);
or U6921 (N_6921,N_5477,N_5832);
nor U6922 (N_6922,N_5387,N_5771);
nor U6923 (N_6923,N_5500,N_5445);
and U6924 (N_6924,N_5878,N_5426);
nor U6925 (N_6925,N_5386,N_5754);
and U6926 (N_6926,N_5255,N_5832);
nand U6927 (N_6927,N_5591,N_5011);
and U6928 (N_6928,N_5707,N_5774);
and U6929 (N_6929,N_5101,N_5955);
or U6930 (N_6930,N_5413,N_5241);
or U6931 (N_6931,N_5490,N_5085);
nand U6932 (N_6932,N_5697,N_5008);
or U6933 (N_6933,N_5584,N_5413);
or U6934 (N_6934,N_5167,N_5621);
or U6935 (N_6935,N_5268,N_5350);
or U6936 (N_6936,N_5748,N_5879);
xnor U6937 (N_6937,N_5428,N_5527);
nand U6938 (N_6938,N_5021,N_5254);
nand U6939 (N_6939,N_5530,N_5046);
and U6940 (N_6940,N_5156,N_5918);
nor U6941 (N_6941,N_5444,N_5681);
nor U6942 (N_6942,N_5850,N_5864);
nor U6943 (N_6943,N_5684,N_5337);
nor U6944 (N_6944,N_5750,N_5395);
and U6945 (N_6945,N_5277,N_5439);
nor U6946 (N_6946,N_5829,N_5406);
and U6947 (N_6947,N_5736,N_5927);
xnor U6948 (N_6948,N_5926,N_5590);
xnor U6949 (N_6949,N_5452,N_5071);
nor U6950 (N_6950,N_5065,N_5784);
nand U6951 (N_6951,N_5357,N_5354);
nand U6952 (N_6952,N_5687,N_5782);
nor U6953 (N_6953,N_5475,N_5261);
and U6954 (N_6954,N_5054,N_5214);
and U6955 (N_6955,N_5478,N_5179);
nand U6956 (N_6956,N_5070,N_5134);
xor U6957 (N_6957,N_5473,N_5739);
or U6958 (N_6958,N_5841,N_5353);
nor U6959 (N_6959,N_5036,N_5456);
xor U6960 (N_6960,N_5500,N_5436);
and U6961 (N_6961,N_5287,N_5678);
nor U6962 (N_6962,N_5741,N_5934);
nor U6963 (N_6963,N_5238,N_5643);
xnor U6964 (N_6964,N_5605,N_5619);
xor U6965 (N_6965,N_5662,N_5807);
or U6966 (N_6966,N_5729,N_5223);
or U6967 (N_6967,N_5233,N_5258);
nor U6968 (N_6968,N_5101,N_5944);
xor U6969 (N_6969,N_5608,N_5977);
nand U6970 (N_6970,N_5654,N_5496);
nand U6971 (N_6971,N_5812,N_5579);
nand U6972 (N_6972,N_5753,N_5219);
nor U6973 (N_6973,N_5535,N_5275);
or U6974 (N_6974,N_5131,N_5781);
or U6975 (N_6975,N_5970,N_5408);
nand U6976 (N_6976,N_5096,N_5203);
xor U6977 (N_6977,N_5346,N_5343);
xnor U6978 (N_6978,N_5305,N_5332);
nor U6979 (N_6979,N_5225,N_5461);
xnor U6980 (N_6980,N_5698,N_5230);
xor U6981 (N_6981,N_5118,N_5663);
xor U6982 (N_6982,N_5743,N_5041);
nor U6983 (N_6983,N_5090,N_5021);
nand U6984 (N_6984,N_5533,N_5366);
xor U6985 (N_6985,N_5330,N_5249);
and U6986 (N_6986,N_5515,N_5789);
xnor U6987 (N_6987,N_5746,N_5300);
nor U6988 (N_6988,N_5510,N_5508);
nor U6989 (N_6989,N_5694,N_5285);
xor U6990 (N_6990,N_5577,N_5236);
nand U6991 (N_6991,N_5140,N_5689);
xnor U6992 (N_6992,N_5304,N_5584);
and U6993 (N_6993,N_5512,N_5385);
and U6994 (N_6994,N_5154,N_5888);
and U6995 (N_6995,N_5672,N_5787);
nand U6996 (N_6996,N_5255,N_5319);
and U6997 (N_6997,N_5156,N_5891);
nand U6998 (N_6998,N_5498,N_5027);
and U6999 (N_6999,N_5984,N_5456);
or U7000 (N_7000,N_6291,N_6779);
nor U7001 (N_7001,N_6127,N_6758);
nand U7002 (N_7002,N_6745,N_6713);
nand U7003 (N_7003,N_6054,N_6123);
and U7004 (N_7004,N_6289,N_6018);
or U7005 (N_7005,N_6964,N_6366);
xnor U7006 (N_7006,N_6064,N_6514);
nor U7007 (N_7007,N_6029,N_6844);
xor U7008 (N_7008,N_6309,N_6489);
or U7009 (N_7009,N_6037,N_6194);
and U7010 (N_7010,N_6626,N_6902);
nand U7011 (N_7011,N_6735,N_6606);
or U7012 (N_7012,N_6683,N_6337);
or U7013 (N_7013,N_6100,N_6004);
nand U7014 (N_7014,N_6015,N_6109);
or U7015 (N_7015,N_6173,N_6768);
xnor U7016 (N_7016,N_6619,N_6988);
or U7017 (N_7017,N_6885,N_6142);
nor U7018 (N_7018,N_6915,N_6012);
nand U7019 (N_7019,N_6655,N_6716);
or U7020 (N_7020,N_6958,N_6536);
or U7021 (N_7021,N_6718,N_6043);
nor U7022 (N_7022,N_6107,N_6339);
nor U7023 (N_7023,N_6263,N_6546);
nor U7024 (N_7024,N_6290,N_6597);
nand U7025 (N_7025,N_6265,N_6368);
xor U7026 (N_7026,N_6464,N_6687);
nand U7027 (N_7027,N_6517,N_6962);
or U7028 (N_7028,N_6350,N_6829);
xor U7029 (N_7029,N_6407,N_6007);
xor U7030 (N_7030,N_6643,N_6056);
or U7031 (N_7031,N_6277,N_6948);
xnor U7032 (N_7032,N_6956,N_6944);
or U7033 (N_7033,N_6845,N_6518);
xor U7034 (N_7034,N_6893,N_6434);
nand U7035 (N_7035,N_6828,N_6761);
nand U7036 (N_7036,N_6231,N_6719);
nand U7037 (N_7037,N_6520,N_6177);
nor U7038 (N_7038,N_6091,N_6787);
nor U7039 (N_7039,N_6651,N_6608);
or U7040 (N_7040,N_6117,N_6225);
and U7041 (N_7041,N_6537,N_6444);
xor U7042 (N_7042,N_6771,N_6542);
or U7043 (N_7043,N_6452,N_6961);
nand U7044 (N_7044,N_6191,N_6299);
xor U7045 (N_7045,N_6180,N_6280);
nand U7046 (N_7046,N_6135,N_6394);
and U7047 (N_7047,N_6121,N_6507);
nand U7048 (N_7048,N_6929,N_6181);
xor U7049 (N_7049,N_6255,N_6087);
nand U7050 (N_7050,N_6752,N_6805);
and U7051 (N_7051,N_6631,N_6302);
and U7052 (N_7052,N_6106,N_6157);
or U7053 (N_7053,N_6044,N_6788);
nand U7054 (N_7054,N_6273,N_6074);
or U7055 (N_7055,N_6101,N_6497);
nand U7056 (N_7056,N_6413,N_6659);
nor U7057 (N_7057,N_6818,N_6021);
nor U7058 (N_7058,N_6780,N_6221);
xnor U7059 (N_7059,N_6529,N_6877);
nand U7060 (N_7060,N_6022,N_6184);
xnor U7061 (N_7061,N_6275,N_6873);
or U7062 (N_7062,N_6859,N_6333);
nor U7063 (N_7063,N_6588,N_6675);
nand U7064 (N_7064,N_6065,N_6389);
and U7065 (N_7065,N_6010,N_6344);
or U7066 (N_7066,N_6623,N_6704);
or U7067 (N_7067,N_6381,N_6865);
nor U7068 (N_7068,N_6459,N_6308);
and U7069 (N_7069,N_6419,N_6693);
nand U7070 (N_7070,N_6611,N_6484);
nand U7071 (N_7071,N_6806,N_6930);
xor U7072 (N_7072,N_6324,N_6025);
or U7073 (N_7073,N_6223,N_6667);
and U7074 (N_7074,N_6269,N_6808);
nor U7075 (N_7075,N_6923,N_6750);
or U7076 (N_7076,N_6951,N_6345);
nand U7077 (N_7077,N_6601,N_6083);
nor U7078 (N_7078,N_6682,N_6454);
or U7079 (N_7079,N_6229,N_6193);
and U7080 (N_7080,N_6851,N_6629);
or U7081 (N_7081,N_6617,N_6285);
nand U7082 (N_7082,N_6460,N_6802);
xnor U7083 (N_7083,N_6813,N_6075);
nand U7084 (N_7084,N_6001,N_6848);
xor U7085 (N_7085,N_6803,N_6421);
nor U7086 (N_7086,N_6531,N_6641);
or U7087 (N_7087,N_6941,N_6110);
xnor U7088 (N_7088,N_6053,N_6932);
and U7089 (N_7089,N_6038,N_6981);
or U7090 (N_7090,N_6039,N_6268);
nor U7091 (N_7091,N_6365,N_6170);
or U7092 (N_7092,N_6028,N_6952);
nand U7093 (N_7093,N_6373,N_6737);
xnor U7094 (N_7094,N_6799,N_6097);
nand U7095 (N_7095,N_6792,N_6842);
xnor U7096 (N_7096,N_6510,N_6816);
or U7097 (N_7097,N_6418,N_6080);
nor U7098 (N_7098,N_6032,N_6662);
and U7099 (N_7099,N_6040,N_6371);
xor U7100 (N_7100,N_6296,N_6111);
or U7101 (N_7101,N_6736,N_6685);
and U7102 (N_7102,N_6436,N_6959);
and U7103 (N_7103,N_6896,N_6971);
nand U7104 (N_7104,N_6831,N_6890);
xor U7105 (N_7105,N_6622,N_6823);
nor U7106 (N_7106,N_6953,N_6041);
xnor U7107 (N_7107,N_6209,N_6156);
and U7108 (N_7108,N_6722,N_6994);
and U7109 (N_7109,N_6329,N_6336);
xnor U7110 (N_7110,N_6585,N_6566);
xnor U7111 (N_7111,N_6487,N_6208);
and U7112 (N_7112,N_6131,N_6774);
and U7113 (N_7113,N_6306,N_6534);
xor U7114 (N_7114,N_6462,N_6702);
and U7115 (N_7115,N_6978,N_6997);
nor U7116 (N_7116,N_6166,N_6378);
nand U7117 (N_7117,N_6319,N_6504);
nand U7118 (N_7118,N_6068,N_6471);
xnor U7119 (N_7119,N_6082,N_6164);
xor U7120 (N_7120,N_6649,N_6133);
nor U7121 (N_7121,N_6599,N_6513);
or U7122 (N_7122,N_6917,N_6179);
nor U7123 (N_7123,N_6925,N_6212);
or U7124 (N_7124,N_6732,N_6690);
or U7125 (N_7125,N_6213,N_6600);
and U7126 (N_7126,N_6526,N_6821);
or U7127 (N_7127,N_6453,N_6232);
or U7128 (N_7128,N_6791,N_6969);
and U7129 (N_7129,N_6063,N_6077);
or U7130 (N_7130,N_6099,N_6402);
xor U7131 (N_7131,N_6415,N_6211);
xor U7132 (N_7132,N_6924,N_6256);
nor U7133 (N_7133,N_6798,N_6440);
and U7134 (N_7134,N_6122,N_6466);
and U7135 (N_7135,N_6343,N_6697);
and U7136 (N_7136,N_6253,N_6559);
nand U7137 (N_7137,N_6363,N_6910);
and U7138 (N_7138,N_6814,N_6618);
xnor U7139 (N_7139,N_6547,N_6246);
xnor U7140 (N_7140,N_6423,N_6238);
xnor U7141 (N_7141,N_6207,N_6695);
or U7142 (N_7142,N_6933,N_6922);
and U7143 (N_7143,N_6137,N_6898);
nor U7144 (N_7144,N_6954,N_6615);
or U7145 (N_7145,N_6605,N_6321);
xnor U7146 (N_7146,N_6642,N_6957);
nor U7147 (N_7147,N_6377,N_6790);
nand U7148 (N_7148,N_6551,N_6867);
and U7149 (N_7149,N_6376,N_6461);
and U7150 (N_7150,N_6432,N_6847);
nand U7151 (N_7151,N_6495,N_6852);
and U7152 (N_7152,N_6351,N_6627);
nor U7153 (N_7153,N_6151,N_6927);
xor U7154 (N_7154,N_6398,N_6721);
xnor U7155 (N_7155,N_6793,N_6195);
nor U7156 (N_7156,N_6201,N_6854);
nand U7157 (N_7157,N_6677,N_6580);
or U7158 (N_7158,N_6125,N_6729);
and U7159 (N_7159,N_6789,N_6202);
xnor U7160 (N_7160,N_6522,N_6086);
nor U7161 (N_7161,N_6476,N_6731);
or U7162 (N_7162,N_6717,N_6680);
or U7163 (N_7163,N_6352,N_6889);
or U7164 (N_7164,N_6769,N_6260);
nand U7165 (N_7165,N_6970,N_6807);
nor U7166 (N_7166,N_6034,N_6668);
and U7167 (N_7167,N_6516,N_6139);
xor U7168 (N_7168,N_6741,N_6553);
nor U7169 (N_7169,N_6616,N_6167);
or U7170 (N_7170,N_6341,N_6017);
or U7171 (N_7171,N_6447,N_6119);
and U7172 (N_7172,N_6115,N_6678);
or U7173 (N_7173,N_6832,N_6382);
and U7174 (N_7174,N_6420,N_6822);
or U7175 (N_7175,N_6215,N_6856);
or U7176 (N_7176,N_6129,N_6408);
and U7177 (N_7177,N_6442,N_6475);
nor U7178 (N_7178,N_6422,N_6846);
or U7179 (N_7179,N_6493,N_6036);
nor U7180 (N_7180,N_6470,N_6488);
nand U7181 (N_7181,N_6491,N_6092);
nand U7182 (N_7182,N_6556,N_6456);
nor U7183 (N_7183,N_6661,N_6590);
nand U7184 (N_7184,N_6767,N_6334);
and U7185 (N_7185,N_6349,N_6955);
or U7186 (N_7186,N_6375,N_6240);
and U7187 (N_7187,N_6163,N_6236);
nand U7188 (N_7188,N_6148,N_6938);
nand U7189 (N_7189,N_6070,N_6786);
xnor U7190 (N_7190,N_6234,N_6384);
and U7191 (N_7191,N_6259,N_6301);
xor U7192 (N_7192,N_6937,N_6120);
nand U7193 (N_7193,N_6742,N_6326);
or U7194 (N_7194,N_6748,N_6498);
or U7195 (N_7195,N_6013,N_6975);
and U7196 (N_7196,N_6328,N_6632);
or U7197 (N_7197,N_6354,N_6250);
nor U7198 (N_7198,N_6689,N_6648);
or U7199 (N_7199,N_6548,N_6950);
nor U7200 (N_7200,N_6228,N_6985);
xor U7201 (N_7201,N_6297,N_6401);
nand U7202 (N_7202,N_6835,N_6132);
and U7203 (N_7203,N_6282,N_6026);
xnor U7204 (N_7204,N_6294,N_6186);
nor U7205 (N_7205,N_6433,N_6663);
nor U7206 (N_7206,N_6380,N_6620);
and U7207 (N_7207,N_6860,N_6102);
nor U7208 (N_7208,N_6149,N_6754);
nand U7209 (N_7209,N_6050,N_6206);
nand U7210 (N_7210,N_6155,N_6593);
xor U7211 (N_7211,N_6411,N_6533);
nand U7212 (N_7212,N_6914,N_6176);
nand U7213 (N_7213,N_6760,N_6314);
or U7214 (N_7214,N_6113,N_6843);
or U7215 (N_7215,N_6499,N_6224);
xor U7216 (N_7216,N_6508,N_6968);
xor U7217 (N_7217,N_6020,N_6869);
or U7218 (N_7218,N_6174,N_6078);
xor U7219 (N_7219,N_6219,N_6490);
xor U7220 (N_7220,N_6200,N_6205);
and U7221 (N_7221,N_6243,N_6909);
or U7222 (N_7222,N_6574,N_6359);
or U7223 (N_7223,N_6185,N_6960);
or U7224 (N_7224,N_6973,N_6839);
or U7225 (N_7225,N_6128,N_6435);
or U7226 (N_7226,N_6670,N_6169);
xor U7227 (N_7227,N_6540,N_6469);
xnor U7228 (N_7228,N_6563,N_6587);
xnor U7229 (N_7229,N_6947,N_6494);
and U7230 (N_7230,N_6126,N_6582);
xnor U7231 (N_7231,N_6059,N_6607);
and U7232 (N_7232,N_6784,N_6819);
nand U7233 (N_7233,N_6226,N_6857);
nand U7234 (N_7234,N_6963,N_6316);
xnor U7235 (N_7235,N_6740,N_6465);
or U7236 (N_7236,N_6257,N_6147);
or U7237 (N_7237,N_6134,N_6136);
nand U7238 (N_7238,N_6372,N_6198);
nor U7239 (N_7239,N_6726,N_6899);
nor U7240 (N_7240,N_6841,N_6654);
xnor U7241 (N_7241,N_6430,N_6781);
and U7242 (N_7242,N_6364,N_6448);
and U7243 (N_7243,N_6438,N_6485);
xor U7244 (N_7244,N_6666,N_6610);
or U7245 (N_7245,N_6390,N_6628);
xnor U7246 (N_7246,N_6239,N_6613);
or U7247 (N_7247,N_6210,N_6313);
nand U7248 (N_7248,N_6458,N_6974);
nand U7249 (N_7249,N_6045,N_6393);
nor U7250 (N_7250,N_6035,N_6332);
xor U7251 (N_7251,N_6323,N_6870);
nand U7252 (N_7252,N_6451,N_6284);
or U7253 (N_7253,N_6227,N_6235);
xnor U7254 (N_7254,N_6369,N_6983);
or U7255 (N_7255,N_6812,N_6995);
or U7256 (N_7256,N_6278,N_6783);
nand U7257 (N_7257,N_6863,N_6303);
nor U7258 (N_7258,N_6358,N_6673);
nor U7259 (N_7259,N_6016,N_6967);
and U7260 (N_7260,N_6160,N_6700);
nand U7261 (N_7261,N_6446,N_6604);
and U7262 (N_7262,N_6698,N_6271);
xnor U7263 (N_7263,N_6990,N_6357);
xnor U7264 (N_7264,N_6984,N_6449);
nand U7265 (N_7265,N_6864,N_6711);
nand U7266 (N_7266,N_6244,N_6385);
nand U7267 (N_7267,N_6576,N_6088);
xnor U7268 (N_7268,N_6886,N_6738);
nand U7269 (N_7269,N_6935,N_6921);
or U7270 (N_7270,N_6425,N_6871);
or U7271 (N_7271,N_6347,N_6108);
xor U7272 (N_7272,N_6501,N_6757);
xnor U7273 (N_7273,N_6320,N_6443);
and U7274 (N_7274,N_6577,N_6809);
and U7275 (N_7275,N_6005,N_6072);
nand U7276 (N_7276,N_6804,N_6006);
or U7277 (N_7277,N_6340,N_6614);
nand U7278 (N_7278,N_6674,N_6424);
nand U7279 (N_7279,N_6178,N_6633);
and U7280 (N_7280,N_6573,N_6230);
or U7281 (N_7281,N_6245,N_6116);
nand U7282 (N_7282,N_6824,N_6248);
nand U7283 (N_7283,N_6753,N_6724);
nand U7284 (N_7284,N_6159,N_6154);
and U7285 (N_7285,N_6400,N_6646);
nor U7286 (N_7286,N_6410,N_6450);
or U7287 (N_7287,N_6705,N_6647);
or U7288 (N_7288,N_6062,N_6901);
and U7289 (N_7289,N_6024,N_6171);
nand U7290 (N_7290,N_6532,N_6908);
xor U7291 (N_7291,N_6067,N_6165);
nor U7292 (N_7292,N_6817,N_6725);
and U7293 (N_7293,N_6966,N_6437);
xor U7294 (N_7294,N_6874,N_6850);
or U7295 (N_7295,N_6298,N_6153);
or U7296 (N_7296,N_6479,N_6557);
nand U7297 (N_7297,N_6706,N_6946);
nand U7298 (N_7298,N_6189,N_6730);
nor U7299 (N_7299,N_6766,N_6478);
nand U7300 (N_7300,N_6635,N_6515);
nand U7301 (N_7301,N_6355,N_6746);
or U7302 (N_7302,N_6999,N_6940);
xor U7303 (N_7303,N_6720,N_6887);
and U7304 (N_7304,N_6891,N_6868);
and U7305 (N_7305,N_6085,N_6307);
nand U7306 (N_7306,N_6318,N_6431);
nand U7307 (N_7307,N_6744,N_6058);
nor U7308 (N_7308,N_6912,N_6103);
nand U7309 (N_7309,N_6942,N_6145);
nand U7310 (N_7310,N_6042,N_6696);
nand U7311 (N_7311,N_6609,N_6405);
or U7312 (N_7312,N_6519,N_6703);
nand U7313 (N_7313,N_6486,N_6892);
or U7314 (N_7314,N_6895,N_6247);
nor U7315 (N_7315,N_6827,N_6777);
nand U7316 (N_7316,N_6342,N_6701);
or U7317 (N_7317,N_6500,N_6778);
xor U7318 (N_7318,N_6882,N_6338);
xnor U7319 (N_7319,N_6217,N_6637);
nor U7320 (N_7320,N_6644,N_6759);
xnor U7321 (N_7321,N_6564,N_6203);
nor U7322 (N_7322,N_6876,N_6233);
nor U7323 (N_7323,N_6567,N_6918);
xnor U7324 (N_7324,N_6114,N_6279);
or U7325 (N_7325,N_6992,N_6688);
and U7326 (N_7326,N_6652,N_6492);
nor U7327 (N_7327,N_6764,N_6412);
xnor U7328 (N_7328,N_6027,N_6237);
or U7329 (N_7329,N_6292,N_6304);
and U7330 (N_7330,N_6482,N_6589);
nand U7331 (N_7331,N_6747,N_6977);
nand U7332 (N_7332,N_6315,N_6911);
xnor U7333 (N_7333,N_6218,N_6562);
nor U7334 (N_7334,N_6763,N_6158);
or U7335 (N_7335,N_6252,N_6653);
or U7336 (N_7336,N_6884,N_6011);
or U7337 (N_7337,N_6672,N_6660);
and U7338 (N_7338,N_6069,N_6055);
or U7339 (N_7339,N_6976,N_6472);
and U7340 (N_7340,N_6140,N_6665);
and U7341 (N_7341,N_6524,N_6266);
or U7342 (N_7342,N_6993,N_6888);
nor U7343 (N_7343,N_6048,N_6270);
nor U7344 (N_7344,N_6676,N_6919);
xor U7345 (N_7345,N_6991,N_6723);
nand U7346 (N_7346,N_6880,N_6739);
nand U7347 (N_7347,N_6710,N_6949);
xor U7348 (N_7348,N_6003,N_6033);
nor U7349 (N_7349,N_6595,N_6503);
or U7350 (N_7350,N_6283,N_6386);
xnor U7351 (N_7351,N_6810,N_6785);
nor U7352 (N_7352,N_6709,N_6441);
or U7353 (N_7353,N_6945,N_6335);
nor U7354 (N_7354,N_6467,N_6090);
xnor U7355 (N_7355,N_6571,N_6249);
and U7356 (N_7356,N_6681,N_6552);
xor U7357 (N_7357,N_6311,N_6658);
nand U7358 (N_7358,N_6794,N_6530);
nor U7359 (N_7359,N_6903,N_6762);
or U7360 (N_7360,N_6776,N_6811);
nor U7361 (N_7361,N_6905,N_6241);
nor U7362 (N_7362,N_6544,N_6391);
xnor U7363 (N_7363,N_6965,N_6047);
or U7364 (N_7364,N_6496,N_6286);
and U7365 (N_7365,N_6192,N_6612);
nand U7366 (N_7366,N_6220,N_6980);
nor U7367 (N_7367,N_6076,N_6775);
or U7368 (N_7368,N_6554,N_6019);
nand U7369 (N_7369,N_6066,N_6686);
xor U7370 (N_7370,N_6162,N_6144);
nor U7371 (N_7371,N_6214,N_6645);
and U7372 (N_7372,N_6071,N_6428);
and U7373 (N_7373,N_6457,N_6348);
nand U7374 (N_7374,N_6861,N_6906);
xnor U7375 (N_7375,N_6715,N_6057);
nor U7376 (N_7376,N_6883,N_6468);
xor U7377 (N_7377,N_6000,N_6124);
nand U7378 (N_7378,N_6800,N_6541);
xnor U7379 (N_7379,N_6679,N_6833);
nor U7380 (N_7380,N_6765,N_6477);
xnor U7381 (N_7381,N_6579,N_6356);
or U7382 (N_7382,N_6404,N_6330);
or U7383 (N_7383,N_6826,N_6743);
or U7384 (N_7384,N_6295,N_6455);
nor U7385 (N_7385,N_6801,N_6555);
xor U7386 (N_7386,N_6782,N_6161);
nand U7387 (N_7387,N_6545,N_6879);
nand U7388 (N_7388,N_6836,N_6288);
and U7389 (N_7389,N_6426,N_6592);
nor U7390 (N_7390,N_6858,N_6527);
xor U7391 (N_7391,N_6853,N_6671);
xnor U7392 (N_7392,N_6094,N_6222);
or U7393 (N_7393,N_6897,N_6361);
nor U7394 (N_7394,N_6657,N_6261);
nand U7395 (N_7395,N_6276,N_6374);
nand U7396 (N_7396,N_6838,N_6692);
or U7397 (N_7397,N_6112,N_6403);
or U7398 (N_7398,N_6150,N_6264);
xor U7399 (N_7399,N_6664,N_6862);
or U7400 (N_7400,N_6712,N_6098);
or U7401 (N_7401,N_6009,N_6928);
and U7402 (N_7402,N_6242,N_6281);
nand U7403 (N_7403,N_6439,N_6581);
nor U7404 (N_7404,N_6797,N_6152);
xnor U7405 (N_7405,N_6322,N_6727);
xor U7406 (N_7406,N_6406,N_6190);
nand U7407 (N_7407,N_6502,N_6998);
nor U7408 (N_7408,N_6815,N_6528);
or U7409 (N_7409,N_6598,N_6849);
xor U7410 (N_7410,N_6300,N_6584);
nor U7411 (N_7411,N_6197,N_6429);
and U7412 (N_7412,N_6168,N_6575);
and U7413 (N_7413,N_6691,N_6093);
xor U7414 (N_7414,N_6987,N_6521);
nor U7415 (N_7415,N_6982,N_6199);
or U7416 (N_7416,N_6525,N_6561);
nand U7417 (N_7417,N_6830,N_6014);
nand U7418 (N_7418,N_6820,N_6603);
nor U7419 (N_7419,N_6293,N_6872);
nor U7420 (N_7420,N_6639,N_6578);
or U7421 (N_7421,N_6511,N_6558);
nand U7422 (N_7422,N_6325,N_6141);
and U7423 (N_7423,N_6770,N_6346);
nand U7424 (N_7424,N_6287,N_6379);
xor U7425 (N_7425,N_6926,N_6638);
nand U7426 (N_7426,N_6772,N_6630);
xnor U7427 (N_7427,N_6512,N_6734);
xor U7428 (N_7428,N_6550,N_6353);
or U7429 (N_7429,N_6931,N_6105);
nor U7430 (N_7430,N_6188,N_6414);
nand U7431 (N_7431,N_6023,N_6370);
or U7432 (N_7432,N_6570,N_6894);
and U7433 (N_7433,N_6907,N_6095);
nor U7434 (N_7434,N_6881,N_6146);
and U7435 (N_7435,N_6262,N_6568);
or U7436 (N_7436,N_6254,N_6473);
nor U7437 (N_7437,N_6416,N_6539);
nand U7438 (N_7438,N_6834,N_6594);
and U7439 (N_7439,N_6104,N_6621);
xnor U7440 (N_7440,N_6187,N_6796);
or U7441 (N_7441,N_6943,N_6360);
xnor U7442 (N_7442,N_6474,N_6182);
xnor U7443 (N_7443,N_6138,N_6640);
or U7444 (N_7444,N_6840,N_6031);
nor U7445 (N_7445,N_6312,N_6979);
nand U7446 (N_7446,N_6397,N_6934);
nor U7447 (N_7447,N_6175,N_6445);
nor U7448 (N_7448,N_6387,N_6543);
xnor U7449 (N_7449,N_6591,N_6272);
nand U7450 (N_7450,N_6396,N_6751);
xor U7451 (N_7451,N_6707,N_6523);
nand U7452 (N_7452,N_6046,N_6096);
xor U7453 (N_7453,N_6388,N_6084);
nor U7454 (N_7454,N_6305,N_6936);
nand U7455 (N_7455,N_6773,N_6258);
xor U7456 (N_7456,N_6383,N_6395);
and U7457 (N_7457,N_6251,N_6008);
nor U7458 (N_7458,N_6060,N_6756);
and U7459 (N_7459,N_6733,N_6392);
xor U7460 (N_7460,N_6939,N_6216);
nand U7461 (N_7461,N_6549,N_6030);
or U7462 (N_7462,N_6052,N_6538);
or U7463 (N_7463,N_6602,N_6427);
and U7464 (N_7464,N_6572,N_6204);
or U7465 (N_7465,N_6081,N_6708);
nand U7466 (N_7466,N_6505,N_6728);
xnor U7467 (N_7467,N_6586,N_6634);
nor U7468 (N_7468,N_6183,N_6051);
nand U7469 (N_7469,N_6118,N_6310);
and U7470 (N_7470,N_6904,N_6920);
xnor U7471 (N_7471,N_6143,N_6972);
nand U7472 (N_7472,N_6274,N_6506);
nor U7473 (N_7473,N_6509,N_6986);
or U7474 (N_7474,N_6327,N_6900);
and U7475 (N_7475,N_6755,N_6694);
and U7476 (N_7476,N_6989,N_6362);
or U7477 (N_7477,N_6656,N_6699);
nor U7478 (N_7478,N_6875,N_6684);
and U7479 (N_7479,N_6130,N_6073);
nor U7480 (N_7480,N_6855,N_6913);
xor U7481 (N_7481,N_6267,N_6866);
or U7482 (N_7482,N_6565,N_6002);
nor U7483 (N_7483,N_6916,N_6399);
and U7484 (N_7484,N_6569,N_6624);
nand U7485 (N_7485,N_6463,N_6172);
nand U7486 (N_7486,N_6560,N_6196);
nand U7487 (N_7487,N_6480,N_6417);
xor U7488 (N_7488,N_6481,N_6878);
nand U7489 (N_7489,N_6650,N_6317);
and U7490 (N_7490,N_6367,N_6483);
or U7491 (N_7491,N_6089,N_6331);
nand U7492 (N_7492,N_6061,N_6996);
xor U7493 (N_7493,N_6636,N_6535);
and U7494 (N_7494,N_6749,N_6825);
nor U7495 (N_7495,N_6583,N_6837);
nand U7496 (N_7496,N_6596,N_6049);
nor U7497 (N_7497,N_6669,N_6795);
and U7498 (N_7498,N_6409,N_6714);
nor U7499 (N_7499,N_6625,N_6079);
or U7500 (N_7500,N_6475,N_6449);
nand U7501 (N_7501,N_6850,N_6891);
nor U7502 (N_7502,N_6671,N_6043);
or U7503 (N_7503,N_6646,N_6252);
or U7504 (N_7504,N_6796,N_6439);
and U7505 (N_7505,N_6592,N_6440);
and U7506 (N_7506,N_6888,N_6975);
nor U7507 (N_7507,N_6222,N_6774);
and U7508 (N_7508,N_6738,N_6700);
xor U7509 (N_7509,N_6651,N_6243);
or U7510 (N_7510,N_6734,N_6259);
or U7511 (N_7511,N_6963,N_6101);
and U7512 (N_7512,N_6061,N_6960);
nand U7513 (N_7513,N_6596,N_6693);
nand U7514 (N_7514,N_6855,N_6337);
or U7515 (N_7515,N_6523,N_6130);
xor U7516 (N_7516,N_6936,N_6926);
nand U7517 (N_7517,N_6542,N_6070);
and U7518 (N_7518,N_6175,N_6823);
or U7519 (N_7519,N_6681,N_6014);
or U7520 (N_7520,N_6684,N_6394);
and U7521 (N_7521,N_6440,N_6228);
nand U7522 (N_7522,N_6324,N_6523);
nor U7523 (N_7523,N_6078,N_6425);
and U7524 (N_7524,N_6440,N_6632);
nor U7525 (N_7525,N_6284,N_6290);
or U7526 (N_7526,N_6779,N_6439);
and U7527 (N_7527,N_6718,N_6340);
and U7528 (N_7528,N_6281,N_6511);
nand U7529 (N_7529,N_6950,N_6823);
nand U7530 (N_7530,N_6115,N_6783);
or U7531 (N_7531,N_6624,N_6954);
or U7532 (N_7532,N_6605,N_6375);
nor U7533 (N_7533,N_6532,N_6661);
and U7534 (N_7534,N_6152,N_6740);
xor U7535 (N_7535,N_6924,N_6486);
nand U7536 (N_7536,N_6664,N_6499);
nand U7537 (N_7537,N_6922,N_6377);
and U7538 (N_7538,N_6858,N_6978);
nor U7539 (N_7539,N_6466,N_6727);
nand U7540 (N_7540,N_6243,N_6633);
nor U7541 (N_7541,N_6779,N_6410);
and U7542 (N_7542,N_6289,N_6371);
xor U7543 (N_7543,N_6077,N_6352);
nand U7544 (N_7544,N_6124,N_6901);
nor U7545 (N_7545,N_6050,N_6259);
and U7546 (N_7546,N_6470,N_6806);
or U7547 (N_7547,N_6128,N_6194);
nor U7548 (N_7548,N_6915,N_6882);
nand U7549 (N_7549,N_6053,N_6214);
and U7550 (N_7550,N_6313,N_6992);
xor U7551 (N_7551,N_6496,N_6541);
xnor U7552 (N_7552,N_6070,N_6469);
xor U7553 (N_7553,N_6805,N_6690);
nor U7554 (N_7554,N_6737,N_6181);
xnor U7555 (N_7555,N_6198,N_6808);
nand U7556 (N_7556,N_6429,N_6790);
and U7557 (N_7557,N_6219,N_6667);
or U7558 (N_7558,N_6825,N_6338);
nor U7559 (N_7559,N_6823,N_6751);
xnor U7560 (N_7560,N_6358,N_6337);
and U7561 (N_7561,N_6694,N_6021);
and U7562 (N_7562,N_6365,N_6226);
and U7563 (N_7563,N_6053,N_6815);
and U7564 (N_7564,N_6728,N_6057);
nand U7565 (N_7565,N_6122,N_6727);
or U7566 (N_7566,N_6616,N_6575);
nor U7567 (N_7567,N_6390,N_6847);
xor U7568 (N_7568,N_6111,N_6118);
and U7569 (N_7569,N_6942,N_6752);
xnor U7570 (N_7570,N_6725,N_6061);
nand U7571 (N_7571,N_6129,N_6028);
xnor U7572 (N_7572,N_6778,N_6438);
or U7573 (N_7573,N_6645,N_6461);
nor U7574 (N_7574,N_6463,N_6366);
or U7575 (N_7575,N_6245,N_6431);
and U7576 (N_7576,N_6843,N_6123);
nand U7577 (N_7577,N_6691,N_6973);
nand U7578 (N_7578,N_6834,N_6232);
nor U7579 (N_7579,N_6018,N_6228);
or U7580 (N_7580,N_6888,N_6764);
nor U7581 (N_7581,N_6787,N_6751);
xor U7582 (N_7582,N_6054,N_6235);
or U7583 (N_7583,N_6782,N_6474);
xor U7584 (N_7584,N_6114,N_6416);
nor U7585 (N_7585,N_6679,N_6197);
or U7586 (N_7586,N_6027,N_6142);
and U7587 (N_7587,N_6872,N_6825);
nand U7588 (N_7588,N_6557,N_6343);
or U7589 (N_7589,N_6801,N_6478);
and U7590 (N_7590,N_6300,N_6603);
and U7591 (N_7591,N_6555,N_6084);
nor U7592 (N_7592,N_6472,N_6936);
xor U7593 (N_7593,N_6376,N_6457);
and U7594 (N_7594,N_6327,N_6509);
nor U7595 (N_7595,N_6487,N_6834);
nor U7596 (N_7596,N_6871,N_6843);
or U7597 (N_7597,N_6212,N_6737);
and U7598 (N_7598,N_6843,N_6709);
xnor U7599 (N_7599,N_6964,N_6027);
xnor U7600 (N_7600,N_6795,N_6620);
or U7601 (N_7601,N_6999,N_6743);
nand U7602 (N_7602,N_6583,N_6054);
xor U7603 (N_7603,N_6895,N_6141);
and U7604 (N_7604,N_6478,N_6021);
nand U7605 (N_7605,N_6477,N_6668);
nor U7606 (N_7606,N_6759,N_6428);
or U7607 (N_7607,N_6794,N_6225);
and U7608 (N_7608,N_6963,N_6952);
nand U7609 (N_7609,N_6293,N_6108);
nand U7610 (N_7610,N_6418,N_6120);
nor U7611 (N_7611,N_6721,N_6373);
and U7612 (N_7612,N_6547,N_6925);
nand U7613 (N_7613,N_6751,N_6859);
xnor U7614 (N_7614,N_6906,N_6865);
nand U7615 (N_7615,N_6714,N_6126);
and U7616 (N_7616,N_6227,N_6030);
or U7617 (N_7617,N_6875,N_6076);
xnor U7618 (N_7618,N_6280,N_6681);
or U7619 (N_7619,N_6000,N_6223);
and U7620 (N_7620,N_6011,N_6851);
nand U7621 (N_7621,N_6281,N_6151);
and U7622 (N_7622,N_6065,N_6884);
and U7623 (N_7623,N_6363,N_6778);
xor U7624 (N_7624,N_6075,N_6798);
xor U7625 (N_7625,N_6080,N_6684);
xnor U7626 (N_7626,N_6214,N_6430);
xor U7627 (N_7627,N_6077,N_6933);
nand U7628 (N_7628,N_6385,N_6825);
nand U7629 (N_7629,N_6559,N_6353);
xnor U7630 (N_7630,N_6665,N_6862);
or U7631 (N_7631,N_6819,N_6630);
xnor U7632 (N_7632,N_6587,N_6876);
and U7633 (N_7633,N_6492,N_6334);
nand U7634 (N_7634,N_6345,N_6914);
or U7635 (N_7635,N_6228,N_6711);
and U7636 (N_7636,N_6199,N_6845);
and U7637 (N_7637,N_6321,N_6153);
and U7638 (N_7638,N_6668,N_6086);
nor U7639 (N_7639,N_6770,N_6309);
xor U7640 (N_7640,N_6481,N_6562);
or U7641 (N_7641,N_6761,N_6721);
nor U7642 (N_7642,N_6201,N_6953);
nand U7643 (N_7643,N_6527,N_6879);
nor U7644 (N_7644,N_6194,N_6473);
nand U7645 (N_7645,N_6020,N_6758);
xnor U7646 (N_7646,N_6006,N_6879);
nor U7647 (N_7647,N_6368,N_6627);
nor U7648 (N_7648,N_6563,N_6244);
xor U7649 (N_7649,N_6917,N_6301);
or U7650 (N_7650,N_6467,N_6205);
xor U7651 (N_7651,N_6079,N_6498);
xor U7652 (N_7652,N_6902,N_6236);
or U7653 (N_7653,N_6775,N_6967);
nor U7654 (N_7654,N_6604,N_6838);
nand U7655 (N_7655,N_6421,N_6594);
xor U7656 (N_7656,N_6481,N_6758);
and U7657 (N_7657,N_6686,N_6221);
nor U7658 (N_7658,N_6393,N_6525);
and U7659 (N_7659,N_6112,N_6500);
or U7660 (N_7660,N_6851,N_6509);
nand U7661 (N_7661,N_6237,N_6174);
or U7662 (N_7662,N_6466,N_6424);
or U7663 (N_7663,N_6332,N_6625);
and U7664 (N_7664,N_6185,N_6739);
or U7665 (N_7665,N_6313,N_6501);
nand U7666 (N_7666,N_6623,N_6527);
xnor U7667 (N_7667,N_6035,N_6389);
nand U7668 (N_7668,N_6590,N_6089);
and U7669 (N_7669,N_6987,N_6939);
nand U7670 (N_7670,N_6379,N_6094);
and U7671 (N_7671,N_6981,N_6032);
and U7672 (N_7672,N_6935,N_6754);
or U7673 (N_7673,N_6513,N_6690);
and U7674 (N_7674,N_6254,N_6175);
xor U7675 (N_7675,N_6789,N_6674);
nor U7676 (N_7676,N_6465,N_6449);
xor U7677 (N_7677,N_6651,N_6266);
and U7678 (N_7678,N_6629,N_6357);
or U7679 (N_7679,N_6255,N_6167);
nor U7680 (N_7680,N_6245,N_6623);
xor U7681 (N_7681,N_6753,N_6915);
nor U7682 (N_7682,N_6527,N_6437);
nand U7683 (N_7683,N_6190,N_6268);
xnor U7684 (N_7684,N_6819,N_6274);
nand U7685 (N_7685,N_6365,N_6034);
xnor U7686 (N_7686,N_6805,N_6366);
nand U7687 (N_7687,N_6294,N_6950);
nand U7688 (N_7688,N_6829,N_6323);
nor U7689 (N_7689,N_6944,N_6497);
nor U7690 (N_7690,N_6315,N_6965);
and U7691 (N_7691,N_6559,N_6217);
or U7692 (N_7692,N_6237,N_6083);
nand U7693 (N_7693,N_6140,N_6313);
or U7694 (N_7694,N_6312,N_6862);
nor U7695 (N_7695,N_6580,N_6978);
xnor U7696 (N_7696,N_6472,N_6315);
nor U7697 (N_7697,N_6875,N_6047);
and U7698 (N_7698,N_6928,N_6217);
and U7699 (N_7699,N_6165,N_6194);
and U7700 (N_7700,N_6293,N_6533);
nor U7701 (N_7701,N_6297,N_6446);
or U7702 (N_7702,N_6785,N_6733);
or U7703 (N_7703,N_6371,N_6359);
xnor U7704 (N_7704,N_6305,N_6849);
nor U7705 (N_7705,N_6519,N_6813);
nand U7706 (N_7706,N_6303,N_6172);
and U7707 (N_7707,N_6784,N_6654);
or U7708 (N_7708,N_6860,N_6080);
nor U7709 (N_7709,N_6129,N_6811);
or U7710 (N_7710,N_6212,N_6159);
and U7711 (N_7711,N_6723,N_6204);
and U7712 (N_7712,N_6018,N_6440);
or U7713 (N_7713,N_6369,N_6587);
or U7714 (N_7714,N_6258,N_6420);
nor U7715 (N_7715,N_6950,N_6639);
nor U7716 (N_7716,N_6908,N_6230);
xor U7717 (N_7717,N_6064,N_6501);
nor U7718 (N_7718,N_6782,N_6546);
and U7719 (N_7719,N_6418,N_6856);
and U7720 (N_7720,N_6406,N_6673);
nor U7721 (N_7721,N_6357,N_6840);
or U7722 (N_7722,N_6897,N_6151);
nor U7723 (N_7723,N_6579,N_6701);
nand U7724 (N_7724,N_6308,N_6083);
nand U7725 (N_7725,N_6272,N_6899);
and U7726 (N_7726,N_6356,N_6715);
nand U7727 (N_7727,N_6998,N_6067);
nand U7728 (N_7728,N_6274,N_6923);
nor U7729 (N_7729,N_6505,N_6524);
and U7730 (N_7730,N_6853,N_6677);
xnor U7731 (N_7731,N_6250,N_6643);
xor U7732 (N_7732,N_6711,N_6705);
and U7733 (N_7733,N_6854,N_6176);
and U7734 (N_7734,N_6168,N_6541);
xor U7735 (N_7735,N_6800,N_6320);
and U7736 (N_7736,N_6889,N_6807);
xor U7737 (N_7737,N_6468,N_6178);
nor U7738 (N_7738,N_6949,N_6531);
nor U7739 (N_7739,N_6847,N_6510);
or U7740 (N_7740,N_6302,N_6411);
xor U7741 (N_7741,N_6196,N_6000);
or U7742 (N_7742,N_6051,N_6449);
and U7743 (N_7743,N_6736,N_6136);
and U7744 (N_7744,N_6827,N_6798);
nand U7745 (N_7745,N_6473,N_6319);
xnor U7746 (N_7746,N_6709,N_6877);
and U7747 (N_7747,N_6193,N_6681);
xnor U7748 (N_7748,N_6876,N_6527);
and U7749 (N_7749,N_6885,N_6066);
and U7750 (N_7750,N_6115,N_6540);
nand U7751 (N_7751,N_6590,N_6338);
nor U7752 (N_7752,N_6068,N_6858);
or U7753 (N_7753,N_6214,N_6400);
or U7754 (N_7754,N_6464,N_6148);
or U7755 (N_7755,N_6131,N_6466);
xor U7756 (N_7756,N_6422,N_6602);
nand U7757 (N_7757,N_6291,N_6076);
or U7758 (N_7758,N_6857,N_6184);
xor U7759 (N_7759,N_6800,N_6201);
and U7760 (N_7760,N_6006,N_6141);
or U7761 (N_7761,N_6001,N_6376);
xor U7762 (N_7762,N_6080,N_6319);
xnor U7763 (N_7763,N_6508,N_6043);
or U7764 (N_7764,N_6138,N_6639);
xnor U7765 (N_7765,N_6001,N_6378);
xor U7766 (N_7766,N_6967,N_6972);
and U7767 (N_7767,N_6691,N_6341);
or U7768 (N_7768,N_6889,N_6301);
xnor U7769 (N_7769,N_6662,N_6266);
and U7770 (N_7770,N_6244,N_6138);
nor U7771 (N_7771,N_6710,N_6674);
and U7772 (N_7772,N_6561,N_6054);
xnor U7773 (N_7773,N_6023,N_6971);
nand U7774 (N_7774,N_6501,N_6729);
nand U7775 (N_7775,N_6326,N_6266);
or U7776 (N_7776,N_6792,N_6491);
nand U7777 (N_7777,N_6937,N_6298);
xnor U7778 (N_7778,N_6790,N_6053);
or U7779 (N_7779,N_6162,N_6128);
nand U7780 (N_7780,N_6094,N_6438);
or U7781 (N_7781,N_6634,N_6576);
nand U7782 (N_7782,N_6036,N_6665);
nand U7783 (N_7783,N_6411,N_6234);
or U7784 (N_7784,N_6162,N_6718);
xnor U7785 (N_7785,N_6156,N_6436);
nor U7786 (N_7786,N_6072,N_6546);
or U7787 (N_7787,N_6166,N_6984);
or U7788 (N_7788,N_6636,N_6484);
xor U7789 (N_7789,N_6278,N_6781);
and U7790 (N_7790,N_6721,N_6271);
xor U7791 (N_7791,N_6495,N_6229);
nand U7792 (N_7792,N_6723,N_6859);
nor U7793 (N_7793,N_6225,N_6632);
or U7794 (N_7794,N_6729,N_6080);
xnor U7795 (N_7795,N_6251,N_6897);
and U7796 (N_7796,N_6949,N_6335);
nand U7797 (N_7797,N_6517,N_6016);
or U7798 (N_7798,N_6196,N_6503);
xor U7799 (N_7799,N_6678,N_6946);
nor U7800 (N_7800,N_6794,N_6868);
xnor U7801 (N_7801,N_6451,N_6218);
or U7802 (N_7802,N_6540,N_6027);
or U7803 (N_7803,N_6586,N_6600);
and U7804 (N_7804,N_6886,N_6381);
or U7805 (N_7805,N_6595,N_6112);
xnor U7806 (N_7806,N_6018,N_6771);
xor U7807 (N_7807,N_6001,N_6557);
or U7808 (N_7808,N_6559,N_6557);
nor U7809 (N_7809,N_6289,N_6335);
or U7810 (N_7810,N_6979,N_6815);
or U7811 (N_7811,N_6196,N_6357);
nand U7812 (N_7812,N_6274,N_6623);
and U7813 (N_7813,N_6534,N_6961);
or U7814 (N_7814,N_6334,N_6898);
nand U7815 (N_7815,N_6970,N_6193);
or U7816 (N_7816,N_6650,N_6494);
nor U7817 (N_7817,N_6615,N_6742);
nor U7818 (N_7818,N_6584,N_6598);
xnor U7819 (N_7819,N_6373,N_6886);
nor U7820 (N_7820,N_6584,N_6990);
nand U7821 (N_7821,N_6951,N_6819);
and U7822 (N_7822,N_6184,N_6807);
nor U7823 (N_7823,N_6406,N_6923);
nand U7824 (N_7824,N_6067,N_6387);
or U7825 (N_7825,N_6765,N_6945);
nor U7826 (N_7826,N_6524,N_6420);
nand U7827 (N_7827,N_6833,N_6791);
or U7828 (N_7828,N_6701,N_6201);
nor U7829 (N_7829,N_6491,N_6888);
or U7830 (N_7830,N_6505,N_6843);
and U7831 (N_7831,N_6933,N_6500);
nor U7832 (N_7832,N_6250,N_6867);
nor U7833 (N_7833,N_6180,N_6388);
nor U7834 (N_7834,N_6496,N_6349);
nand U7835 (N_7835,N_6012,N_6258);
nor U7836 (N_7836,N_6123,N_6969);
nand U7837 (N_7837,N_6939,N_6093);
nand U7838 (N_7838,N_6014,N_6533);
nor U7839 (N_7839,N_6407,N_6495);
and U7840 (N_7840,N_6683,N_6215);
nor U7841 (N_7841,N_6690,N_6438);
and U7842 (N_7842,N_6631,N_6127);
xnor U7843 (N_7843,N_6435,N_6650);
nand U7844 (N_7844,N_6435,N_6908);
nor U7845 (N_7845,N_6709,N_6069);
xnor U7846 (N_7846,N_6219,N_6233);
nor U7847 (N_7847,N_6194,N_6420);
nand U7848 (N_7848,N_6896,N_6236);
xor U7849 (N_7849,N_6923,N_6424);
nand U7850 (N_7850,N_6571,N_6529);
xor U7851 (N_7851,N_6505,N_6992);
nor U7852 (N_7852,N_6364,N_6287);
or U7853 (N_7853,N_6637,N_6351);
and U7854 (N_7854,N_6198,N_6729);
nor U7855 (N_7855,N_6872,N_6097);
nor U7856 (N_7856,N_6469,N_6746);
or U7857 (N_7857,N_6231,N_6826);
or U7858 (N_7858,N_6129,N_6682);
or U7859 (N_7859,N_6512,N_6706);
xnor U7860 (N_7860,N_6903,N_6972);
and U7861 (N_7861,N_6466,N_6757);
or U7862 (N_7862,N_6011,N_6621);
nor U7863 (N_7863,N_6260,N_6773);
or U7864 (N_7864,N_6177,N_6661);
xor U7865 (N_7865,N_6870,N_6646);
nand U7866 (N_7866,N_6909,N_6022);
xnor U7867 (N_7867,N_6706,N_6639);
nand U7868 (N_7868,N_6287,N_6826);
or U7869 (N_7869,N_6395,N_6160);
or U7870 (N_7870,N_6819,N_6376);
xor U7871 (N_7871,N_6160,N_6852);
and U7872 (N_7872,N_6213,N_6373);
nor U7873 (N_7873,N_6833,N_6577);
or U7874 (N_7874,N_6477,N_6909);
nand U7875 (N_7875,N_6280,N_6117);
nand U7876 (N_7876,N_6927,N_6144);
or U7877 (N_7877,N_6733,N_6363);
or U7878 (N_7878,N_6877,N_6489);
or U7879 (N_7879,N_6249,N_6163);
xor U7880 (N_7880,N_6972,N_6926);
and U7881 (N_7881,N_6472,N_6629);
nand U7882 (N_7882,N_6273,N_6710);
xor U7883 (N_7883,N_6028,N_6464);
nor U7884 (N_7884,N_6072,N_6037);
nor U7885 (N_7885,N_6905,N_6522);
or U7886 (N_7886,N_6552,N_6522);
and U7887 (N_7887,N_6004,N_6247);
nand U7888 (N_7888,N_6650,N_6353);
or U7889 (N_7889,N_6787,N_6434);
xor U7890 (N_7890,N_6517,N_6046);
xor U7891 (N_7891,N_6360,N_6656);
nand U7892 (N_7892,N_6407,N_6602);
or U7893 (N_7893,N_6466,N_6849);
xnor U7894 (N_7894,N_6876,N_6283);
or U7895 (N_7895,N_6126,N_6339);
xor U7896 (N_7896,N_6373,N_6957);
nand U7897 (N_7897,N_6414,N_6447);
nand U7898 (N_7898,N_6831,N_6911);
and U7899 (N_7899,N_6667,N_6578);
nand U7900 (N_7900,N_6809,N_6763);
xor U7901 (N_7901,N_6140,N_6351);
nand U7902 (N_7902,N_6090,N_6166);
and U7903 (N_7903,N_6786,N_6002);
nor U7904 (N_7904,N_6460,N_6792);
nand U7905 (N_7905,N_6476,N_6716);
xor U7906 (N_7906,N_6613,N_6336);
nor U7907 (N_7907,N_6087,N_6743);
or U7908 (N_7908,N_6022,N_6502);
and U7909 (N_7909,N_6015,N_6164);
and U7910 (N_7910,N_6010,N_6857);
xnor U7911 (N_7911,N_6864,N_6071);
nand U7912 (N_7912,N_6073,N_6872);
or U7913 (N_7913,N_6977,N_6304);
nand U7914 (N_7914,N_6823,N_6073);
xnor U7915 (N_7915,N_6396,N_6765);
xnor U7916 (N_7916,N_6665,N_6317);
nand U7917 (N_7917,N_6258,N_6482);
nand U7918 (N_7918,N_6278,N_6832);
xor U7919 (N_7919,N_6051,N_6899);
or U7920 (N_7920,N_6764,N_6791);
and U7921 (N_7921,N_6880,N_6515);
and U7922 (N_7922,N_6885,N_6255);
nand U7923 (N_7923,N_6530,N_6000);
or U7924 (N_7924,N_6340,N_6147);
nor U7925 (N_7925,N_6301,N_6870);
nor U7926 (N_7926,N_6633,N_6100);
xor U7927 (N_7927,N_6186,N_6296);
nand U7928 (N_7928,N_6476,N_6408);
xor U7929 (N_7929,N_6778,N_6607);
or U7930 (N_7930,N_6995,N_6680);
nor U7931 (N_7931,N_6047,N_6450);
nor U7932 (N_7932,N_6926,N_6401);
nor U7933 (N_7933,N_6044,N_6382);
or U7934 (N_7934,N_6067,N_6485);
and U7935 (N_7935,N_6306,N_6189);
and U7936 (N_7936,N_6271,N_6354);
and U7937 (N_7937,N_6690,N_6726);
nor U7938 (N_7938,N_6143,N_6130);
nand U7939 (N_7939,N_6467,N_6348);
nor U7940 (N_7940,N_6700,N_6424);
or U7941 (N_7941,N_6786,N_6696);
xnor U7942 (N_7942,N_6781,N_6213);
or U7943 (N_7943,N_6498,N_6801);
nand U7944 (N_7944,N_6166,N_6913);
xor U7945 (N_7945,N_6082,N_6752);
or U7946 (N_7946,N_6161,N_6624);
nand U7947 (N_7947,N_6163,N_6547);
xnor U7948 (N_7948,N_6388,N_6100);
or U7949 (N_7949,N_6907,N_6089);
nor U7950 (N_7950,N_6489,N_6345);
xor U7951 (N_7951,N_6362,N_6335);
xor U7952 (N_7952,N_6224,N_6219);
nor U7953 (N_7953,N_6529,N_6330);
and U7954 (N_7954,N_6606,N_6743);
xor U7955 (N_7955,N_6411,N_6836);
or U7956 (N_7956,N_6076,N_6126);
and U7957 (N_7957,N_6362,N_6624);
nor U7958 (N_7958,N_6774,N_6534);
nor U7959 (N_7959,N_6414,N_6058);
or U7960 (N_7960,N_6439,N_6826);
nand U7961 (N_7961,N_6478,N_6151);
nor U7962 (N_7962,N_6860,N_6083);
nand U7963 (N_7963,N_6778,N_6722);
or U7964 (N_7964,N_6805,N_6901);
or U7965 (N_7965,N_6206,N_6761);
nand U7966 (N_7966,N_6629,N_6367);
nor U7967 (N_7967,N_6989,N_6816);
or U7968 (N_7968,N_6137,N_6464);
nand U7969 (N_7969,N_6602,N_6188);
nor U7970 (N_7970,N_6698,N_6288);
xnor U7971 (N_7971,N_6216,N_6708);
xnor U7972 (N_7972,N_6259,N_6521);
nor U7973 (N_7973,N_6981,N_6791);
and U7974 (N_7974,N_6337,N_6946);
nor U7975 (N_7975,N_6776,N_6995);
nand U7976 (N_7976,N_6582,N_6398);
xnor U7977 (N_7977,N_6807,N_6428);
and U7978 (N_7978,N_6209,N_6017);
nand U7979 (N_7979,N_6211,N_6784);
nor U7980 (N_7980,N_6665,N_6457);
nand U7981 (N_7981,N_6943,N_6164);
xor U7982 (N_7982,N_6945,N_6801);
xnor U7983 (N_7983,N_6159,N_6193);
xnor U7984 (N_7984,N_6751,N_6582);
nor U7985 (N_7985,N_6121,N_6799);
nand U7986 (N_7986,N_6337,N_6399);
and U7987 (N_7987,N_6565,N_6477);
and U7988 (N_7988,N_6190,N_6322);
nand U7989 (N_7989,N_6389,N_6550);
nand U7990 (N_7990,N_6422,N_6956);
and U7991 (N_7991,N_6362,N_6880);
nor U7992 (N_7992,N_6565,N_6420);
or U7993 (N_7993,N_6624,N_6108);
nand U7994 (N_7994,N_6325,N_6285);
nand U7995 (N_7995,N_6918,N_6810);
nand U7996 (N_7996,N_6063,N_6996);
and U7997 (N_7997,N_6606,N_6280);
nand U7998 (N_7998,N_6217,N_6987);
xor U7999 (N_7999,N_6456,N_6484);
nor U8000 (N_8000,N_7885,N_7715);
and U8001 (N_8001,N_7433,N_7208);
or U8002 (N_8002,N_7414,N_7207);
or U8003 (N_8003,N_7301,N_7920);
nor U8004 (N_8004,N_7965,N_7701);
nand U8005 (N_8005,N_7387,N_7108);
nor U8006 (N_8006,N_7296,N_7825);
xnor U8007 (N_8007,N_7032,N_7751);
and U8008 (N_8008,N_7412,N_7114);
nand U8009 (N_8009,N_7709,N_7667);
xor U8010 (N_8010,N_7502,N_7256);
xnor U8011 (N_8011,N_7326,N_7214);
and U8012 (N_8012,N_7453,N_7764);
nor U8013 (N_8013,N_7640,N_7641);
and U8014 (N_8014,N_7394,N_7507);
xnor U8015 (N_8015,N_7887,N_7959);
nor U8016 (N_8016,N_7355,N_7639);
nand U8017 (N_8017,N_7204,N_7197);
nor U8018 (N_8018,N_7698,N_7379);
or U8019 (N_8019,N_7949,N_7606);
xnor U8020 (N_8020,N_7378,N_7155);
nand U8021 (N_8021,N_7141,N_7727);
nor U8022 (N_8022,N_7780,N_7110);
or U8023 (N_8023,N_7788,N_7921);
and U8024 (N_8024,N_7358,N_7315);
and U8025 (N_8025,N_7448,N_7418);
nand U8026 (N_8026,N_7305,N_7392);
nor U8027 (N_8027,N_7483,N_7468);
nand U8028 (N_8028,N_7530,N_7730);
or U8029 (N_8029,N_7390,N_7362);
nand U8030 (N_8030,N_7031,N_7400);
nor U8031 (N_8031,N_7829,N_7045);
xor U8032 (N_8032,N_7983,N_7666);
xnor U8033 (N_8033,N_7842,N_7810);
nor U8034 (N_8034,N_7516,N_7515);
and U8035 (N_8035,N_7747,N_7773);
or U8036 (N_8036,N_7374,N_7377);
and U8037 (N_8037,N_7619,N_7932);
nand U8038 (N_8038,N_7153,N_7271);
nand U8039 (N_8039,N_7977,N_7323);
nor U8040 (N_8040,N_7503,N_7867);
or U8041 (N_8041,N_7524,N_7465);
or U8042 (N_8042,N_7156,N_7350);
and U8043 (N_8043,N_7955,N_7783);
xnor U8044 (N_8044,N_7703,N_7725);
or U8045 (N_8045,N_7984,N_7405);
nand U8046 (N_8046,N_7539,N_7324);
xnor U8047 (N_8047,N_7275,N_7840);
or U8048 (N_8048,N_7099,N_7508);
nor U8049 (N_8049,N_7929,N_7707);
nor U8050 (N_8050,N_7196,N_7924);
or U8051 (N_8051,N_7257,N_7230);
and U8052 (N_8052,N_7423,N_7716);
nor U8053 (N_8053,N_7091,N_7813);
and U8054 (N_8054,N_7556,N_7946);
xor U8055 (N_8055,N_7778,N_7149);
and U8056 (N_8056,N_7118,N_7664);
nand U8057 (N_8057,N_7314,N_7564);
nor U8058 (N_8058,N_7679,N_7452);
nand U8059 (N_8059,N_7368,N_7280);
or U8060 (N_8060,N_7660,N_7767);
nor U8061 (N_8061,N_7759,N_7522);
and U8062 (N_8062,N_7923,N_7426);
and U8063 (N_8063,N_7194,N_7389);
nor U8064 (N_8064,N_7839,N_7056);
xor U8065 (N_8065,N_7163,N_7854);
xor U8066 (N_8066,N_7001,N_7501);
nand U8067 (N_8067,N_7478,N_7025);
or U8068 (N_8068,N_7222,N_7677);
nand U8069 (N_8069,N_7816,N_7781);
nor U8070 (N_8070,N_7688,N_7255);
nand U8071 (N_8071,N_7450,N_7051);
xor U8072 (N_8072,N_7057,N_7279);
nand U8073 (N_8073,N_7420,N_7457);
or U8074 (N_8074,N_7048,N_7859);
or U8075 (N_8075,N_7933,N_7916);
nor U8076 (N_8076,N_7500,N_7439);
xor U8077 (N_8077,N_7819,N_7321);
nor U8078 (N_8078,N_7975,N_7003);
xnor U8079 (N_8079,N_7901,N_7239);
nand U8080 (N_8080,N_7444,N_7659);
nand U8081 (N_8081,N_7541,N_7283);
nand U8082 (N_8082,N_7080,N_7729);
and U8083 (N_8083,N_7352,N_7934);
nand U8084 (N_8084,N_7732,N_7513);
or U8085 (N_8085,N_7310,N_7528);
and U8086 (N_8086,N_7891,N_7008);
xnor U8087 (N_8087,N_7202,N_7333);
nor U8088 (N_8088,N_7168,N_7044);
nor U8089 (N_8089,N_7122,N_7771);
and U8090 (N_8090,N_7436,N_7154);
nor U8091 (N_8091,N_7160,N_7776);
or U8092 (N_8092,N_7259,N_7079);
nor U8093 (N_8093,N_7179,N_7769);
or U8094 (N_8094,N_7061,N_7096);
xor U8095 (N_8095,N_7325,N_7753);
xnor U8096 (N_8096,N_7422,N_7894);
and U8097 (N_8097,N_7415,N_7672);
or U8098 (N_8098,N_7888,N_7630);
nor U8099 (N_8099,N_7177,N_7908);
xnor U8100 (N_8100,N_7713,N_7724);
and U8101 (N_8101,N_7629,N_7049);
or U8102 (N_8102,N_7437,N_7055);
nand U8103 (N_8103,N_7237,N_7077);
nand U8104 (N_8104,N_7095,N_7477);
nand U8105 (N_8105,N_7957,N_7951);
and U8106 (N_8106,N_7600,N_7135);
xnor U8107 (N_8107,N_7058,N_7624);
and U8108 (N_8108,N_7419,N_7429);
xor U8109 (N_8109,N_7559,N_7602);
xnor U8110 (N_8110,N_7488,N_7900);
nor U8111 (N_8111,N_7388,N_7763);
nor U8112 (N_8112,N_7313,N_7073);
nand U8113 (N_8113,N_7584,N_7183);
nor U8114 (N_8114,N_7798,N_7789);
or U8115 (N_8115,N_7143,N_7626);
nor U8116 (N_8116,N_7219,N_7342);
nor U8117 (N_8117,N_7004,N_7790);
xnor U8118 (N_8118,N_7245,N_7066);
nand U8119 (N_8119,N_7112,N_7162);
and U8120 (N_8120,N_7517,N_7953);
nor U8121 (N_8121,N_7235,N_7650);
nor U8122 (N_8122,N_7950,N_7131);
or U8123 (N_8123,N_7871,N_7070);
nor U8124 (N_8124,N_7801,N_7735);
or U8125 (N_8125,N_7292,N_7944);
nor U8126 (N_8126,N_7111,N_7647);
xor U8127 (N_8127,N_7895,N_7940);
xor U8128 (N_8128,N_7519,N_7613);
and U8129 (N_8129,N_7571,N_7100);
nand U8130 (N_8130,N_7968,N_7527);
or U8131 (N_8131,N_7126,N_7481);
or U8132 (N_8132,N_7775,N_7307);
and U8133 (N_8133,N_7892,N_7733);
xor U8134 (N_8134,N_7897,N_7808);
nor U8135 (N_8135,N_7213,N_7147);
nor U8136 (N_8136,N_7329,N_7845);
nor U8137 (N_8137,N_7399,N_7708);
or U8138 (N_8138,N_7263,N_7142);
xor U8139 (N_8139,N_7391,N_7912);
and U8140 (N_8140,N_7546,N_7364);
xor U8141 (N_8141,N_7037,N_7124);
or U8142 (N_8142,N_7806,N_7942);
or U8143 (N_8143,N_7490,N_7140);
nand U8144 (N_8144,N_7148,N_7996);
or U8145 (N_8145,N_7286,N_7473);
or U8146 (N_8146,N_7447,N_7675);
nor U8147 (N_8147,N_7351,N_7869);
and U8148 (N_8148,N_7749,N_7532);
nand U8149 (N_8149,N_7739,N_7621);
nor U8150 (N_8150,N_7841,N_7172);
nand U8151 (N_8151,N_7756,N_7475);
nor U8152 (N_8152,N_7435,N_7247);
and U8153 (N_8153,N_7910,N_7631);
nand U8154 (N_8154,N_7171,N_7694);
and U8155 (N_8155,N_7898,N_7252);
or U8156 (N_8156,N_7879,N_7896);
or U8157 (N_8157,N_7234,N_7565);
nand U8158 (N_8158,N_7577,N_7434);
nand U8159 (N_8159,N_7590,N_7697);
nor U8160 (N_8160,N_7406,N_7480);
and U8161 (N_8161,N_7890,N_7521);
or U8162 (N_8162,N_7087,N_7467);
nand U8163 (N_8163,N_7381,N_7159);
nand U8164 (N_8164,N_7327,N_7088);
nand U8165 (N_8165,N_7092,N_7121);
xnor U8166 (N_8166,N_7766,N_7462);
nor U8167 (N_8167,N_7760,N_7711);
nand U8168 (N_8168,N_7486,N_7529);
or U8169 (N_8169,N_7979,N_7623);
nand U8170 (N_8170,N_7016,N_7236);
nand U8171 (N_8171,N_7262,N_7687);
or U8172 (N_8172,N_7880,N_7047);
nor U8173 (N_8173,N_7007,N_7410);
and U8174 (N_8174,N_7827,N_7791);
xor U8175 (N_8175,N_7928,N_7385);
and U8176 (N_8176,N_7525,N_7714);
xnor U8177 (N_8177,N_7846,N_7877);
xor U8178 (N_8178,N_7855,N_7557);
xnor U8179 (N_8179,N_7233,N_7992);
nand U8180 (N_8180,N_7874,N_7266);
xor U8181 (N_8181,N_7015,N_7134);
or U8182 (N_8182,N_7925,N_7312);
nor U8183 (N_8183,N_7914,N_7611);
or U8184 (N_8184,N_7591,N_7568);
nand U8185 (N_8185,N_7241,N_7669);
xnor U8186 (N_8186,N_7268,N_7186);
nor U8187 (N_8187,N_7570,N_7344);
nor U8188 (N_8188,N_7978,N_7594);
or U8189 (N_8189,N_7881,N_7402);
nor U8190 (N_8190,N_7030,N_7821);
or U8191 (N_8191,N_7216,N_7913);
and U8192 (N_8192,N_7098,N_7768);
xor U8193 (N_8193,N_7603,N_7548);
or U8194 (N_8194,N_7523,N_7856);
xor U8195 (N_8195,N_7661,N_7620);
nand U8196 (N_8196,N_7765,N_7097);
and U8197 (N_8197,N_7017,N_7461);
and U8198 (N_8198,N_7440,N_7123);
xnor U8199 (N_8199,N_7248,N_7253);
nand U8200 (N_8200,N_7982,N_7549);
nand U8201 (N_8201,N_7199,N_7614);
nor U8202 (N_8202,N_7165,N_7533);
nor U8203 (N_8203,N_7864,N_7947);
or U8204 (N_8204,N_7618,N_7662);
nand U8205 (N_8205,N_7023,N_7634);
or U8206 (N_8206,N_7592,N_7962);
xor U8207 (N_8207,N_7225,N_7157);
nand U8208 (N_8208,N_7849,N_7930);
and U8209 (N_8209,N_7474,N_7460);
xnor U8210 (N_8210,N_7282,N_7258);
xnor U8211 (N_8211,N_7671,N_7628);
or U8212 (N_8212,N_7065,N_7361);
nand U8213 (N_8213,N_7341,N_7396);
or U8214 (N_8214,N_7064,N_7411);
xor U8215 (N_8215,N_7884,N_7021);
xnor U8216 (N_8216,N_7089,N_7700);
and U8217 (N_8217,N_7745,N_7356);
xor U8218 (N_8218,N_7642,N_7260);
nand U8219 (N_8219,N_7941,N_7328);
and U8220 (N_8220,N_7685,N_7693);
or U8221 (N_8221,N_7824,N_7334);
nand U8222 (N_8222,N_7487,N_7288);
nand U8223 (N_8223,N_7779,N_7425);
xnor U8224 (N_8224,N_7536,N_7980);
nor U8225 (N_8225,N_7710,N_7298);
and U8226 (N_8226,N_7303,N_7802);
nand U8227 (N_8227,N_7878,N_7543);
or U8228 (N_8228,N_7853,N_7970);
nand U8229 (N_8229,N_7935,N_7598);
xnor U8230 (N_8230,N_7084,N_7404);
and U8231 (N_8231,N_7883,N_7408);
nor U8232 (N_8232,N_7649,N_7251);
nand U8233 (N_8233,N_7309,N_7917);
nor U8234 (N_8234,N_7013,N_7445);
nand U8235 (N_8235,N_7876,N_7347);
nor U8236 (N_8236,N_7482,N_7318);
and U8237 (N_8237,N_7206,N_7063);
nor U8238 (N_8238,N_7865,N_7109);
xor U8239 (N_8239,N_7033,N_7812);
or U8240 (N_8240,N_7012,N_7043);
or U8241 (N_8241,N_7862,N_7269);
nor U8242 (N_8242,N_7542,N_7998);
and U8243 (N_8243,N_7873,N_7201);
and U8244 (N_8244,N_7428,N_7952);
nand U8245 (N_8245,N_7755,N_7691);
or U8246 (N_8246,N_7062,N_7299);
or U8247 (N_8247,N_7971,N_7441);
xor U8248 (N_8248,N_7526,N_7999);
xor U8249 (N_8249,N_7491,N_7985);
nand U8250 (N_8250,N_7608,N_7981);
and U8251 (N_8251,N_7615,N_7178);
nor U8252 (N_8252,N_7116,N_7136);
nand U8253 (N_8253,N_7242,N_7376);
or U8254 (N_8254,N_7866,N_7297);
and U8255 (N_8255,N_7627,N_7102);
and U8256 (N_8256,N_7586,N_7692);
xor U8257 (N_8257,N_7676,N_7146);
or U8258 (N_8258,N_7567,N_7550);
nor U8259 (N_8259,N_7416,N_7169);
nor U8260 (N_8260,N_7834,N_7553);
nand U8261 (N_8261,N_7072,N_7616);
xor U8262 (N_8262,N_7345,N_7195);
or U8263 (N_8263,N_7674,N_7238);
nor U8264 (N_8264,N_7939,N_7181);
and U8265 (N_8265,N_7758,N_7218);
nand U8266 (N_8266,N_7024,N_7188);
or U8267 (N_8267,N_7166,N_7086);
and U8268 (N_8268,N_7814,N_7720);
nand U8269 (N_8269,N_7330,N_7050);
or U8270 (N_8270,N_7499,N_7074);
nand U8271 (N_8271,N_7451,N_7212);
nor U8272 (N_8272,N_7994,N_7466);
or U8273 (N_8273,N_7265,N_7651);
xnor U8274 (N_8274,N_7200,N_7987);
xnor U8275 (N_8275,N_7117,N_7316);
nor U8276 (N_8276,N_7370,N_7289);
and U8277 (N_8277,N_7384,N_7961);
nand U8278 (N_8278,N_7078,N_7607);
and U8279 (N_8279,N_7903,N_7860);
nor U8280 (N_8280,N_7966,N_7656);
xnor U8281 (N_8281,N_7844,N_7706);
nor U8282 (N_8282,N_7906,N_7636);
or U8283 (N_8283,N_7909,N_7511);
or U8284 (N_8284,N_7250,N_7489);
or U8285 (N_8285,N_7028,N_7438);
and U8286 (N_8286,N_7005,N_7907);
and U8287 (N_8287,N_7538,N_7742);
xor U8288 (N_8288,N_7902,N_7340);
nand U8289 (N_8289,N_7609,N_7723);
or U8290 (N_8290,N_7772,N_7161);
or U8291 (N_8291,N_7432,N_7833);
nand U8292 (N_8292,N_7354,N_7743);
and U8293 (N_8293,N_7974,N_7366);
nand U8294 (N_8294,N_7915,N_7454);
or U8295 (N_8295,N_7803,N_7304);
xnor U8296 (N_8296,N_7809,N_7203);
xnor U8297 (N_8297,N_7562,N_7799);
or U8298 (N_8298,N_7848,N_7637);
or U8299 (N_8299,N_7800,N_7128);
and U8300 (N_8300,N_7997,N_7823);
or U8301 (N_8301,N_7311,N_7964);
and U8302 (N_8302,N_7872,N_7430);
or U8303 (N_8303,N_7040,N_7363);
nor U8304 (N_8304,N_7119,N_7645);
nand U8305 (N_8305,N_7011,N_7596);
and U8306 (N_8306,N_7835,N_7815);
nand U8307 (N_8307,N_7287,N_7520);
and U8308 (N_8308,N_7223,N_7851);
xnor U8309 (N_8309,N_7176,N_7284);
nand U8310 (N_8310,N_7270,N_7699);
or U8311 (N_8311,N_7371,N_7741);
xnor U8312 (N_8312,N_7215,N_7217);
and U8313 (N_8313,N_7658,N_7348);
or U8314 (N_8314,N_7331,N_7882);
nor U8315 (N_8315,N_7459,N_7372);
nand U8316 (N_8316,N_7817,N_7076);
nor U8317 (N_8317,N_7278,N_7495);
and U8318 (N_8318,N_7211,N_7173);
nand U8319 (N_8319,N_7139,N_7332);
xnor U8320 (N_8320,N_7456,N_7837);
or U8321 (N_8321,N_7752,N_7512);
and U8322 (N_8322,N_7943,N_7967);
nand U8323 (N_8323,N_7681,N_7187);
and U8324 (N_8324,N_7684,N_7736);
and U8325 (N_8325,N_7811,N_7551);
xor U8326 (N_8326,N_7795,N_7035);
xnor U8327 (N_8327,N_7680,N_7617);
and U8328 (N_8328,N_7805,N_7740);
or U8329 (N_8329,N_7053,N_7471);
xnor U8330 (N_8330,N_7663,N_7861);
nand U8331 (N_8331,N_7132,N_7518);
nand U8332 (N_8332,N_7514,N_7638);
nand U8333 (N_8333,N_7382,N_7277);
xor U8334 (N_8334,N_7373,N_7020);
nand U8335 (N_8335,N_7113,N_7285);
nand U8336 (N_8336,N_7427,N_7145);
nor U8337 (N_8337,N_7678,N_7104);
xnor U8338 (N_8338,N_7101,N_7386);
and U8339 (N_8339,N_7583,N_7317);
xnor U8340 (N_8340,N_7417,N_7643);
xor U8341 (N_8341,N_7726,N_7174);
or U8342 (N_8342,N_7682,N_7375);
xor U8343 (N_8343,N_7774,N_7308);
or U8344 (N_8344,N_7744,N_7130);
or U8345 (N_8345,N_7762,N_7972);
nor U8346 (N_8346,N_7221,N_7424);
and U8347 (N_8347,N_7610,N_7272);
nor U8348 (N_8348,N_7039,N_7449);
xor U8349 (N_8349,N_7267,N_7654);
xnor U8350 (N_8350,N_7818,N_7127);
nor U8351 (N_8351,N_7357,N_7353);
and U8352 (N_8352,N_7976,N_7261);
or U8353 (N_8353,N_7988,N_7464);
nand U8354 (N_8354,N_7785,N_7938);
or U8355 (N_8355,N_7446,N_7041);
nor U8356 (N_8356,N_7734,N_7249);
nand U8357 (N_8357,N_7995,N_7403);
nor U8358 (N_8358,N_7504,N_7338);
or U8359 (N_8359,N_7232,N_7843);
nand U8360 (N_8360,N_7264,N_7797);
or U8361 (N_8361,N_7455,N_7281);
nand U8362 (N_8362,N_7973,N_7652);
nor U8363 (N_8363,N_7863,N_7210);
xor U8364 (N_8364,N_7018,N_7068);
xor U8365 (N_8365,N_7137,N_7254);
xor U8366 (N_8366,N_7822,N_7632);
nand U8367 (N_8367,N_7804,N_7576);
and U8368 (N_8368,N_7198,N_7721);
nand U8369 (N_8369,N_7274,N_7306);
xor U8370 (N_8370,N_7657,N_7034);
and U8371 (N_8371,N_7138,N_7052);
nand U8372 (N_8372,N_7850,N_7991);
or U8373 (N_8373,N_7604,N_7605);
and U8374 (N_8374,N_7106,N_7082);
nor U8375 (N_8375,N_7151,N_7227);
or U8376 (N_8376,N_7534,N_7060);
nand U8377 (N_8377,N_7580,N_7494);
nand U8378 (N_8378,N_7026,N_7537);
nor U8379 (N_8379,N_7493,N_7209);
or U8380 (N_8380,N_7722,N_7847);
nor U8381 (N_8381,N_7807,N_7831);
nand U8382 (N_8382,N_7936,N_7367);
nor U8383 (N_8383,N_7746,N_7343);
xnor U8384 (N_8384,N_7226,N_7793);
or U8385 (N_8385,N_7828,N_7717);
nand U8386 (N_8386,N_7931,N_7360);
xor U8387 (N_8387,N_7963,N_7545);
and U8388 (N_8388,N_7830,N_7622);
nor U8389 (N_8389,N_7597,N_7273);
xor U8390 (N_8390,N_7555,N_7094);
or U8391 (N_8391,N_7046,N_7969);
nor U8392 (N_8392,N_7653,N_7852);
or U8393 (N_8393,N_7673,N_7359);
nand U8394 (N_8394,N_7000,N_7152);
xor U8395 (N_8395,N_7335,N_7820);
nor U8396 (N_8396,N_7421,N_7191);
and U8397 (N_8397,N_7686,N_7566);
nand U8398 (N_8398,N_7059,N_7719);
nand U8399 (N_8399,N_7190,N_7506);
nand U8400 (N_8400,N_7893,N_7244);
nand U8401 (N_8401,N_7192,N_7067);
and U8402 (N_8402,N_7240,N_7081);
nand U8403 (N_8403,N_7886,N_7243);
xor U8404 (N_8404,N_7458,N_7105);
or U8405 (N_8405,N_7705,N_7397);
and U8406 (N_8406,N_7593,N_7349);
nand U8407 (N_8407,N_7993,N_7167);
nand U8408 (N_8408,N_7069,N_7540);
or U8409 (N_8409,N_7071,N_7737);
nand U8410 (N_8410,N_7761,N_7569);
or U8411 (N_8411,N_7150,N_7784);
or U8412 (N_8412,N_7728,N_7409);
xor U8413 (N_8413,N_7782,N_7958);
or U8414 (N_8414,N_7560,N_7588);
or U8415 (N_8415,N_7125,N_7413);
xnor U8416 (N_8416,N_7479,N_7683);
and U8417 (N_8417,N_7291,N_7754);
and U8418 (N_8418,N_7510,N_7010);
and U8419 (N_8419,N_7498,N_7919);
nand U8420 (N_8420,N_7144,N_7575);
nor U8421 (N_8421,N_7319,N_7470);
xnor U8422 (N_8422,N_7103,N_7295);
nor U8423 (N_8423,N_7009,N_7646);
nand U8424 (N_8424,N_7612,N_7574);
nor U8425 (N_8425,N_7369,N_7904);
nand U8426 (N_8426,N_7184,N_7561);
and U8427 (N_8427,N_7294,N_7563);
nor U8428 (N_8428,N_7246,N_7648);
xor U8429 (N_8429,N_7476,N_7029);
and U8430 (N_8430,N_7712,N_7189);
or U8431 (N_8431,N_7702,N_7276);
or U8432 (N_8432,N_7164,N_7670);
or U8433 (N_8433,N_7175,N_7365);
and U8434 (N_8434,N_7937,N_7180);
nand U8435 (N_8435,N_7485,N_7129);
or U8436 (N_8436,N_7085,N_7731);
or U8437 (N_8437,N_7042,N_7558);
or U8438 (N_8438,N_7182,N_7075);
nor U8439 (N_8439,N_7229,N_7472);
xor U8440 (N_8440,N_7220,N_7302);
xor U8441 (N_8441,N_7552,N_7133);
nand U8442 (N_8442,N_7492,N_7038);
nor U8443 (N_8443,N_7792,N_7770);
nor U8444 (N_8444,N_7544,N_7115);
xnor U8445 (N_8445,N_7750,N_7554);
and U8446 (N_8446,N_7442,N_7228);
nor U8447 (N_8447,N_7899,N_7870);
nor U8448 (N_8448,N_7339,N_7836);
xor U8449 (N_8449,N_7393,N_7911);
or U8450 (N_8450,N_7858,N_7573);
nor U8451 (N_8451,N_7625,N_7158);
or U8452 (N_8452,N_7786,N_7838);
nor U8453 (N_8453,N_7601,N_7585);
nand U8454 (N_8454,N_7547,N_7579);
nand U8455 (N_8455,N_7794,N_7695);
nor U8456 (N_8456,N_7290,N_7589);
xnor U8457 (N_8457,N_7300,N_7395);
nor U8458 (N_8458,N_7905,N_7401);
or U8459 (N_8459,N_7927,N_7572);
nand U8460 (N_8460,N_7535,N_7655);
xnor U8461 (N_8461,N_7696,N_7170);
xnor U8462 (N_8462,N_7704,N_7690);
and U8463 (N_8463,N_7578,N_7926);
xor U8464 (N_8464,N_7531,N_7826);
or U8465 (N_8465,N_7380,N_7107);
nand U8466 (N_8466,N_7582,N_7463);
nand U8467 (N_8467,N_7948,N_7336);
and U8468 (N_8468,N_7889,N_7777);
and U8469 (N_8469,N_7787,N_7185);
nand U8470 (N_8470,N_7120,N_7738);
nor U8471 (N_8471,N_7224,N_7006);
xor U8472 (N_8472,N_7320,N_7644);
or U8473 (N_8473,N_7796,N_7665);
xor U8474 (N_8474,N_7054,N_7002);
nand U8475 (N_8475,N_7014,N_7036);
nand U8476 (N_8476,N_7956,N_7875);
nor U8477 (N_8477,N_7027,N_7718);
and U8478 (N_8478,N_7469,N_7918);
nand U8479 (N_8479,N_7509,N_7497);
nand U8480 (N_8480,N_7322,N_7922);
or U8481 (N_8481,N_7990,N_7868);
xnor U8482 (N_8482,N_7505,N_7398);
and U8483 (N_8483,N_7832,N_7748);
nand U8484 (N_8484,N_7022,N_7083);
nand U8485 (N_8485,N_7986,N_7346);
and U8486 (N_8486,N_7231,N_7757);
nand U8487 (N_8487,N_7587,N_7945);
and U8488 (N_8488,N_7407,N_7205);
xnor U8489 (N_8489,N_7668,N_7383);
nand U8490 (N_8490,N_7431,N_7954);
nand U8491 (N_8491,N_7595,N_7635);
nand U8492 (N_8492,N_7093,N_7293);
nor U8493 (N_8493,N_7960,N_7689);
nor U8494 (N_8494,N_7090,N_7496);
nor U8495 (N_8495,N_7484,N_7581);
nor U8496 (N_8496,N_7443,N_7337);
nand U8497 (N_8497,N_7599,N_7857);
xnor U8498 (N_8498,N_7193,N_7633);
and U8499 (N_8499,N_7989,N_7019);
nand U8500 (N_8500,N_7702,N_7630);
nor U8501 (N_8501,N_7095,N_7130);
xor U8502 (N_8502,N_7795,N_7323);
and U8503 (N_8503,N_7056,N_7112);
or U8504 (N_8504,N_7386,N_7389);
or U8505 (N_8505,N_7990,N_7614);
or U8506 (N_8506,N_7976,N_7932);
and U8507 (N_8507,N_7099,N_7161);
and U8508 (N_8508,N_7494,N_7428);
nand U8509 (N_8509,N_7342,N_7184);
and U8510 (N_8510,N_7867,N_7649);
xor U8511 (N_8511,N_7817,N_7892);
and U8512 (N_8512,N_7597,N_7844);
and U8513 (N_8513,N_7296,N_7835);
xor U8514 (N_8514,N_7577,N_7496);
nand U8515 (N_8515,N_7196,N_7274);
nand U8516 (N_8516,N_7279,N_7326);
xor U8517 (N_8517,N_7136,N_7639);
or U8518 (N_8518,N_7385,N_7087);
or U8519 (N_8519,N_7149,N_7673);
xor U8520 (N_8520,N_7509,N_7411);
or U8521 (N_8521,N_7099,N_7095);
nor U8522 (N_8522,N_7448,N_7288);
nor U8523 (N_8523,N_7020,N_7527);
nor U8524 (N_8524,N_7028,N_7052);
and U8525 (N_8525,N_7368,N_7616);
or U8526 (N_8526,N_7405,N_7409);
nor U8527 (N_8527,N_7278,N_7308);
xor U8528 (N_8528,N_7659,N_7692);
nand U8529 (N_8529,N_7313,N_7647);
nand U8530 (N_8530,N_7690,N_7879);
nand U8531 (N_8531,N_7125,N_7186);
nor U8532 (N_8532,N_7243,N_7708);
or U8533 (N_8533,N_7167,N_7397);
or U8534 (N_8534,N_7037,N_7680);
and U8535 (N_8535,N_7095,N_7472);
or U8536 (N_8536,N_7160,N_7169);
nand U8537 (N_8537,N_7859,N_7588);
or U8538 (N_8538,N_7468,N_7265);
or U8539 (N_8539,N_7321,N_7670);
xnor U8540 (N_8540,N_7377,N_7551);
nor U8541 (N_8541,N_7446,N_7686);
nand U8542 (N_8542,N_7231,N_7002);
or U8543 (N_8543,N_7274,N_7551);
and U8544 (N_8544,N_7585,N_7655);
or U8545 (N_8545,N_7955,N_7662);
nand U8546 (N_8546,N_7857,N_7156);
nor U8547 (N_8547,N_7843,N_7447);
nor U8548 (N_8548,N_7299,N_7889);
nor U8549 (N_8549,N_7075,N_7900);
or U8550 (N_8550,N_7239,N_7104);
and U8551 (N_8551,N_7045,N_7055);
or U8552 (N_8552,N_7732,N_7997);
xor U8553 (N_8553,N_7981,N_7116);
or U8554 (N_8554,N_7437,N_7376);
and U8555 (N_8555,N_7453,N_7611);
nor U8556 (N_8556,N_7658,N_7061);
nand U8557 (N_8557,N_7397,N_7164);
xnor U8558 (N_8558,N_7025,N_7811);
and U8559 (N_8559,N_7145,N_7232);
xnor U8560 (N_8560,N_7980,N_7732);
nand U8561 (N_8561,N_7822,N_7407);
or U8562 (N_8562,N_7842,N_7290);
xnor U8563 (N_8563,N_7081,N_7912);
xnor U8564 (N_8564,N_7195,N_7538);
and U8565 (N_8565,N_7950,N_7166);
nor U8566 (N_8566,N_7646,N_7605);
nor U8567 (N_8567,N_7488,N_7679);
xor U8568 (N_8568,N_7438,N_7607);
nand U8569 (N_8569,N_7318,N_7249);
or U8570 (N_8570,N_7351,N_7064);
xor U8571 (N_8571,N_7757,N_7764);
nand U8572 (N_8572,N_7689,N_7623);
and U8573 (N_8573,N_7014,N_7483);
or U8574 (N_8574,N_7782,N_7983);
xor U8575 (N_8575,N_7896,N_7379);
nand U8576 (N_8576,N_7028,N_7037);
or U8577 (N_8577,N_7761,N_7229);
or U8578 (N_8578,N_7792,N_7027);
or U8579 (N_8579,N_7553,N_7089);
nand U8580 (N_8580,N_7271,N_7553);
and U8581 (N_8581,N_7969,N_7442);
xnor U8582 (N_8582,N_7868,N_7187);
or U8583 (N_8583,N_7978,N_7456);
or U8584 (N_8584,N_7161,N_7272);
nand U8585 (N_8585,N_7622,N_7274);
and U8586 (N_8586,N_7995,N_7679);
xor U8587 (N_8587,N_7358,N_7215);
nand U8588 (N_8588,N_7942,N_7934);
or U8589 (N_8589,N_7499,N_7819);
xnor U8590 (N_8590,N_7746,N_7493);
nand U8591 (N_8591,N_7078,N_7972);
nor U8592 (N_8592,N_7452,N_7478);
xor U8593 (N_8593,N_7024,N_7141);
or U8594 (N_8594,N_7821,N_7244);
nand U8595 (N_8595,N_7961,N_7300);
nand U8596 (N_8596,N_7342,N_7387);
or U8597 (N_8597,N_7484,N_7472);
nor U8598 (N_8598,N_7357,N_7554);
xor U8599 (N_8599,N_7590,N_7839);
or U8600 (N_8600,N_7961,N_7615);
nor U8601 (N_8601,N_7163,N_7502);
xor U8602 (N_8602,N_7949,N_7177);
nand U8603 (N_8603,N_7129,N_7440);
nand U8604 (N_8604,N_7430,N_7776);
nor U8605 (N_8605,N_7021,N_7727);
and U8606 (N_8606,N_7573,N_7644);
xnor U8607 (N_8607,N_7049,N_7155);
and U8608 (N_8608,N_7419,N_7967);
or U8609 (N_8609,N_7347,N_7825);
xnor U8610 (N_8610,N_7471,N_7088);
or U8611 (N_8611,N_7592,N_7431);
xor U8612 (N_8612,N_7479,N_7463);
or U8613 (N_8613,N_7573,N_7791);
nand U8614 (N_8614,N_7209,N_7473);
xnor U8615 (N_8615,N_7879,N_7815);
or U8616 (N_8616,N_7434,N_7462);
and U8617 (N_8617,N_7217,N_7419);
or U8618 (N_8618,N_7323,N_7129);
xor U8619 (N_8619,N_7540,N_7421);
nand U8620 (N_8620,N_7799,N_7886);
and U8621 (N_8621,N_7438,N_7948);
xnor U8622 (N_8622,N_7466,N_7576);
or U8623 (N_8623,N_7389,N_7879);
nor U8624 (N_8624,N_7741,N_7782);
and U8625 (N_8625,N_7174,N_7894);
xnor U8626 (N_8626,N_7243,N_7849);
nor U8627 (N_8627,N_7720,N_7381);
nor U8628 (N_8628,N_7323,N_7627);
nand U8629 (N_8629,N_7385,N_7302);
or U8630 (N_8630,N_7741,N_7522);
nor U8631 (N_8631,N_7995,N_7357);
xor U8632 (N_8632,N_7676,N_7988);
and U8633 (N_8633,N_7903,N_7690);
nand U8634 (N_8634,N_7607,N_7436);
nand U8635 (N_8635,N_7976,N_7871);
nand U8636 (N_8636,N_7577,N_7563);
or U8637 (N_8637,N_7527,N_7740);
nand U8638 (N_8638,N_7811,N_7526);
nor U8639 (N_8639,N_7244,N_7046);
xnor U8640 (N_8640,N_7044,N_7669);
and U8641 (N_8641,N_7041,N_7518);
xor U8642 (N_8642,N_7101,N_7143);
and U8643 (N_8643,N_7658,N_7463);
and U8644 (N_8644,N_7037,N_7281);
xnor U8645 (N_8645,N_7544,N_7400);
and U8646 (N_8646,N_7909,N_7041);
nand U8647 (N_8647,N_7329,N_7250);
or U8648 (N_8648,N_7318,N_7614);
and U8649 (N_8649,N_7906,N_7759);
nand U8650 (N_8650,N_7271,N_7969);
or U8651 (N_8651,N_7202,N_7679);
xnor U8652 (N_8652,N_7618,N_7578);
nor U8653 (N_8653,N_7598,N_7508);
or U8654 (N_8654,N_7186,N_7237);
nor U8655 (N_8655,N_7944,N_7251);
and U8656 (N_8656,N_7082,N_7591);
xor U8657 (N_8657,N_7304,N_7005);
and U8658 (N_8658,N_7499,N_7988);
xnor U8659 (N_8659,N_7752,N_7539);
nor U8660 (N_8660,N_7910,N_7487);
or U8661 (N_8661,N_7720,N_7654);
and U8662 (N_8662,N_7492,N_7971);
xor U8663 (N_8663,N_7125,N_7512);
nand U8664 (N_8664,N_7582,N_7146);
nor U8665 (N_8665,N_7139,N_7344);
and U8666 (N_8666,N_7971,N_7633);
or U8667 (N_8667,N_7608,N_7572);
or U8668 (N_8668,N_7835,N_7677);
xor U8669 (N_8669,N_7167,N_7834);
nor U8670 (N_8670,N_7094,N_7522);
nand U8671 (N_8671,N_7548,N_7764);
or U8672 (N_8672,N_7300,N_7241);
xor U8673 (N_8673,N_7795,N_7691);
nor U8674 (N_8674,N_7209,N_7289);
nor U8675 (N_8675,N_7740,N_7928);
or U8676 (N_8676,N_7272,N_7010);
nand U8677 (N_8677,N_7529,N_7736);
nand U8678 (N_8678,N_7531,N_7264);
xor U8679 (N_8679,N_7771,N_7145);
and U8680 (N_8680,N_7840,N_7802);
and U8681 (N_8681,N_7466,N_7512);
nand U8682 (N_8682,N_7996,N_7238);
nand U8683 (N_8683,N_7942,N_7465);
xnor U8684 (N_8684,N_7994,N_7827);
xor U8685 (N_8685,N_7527,N_7296);
and U8686 (N_8686,N_7406,N_7877);
nor U8687 (N_8687,N_7686,N_7757);
nor U8688 (N_8688,N_7177,N_7445);
nor U8689 (N_8689,N_7573,N_7181);
and U8690 (N_8690,N_7262,N_7026);
nor U8691 (N_8691,N_7501,N_7097);
xnor U8692 (N_8692,N_7665,N_7442);
or U8693 (N_8693,N_7974,N_7973);
and U8694 (N_8694,N_7467,N_7650);
and U8695 (N_8695,N_7593,N_7650);
or U8696 (N_8696,N_7799,N_7663);
nor U8697 (N_8697,N_7220,N_7899);
or U8698 (N_8698,N_7175,N_7661);
or U8699 (N_8699,N_7389,N_7656);
nor U8700 (N_8700,N_7736,N_7623);
or U8701 (N_8701,N_7924,N_7090);
nand U8702 (N_8702,N_7676,N_7620);
nor U8703 (N_8703,N_7673,N_7347);
nor U8704 (N_8704,N_7414,N_7619);
or U8705 (N_8705,N_7072,N_7581);
and U8706 (N_8706,N_7538,N_7379);
xnor U8707 (N_8707,N_7951,N_7095);
xor U8708 (N_8708,N_7846,N_7964);
or U8709 (N_8709,N_7307,N_7470);
xnor U8710 (N_8710,N_7445,N_7081);
nor U8711 (N_8711,N_7823,N_7730);
and U8712 (N_8712,N_7592,N_7499);
nand U8713 (N_8713,N_7316,N_7458);
nand U8714 (N_8714,N_7631,N_7255);
xnor U8715 (N_8715,N_7811,N_7019);
or U8716 (N_8716,N_7856,N_7968);
nand U8717 (N_8717,N_7273,N_7123);
or U8718 (N_8718,N_7061,N_7278);
nand U8719 (N_8719,N_7326,N_7928);
nand U8720 (N_8720,N_7288,N_7828);
or U8721 (N_8721,N_7753,N_7026);
nor U8722 (N_8722,N_7039,N_7165);
nand U8723 (N_8723,N_7276,N_7763);
and U8724 (N_8724,N_7472,N_7551);
or U8725 (N_8725,N_7617,N_7602);
and U8726 (N_8726,N_7300,N_7166);
xnor U8727 (N_8727,N_7434,N_7852);
or U8728 (N_8728,N_7429,N_7482);
or U8729 (N_8729,N_7791,N_7178);
and U8730 (N_8730,N_7839,N_7543);
or U8731 (N_8731,N_7160,N_7124);
nor U8732 (N_8732,N_7167,N_7057);
or U8733 (N_8733,N_7436,N_7718);
or U8734 (N_8734,N_7566,N_7285);
xor U8735 (N_8735,N_7393,N_7549);
nor U8736 (N_8736,N_7502,N_7360);
and U8737 (N_8737,N_7064,N_7201);
and U8738 (N_8738,N_7229,N_7779);
or U8739 (N_8739,N_7891,N_7116);
and U8740 (N_8740,N_7952,N_7425);
nand U8741 (N_8741,N_7992,N_7569);
or U8742 (N_8742,N_7711,N_7933);
nand U8743 (N_8743,N_7935,N_7168);
xor U8744 (N_8744,N_7033,N_7069);
nor U8745 (N_8745,N_7817,N_7889);
or U8746 (N_8746,N_7825,N_7109);
nor U8747 (N_8747,N_7220,N_7849);
xor U8748 (N_8748,N_7913,N_7846);
or U8749 (N_8749,N_7455,N_7864);
xor U8750 (N_8750,N_7132,N_7368);
nor U8751 (N_8751,N_7052,N_7117);
or U8752 (N_8752,N_7941,N_7420);
xor U8753 (N_8753,N_7694,N_7144);
and U8754 (N_8754,N_7041,N_7779);
and U8755 (N_8755,N_7653,N_7941);
nand U8756 (N_8756,N_7530,N_7819);
nor U8757 (N_8757,N_7678,N_7503);
xor U8758 (N_8758,N_7699,N_7612);
or U8759 (N_8759,N_7921,N_7812);
xor U8760 (N_8760,N_7955,N_7785);
and U8761 (N_8761,N_7228,N_7706);
nand U8762 (N_8762,N_7063,N_7966);
nor U8763 (N_8763,N_7803,N_7420);
or U8764 (N_8764,N_7115,N_7446);
nor U8765 (N_8765,N_7528,N_7076);
nor U8766 (N_8766,N_7318,N_7455);
and U8767 (N_8767,N_7552,N_7040);
nand U8768 (N_8768,N_7776,N_7476);
nand U8769 (N_8769,N_7438,N_7913);
xnor U8770 (N_8770,N_7675,N_7604);
or U8771 (N_8771,N_7745,N_7853);
xnor U8772 (N_8772,N_7543,N_7558);
and U8773 (N_8773,N_7855,N_7663);
nand U8774 (N_8774,N_7520,N_7321);
or U8775 (N_8775,N_7610,N_7155);
nor U8776 (N_8776,N_7196,N_7794);
nor U8777 (N_8777,N_7648,N_7914);
nor U8778 (N_8778,N_7806,N_7756);
nor U8779 (N_8779,N_7794,N_7555);
nor U8780 (N_8780,N_7844,N_7604);
nand U8781 (N_8781,N_7199,N_7039);
xor U8782 (N_8782,N_7874,N_7367);
nor U8783 (N_8783,N_7056,N_7343);
nand U8784 (N_8784,N_7834,N_7769);
or U8785 (N_8785,N_7893,N_7882);
nor U8786 (N_8786,N_7158,N_7598);
or U8787 (N_8787,N_7996,N_7432);
and U8788 (N_8788,N_7065,N_7478);
or U8789 (N_8789,N_7634,N_7496);
nand U8790 (N_8790,N_7837,N_7265);
nor U8791 (N_8791,N_7404,N_7130);
xnor U8792 (N_8792,N_7182,N_7002);
and U8793 (N_8793,N_7085,N_7061);
nor U8794 (N_8794,N_7653,N_7705);
or U8795 (N_8795,N_7867,N_7992);
and U8796 (N_8796,N_7554,N_7620);
or U8797 (N_8797,N_7998,N_7683);
nor U8798 (N_8798,N_7856,N_7402);
xor U8799 (N_8799,N_7435,N_7959);
and U8800 (N_8800,N_7962,N_7744);
xor U8801 (N_8801,N_7570,N_7031);
nor U8802 (N_8802,N_7136,N_7399);
xnor U8803 (N_8803,N_7178,N_7259);
and U8804 (N_8804,N_7852,N_7101);
and U8805 (N_8805,N_7099,N_7176);
or U8806 (N_8806,N_7928,N_7901);
and U8807 (N_8807,N_7205,N_7749);
nand U8808 (N_8808,N_7584,N_7734);
nand U8809 (N_8809,N_7687,N_7550);
xor U8810 (N_8810,N_7060,N_7998);
nor U8811 (N_8811,N_7806,N_7298);
nor U8812 (N_8812,N_7610,N_7149);
nand U8813 (N_8813,N_7995,N_7672);
xnor U8814 (N_8814,N_7382,N_7050);
xor U8815 (N_8815,N_7086,N_7382);
and U8816 (N_8816,N_7983,N_7107);
nor U8817 (N_8817,N_7226,N_7374);
or U8818 (N_8818,N_7715,N_7880);
or U8819 (N_8819,N_7084,N_7915);
xnor U8820 (N_8820,N_7125,N_7104);
nor U8821 (N_8821,N_7165,N_7148);
nor U8822 (N_8822,N_7917,N_7528);
xnor U8823 (N_8823,N_7896,N_7566);
and U8824 (N_8824,N_7119,N_7551);
and U8825 (N_8825,N_7170,N_7114);
and U8826 (N_8826,N_7453,N_7950);
and U8827 (N_8827,N_7529,N_7885);
nand U8828 (N_8828,N_7484,N_7153);
xor U8829 (N_8829,N_7937,N_7486);
nand U8830 (N_8830,N_7881,N_7531);
nand U8831 (N_8831,N_7321,N_7946);
nor U8832 (N_8832,N_7481,N_7812);
nor U8833 (N_8833,N_7839,N_7136);
nor U8834 (N_8834,N_7241,N_7793);
or U8835 (N_8835,N_7566,N_7385);
xnor U8836 (N_8836,N_7199,N_7293);
and U8837 (N_8837,N_7798,N_7521);
xor U8838 (N_8838,N_7762,N_7978);
or U8839 (N_8839,N_7602,N_7035);
and U8840 (N_8840,N_7147,N_7496);
or U8841 (N_8841,N_7449,N_7657);
nand U8842 (N_8842,N_7865,N_7478);
xnor U8843 (N_8843,N_7357,N_7534);
and U8844 (N_8844,N_7720,N_7610);
and U8845 (N_8845,N_7003,N_7126);
xnor U8846 (N_8846,N_7065,N_7170);
and U8847 (N_8847,N_7393,N_7991);
or U8848 (N_8848,N_7040,N_7901);
nand U8849 (N_8849,N_7203,N_7783);
nor U8850 (N_8850,N_7395,N_7853);
and U8851 (N_8851,N_7113,N_7167);
and U8852 (N_8852,N_7403,N_7896);
or U8853 (N_8853,N_7676,N_7650);
nor U8854 (N_8854,N_7514,N_7277);
and U8855 (N_8855,N_7380,N_7922);
xnor U8856 (N_8856,N_7772,N_7450);
xnor U8857 (N_8857,N_7894,N_7135);
and U8858 (N_8858,N_7470,N_7443);
nand U8859 (N_8859,N_7775,N_7940);
nand U8860 (N_8860,N_7650,N_7380);
xnor U8861 (N_8861,N_7930,N_7323);
or U8862 (N_8862,N_7685,N_7716);
or U8863 (N_8863,N_7400,N_7156);
xnor U8864 (N_8864,N_7203,N_7796);
nand U8865 (N_8865,N_7538,N_7907);
or U8866 (N_8866,N_7615,N_7191);
nor U8867 (N_8867,N_7186,N_7442);
and U8868 (N_8868,N_7994,N_7380);
or U8869 (N_8869,N_7893,N_7381);
or U8870 (N_8870,N_7370,N_7680);
and U8871 (N_8871,N_7842,N_7730);
nand U8872 (N_8872,N_7947,N_7455);
nor U8873 (N_8873,N_7098,N_7854);
xor U8874 (N_8874,N_7617,N_7051);
or U8875 (N_8875,N_7473,N_7862);
nor U8876 (N_8876,N_7590,N_7041);
or U8877 (N_8877,N_7270,N_7813);
xnor U8878 (N_8878,N_7739,N_7485);
nor U8879 (N_8879,N_7086,N_7264);
and U8880 (N_8880,N_7275,N_7241);
and U8881 (N_8881,N_7541,N_7427);
and U8882 (N_8882,N_7150,N_7323);
or U8883 (N_8883,N_7356,N_7334);
nor U8884 (N_8884,N_7664,N_7409);
and U8885 (N_8885,N_7332,N_7350);
nor U8886 (N_8886,N_7106,N_7552);
or U8887 (N_8887,N_7489,N_7542);
xor U8888 (N_8888,N_7469,N_7352);
and U8889 (N_8889,N_7435,N_7143);
and U8890 (N_8890,N_7443,N_7740);
and U8891 (N_8891,N_7719,N_7609);
nor U8892 (N_8892,N_7229,N_7244);
or U8893 (N_8893,N_7346,N_7707);
nand U8894 (N_8894,N_7335,N_7134);
nand U8895 (N_8895,N_7965,N_7229);
nand U8896 (N_8896,N_7118,N_7148);
and U8897 (N_8897,N_7757,N_7521);
or U8898 (N_8898,N_7814,N_7207);
and U8899 (N_8899,N_7123,N_7740);
nand U8900 (N_8900,N_7468,N_7195);
nand U8901 (N_8901,N_7654,N_7697);
and U8902 (N_8902,N_7212,N_7340);
nor U8903 (N_8903,N_7850,N_7806);
xor U8904 (N_8904,N_7002,N_7118);
nand U8905 (N_8905,N_7159,N_7872);
or U8906 (N_8906,N_7076,N_7109);
or U8907 (N_8907,N_7246,N_7322);
and U8908 (N_8908,N_7171,N_7259);
nor U8909 (N_8909,N_7078,N_7761);
nand U8910 (N_8910,N_7790,N_7888);
and U8911 (N_8911,N_7371,N_7164);
nor U8912 (N_8912,N_7502,N_7400);
and U8913 (N_8913,N_7733,N_7428);
xor U8914 (N_8914,N_7790,N_7243);
nand U8915 (N_8915,N_7921,N_7958);
or U8916 (N_8916,N_7325,N_7272);
xnor U8917 (N_8917,N_7236,N_7561);
or U8918 (N_8918,N_7810,N_7679);
and U8919 (N_8919,N_7448,N_7609);
nand U8920 (N_8920,N_7025,N_7279);
and U8921 (N_8921,N_7818,N_7412);
and U8922 (N_8922,N_7217,N_7932);
nand U8923 (N_8923,N_7401,N_7544);
or U8924 (N_8924,N_7397,N_7816);
or U8925 (N_8925,N_7158,N_7449);
xor U8926 (N_8926,N_7592,N_7576);
and U8927 (N_8927,N_7585,N_7511);
nor U8928 (N_8928,N_7028,N_7553);
xnor U8929 (N_8929,N_7133,N_7365);
xnor U8930 (N_8930,N_7478,N_7257);
or U8931 (N_8931,N_7277,N_7720);
xnor U8932 (N_8932,N_7138,N_7420);
nand U8933 (N_8933,N_7884,N_7429);
nand U8934 (N_8934,N_7014,N_7681);
nand U8935 (N_8935,N_7598,N_7847);
or U8936 (N_8936,N_7458,N_7210);
nor U8937 (N_8937,N_7968,N_7168);
or U8938 (N_8938,N_7294,N_7286);
nand U8939 (N_8939,N_7032,N_7082);
or U8940 (N_8940,N_7986,N_7994);
nor U8941 (N_8941,N_7278,N_7985);
and U8942 (N_8942,N_7513,N_7521);
or U8943 (N_8943,N_7441,N_7966);
nor U8944 (N_8944,N_7294,N_7463);
nand U8945 (N_8945,N_7244,N_7850);
xnor U8946 (N_8946,N_7075,N_7460);
nand U8947 (N_8947,N_7540,N_7668);
and U8948 (N_8948,N_7155,N_7020);
nor U8949 (N_8949,N_7221,N_7974);
or U8950 (N_8950,N_7473,N_7141);
nor U8951 (N_8951,N_7424,N_7026);
or U8952 (N_8952,N_7935,N_7195);
and U8953 (N_8953,N_7246,N_7825);
xnor U8954 (N_8954,N_7757,N_7893);
xor U8955 (N_8955,N_7153,N_7950);
nor U8956 (N_8956,N_7696,N_7191);
and U8957 (N_8957,N_7589,N_7542);
nand U8958 (N_8958,N_7703,N_7862);
nor U8959 (N_8959,N_7973,N_7212);
and U8960 (N_8960,N_7740,N_7617);
xnor U8961 (N_8961,N_7047,N_7110);
nand U8962 (N_8962,N_7293,N_7901);
or U8963 (N_8963,N_7610,N_7840);
nor U8964 (N_8964,N_7446,N_7458);
xor U8965 (N_8965,N_7491,N_7806);
or U8966 (N_8966,N_7081,N_7596);
or U8967 (N_8967,N_7813,N_7720);
nand U8968 (N_8968,N_7704,N_7492);
nor U8969 (N_8969,N_7015,N_7548);
nor U8970 (N_8970,N_7794,N_7288);
nor U8971 (N_8971,N_7097,N_7769);
xnor U8972 (N_8972,N_7715,N_7558);
xnor U8973 (N_8973,N_7440,N_7362);
nor U8974 (N_8974,N_7994,N_7314);
and U8975 (N_8975,N_7056,N_7704);
nor U8976 (N_8976,N_7340,N_7208);
nand U8977 (N_8977,N_7259,N_7642);
nor U8978 (N_8978,N_7079,N_7912);
nor U8979 (N_8979,N_7367,N_7952);
or U8980 (N_8980,N_7966,N_7061);
and U8981 (N_8981,N_7269,N_7611);
or U8982 (N_8982,N_7701,N_7819);
nand U8983 (N_8983,N_7154,N_7058);
or U8984 (N_8984,N_7482,N_7220);
and U8985 (N_8985,N_7722,N_7107);
and U8986 (N_8986,N_7661,N_7248);
or U8987 (N_8987,N_7474,N_7334);
nand U8988 (N_8988,N_7901,N_7411);
xor U8989 (N_8989,N_7374,N_7398);
or U8990 (N_8990,N_7085,N_7746);
nor U8991 (N_8991,N_7553,N_7640);
xor U8992 (N_8992,N_7640,N_7658);
and U8993 (N_8993,N_7483,N_7721);
xnor U8994 (N_8994,N_7846,N_7103);
or U8995 (N_8995,N_7366,N_7265);
or U8996 (N_8996,N_7265,N_7738);
xor U8997 (N_8997,N_7657,N_7889);
and U8998 (N_8998,N_7421,N_7706);
or U8999 (N_8999,N_7001,N_7219);
or U9000 (N_9000,N_8026,N_8676);
and U9001 (N_9001,N_8841,N_8797);
xor U9002 (N_9002,N_8873,N_8205);
nor U9003 (N_9003,N_8192,N_8451);
xor U9004 (N_9004,N_8601,N_8561);
xnor U9005 (N_9005,N_8622,N_8189);
and U9006 (N_9006,N_8737,N_8777);
nor U9007 (N_9007,N_8748,N_8498);
nor U9008 (N_9008,N_8068,N_8190);
or U9009 (N_9009,N_8655,N_8636);
and U9010 (N_9010,N_8215,N_8755);
or U9011 (N_9011,N_8317,N_8268);
nor U9012 (N_9012,N_8140,N_8202);
nor U9013 (N_9013,N_8828,N_8400);
xnor U9014 (N_9014,N_8009,N_8106);
and U9015 (N_9015,N_8596,N_8639);
nor U9016 (N_9016,N_8866,N_8057);
nand U9017 (N_9017,N_8193,N_8604);
or U9018 (N_9018,N_8666,N_8844);
nor U9019 (N_9019,N_8997,N_8659);
xnor U9020 (N_9020,N_8910,N_8480);
or U9021 (N_9021,N_8888,N_8329);
nor U9022 (N_9022,N_8459,N_8078);
nor U9023 (N_9023,N_8827,N_8074);
nand U9024 (N_9024,N_8183,N_8819);
nor U9025 (N_9025,N_8590,N_8710);
nor U9026 (N_9026,N_8124,N_8924);
and U9027 (N_9027,N_8226,N_8243);
or U9028 (N_9028,N_8879,N_8449);
nor U9029 (N_9029,N_8346,N_8641);
or U9030 (N_9030,N_8709,N_8892);
nand U9031 (N_9031,N_8385,N_8514);
and U9032 (N_9032,N_8576,N_8436);
nand U9033 (N_9033,N_8107,N_8743);
or U9034 (N_9034,N_8220,N_8468);
xor U9035 (N_9035,N_8472,N_8266);
and U9036 (N_9036,N_8904,N_8146);
nor U9037 (N_9037,N_8988,N_8328);
and U9038 (N_9038,N_8184,N_8872);
nor U9039 (N_9039,N_8450,N_8500);
xor U9040 (N_9040,N_8363,N_8377);
and U9041 (N_9041,N_8851,N_8335);
nand U9042 (N_9042,N_8130,N_8847);
xnor U9043 (N_9043,N_8548,N_8390);
xor U9044 (N_9044,N_8303,N_8764);
nor U9045 (N_9045,N_8504,N_8017);
nand U9046 (N_9046,N_8355,N_8144);
xnor U9047 (N_9047,N_8409,N_8447);
nor U9048 (N_9048,N_8261,N_8383);
nor U9049 (N_9049,N_8034,N_8875);
and U9050 (N_9050,N_8570,N_8458);
nor U9051 (N_9051,N_8552,N_8929);
nand U9052 (N_9052,N_8065,N_8413);
nor U9053 (N_9053,N_8248,N_8726);
nor U9054 (N_9054,N_8059,N_8652);
nand U9055 (N_9055,N_8476,N_8595);
and U9056 (N_9056,N_8708,N_8671);
xor U9057 (N_9057,N_8406,N_8286);
nor U9058 (N_9058,N_8396,N_8922);
or U9059 (N_9059,N_8153,N_8959);
or U9060 (N_9060,N_8420,N_8923);
nand U9061 (N_9061,N_8496,N_8501);
nand U9062 (N_9062,N_8740,N_8375);
xnor U9063 (N_9063,N_8485,N_8817);
or U9064 (N_9064,N_8244,N_8826);
and U9065 (N_9065,N_8667,N_8914);
or U9066 (N_9066,N_8908,N_8632);
xnor U9067 (N_9067,N_8234,N_8766);
nor U9068 (N_9068,N_8209,N_8663);
or U9069 (N_9069,N_8265,N_8233);
xnor U9070 (N_9070,N_8158,N_8870);
nor U9071 (N_9071,N_8661,N_8672);
or U9072 (N_9072,N_8763,N_8316);
or U9073 (N_9073,N_8166,N_8120);
or U9074 (N_9074,N_8195,N_8857);
or U9075 (N_9075,N_8259,N_8991);
and U9076 (N_9076,N_8681,N_8211);
and U9077 (N_9077,N_8264,N_8599);
xor U9078 (N_9078,N_8818,N_8643);
nand U9079 (N_9079,N_8654,N_8691);
nor U9080 (N_9080,N_8114,N_8855);
nor U9081 (N_9081,N_8462,N_8674);
nand U9082 (N_9082,N_8007,N_8101);
xor U9083 (N_9083,N_8902,N_8370);
xnor U9084 (N_9084,N_8055,N_8619);
and U9085 (N_9085,N_8711,N_8582);
or U9086 (N_9086,N_8275,N_8644);
and U9087 (N_9087,N_8372,N_8814);
nand U9088 (N_9088,N_8803,N_8810);
or U9089 (N_9089,N_8906,N_8345);
or U9090 (N_9090,N_8706,N_8037);
nor U9091 (N_9091,N_8634,N_8031);
nand U9092 (N_9092,N_8418,N_8829);
xnor U9093 (N_9093,N_8430,N_8796);
nand U9094 (N_9094,N_8069,N_8925);
nor U9095 (N_9095,N_8798,N_8288);
and U9096 (N_9096,N_8966,N_8327);
or U9097 (N_9097,N_8394,N_8566);
and U9098 (N_9098,N_8794,N_8675);
or U9099 (N_9099,N_8044,N_8555);
nand U9100 (N_9100,N_8313,N_8276);
nor U9101 (N_9101,N_8678,N_8035);
and U9102 (N_9102,N_8607,N_8371);
nor U9103 (N_9103,N_8123,N_8869);
nor U9104 (N_9104,N_8445,N_8089);
xnor U9105 (N_9105,N_8664,N_8121);
and U9106 (N_9106,N_8992,N_8522);
and U9107 (N_9107,N_8884,N_8323);
xnor U9108 (N_9108,N_8860,N_8455);
or U9109 (N_9109,N_8949,N_8615);
xnor U9110 (N_9110,N_8048,N_8386);
and U9111 (N_9111,N_8887,N_8544);
nor U9112 (N_9112,N_8573,N_8315);
and U9113 (N_9113,N_8354,N_8614);
and U9114 (N_9114,N_8142,N_8612);
xor U9115 (N_9115,N_8159,N_8493);
xor U9116 (N_9116,N_8568,N_8983);
nor U9117 (N_9117,N_8033,N_8403);
xnor U9118 (N_9118,N_8537,N_8361);
nand U9119 (N_9119,N_8094,N_8297);
nor U9120 (N_9120,N_8882,N_8310);
xnor U9121 (N_9121,N_8163,N_8405);
xnor U9122 (N_9122,N_8520,N_8252);
xor U9123 (N_9123,N_8382,N_8024);
or U9124 (N_9124,N_8347,N_8648);
nor U9125 (N_9125,N_8953,N_8481);
nor U9126 (N_9126,N_8425,N_8968);
nand U9127 (N_9127,N_8032,N_8433);
and U9128 (N_9128,N_8350,N_8199);
and U9129 (N_9129,N_8277,N_8490);
and U9130 (N_9130,N_8981,N_8137);
and U9131 (N_9131,N_8314,N_8115);
xnor U9132 (N_9132,N_8407,N_8917);
and U9133 (N_9133,N_8630,N_8208);
nand U9134 (N_9134,N_8918,N_8896);
xor U9135 (N_9135,N_8129,N_8658);
xnor U9136 (N_9136,N_8242,N_8541);
nor U9137 (N_9137,N_8721,N_8127);
and U9138 (N_9138,N_8526,N_8756);
xor U9139 (N_9139,N_8754,N_8172);
nand U9140 (N_9140,N_8954,N_8986);
nor U9141 (N_9141,N_8509,N_8728);
and U9142 (N_9142,N_8686,N_8185);
xor U9143 (N_9143,N_8649,N_8856);
nor U9144 (N_9144,N_8408,N_8730);
xnor U9145 (N_9145,N_8811,N_8943);
nand U9146 (N_9146,N_8003,N_8011);
and U9147 (N_9147,N_8285,N_8367);
nand U9148 (N_9148,N_8625,N_8744);
and U9149 (N_9149,N_8359,N_8998);
or U9150 (N_9150,N_8876,N_8830);
or U9151 (N_9151,N_8016,N_8928);
nand U9152 (N_9152,N_8699,N_8132);
xnor U9153 (N_9153,N_8296,N_8562);
xor U9154 (N_9154,N_8502,N_8467);
nand U9155 (N_9155,N_8336,N_8182);
nor U9156 (N_9156,N_8095,N_8116);
xor U9157 (N_9157,N_8119,N_8284);
nor U9158 (N_9158,N_8045,N_8871);
xor U9159 (N_9159,N_8201,N_8402);
xor U9160 (N_9160,N_8442,N_8391);
nand U9161 (N_9161,N_8203,N_8160);
xor U9162 (N_9162,N_8683,N_8427);
nor U9163 (N_9163,N_8001,N_8752);
or U9164 (N_9164,N_8088,N_8344);
xnor U9165 (N_9165,N_8046,N_8858);
nand U9166 (N_9166,N_8196,N_8489);
or U9167 (N_9167,N_8452,N_8620);
or U9168 (N_9168,N_8687,N_8010);
xnor U9169 (N_9169,N_8495,N_8369);
nor U9170 (N_9170,N_8042,N_8004);
nor U9171 (N_9171,N_8657,N_8602);
nor U9172 (N_9172,N_8969,N_8099);
nand U9173 (N_9173,N_8753,N_8337);
and U9174 (N_9174,N_8230,N_8030);
and U9175 (N_9175,N_8979,N_8843);
nand U9176 (N_9176,N_8349,N_8019);
or U9177 (N_9177,N_8150,N_8679);
nor U9178 (N_9178,N_8613,N_8577);
nor U9179 (N_9179,N_8651,N_8389);
or U9180 (N_9180,N_8618,N_8025);
nor U9181 (N_9181,N_8175,N_8374);
and U9182 (N_9182,N_8174,N_8775);
xor U9183 (N_9183,N_8885,N_8169);
and U9184 (N_9184,N_8536,N_8318);
or U9185 (N_9185,N_8513,N_8916);
nor U9186 (N_9186,N_8254,N_8880);
and U9187 (N_9187,N_8718,N_8801);
nor U9188 (N_9188,N_8889,N_8850);
and U9189 (N_9189,N_8028,N_8720);
or U9190 (N_9190,N_8538,N_8881);
and U9191 (N_9191,N_8689,N_8603);
xor U9192 (N_9192,N_8974,N_8308);
nor U9193 (N_9193,N_8834,N_8125);
and U9194 (N_9194,N_8897,N_8593);
and U9195 (N_9195,N_8795,N_8353);
or U9196 (N_9196,N_8417,N_8176);
nor U9197 (N_9197,N_8907,N_8940);
and U9198 (N_9198,N_8746,N_8149);
or U9199 (N_9199,N_8584,N_8020);
and U9200 (N_9200,N_8157,N_8499);
or U9201 (N_9201,N_8384,N_8839);
nand U9202 (N_9202,N_8168,N_8274);
xnor U9203 (N_9203,N_8151,N_8776);
and U9204 (N_9204,N_8682,N_8825);
or U9205 (N_9205,N_8426,N_8668);
nor U9206 (N_9206,N_8006,N_8198);
and U9207 (N_9207,N_8993,N_8236);
and U9208 (N_9208,N_8861,N_8180);
nor U9209 (N_9209,N_8022,N_8950);
or U9210 (N_9210,N_8269,N_8240);
nor U9211 (N_9211,N_8883,N_8719);
xor U9212 (N_9212,N_8808,N_8479);
and U9213 (N_9213,N_8491,N_8945);
xor U9214 (N_9214,N_8111,N_8791);
or U9215 (N_9215,N_8765,N_8271);
nand U9216 (N_9216,N_8066,N_8574);
or U9217 (N_9217,N_8340,N_8564);
nand U9218 (N_9218,N_8802,N_8809);
nor U9219 (N_9219,N_8267,N_8645);
nand U9220 (N_9220,N_8964,N_8005);
nand U9221 (N_9221,N_8926,N_8342);
nor U9222 (N_9222,N_8633,N_8348);
nor U9223 (N_9223,N_8488,N_8854);
nor U9224 (N_9224,N_8126,N_8145);
nor U9225 (N_9225,N_8283,N_8747);
nor U9226 (N_9226,N_8932,N_8665);
nand U9227 (N_9227,N_8813,N_8131);
and U9228 (N_9228,N_8421,N_8191);
or U9229 (N_9229,N_8014,N_8696);
and U9230 (N_9230,N_8250,N_8294);
or U9231 (N_9231,N_8581,N_8903);
nor U9232 (N_9232,N_8650,N_8038);
xnor U9233 (N_9233,N_8735,N_8669);
or U9234 (N_9234,N_8788,N_8996);
xor U9235 (N_9235,N_8260,N_8487);
and U9236 (N_9236,N_8840,N_8300);
nand U9237 (N_9237,N_8431,N_8521);
nand U9238 (N_9238,N_8936,N_8626);
or U9239 (N_9239,N_8097,N_8967);
or U9240 (N_9240,N_8093,N_8523);
nand U9241 (N_9241,N_8291,N_8104);
nor U9242 (N_9242,N_8213,N_8225);
nor U9243 (N_9243,N_8760,N_8734);
nand U9244 (N_9244,N_8585,N_8423);
nor U9245 (N_9245,N_8905,N_8703);
or U9246 (N_9246,N_8262,N_8771);
nor U9247 (N_9247,N_8617,N_8510);
and U9248 (N_9248,N_8051,N_8571);
nand U9249 (N_9249,N_8729,N_8334);
or U9250 (N_9250,N_8608,N_8783);
xor U9251 (N_9251,N_8273,N_8432);
nor U9252 (N_9252,N_8098,N_8457);
nor U9253 (N_9253,N_8698,N_8768);
nand U9254 (N_9254,N_8133,N_8660);
nand U9255 (N_9255,N_8990,N_8102);
or U9256 (N_9256,N_8036,N_8781);
nand U9257 (N_9257,N_8656,N_8978);
nand U9258 (N_9258,N_8219,N_8836);
nand U9259 (N_9259,N_8280,N_8404);
xor U9260 (N_9260,N_8890,N_8422);
nor U9261 (N_9261,N_8217,N_8227);
nand U9262 (N_9262,N_8087,N_8832);
nand U9263 (N_9263,N_8517,N_8930);
and U9264 (N_9264,N_8039,N_8773);
or U9265 (N_9265,N_8623,N_8567);
nor U9266 (N_9266,N_8960,N_8257);
and U9267 (N_9267,N_8272,N_8064);
or U9268 (N_9268,N_8021,N_8563);
or U9269 (N_9269,N_8662,N_8255);
or U9270 (N_9270,N_8725,N_8238);
nand U9271 (N_9271,N_8118,N_8694);
nand U9272 (N_9272,N_8973,N_8982);
xor U9273 (N_9273,N_8343,N_8944);
nand U9274 (N_9274,N_8164,N_8440);
and U9275 (N_9275,N_8901,N_8712);
or U9276 (N_9276,N_8782,N_8415);
and U9277 (N_9277,N_8456,N_8070);
nor U9278 (N_9278,N_8739,N_8597);
xor U9279 (N_9279,N_8551,N_8886);
nor U9280 (N_9280,N_8519,N_8441);
nor U9281 (N_9281,N_8939,N_8084);
xor U9282 (N_9282,N_8898,N_8148);
or U9283 (N_9283,N_8282,N_8583);
or U9284 (N_9284,N_8942,N_8780);
nand U9285 (N_9285,N_8987,N_8387);
nor U9286 (N_9286,N_8351,N_8961);
nand U9287 (N_9287,N_8061,N_8793);
nor U9288 (N_9288,N_8197,N_8256);
xor U9289 (N_9289,N_8155,N_8330);
or U9290 (N_9290,N_8690,N_8492);
nor U9291 (N_9291,N_8995,N_8779);
nand U9292 (N_9292,N_8043,N_8444);
or U9293 (N_9293,N_8933,N_8008);
nand U9294 (N_9294,N_8484,N_8688);
and U9295 (N_9295,N_8002,N_8076);
nor U9296 (N_9296,N_8304,N_8053);
xor U9297 (N_9297,N_8647,N_8716);
or U9298 (N_9298,N_8128,N_8532);
nor U9299 (N_9299,N_8471,N_8535);
or U9300 (N_9300,N_8322,N_8470);
nand U9301 (N_9301,N_8429,N_8846);
or U9302 (N_9302,N_8122,N_8139);
xnor U9303 (N_9303,N_8948,N_8392);
or U9304 (N_9304,N_8477,N_8963);
nor U9305 (N_9305,N_8062,N_8278);
xnor U9306 (N_9306,N_8999,N_8842);
and U9307 (N_9307,N_8309,N_8287);
nor U9308 (N_9308,N_8799,N_8772);
or U9309 (N_9309,N_8388,N_8245);
or U9310 (N_9310,N_8543,N_8077);
nor U9311 (N_9311,N_8741,N_8692);
xnor U9312 (N_9312,N_8539,N_8865);
nand U9313 (N_9313,N_8165,N_8326);
nor U9314 (N_9314,N_8235,N_8864);
nand U9315 (N_9315,N_8970,N_8241);
or U9316 (N_9316,N_8237,N_8357);
and U9317 (N_9317,N_8306,N_8722);
and U9318 (N_9318,N_8587,N_8732);
nor U9319 (N_9319,N_8971,N_8338);
and U9320 (N_9320,N_8414,N_8082);
nor U9321 (N_9321,N_8770,N_8727);
xnor U9322 (N_9322,N_8437,N_8497);
xnor U9323 (N_9323,N_8774,N_8767);
nor U9324 (N_9324,N_8673,N_8453);
xnor U9325 (N_9325,N_8224,N_8073);
xnor U9326 (N_9326,N_8554,N_8154);
nor U9327 (N_9327,N_8786,N_8849);
or U9328 (N_9328,N_8319,N_8919);
nor U9329 (N_9329,N_8463,N_8207);
xor U9330 (N_9330,N_8279,N_8937);
xor U9331 (N_9331,N_8815,N_8047);
nor U9332 (N_9332,N_8934,N_8320);
and U9333 (N_9333,N_8640,N_8141);
and U9334 (N_9334,N_8909,N_8560);
and U9335 (N_9335,N_8222,N_8938);
or U9336 (N_9336,N_8745,N_8258);
or U9337 (N_9337,N_8707,N_8540);
xor U9338 (N_9338,N_8096,N_8446);
nand U9339 (N_9339,N_8697,N_8460);
nor U9340 (N_9340,N_8578,N_8972);
xor U9341 (N_9341,N_8931,N_8506);
nand U9342 (N_9342,N_8511,N_8616);
nand U9343 (N_9343,N_8598,N_8704);
and U9344 (N_9344,N_8435,N_8547);
or U9345 (N_9345,N_8920,N_8181);
xnor U9346 (N_9346,N_8134,N_8758);
or U9347 (N_9347,N_8247,N_8605);
nand U9348 (N_9348,N_8913,N_8863);
nor U9349 (N_9349,N_8862,N_8516);
xnor U9350 (N_9350,N_8610,N_8528);
nor U9351 (N_9351,N_8352,N_8281);
nand U9352 (N_9352,N_8638,N_8534);
nor U9353 (N_9353,N_8290,N_8977);
nand U9354 (N_9354,N_8733,N_8980);
nand U9355 (N_9355,N_8298,N_8063);
or U9356 (N_9356,N_8805,N_8529);
nand U9357 (N_9357,N_8549,N_8067);
nor U9358 (N_9358,N_8778,N_8812);
nand U9359 (N_9359,N_8364,N_8816);
xnor U9360 (N_9360,N_8989,N_8398);
nand U9361 (N_9361,N_8356,N_8759);
and U9362 (N_9362,N_8465,N_8976);
nor U9363 (N_9363,N_8381,N_8994);
xor U9364 (N_9364,N_8899,N_8751);
or U9365 (N_9365,N_8695,N_8138);
nor U9366 (N_9366,N_8822,N_8820);
nand U9367 (N_9367,N_8731,N_8680);
xor U9368 (N_9368,N_8360,N_8027);
or U9369 (N_9369,N_8325,N_8579);
nand U9370 (N_9370,N_8443,N_8056);
and U9371 (N_9371,N_8013,N_8307);
nor U9372 (N_9372,N_8419,N_8724);
xnor U9373 (N_9373,N_8503,N_8946);
and U9374 (N_9374,N_8527,N_8079);
and U9375 (N_9375,N_8915,N_8410);
nor U9376 (N_9376,N_8210,N_8214);
and U9377 (N_9377,N_8092,N_8556);
xnor U9378 (N_9378,N_8845,N_8800);
and U9379 (N_9379,N_8592,N_8081);
nand U9380 (N_9380,N_8117,N_8693);
nor U9381 (N_9381,N_8401,N_8941);
xor U9382 (N_9382,N_8263,N_8321);
or U9383 (N_9383,N_8221,N_8545);
or U9384 (N_9384,N_8058,N_8161);
nand U9385 (N_9385,N_8110,N_8677);
xor U9386 (N_9386,N_8289,N_8685);
and U9387 (N_9387,N_8962,N_8512);
nand U9388 (N_9388,N_8050,N_8738);
nor U9389 (N_9389,N_8769,N_8804);
nand U9390 (N_9390,N_8821,N_8553);
nand U9391 (N_9391,N_8393,N_8478);
or U9392 (N_9392,N_8507,N_8473);
xor U9393 (N_9393,N_8787,N_8723);
or U9394 (N_9394,N_8984,N_8448);
nor U9395 (N_9395,N_8469,N_8293);
xnor U9396 (N_9396,N_8186,N_8380);
or U9397 (N_9397,N_8376,N_8893);
xnor U9398 (N_9398,N_8807,N_8434);
and U9399 (N_9399,N_8831,N_8609);
or U9400 (N_9400,N_8670,N_8103);
xnor U9401 (N_9401,N_8867,N_8628);
nor U9402 (N_9402,N_8653,N_8424);
nor U9403 (N_9403,N_8715,N_8086);
xnor U9404 (N_9404,N_8112,N_8249);
or U9405 (N_9405,N_8790,N_8464);
or U9406 (N_9406,N_8331,N_8223);
nand U9407 (N_9407,N_8075,N_8105);
or U9408 (N_9408,N_8108,N_8606);
and U9409 (N_9409,N_8200,N_8591);
and U9410 (N_9410,N_8789,N_8515);
nand U9411 (N_9411,N_8312,N_8594);
nor U9412 (N_9412,N_8412,N_8550);
xnor U9413 (N_9413,N_8785,N_8957);
xnor U9414 (N_9414,N_8806,N_8299);
nand U9415 (N_9415,N_8171,N_8177);
nor U9416 (N_9416,N_8702,N_8700);
and U9417 (N_9417,N_8023,N_8188);
and U9418 (N_9418,N_8365,N_8399);
and U9419 (N_9419,N_8486,N_8218);
xnor U9420 (N_9420,N_8167,N_8204);
nand U9421 (N_9421,N_8611,N_8838);
xor U9422 (N_9422,N_8428,N_8332);
or U9423 (N_9423,N_8878,N_8466);
and U9424 (N_9424,N_8091,N_8580);
nor U9425 (N_9425,N_8378,N_8530);
and U9426 (N_9426,N_8921,N_8947);
xor U9427 (N_9427,N_8178,N_8588);
nor U9428 (N_9428,N_8642,N_8736);
nor U9429 (N_9429,N_8333,N_8524);
and U9430 (N_9430,N_8018,N_8270);
or U9431 (N_9431,N_8874,N_8557);
and U9432 (N_9432,N_8109,N_8295);
xnor U9433 (N_9433,N_8952,N_8635);
or U9434 (N_9434,N_8071,N_8631);
xor U9435 (N_9435,N_8113,N_8041);
nand U9436 (N_9436,N_8085,N_8701);
or U9437 (N_9437,N_8955,N_8341);
xor U9438 (N_9438,N_8868,N_8373);
or U9439 (N_9439,N_8362,N_8216);
xor U9440 (N_9440,N_8757,N_8135);
and U9441 (N_9441,N_8531,N_8912);
xnor U9442 (N_9442,N_8232,N_8600);
nor U9443 (N_9443,N_8572,N_8156);
nor U9444 (N_9444,N_8305,N_8461);
or U9445 (N_9445,N_8368,N_8012);
and U9446 (N_9446,N_8083,N_8894);
or U9447 (N_9447,N_8891,N_8179);
or U9448 (N_9448,N_8054,N_8147);
nor U9449 (N_9449,N_8170,N_8482);
or U9450 (N_9450,N_8935,N_8558);
or U9451 (N_9451,N_8302,N_8525);
nand U9452 (N_9452,N_8956,N_8761);
xor U9453 (N_9453,N_8397,N_8251);
nand U9454 (N_9454,N_8040,N_8629);
nor U9455 (N_9455,N_8438,N_8090);
xor U9456 (N_9456,N_8714,N_8416);
nand U9457 (N_9457,N_8162,N_8015);
nand U9458 (N_9458,N_8439,N_8358);
xnor U9459 (N_9459,N_8833,N_8366);
and U9460 (N_9460,N_8231,N_8637);
nor U9461 (N_9461,N_8253,N_8080);
or U9462 (N_9462,N_8837,N_8029);
or U9463 (N_9463,N_8624,N_8852);
nand U9464 (N_9464,N_8152,N_8927);
nand U9465 (N_9465,N_8717,N_8533);
nor U9466 (N_9466,N_8494,N_8505);
nand U9467 (N_9467,N_8911,N_8762);
nand U9468 (N_9468,N_8542,N_8848);
nor U9469 (N_9469,N_8713,N_8173);
xor U9470 (N_9470,N_8749,N_8575);
or U9471 (N_9471,N_8206,N_8475);
xnor U9472 (N_9472,N_8853,N_8750);
xor U9473 (N_9473,N_8049,N_8621);
or U9474 (N_9474,N_8824,N_8292);
or U9475 (N_9475,N_8395,N_8474);
or U9476 (N_9476,N_8784,N_8705);
or U9477 (N_9477,N_8895,N_8792);
and U9478 (N_9478,N_8072,N_8229);
nand U9479 (N_9479,N_8339,N_8565);
nand U9480 (N_9480,N_8228,N_8742);
and U9481 (N_9481,N_8877,N_8965);
xnor U9482 (N_9482,N_8212,N_8975);
nor U9483 (N_9483,N_8646,N_8589);
nor U9484 (N_9484,N_8000,N_8246);
and U9485 (N_9485,N_8586,N_8859);
xor U9486 (N_9486,N_8823,N_8518);
and U9487 (N_9487,N_8379,N_8324);
nor U9488 (N_9488,N_8060,N_8143);
or U9489 (N_9489,N_8900,N_8958);
nand U9490 (N_9490,N_8627,N_8301);
xnor U9491 (N_9491,N_8187,N_8483);
xor U9492 (N_9492,N_8136,N_8684);
nand U9493 (N_9493,N_8411,N_8835);
and U9494 (N_9494,N_8569,N_8454);
nand U9495 (N_9495,N_8546,N_8951);
and U9496 (N_9496,N_8100,N_8311);
nor U9497 (N_9497,N_8239,N_8985);
nand U9498 (N_9498,N_8194,N_8508);
and U9499 (N_9499,N_8052,N_8559);
nand U9500 (N_9500,N_8498,N_8709);
and U9501 (N_9501,N_8889,N_8047);
nor U9502 (N_9502,N_8790,N_8162);
nor U9503 (N_9503,N_8675,N_8246);
xor U9504 (N_9504,N_8522,N_8907);
nand U9505 (N_9505,N_8969,N_8501);
nand U9506 (N_9506,N_8855,N_8155);
xor U9507 (N_9507,N_8044,N_8825);
nand U9508 (N_9508,N_8829,N_8624);
and U9509 (N_9509,N_8965,N_8181);
and U9510 (N_9510,N_8835,N_8355);
xor U9511 (N_9511,N_8511,N_8102);
or U9512 (N_9512,N_8540,N_8910);
xor U9513 (N_9513,N_8733,N_8803);
nor U9514 (N_9514,N_8279,N_8001);
and U9515 (N_9515,N_8633,N_8929);
nand U9516 (N_9516,N_8918,N_8429);
or U9517 (N_9517,N_8605,N_8282);
or U9518 (N_9518,N_8418,N_8213);
and U9519 (N_9519,N_8246,N_8520);
nand U9520 (N_9520,N_8721,N_8027);
and U9521 (N_9521,N_8203,N_8951);
or U9522 (N_9522,N_8372,N_8913);
nor U9523 (N_9523,N_8110,N_8416);
nand U9524 (N_9524,N_8370,N_8796);
xor U9525 (N_9525,N_8420,N_8458);
nor U9526 (N_9526,N_8855,N_8975);
xnor U9527 (N_9527,N_8064,N_8654);
nor U9528 (N_9528,N_8186,N_8011);
nand U9529 (N_9529,N_8907,N_8200);
or U9530 (N_9530,N_8696,N_8143);
nor U9531 (N_9531,N_8946,N_8569);
nor U9532 (N_9532,N_8054,N_8768);
or U9533 (N_9533,N_8763,N_8862);
and U9534 (N_9534,N_8841,N_8431);
xnor U9535 (N_9535,N_8382,N_8810);
or U9536 (N_9536,N_8217,N_8349);
or U9537 (N_9537,N_8261,N_8994);
nand U9538 (N_9538,N_8096,N_8768);
nor U9539 (N_9539,N_8439,N_8046);
nor U9540 (N_9540,N_8540,N_8026);
xnor U9541 (N_9541,N_8962,N_8807);
xnor U9542 (N_9542,N_8860,N_8142);
nor U9543 (N_9543,N_8243,N_8551);
or U9544 (N_9544,N_8503,N_8528);
xor U9545 (N_9545,N_8829,N_8539);
nand U9546 (N_9546,N_8094,N_8301);
or U9547 (N_9547,N_8137,N_8727);
or U9548 (N_9548,N_8013,N_8273);
or U9549 (N_9549,N_8842,N_8665);
xnor U9550 (N_9550,N_8707,N_8783);
nand U9551 (N_9551,N_8571,N_8812);
nand U9552 (N_9552,N_8281,N_8004);
xnor U9553 (N_9553,N_8045,N_8355);
nand U9554 (N_9554,N_8565,N_8937);
and U9555 (N_9555,N_8954,N_8905);
nand U9556 (N_9556,N_8267,N_8218);
xor U9557 (N_9557,N_8259,N_8293);
and U9558 (N_9558,N_8470,N_8189);
xor U9559 (N_9559,N_8946,N_8504);
or U9560 (N_9560,N_8489,N_8856);
xnor U9561 (N_9561,N_8231,N_8521);
and U9562 (N_9562,N_8315,N_8400);
nor U9563 (N_9563,N_8860,N_8084);
and U9564 (N_9564,N_8221,N_8244);
nor U9565 (N_9565,N_8003,N_8795);
nor U9566 (N_9566,N_8864,N_8708);
nor U9567 (N_9567,N_8812,N_8301);
nand U9568 (N_9568,N_8443,N_8390);
xnor U9569 (N_9569,N_8747,N_8615);
xnor U9570 (N_9570,N_8407,N_8528);
and U9571 (N_9571,N_8959,N_8154);
or U9572 (N_9572,N_8123,N_8124);
nand U9573 (N_9573,N_8983,N_8647);
nor U9574 (N_9574,N_8972,N_8683);
xnor U9575 (N_9575,N_8497,N_8157);
nand U9576 (N_9576,N_8770,N_8525);
nand U9577 (N_9577,N_8840,N_8959);
nor U9578 (N_9578,N_8920,N_8266);
nand U9579 (N_9579,N_8424,N_8201);
or U9580 (N_9580,N_8076,N_8126);
xnor U9581 (N_9581,N_8690,N_8626);
nor U9582 (N_9582,N_8396,N_8717);
nand U9583 (N_9583,N_8030,N_8887);
and U9584 (N_9584,N_8715,N_8626);
and U9585 (N_9585,N_8655,N_8280);
or U9586 (N_9586,N_8863,N_8975);
nor U9587 (N_9587,N_8629,N_8188);
nor U9588 (N_9588,N_8928,N_8111);
or U9589 (N_9589,N_8294,N_8969);
and U9590 (N_9590,N_8112,N_8202);
and U9591 (N_9591,N_8789,N_8489);
nor U9592 (N_9592,N_8213,N_8993);
nand U9593 (N_9593,N_8995,N_8584);
nand U9594 (N_9594,N_8022,N_8553);
nor U9595 (N_9595,N_8947,N_8486);
xnor U9596 (N_9596,N_8282,N_8323);
nand U9597 (N_9597,N_8054,N_8139);
xnor U9598 (N_9598,N_8956,N_8379);
xnor U9599 (N_9599,N_8083,N_8074);
nor U9600 (N_9600,N_8421,N_8014);
or U9601 (N_9601,N_8957,N_8358);
nand U9602 (N_9602,N_8936,N_8019);
xnor U9603 (N_9603,N_8689,N_8450);
and U9604 (N_9604,N_8228,N_8820);
nor U9605 (N_9605,N_8462,N_8375);
nor U9606 (N_9606,N_8034,N_8307);
and U9607 (N_9607,N_8810,N_8432);
nand U9608 (N_9608,N_8779,N_8900);
xor U9609 (N_9609,N_8174,N_8884);
xor U9610 (N_9610,N_8734,N_8940);
or U9611 (N_9611,N_8947,N_8968);
and U9612 (N_9612,N_8056,N_8272);
xnor U9613 (N_9613,N_8538,N_8960);
nand U9614 (N_9614,N_8044,N_8059);
xor U9615 (N_9615,N_8313,N_8007);
or U9616 (N_9616,N_8386,N_8226);
and U9617 (N_9617,N_8766,N_8907);
xor U9618 (N_9618,N_8261,N_8640);
and U9619 (N_9619,N_8374,N_8049);
xnor U9620 (N_9620,N_8577,N_8931);
xnor U9621 (N_9621,N_8844,N_8098);
xor U9622 (N_9622,N_8624,N_8989);
nand U9623 (N_9623,N_8594,N_8921);
or U9624 (N_9624,N_8515,N_8923);
or U9625 (N_9625,N_8410,N_8946);
nor U9626 (N_9626,N_8982,N_8614);
and U9627 (N_9627,N_8557,N_8202);
nand U9628 (N_9628,N_8608,N_8471);
xnor U9629 (N_9629,N_8535,N_8620);
or U9630 (N_9630,N_8210,N_8720);
nor U9631 (N_9631,N_8080,N_8018);
nand U9632 (N_9632,N_8897,N_8280);
nor U9633 (N_9633,N_8575,N_8220);
or U9634 (N_9634,N_8683,N_8328);
xor U9635 (N_9635,N_8749,N_8499);
nor U9636 (N_9636,N_8383,N_8380);
nand U9637 (N_9637,N_8919,N_8584);
nor U9638 (N_9638,N_8447,N_8173);
nand U9639 (N_9639,N_8015,N_8950);
or U9640 (N_9640,N_8228,N_8296);
or U9641 (N_9641,N_8675,N_8149);
and U9642 (N_9642,N_8485,N_8303);
nand U9643 (N_9643,N_8776,N_8263);
nor U9644 (N_9644,N_8519,N_8401);
xor U9645 (N_9645,N_8542,N_8207);
nand U9646 (N_9646,N_8037,N_8365);
or U9647 (N_9647,N_8558,N_8317);
or U9648 (N_9648,N_8876,N_8606);
nor U9649 (N_9649,N_8247,N_8095);
and U9650 (N_9650,N_8846,N_8941);
xor U9651 (N_9651,N_8260,N_8962);
nand U9652 (N_9652,N_8468,N_8978);
and U9653 (N_9653,N_8968,N_8894);
or U9654 (N_9654,N_8594,N_8745);
or U9655 (N_9655,N_8254,N_8156);
and U9656 (N_9656,N_8772,N_8878);
nand U9657 (N_9657,N_8653,N_8927);
and U9658 (N_9658,N_8774,N_8960);
xnor U9659 (N_9659,N_8507,N_8820);
nor U9660 (N_9660,N_8957,N_8192);
nor U9661 (N_9661,N_8501,N_8716);
xor U9662 (N_9662,N_8522,N_8889);
nor U9663 (N_9663,N_8827,N_8378);
and U9664 (N_9664,N_8870,N_8627);
nand U9665 (N_9665,N_8527,N_8771);
and U9666 (N_9666,N_8049,N_8358);
and U9667 (N_9667,N_8717,N_8085);
nor U9668 (N_9668,N_8117,N_8114);
nor U9669 (N_9669,N_8274,N_8082);
nor U9670 (N_9670,N_8097,N_8550);
nand U9671 (N_9671,N_8927,N_8888);
and U9672 (N_9672,N_8532,N_8055);
nor U9673 (N_9673,N_8335,N_8067);
or U9674 (N_9674,N_8968,N_8398);
xor U9675 (N_9675,N_8859,N_8857);
xnor U9676 (N_9676,N_8029,N_8739);
nand U9677 (N_9677,N_8405,N_8377);
or U9678 (N_9678,N_8128,N_8130);
and U9679 (N_9679,N_8971,N_8576);
nand U9680 (N_9680,N_8486,N_8630);
or U9681 (N_9681,N_8860,N_8332);
xor U9682 (N_9682,N_8414,N_8300);
and U9683 (N_9683,N_8668,N_8765);
or U9684 (N_9684,N_8338,N_8127);
or U9685 (N_9685,N_8671,N_8440);
nand U9686 (N_9686,N_8595,N_8939);
and U9687 (N_9687,N_8261,N_8721);
nand U9688 (N_9688,N_8590,N_8811);
or U9689 (N_9689,N_8326,N_8693);
nand U9690 (N_9690,N_8396,N_8428);
xnor U9691 (N_9691,N_8342,N_8053);
xor U9692 (N_9692,N_8793,N_8792);
or U9693 (N_9693,N_8939,N_8614);
xnor U9694 (N_9694,N_8459,N_8464);
or U9695 (N_9695,N_8786,N_8177);
nand U9696 (N_9696,N_8982,N_8027);
and U9697 (N_9697,N_8536,N_8241);
xnor U9698 (N_9698,N_8445,N_8745);
or U9699 (N_9699,N_8194,N_8846);
nand U9700 (N_9700,N_8527,N_8571);
nand U9701 (N_9701,N_8218,N_8110);
nor U9702 (N_9702,N_8483,N_8853);
or U9703 (N_9703,N_8511,N_8233);
nand U9704 (N_9704,N_8131,N_8547);
or U9705 (N_9705,N_8751,N_8245);
nand U9706 (N_9706,N_8906,N_8705);
or U9707 (N_9707,N_8959,N_8452);
or U9708 (N_9708,N_8681,N_8398);
and U9709 (N_9709,N_8860,N_8327);
or U9710 (N_9710,N_8332,N_8191);
or U9711 (N_9711,N_8377,N_8617);
nor U9712 (N_9712,N_8481,N_8243);
nor U9713 (N_9713,N_8657,N_8061);
nand U9714 (N_9714,N_8489,N_8772);
nor U9715 (N_9715,N_8939,N_8324);
xor U9716 (N_9716,N_8073,N_8663);
and U9717 (N_9717,N_8423,N_8954);
or U9718 (N_9718,N_8413,N_8030);
nand U9719 (N_9719,N_8343,N_8985);
nor U9720 (N_9720,N_8417,N_8862);
xnor U9721 (N_9721,N_8222,N_8785);
and U9722 (N_9722,N_8862,N_8490);
nor U9723 (N_9723,N_8727,N_8079);
or U9724 (N_9724,N_8939,N_8843);
and U9725 (N_9725,N_8381,N_8899);
and U9726 (N_9726,N_8515,N_8780);
nor U9727 (N_9727,N_8610,N_8952);
or U9728 (N_9728,N_8833,N_8664);
xor U9729 (N_9729,N_8477,N_8146);
or U9730 (N_9730,N_8731,N_8555);
or U9731 (N_9731,N_8917,N_8206);
nand U9732 (N_9732,N_8409,N_8494);
nor U9733 (N_9733,N_8994,N_8608);
or U9734 (N_9734,N_8602,N_8196);
or U9735 (N_9735,N_8485,N_8655);
xnor U9736 (N_9736,N_8938,N_8463);
nor U9737 (N_9737,N_8390,N_8804);
nand U9738 (N_9738,N_8183,N_8847);
nor U9739 (N_9739,N_8910,N_8610);
or U9740 (N_9740,N_8992,N_8893);
nand U9741 (N_9741,N_8918,N_8344);
or U9742 (N_9742,N_8904,N_8471);
nand U9743 (N_9743,N_8686,N_8880);
or U9744 (N_9744,N_8428,N_8371);
nor U9745 (N_9745,N_8667,N_8353);
and U9746 (N_9746,N_8314,N_8365);
nand U9747 (N_9747,N_8893,N_8779);
or U9748 (N_9748,N_8418,N_8933);
nor U9749 (N_9749,N_8428,N_8293);
nand U9750 (N_9750,N_8877,N_8090);
or U9751 (N_9751,N_8280,N_8502);
xor U9752 (N_9752,N_8752,N_8940);
or U9753 (N_9753,N_8642,N_8273);
nand U9754 (N_9754,N_8359,N_8996);
or U9755 (N_9755,N_8656,N_8520);
nand U9756 (N_9756,N_8619,N_8293);
nand U9757 (N_9757,N_8873,N_8378);
nand U9758 (N_9758,N_8620,N_8597);
nand U9759 (N_9759,N_8030,N_8808);
xor U9760 (N_9760,N_8276,N_8486);
nor U9761 (N_9761,N_8408,N_8272);
and U9762 (N_9762,N_8145,N_8691);
nand U9763 (N_9763,N_8677,N_8572);
nand U9764 (N_9764,N_8973,N_8625);
xor U9765 (N_9765,N_8562,N_8452);
xnor U9766 (N_9766,N_8336,N_8248);
nor U9767 (N_9767,N_8377,N_8375);
nand U9768 (N_9768,N_8781,N_8418);
xnor U9769 (N_9769,N_8296,N_8684);
or U9770 (N_9770,N_8441,N_8567);
nand U9771 (N_9771,N_8378,N_8180);
or U9772 (N_9772,N_8420,N_8600);
nand U9773 (N_9773,N_8298,N_8452);
nor U9774 (N_9774,N_8522,N_8537);
nand U9775 (N_9775,N_8454,N_8993);
or U9776 (N_9776,N_8441,N_8772);
nor U9777 (N_9777,N_8499,N_8063);
xor U9778 (N_9778,N_8516,N_8131);
or U9779 (N_9779,N_8427,N_8369);
xnor U9780 (N_9780,N_8268,N_8485);
or U9781 (N_9781,N_8787,N_8914);
and U9782 (N_9782,N_8865,N_8784);
xor U9783 (N_9783,N_8590,N_8164);
xor U9784 (N_9784,N_8580,N_8797);
nor U9785 (N_9785,N_8605,N_8657);
nor U9786 (N_9786,N_8346,N_8173);
nor U9787 (N_9787,N_8715,N_8140);
nor U9788 (N_9788,N_8045,N_8943);
or U9789 (N_9789,N_8593,N_8980);
or U9790 (N_9790,N_8766,N_8963);
nand U9791 (N_9791,N_8135,N_8980);
nand U9792 (N_9792,N_8555,N_8914);
and U9793 (N_9793,N_8387,N_8177);
or U9794 (N_9794,N_8324,N_8391);
xnor U9795 (N_9795,N_8249,N_8469);
nand U9796 (N_9796,N_8358,N_8861);
nand U9797 (N_9797,N_8760,N_8782);
or U9798 (N_9798,N_8334,N_8656);
nor U9799 (N_9799,N_8941,N_8905);
or U9800 (N_9800,N_8986,N_8474);
and U9801 (N_9801,N_8065,N_8101);
nand U9802 (N_9802,N_8259,N_8956);
and U9803 (N_9803,N_8818,N_8907);
nor U9804 (N_9804,N_8375,N_8785);
nand U9805 (N_9805,N_8946,N_8512);
xor U9806 (N_9806,N_8001,N_8256);
or U9807 (N_9807,N_8733,N_8986);
xor U9808 (N_9808,N_8875,N_8348);
and U9809 (N_9809,N_8362,N_8114);
xor U9810 (N_9810,N_8128,N_8421);
nor U9811 (N_9811,N_8396,N_8406);
nor U9812 (N_9812,N_8994,N_8717);
nor U9813 (N_9813,N_8600,N_8605);
nand U9814 (N_9814,N_8187,N_8669);
nor U9815 (N_9815,N_8364,N_8941);
xor U9816 (N_9816,N_8601,N_8964);
and U9817 (N_9817,N_8642,N_8277);
xor U9818 (N_9818,N_8304,N_8497);
xor U9819 (N_9819,N_8188,N_8346);
nand U9820 (N_9820,N_8809,N_8791);
or U9821 (N_9821,N_8149,N_8642);
nand U9822 (N_9822,N_8076,N_8234);
or U9823 (N_9823,N_8531,N_8056);
or U9824 (N_9824,N_8236,N_8358);
and U9825 (N_9825,N_8987,N_8335);
xnor U9826 (N_9826,N_8585,N_8846);
xnor U9827 (N_9827,N_8469,N_8119);
or U9828 (N_9828,N_8049,N_8406);
or U9829 (N_9829,N_8004,N_8850);
xnor U9830 (N_9830,N_8800,N_8837);
nor U9831 (N_9831,N_8878,N_8419);
and U9832 (N_9832,N_8181,N_8986);
or U9833 (N_9833,N_8416,N_8796);
xnor U9834 (N_9834,N_8311,N_8961);
and U9835 (N_9835,N_8381,N_8561);
nand U9836 (N_9836,N_8634,N_8216);
xor U9837 (N_9837,N_8839,N_8612);
xor U9838 (N_9838,N_8359,N_8470);
xnor U9839 (N_9839,N_8445,N_8412);
xnor U9840 (N_9840,N_8005,N_8568);
nand U9841 (N_9841,N_8231,N_8816);
and U9842 (N_9842,N_8109,N_8218);
nor U9843 (N_9843,N_8594,N_8666);
or U9844 (N_9844,N_8151,N_8722);
or U9845 (N_9845,N_8640,N_8625);
xor U9846 (N_9846,N_8806,N_8289);
and U9847 (N_9847,N_8649,N_8803);
xor U9848 (N_9848,N_8750,N_8303);
nor U9849 (N_9849,N_8400,N_8565);
xor U9850 (N_9850,N_8581,N_8479);
nand U9851 (N_9851,N_8483,N_8043);
xnor U9852 (N_9852,N_8414,N_8913);
and U9853 (N_9853,N_8984,N_8969);
nand U9854 (N_9854,N_8919,N_8968);
nand U9855 (N_9855,N_8701,N_8088);
or U9856 (N_9856,N_8095,N_8490);
nor U9857 (N_9857,N_8983,N_8519);
or U9858 (N_9858,N_8698,N_8309);
nor U9859 (N_9859,N_8771,N_8620);
and U9860 (N_9860,N_8608,N_8388);
nand U9861 (N_9861,N_8865,N_8739);
nor U9862 (N_9862,N_8186,N_8383);
or U9863 (N_9863,N_8817,N_8685);
nor U9864 (N_9864,N_8828,N_8964);
nand U9865 (N_9865,N_8637,N_8232);
and U9866 (N_9866,N_8115,N_8075);
nand U9867 (N_9867,N_8475,N_8910);
or U9868 (N_9868,N_8785,N_8581);
nand U9869 (N_9869,N_8277,N_8993);
nand U9870 (N_9870,N_8172,N_8339);
nor U9871 (N_9871,N_8880,N_8016);
nand U9872 (N_9872,N_8187,N_8420);
or U9873 (N_9873,N_8112,N_8470);
and U9874 (N_9874,N_8864,N_8529);
nand U9875 (N_9875,N_8521,N_8492);
or U9876 (N_9876,N_8848,N_8979);
nor U9877 (N_9877,N_8160,N_8946);
nor U9878 (N_9878,N_8102,N_8427);
nor U9879 (N_9879,N_8576,N_8459);
or U9880 (N_9880,N_8220,N_8526);
and U9881 (N_9881,N_8791,N_8333);
and U9882 (N_9882,N_8712,N_8123);
xor U9883 (N_9883,N_8441,N_8187);
nor U9884 (N_9884,N_8795,N_8347);
nor U9885 (N_9885,N_8923,N_8728);
and U9886 (N_9886,N_8924,N_8979);
or U9887 (N_9887,N_8626,N_8164);
nor U9888 (N_9888,N_8911,N_8880);
nor U9889 (N_9889,N_8020,N_8664);
nor U9890 (N_9890,N_8374,N_8250);
nor U9891 (N_9891,N_8228,N_8210);
nand U9892 (N_9892,N_8106,N_8170);
and U9893 (N_9893,N_8433,N_8683);
and U9894 (N_9894,N_8557,N_8354);
nor U9895 (N_9895,N_8375,N_8842);
nor U9896 (N_9896,N_8293,N_8946);
xnor U9897 (N_9897,N_8950,N_8828);
or U9898 (N_9898,N_8594,N_8959);
nor U9899 (N_9899,N_8004,N_8791);
and U9900 (N_9900,N_8243,N_8946);
nand U9901 (N_9901,N_8769,N_8485);
or U9902 (N_9902,N_8076,N_8787);
or U9903 (N_9903,N_8321,N_8268);
or U9904 (N_9904,N_8927,N_8316);
nand U9905 (N_9905,N_8149,N_8605);
nor U9906 (N_9906,N_8985,N_8559);
and U9907 (N_9907,N_8148,N_8151);
nor U9908 (N_9908,N_8144,N_8110);
nor U9909 (N_9909,N_8693,N_8490);
and U9910 (N_9910,N_8856,N_8860);
xnor U9911 (N_9911,N_8689,N_8423);
nand U9912 (N_9912,N_8337,N_8833);
xnor U9913 (N_9913,N_8892,N_8256);
and U9914 (N_9914,N_8133,N_8763);
nand U9915 (N_9915,N_8951,N_8649);
xor U9916 (N_9916,N_8612,N_8382);
nor U9917 (N_9917,N_8068,N_8755);
and U9918 (N_9918,N_8545,N_8841);
and U9919 (N_9919,N_8165,N_8978);
and U9920 (N_9920,N_8760,N_8772);
or U9921 (N_9921,N_8311,N_8043);
and U9922 (N_9922,N_8609,N_8201);
xor U9923 (N_9923,N_8905,N_8787);
xnor U9924 (N_9924,N_8254,N_8889);
or U9925 (N_9925,N_8896,N_8476);
and U9926 (N_9926,N_8371,N_8220);
and U9927 (N_9927,N_8303,N_8664);
and U9928 (N_9928,N_8976,N_8648);
xnor U9929 (N_9929,N_8450,N_8877);
nor U9930 (N_9930,N_8122,N_8865);
or U9931 (N_9931,N_8688,N_8546);
and U9932 (N_9932,N_8441,N_8047);
nand U9933 (N_9933,N_8595,N_8483);
or U9934 (N_9934,N_8191,N_8646);
nand U9935 (N_9935,N_8106,N_8242);
and U9936 (N_9936,N_8689,N_8584);
nand U9937 (N_9937,N_8932,N_8382);
nor U9938 (N_9938,N_8583,N_8777);
nor U9939 (N_9939,N_8007,N_8133);
nand U9940 (N_9940,N_8293,N_8578);
nor U9941 (N_9941,N_8657,N_8455);
xnor U9942 (N_9942,N_8163,N_8906);
xnor U9943 (N_9943,N_8964,N_8511);
nand U9944 (N_9944,N_8430,N_8548);
xnor U9945 (N_9945,N_8312,N_8038);
or U9946 (N_9946,N_8242,N_8269);
xnor U9947 (N_9947,N_8825,N_8982);
and U9948 (N_9948,N_8758,N_8277);
nor U9949 (N_9949,N_8000,N_8995);
nor U9950 (N_9950,N_8750,N_8690);
xnor U9951 (N_9951,N_8827,N_8896);
xnor U9952 (N_9952,N_8855,N_8857);
nand U9953 (N_9953,N_8569,N_8638);
nor U9954 (N_9954,N_8669,N_8804);
nand U9955 (N_9955,N_8335,N_8148);
or U9956 (N_9956,N_8320,N_8650);
or U9957 (N_9957,N_8863,N_8849);
xor U9958 (N_9958,N_8636,N_8353);
or U9959 (N_9959,N_8110,N_8683);
xnor U9960 (N_9960,N_8144,N_8902);
nor U9961 (N_9961,N_8866,N_8762);
nor U9962 (N_9962,N_8092,N_8035);
or U9963 (N_9963,N_8464,N_8658);
and U9964 (N_9964,N_8209,N_8109);
nor U9965 (N_9965,N_8956,N_8582);
xnor U9966 (N_9966,N_8152,N_8962);
and U9967 (N_9967,N_8067,N_8751);
nor U9968 (N_9968,N_8601,N_8138);
nor U9969 (N_9969,N_8211,N_8031);
xnor U9970 (N_9970,N_8866,N_8596);
xor U9971 (N_9971,N_8557,N_8568);
xor U9972 (N_9972,N_8062,N_8148);
nand U9973 (N_9973,N_8560,N_8673);
or U9974 (N_9974,N_8600,N_8510);
nand U9975 (N_9975,N_8582,N_8944);
and U9976 (N_9976,N_8081,N_8491);
nand U9977 (N_9977,N_8942,N_8796);
nor U9978 (N_9978,N_8083,N_8728);
nand U9979 (N_9979,N_8987,N_8353);
or U9980 (N_9980,N_8663,N_8645);
xnor U9981 (N_9981,N_8823,N_8485);
nor U9982 (N_9982,N_8783,N_8753);
nor U9983 (N_9983,N_8787,N_8678);
nor U9984 (N_9984,N_8782,N_8422);
or U9985 (N_9985,N_8563,N_8204);
and U9986 (N_9986,N_8003,N_8617);
xor U9987 (N_9987,N_8398,N_8841);
xnor U9988 (N_9988,N_8707,N_8123);
nor U9989 (N_9989,N_8397,N_8328);
or U9990 (N_9990,N_8837,N_8874);
and U9991 (N_9991,N_8868,N_8840);
or U9992 (N_9992,N_8529,N_8185);
and U9993 (N_9993,N_8854,N_8808);
or U9994 (N_9994,N_8730,N_8281);
nor U9995 (N_9995,N_8987,N_8622);
and U9996 (N_9996,N_8066,N_8280);
and U9997 (N_9997,N_8492,N_8916);
nand U9998 (N_9998,N_8755,N_8781);
nand U9999 (N_9999,N_8511,N_8142);
or U10000 (N_10000,N_9199,N_9542);
xnor U10001 (N_10001,N_9053,N_9195);
nor U10002 (N_10002,N_9984,N_9055);
or U10003 (N_10003,N_9746,N_9952);
nor U10004 (N_10004,N_9016,N_9694);
xor U10005 (N_10005,N_9044,N_9815);
nor U10006 (N_10006,N_9159,N_9413);
nor U10007 (N_10007,N_9294,N_9616);
or U10008 (N_10008,N_9477,N_9880);
and U10009 (N_10009,N_9622,N_9111);
nor U10010 (N_10010,N_9029,N_9783);
and U10011 (N_10011,N_9970,N_9757);
xor U10012 (N_10012,N_9104,N_9089);
and U10013 (N_10013,N_9212,N_9866);
nor U10014 (N_10014,N_9310,N_9998);
nand U10015 (N_10015,N_9821,N_9057);
xor U10016 (N_10016,N_9000,N_9283);
nor U10017 (N_10017,N_9606,N_9278);
xnor U10018 (N_10018,N_9877,N_9617);
nor U10019 (N_10019,N_9560,N_9767);
and U10020 (N_10020,N_9474,N_9811);
or U10021 (N_10021,N_9657,N_9682);
nand U10022 (N_10022,N_9257,N_9013);
and U10023 (N_10023,N_9108,N_9752);
and U10024 (N_10024,N_9393,N_9776);
and U10025 (N_10025,N_9087,N_9434);
xor U10026 (N_10026,N_9962,N_9589);
nand U10027 (N_10027,N_9018,N_9848);
nand U10028 (N_10028,N_9178,N_9058);
xnor U10029 (N_10029,N_9748,N_9620);
nand U10030 (N_10030,N_9336,N_9530);
and U10031 (N_10031,N_9100,N_9714);
nand U10032 (N_10032,N_9960,N_9595);
and U10033 (N_10033,N_9325,N_9750);
nand U10034 (N_10034,N_9311,N_9799);
nand U10035 (N_10035,N_9677,N_9295);
and U10036 (N_10036,N_9569,N_9365);
nor U10037 (N_10037,N_9581,N_9446);
and U10038 (N_10038,N_9771,N_9025);
nor U10039 (N_10039,N_9741,N_9071);
or U10040 (N_10040,N_9476,N_9399);
and U10041 (N_10041,N_9534,N_9461);
nand U10042 (N_10042,N_9355,N_9395);
and U10043 (N_10043,N_9743,N_9472);
or U10044 (N_10044,N_9964,N_9286);
or U10045 (N_10045,N_9133,N_9538);
nand U10046 (N_10046,N_9322,N_9320);
nor U10047 (N_10047,N_9500,N_9402);
nor U10048 (N_10048,N_9379,N_9838);
nand U10049 (N_10049,N_9759,N_9908);
or U10050 (N_10050,N_9234,N_9239);
and U10051 (N_10051,N_9463,N_9011);
or U10052 (N_10052,N_9307,N_9897);
and U10053 (N_10053,N_9468,N_9818);
nor U10054 (N_10054,N_9223,N_9527);
nand U10055 (N_10055,N_9823,N_9408);
and U10056 (N_10056,N_9571,N_9782);
nor U10057 (N_10057,N_9374,N_9705);
nand U10058 (N_10058,N_9174,N_9966);
and U10059 (N_10059,N_9600,N_9593);
nand U10060 (N_10060,N_9351,N_9774);
and U10061 (N_10061,N_9906,N_9037);
or U10062 (N_10062,N_9301,N_9331);
xnor U10063 (N_10063,N_9574,N_9202);
xor U10064 (N_10064,N_9482,N_9917);
nor U10065 (N_10065,N_9932,N_9891);
nor U10066 (N_10066,N_9192,N_9441);
and U10067 (N_10067,N_9364,N_9047);
nor U10068 (N_10068,N_9819,N_9352);
xnor U10069 (N_10069,N_9868,N_9388);
and U10070 (N_10070,N_9885,N_9222);
or U10071 (N_10071,N_9024,N_9656);
or U10072 (N_10072,N_9967,N_9489);
xnor U10073 (N_10073,N_9665,N_9471);
or U10074 (N_10074,N_9856,N_9997);
nor U10075 (N_10075,N_9221,N_9158);
nand U10076 (N_10076,N_9084,N_9603);
nand U10077 (N_10077,N_9840,N_9807);
nor U10078 (N_10078,N_9288,N_9266);
or U10079 (N_10079,N_9640,N_9503);
and U10080 (N_10080,N_9319,N_9430);
nor U10081 (N_10081,N_9107,N_9899);
nand U10082 (N_10082,N_9973,N_9834);
nand U10083 (N_10083,N_9380,N_9141);
nor U10084 (N_10084,N_9117,N_9654);
or U10085 (N_10085,N_9719,N_9685);
nor U10086 (N_10086,N_9812,N_9465);
nor U10087 (N_10087,N_9647,N_9337);
nand U10088 (N_10088,N_9568,N_9988);
nand U10089 (N_10089,N_9762,N_9933);
nand U10090 (N_10090,N_9959,N_9918);
and U10091 (N_10091,N_9761,N_9710);
and U10092 (N_10092,N_9144,N_9299);
xnor U10093 (N_10093,N_9314,N_9069);
and U10094 (N_10094,N_9995,N_9781);
xnor U10095 (N_10095,N_9093,N_9930);
xor U10096 (N_10096,N_9232,N_9189);
xor U10097 (N_10097,N_9258,N_9638);
or U10098 (N_10098,N_9550,N_9254);
nand U10099 (N_10099,N_9562,N_9733);
and U10100 (N_10100,N_9711,N_9666);
nor U10101 (N_10101,N_9553,N_9376);
xnor U10102 (N_10102,N_9367,N_9464);
nand U10103 (N_10103,N_9173,N_9923);
nand U10104 (N_10104,N_9318,N_9080);
nand U10105 (N_10105,N_9241,N_9925);
nor U10106 (N_10106,N_9936,N_9006);
nor U10107 (N_10107,N_9371,N_9479);
nor U10108 (N_10108,N_9113,N_9309);
nor U10109 (N_10109,N_9884,N_9305);
xnor U10110 (N_10110,N_9172,N_9440);
xnor U10111 (N_10111,N_9341,N_9516);
and U10112 (N_10112,N_9313,N_9914);
nor U10113 (N_10113,N_9456,N_9700);
xor U10114 (N_10114,N_9297,N_9533);
xnor U10115 (N_10115,N_9378,N_9801);
xnor U10116 (N_10116,N_9846,N_9233);
nor U10117 (N_10117,N_9122,N_9974);
nor U10118 (N_10118,N_9484,N_9702);
nor U10119 (N_10119,N_9033,N_9354);
nor U10120 (N_10120,N_9728,N_9680);
xor U10121 (N_10121,N_9327,N_9594);
nand U10122 (N_10122,N_9109,N_9428);
or U10123 (N_10123,N_9835,N_9391);
xnor U10124 (N_10124,N_9583,N_9343);
xnor U10125 (N_10125,N_9804,N_9602);
xor U10126 (N_10126,N_9153,N_9177);
and U10127 (N_10127,N_9439,N_9887);
and U10128 (N_10128,N_9727,N_9264);
and U10129 (N_10129,N_9422,N_9253);
nand U10130 (N_10130,N_9131,N_9099);
nand U10131 (N_10131,N_9851,N_9892);
or U10132 (N_10132,N_9675,N_9853);
nand U10133 (N_10133,N_9777,N_9809);
nor U10134 (N_10134,N_9123,N_9490);
or U10135 (N_10135,N_9734,N_9870);
and U10136 (N_10136,N_9458,N_9546);
nand U10137 (N_10137,N_9027,N_9163);
or U10138 (N_10138,N_9949,N_9921);
nand U10139 (N_10139,N_9849,N_9514);
or U10140 (N_10140,N_9206,N_9034);
xnor U10141 (N_10141,N_9911,N_9340);
xnor U10142 (N_10142,N_9041,N_9825);
or U10143 (N_10143,N_9878,N_9764);
and U10144 (N_10144,N_9971,N_9115);
xnor U10145 (N_10145,N_9986,N_9448);
or U10146 (N_10146,N_9713,N_9788);
xor U10147 (N_10147,N_9779,N_9097);
or U10148 (N_10148,N_9180,N_9416);
nand U10149 (N_10149,N_9999,N_9709);
nor U10150 (N_10150,N_9769,N_9551);
nand U10151 (N_10151,N_9447,N_9548);
nor U10152 (N_10152,N_9910,N_9085);
or U10153 (N_10153,N_9052,N_9614);
nand U10154 (N_10154,N_9704,N_9338);
nand U10155 (N_10155,N_9086,N_9857);
or U10156 (N_10156,N_9633,N_9867);
xnor U10157 (N_10157,N_9247,N_9142);
and U10158 (N_10158,N_9648,N_9755);
or U10159 (N_10159,N_9631,N_9604);
nand U10160 (N_10160,N_9082,N_9237);
and U10161 (N_10161,N_9738,N_9147);
nand U10162 (N_10162,N_9907,N_9356);
nand U10163 (N_10163,N_9487,N_9929);
or U10164 (N_10164,N_9865,N_9420);
and U10165 (N_10165,N_9187,N_9235);
and U10166 (N_10166,N_9671,N_9976);
xor U10167 (N_10167,N_9164,N_9658);
or U10168 (N_10168,N_9676,N_9483);
and U10169 (N_10169,N_9020,N_9268);
xor U10170 (N_10170,N_9717,N_9270);
xor U10171 (N_10171,N_9035,N_9506);
xor U10172 (N_10172,N_9160,N_9968);
nor U10173 (N_10173,N_9893,N_9394);
nor U10174 (N_10174,N_9813,N_9475);
and U10175 (N_10175,N_9599,N_9276);
nand U10176 (N_10176,N_9359,N_9040);
nor U10177 (N_10177,N_9512,N_9522);
or U10178 (N_10178,N_9135,N_9580);
and U10179 (N_10179,N_9635,N_9398);
or U10180 (N_10180,N_9207,N_9118);
and U10181 (N_10181,N_9150,N_9888);
nand U10182 (N_10182,N_9363,N_9768);
and U10183 (N_10183,N_9121,N_9498);
nor U10184 (N_10184,N_9358,N_9156);
or U10185 (N_10185,N_9050,N_9065);
nor U10186 (N_10186,N_9260,N_9944);
nand U10187 (N_10187,N_9170,N_9735);
nor U10188 (N_10188,N_9256,N_9438);
xnor U10189 (N_10189,N_9280,N_9443);
nor U10190 (N_10190,N_9238,N_9820);
or U10191 (N_10191,N_9598,N_9674);
xnor U10192 (N_10192,N_9154,N_9397);
or U10193 (N_10193,N_9725,N_9308);
nor U10194 (N_10194,N_9655,N_9060);
or U10195 (N_10195,N_9218,N_9077);
nor U10196 (N_10196,N_9136,N_9566);
xnor U10197 (N_10197,N_9303,N_9555);
or U10198 (N_10198,N_9271,N_9753);
xnor U10199 (N_10199,N_9196,N_9003);
xnor U10200 (N_10200,N_9272,N_9083);
nand U10201 (N_10201,N_9149,N_9789);
and U10202 (N_10202,N_9756,N_9185);
or U10203 (N_10203,N_9822,N_9990);
xor U10204 (N_10204,N_9227,N_9491);
nand U10205 (N_10205,N_9079,N_9766);
nor U10206 (N_10206,N_9072,N_9208);
and U10207 (N_10207,N_9537,N_9396);
nand U10208 (N_10208,N_9520,N_9883);
nor U10209 (N_10209,N_9942,N_9197);
nand U10210 (N_10210,N_9210,N_9216);
or U10211 (N_10211,N_9745,N_9132);
xor U10212 (N_10212,N_9444,N_9151);
nor U10213 (N_10213,N_9670,N_9882);
nand U10214 (N_10214,N_9179,N_9146);
nor U10215 (N_10215,N_9102,N_9977);
and U10216 (N_10216,N_9316,N_9559);
nand U10217 (N_10217,N_9261,N_9827);
nand U10218 (N_10218,N_9507,N_9695);
and U10219 (N_10219,N_9576,N_9852);
and U10220 (N_10220,N_9505,N_9019);
xor U10221 (N_10221,N_9112,N_9532);
nand U10222 (N_10222,N_9703,N_9333);
xnor U10223 (N_10223,N_9161,N_9722);
xor U10224 (N_10224,N_9412,N_9833);
nand U10225 (N_10225,N_9454,N_9424);
xnor U10226 (N_10226,N_9690,N_9592);
nand U10227 (N_10227,N_9611,N_9610);
nor U10228 (N_10228,N_9961,N_9262);
nor U10229 (N_10229,N_9431,N_9074);
xnor U10230 (N_10230,N_9947,N_9090);
xor U10231 (N_10231,N_9526,N_9517);
xor U10232 (N_10232,N_9720,N_9850);
xnor U10233 (N_10233,N_9826,N_9134);
xor U10234 (N_10234,N_9950,N_9513);
nor U10235 (N_10235,N_9978,N_9552);
xor U10236 (N_10236,N_9404,N_9637);
and U10237 (N_10237,N_9110,N_9708);
xnor U10238 (N_10238,N_9284,N_9392);
or U10239 (N_10239,N_9073,N_9693);
xor U10240 (N_10240,N_9228,N_9903);
nand U10241 (N_10241,N_9473,N_9148);
nand U10242 (N_10242,N_9101,N_9323);
xnor U10243 (N_10243,N_9059,N_9528);
nor U10244 (N_10244,N_9747,N_9860);
and U10245 (N_10245,N_9591,N_9778);
and U10246 (N_10246,N_9858,N_9525);
xnor U10247 (N_10247,N_9433,N_9401);
nand U10248 (N_10248,N_9678,N_9524);
nor U10249 (N_10249,N_9895,N_9641);
and U10250 (N_10250,N_9429,N_9415);
or U10251 (N_10251,N_9051,N_9608);
xor U10252 (N_10252,N_9017,N_9829);
nor U10253 (N_10253,N_9935,N_9467);
xnor U10254 (N_10254,N_9014,N_9138);
nand U10255 (N_10255,N_9282,N_9837);
and U10256 (N_10256,N_9924,N_9855);
xnor U10257 (N_10257,N_9381,N_9938);
and U10258 (N_10258,N_9981,N_9493);
or U10259 (N_10259,N_9502,N_9230);
xnor U10260 (N_10260,N_9549,N_9008);
xor U10261 (N_10261,N_9066,N_9469);
nor U10262 (N_10262,N_9578,N_9347);
and U10263 (N_10263,N_9605,N_9830);
nand U10264 (N_10264,N_9405,N_9321);
and U10265 (N_10265,N_9031,N_9499);
xnor U10266 (N_10266,N_9445,N_9492);
xor U10267 (N_10267,N_9902,N_9417);
xnor U10268 (N_10268,N_9645,N_9758);
nand U10269 (N_10269,N_9784,N_9958);
xor U10270 (N_10270,N_9361,N_9712);
nand U10271 (N_10271,N_9863,N_9689);
or U10272 (N_10272,N_9688,N_9561);
nor U10273 (N_10273,N_9890,N_9383);
xor U10274 (N_10274,N_9010,N_9511);
nand U10275 (N_10275,N_9824,N_9406);
nand U10276 (N_10276,N_9803,N_9466);
and U10277 (N_10277,N_9194,N_9400);
or U10278 (N_10278,N_9535,N_9353);
or U10279 (N_10279,N_9937,N_9248);
xnor U10280 (N_10280,N_9198,N_9558);
and U10281 (N_10281,N_9162,N_9718);
xor U10282 (N_10282,N_9274,N_9975);
or U10283 (N_10283,N_9168,N_9231);
xor U10284 (N_10284,N_9630,N_9531);
and U10285 (N_10285,N_9012,N_9368);
nor U10286 (N_10286,N_9488,N_9296);
xnor U10287 (N_10287,N_9106,N_9350);
nand U10288 (N_10288,N_9504,N_9165);
nand U10289 (N_10289,N_9565,N_9817);
and U10290 (N_10290,N_9715,N_9991);
nor U10291 (N_10291,N_9387,N_9686);
and U10292 (N_10292,N_9965,N_9729);
nand U10293 (N_10293,N_9459,N_9009);
nor U10294 (N_10294,N_9203,N_9171);
and U10295 (N_10295,N_9273,N_9796);
nand U10296 (N_10296,N_9518,N_9544);
xor U10297 (N_10297,N_9847,N_9201);
nor U10298 (N_10298,N_9623,N_9983);
nor U10299 (N_10299,N_9864,N_9931);
and U10300 (N_10300,N_9030,N_9453);
nor U10301 (N_10301,N_9114,N_9618);
nor U10302 (N_10302,N_9026,N_9214);
xnor U10303 (N_10303,N_9760,N_9423);
and U10304 (N_10304,N_9332,N_9668);
nand U10305 (N_10305,N_9841,N_9795);
nand U10306 (N_10306,N_9786,N_9844);
nor U10307 (N_10307,N_9798,N_9845);
nor U10308 (N_10308,N_9259,N_9979);
and U10309 (N_10309,N_9426,N_9628);
and U10310 (N_10310,N_9881,N_9765);
and U10311 (N_10311,N_9495,N_9805);
xnor U10312 (N_10312,N_9501,N_9780);
nand U10313 (N_10313,N_9128,N_9244);
and U10314 (N_10314,N_9486,N_9269);
xnor U10315 (N_10315,N_9349,N_9775);
nor U10316 (N_10316,N_9963,N_9792);
or U10317 (N_10317,N_9176,N_9127);
nand U10318 (N_10318,N_9157,N_9669);
xnor U10319 (N_10319,N_9389,N_9063);
xnor U10320 (N_10320,N_9442,N_9816);
or U10321 (N_10321,N_9373,N_9224);
or U10322 (N_10322,N_9457,N_9872);
or U10323 (N_10323,N_9831,N_9229);
and U10324 (N_10324,N_9586,N_9450);
xnor U10325 (N_10325,N_9225,N_9994);
nand U10326 (N_10326,N_9992,N_9624);
nand U10327 (N_10327,N_9679,N_9478);
and U10328 (N_10328,N_9683,N_9627);
nor U10329 (N_10329,N_9739,N_9707);
nand U10330 (N_10330,N_9190,N_9793);
nor U10331 (N_10331,N_9904,N_9091);
or U10332 (N_10332,N_9545,N_9357);
and U10333 (N_10333,N_9724,N_9455);
and U10334 (N_10334,N_9873,N_9653);
nor U10335 (N_10335,N_9875,N_9510);
and U10336 (N_10336,N_9951,N_9167);
and U10337 (N_10337,N_9421,N_9183);
and U10338 (N_10338,N_9103,N_9279);
and U10339 (N_10339,N_9732,N_9362);
and U10340 (N_10340,N_9001,N_9480);
or U10341 (N_10341,N_9621,N_9054);
xor U10342 (N_10342,N_9905,N_9191);
nand U10343 (N_10343,N_9096,N_9081);
nand U10344 (N_10344,N_9706,N_9042);
nand U10345 (N_10345,N_9579,N_9411);
and U10346 (N_10346,N_9806,N_9912);
and U10347 (N_10347,N_9889,N_9263);
and U10348 (N_10348,N_9632,N_9539);
nor U10349 (N_10349,N_9215,N_9650);
nand U10350 (N_10350,N_9032,N_9140);
nand U10351 (N_10351,N_9245,N_9219);
nand U10352 (N_10352,N_9088,N_9808);
and U10353 (N_10353,N_9927,N_9265);
and U10354 (N_10354,N_9521,N_9554);
and U10355 (N_10355,N_9312,N_9763);
nor U10356 (N_10356,N_9585,N_9129);
nand U10357 (N_10357,N_9384,N_9175);
xor U10358 (N_10358,N_9291,N_9497);
or U10359 (N_10359,N_9036,N_9220);
and U10360 (N_10360,N_9372,N_9943);
or U10361 (N_10361,N_9414,N_9701);
xor U10362 (N_10362,N_9800,N_9920);
nor U10363 (N_10363,N_9095,N_9615);
and U10364 (N_10364,N_9660,N_9543);
or U10365 (N_10365,N_9980,N_9425);
xnor U10366 (N_10366,N_9723,N_9957);
or U10367 (N_10367,N_9540,N_9125);
nand U10368 (N_10368,N_9567,N_9346);
nor U10369 (N_10369,N_9246,N_9344);
or U10370 (N_10370,N_9049,N_9590);
and U10371 (N_10371,N_9646,N_9730);
or U10372 (N_10372,N_9452,N_9289);
xnor U10373 (N_10373,N_9120,N_9787);
nor U10374 (N_10374,N_9587,N_9664);
or U10375 (N_10375,N_9205,N_9370);
nor U10376 (N_10376,N_9919,N_9076);
nor U10377 (N_10377,N_9005,N_9588);
nand U10378 (N_10378,N_9330,N_9427);
nand U10379 (N_10379,N_9302,N_9754);
xor U10380 (N_10380,N_9298,N_9240);
or U10381 (N_10381,N_9326,N_9915);
or U10382 (N_10382,N_9629,N_9437);
nand U10383 (N_10383,N_9068,N_9744);
xnor U10384 (N_10384,N_9900,N_9304);
or U10385 (N_10385,N_9557,N_9691);
or U10386 (N_10386,N_9573,N_9048);
nor U10387 (N_10387,N_9075,N_9619);
nand U10388 (N_10388,N_9625,N_9896);
or U10389 (N_10389,N_9249,N_9987);
and U10390 (N_10390,N_9460,N_9038);
nor U10391 (N_10391,N_9989,N_9993);
and U10392 (N_10392,N_9064,N_9105);
xnor U10393 (N_10393,N_9021,N_9751);
and U10394 (N_10394,N_9861,N_9596);
nand U10395 (N_10395,N_9577,N_9281);
or U10396 (N_10396,N_9267,N_9785);
xnor U10397 (N_10397,N_9403,N_9901);
and U10398 (N_10398,N_9386,N_9143);
nand U10399 (N_10399,N_9334,N_9366);
or U10400 (N_10400,N_9382,N_9290);
nand U10401 (N_10401,N_9854,N_9092);
and U10402 (N_10402,N_9409,N_9547);
nor U10403 (N_10403,N_9285,N_9582);
or U10404 (N_10404,N_9939,N_9662);
nand U10405 (N_10405,N_9390,N_9200);
nand U10406 (N_10406,N_9070,N_9494);
nor U10407 (N_10407,N_9345,N_9697);
and U10408 (N_10408,N_9335,N_9661);
nor U10409 (N_10409,N_9874,N_9955);
and U10410 (N_10410,N_9842,N_9859);
or U10411 (N_10411,N_9002,N_9242);
xnor U10412 (N_10412,N_9342,N_9023);
nor U10413 (N_10413,N_9300,N_9721);
nor U10414 (N_10414,N_9509,N_9226);
nand U10415 (N_10415,N_9007,N_9287);
nor U10416 (N_10416,N_9996,N_9740);
and U10417 (N_10417,N_9663,N_9687);
and U10418 (N_10418,N_9410,N_9209);
xnor U10419 (N_10419,N_9022,N_9916);
nand U10420 (N_10420,N_9435,N_9251);
xor U10421 (N_10421,N_9649,N_9797);
nor U10422 (N_10422,N_9644,N_9056);
xor U10423 (N_10423,N_9948,N_9651);
nand U10424 (N_10424,N_9563,N_9982);
or U10425 (N_10425,N_9126,N_9275);
nor U10426 (N_10426,N_9315,N_9575);
or U10427 (N_10427,N_9794,N_9810);
xnor U10428 (N_10428,N_9124,N_9659);
or U10429 (N_10429,N_9119,N_9692);
nand U10430 (N_10430,N_9913,N_9876);
or U10431 (N_10431,N_9564,N_9731);
or U10432 (N_10432,N_9922,N_9169);
xor U10433 (N_10433,N_9451,N_9934);
or U10434 (N_10434,N_9802,N_9317);
nand U10435 (N_10435,N_9449,N_9770);
and U10436 (N_10436,N_9204,N_9039);
and U10437 (N_10437,N_9255,N_9211);
and U10438 (N_10438,N_9004,N_9737);
nor U10439 (N_10439,N_9684,N_9832);
and U10440 (N_10440,N_9672,N_9293);
nor U10441 (N_10441,N_9462,N_9329);
and U10442 (N_10442,N_9909,N_9607);
xnor U10443 (N_10443,N_9597,N_9945);
nand U10444 (N_10444,N_9130,N_9626);
xnor U10445 (N_10445,N_9184,N_9250);
nor U10446 (N_10446,N_9613,N_9015);
and U10447 (N_10447,N_9375,N_9152);
nor U10448 (N_10448,N_9953,N_9377);
or U10449 (N_10449,N_9252,N_9098);
xnor U10450 (N_10450,N_9941,N_9584);
xor U10451 (N_10451,N_9940,N_9879);
or U10452 (N_10452,N_9673,N_9667);
or U10453 (N_10453,N_9736,N_9972);
xnor U10454 (N_10454,N_9496,N_9699);
nand U10455 (N_10455,N_9572,N_9698);
and U10456 (N_10456,N_9836,N_9642);
xor U10457 (N_10457,N_9681,N_9643);
nor U10458 (N_10458,N_9481,N_9116);
xnor U10459 (N_10459,N_9869,N_9306);
nand U10460 (N_10460,N_9155,N_9277);
nand U10461 (N_10461,N_9839,N_9186);
xor U10462 (N_10462,N_9926,N_9360);
nor U10463 (N_10463,N_9814,N_9862);
and U10464 (N_10464,N_9193,N_9137);
nand U10465 (N_10465,N_9536,N_9716);
xnor U10466 (N_10466,N_9556,N_9418);
and U10467 (N_10467,N_9898,N_9529);
xnor U10468 (N_10468,N_9541,N_9601);
nand U10469 (N_10469,N_9166,N_9696);
nand U10470 (N_10470,N_9828,N_9046);
nor U10471 (N_10471,N_9243,N_9508);
and U10472 (N_10472,N_9886,N_9470);
and U10473 (N_10473,N_9028,N_9062);
nor U10474 (N_10474,N_9432,N_9339);
nor U10475 (N_10475,N_9985,N_9612);
and U10476 (N_10476,N_9609,N_9742);
nor U10477 (N_10477,N_9954,N_9485);
nand U10478 (N_10478,N_9061,N_9419);
nand U10479 (N_10479,N_9772,N_9843);
nand U10480 (N_10480,N_9213,N_9385);
or U10481 (N_10481,N_9188,N_9790);
nand U10482 (N_10482,N_9067,N_9043);
xor U10483 (N_10483,N_9436,N_9871);
nand U10484 (N_10484,N_9519,N_9791);
and U10485 (N_10485,N_9078,N_9639);
nand U10486 (N_10486,N_9182,N_9181);
xnor U10487 (N_10487,N_9652,N_9636);
nand U10488 (N_10488,N_9145,N_9749);
nand U10489 (N_10489,N_9348,N_9328);
nor U10490 (N_10490,N_9045,N_9324);
or U10491 (N_10491,N_9946,N_9217);
nand U10492 (N_10492,N_9515,N_9139);
or U10493 (N_10493,N_9773,N_9956);
and U10494 (N_10494,N_9928,N_9094);
and U10495 (N_10495,N_9894,N_9369);
and U10496 (N_10496,N_9292,N_9969);
xnor U10497 (N_10497,N_9236,N_9634);
or U10498 (N_10498,N_9407,N_9570);
nand U10499 (N_10499,N_9523,N_9726);
nand U10500 (N_10500,N_9223,N_9318);
nor U10501 (N_10501,N_9240,N_9966);
nor U10502 (N_10502,N_9392,N_9689);
nand U10503 (N_10503,N_9823,N_9971);
xnor U10504 (N_10504,N_9087,N_9230);
or U10505 (N_10505,N_9650,N_9223);
xor U10506 (N_10506,N_9728,N_9692);
or U10507 (N_10507,N_9724,N_9750);
xor U10508 (N_10508,N_9560,N_9290);
xor U10509 (N_10509,N_9594,N_9087);
nor U10510 (N_10510,N_9981,N_9948);
and U10511 (N_10511,N_9395,N_9790);
nor U10512 (N_10512,N_9135,N_9499);
or U10513 (N_10513,N_9119,N_9793);
and U10514 (N_10514,N_9207,N_9274);
or U10515 (N_10515,N_9716,N_9740);
or U10516 (N_10516,N_9200,N_9956);
xor U10517 (N_10517,N_9812,N_9089);
xnor U10518 (N_10518,N_9423,N_9388);
or U10519 (N_10519,N_9272,N_9114);
or U10520 (N_10520,N_9436,N_9617);
or U10521 (N_10521,N_9261,N_9529);
and U10522 (N_10522,N_9679,N_9063);
and U10523 (N_10523,N_9593,N_9969);
nor U10524 (N_10524,N_9203,N_9443);
nor U10525 (N_10525,N_9424,N_9781);
xnor U10526 (N_10526,N_9520,N_9954);
and U10527 (N_10527,N_9917,N_9455);
nand U10528 (N_10528,N_9092,N_9366);
and U10529 (N_10529,N_9096,N_9981);
and U10530 (N_10530,N_9582,N_9345);
xor U10531 (N_10531,N_9184,N_9878);
nand U10532 (N_10532,N_9345,N_9076);
xor U10533 (N_10533,N_9643,N_9923);
nand U10534 (N_10534,N_9670,N_9929);
and U10535 (N_10535,N_9742,N_9006);
xnor U10536 (N_10536,N_9322,N_9303);
nand U10537 (N_10537,N_9201,N_9760);
xnor U10538 (N_10538,N_9947,N_9895);
or U10539 (N_10539,N_9430,N_9530);
and U10540 (N_10540,N_9243,N_9881);
or U10541 (N_10541,N_9130,N_9934);
nand U10542 (N_10542,N_9920,N_9495);
xor U10543 (N_10543,N_9294,N_9893);
nand U10544 (N_10544,N_9602,N_9834);
xnor U10545 (N_10545,N_9248,N_9684);
nand U10546 (N_10546,N_9220,N_9640);
and U10547 (N_10547,N_9491,N_9850);
and U10548 (N_10548,N_9411,N_9787);
or U10549 (N_10549,N_9647,N_9474);
or U10550 (N_10550,N_9664,N_9908);
nand U10551 (N_10551,N_9322,N_9534);
or U10552 (N_10552,N_9271,N_9138);
nor U10553 (N_10553,N_9058,N_9205);
nand U10554 (N_10554,N_9810,N_9243);
and U10555 (N_10555,N_9566,N_9473);
xnor U10556 (N_10556,N_9657,N_9791);
or U10557 (N_10557,N_9640,N_9636);
nand U10558 (N_10558,N_9754,N_9261);
and U10559 (N_10559,N_9423,N_9536);
or U10560 (N_10560,N_9057,N_9548);
or U10561 (N_10561,N_9664,N_9185);
nor U10562 (N_10562,N_9273,N_9264);
xor U10563 (N_10563,N_9538,N_9954);
nand U10564 (N_10564,N_9161,N_9999);
xnor U10565 (N_10565,N_9458,N_9422);
and U10566 (N_10566,N_9216,N_9910);
xnor U10567 (N_10567,N_9742,N_9820);
nand U10568 (N_10568,N_9686,N_9828);
or U10569 (N_10569,N_9805,N_9620);
or U10570 (N_10570,N_9011,N_9891);
and U10571 (N_10571,N_9111,N_9598);
nand U10572 (N_10572,N_9013,N_9373);
or U10573 (N_10573,N_9133,N_9192);
and U10574 (N_10574,N_9232,N_9022);
nor U10575 (N_10575,N_9359,N_9429);
or U10576 (N_10576,N_9205,N_9954);
or U10577 (N_10577,N_9095,N_9144);
nand U10578 (N_10578,N_9248,N_9160);
xor U10579 (N_10579,N_9289,N_9521);
nand U10580 (N_10580,N_9461,N_9153);
nor U10581 (N_10581,N_9947,N_9001);
or U10582 (N_10582,N_9239,N_9505);
and U10583 (N_10583,N_9924,N_9555);
or U10584 (N_10584,N_9933,N_9139);
nor U10585 (N_10585,N_9405,N_9579);
or U10586 (N_10586,N_9885,N_9756);
or U10587 (N_10587,N_9308,N_9564);
xnor U10588 (N_10588,N_9806,N_9230);
and U10589 (N_10589,N_9179,N_9423);
nor U10590 (N_10590,N_9243,N_9229);
and U10591 (N_10591,N_9874,N_9659);
or U10592 (N_10592,N_9063,N_9696);
or U10593 (N_10593,N_9128,N_9591);
nor U10594 (N_10594,N_9183,N_9572);
xnor U10595 (N_10595,N_9259,N_9739);
nand U10596 (N_10596,N_9825,N_9705);
and U10597 (N_10597,N_9485,N_9219);
nand U10598 (N_10598,N_9043,N_9712);
nor U10599 (N_10599,N_9605,N_9203);
or U10600 (N_10600,N_9162,N_9971);
nor U10601 (N_10601,N_9607,N_9088);
and U10602 (N_10602,N_9855,N_9374);
nand U10603 (N_10603,N_9891,N_9721);
or U10604 (N_10604,N_9543,N_9443);
nor U10605 (N_10605,N_9765,N_9459);
and U10606 (N_10606,N_9070,N_9952);
nand U10607 (N_10607,N_9586,N_9740);
xnor U10608 (N_10608,N_9686,N_9428);
and U10609 (N_10609,N_9920,N_9926);
or U10610 (N_10610,N_9810,N_9854);
nand U10611 (N_10611,N_9418,N_9316);
nand U10612 (N_10612,N_9837,N_9375);
xnor U10613 (N_10613,N_9724,N_9950);
xnor U10614 (N_10614,N_9922,N_9981);
xor U10615 (N_10615,N_9741,N_9181);
xor U10616 (N_10616,N_9593,N_9863);
nor U10617 (N_10617,N_9164,N_9543);
and U10618 (N_10618,N_9880,N_9850);
nor U10619 (N_10619,N_9252,N_9118);
nor U10620 (N_10620,N_9475,N_9831);
or U10621 (N_10621,N_9404,N_9395);
nand U10622 (N_10622,N_9270,N_9108);
and U10623 (N_10623,N_9602,N_9561);
or U10624 (N_10624,N_9584,N_9339);
nand U10625 (N_10625,N_9616,N_9290);
nor U10626 (N_10626,N_9952,N_9908);
or U10627 (N_10627,N_9774,N_9482);
nand U10628 (N_10628,N_9324,N_9728);
or U10629 (N_10629,N_9333,N_9563);
nor U10630 (N_10630,N_9324,N_9826);
xnor U10631 (N_10631,N_9732,N_9750);
nand U10632 (N_10632,N_9209,N_9445);
or U10633 (N_10633,N_9745,N_9223);
nand U10634 (N_10634,N_9042,N_9022);
xor U10635 (N_10635,N_9257,N_9698);
and U10636 (N_10636,N_9316,N_9821);
nand U10637 (N_10637,N_9958,N_9000);
and U10638 (N_10638,N_9593,N_9835);
xor U10639 (N_10639,N_9408,N_9701);
and U10640 (N_10640,N_9033,N_9889);
and U10641 (N_10641,N_9182,N_9416);
or U10642 (N_10642,N_9339,N_9456);
xor U10643 (N_10643,N_9276,N_9144);
nand U10644 (N_10644,N_9034,N_9283);
xor U10645 (N_10645,N_9979,N_9178);
nand U10646 (N_10646,N_9318,N_9332);
xnor U10647 (N_10647,N_9610,N_9974);
xnor U10648 (N_10648,N_9725,N_9880);
and U10649 (N_10649,N_9607,N_9351);
nand U10650 (N_10650,N_9106,N_9745);
nor U10651 (N_10651,N_9554,N_9119);
or U10652 (N_10652,N_9490,N_9966);
or U10653 (N_10653,N_9860,N_9807);
or U10654 (N_10654,N_9159,N_9111);
and U10655 (N_10655,N_9113,N_9523);
and U10656 (N_10656,N_9525,N_9461);
xnor U10657 (N_10657,N_9896,N_9895);
and U10658 (N_10658,N_9132,N_9452);
and U10659 (N_10659,N_9024,N_9986);
nand U10660 (N_10660,N_9585,N_9793);
nor U10661 (N_10661,N_9663,N_9860);
and U10662 (N_10662,N_9534,N_9656);
nand U10663 (N_10663,N_9638,N_9156);
and U10664 (N_10664,N_9884,N_9494);
and U10665 (N_10665,N_9562,N_9632);
or U10666 (N_10666,N_9310,N_9789);
nand U10667 (N_10667,N_9223,N_9455);
xnor U10668 (N_10668,N_9385,N_9002);
nor U10669 (N_10669,N_9090,N_9440);
and U10670 (N_10670,N_9743,N_9281);
or U10671 (N_10671,N_9872,N_9340);
nor U10672 (N_10672,N_9168,N_9240);
nand U10673 (N_10673,N_9673,N_9804);
nand U10674 (N_10674,N_9928,N_9728);
nor U10675 (N_10675,N_9436,N_9227);
nand U10676 (N_10676,N_9009,N_9272);
nor U10677 (N_10677,N_9835,N_9032);
and U10678 (N_10678,N_9034,N_9740);
nor U10679 (N_10679,N_9609,N_9652);
and U10680 (N_10680,N_9762,N_9989);
or U10681 (N_10681,N_9408,N_9996);
nor U10682 (N_10682,N_9392,N_9700);
and U10683 (N_10683,N_9637,N_9518);
nand U10684 (N_10684,N_9224,N_9180);
xor U10685 (N_10685,N_9641,N_9056);
nand U10686 (N_10686,N_9079,N_9095);
xnor U10687 (N_10687,N_9224,N_9645);
nor U10688 (N_10688,N_9655,N_9391);
nor U10689 (N_10689,N_9936,N_9636);
nand U10690 (N_10690,N_9763,N_9336);
and U10691 (N_10691,N_9819,N_9696);
or U10692 (N_10692,N_9103,N_9256);
nor U10693 (N_10693,N_9528,N_9994);
nor U10694 (N_10694,N_9561,N_9810);
nor U10695 (N_10695,N_9674,N_9093);
nand U10696 (N_10696,N_9726,N_9599);
and U10697 (N_10697,N_9330,N_9685);
and U10698 (N_10698,N_9556,N_9764);
or U10699 (N_10699,N_9915,N_9533);
xor U10700 (N_10700,N_9209,N_9414);
and U10701 (N_10701,N_9323,N_9350);
and U10702 (N_10702,N_9922,N_9662);
or U10703 (N_10703,N_9350,N_9851);
and U10704 (N_10704,N_9849,N_9586);
and U10705 (N_10705,N_9568,N_9095);
nand U10706 (N_10706,N_9355,N_9410);
nand U10707 (N_10707,N_9735,N_9377);
nand U10708 (N_10708,N_9219,N_9390);
nor U10709 (N_10709,N_9475,N_9009);
xor U10710 (N_10710,N_9452,N_9886);
nor U10711 (N_10711,N_9464,N_9542);
and U10712 (N_10712,N_9530,N_9321);
xnor U10713 (N_10713,N_9316,N_9328);
nor U10714 (N_10714,N_9243,N_9893);
xor U10715 (N_10715,N_9407,N_9926);
nand U10716 (N_10716,N_9666,N_9552);
and U10717 (N_10717,N_9532,N_9448);
and U10718 (N_10718,N_9331,N_9498);
nor U10719 (N_10719,N_9729,N_9822);
xnor U10720 (N_10720,N_9637,N_9567);
and U10721 (N_10721,N_9489,N_9252);
nand U10722 (N_10722,N_9522,N_9857);
and U10723 (N_10723,N_9048,N_9495);
and U10724 (N_10724,N_9999,N_9692);
or U10725 (N_10725,N_9926,N_9901);
or U10726 (N_10726,N_9705,N_9029);
nor U10727 (N_10727,N_9421,N_9288);
nand U10728 (N_10728,N_9174,N_9221);
and U10729 (N_10729,N_9871,N_9968);
nor U10730 (N_10730,N_9075,N_9702);
nand U10731 (N_10731,N_9438,N_9903);
and U10732 (N_10732,N_9988,N_9778);
nor U10733 (N_10733,N_9579,N_9134);
xnor U10734 (N_10734,N_9006,N_9985);
nand U10735 (N_10735,N_9976,N_9503);
xor U10736 (N_10736,N_9327,N_9516);
nand U10737 (N_10737,N_9492,N_9991);
and U10738 (N_10738,N_9051,N_9867);
nand U10739 (N_10739,N_9773,N_9383);
or U10740 (N_10740,N_9720,N_9246);
xnor U10741 (N_10741,N_9568,N_9127);
nor U10742 (N_10742,N_9483,N_9247);
xor U10743 (N_10743,N_9674,N_9972);
and U10744 (N_10744,N_9935,N_9135);
xor U10745 (N_10745,N_9513,N_9329);
or U10746 (N_10746,N_9628,N_9003);
xnor U10747 (N_10747,N_9117,N_9873);
xor U10748 (N_10748,N_9519,N_9284);
or U10749 (N_10749,N_9565,N_9592);
and U10750 (N_10750,N_9981,N_9829);
nor U10751 (N_10751,N_9359,N_9233);
nand U10752 (N_10752,N_9459,N_9795);
or U10753 (N_10753,N_9325,N_9155);
nor U10754 (N_10754,N_9966,N_9649);
nor U10755 (N_10755,N_9797,N_9248);
and U10756 (N_10756,N_9746,N_9345);
and U10757 (N_10757,N_9189,N_9602);
and U10758 (N_10758,N_9977,N_9649);
or U10759 (N_10759,N_9245,N_9131);
and U10760 (N_10760,N_9442,N_9102);
xor U10761 (N_10761,N_9674,N_9592);
xor U10762 (N_10762,N_9119,N_9513);
nand U10763 (N_10763,N_9067,N_9806);
nor U10764 (N_10764,N_9181,N_9948);
xnor U10765 (N_10765,N_9153,N_9488);
or U10766 (N_10766,N_9592,N_9782);
and U10767 (N_10767,N_9176,N_9319);
or U10768 (N_10768,N_9186,N_9509);
nor U10769 (N_10769,N_9867,N_9055);
or U10770 (N_10770,N_9002,N_9057);
nor U10771 (N_10771,N_9783,N_9796);
xor U10772 (N_10772,N_9141,N_9280);
nor U10773 (N_10773,N_9340,N_9847);
or U10774 (N_10774,N_9825,N_9460);
xor U10775 (N_10775,N_9908,N_9553);
or U10776 (N_10776,N_9879,N_9113);
and U10777 (N_10777,N_9676,N_9337);
nand U10778 (N_10778,N_9614,N_9540);
xnor U10779 (N_10779,N_9542,N_9825);
or U10780 (N_10780,N_9959,N_9878);
xor U10781 (N_10781,N_9579,N_9816);
or U10782 (N_10782,N_9093,N_9071);
nor U10783 (N_10783,N_9736,N_9745);
xor U10784 (N_10784,N_9356,N_9953);
xnor U10785 (N_10785,N_9983,N_9081);
nor U10786 (N_10786,N_9412,N_9508);
and U10787 (N_10787,N_9053,N_9323);
nor U10788 (N_10788,N_9186,N_9755);
xor U10789 (N_10789,N_9196,N_9467);
and U10790 (N_10790,N_9993,N_9285);
or U10791 (N_10791,N_9984,N_9006);
xnor U10792 (N_10792,N_9008,N_9260);
xnor U10793 (N_10793,N_9178,N_9532);
or U10794 (N_10794,N_9753,N_9428);
nor U10795 (N_10795,N_9562,N_9885);
nand U10796 (N_10796,N_9801,N_9829);
or U10797 (N_10797,N_9750,N_9183);
nand U10798 (N_10798,N_9179,N_9061);
and U10799 (N_10799,N_9069,N_9000);
or U10800 (N_10800,N_9777,N_9467);
or U10801 (N_10801,N_9518,N_9016);
and U10802 (N_10802,N_9150,N_9793);
nand U10803 (N_10803,N_9077,N_9087);
nand U10804 (N_10804,N_9823,N_9975);
nor U10805 (N_10805,N_9333,N_9362);
xor U10806 (N_10806,N_9471,N_9611);
xor U10807 (N_10807,N_9895,N_9317);
or U10808 (N_10808,N_9105,N_9864);
nand U10809 (N_10809,N_9014,N_9521);
or U10810 (N_10810,N_9145,N_9177);
nand U10811 (N_10811,N_9415,N_9754);
nand U10812 (N_10812,N_9488,N_9008);
xor U10813 (N_10813,N_9275,N_9403);
nor U10814 (N_10814,N_9314,N_9509);
and U10815 (N_10815,N_9191,N_9113);
xnor U10816 (N_10816,N_9778,N_9421);
xnor U10817 (N_10817,N_9280,N_9610);
xor U10818 (N_10818,N_9589,N_9210);
xor U10819 (N_10819,N_9228,N_9718);
nor U10820 (N_10820,N_9456,N_9656);
xor U10821 (N_10821,N_9069,N_9858);
xnor U10822 (N_10822,N_9343,N_9339);
or U10823 (N_10823,N_9868,N_9136);
xnor U10824 (N_10824,N_9654,N_9293);
or U10825 (N_10825,N_9756,N_9915);
xnor U10826 (N_10826,N_9559,N_9425);
and U10827 (N_10827,N_9582,N_9226);
nor U10828 (N_10828,N_9892,N_9320);
nor U10829 (N_10829,N_9581,N_9792);
and U10830 (N_10830,N_9221,N_9241);
or U10831 (N_10831,N_9907,N_9660);
or U10832 (N_10832,N_9312,N_9144);
xnor U10833 (N_10833,N_9368,N_9311);
nand U10834 (N_10834,N_9785,N_9234);
nand U10835 (N_10835,N_9175,N_9032);
xnor U10836 (N_10836,N_9828,N_9727);
nand U10837 (N_10837,N_9745,N_9783);
or U10838 (N_10838,N_9686,N_9018);
xnor U10839 (N_10839,N_9443,N_9493);
and U10840 (N_10840,N_9309,N_9463);
or U10841 (N_10841,N_9523,N_9965);
nor U10842 (N_10842,N_9411,N_9687);
and U10843 (N_10843,N_9390,N_9156);
or U10844 (N_10844,N_9907,N_9255);
xor U10845 (N_10845,N_9784,N_9918);
xor U10846 (N_10846,N_9336,N_9166);
nor U10847 (N_10847,N_9718,N_9328);
or U10848 (N_10848,N_9983,N_9437);
or U10849 (N_10849,N_9998,N_9313);
xnor U10850 (N_10850,N_9958,N_9633);
nor U10851 (N_10851,N_9463,N_9607);
or U10852 (N_10852,N_9774,N_9928);
xnor U10853 (N_10853,N_9173,N_9799);
xor U10854 (N_10854,N_9174,N_9181);
xor U10855 (N_10855,N_9702,N_9078);
nand U10856 (N_10856,N_9219,N_9277);
and U10857 (N_10857,N_9265,N_9994);
nand U10858 (N_10858,N_9060,N_9070);
or U10859 (N_10859,N_9102,N_9824);
or U10860 (N_10860,N_9817,N_9289);
xor U10861 (N_10861,N_9547,N_9294);
and U10862 (N_10862,N_9027,N_9970);
and U10863 (N_10863,N_9838,N_9200);
nand U10864 (N_10864,N_9141,N_9317);
nor U10865 (N_10865,N_9020,N_9880);
xor U10866 (N_10866,N_9417,N_9239);
or U10867 (N_10867,N_9479,N_9642);
nor U10868 (N_10868,N_9235,N_9741);
xor U10869 (N_10869,N_9426,N_9070);
or U10870 (N_10870,N_9200,N_9742);
xnor U10871 (N_10871,N_9880,N_9166);
nor U10872 (N_10872,N_9613,N_9685);
nand U10873 (N_10873,N_9919,N_9208);
nor U10874 (N_10874,N_9387,N_9809);
or U10875 (N_10875,N_9056,N_9633);
and U10876 (N_10876,N_9885,N_9773);
or U10877 (N_10877,N_9029,N_9943);
nand U10878 (N_10878,N_9292,N_9127);
and U10879 (N_10879,N_9843,N_9357);
nor U10880 (N_10880,N_9270,N_9412);
nand U10881 (N_10881,N_9800,N_9003);
nor U10882 (N_10882,N_9710,N_9414);
or U10883 (N_10883,N_9666,N_9971);
nand U10884 (N_10884,N_9465,N_9016);
or U10885 (N_10885,N_9592,N_9512);
nand U10886 (N_10886,N_9160,N_9622);
nand U10887 (N_10887,N_9484,N_9548);
nand U10888 (N_10888,N_9914,N_9853);
xor U10889 (N_10889,N_9715,N_9882);
nand U10890 (N_10890,N_9038,N_9873);
or U10891 (N_10891,N_9425,N_9238);
nand U10892 (N_10892,N_9672,N_9283);
or U10893 (N_10893,N_9596,N_9394);
nand U10894 (N_10894,N_9053,N_9710);
or U10895 (N_10895,N_9826,N_9348);
xnor U10896 (N_10896,N_9576,N_9191);
and U10897 (N_10897,N_9085,N_9294);
or U10898 (N_10898,N_9701,N_9237);
nor U10899 (N_10899,N_9830,N_9755);
or U10900 (N_10900,N_9768,N_9051);
nor U10901 (N_10901,N_9996,N_9958);
nand U10902 (N_10902,N_9184,N_9571);
nor U10903 (N_10903,N_9689,N_9249);
or U10904 (N_10904,N_9774,N_9040);
nand U10905 (N_10905,N_9736,N_9773);
and U10906 (N_10906,N_9932,N_9965);
or U10907 (N_10907,N_9726,N_9313);
and U10908 (N_10908,N_9612,N_9077);
nor U10909 (N_10909,N_9947,N_9039);
and U10910 (N_10910,N_9518,N_9494);
nand U10911 (N_10911,N_9299,N_9913);
xnor U10912 (N_10912,N_9457,N_9450);
and U10913 (N_10913,N_9921,N_9505);
or U10914 (N_10914,N_9391,N_9950);
or U10915 (N_10915,N_9742,N_9304);
nor U10916 (N_10916,N_9966,N_9767);
xor U10917 (N_10917,N_9725,N_9062);
nor U10918 (N_10918,N_9133,N_9304);
or U10919 (N_10919,N_9863,N_9718);
and U10920 (N_10920,N_9717,N_9139);
xor U10921 (N_10921,N_9238,N_9427);
nand U10922 (N_10922,N_9781,N_9886);
nand U10923 (N_10923,N_9548,N_9309);
nand U10924 (N_10924,N_9671,N_9329);
nand U10925 (N_10925,N_9701,N_9647);
and U10926 (N_10926,N_9355,N_9731);
and U10927 (N_10927,N_9843,N_9808);
nor U10928 (N_10928,N_9063,N_9225);
xnor U10929 (N_10929,N_9942,N_9601);
or U10930 (N_10930,N_9736,N_9455);
xor U10931 (N_10931,N_9740,N_9552);
nand U10932 (N_10932,N_9918,N_9208);
nor U10933 (N_10933,N_9431,N_9203);
nor U10934 (N_10934,N_9341,N_9078);
nor U10935 (N_10935,N_9864,N_9469);
or U10936 (N_10936,N_9261,N_9522);
or U10937 (N_10937,N_9429,N_9220);
nor U10938 (N_10938,N_9561,N_9881);
xnor U10939 (N_10939,N_9917,N_9072);
and U10940 (N_10940,N_9191,N_9642);
or U10941 (N_10941,N_9644,N_9185);
nand U10942 (N_10942,N_9111,N_9744);
xnor U10943 (N_10943,N_9757,N_9880);
or U10944 (N_10944,N_9981,N_9108);
and U10945 (N_10945,N_9903,N_9203);
nand U10946 (N_10946,N_9247,N_9347);
nor U10947 (N_10947,N_9632,N_9034);
xor U10948 (N_10948,N_9730,N_9772);
nand U10949 (N_10949,N_9517,N_9866);
xor U10950 (N_10950,N_9230,N_9697);
nand U10951 (N_10951,N_9875,N_9607);
nor U10952 (N_10952,N_9114,N_9842);
xnor U10953 (N_10953,N_9418,N_9886);
or U10954 (N_10954,N_9129,N_9316);
nand U10955 (N_10955,N_9708,N_9550);
nand U10956 (N_10956,N_9373,N_9249);
and U10957 (N_10957,N_9502,N_9523);
xor U10958 (N_10958,N_9118,N_9412);
nand U10959 (N_10959,N_9402,N_9935);
and U10960 (N_10960,N_9469,N_9553);
or U10961 (N_10961,N_9411,N_9784);
and U10962 (N_10962,N_9453,N_9917);
or U10963 (N_10963,N_9472,N_9560);
or U10964 (N_10964,N_9374,N_9822);
or U10965 (N_10965,N_9787,N_9008);
or U10966 (N_10966,N_9422,N_9774);
xor U10967 (N_10967,N_9296,N_9725);
nand U10968 (N_10968,N_9393,N_9028);
nor U10969 (N_10969,N_9381,N_9638);
nand U10970 (N_10970,N_9742,N_9571);
or U10971 (N_10971,N_9261,N_9464);
xnor U10972 (N_10972,N_9502,N_9789);
nand U10973 (N_10973,N_9741,N_9126);
nor U10974 (N_10974,N_9052,N_9784);
nor U10975 (N_10975,N_9743,N_9634);
or U10976 (N_10976,N_9783,N_9687);
nand U10977 (N_10977,N_9434,N_9090);
and U10978 (N_10978,N_9680,N_9762);
or U10979 (N_10979,N_9748,N_9296);
or U10980 (N_10980,N_9617,N_9115);
nand U10981 (N_10981,N_9917,N_9728);
and U10982 (N_10982,N_9770,N_9012);
nor U10983 (N_10983,N_9829,N_9222);
nor U10984 (N_10984,N_9433,N_9108);
xnor U10985 (N_10985,N_9735,N_9981);
and U10986 (N_10986,N_9747,N_9946);
or U10987 (N_10987,N_9718,N_9286);
or U10988 (N_10988,N_9805,N_9100);
nand U10989 (N_10989,N_9935,N_9016);
nor U10990 (N_10990,N_9418,N_9564);
xnor U10991 (N_10991,N_9082,N_9709);
nor U10992 (N_10992,N_9295,N_9512);
nor U10993 (N_10993,N_9037,N_9737);
and U10994 (N_10994,N_9873,N_9851);
and U10995 (N_10995,N_9284,N_9999);
nand U10996 (N_10996,N_9873,N_9521);
nor U10997 (N_10997,N_9727,N_9108);
and U10998 (N_10998,N_9389,N_9910);
xnor U10999 (N_10999,N_9505,N_9967);
and U11000 (N_11000,N_10165,N_10535);
nor U11001 (N_11001,N_10602,N_10764);
nor U11002 (N_11002,N_10003,N_10903);
nand U11003 (N_11003,N_10448,N_10643);
nand U11004 (N_11004,N_10388,N_10335);
nor U11005 (N_11005,N_10005,N_10672);
and U11006 (N_11006,N_10073,N_10329);
nand U11007 (N_11007,N_10317,N_10596);
nor U11008 (N_11008,N_10196,N_10600);
and U11009 (N_11009,N_10563,N_10195);
nor U11010 (N_11010,N_10557,N_10298);
and U11011 (N_11011,N_10280,N_10931);
or U11012 (N_11012,N_10149,N_10978);
and U11013 (N_11013,N_10257,N_10450);
nor U11014 (N_11014,N_10034,N_10309);
nand U11015 (N_11015,N_10876,N_10191);
nand U11016 (N_11016,N_10033,N_10733);
and U11017 (N_11017,N_10731,N_10820);
or U11018 (N_11018,N_10341,N_10015);
and U11019 (N_11019,N_10251,N_10702);
xnor U11020 (N_11020,N_10669,N_10480);
nor U11021 (N_11021,N_10841,N_10118);
xor U11022 (N_11022,N_10908,N_10681);
or U11023 (N_11023,N_10741,N_10549);
or U11024 (N_11024,N_10048,N_10942);
or U11025 (N_11025,N_10293,N_10456);
xor U11026 (N_11026,N_10119,N_10113);
xor U11027 (N_11027,N_10246,N_10453);
and U11028 (N_11028,N_10881,N_10553);
or U11029 (N_11029,N_10849,N_10943);
nand U11030 (N_11030,N_10086,N_10355);
and U11031 (N_11031,N_10124,N_10805);
or U11032 (N_11032,N_10787,N_10188);
nand U11033 (N_11033,N_10577,N_10268);
nor U11034 (N_11034,N_10956,N_10834);
and U11035 (N_11035,N_10700,N_10387);
xnor U11036 (N_11036,N_10830,N_10499);
and U11037 (N_11037,N_10373,N_10862);
or U11038 (N_11038,N_10079,N_10590);
nor U11039 (N_11039,N_10366,N_10140);
and U11040 (N_11040,N_10069,N_10856);
nor U11041 (N_11041,N_10305,N_10888);
nor U11042 (N_11042,N_10239,N_10714);
nand U11043 (N_11043,N_10249,N_10502);
nand U11044 (N_11044,N_10259,N_10601);
xor U11045 (N_11045,N_10980,N_10695);
or U11046 (N_11046,N_10569,N_10458);
nor U11047 (N_11047,N_10482,N_10773);
and U11048 (N_11048,N_10099,N_10029);
and U11049 (N_11049,N_10804,N_10679);
xnor U11050 (N_11050,N_10904,N_10476);
nand U11051 (N_11051,N_10678,N_10272);
nand U11052 (N_11052,N_10997,N_10279);
and U11053 (N_11053,N_10248,N_10181);
nand U11054 (N_11054,N_10582,N_10220);
or U11055 (N_11055,N_10746,N_10004);
and U11056 (N_11056,N_10779,N_10639);
nand U11057 (N_11057,N_10545,N_10342);
and U11058 (N_11058,N_10505,N_10556);
nor U11059 (N_11059,N_10211,N_10288);
or U11060 (N_11060,N_10981,N_10972);
nor U11061 (N_11061,N_10433,N_10047);
or U11062 (N_11062,N_10863,N_10066);
nor U11063 (N_11063,N_10250,N_10411);
and U11064 (N_11064,N_10243,N_10708);
xor U11065 (N_11065,N_10656,N_10735);
nand U11066 (N_11066,N_10800,N_10889);
nor U11067 (N_11067,N_10906,N_10833);
or U11068 (N_11068,N_10712,N_10912);
nand U11069 (N_11069,N_10621,N_10114);
nand U11070 (N_11070,N_10706,N_10854);
or U11071 (N_11071,N_10893,N_10543);
and U11072 (N_11072,N_10444,N_10216);
xor U11073 (N_11073,N_10096,N_10595);
and U11074 (N_11074,N_10218,N_10056);
or U11075 (N_11075,N_10438,N_10281);
nand U11076 (N_11076,N_10348,N_10057);
nor U11077 (N_11077,N_10959,N_10691);
nand U11078 (N_11078,N_10657,N_10055);
nand U11079 (N_11079,N_10921,N_10913);
or U11080 (N_11080,N_10219,N_10996);
and U11081 (N_11081,N_10283,N_10848);
nand U11082 (N_11082,N_10423,N_10585);
nand U11083 (N_11083,N_10197,N_10562);
or U11084 (N_11084,N_10263,N_10721);
and U11085 (N_11085,N_10891,N_10137);
xor U11086 (N_11086,N_10973,N_10724);
or U11087 (N_11087,N_10227,N_10007);
and U11088 (N_11088,N_10175,N_10457);
or U11089 (N_11089,N_10103,N_10513);
nor U11090 (N_11090,N_10430,N_10950);
nand U11091 (N_11091,N_10240,N_10021);
nor U11092 (N_11092,N_10794,N_10937);
nand U11093 (N_11093,N_10770,N_10995);
or U11094 (N_11094,N_10353,N_10381);
nor U11095 (N_11095,N_10983,N_10971);
nand U11096 (N_11096,N_10238,N_10842);
or U11097 (N_11097,N_10707,N_10000);
or U11098 (N_11098,N_10870,N_10551);
nand U11099 (N_11099,N_10372,N_10190);
or U11100 (N_11100,N_10696,N_10436);
nor U11101 (N_11101,N_10327,N_10187);
nand U11102 (N_11102,N_10117,N_10910);
nand U11103 (N_11103,N_10151,N_10840);
nand U11104 (N_11104,N_10396,N_10132);
xnor U11105 (N_11105,N_10414,N_10415);
xor U11106 (N_11106,N_10336,N_10624);
and U11107 (N_11107,N_10442,N_10258);
xor U11108 (N_11108,N_10485,N_10736);
nor U11109 (N_11109,N_10075,N_10939);
xnor U11110 (N_11110,N_10088,N_10084);
nand U11111 (N_11111,N_10674,N_10801);
and U11112 (N_11112,N_10122,N_10198);
nor U11113 (N_11113,N_10019,N_10785);
nand U11114 (N_11114,N_10161,N_10732);
or U11115 (N_11115,N_10920,N_10107);
and U11116 (N_11116,N_10895,N_10362);
and U11117 (N_11117,N_10711,N_10429);
or U11118 (N_11118,N_10665,N_10166);
xor U11119 (N_11119,N_10659,N_10914);
nor U11120 (N_11120,N_10496,N_10509);
nand U11121 (N_11121,N_10559,N_10802);
nor U11122 (N_11122,N_10169,N_10441);
or U11123 (N_11123,N_10291,N_10857);
nand U11124 (N_11124,N_10953,N_10323);
and U11125 (N_11125,N_10526,N_10793);
xor U11126 (N_11126,N_10528,N_10072);
or U11127 (N_11127,N_10725,N_10233);
nand U11128 (N_11128,N_10338,N_10177);
xor U11129 (N_11129,N_10992,N_10874);
nor U11130 (N_11130,N_10717,N_10269);
nor U11131 (N_11131,N_10946,N_10286);
xnor U11132 (N_11132,N_10580,N_10466);
and U11133 (N_11133,N_10176,N_10858);
and U11134 (N_11134,N_10040,N_10765);
nor U11135 (N_11135,N_10811,N_10558);
nor U11136 (N_11136,N_10383,N_10748);
or U11137 (N_11137,N_10941,N_10809);
nor U11138 (N_11138,N_10852,N_10527);
nand U11139 (N_11139,N_10630,N_10352);
nand U11140 (N_11140,N_10028,N_10835);
nor U11141 (N_11141,N_10449,N_10924);
and U11142 (N_11142,N_10407,N_10470);
nand U11143 (N_11143,N_10092,N_10483);
nand U11144 (N_11144,N_10310,N_10018);
or U11145 (N_11145,N_10367,N_10247);
xor U11146 (N_11146,N_10264,N_10478);
nand U11147 (N_11147,N_10756,N_10202);
xnor U11148 (N_11148,N_10544,N_10306);
nand U11149 (N_11149,N_10928,N_10797);
or U11150 (N_11150,N_10186,N_10302);
or U11151 (N_11151,N_10587,N_10481);
nand U11152 (N_11152,N_10767,N_10803);
nor U11153 (N_11153,N_10668,N_10168);
or U11154 (N_11154,N_10548,N_10789);
and U11155 (N_11155,N_10667,N_10235);
nand U11156 (N_11156,N_10322,N_10518);
nor U11157 (N_11157,N_10012,N_10185);
nor U11158 (N_11158,N_10445,N_10212);
nor U11159 (N_11159,N_10333,N_10579);
or U11160 (N_11160,N_10345,N_10008);
nand U11161 (N_11161,N_10963,N_10892);
or U11162 (N_11162,N_10693,N_10147);
xnor U11163 (N_11163,N_10573,N_10699);
or U11164 (N_11164,N_10490,N_10230);
nand U11165 (N_11165,N_10087,N_10522);
or U11166 (N_11166,N_10964,N_10262);
or U11167 (N_11167,N_10357,N_10645);
nor U11168 (N_11168,N_10347,N_10022);
and U11169 (N_11169,N_10753,N_10917);
and U11170 (N_11170,N_10360,N_10395);
nand U11171 (N_11171,N_10215,N_10465);
or U11172 (N_11172,N_10821,N_10989);
and U11173 (N_11173,N_10455,N_10402);
nor U11174 (N_11174,N_10027,N_10815);
nand U11175 (N_11175,N_10823,N_10845);
nor U11176 (N_11176,N_10163,N_10990);
and U11177 (N_11177,N_10918,N_10783);
and U11178 (N_11178,N_10358,N_10726);
and U11179 (N_11179,N_10976,N_10653);
and U11180 (N_11180,N_10900,N_10617);
or U11181 (N_11181,N_10439,N_10564);
xor U11182 (N_11182,N_10651,N_10267);
xnor U11183 (N_11183,N_10515,N_10541);
or U11184 (N_11184,N_10546,N_10300);
nand U11185 (N_11185,N_10339,N_10214);
nor U11186 (N_11186,N_10615,N_10053);
nand U11187 (N_11187,N_10762,N_10153);
and U11188 (N_11188,N_10207,N_10299);
nand U11189 (N_11189,N_10713,N_10241);
xnor U11190 (N_11190,N_10328,N_10192);
or U11191 (N_11191,N_10504,N_10728);
xnor U11192 (N_11192,N_10330,N_10744);
and U11193 (N_11193,N_10390,N_10663);
nand U11194 (N_11194,N_10795,N_10616);
and U11195 (N_11195,N_10666,N_10266);
and U11196 (N_11196,N_10619,N_10560);
and U11197 (N_11197,N_10882,N_10897);
nand U11198 (N_11198,N_10193,N_10832);
and U11199 (N_11199,N_10957,N_10974);
nand U11200 (N_11200,N_10958,N_10567);
nor U11201 (N_11201,N_10319,N_10303);
or U11202 (N_11202,N_10688,N_10968);
xnor U11203 (N_11203,N_10135,N_10393);
or U11204 (N_11204,N_10627,N_10510);
nor U11205 (N_11205,N_10772,N_10098);
or U11206 (N_11206,N_10723,N_10822);
and U11207 (N_11207,N_10861,N_10816);
nor U11208 (N_11208,N_10568,N_10745);
and U11209 (N_11209,N_10460,N_10253);
and U11210 (N_11210,N_10799,N_10986);
xnor U11211 (N_11211,N_10575,N_10925);
or U11212 (N_11212,N_10182,N_10083);
nor U11213 (N_11213,N_10649,N_10947);
nor U11214 (N_11214,N_10002,N_10063);
nor U11215 (N_11215,N_10422,N_10884);
nand U11216 (N_11216,N_10231,N_10592);
nor U11217 (N_11217,N_10487,N_10189);
or U11218 (N_11218,N_10778,N_10419);
nor U11219 (N_11219,N_10781,N_10749);
and U11220 (N_11220,N_10539,N_10447);
xor U11221 (N_11221,N_10226,N_10818);
and U11222 (N_11222,N_10705,N_10593);
or U11223 (N_11223,N_10343,N_10529);
nand U11224 (N_11224,N_10375,N_10684);
xor U11225 (N_11225,N_10134,N_10059);
and U11226 (N_11226,N_10125,N_10637);
or U11227 (N_11227,N_10632,N_10318);
xnor U11228 (N_11228,N_10332,N_10346);
or U11229 (N_11229,N_10364,N_10780);
nor U11230 (N_11230,N_10911,N_10324);
and U11231 (N_11231,N_10452,N_10829);
nor U11232 (N_11232,N_10400,N_10727);
nand U11233 (N_11233,N_10013,N_10225);
or U11234 (N_11234,N_10493,N_10042);
or U11235 (N_11235,N_10065,N_10109);
and U11236 (N_11236,N_10256,N_10909);
nand U11237 (N_11237,N_10320,N_10853);
or U11238 (N_11238,N_10392,N_10289);
nor U11239 (N_11239,N_10127,N_10060);
nand U11240 (N_11240,N_10171,N_10474);
nand U11241 (N_11241,N_10363,N_10839);
nor U11242 (N_11242,N_10229,N_10044);
nand U11243 (N_11243,N_10960,N_10097);
and U11244 (N_11244,N_10111,N_10807);
nor U11245 (N_11245,N_10473,N_10877);
xor U11246 (N_11246,N_10650,N_10454);
xnor U11247 (N_11247,N_10277,N_10661);
xnor U11248 (N_11248,N_10150,N_10790);
or U11249 (N_11249,N_10254,N_10143);
xnor U11250 (N_11250,N_10867,N_10144);
xor U11251 (N_11251,N_10316,N_10993);
or U11252 (N_11252,N_10704,N_10041);
nor U11253 (N_11253,N_10697,N_10312);
xor U11254 (N_11254,N_10039,N_10091);
nand U11255 (N_11255,N_10782,N_10718);
or U11256 (N_11256,N_10110,N_10572);
or U11257 (N_11257,N_10275,N_10570);
xor U11258 (N_11258,N_10915,N_10424);
or U11259 (N_11259,N_10951,N_10106);
and U11260 (N_11260,N_10136,N_10294);
and U11261 (N_11261,N_10244,N_10301);
and U11262 (N_11262,N_10826,N_10652);
or U11263 (N_11263,N_10885,N_10866);
nor U11264 (N_11264,N_10497,N_10500);
and U11265 (N_11265,N_10164,N_10644);
xor U11266 (N_11266,N_10965,N_10133);
or U11267 (N_11267,N_10475,N_10070);
nand U11268 (N_11268,N_10094,N_10417);
xnor U11269 (N_11269,N_10922,N_10156);
and U11270 (N_11270,N_10880,N_10677);
or U11271 (N_11271,N_10359,N_10058);
xnor U11272 (N_11272,N_10896,N_10844);
nand U11273 (N_11273,N_10750,N_10524);
nor U11274 (N_11274,N_10507,N_10154);
or U11275 (N_11275,N_10203,N_10081);
nand U11276 (N_11276,N_10126,N_10213);
or U11277 (N_11277,N_10584,N_10610);
xor U11278 (N_11278,N_10670,N_10631);
xor U11279 (N_11279,N_10872,N_10488);
nor U11280 (N_11280,N_10371,N_10817);
or U11281 (N_11281,N_10308,N_10599);
nand U11282 (N_11282,N_10382,N_10720);
xor U11283 (N_11283,N_10537,N_10090);
and U11284 (N_11284,N_10418,N_10634);
and U11285 (N_11285,N_10228,N_10952);
nor U11286 (N_11286,N_10128,N_10855);
or U11287 (N_11287,N_10542,N_10222);
nor U11288 (N_11288,N_10581,N_10641);
xnor U11289 (N_11289,N_10934,N_10970);
and U11290 (N_11290,N_10686,N_10552);
nand U11291 (N_11291,N_10385,N_10451);
nand U11292 (N_11292,N_10949,N_10771);
nor U11293 (N_11293,N_10167,N_10123);
xor U11294 (N_11294,N_10217,N_10242);
xnor U11295 (N_11295,N_10080,N_10378);
xor U11296 (N_11296,N_10139,N_10221);
nand U11297 (N_11297,N_10759,N_10403);
or U11298 (N_11298,N_10533,N_10612);
or U11299 (N_11299,N_10998,N_10658);
or U11300 (N_11300,N_10479,N_10204);
nand U11301 (N_11301,N_10729,N_10273);
nor U11302 (N_11302,N_10032,N_10016);
xnor U11303 (N_11303,N_10089,N_10991);
xor U11304 (N_11304,N_10873,N_10287);
xnor U11305 (N_11305,N_10969,N_10443);
and U11306 (N_11306,N_10682,N_10685);
and U11307 (N_11307,N_10907,N_10886);
nor U11308 (N_11308,N_10337,N_10565);
nor U11309 (N_11309,N_10174,N_10927);
and U11310 (N_11310,N_10102,N_10623);
or U11311 (N_11311,N_10232,N_10523);
nand U11312 (N_11312,N_10586,N_10977);
and U11313 (N_11313,N_10709,N_10825);
xnor U11314 (N_11314,N_10796,N_10916);
nand U11315 (N_11315,N_10890,N_10923);
or U11316 (N_11316,N_10605,N_10270);
nand U11317 (N_11317,N_10408,N_10571);
and U11318 (N_11318,N_10369,N_10798);
xnor U11319 (N_11319,N_10664,N_10967);
and U11320 (N_11320,N_10416,N_10010);
xor U11321 (N_11321,N_10112,N_10325);
nand U11322 (N_11322,N_10680,N_10660);
and U11323 (N_11323,N_10437,N_10598);
and U11324 (N_11324,N_10142,N_10374);
nor U11325 (N_11325,N_10101,N_10766);
nor U11326 (N_11326,N_10503,N_10351);
xnor U11327 (N_11327,N_10052,N_10626);
and U11328 (N_11328,N_10646,N_10394);
nand U11329 (N_11329,N_10105,N_10608);
nor U11330 (N_11330,N_10859,N_10905);
nor U11331 (N_11331,N_10494,N_10550);
nor U11332 (N_11332,N_10607,N_10078);
and U11333 (N_11333,N_10183,N_10935);
and U11334 (N_11334,N_10271,N_10391);
nand U11335 (N_11335,N_10987,N_10954);
nor U11336 (N_11336,N_10030,N_10994);
or U11337 (N_11337,N_10206,N_10932);
nor U11338 (N_11338,N_10531,N_10426);
or U11339 (N_11339,N_10389,N_10314);
and U11340 (N_11340,N_10326,N_10847);
or U11341 (N_11341,N_10498,N_10810);
nor U11342 (N_11342,N_10647,N_10440);
or U11343 (N_11343,N_10376,N_10609);
nor U11344 (N_11344,N_10331,N_10236);
or U11345 (N_11345,N_10566,N_10878);
xor U11346 (N_11346,N_10349,N_10690);
or U11347 (N_11347,N_10199,N_10739);
or U11348 (N_11348,N_10521,N_10082);
nand U11349 (N_11349,N_10014,N_10938);
nand U11350 (N_11350,N_10701,N_10827);
xor U11351 (N_11351,N_10622,N_10945);
or U11352 (N_11352,N_10129,N_10633);
and U11353 (N_11353,N_10282,N_10648);
nor U11354 (N_11354,N_10869,N_10525);
nand U11355 (N_11355,N_10901,N_10121);
and U11356 (N_11356,N_10074,N_10285);
nor U11357 (N_11357,N_10636,N_10763);
nor U11358 (N_11358,N_10520,N_10988);
nand U11359 (N_11359,N_10806,N_10758);
or U11360 (N_11360,N_10208,N_10296);
xor U11361 (N_11361,N_10412,N_10062);
and U11362 (N_11362,N_10006,N_10514);
nor U11363 (N_11363,N_10141,N_10170);
nor U11364 (N_11364,N_10620,N_10757);
nand U11365 (N_11365,N_10640,N_10824);
or U11366 (N_11366,N_10671,N_10477);
nand U11367 (N_11367,N_10591,N_10675);
or U11368 (N_11368,N_10694,N_10734);
xor U11369 (N_11369,N_10583,N_10768);
or U11370 (N_11370,N_10962,N_10252);
nor U11371 (N_11371,N_10597,N_10162);
and U11372 (N_11372,N_10940,N_10274);
or U11373 (N_11373,N_10077,N_10589);
and U11374 (N_11374,N_10031,N_10157);
xor U11375 (N_11375,N_10155,N_10410);
xnor U11376 (N_11376,N_10145,N_10606);
nor U11377 (N_11377,N_10929,N_10061);
xor U11378 (N_11378,N_10838,N_10464);
or U11379 (N_11379,N_10100,N_10009);
xor U11380 (N_11380,N_10011,N_10446);
xor U11381 (N_11381,N_10613,N_10205);
nor U11382 (N_11382,N_10740,N_10655);
and U11383 (N_11383,N_10472,N_10761);
xnor U11384 (N_11384,N_10982,N_10344);
nor U11385 (N_11385,N_10836,N_10754);
nor U11386 (N_11386,N_10260,N_10340);
and U11387 (N_11387,N_10026,N_10370);
or U11388 (N_11388,N_10898,N_10290);
or U11389 (N_11389,N_10777,N_10201);
nor U11390 (N_11390,N_10051,N_10628);
xor U11391 (N_11391,N_10828,N_10561);
and U11392 (N_11392,N_10130,N_10755);
nor U11393 (N_11393,N_10819,N_10315);
and U11394 (N_11394,N_10933,N_10519);
nand U11395 (N_11395,N_10049,N_10875);
nor U11396 (N_11396,N_10791,N_10846);
xor U11397 (N_11397,N_10307,N_10085);
nor U11398 (N_11398,N_10409,N_10108);
nand U11399 (N_11399,N_10698,N_10471);
or U11400 (N_11400,N_10948,N_10462);
xnor U11401 (N_11401,N_10413,N_10261);
nand U11402 (N_11402,N_10899,N_10304);
nor U11403 (N_11403,N_10463,N_10554);
and U11404 (N_11404,N_10116,N_10966);
xnor U11405 (N_11405,N_10334,N_10361);
nor U11406 (N_11406,N_10851,N_10692);
or U11407 (N_11407,N_10883,N_10160);
nor U11408 (N_11408,N_10625,N_10321);
and U11409 (N_11409,N_10401,N_10831);
and U11410 (N_11410,N_10313,N_10689);
and U11411 (N_11411,N_10534,N_10420);
nand U11412 (N_11412,N_10431,N_10276);
xor U11413 (N_11413,N_10435,N_10377);
nand U11414 (N_11414,N_10104,N_10071);
or U11415 (N_11415,N_10354,N_10769);
nand U11416 (N_11416,N_10210,N_10045);
or U11417 (N_11417,N_10486,N_10588);
nor U11418 (N_11418,N_10237,N_10278);
xnor U11419 (N_11419,N_10719,N_10574);
nor U11420 (N_11420,N_10638,N_10295);
nor U11421 (N_11421,N_10432,N_10635);
nand U11422 (N_11422,N_10629,N_10985);
and U11423 (N_11423,N_10979,N_10035);
xor U11424 (N_11424,N_10025,N_10611);
and U11425 (N_11425,N_10642,N_10023);
nor U11426 (N_11426,N_10747,N_10148);
and U11427 (N_11427,N_10930,N_10038);
nand U11428 (N_11428,N_10428,N_10265);
and U11429 (N_11429,N_10865,N_10489);
nand U11430 (N_11430,N_10173,N_10555);
or U11431 (N_11431,N_10730,N_10434);
and U11432 (N_11432,N_10926,N_10676);
or U11433 (N_11433,N_10501,N_10200);
xnor U11434 (N_11434,N_10506,N_10530);
nand U11435 (N_11435,N_10540,N_10397);
xnor U11436 (N_11436,N_10095,N_10813);
and U11437 (N_11437,N_10703,N_10037);
nor U11438 (N_11438,N_10120,N_10814);
xor U11439 (N_11439,N_10380,N_10398);
xor U11440 (N_11440,N_10495,N_10517);
nor U11441 (N_11441,N_10001,N_10784);
nand U11442 (N_11442,N_10512,N_10860);
or U11443 (N_11443,N_10999,N_10158);
nand U11444 (N_11444,N_10752,N_10716);
or U11445 (N_11445,N_10297,N_10245);
xnor U11446 (N_11446,N_10654,N_10404);
xnor U11447 (N_11447,N_10365,N_10255);
nor U11448 (N_11448,N_10683,N_10975);
nor U11449 (N_11449,N_10837,N_10224);
and U11450 (N_11450,N_10152,N_10738);
and U11451 (N_11451,N_10068,N_10508);
or U11452 (N_11452,N_10868,N_10020);
nor U11453 (N_11453,N_10751,N_10843);
xnor U11454 (N_11454,N_10050,N_10054);
and U11455 (N_11455,N_10209,N_10776);
nand U11456 (N_11456,N_10491,N_10194);
or U11457 (N_11457,N_10076,N_10808);
nor U11458 (N_11458,N_10722,N_10469);
nor U11459 (N_11459,N_10384,N_10046);
and U11460 (N_11460,N_10604,N_10944);
nor U11461 (N_11461,N_10792,N_10406);
nor U11462 (N_11462,N_10603,N_10662);
or U11463 (N_11463,N_10064,N_10710);
or U11464 (N_11464,N_10687,N_10775);
or U11465 (N_11465,N_10368,N_10871);
or U11466 (N_11466,N_10036,N_10379);
xnor U11467 (N_11467,N_10234,N_10024);
xor U11468 (N_11468,N_10594,N_10421);
nand U11469 (N_11469,N_10715,N_10138);
xnor U11470 (N_11470,N_10737,N_10427);
nand U11471 (N_11471,N_10984,N_10578);
nor U11472 (N_11472,N_10532,N_10284);
nor U11473 (N_11473,N_10180,N_10484);
or U11474 (N_11474,N_10468,N_10405);
xnor U11475 (N_11475,N_10356,N_10673);
and U11476 (N_11476,N_10516,N_10311);
nand U11477 (N_11477,N_10894,N_10350);
nand U11478 (N_11478,N_10399,N_10179);
or U11479 (N_11479,N_10093,N_10461);
and U11480 (N_11480,N_10223,N_10760);
nand U11481 (N_11481,N_10538,N_10774);
and U11482 (N_11482,N_10614,N_10425);
nand U11483 (N_11483,N_10864,N_10887);
or U11484 (N_11484,N_10492,N_10146);
nand U11485 (N_11485,N_10812,N_10902);
xor U11486 (N_11486,N_10743,N_10017);
or U11487 (N_11487,N_10955,N_10459);
nand U11488 (N_11488,N_10536,N_10879);
nand U11489 (N_11489,N_10386,N_10511);
nor U11490 (N_11490,N_10184,N_10178);
nand U11491 (N_11491,N_10547,N_10850);
xnor U11492 (N_11492,N_10131,N_10961);
or U11493 (N_11493,N_10936,N_10618);
nand U11494 (N_11494,N_10786,N_10788);
nand U11495 (N_11495,N_10115,N_10576);
and U11496 (N_11496,N_10159,N_10919);
nand U11497 (N_11497,N_10292,N_10467);
xnor U11498 (N_11498,N_10067,N_10172);
nand U11499 (N_11499,N_10742,N_10043);
xor U11500 (N_11500,N_10599,N_10354);
and U11501 (N_11501,N_10950,N_10676);
nand U11502 (N_11502,N_10422,N_10974);
and U11503 (N_11503,N_10545,N_10582);
nand U11504 (N_11504,N_10211,N_10524);
nor U11505 (N_11505,N_10959,N_10660);
xor U11506 (N_11506,N_10624,N_10652);
nand U11507 (N_11507,N_10719,N_10939);
or U11508 (N_11508,N_10286,N_10244);
xor U11509 (N_11509,N_10734,N_10013);
nor U11510 (N_11510,N_10546,N_10370);
or U11511 (N_11511,N_10970,N_10000);
nand U11512 (N_11512,N_10468,N_10346);
and U11513 (N_11513,N_10162,N_10552);
nor U11514 (N_11514,N_10541,N_10855);
or U11515 (N_11515,N_10970,N_10391);
nand U11516 (N_11516,N_10882,N_10994);
xnor U11517 (N_11517,N_10332,N_10749);
or U11518 (N_11518,N_10436,N_10290);
or U11519 (N_11519,N_10624,N_10339);
or U11520 (N_11520,N_10245,N_10480);
nor U11521 (N_11521,N_10790,N_10934);
xor U11522 (N_11522,N_10378,N_10348);
and U11523 (N_11523,N_10699,N_10507);
xnor U11524 (N_11524,N_10915,N_10979);
or U11525 (N_11525,N_10621,N_10063);
nor U11526 (N_11526,N_10916,N_10222);
nand U11527 (N_11527,N_10716,N_10131);
or U11528 (N_11528,N_10582,N_10728);
or U11529 (N_11529,N_10910,N_10577);
nor U11530 (N_11530,N_10346,N_10582);
and U11531 (N_11531,N_10498,N_10991);
xnor U11532 (N_11532,N_10696,N_10234);
and U11533 (N_11533,N_10941,N_10471);
nor U11534 (N_11534,N_10439,N_10018);
or U11535 (N_11535,N_10814,N_10589);
nor U11536 (N_11536,N_10708,N_10522);
and U11537 (N_11537,N_10350,N_10383);
and U11538 (N_11538,N_10539,N_10114);
xnor U11539 (N_11539,N_10159,N_10905);
and U11540 (N_11540,N_10478,N_10915);
or U11541 (N_11541,N_10660,N_10731);
and U11542 (N_11542,N_10926,N_10028);
and U11543 (N_11543,N_10069,N_10714);
xnor U11544 (N_11544,N_10512,N_10967);
and U11545 (N_11545,N_10371,N_10080);
and U11546 (N_11546,N_10740,N_10659);
or U11547 (N_11547,N_10306,N_10078);
and U11548 (N_11548,N_10295,N_10068);
nand U11549 (N_11549,N_10746,N_10522);
nor U11550 (N_11550,N_10315,N_10001);
xor U11551 (N_11551,N_10960,N_10940);
and U11552 (N_11552,N_10285,N_10836);
nor U11553 (N_11553,N_10550,N_10653);
or U11554 (N_11554,N_10988,N_10125);
nor U11555 (N_11555,N_10799,N_10166);
and U11556 (N_11556,N_10436,N_10376);
xnor U11557 (N_11557,N_10153,N_10268);
and U11558 (N_11558,N_10353,N_10841);
xnor U11559 (N_11559,N_10814,N_10276);
nor U11560 (N_11560,N_10196,N_10418);
and U11561 (N_11561,N_10144,N_10417);
or U11562 (N_11562,N_10534,N_10174);
xor U11563 (N_11563,N_10054,N_10491);
and U11564 (N_11564,N_10186,N_10069);
nor U11565 (N_11565,N_10303,N_10839);
xnor U11566 (N_11566,N_10175,N_10858);
or U11567 (N_11567,N_10116,N_10226);
nor U11568 (N_11568,N_10506,N_10667);
xor U11569 (N_11569,N_10312,N_10798);
nand U11570 (N_11570,N_10966,N_10233);
nor U11571 (N_11571,N_10974,N_10519);
xor U11572 (N_11572,N_10842,N_10778);
and U11573 (N_11573,N_10308,N_10922);
nand U11574 (N_11574,N_10728,N_10934);
xnor U11575 (N_11575,N_10060,N_10933);
and U11576 (N_11576,N_10989,N_10666);
nor U11577 (N_11577,N_10108,N_10450);
xor U11578 (N_11578,N_10487,N_10003);
or U11579 (N_11579,N_10145,N_10493);
xor U11580 (N_11580,N_10975,N_10525);
nand U11581 (N_11581,N_10920,N_10616);
nor U11582 (N_11582,N_10317,N_10407);
nand U11583 (N_11583,N_10588,N_10697);
xnor U11584 (N_11584,N_10610,N_10236);
nor U11585 (N_11585,N_10104,N_10504);
xnor U11586 (N_11586,N_10596,N_10422);
nor U11587 (N_11587,N_10987,N_10414);
or U11588 (N_11588,N_10919,N_10441);
nor U11589 (N_11589,N_10399,N_10329);
nor U11590 (N_11590,N_10580,N_10219);
nor U11591 (N_11591,N_10193,N_10002);
xor U11592 (N_11592,N_10447,N_10330);
xor U11593 (N_11593,N_10903,N_10759);
nand U11594 (N_11594,N_10444,N_10015);
xor U11595 (N_11595,N_10615,N_10039);
nor U11596 (N_11596,N_10226,N_10550);
nand U11597 (N_11597,N_10014,N_10423);
xnor U11598 (N_11598,N_10915,N_10295);
and U11599 (N_11599,N_10003,N_10793);
nor U11600 (N_11600,N_10841,N_10287);
and U11601 (N_11601,N_10154,N_10714);
and U11602 (N_11602,N_10057,N_10637);
and U11603 (N_11603,N_10904,N_10009);
and U11604 (N_11604,N_10895,N_10643);
nor U11605 (N_11605,N_10257,N_10356);
nand U11606 (N_11606,N_10242,N_10661);
nor U11607 (N_11607,N_10778,N_10213);
xnor U11608 (N_11608,N_10852,N_10229);
xor U11609 (N_11609,N_10836,N_10488);
or U11610 (N_11610,N_10414,N_10200);
or U11611 (N_11611,N_10409,N_10076);
nor U11612 (N_11612,N_10307,N_10679);
or U11613 (N_11613,N_10875,N_10237);
nand U11614 (N_11614,N_10210,N_10178);
and U11615 (N_11615,N_10462,N_10192);
nand U11616 (N_11616,N_10070,N_10756);
or U11617 (N_11617,N_10263,N_10684);
xnor U11618 (N_11618,N_10412,N_10620);
xnor U11619 (N_11619,N_10744,N_10022);
and U11620 (N_11620,N_10601,N_10862);
or U11621 (N_11621,N_10634,N_10969);
and U11622 (N_11622,N_10602,N_10340);
and U11623 (N_11623,N_10885,N_10249);
or U11624 (N_11624,N_10026,N_10263);
nand U11625 (N_11625,N_10613,N_10696);
nor U11626 (N_11626,N_10346,N_10140);
or U11627 (N_11627,N_10453,N_10828);
or U11628 (N_11628,N_10457,N_10701);
xnor U11629 (N_11629,N_10821,N_10203);
xnor U11630 (N_11630,N_10427,N_10364);
or U11631 (N_11631,N_10994,N_10327);
and U11632 (N_11632,N_10242,N_10214);
xnor U11633 (N_11633,N_10938,N_10370);
nand U11634 (N_11634,N_10243,N_10082);
nor U11635 (N_11635,N_10423,N_10187);
and U11636 (N_11636,N_10155,N_10306);
and U11637 (N_11637,N_10391,N_10971);
xnor U11638 (N_11638,N_10589,N_10849);
nor U11639 (N_11639,N_10565,N_10487);
or U11640 (N_11640,N_10395,N_10143);
nor U11641 (N_11641,N_10885,N_10523);
nand U11642 (N_11642,N_10164,N_10315);
xnor U11643 (N_11643,N_10269,N_10291);
or U11644 (N_11644,N_10040,N_10970);
or U11645 (N_11645,N_10850,N_10857);
xnor U11646 (N_11646,N_10481,N_10332);
nor U11647 (N_11647,N_10107,N_10214);
nor U11648 (N_11648,N_10823,N_10095);
nor U11649 (N_11649,N_10062,N_10028);
nor U11650 (N_11650,N_10211,N_10098);
nor U11651 (N_11651,N_10802,N_10255);
nor U11652 (N_11652,N_10719,N_10163);
nand U11653 (N_11653,N_10360,N_10692);
or U11654 (N_11654,N_10067,N_10796);
or U11655 (N_11655,N_10366,N_10288);
and U11656 (N_11656,N_10116,N_10237);
nand U11657 (N_11657,N_10980,N_10510);
nand U11658 (N_11658,N_10268,N_10355);
xor U11659 (N_11659,N_10084,N_10808);
nand U11660 (N_11660,N_10441,N_10879);
and U11661 (N_11661,N_10554,N_10549);
nand U11662 (N_11662,N_10059,N_10029);
nand U11663 (N_11663,N_10171,N_10991);
and U11664 (N_11664,N_10676,N_10235);
or U11665 (N_11665,N_10013,N_10712);
nor U11666 (N_11666,N_10443,N_10580);
and U11667 (N_11667,N_10056,N_10909);
xor U11668 (N_11668,N_10955,N_10104);
nand U11669 (N_11669,N_10621,N_10513);
nand U11670 (N_11670,N_10048,N_10631);
nand U11671 (N_11671,N_10011,N_10018);
xnor U11672 (N_11672,N_10925,N_10758);
xor U11673 (N_11673,N_10129,N_10451);
and U11674 (N_11674,N_10919,N_10632);
nor U11675 (N_11675,N_10686,N_10114);
and U11676 (N_11676,N_10625,N_10035);
nor U11677 (N_11677,N_10830,N_10417);
nor U11678 (N_11678,N_10780,N_10209);
nor U11679 (N_11679,N_10237,N_10646);
nand U11680 (N_11680,N_10702,N_10630);
and U11681 (N_11681,N_10212,N_10914);
xor U11682 (N_11682,N_10151,N_10314);
and U11683 (N_11683,N_10856,N_10773);
nand U11684 (N_11684,N_10042,N_10445);
nor U11685 (N_11685,N_10123,N_10085);
or U11686 (N_11686,N_10705,N_10706);
and U11687 (N_11687,N_10129,N_10037);
nor U11688 (N_11688,N_10399,N_10316);
or U11689 (N_11689,N_10419,N_10796);
nand U11690 (N_11690,N_10128,N_10281);
xor U11691 (N_11691,N_10508,N_10938);
or U11692 (N_11692,N_10803,N_10495);
or U11693 (N_11693,N_10751,N_10136);
xnor U11694 (N_11694,N_10618,N_10734);
nand U11695 (N_11695,N_10603,N_10793);
nor U11696 (N_11696,N_10138,N_10207);
and U11697 (N_11697,N_10600,N_10016);
or U11698 (N_11698,N_10430,N_10345);
nand U11699 (N_11699,N_10490,N_10120);
xor U11700 (N_11700,N_10026,N_10874);
nand U11701 (N_11701,N_10215,N_10943);
xor U11702 (N_11702,N_10820,N_10895);
or U11703 (N_11703,N_10390,N_10004);
or U11704 (N_11704,N_10317,N_10760);
nor U11705 (N_11705,N_10699,N_10394);
and U11706 (N_11706,N_10042,N_10661);
or U11707 (N_11707,N_10924,N_10448);
xor U11708 (N_11708,N_10521,N_10395);
nand U11709 (N_11709,N_10154,N_10089);
or U11710 (N_11710,N_10233,N_10870);
or U11711 (N_11711,N_10811,N_10509);
xor U11712 (N_11712,N_10370,N_10131);
nor U11713 (N_11713,N_10127,N_10491);
or U11714 (N_11714,N_10109,N_10487);
and U11715 (N_11715,N_10256,N_10650);
xor U11716 (N_11716,N_10486,N_10401);
xnor U11717 (N_11717,N_10773,N_10334);
nand U11718 (N_11718,N_10652,N_10761);
and U11719 (N_11719,N_10579,N_10624);
nor U11720 (N_11720,N_10458,N_10095);
nor U11721 (N_11721,N_10503,N_10657);
and U11722 (N_11722,N_10928,N_10234);
nand U11723 (N_11723,N_10276,N_10703);
nand U11724 (N_11724,N_10664,N_10446);
nor U11725 (N_11725,N_10365,N_10107);
xor U11726 (N_11726,N_10072,N_10521);
and U11727 (N_11727,N_10762,N_10550);
nand U11728 (N_11728,N_10309,N_10360);
and U11729 (N_11729,N_10884,N_10385);
xor U11730 (N_11730,N_10545,N_10965);
and U11731 (N_11731,N_10613,N_10253);
xor U11732 (N_11732,N_10030,N_10226);
or U11733 (N_11733,N_10718,N_10692);
or U11734 (N_11734,N_10149,N_10503);
and U11735 (N_11735,N_10447,N_10243);
xnor U11736 (N_11736,N_10832,N_10553);
and U11737 (N_11737,N_10650,N_10652);
and U11738 (N_11738,N_10493,N_10469);
or U11739 (N_11739,N_10949,N_10408);
nand U11740 (N_11740,N_10738,N_10388);
or U11741 (N_11741,N_10370,N_10442);
nand U11742 (N_11742,N_10833,N_10209);
xor U11743 (N_11743,N_10630,N_10347);
or U11744 (N_11744,N_10862,N_10726);
or U11745 (N_11745,N_10680,N_10892);
nand U11746 (N_11746,N_10790,N_10159);
nand U11747 (N_11747,N_10362,N_10466);
or U11748 (N_11748,N_10163,N_10026);
nand U11749 (N_11749,N_10325,N_10308);
nor U11750 (N_11750,N_10789,N_10426);
nand U11751 (N_11751,N_10516,N_10650);
nor U11752 (N_11752,N_10058,N_10675);
nor U11753 (N_11753,N_10883,N_10111);
nor U11754 (N_11754,N_10551,N_10411);
xnor U11755 (N_11755,N_10499,N_10752);
and U11756 (N_11756,N_10807,N_10508);
nand U11757 (N_11757,N_10487,N_10375);
nand U11758 (N_11758,N_10806,N_10179);
nand U11759 (N_11759,N_10673,N_10466);
xnor U11760 (N_11760,N_10923,N_10311);
or U11761 (N_11761,N_10004,N_10045);
and U11762 (N_11762,N_10730,N_10729);
nand U11763 (N_11763,N_10964,N_10898);
and U11764 (N_11764,N_10258,N_10938);
and U11765 (N_11765,N_10235,N_10006);
xnor U11766 (N_11766,N_10348,N_10186);
and U11767 (N_11767,N_10424,N_10960);
nand U11768 (N_11768,N_10445,N_10466);
nand U11769 (N_11769,N_10872,N_10353);
or U11770 (N_11770,N_10859,N_10922);
or U11771 (N_11771,N_10258,N_10612);
or U11772 (N_11772,N_10943,N_10315);
nand U11773 (N_11773,N_10287,N_10372);
nor U11774 (N_11774,N_10733,N_10551);
xnor U11775 (N_11775,N_10242,N_10578);
xnor U11776 (N_11776,N_10500,N_10125);
xor U11777 (N_11777,N_10737,N_10043);
and U11778 (N_11778,N_10412,N_10455);
nor U11779 (N_11779,N_10871,N_10551);
nand U11780 (N_11780,N_10908,N_10261);
and U11781 (N_11781,N_10508,N_10426);
nor U11782 (N_11782,N_10852,N_10790);
nand U11783 (N_11783,N_10239,N_10558);
nor U11784 (N_11784,N_10694,N_10871);
nor U11785 (N_11785,N_10254,N_10599);
xnor U11786 (N_11786,N_10162,N_10608);
xnor U11787 (N_11787,N_10791,N_10933);
and U11788 (N_11788,N_10732,N_10459);
nand U11789 (N_11789,N_10452,N_10413);
or U11790 (N_11790,N_10636,N_10422);
and U11791 (N_11791,N_10955,N_10166);
and U11792 (N_11792,N_10060,N_10984);
xnor U11793 (N_11793,N_10155,N_10138);
nand U11794 (N_11794,N_10847,N_10396);
xor U11795 (N_11795,N_10451,N_10838);
nand U11796 (N_11796,N_10917,N_10769);
nor U11797 (N_11797,N_10126,N_10999);
or U11798 (N_11798,N_10476,N_10392);
or U11799 (N_11799,N_10783,N_10834);
or U11800 (N_11800,N_10671,N_10300);
or U11801 (N_11801,N_10714,N_10640);
and U11802 (N_11802,N_10038,N_10419);
xnor U11803 (N_11803,N_10562,N_10563);
xor U11804 (N_11804,N_10022,N_10395);
xor U11805 (N_11805,N_10704,N_10805);
nor U11806 (N_11806,N_10806,N_10081);
and U11807 (N_11807,N_10862,N_10651);
and U11808 (N_11808,N_10048,N_10341);
and U11809 (N_11809,N_10290,N_10783);
xnor U11810 (N_11810,N_10767,N_10829);
or U11811 (N_11811,N_10948,N_10717);
xnor U11812 (N_11812,N_10863,N_10300);
nor U11813 (N_11813,N_10036,N_10213);
xor U11814 (N_11814,N_10745,N_10108);
xor U11815 (N_11815,N_10535,N_10823);
nand U11816 (N_11816,N_10302,N_10261);
xnor U11817 (N_11817,N_10780,N_10184);
xnor U11818 (N_11818,N_10315,N_10324);
xor U11819 (N_11819,N_10400,N_10186);
nand U11820 (N_11820,N_10132,N_10458);
xnor U11821 (N_11821,N_10116,N_10921);
xor U11822 (N_11822,N_10553,N_10129);
nand U11823 (N_11823,N_10206,N_10315);
nand U11824 (N_11824,N_10842,N_10769);
and U11825 (N_11825,N_10354,N_10343);
nor U11826 (N_11826,N_10333,N_10814);
xor U11827 (N_11827,N_10096,N_10365);
xor U11828 (N_11828,N_10001,N_10245);
nand U11829 (N_11829,N_10656,N_10232);
nor U11830 (N_11830,N_10760,N_10728);
and U11831 (N_11831,N_10675,N_10666);
nor U11832 (N_11832,N_10638,N_10089);
nand U11833 (N_11833,N_10630,N_10525);
nand U11834 (N_11834,N_10312,N_10439);
xor U11835 (N_11835,N_10127,N_10293);
or U11836 (N_11836,N_10713,N_10643);
xor U11837 (N_11837,N_10706,N_10991);
nand U11838 (N_11838,N_10842,N_10817);
or U11839 (N_11839,N_10542,N_10948);
nor U11840 (N_11840,N_10961,N_10814);
or U11841 (N_11841,N_10427,N_10940);
xnor U11842 (N_11842,N_10097,N_10062);
nand U11843 (N_11843,N_10775,N_10330);
nand U11844 (N_11844,N_10850,N_10167);
nand U11845 (N_11845,N_10970,N_10962);
nand U11846 (N_11846,N_10105,N_10131);
nor U11847 (N_11847,N_10319,N_10450);
nand U11848 (N_11848,N_10740,N_10410);
nand U11849 (N_11849,N_10253,N_10892);
and U11850 (N_11850,N_10967,N_10424);
or U11851 (N_11851,N_10327,N_10046);
nand U11852 (N_11852,N_10975,N_10419);
and U11853 (N_11853,N_10104,N_10777);
and U11854 (N_11854,N_10522,N_10782);
nor U11855 (N_11855,N_10291,N_10546);
nand U11856 (N_11856,N_10208,N_10889);
and U11857 (N_11857,N_10997,N_10444);
nand U11858 (N_11858,N_10933,N_10900);
nand U11859 (N_11859,N_10017,N_10175);
nor U11860 (N_11860,N_10848,N_10924);
and U11861 (N_11861,N_10371,N_10884);
and U11862 (N_11862,N_10023,N_10228);
or U11863 (N_11863,N_10750,N_10497);
and U11864 (N_11864,N_10397,N_10531);
or U11865 (N_11865,N_10820,N_10586);
nand U11866 (N_11866,N_10890,N_10379);
nand U11867 (N_11867,N_10119,N_10553);
nand U11868 (N_11868,N_10574,N_10161);
nor U11869 (N_11869,N_10849,N_10040);
xor U11870 (N_11870,N_10397,N_10891);
xor U11871 (N_11871,N_10290,N_10534);
or U11872 (N_11872,N_10031,N_10867);
nand U11873 (N_11873,N_10341,N_10186);
nand U11874 (N_11874,N_10480,N_10966);
nor U11875 (N_11875,N_10598,N_10699);
and U11876 (N_11876,N_10127,N_10465);
nor U11877 (N_11877,N_10497,N_10175);
and U11878 (N_11878,N_10574,N_10500);
or U11879 (N_11879,N_10056,N_10907);
nand U11880 (N_11880,N_10113,N_10593);
xnor U11881 (N_11881,N_10179,N_10069);
nor U11882 (N_11882,N_10519,N_10382);
nand U11883 (N_11883,N_10427,N_10587);
and U11884 (N_11884,N_10129,N_10371);
nor U11885 (N_11885,N_10744,N_10211);
nor U11886 (N_11886,N_10560,N_10545);
or U11887 (N_11887,N_10203,N_10695);
xnor U11888 (N_11888,N_10192,N_10794);
and U11889 (N_11889,N_10502,N_10072);
xnor U11890 (N_11890,N_10786,N_10076);
nor U11891 (N_11891,N_10324,N_10595);
nor U11892 (N_11892,N_10192,N_10150);
nor U11893 (N_11893,N_10979,N_10091);
nor U11894 (N_11894,N_10721,N_10449);
or U11895 (N_11895,N_10255,N_10994);
and U11896 (N_11896,N_10160,N_10336);
or U11897 (N_11897,N_10745,N_10965);
and U11898 (N_11898,N_10983,N_10818);
xnor U11899 (N_11899,N_10715,N_10574);
nand U11900 (N_11900,N_10039,N_10348);
xor U11901 (N_11901,N_10055,N_10969);
nor U11902 (N_11902,N_10120,N_10517);
and U11903 (N_11903,N_10894,N_10475);
xnor U11904 (N_11904,N_10753,N_10203);
xor U11905 (N_11905,N_10249,N_10550);
nor U11906 (N_11906,N_10031,N_10439);
nand U11907 (N_11907,N_10818,N_10290);
or U11908 (N_11908,N_10597,N_10237);
xnor U11909 (N_11909,N_10845,N_10495);
nor U11910 (N_11910,N_10588,N_10105);
or U11911 (N_11911,N_10387,N_10310);
nor U11912 (N_11912,N_10477,N_10418);
nor U11913 (N_11913,N_10842,N_10532);
nor U11914 (N_11914,N_10452,N_10403);
nor U11915 (N_11915,N_10413,N_10900);
and U11916 (N_11916,N_10851,N_10447);
nor U11917 (N_11917,N_10535,N_10689);
nor U11918 (N_11918,N_10378,N_10595);
and U11919 (N_11919,N_10199,N_10426);
and U11920 (N_11920,N_10120,N_10067);
or U11921 (N_11921,N_10971,N_10652);
nor U11922 (N_11922,N_10073,N_10480);
nor U11923 (N_11923,N_10481,N_10590);
nor U11924 (N_11924,N_10737,N_10927);
and U11925 (N_11925,N_10992,N_10543);
and U11926 (N_11926,N_10220,N_10195);
nand U11927 (N_11927,N_10094,N_10680);
xor U11928 (N_11928,N_10674,N_10851);
nand U11929 (N_11929,N_10679,N_10125);
or U11930 (N_11930,N_10307,N_10351);
and U11931 (N_11931,N_10454,N_10611);
and U11932 (N_11932,N_10431,N_10103);
nor U11933 (N_11933,N_10776,N_10569);
nand U11934 (N_11934,N_10370,N_10307);
nor U11935 (N_11935,N_10620,N_10869);
xnor U11936 (N_11936,N_10140,N_10332);
or U11937 (N_11937,N_10835,N_10619);
nand U11938 (N_11938,N_10946,N_10154);
and U11939 (N_11939,N_10442,N_10588);
and U11940 (N_11940,N_10479,N_10794);
or U11941 (N_11941,N_10562,N_10940);
nand U11942 (N_11942,N_10765,N_10984);
nand U11943 (N_11943,N_10547,N_10562);
and U11944 (N_11944,N_10071,N_10807);
nor U11945 (N_11945,N_10003,N_10225);
or U11946 (N_11946,N_10560,N_10154);
nor U11947 (N_11947,N_10944,N_10453);
and U11948 (N_11948,N_10944,N_10073);
and U11949 (N_11949,N_10128,N_10771);
nor U11950 (N_11950,N_10588,N_10426);
and U11951 (N_11951,N_10493,N_10955);
nand U11952 (N_11952,N_10079,N_10510);
nand U11953 (N_11953,N_10674,N_10737);
and U11954 (N_11954,N_10599,N_10826);
or U11955 (N_11955,N_10611,N_10640);
nand U11956 (N_11956,N_10640,N_10656);
xor U11957 (N_11957,N_10627,N_10029);
nand U11958 (N_11958,N_10013,N_10755);
nand U11959 (N_11959,N_10512,N_10568);
xnor U11960 (N_11960,N_10619,N_10469);
nand U11961 (N_11961,N_10914,N_10263);
nor U11962 (N_11962,N_10173,N_10823);
xnor U11963 (N_11963,N_10945,N_10217);
nor U11964 (N_11964,N_10980,N_10668);
nand U11965 (N_11965,N_10533,N_10282);
nor U11966 (N_11966,N_10274,N_10152);
or U11967 (N_11967,N_10310,N_10844);
or U11968 (N_11968,N_10333,N_10344);
or U11969 (N_11969,N_10829,N_10874);
xnor U11970 (N_11970,N_10898,N_10839);
nand U11971 (N_11971,N_10831,N_10219);
xnor U11972 (N_11972,N_10045,N_10461);
or U11973 (N_11973,N_10255,N_10266);
nor U11974 (N_11974,N_10791,N_10833);
nor U11975 (N_11975,N_10469,N_10136);
nor U11976 (N_11976,N_10499,N_10771);
and U11977 (N_11977,N_10121,N_10628);
and U11978 (N_11978,N_10594,N_10514);
or U11979 (N_11979,N_10570,N_10003);
nor U11980 (N_11980,N_10752,N_10973);
nor U11981 (N_11981,N_10424,N_10617);
or U11982 (N_11982,N_10110,N_10075);
and U11983 (N_11983,N_10299,N_10615);
xor U11984 (N_11984,N_10103,N_10340);
xnor U11985 (N_11985,N_10431,N_10936);
and U11986 (N_11986,N_10641,N_10063);
nor U11987 (N_11987,N_10261,N_10385);
nor U11988 (N_11988,N_10103,N_10559);
and U11989 (N_11989,N_10093,N_10525);
and U11990 (N_11990,N_10474,N_10389);
or U11991 (N_11991,N_10353,N_10820);
and U11992 (N_11992,N_10318,N_10715);
nand U11993 (N_11993,N_10928,N_10745);
nand U11994 (N_11994,N_10498,N_10554);
and U11995 (N_11995,N_10082,N_10959);
or U11996 (N_11996,N_10824,N_10886);
xor U11997 (N_11997,N_10115,N_10754);
and U11998 (N_11998,N_10099,N_10160);
xor U11999 (N_11999,N_10054,N_10929);
xnor U12000 (N_12000,N_11904,N_11957);
nor U12001 (N_12001,N_11881,N_11022);
and U12002 (N_12002,N_11706,N_11730);
and U12003 (N_12003,N_11675,N_11654);
nor U12004 (N_12004,N_11603,N_11921);
nand U12005 (N_12005,N_11451,N_11703);
and U12006 (N_12006,N_11089,N_11508);
nor U12007 (N_12007,N_11587,N_11344);
xor U12008 (N_12008,N_11059,N_11004);
or U12009 (N_12009,N_11725,N_11506);
or U12010 (N_12010,N_11563,N_11140);
and U12011 (N_12011,N_11607,N_11191);
nor U12012 (N_12012,N_11003,N_11822);
or U12013 (N_12013,N_11204,N_11057);
and U12014 (N_12014,N_11320,N_11115);
or U12015 (N_12015,N_11394,N_11181);
xnor U12016 (N_12016,N_11061,N_11544);
or U12017 (N_12017,N_11727,N_11783);
xor U12018 (N_12018,N_11826,N_11509);
or U12019 (N_12019,N_11153,N_11653);
nand U12020 (N_12020,N_11933,N_11348);
xor U12021 (N_12021,N_11273,N_11880);
nand U12022 (N_12022,N_11321,N_11310);
nor U12023 (N_12023,N_11131,N_11757);
or U12024 (N_12024,N_11923,N_11533);
or U12025 (N_12025,N_11298,N_11839);
nand U12026 (N_12026,N_11358,N_11854);
or U12027 (N_12027,N_11700,N_11389);
nor U12028 (N_12028,N_11135,N_11821);
and U12029 (N_12029,N_11091,N_11866);
nand U12030 (N_12030,N_11044,N_11278);
xor U12031 (N_12031,N_11827,N_11522);
xnor U12032 (N_12032,N_11788,N_11773);
and U12033 (N_12033,N_11211,N_11376);
nor U12034 (N_12034,N_11173,N_11023);
or U12035 (N_12035,N_11926,N_11980);
nor U12036 (N_12036,N_11184,N_11843);
nor U12037 (N_12037,N_11097,N_11805);
xnor U12038 (N_12038,N_11218,N_11391);
nand U12039 (N_12039,N_11373,N_11058);
and U12040 (N_12040,N_11951,N_11034);
and U12041 (N_12041,N_11581,N_11311);
nor U12042 (N_12042,N_11152,N_11400);
and U12043 (N_12043,N_11448,N_11415);
and U12044 (N_12044,N_11909,N_11802);
and U12045 (N_12045,N_11914,N_11844);
nor U12046 (N_12046,N_11610,N_11285);
nor U12047 (N_12047,N_11535,N_11574);
or U12048 (N_12048,N_11417,N_11196);
nor U12049 (N_12049,N_11493,N_11227);
nand U12050 (N_12050,N_11225,N_11998);
or U12051 (N_12051,N_11371,N_11553);
xor U12052 (N_12052,N_11812,N_11685);
or U12053 (N_12053,N_11962,N_11717);
nor U12054 (N_12054,N_11289,N_11069);
xnor U12055 (N_12055,N_11288,N_11944);
or U12056 (N_12056,N_11476,N_11531);
xnor U12057 (N_12057,N_11918,N_11324);
xor U12058 (N_12058,N_11720,N_11546);
xnor U12059 (N_12059,N_11609,N_11659);
or U12060 (N_12060,N_11830,N_11224);
nor U12061 (N_12061,N_11965,N_11862);
nand U12062 (N_12062,N_11429,N_11616);
nor U12063 (N_12063,N_11838,N_11269);
and U12064 (N_12064,N_11316,N_11172);
xor U12065 (N_12065,N_11635,N_11449);
or U12066 (N_12066,N_11092,N_11375);
nor U12067 (N_12067,N_11083,N_11006);
nand U12068 (N_12068,N_11698,N_11354);
nor U12069 (N_12069,N_11947,N_11431);
or U12070 (N_12070,N_11591,N_11833);
and U12071 (N_12071,N_11967,N_11814);
and U12072 (N_12072,N_11657,N_11895);
or U12073 (N_12073,N_11979,N_11537);
and U12074 (N_12074,N_11467,N_11643);
and U12075 (N_12075,N_11193,N_11859);
nor U12076 (N_12076,N_11699,N_11768);
nor U12077 (N_12077,N_11786,N_11398);
nand U12078 (N_12078,N_11548,N_11987);
nand U12079 (N_12079,N_11636,N_11108);
nand U12080 (N_12080,N_11529,N_11223);
nand U12081 (N_12081,N_11236,N_11632);
nor U12082 (N_12082,N_11887,N_11744);
and U12083 (N_12083,N_11575,N_11337);
nand U12084 (N_12084,N_11586,N_11490);
or U12085 (N_12085,N_11021,N_11498);
nand U12086 (N_12086,N_11105,N_11286);
xor U12087 (N_12087,N_11060,N_11229);
nand U12088 (N_12088,N_11713,N_11627);
nand U12089 (N_12089,N_11972,N_11035);
nor U12090 (N_12090,N_11145,N_11040);
or U12091 (N_12091,N_11526,N_11365);
xor U12092 (N_12092,N_11828,N_11290);
xnor U12093 (N_12093,N_11284,N_11538);
or U12094 (N_12094,N_11195,N_11599);
nand U12095 (N_12095,N_11729,N_11680);
xnor U12096 (N_12096,N_11272,N_11855);
or U12097 (N_12097,N_11074,N_11455);
nor U12098 (N_12098,N_11569,N_11712);
nand U12099 (N_12099,N_11361,N_11882);
and U12100 (N_12100,N_11129,N_11048);
nor U12101 (N_12101,N_11495,N_11112);
xnor U12102 (N_12102,N_11463,N_11994);
and U12103 (N_12103,N_11403,N_11641);
xnor U12104 (N_12104,N_11602,N_11510);
or U12105 (N_12105,N_11953,N_11169);
nor U12106 (N_12106,N_11910,N_11249);
xor U12107 (N_12107,N_11749,N_11670);
and U12108 (N_12108,N_11428,N_11435);
nand U12109 (N_12109,N_11939,N_11948);
nor U12110 (N_12110,N_11160,N_11010);
and U12111 (N_12111,N_11125,N_11268);
and U12112 (N_12112,N_11293,N_11307);
nor U12113 (N_12113,N_11488,N_11343);
nor U12114 (N_12114,N_11751,N_11017);
and U12115 (N_12115,N_11379,N_11634);
nand U12116 (N_12116,N_11138,N_11836);
nand U12117 (N_12117,N_11494,N_11246);
or U12118 (N_12118,N_11663,N_11304);
and U12119 (N_12119,N_11582,N_11327);
xor U12120 (N_12120,N_11710,N_11103);
or U12121 (N_12121,N_11033,N_11254);
nor U12122 (N_12122,N_11955,N_11232);
nand U12123 (N_12123,N_11850,N_11540);
or U12124 (N_12124,N_11666,N_11432);
nand U12125 (N_12125,N_11928,N_11758);
xor U12126 (N_12126,N_11804,N_11792);
nand U12127 (N_12127,N_11157,N_11491);
xor U12128 (N_12128,N_11925,N_11356);
nand U12129 (N_12129,N_11256,N_11199);
nor U12130 (N_12130,N_11963,N_11355);
nand U12131 (N_12131,N_11752,N_11385);
and U12132 (N_12132,N_11917,N_11203);
nor U12133 (N_12133,N_11228,N_11848);
nand U12134 (N_12134,N_11572,N_11560);
or U12135 (N_12135,N_11566,N_11088);
or U12136 (N_12136,N_11071,N_11949);
xnor U12137 (N_12137,N_11772,N_11280);
and U12138 (N_12138,N_11077,N_11978);
and U12139 (N_12139,N_11565,N_11576);
and U12140 (N_12140,N_11913,N_11894);
and U12141 (N_12141,N_11990,N_11483);
nor U12142 (N_12142,N_11890,N_11983);
and U12143 (N_12143,N_11942,N_11420);
nand U12144 (N_12144,N_11043,N_11469);
nand U12145 (N_12145,N_11513,N_11511);
or U12146 (N_12146,N_11200,N_11002);
and U12147 (N_12147,N_11601,N_11167);
nor U12148 (N_12148,N_11604,N_11845);
xor U12149 (N_12149,N_11276,N_11724);
xor U12150 (N_12150,N_11339,N_11111);
xnor U12151 (N_12151,N_11456,N_11785);
and U12152 (N_12152,N_11381,N_11208);
nor U12153 (N_12153,N_11096,N_11564);
or U12154 (N_12154,N_11243,N_11263);
xnor U12155 (N_12155,N_11387,N_11704);
nor U12156 (N_12156,N_11642,N_11212);
nor U12157 (N_12157,N_11613,N_11350);
nand U12158 (N_12158,N_11555,N_11693);
and U12159 (N_12159,N_11308,N_11931);
and U12160 (N_12160,N_11534,N_11958);
nor U12161 (N_12161,N_11150,N_11718);
nand U12162 (N_12162,N_11611,N_11815);
or U12163 (N_12163,N_11527,N_11501);
or U12164 (N_12164,N_11924,N_11440);
and U12165 (N_12165,N_11341,N_11771);
or U12166 (N_12166,N_11745,N_11045);
or U12167 (N_12167,N_11027,N_11852);
nand U12168 (N_12168,N_11128,N_11794);
nand U12169 (N_12169,N_11168,N_11543);
nor U12170 (N_12170,N_11347,N_11774);
nand U12171 (N_12171,N_11639,N_11452);
or U12172 (N_12172,N_11072,N_11335);
and U12173 (N_12173,N_11334,N_11776);
and U12174 (N_12174,N_11110,N_11971);
nor U12175 (N_12175,N_11433,N_11831);
nor U12176 (N_12176,N_11738,N_11661);
nand U12177 (N_12177,N_11446,N_11364);
nand U12178 (N_12178,N_11662,N_11479);
nor U12179 (N_12179,N_11192,N_11179);
nand U12180 (N_12180,N_11550,N_11976);
or U12181 (N_12181,N_11580,N_11408);
and U12182 (N_12182,N_11665,N_11049);
nand U12183 (N_12183,N_11042,N_11719);
and U12184 (N_12184,N_11419,N_11331);
nor U12185 (N_12185,N_11098,N_11041);
nor U12186 (N_12186,N_11888,N_11655);
nor U12187 (N_12187,N_11360,N_11697);
xnor U12188 (N_12188,N_11711,N_11902);
or U12189 (N_12189,N_11791,N_11899);
nand U12190 (N_12190,N_11945,N_11250);
xor U12191 (N_12191,N_11143,N_11161);
and U12192 (N_12192,N_11399,N_11528);
and U12193 (N_12193,N_11127,N_11282);
xor U12194 (N_12194,N_11743,N_11595);
and U12195 (N_12195,N_11158,N_11062);
nand U12196 (N_12196,N_11742,N_11038);
nor U12197 (N_12197,N_11996,N_11251);
nor U12198 (N_12198,N_11608,N_11715);
or U12199 (N_12199,N_11545,N_11741);
nor U12200 (N_12200,N_11001,N_11472);
nand U12201 (N_12201,N_11934,N_11916);
and U12202 (N_12202,N_11294,N_11064);
nor U12203 (N_12203,N_11695,N_11261);
xor U12204 (N_12204,N_11146,N_11504);
or U12205 (N_12205,N_11221,N_11906);
and U12206 (N_12206,N_11012,N_11935);
nand U12207 (N_12207,N_11011,N_11633);
xor U12208 (N_12208,N_11851,N_11780);
nand U12209 (N_12209,N_11974,N_11075);
nand U12210 (N_12210,N_11739,N_11301);
or U12211 (N_12211,N_11305,N_11877);
nand U12212 (N_12212,N_11405,N_11952);
xor U12213 (N_12213,N_11919,N_11484);
nand U12214 (N_12214,N_11325,N_11824);
nand U12215 (N_12215,N_11026,N_11300);
or U12216 (N_12216,N_11518,N_11406);
nor U12217 (N_12217,N_11692,N_11648);
or U12218 (N_12218,N_11466,N_11872);
nand U12219 (N_12219,N_11702,N_11503);
nor U12220 (N_12220,N_11922,N_11619);
and U12221 (N_12221,N_11318,N_11541);
and U12222 (N_12222,N_11076,N_11136);
nor U12223 (N_12223,N_11194,N_11297);
nand U12224 (N_12224,N_11829,N_11082);
or U12225 (N_12225,N_11502,N_11482);
nor U12226 (N_12226,N_11592,N_11559);
nor U12227 (N_12227,N_11411,N_11800);
and U12228 (N_12228,N_11823,N_11891);
xor U12229 (N_12229,N_11690,N_11015);
and U12230 (N_12230,N_11521,N_11209);
or U12231 (N_12231,N_11789,N_11000);
xnor U12232 (N_12232,N_11622,N_11864);
nand U12233 (N_12233,N_11468,N_11927);
xnor U12234 (N_12234,N_11068,N_11940);
and U12235 (N_12235,N_11287,N_11257);
xor U12236 (N_12236,N_11686,N_11631);
xnor U12237 (N_12237,N_11231,N_11312);
nor U12238 (N_12238,N_11803,N_11733);
xnor U12239 (N_12239,N_11763,N_11073);
or U12240 (N_12240,N_11530,N_11264);
and U12241 (N_12241,N_11445,N_11556);
or U12242 (N_12242,N_11860,N_11409);
nor U12243 (N_12243,N_11943,N_11233);
xor U12244 (N_12244,N_11107,N_11929);
and U12245 (N_12245,N_11995,N_11628);
nor U12246 (N_12246,N_11999,N_11645);
xnor U12247 (N_12247,N_11517,N_11746);
nor U12248 (N_12248,N_11677,N_11853);
xnor U12249 (N_12249,N_11694,N_11968);
nor U12250 (N_12250,N_11121,N_11147);
or U12251 (N_12251,N_11245,N_11753);
or U12252 (N_12252,N_11081,N_11732);
nor U12253 (N_12253,N_11497,N_11395);
and U12254 (N_12254,N_11322,N_11593);
or U12255 (N_12255,N_11104,N_11903);
and U12256 (N_12256,N_11606,N_11879);
and U12257 (N_12257,N_11215,N_11539);
nand U12258 (N_12258,N_11116,N_11039);
and U12259 (N_12259,N_11801,N_11422);
nand U12260 (N_12260,N_11915,N_11182);
nor U12261 (N_12261,N_11007,N_11667);
and U12262 (N_12262,N_11647,N_11051);
nand U12263 (N_12263,N_11874,N_11018);
nor U12264 (N_12264,N_11120,N_11876);
or U12265 (N_12265,N_11013,N_11137);
xor U12266 (N_12266,N_11477,N_11410);
xnor U12267 (N_12267,N_11180,N_11835);
nor U12268 (N_12268,N_11134,N_11912);
and U12269 (N_12269,N_11937,N_11333);
nor U12270 (N_12270,N_11795,N_11177);
nand U12271 (N_12271,N_11867,N_11683);
or U12272 (N_12272,N_11554,N_11977);
xor U12273 (N_12273,N_11857,N_11016);
or U12274 (N_12274,N_11736,N_11352);
xnor U12275 (N_12275,N_11470,N_11597);
and U12276 (N_12276,N_11418,N_11148);
nand U12277 (N_12277,N_11412,N_11779);
or U12278 (N_12278,N_11676,N_11106);
xnor U12279 (N_12279,N_11817,N_11840);
nor U12280 (N_12280,N_11067,N_11054);
nor U12281 (N_12281,N_11651,N_11434);
or U12282 (N_12282,N_11590,N_11464);
xor U12283 (N_12283,N_11809,N_11551);
and U12284 (N_12284,N_11542,N_11270);
or U12285 (N_12285,N_11781,N_11640);
xnor U12286 (N_12286,N_11100,N_11142);
nor U12287 (N_12287,N_11413,N_11870);
nand U12288 (N_12288,N_11426,N_11512);
xor U12289 (N_12289,N_11873,N_11793);
or U12290 (N_12290,N_11079,N_11485);
nor U12291 (N_12291,N_11423,N_11578);
or U12292 (N_12292,N_11799,N_11349);
nand U12293 (N_12293,N_11846,N_11709);
nand U12294 (N_12294,N_11295,N_11638);
or U12295 (N_12295,N_11317,N_11367);
xor U12296 (N_12296,N_11883,N_11296);
xnor U12297 (N_12297,N_11784,N_11032);
and U12298 (N_12298,N_11213,N_11900);
nor U12299 (N_12299,N_11357,N_11154);
xnor U12300 (N_12300,N_11388,N_11244);
or U12301 (N_12301,N_11570,N_11523);
and U12302 (N_12302,N_11637,N_11187);
xnor U12303 (N_12303,N_11624,N_11271);
and U12304 (N_12304,N_11056,N_11691);
xnor U12305 (N_12305,N_11407,N_11053);
or U12306 (N_12306,N_11811,N_11579);
or U12307 (N_12307,N_11281,N_11989);
or U12308 (N_12308,N_11668,N_11178);
or U12309 (N_12309,N_11562,N_11283);
or U12310 (N_12310,N_11372,N_11351);
xor U12311 (N_12311,N_11920,N_11340);
nand U12312 (N_12312,N_11726,N_11197);
nand U12313 (N_12313,N_11353,N_11847);
nor U12314 (N_12314,N_11505,N_11630);
nand U12315 (N_12315,N_11070,N_11532);
nand U12316 (N_12316,N_11658,N_11474);
and U12317 (N_12317,N_11600,N_11707);
and U12318 (N_12318,N_11722,N_11369);
nor U12319 (N_12319,N_11889,N_11901);
nand U12320 (N_12320,N_11790,N_11892);
and U12321 (N_12321,N_11731,N_11973);
and U12322 (N_12322,N_11362,N_11465);
nor U12323 (N_12323,N_11893,N_11760);
nor U12324 (N_12324,N_11868,N_11392);
or U12325 (N_12325,N_11166,N_11222);
nor U12326 (N_12326,N_11066,N_11671);
nand U12327 (N_12327,N_11858,N_11626);
nor U12328 (N_12328,N_11520,N_11119);
nor U12329 (N_12329,N_11037,N_11226);
or U12330 (N_12330,N_11778,N_11629);
nor U12331 (N_12331,N_11237,N_11583);
and U12332 (N_12332,N_11863,N_11620);
nor U12333 (N_12333,N_11252,N_11370);
xnor U12334 (N_12334,N_11766,N_11338);
xnor U12335 (N_12335,N_11437,N_11315);
and U12336 (N_12336,N_11374,N_11234);
nor U12337 (N_12337,N_11087,N_11235);
nand U12338 (N_12338,N_11991,N_11478);
nand U12339 (N_12339,N_11139,N_11216);
nand U12340 (N_12340,N_11302,N_11065);
or U12341 (N_12341,N_11239,N_11303);
xor U12342 (N_12342,N_11721,N_11210);
nor U12343 (N_12343,N_11480,N_11292);
and U12344 (N_12344,N_11008,N_11567);
xnor U12345 (N_12345,N_11176,N_11740);
or U12346 (N_12346,N_11825,N_11798);
nand U12347 (N_12347,N_11424,N_11306);
nand U12348 (N_12348,N_11363,N_11819);
or U12349 (N_12349,N_11761,N_11625);
nand U12350 (N_12350,N_11808,N_11930);
or U12351 (N_12351,N_11897,N_11214);
nor U12352 (N_12352,N_11240,N_11605);
xor U12353 (N_12353,N_11093,N_11291);
and U12354 (N_12354,N_11009,N_11346);
and U12355 (N_12355,N_11524,N_11101);
and U12356 (N_12356,N_11085,N_11557);
or U12357 (N_12357,N_11907,N_11756);
and U12358 (N_12358,N_11368,N_11806);
nor U12359 (N_12359,N_11869,N_11684);
nand U12360 (N_12360,N_11688,N_11674);
nand U12361 (N_12361,N_11047,N_11441);
and U12362 (N_12362,N_11764,N_11765);
nor U12363 (N_12363,N_11220,N_11486);
and U12364 (N_12364,N_11267,N_11961);
nor U12365 (N_12365,N_11171,N_11382);
xor U12366 (N_12366,N_11617,N_11820);
xor U12367 (N_12367,N_11207,N_11313);
nor U12368 (N_12368,N_11095,N_11842);
or U12369 (N_12369,N_11767,N_11734);
xor U12370 (N_12370,N_11938,N_11810);
or U12371 (N_12371,N_11614,N_11132);
xnor U12372 (N_12372,N_11573,N_11500);
or U12373 (N_12373,N_11737,N_11242);
or U12374 (N_12374,N_11427,N_11716);
and U12375 (N_12375,N_11314,N_11886);
or U12376 (N_12376,N_11299,N_11936);
nor U12377 (N_12377,N_11701,N_11198);
nand U12378 (N_12378,N_11025,N_11777);
or U12379 (N_12379,N_11959,N_11813);
xor U12380 (N_12380,N_11024,N_11460);
nor U12381 (N_12381,N_11568,N_11393);
or U12382 (N_12382,N_11818,N_11487);
and U12383 (N_12383,N_11328,N_11019);
nor U12384 (N_12384,N_11841,N_11461);
xnor U12385 (N_12385,N_11549,N_11028);
xnor U12386 (N_12386,N_11086,N_11036);
xor U12387 (N_12387,N_11769,N_11885);
nand U12388 (N_12388,N_11439,N_11552);
xnor U12389 (N_12389,N_11063,N_11911);
or U12390 (N_12390,N_11163,N_11672);
nor U12391 (N_12391,N_11050,N_11673);
nor U12392 (N_12392,N_11770,N_11031);
nor U12393 (N_12393,N_11705,N_11133);
nor U12394 (N_12394,N_11832,N_11970);
xor U12395 (N_12395,N_11384,N_11997);
nand U12396 (N_12396,N_11588,N_11190);
or U12397 (N_12397,N_11589,N_11046);
nand U12398 (N_12398,N_11941,N_11507);
nor U12399 (N_12399,N_11265,N_11975);
and U12400 (N_12400,N_11094,N_11787);
xnor U12401 (N_12401,N_11982,N_11782);
or U12402 (N_12402,N_11515,N_11122);
xor U12403 (N_12403,N_11837,N_11908);
nor U12404 (N_12404,N_11669,N_11946);
xor U12405 (N_12405,N_11481,N_11155);
nand U12406 (N_12406,N_11124,N_11330);
xor U12407 (N_12407,N_11113,N_11165);
and U12408 (N_12408,N_11453,N_11144);
or U12409 (N_12409,N_11596,N_11402);
or U12410 (N_12410,N_11259,N_11030);
nand U12411 (N_12411,N_11390,N_11856);
xnor U12412 (N_12412,N_11117,N_11547);
or U12413 (N_12413,N_11689,N_11898);
nand U12414 (N_12414,N_11450,N_11954);
or U12415 (N_12415,N_11020,N_11561);
nor U12416 (N_12416,N_11679,N_11747);
or U12417 (N_12417,N_11055,N_11594);
nand U12418 (N_12418,N_11217,N_11681);
nand U12419 (N_12419,N_11279,N_11201);
nor U12420 (N_12420,N_11149,N_11932);
nor U12421 (N_12421,N_11618,N_11816);
xnor U12422 (N_12422,N_11585,N_11090);
xor U12423 (N_12423,N_11359,N_11558);
nand U12424 (N_12424,N_11966,N_11005);
xor U12425 (N_12425,N_11189,N_11988);
nor U12426 (N_12426,N_11396,N_11183);
and U12427 (N_12427,N_11253,N_11262);
or U12428 (N_12428,N_11156,N_11577);
nand U12429 (N_12429,N_11458,N_11170);
nor U12430 (N_12430,N_11319,N_11985);
and U12431 (N_12431,N_11436,N_11238);
and U12432 (N_12432,N_11878,N_11646);
nand U12433 (N_12433,N_11584,N_11366);
nor U12434 (N_12434,N_11206,N_11598);
or U12435 (N_12435,N_11438,N_11164);
nor U12436 (N_12436,N_11457,N_11536);
xor U12437 (N_12437,N_11219,N_11447);
or U12438 (N_12438,N_11499,N_11099);
xnor U12439 (N_12439,N_11014,N_11992);
nor U12440 (N_12440,N_11443,N_11492);
and U12441 (N_12441,N_11723,N_11188);
xor U12442 (N_12442,N_11644,N_11430);
xnor U12443 (N_12443,N_11130,N_11248);
and U12444 (N_12444,N_11986,N_11687);
nand U12445 (N_12445,N_11151,N_11884);
nand U12446 (N_12446,N_11462,N_11230);
nor U12447 (N_12447,N_11102,N_11380);
nand U12448 (N_12448,N_11652,N_11141);
nand U12449 (N_12449,N_11797,N_11404);
nor U12450 (N_12450,N_11397,N_11623);
nor U12451 (N_12451,N_11274,N_11621);
xor U12452 (N_12452,N_11080,N_11759);
xor U12453 (N_12453,N_11525,N_11332);
xor U12454 (N_12454,N_11185,N_11084);
nor U12455 (N_12455,N_11258,N_11454);
or U12456 (N_12456,N_11175,N_11981);
and U12457 (N_12457,N_11993,N_11960);
and U12458 (N_12458,N_11255,N_11660);
nand U12459 (N_12459,N_11471,N_11473);
nor U12460 (N_12460,N_11650,N_11984);
and U12461 (N_12461,N_11696,N_11871);
nand U12462 (N_12462,N_11612,N_11748);
xnor U12463 (N_12463,N_11416,N_11496);
xor U12464 (N_12464,N_11421,N_11755);
nor U12465 (N_12465,N_11796,N_11377);
xnor U12466 (N_12466,N_11875,N_11571);
or U12467 (N_12467,N_11762,N_11865);
and U12468 (N_12468,N_11401,N_11266);
or U12469 (N_12469,N_11326,N_11052);
xor U12470 (N_12470,N_11656,N_11708);
or U12471 (N_12471,N_11682,N_11123);
and U12472 (N_12472,N_11649,N_11459);
or U12473 (N_12473,N_11444,N_11277);
nand U12474 (N_12474,N_11174,N_11475);
or U12475 (N_12475,N_11247,N_11442);
and U12476 (N_12476,N_11754,N_11425);
xnor U12477 (N_12477,N_11969,N_11241);
and U12478 (N_12478,N_11956,N_11078);
nand U12479 (N_12479,N_11514,N_11735);
and U12480 (N_12480,N_11678,N_11309);
xor U12481 (N_12481,N_11029,N_11807);
and U12482 (N_12482,N_11342,N_11489);
nor U12483 (N_12483,N_11336,N_11126);
and U12484 (N_12484,N_11950,N_11159);
xnor U12485 (N_12485,N_11861,N_11750);
nor U12486 (N_12486,N_11260,N_11386);
nand U12487 (N_12487,N_11329,N_11275);
nand U12488 (N_12488,N_11383,N_11849);
nand U12489 (N_12489,N_11714,N_11205);
xnor U12490 (N_12490,N_11516,N_11728);
or U12491 (N_12491,N_11834,N_11615);
or U12492 (N_12492,N_11775,N_11905);
and U12493 (N_12493,N_11114,N_11519);
or U12494 (N_12494,N_11345,N_11414);
nor U12495 (N_12495,N_11964,N_11202);
nand U12496 (N_12496,N_11323,N_11109);
or U12497 (N_12497,N_11162,N_11186);
nand U12498 (N_12498,N_11118,N_11896);
or U12499 (N_12499,N_11664,N_11378);
xor U12500 (N_12500,N_11301,N_11756);
xnor U12501 (N_12501,N_11793,N_11593);
nor U12502 (N_12502,N_11097,N_11088);
xnor U12503 (N_12503,N_11972,N_11475);
or U12504 (N_12504,N_11439,N_11551);
and U12505 (N_12505,N_11037,N_11549);
or U12506 (N_12506,N_11114,N_11666);
xnor U12507 (N_12507,N_11086,N_11269);
nor U12508 (N_12508,N_11195,N_11747);
or U12509 (N_12509,N_11448,N_11839);
or U12510 (N_12510,N_11666,N_11813);
nor U12511 (N_12511,N_11016,N_11831);
or U12512 (N_12512,N_11156,N_11983);
nand U12513 (N_12513,N_11620,N_11442);
and U12514 (N_12514,N_11018,N_11879);
and U12515 (N_12515,N_11634,N_11340);
xnor U12516 (N_12516,N_11696,N_11266);
nand U12517 (N_12517,N_11535,N_11339);
nand U12518 (N_12518,N_11651,N_11493);
or U12519 (N_12519,N_11032,N_11750);
or U12520 (N_12520,N_11135,N_11830);
and U12521 (N_12521,N_11803,N_11907);
xor U12522 (N_12522,N_11246,N_11563);
nor U12523 (N_12523,N_11221,N_11029);
xnor U12524 (N_12524,N_11892,N_11331);
and U12525 (N_12525,N_11004,N_11861);
xor U12526 (N_12526,N_11610,N_11979);
nand U12527 (N_12527,N_11951,N_11494);
xor U12528 (N_12528,N_11122,N_11862);
and U12529 (N_12529,N_11623,N_11420);
nor U12530 (N_12530,N_11356,N_11552);
and U12531 (N_12531,N_11821,N_11663);
nand U12532 (N_12532,N_11701,N_11773);
nor U12533 (N_12533,N_11390,N_11447);
and U12534 (N_12534,N_11867,N_11629);
or U12535 (N_12535,N_11719,N_11519);
nand U12536 (N_12536,N_11877,N_11776);
xor U12537 (N_12537,N_11550,N_11119);
nor U12538 (N_12538,N_11762,N_11777);
nor U12539 (N_12539,N_11430,N_11425);
nor U12540 (N_12540,N_11810,N_11379);
nor U12541 (N_12541,N_11510,N_11269);
xor U12542 (N_12542,N_11759,N_11550);
and U12543 (N_12543,N_11409,N_11376);
xnor U12544 (N_12544,N_11398,N_11525);
and U12545 (N_12545,N_11919,N_11564);
and U12546 (N_12546,N_11889,N_11972);
and U12547 (N_12547,N_11425,N_11526);
nor U12548 (N_12548,N_11821,N_11427);
and U12549 (N_12549,N_11973,N_11537);
or U12550 (N_12550,N_11598,N_11969);
or U12551 (N_12551,N_11304,N_11857);
nor U12552 (N_12552,N_11182,N_11460);
and U12553 (N_12553,N_11812,N_11013);
nor U12554 (N_12554,N_11130,N_11101);
xor U12555 (N_12555,N_11559,N_11286);
nand U12556 (N_12556,N_11200,N_11843);
xor U12557 (N_12557,N_11219,N_11256);
and U12558 (N_12558,N_11637,N_11848);
xor U12559 (N_12559,N_11610,N_11799);
and U12560 (N_12560,N_11160,N_11497);
nand U12561 (N_12561,N_11956,N_11345);
nand U12562 (N_12562,N_11239,N_11595);
nand U12563 (N_12563,N_11352,N_11643);
nor U12564 (N_12564,N_11155,N_11779);
or U12565 (N_12565,N_11010,N_11556);
nand U12566 (N_12566,N_11400,N_11062);
and U12567 (N_12567,N_11727,N_11475);
and U12568 (N_12568,N_11552,N_11581);
and U12569 (N_12569,N_11180,N_11233);
nand U12570 (N_12570,N_11031,N_11203);
or U12571 (N_12571,N_11003,N_11846);
and U12572 (N_12572,N_11156,N_11822);
and U12573 (N_12573,N_11902,N_11831);
xor U12574 (N_12574,N_11521,N_11249);
nand U12575 (N_12575,N_11934,N_11017);
and U12576 (N_12576,N_11873,N_11540);
nand U12577 (N_12577,N_11525,N_11550);
or U12578 (N_12578,N_11072,N_11109);
nand U12579 (N_12579,N_11826,N_11706);
xor U12580 (N_12580,N_11708,N_11630);
nor U12581 (N_12581,N_11616,N_11642);
nand U12582 (N_12582,N_11954,N_11483);
or U12583 (N_12583,N_11997,N_11626);
or U12584 (N_12584,N_11744,N_11823);
nor U12585 (N_12585,N_11617,N_11542);
xnor U12586 (N_12586,N_11458,N_11870);
nor U12587 (N_12587,N_11149,N_11974);
or U12588 (N_12588,N_11706,N_11393);
xor U12589 (N_12589,N_11787,N_11292);
xor U12590 (N_12590,N_11511,N_11866);
nor U12591 (N_12591,N_11919,N_11897);
nand U12592 (N_12592,N_11253,N_11440);
and U12593 (N_12593,N_11956,N_11757);
or U12594 (N_12594,N_11795,N_11011);
and U12595 (N_12595,N_11646,N_11764);
nand U12596 (N_12596,N_11114,N_11569);
nand U12597 (N_12597,N_11730,N_11331);
and U12598 (N_12598,N_11315,N_11753);
nand U12599 (N_12599,N_11249,N_11955);
nor U12600 (N_12600,N_11642,N_11237);
or U12601 (N_12601,N_11981,N_11688);
and U12602 (N_12602,N_11960,N_11997);
nand U12603 (N_12603,N_11758,N_11694);
xor U12604 (N_12604,N_11433,N_11809);
nand U12605 (N_12605,N_11029,N_11271);
nand U12606 (N_12606,N_11722,N_11180);
xor U12607 (N_12607,N_11761,N_11454);
nand U12608 (N_12608,N_11814,N_11171);
or U12609 (N_12609,N_11508,N_11174);
nor U12610 (N_12610,N_11392,N_11065);
or U12611 (N_12611,N_11030,N_11399);
or U12612 (N_12612,N_11998,N_11105);
and U12613 (N_12613,N_11327,N_11044);
nand U12614 (N_12614,N_11739,N_11235);
or U12615 (N_12615,N_11632,N_11637);
or U12616 (N_12616,N_11959,N_11841);
xnor U12617 (N_12617,N_11704,N_11265);
nand U12618 (N_12618,N_11095,N_11817);
nor U12619 (N_12619,N_11437,N_11239);
xnor U12620 (N_12620,N_11439,N_11103);
nor U12621 (N_12621,N_11102,N_11996);
nor U12622 (N_12622,N_11510,N_11292);
nor U12623 (N_12623,N_11088,N_11964);
xnor U12624 (N_12624,N_11019,N_11300);
and U12625 (N_12625,N_11884,N_11007);
nand U12626 (N_12626,N_11796,N_11451);
nor U12627 (N_12627,N_11717,N_11700);
nand U12628 (N_12628,N_11424,N_11797);
xor U12629 (N_12629,N_11803,N_11549);
nand U12630 (N_12630,N_11762,N_11485);
nor U12631 (N_12631,N_11277,N_11105);
xnor U12632 (N_12632,N_11465,N_11685);
or U12633 (N_12633,N_11165,N_11740);
or U12634 (N_12634,N_11306,N_11165);
nor U12635 (N_12635,N_11309,N_11444);
xor U12636 (N_12636,N_11581,N_11414);
or U12637 (N_12637,N_11651,N_11187);
xor U12638 (N_12638,N_11675,N_11075);
nor U12639 (N_12639,N_11513,N_11068);
nor U12640 (N_12640,N_11175,N_11098);
xnor U12641 (N_12641,N_11889,N_11337);
or U12642 (N_12642,N_11172,N_11449);
or U12643 (N_12643,N_11503,N_11415);
or U12644 (N_12644,N_11205,N_11411);
xor U12645 (N_12645,N_11695,N_11192);
or U12646 (N_12646,N_11991,N_11264);
xor U12647 (N_12647,N_11606,N_11597);
and U12648 (N_12648,N_11481,N_11116);
nor U12649 (N_12649,N_11586,N_11289);
nor U12650 (N_12650,N_11527,N_11596);
nor U12651 (N_12651,N_11619,N_11975);
or U12652 (N_12652,N_11558,N_11703);
nor U12653 (N_12653,N_11203,N_11824);
and U12654 (N_12654,N_11878,N_11958);
xor U12655 (N_12655,N_11760,N_11052);
nand U12656 (N_12656,N_11240,N_11893);
nor U12657 (N_12657,N_11063,N_11817);
nor U12658 (N_12658,N_11794,N_11323);
and U12659 (N_12659,N_11477,N_11089);
or U12660 (N_12660,N_11608,N_11026);
xor U12661 (N_12661,N_11218,N_11876);
xor U12662 (N_12662,N_11606,N_11032);
nand U12663 (N_12663,N_11368,N_11860);
or U12664 (N_12664,N_11188,N_11517);
xor U12665 (N_12665,N_11525,N_11206);
nor U12666 (N_12666,N_11244,N_11492);
nand U12667 (N_12667,N_11806,N_11734);
xor U12668 (N_12668,N_11481,N_11141);
xor U12669 (N_12669,N_11087,N_11990);
xnor U12670 (N_12670,N_11058,N_11006);
xor U12671 (N_12671,N_11762,N_11254);
nor U12672 (N_12672,N_11465,N_11740);
nor U12673 (N_12673,N_11826,N_11460);
or U12674 (N_12674,N_11563,N_11210);
xor U12675 (N_12675,N_11755,N_11808);
and U12676 (N_12676,N_11094,N_11216);
or U12677 (N_12677,N_11637,N_11541);
and U12678 (N_12678,N_11255,N_11726);
xnor U12679 (N_12679,N_11892,N_11041);
xor U12680 (N_12680,N_11550,N_11786);
xnor U12681 (N_12681,N_11590,N_11489);
or U12682 (N_12682,N_11407,N_11252);
or U12683 (N_12683,N_11134,N_11388);
xor U12684 (N_12684,N_11966,N_11334);
or U12685 (N_12685,N_11467,N_11440);
nor U12686 (N_12686,N_11655,N_11867);
nor U12687 (N_12687,N_11020,N_11825);
and U12688 (N_12688,N_11061,N_11613);
nand U12689 (N_12689,N_11649,N_11991);
xnor U12690 (N_12690,N_11234,N_11687);
xor U12691 (N_12691,N_11806,N_11248);
or U12692 (N_12692,N_11710,N_11388);
or U12693 (N_12693,N_11841,N_11773);
nor U12694 (N_12694,N_11302,N_11990);
and U12695 (N_12695,N_11540,N_11729);
nand U12696 (N_12696,N_11972,N_11397);
nand U12697 (N_12697,N_11027,N_11082);
or U12698 (N_12698,N_11310,N_11568);
nor U12699 (N_12699,N_11059,N_11419);
xor U12700 (N_12700,N_11070,N_11810);
or U12701 (N_12701,N_11673,N_11374);
and U12702 (N_12702,N_11872,N_11635);
and U12703 (N_12703,N_11883,N_11345);
and U12704 (N_12704,N_11882,N_11980);
nor U12705 (N_12705,N_11416,N_11794);
nor U12706 (N_12706,N_11796,N_11633);
nand U12707 (N_12707,N_11009,N_11827);
nor U12708 (N_12708,N_11396,N_11493);
nor U12709 (N_12709,N_11904,N_11641);
and U12710 (N_12710,N_11310,N_11357);
and U12711 (N_12711,N_11390,N_11817);
or U12712 (N_12712,N_11005,N_11791);
or U12713 (N_12713,N_11835,N_11613);
nand U12714 (N_12714,N_11066,N_11589);
and U12715 (N_12715,N_11612,N_11658);
or U12716 (N_12716,N_11194,N_11834);
xnor U12717 (N_12717,N_11856,N_11692);
and U12718 (N_12718,N_11391,N_11695);
and U12719 (N_12719,N_11581,N_11059);
nor U12720 (N_12720,N_11807,N_11196);
nor U12721 (N_12721,N_11290,N_11263);
nand U12722 (N_12722,N_11417,N_11336);
and U12723 (N_12723,N_11131,N_11728);
and U12724 (N_12724,N_11046,N_11764);
xnor U12725 (N_12725,N_11515,N_11189);
xor U12726 (N_12726,N_11923,N_11048);
xor U12727 (N_12727,N_11421,N_11693);
nand U12728 (N_12728,N_11252,N_11776);
nand U12729 (N_12729,N_11118,N_11948);
nor U12730 (N_12730,N_11161,N_11273);
or U12731 (N_12731,N_11417,N_11739);
nand U12732 (N_12732,N_11985,N_11377);
nor U12733 (N_12733,N_11743,N_11783);
nor U12734 (N_12734,N_11539,N_11152);
or U12735 (N_12735,N_11982,N_11967);
nor U12736 (N_12736,N_11176,N_11180);
nor U12737 (N_12737,N_11516,N_11651);
nor U12738 (N_12738,N_11616,N_11568);
nand U12739 (N_12739,N_11005,N_11187);
and U12740 (N_12740,N_11155,N_11124);
and U12741 (N_12741,N_11217,N_11189);
and U12742 (N_12742,N_11255,N_11053);
or U12743 (N_12743,N_11867,N_11897);
nor U12744 (N_12744,N_11451,N_11349);
or U12745 (N_12745,N_11851,N_11265);
and U12746 (N_12746,N_11160,N_11930);
nor U12747 (N_12747,N_11874,N_11430);
nor U12748 (N_12748,N_11918,N_11786);
and U12749 (N_12749,N_11604,N_11030);
or U12750 (N_12750,N_11043,N_11547);
or U12751 (N_12751,N_11191,N_11089);
or U12752 (N_12752,N_11841,N_11748);
nor U12753 (N_12753,N_11659,N_11367);
nor U12754 (N_12754,N_11956,N_11898);
and U12755 (N_12755,N_11937,N_11533);
or U12756 (N_12756,N_11473,N_11004);
xor U12757 (N_12757,N_11053,N_11844);
nor U12758 (N_12758,N_11335,N_11988);
nand U12759 (N_12759,N_11807,N_11760);
and U12760 (N_12760,N_11179,N_11992);
nor U12761 (N_12761,N_11346,N_11823);
and U12762 (N_12762,N_11157,N_11016);
or U12763 (N_12763,N_11986,N_11212);
nand U12764 (N_12764,N_11489,N_11816);
nand U12765 (N_12765,N_11535,N_11422);
nor U12766 (N_12766,N_11976,N_11056);
nor U12767 (N_12767,N_11688,N_11367);
and U12768 (N_12768,N_11820,N_11774);
nand U12769 (N_12769,N_11881,N_11411);
nor U12770 (N_12770,N_11873,N_11064);
and U12771 (N_12771,N_11272,N_11419);
nor U12772 (N_12772,N_11193,N_11036);
or U12773 (N_12773,N_11388,N_11501);
nor U12774 (N_12774,N_11099,N_11166);
nor U12775 (N_12775,N_11658,N_11958);
or U12776 (N_12776,N_11854,N_11172);
nor U12777 (N_12777,N_11738,N_11813);
xor U12778 (N_12778,N_11610,N_11097);
xor U12779 (N_12779,N_11896,N_11699);
xor U12780 (N_12780,N_11215,N_11511);
and U12781 (N_12781,N_11930,N_11412);
and U12782 (N_12782,N_11855,N_11853);
xnor U12783 (N_12783,N_11604,N_11643);
or U12784 (N_12784,N_11683,N_11286);
xor U12785 (N_12785,N_11529,N_11433);
nor U12786 (N_12786,N_11376,N_11757);
nor U12787 (N_12787,N_11284,N_11430);
nor U12788 (N_12788,N_11745,N_11829);
nand U12789 (N_12789,N_11939,N_11721);
nand U12790 (N_12790,N_11347,N_11578);
xor U12791 (N_12791,N_11040,N_11491);
xnor U12792 (N_12792,N_11949,N_11358);
and U12793 (N_12793,N_11002,N_11791);
xnor U12794 (N_12794,N_11052,N_11037);
nor U12795 (N_12795,N_11780,N_11421);
and U12796 (N_12796,N_11436,N_11440);
or U12797 (N_12797,N_11635,N_11947);
nor U12798 (N_12798,N_11390,N_11263);
nand U12799 (N_12799,N_11904,N_11572);
or U12800 (N_12800,N_11527,N_11022);
nor U12801 (N_12801,N_11340,N_11572);
and U12802 (N_12802,N_11311,N_11894);
xnor U12803 (N_12803,N_11052,N_11450);
nor U12804 (N_12804,N_11076,N_11862);
and U12805 (N_12805,N_11174,N_11635);
or U12806 (N_12806,N_11089,N_11258);
nand U12807 (N_12807,N_11400,N_11002);
nand U12808 (N_12808,N_11354,N_11321);
or U12809 (N_12809,N_11026,N_11173);
or U12810 (N_12810,N_11079,N_11772);
nand U12811 (N_12811,N_11708,N_11704);
or U12812 (N_12812,N_11194,N_11626);
nor U12813 (N_12813,N_11221,N_11064);
or U12814 (N_12814,N_11285,N_11830);
or U12815 (N_12815,N_11393,N_11989);
xnor U12816 (N_12816,N_11436,N_11074);
and U12817 (N_12817,N_11368,N_11660);
xor U12818 (N_12818,N_11404,N_11657);
and U12819 (N_12819,N_11713,N_11530);
or U12820 (N_12820,N_11235,N_11881);
xor U12821 (N_12821,N_11855,N_11745);
nand U12822 (N_12822,N_11955,N_11105);
nand U12823 (N_12823,N_11077,N_11379);
xor U12824 (N_12824,N_11986,N_11082);
or U12825 (N_12825,N_11650,N_11218);
and U12826 (N_12826,N_11175,N_11400);
or U12827 (N_12827,N_11420,N_11545);
or U12828 (N_12828,N_11276,N_11547);
nand U12829 (N_12829,N_11947,N_11246);
xor U12830 (N_12830,N_11904,N_11509);
nor U12831 (N_12831,N_11064,N_11053);
or U12832 (N_12832,N_11601,N_11681);
and U12833 (N_12833,N_11050,N_11364);
xor U12834 (N_12834,N_11650,N_11544);
nand U12835 (N_12835,N_11627,N_11603);
and U12836 (N_12836,N_11690,N_11269);
or U12837 (N_12837,N_11185,N_11238);
nand U12838 (N_12838,N_11367,N_11168);
nor U12839 (N_12839,N_11377,N_11086);
nand U12840 (N_12840,N_11020,N_11739);
or U12841 (N_12841,N_11794,N_11067);
and U12842 (N_12842,N_11798,N_11733);
nand U12843 (N_12843,N_11088,N_11031);
xnor U12844 (N_12844,N_11599,N_11814);
xnor U12845 (N_12845,N_11255,N_11608);
nand U12846 (N_12846,N_11958,N_11942);
nand U12847 (N_12847,N_11709,N_11918);
nand U12848 (N_12848,N_11985,N_11063);
nor U12849 (N_12849,N_11335,N_11669);
or U12850 (N_12850,N_11678,N_11639);
and U12851 (N_12851,N_11368,N_11223);
and U12852 (N_12852,N_11922,N_11241);
or U12853 (N_12853,N_11969,N_11731);
nand U12854 (N_12854,N_11842,N_11847);
nor U12855 (N_12855,N_11945,N_11847);
or U12856 (N_12856,N_11432,N_11121);
or U12857 (N_12857,N_11285,N_11117);
nor U12858 (N_12858,N_11737,N_11750);
or U12859 (N_12859,N_11112,N_11016);
nor U12860 (N_12860,N_11648,N_11231);
xor U12861 (N_12861,N_11784,N_11952);
nand U12862 (N_12862,N_11716,N_11263);
nand U12863 (N_12863,N_11790,N_11357);
and U12864 (N_12864,N_11608,N_11046);
nand U12865 (N_12865,N_11211,N_11986);
and U12866 (N_12866,N_11257,N_11756);
nand U12867 (N_12867,N_11928,N_11325);
nor U12868 (N_12868,N_11109,N_11991);
and U12869 (N_12869,N_11148,N_11600);
xnor U12870 (N_12870,N_11097,N_11971);
xnor U12871 (N_12871,N_11619,N_11253);
nand U12872 (N_12872,N_11776,N_11814);
and U12873 (N_12873,N_11238,N_11229);
nor U12874 (N_12874,N_11490,N_11540);
nand U12875 (N_12875,N_11432,N_11471);
nand U12876 (N_12876,N_11813,N_11056);
or U12877 (N_12877,N_11826,N_11187);
xnor U12878 (N_12878,N_11470,N_11326);
nor U12879 (N_12879,N_11474,N_11096);
nand U12880 (N_12880,N_11888,N_11944);
xor U12881 (N_12881,N_11652,N_11423);
or U12882 (N_12882,N_11808,N_11836);
nand U12883 (N_12883,N_11281,N_11516);
xnor U12884 (N_12884,N_11031,N_11678);
or U12885 (N_12885,N_11972,N_11947);
and U12886 (N_12886,N_11121,N_11030);
nand U12887 (N_12887,N_11487,N_11278);
xnor U12888 (N_12888,N_11921,N_11090);
nand U12889 (N_12889,N_11953,N_11237);
nand U12890 (N_12890,N_11300,N_11477);
xor U12891 (N_12891,N_11749,N_11168);
nor U12892 (N_12892,N_11799,N_11559);
and U12893 (N_12893,N_11027,N_11098);
xor U12894 (N_12894,N_11437,N_11104);
nand U12895 (N_12895,N_11698,N_11377);
xor U12896 (N_12896,N_11746,N_11245);
or U12897 (N_12897,N_11717,N_11852);
nand U12898 (N_12898,N_11686,N_11524);
nand U12899 (N_12899,N_11779,N_11176);
and U12900 (N_12900,N_11143,N_11320);
or U12901 (N_12901,N_11205,N_11539);
nor U12902 (N_12902,N_11688,N_11085);
nand U12903 (N_12903,N_11702,N_11164);
or U12904 (N_12904,N_11410,N_11964);
nor U12905 (N_12905,N_11027,N_11868);
and U12906 (N_12906,N_11948,N_11327);
nand U12907 (N_12907,N_11040,N_11298);
nand U12908 (N_12908,N_11335,N_11636);
or U12909 (N_12909,N_11636,N_11501);
and U12910 (N_12910,N_11041,N_11774);
or U12911 (N_12911,N_11518,N_11526);
or U12912 (N_12912,N_11717,N_11816);
xnor U12913 (N_12913,N_11848,N_11835);
nor U12914 (N_12914,N_11763,N_11119);
nand U12915 (N_12915,N_11305,N_11604);
nor U12916 (N_12916,N_11780,N_11685);
or U12917 (N_12917,N_11471,N_11249);
nand U12918 (N_12918,N_11455,N_11398);
nor U12919 (N_12919,N_11527,N_11236);
xor U12920 (N_12920,N_11565,N_11522);
nor U12921 (N_12921,N_11376,N_11103);
or U12922 (N_12922,N_11663,N_11112);
xnor U12923 (N_12923,N_11619,N_11936);
xor U12924 (N_12924,N_11935,N_11194);
and U12925 (N_12925,N_11012,N_11304);
or U12926 (N_12926,N_11156,N_11842);
nand U12927 (N_12927,N_11252,N_11599);
nor U12928 (N_12928,N_11016,N_11310);
or U12929 (N_12929,N_11155,N_11834);
nand U12930 (N_12930,N_11763,N_11236);
or U12931 (N_12931,N_11350,N_11363);
nand U12932 (N_12932,N_11217,N_11415);
and U12933 (N_12933,N_11952,N_11383);
nand U12934 (N_12934,N_11097,N_11641);
and U12935 (N_12935,N_11003,N_11574);
and U12936 (N_12936,N_11986,N_11743);
or U12937 (N_12937,N_11158,N_11265);
nand U12938 (N_12938,N_11262,N_11368);
and U12939 (N_12939,N_11792,N_11364);
nand U12940 (N_12940,N_11482,N_11785);
or U12941 (N_12941,N_11650,N_11633);
and U12942 (N_12942,N_11660,N_11171);
nor U12943 (N_12943,N_11465,N_11455);
nand U12944 (N_12944,N_11636,N_11706);
nor U12945 (N_12945,N_11172,N_11905);
nor U12946 (N_12946,N_11288,N_11375);
nand U12947 (N_12947,N_11910,N_11571);
nor U12948 (N_12948,N_11192,N_11873);
or U12949 (N_12949,N_11816,N_11065);
nand U12950 (N_12950,N_11484,N_11638);
nor U12951 (N_12951,N_11558,N_11570);
or U12952 (N_12952,N_11051,N_11893);
xor U12953 (N_12953,N_11739,N_11298);
nor U12954 (N_12954,N_11753,N_11756);
nand U12955 (N_12955,N_11250,N_11457);
nor U12956 (N_12956,N_11572,N_11760);
and U12957 (N_12957,N_11287,N_11058);
or U12958 (N_12958,N_11857,N_11424);
nand U12959 (N_12959,N_11002,N_11905);
and U12960 (N_12960,N_11018,N_11206);
xnor U12961 (N_12961,N_11673,N_11192);
xnor U12962 (N_12962,N_11798,N_11989);
or U12963 (N_12963,N_11033,N_11124);
xor U12964 (N_12964,N_11532,N_11322);
nand U12965 (N_12965,N_11449,N_11973);
xor U12966 (N_12966,N_11431,N_11441);
and U12967 (N_12967,N_11699,N_11471);
nand U12968 (N_12968,N_11991,N_11636);
nor U12969 (N_12969,N_11815,N_11496);
xor U12970 (N_12970,N_11035,N_11875);
and U12971 (N_12971,N_11108,N_11978);
xnor U12972 (N_12972,N_11874,N_11137);
and U12973 (N_12973,N_11077,N_11709);
or U12974 (N_12974,N_11096,N_11906);
nor U12975 (N_12975,N_11452,N_11291);
nand U12976 (N_12976,N_11492,N_11304);
xor U12977 (N_12977,N_11941,N_11783);
xor U12978 (N_12978,N_11786,N_11489);
or U12979 (N_12979,N_11383,N_11284);
nor U12980 (N_12980,N_11203,N_11229);
nor U12981 (N_12981,N_11055,N_11873);
xnor U12982 (N_12982,N_11170,N_11800);
nor U12983 (N_12983,N_11325,N_11415);
xnor U12984 (N_12984,N_11750,N_11869);
or U12985 (N_12985,N_11911,N_11212);
xor U12986 (N_12986,N_11318,N_11310);
xnor U12987 (N_12987,N_11215,N_11362);
nand U12988 (N_12988,N_11500,N_11658);
xnor U12989 (N_12989,N_11914,N_11150);
nand U12990 (N_12990,N_11870,N_11175);
and U12991 (N_12991,N_11123,N_11744);
xor U12992 (N_12992,N_11303,N_11678);
and U12993 (N_12993,N_11552,N_11418);
nand U12994 (N_12994,N_11900,N_11841);
and U12995 (N_12995,N_11926,N_11915);
nand U12996 (N_12996,N_11376,N_11207);
nor U12997 (N_12997,N_11170,N_11657);
and U12998 (N_12998,N_11630,N_11620);
or U12999 (N_12999,N_11851,N_11085);
and U13000 (N_13000,N_12152,N_12372);
nand U13001 (N_13001,N_12050,N_12027);
xnor U13002 (N_13002,N_12658,N_12205);
or U13003 (N_13003,N_12905,N_12178);
nand U13004 (N_13004,N_12904,N_12528);
nor U13005 (N_13005,N_12560,N_12532);
or U13006 (N_13006,N_12491,N_12717);
or U13007 (N_13007,N_12111,N_12991);
and U13008 (N_13008,N_12595,N_12237);
nor U13009 (N_13009,N_12192,N_12547);
xor U13010 (N_13010,N_12594,N_12196);
and U13011 (N_13011,N_12011,N_12106);
nor U13012 (N_13012,N_12356,N_12202);
xnor U13013 (N_13013,N_12749,N_12033);
and U13014 (N_13014,N_12423,N_12929);
nand U13015 (N_13015,N_12863,N_12030);
nor U13016 (N_13016,N_12850,N_12910);
nand U13017 (N_13017,N_12557,N_12129);
or U13018 (N_13018,N_12825,N_12627);
nand U13019 (N_13019,N_12930,N_12156);
nor U13020 (N_13020,N_12181,N_12988);
xor U13021 (N_13021,N_12374,N_12611);
nand U13022 (N_13022,N_12674,N_12389);
nor U13023 (N_13023,N_12274,N_12698);
nor U13024 (N_13024,N_12358,N_12780);
nand U13025 (N_13025,N_12117,N_12441);
xor U13026 (N_13026,N_12729,N_12644);
nand U13027 (N_13027,N_12250,N_12428);
xor U13028 (N_13028,N_12853,N_12385);
and U13029 (N_13029,N_12555,N_12899);
nor U13030 (N_13030,N_12967,N_12818);
and U13031 (N_13031,N_12999,N_12455);
nand U13032 (N_13032,N_12490,N_12576);
nand U13033 (N_13033,N_12266,N_12151);
xor U13034 (N_13034,N_12961,N_12221);
and U13035 (N_13035,N_12477,N_12494);
nand U13036 (N_13036,N_12907,N_12665);
and U13037 (N_13037,N_12251,N_12878);
and U13038 (N_13038,N_12656,N_12283);
or U13039 (N_13039,N_12335,N_12341);
nand U13040 (N_13040,N_12783,N_12429);
nand U13041 (N_13041,N_12599,N_12330);
or U13042 (N_13042,N_12210,N_12767);
xor U13043 (N_13043,N_12261,N_12233);
and U13044 (N_13044,N_12482,N_12650);
nand U13045 (N_13045,N_12727,N_12831);
nor U13046 (N_13046,N_12039,N_12420);
nor U13047 (N_13047,N_12924,N_12636);
nor U13048 (N_13048,N_12474,N_12996);
nand U13049 (N_13049,N_12125,N_12365);
nor U13050 (N_13050,N_12220,N_12229);
or U13051 (N_13051,N_12077,N_12896);
and U13052 (N_13052,N_12931,N_12579);
nor U13053 (N_13053,N_12406,N_12206);
and U13054 (N_13054,N_12254,N_12268);
or U13055 (N_13055,N_12433,N_12091);
or U13056 (N_13056,N_12239,N_12327);
nor U13057 (N_13057,N_12223,N_12244);
and U13058 (N_13058,N_12546,N_12195);
xnor U13059 (N_13059,N_12504,N_12508);
or U13060 (N_13060,N_12689,N_12534);
or U13061 (N_13061,N_12549,N_12666);
nor U13062 (N_13062,N_12753,N_12982);
and U13063 (N_13063,N_12119,N_12848);
and U13064 (N_13064,N_12804,N_12940);
xnor U13065 (N_13065,N_12681,N_12969);
nor U13066 (N_13066,N_12049,N_12367);
or U13067 (N_13067,N_12760,N_12062);
or U13068 (N_13068,N_12492,N_12165);
xor U13069 (N_13069,N_12144,N_12866);
and U13070 (N_13070,N_12438,N_12874);
xnor U13071 (N_13071,N_12018,N_12216);
or U13072 (N_13072,N_12883,N_12769);
nand U13073 (N_13073,N_12044,N_12805);
xor U13074 (N_13074,N_12456,N_12460);
nor U13075 (N_13075,N_12746,N_12628);
nand U13076 (N_13076,N_12065,N_12744);
nor U13077 (N_13077,N_12885,N_12103);
nor U13078 (N_13078,N_12126,N_12703);
nor U13079 (N_13079,N_12097,N_12677);
nand U13080 (N_13080,N_12522,N_12709);
nor U13081 (N_13081,N_12149,N_12431);
nor U13082 (N_13082,N_12836,N_12912);
xor U13083 (N_13083,N_12445,N_12481);
nand U13084 (N_13084,N_12775,N_12123);
nand U13085 (N_13085,N_12314,N_12046);
or U13086 (N_13086,N_12197,N_12473);
and U13087 (N_13087,N_12407,N_12037);
and U13088 (N_13088,N_12212,N_12166);
xor U13089 (N_13089,N_12034,N_12222);
or U13090 (N_13090,N_12278,N_12059);
and U13091 (N_13091,N_12148,N_12190);
nor U13092 (N_13092,N_12021,N_12104);
nor U13093 (N_13093,N_12626,N_12937);
or U13094 (N_13094,N_12979,N_12102);
nor U13095 (N_13095,N_12082,N_12919);
xor U13096 (N_13096,N_12138,N_12112);
nand U13097 (N_13097,N_12732,N_12000);
and U13098 (N_13098,N_12282,N_12502);
nor U13099 (N_13099,N_12544,N_12267);
or U13100 (N_13100,N_12364,N_12234);
xnor U13101 (N_13101,N_12630,N_12519);
nand U13102 (N_13102,N_12993,N_12252);
nor U13103 (N_13103,N_12830,N_12068);
or U13104 (N_13104,N_12609,N_12755);
nand U13105 (N_13105,N_12213,N_12003);
or U13106 (N_13106,N_12672,N_12277);
nand U13107 (N_13107,N_12561,N_12862);
nor U13108 (N_13108,N_12956,N_12713);
nand U13109 (N_13109,N_12260,N_12770);
and U13110 (N_13110,N_12575,N_12326);
nor U13111 (N_13111,N_12908,N_12435);
and U13112 (N_13112,N_12370,N_12724);
or U13113 (N_13113,N_12621,N_12484);
xor U13114 (N_13114,N_12110,N_12935);
or U13115 (N_13115,N_12538,N_12387);
xor U13116 (N_13116,N_12946,N_12694);
nor U13117 (N_13117,N_12458,N_12145);
or U13118 (N_13118,N_12376,N_12923);
nand U13119 (N_13119,N_12301,N_12699);
xor U13120 (N_13120,N_12584,N_12624);
and U13121 (N_13121,N_12600,N_12945);
or U13122 (N_13122,N_12828,N_12478);
and U13123 (N_13123,N_12401,N_12130);
nand U13124 (N_13124,N_12900,N_12357);
nand U13125 (N_13125,N_12155,N_12537);
xnor U13126 (N_13126,N_12093,N_12486);
nand U13127 (N_13127,N_12936,N_12868);
and U13128 (N_13128,N_12096,N_12392);
nand U13129 (N_13129,N_12015,N_12757);
nor U13130 (N_13130,N_12410,N_12224);
xnor U13131 (N_13131,N_12006,N_12147);
or U13132 (N_13132,N_12328,N_12101);
and U13133 (N_13133,N_12324,N_12997);
xor U13134 (N_13134,N_12132,N_12078);
nor U13135 (N_13135,N_12023,N_12386);
and U13136 (N_13136,N_12291,N_12084);
and U13137 (N_13137,N_12207,N_12542);
xor U13138 (N_13138,N_12901,N_12667);
or U13139 (N_13139,N_12395,N_12648);
nor U13140 (N_13140,N_12976,N_12625);
or U13141 (N_13141,N_12161,N_12142);
and U13142 (N_13142,N_12531,N_12399);
and U13143 (N_13143,N_12005,N_12512);
nand U13144 (N_13144,N_12758,N_12742);
nand U13145 (N_13145,N_12487,N_12054);
nand U13146 (N_13146,N_12682,N_12779);
xor U13147 (N_13147,N_12158,N_12629);
nand U13148 (N_13148,N_12657,N_12505);
nor U13149 (N_13149,N_12743,N_12099);
xor U13150 (N_13150,N_12568,N_12285);
or U13151 (N_13151,N_12641,N_12163);
xor U13152 (N_13152,N_12655,N_12943);
nand U13153 (N_13153,N_12340,N_12897);
xnor U13154 (N_13154,N_12025,N_12995);
and U13155 (N_13155,N_12128,N_12057);
and U13156 (N_13156,N_12638,N_12871);
nor U13157 (N_13157,N_12289,N_12334);
and U13158 (N_13158,N_12041,N_12659);
nand U13159 (N_13159,N_12001,N_12447);
or U13160 (N_13160,N_12735,N_12766);
xnor U13161 (N_13161,N_12020,N_12619);
and U13162 (N_13162,N_12829,N_12708);
nand U13163 (N_13163,N_12509,N_12719);
or U13164 (N_13164,N_12368,N_12499);
nor U13165 (N_13165,N_12591,N_12517);
xnor U13166 (N_13166,N_12247,N_12610);
xnor U13167 (N_13167,N_12095,N_12845);
xor U13168 (N_13168,N_12759,N_12418);
nor U13169 (N_13169,N_12596,N_12498);
xor U13170 (N_13170,N_12772,N_12986);
nand U13171 (N_13171,N_12182,N_12823);
and U13172 (N_13172,N_12564,N_12405);
nand U13173 (N_13173,N_12331,N_12318);
and U13174 (N_13174,N_12605,N_12715);
or U13175 (N_13175,N_12857,N_12462);
xor U13176 (N_13176,N_12738,N_12243);
xor U13177 (N_13177,N_12660,N_12043);
nor U13178 (N_13178,N_12211,N_12572);
nand U13179 (N_13179,N_12664,N_12839);
or U13180 (N_13180,N_12651,N_12606);
and U13181 (N_13181,N_12457,N_12920);
xnor U13182 (N_13182,N_12990,N_12194);
nor U13183 (N_13183,N_12061,N_12977);
xor U13184 (N_13184,N_12203,N_12683);
and U13185 (N_13185,N_12565,N_12279);
nand U13186 (N_13186,N_12157,N_12747);
nand U13187 (N_13187,N_12762,N_12799);
or U13188 (N_13188,N_12721,N_12942);
xor U13189 (N_13189,N_12860,N_12796);
or U13190 (N_13190,N_12476,N_12362);
nand U13191 (N_13191,N_12443,N_12284);
nand U13192 (N_13192,N_12789,N_12360);
xnor U13193 (N_13193,N_12493,N_12671);
and U13194 (N_13194,N_12852,N_12613);
or U13195 (N_13195,N_12019,N_12412);
and U13196 (N_13196,N_12135,N_12134);
nor U13197 (N_13197,N_12464,N_12972);
xor U13198 (N_13198,N_12242,N_12649);
and U13199 (N_13199,N_12179,N_12470);
nor U13200 (N_13200,N_12741,N_12696);
nor U13201 (N_13201,N_12847,N_12807);
nor U13202 (N_13202,N_12336,N_12892);
xnor U13203 (N_13203,N_12926,N_12914);
xnor U13204 (N_13204,N_12167,N_12026);
nor U13205 (N_13205,N_12329,N_12844);
and U13206 (N_13206,N_12425,N_12631);
or U13207 (N_13207,N_12204,N_12922);
and U13208 (N_13208,N_12246,N_12814);
nand U13209 (N_13209,N_12238,N_12558);
or U13210 (N_13210,N_12140,N_12098);
or U13211 (N_13211,N_12058,N_12562);
nand U13212 (N_13212,N_12984,N_12422);
and U13213 (N_13213,N_12583,N_12589);
xnor U13214 (N_13214,N_12894,N_12983);
nand U13215 (N_13215,N_12645,N_12468);
xnor U13216 (N_13216,N_12618,N_12052);
nor U13217 (N_13217,N_12307,N_12380);
nand U13218 (N_13218,N_12784,N_12551);
or U13219 (N_13219,N_12373,N_12465);
nand U13220 (N_13220,N_12859,N_12765);
nand U13221 (N_13221,N_12797,N_12716);
or U13222 (N_13222,N_12722,N_12520);
or U13223 (N_13223,N_12075,N_12409);
and U13224 (N_13224,N_12957,N_12245);
and U13225 (N_13225,N_12343,N_12950);
xnor U13226 (N_13226,N_12559,N_12236);
nand U13227 (N_13227,N_12550,N_12933);
and U13228 (N_13228,N_12603,N_12578);
nand U13229 (N_13229,N_12515,N_12320);
nand U13230 (N_13230,N_12017,N_12281);
and U13231 (N_13231,N_12824,N_12426);
and U13232 (N_13232,N_12060,N_12678);
nand U13233 (N_13233,N_12288,N_12706);
or U13234 (N_13234,N_12835,N_12903);
and U13235 (N_13235,N_12571,N_12411);
nand U13236 (N_13236,N_12662,N_12529);
xor U13237 (N_13237,N_12230,N_12653);
xor U13238 (N_13238,N_12469,N_12339);
and U13239 (N_13239,N_12815,N_12918);
nor U13240 (N_13240,N_12186,N_12856);
and U13241 (N_13241,N_12014,N_12734);
nor U13242 (N_13242,N_12858,N_12604);
nand U13243 (N_13243,N_12688,N_12171);
or U13244 (N_13244,N_12094,N_12371);
and U13245 (N_13245,N_12566,N_12394);
and U13246 (N_13246,N_12120,N_12042);
xnor U13247 (N_13247,N_12820,N_12841);
or U13248 (N_13248,N_12241,N_12726);
and U13249 (N_13249,N_12002,N_12507);
and U13250 (N_13250,N_12752,N_12116);
and U13251 (N_13251,N_12881,N_12524);
xnor U13252 (N_13252,N_12773,N_12353);
xnor U13253 (N_13253,N_12834,N_12137);
and U13254 (N_13254,N_12276,N_12518);
nand U13255 (N_13255,N_12113,N_12055);
nand U13256 (N_13256,N_12813,N_12781);
and U13257 (N_13257,N_12275,N_12887);
nor U13258 (N_13258,N_12180,N_12310);
nand U13259 (N_13259,N_12676,N_12416);
and U13260 (N_13260,N_12258,N_12304);
or U13261 (N_13261,N_12016,N_12122);
nand U13262 (N_13262,N_12654,N_12293);
and U13263 (N_13263,N_12840,N_12467);
or U13264 (N_13264,N_12612,N_12963);
and U13265 (N_13265,N_12865,N_12338);
and U13266 (N_13266,N_12793,N_12436);
nand U13267 (N_13267,N_12777,N_12483);
nand U13268 (N_13268,N_12442,N_12527);
or U13269 (N_13269,N_12553,N_12168);
or U13270 (N_13270,N_12427,N_12215);
nand U13271 (N_13271,N_12185,N_12174);
nand U13272 (N_13272,N_12615,N_12861);
or U13273 (N_13273,N_12637,N_12500);
xor U13274 (N_13274,N_12540,N_12927);
and U13275 (N_13275,N_12700,N_12105);
nor U13276 (N_13276,N_12240,N_12915);
nand U13277 (N_13277,N_12714,N_12567);
xnor U13278 (N_13278,N_12346,N_12071);
or U13279 (N_13279,N_12286,N_12227);
or U13280 (N_13280,N_12088,N_12306);
xnor U13281 (N_13281,N_12375,N_12439);
xor U13282 (N_13282,N_12882,N_12748);
xor U13283 (N_13283,N_12782,N_12430);
nor U13284 (N_13284,N_12256,N_12292);
nand U13285 (N_13285,N_12846,N_12309);
nor U13286 (N_13286,N_12146,N_12255);
xnor U13287 (N_13287,N_12987,N_12728);
and U13288 (N_13288,N_12925,N_12763);
nor U13289 (N_13289,N_12889,N_12315);
nand U13290 (N_13290,N_12786,N_12459);
or U13291 (N_13291,N_12843,N_12086);
or U13292 (N_13292,N_12994,N_12622);
and U13293 (N_13293,N_12479,N_12536);
or U13294 (N_13294,N_12109,N_12970);
or U13295 (N_13295,N_12022,N_12488);
and U13296 (N_13296,N_12952,N_12898);
nand U13297 (N_13297,N_12806,N_12890);
nand U13298 (N_13298,N_12842,N_12377);
or U13299 (N_13299,N_12217,N_12087);
nand U13300 (N_13300,N_12177,N_12415);
and U13301 (N_13301,N_12740,N_12249);
nand U13302 (N_13302,N_12063,N_12776);
xnor U13303 (N_13303,N_12691,N_12495);
nand U13304 (N_13304,N_12880,N_12838);
or U13305 (N_13305,N_12219,N_12774);
and U13306 (N_13306,N_12798,N_12642);
nand U13307 (N_13307,N_12962,N_12960);
and U13308 (N_13308,N_12640,N_12208);
xnor U13309 (N_13309,N_12802,N_12349);
nand U13310 (N_13310,N_12351,N_12663);
or U13311 (N_13311,N_12200,N_12073);
nand U13312 (N_13312,N_12643,N_12964);
xnor U13313 (N_13313,N_12928,N_12879);
nor U13314 (N_13314,N_12556,N_12833);
nand U13315 (N_13315,N_12697,N_12201);
xnor U13316 (N_13316,N_12010,N_12620);
nand U13317 (N_13317,N_12391,N_12383);
or U13318 (N_13318,N_12297,N_12031);
or U13319 (N_13319,N_12647,N_12670);
nand U13320 (N_13320,N_12723,N_12809);
or U13321 (N_13321,N_12958,N_12390);
xor U13322 (N_13322,N_12736,N_12264);
nand U13323 (N_13323,N_12272,N_12989);
xor U13324 (N_13324,N_12811,N_12695);
and U13325 (N_13325,N_12127,N_12601);
nand U13326 (N_13326,N_12702,N_12849);
xnor U13327 (N_13327,N_12398,N_12693);
xor U13328 (N_13328,N_12535,N_12573);
nand U13329 (N_13329,N_12563,N_12543);
nand U13330 (N_13330,N_12248,N_12633);
nand U13331 (N_13331,N_12554,N_12705);
nor U13332 (N_13332,N_12669,N_12616);
or U13333 (N_13333,N_12303,N_12257);
xor U13334 (N_13334,N_12108,N_12253);
nor U13335 (N_13335,N_12322,N_12974);
xnor U13336 (N_13336,N_12004,N_12617);
xor U13337 (N_13337,N_12581,N_12029);
and U13338 (N_13338,N_12232,N_12294);
or U13339 (N_13339,N_12751,N_12819);
xnor U13340 (N_13340,N_12100,N_12745);
or U13341 (N_13341,N_12541,N_12143);
or U13342 (N_13342,N_12263,N_12090);
and U13343 (N_13343,N_12271,N_12737);
and U13344 (N_13344,N_12333,N_12066);
xor U13345 (N_13345,N_12981,N_12837);
nor U13346 (N_13346,N_12822,N_12440);
and U13347 (N_13347,N_12235,N_12184);
or U13348 (N_13348,N_12189,N_12345);
nand U13349 (N_13349,N_12718,N_12506);
and U13350 (N_13350,N_12877,N_12154);
or U13351 (N_13351,N_12397,N_12051);
nand U13352 (N_13352,N_12570,N_12139);
nand U13353 (N_13353,N_12298,N_12175);
and U13354 (N_13354,N_12354,N_12545);
nor U13355 (N_13355,N_12472,N_12413);
or U13356 (N_13356,N_12593,N_12539);
nand U13357 (N_13357,N_12602,N_12585);
and U13358 (N_13358,N_12720,N_12449);
nand U13359 (N_13359,N_12038,N_12821);
and U13360 (N_13360,N_12854,N_12971);
and U13361 (N_13361,N_12909,N_12299);
and U13362 (N_13362,N_12872,N_12975);
nand U13363 (N_13363,N_12712,N_12218);
and U13364 (N_13364,N_12199,N_12265);
nor U13365 (N_13365,N_12521,N_12081);
nand U13366 (N_13366,N_12684,N_12598);
nor U13367 (N_13367,N_12590,N_12827);
xor U13368 (N_13368,N_12580,N_12704);
xor U13369 (N_13369,N_12574,N_12870);
xnor U13370 (N_13370,N_12998,N_12414);
nor U13371 (N_13371,N_12686,N_12707);
and U13372 (N_13372,N_12685,N_12652);
xor U13373 (N_13373,N_12973,N_12516);
xnor U13374 (N_13374,N_12750,N_12141);
nand U13375 (N_13375,N_12803,N_12417);
nand U13376 (N_13376,N_12121,N_12533);
or U13377 (N_13377,N_12454,N_12463);
nand U13378 (N_13378,N_12635,N_12771);
xnor U13379 (N_13379,N_12947,N_12503);
nor U13380 (N_13380,N_12036,N_12992);
or U13381 (N_13381,N_12968,N_12668);
and U13382 (N_13382,N_12347,N_12136);
nand U13383 (N_13383,N_12812,N_12270);
or U13384 (N_13384,N_12592,N_12312);
xor U13385 (N_13385,N_12290,N_12188);
and U13386 (N_13386,N_12949,N_12225);
or U13387 (N_13387,N_12404,N_12118);
xnor U13388 (N_13388,N_12756,N_12954);
xor U13389 (N_13389,N_12785,N_12980);
or U13390 (N_13390,N_12089,N_12496);
nand U13391 (N_13391,N_12466,N_12150);
nor U13392 (N_13392,N_12959,N_12893);
xor U13393 (N_13393,N_12679,N_12342);
nand U13394 (N_13394,N_12434,N_12768);
or U13395 (N_13395,N_12193,N_12906);
and U13396 (N_13396,N_12164,N_12733);
and U13397 (N_13397,N_12067,N_12739);
xor U13398 (N_13398,N_12754,N_12032);
or U13399 (N_13399,N_12944,N_12384);
xnor U13400 (N_13400,N_12092,N_12191);
nor U13401 (N_13401,N_12419,N_12396);
and U13402 (N_13402,N_12424,N_12361);
or U13403 (N_13403,N_12526,N_12913);
nand U13404 (N_13404,N_12064,N_12586);
xor U13405 (N_13405,N_12808,N_12160);
and U13406 (N_13406,N_12891,N_12902);
or U13407 (N_13407,N_12296,N_12884);
nor U13408 (N_13408,N_12169,N_12608);
xnor U13409 (N_13409,N_12226,N_12269);
or U13410 (N_13410,N_12582,N_12461);
nor U13411 (N_13411,N_12939,N_12437);
nand U13412 (N_13412,N_12480,N_12114);
nor U13413 (N_13413,N_12730,N_12587);
nor U13414 (N_13414,N_12778,N_12083);
and U13415 (N_13415,N_12895,N_12305);
nor U13416 (N_13416,N_12795,N_12170);
and U13417 (N_13417,N_12366,N_12382);
xnor U13418 (N_13418,N_12951,N_12597);
or U13419 (N_13419,N_12209,N_12888);
or U13420 (N_13420,N_12378,N_12323);
and U13421 (N_13421,N_12875,N_12725);
nand U13422 (N_13422,N_12007,N_12325);
and U13423 (N_13423,N_12731,N_12869);
or U13424 (N_13424,N_12408,N_12965);
and U13425 (N_13425,N_12183,N_12173);
and U13426 (N_13426,N_12794,N_12316);
xnor U13427 (N_13427,N_12826,N_12363);
or U13428 (N_13428,N_12639,N_12280);
nand U13429 (N_13429,N_12402,N_12867);
xor U13430 (N_13430,N_12337,N_12788);
and U13431 (N_13431,N_12444,N_12344);
and U13432 (N_13432,N_12053,N_12810);
nand U13433 (N_13433,N_12317,N_12450);
or U13434 (N_13434,N_12953,N_12917);
nor U13435 (N_13435,N_12485,N_12024);
nor U13436 (N_13436,N_12510,N_12159);
or U13437 (N_13437,N_12047,N_12941);
or U13438 (N_13438,N_12079,N_12311);
nor U13439 (N_13439,N_12153,N_12632);
and U13440 (N_13440,N_12985,N_12355);
nand U13441 (N_13441,N_12045,N_12332);
and U13442 (N_13442,N_12228,N_12056);
xnor U13443 (N_13443,N_12787,N_12012);
or U13444 (N_13444,N_12214,N_12548);
nor U13445 (N_13445,N_12801,N_12911);
xor U13446 (N_13446,N_12133,N_12076);
nand U13447 (N_13447,N_12687,N_12489);
nand U13448 (N_13448,N_12471,N_12231);
nand U13449 (N_13449,N_12511,N_12313);
nand U13450 (N_13450,N_12432,N_12701);
nor U13451 (N_13451,N_12131,N_12817);
xor U13452 (N_13452,N_12623,N_12388);
nand U13453 (N_13453,N_12259,N_12028);
or U13454 (N_13454,N_12569,N_12369);
and U13455 (N_13455,N_12302,N_12851);
and U13456 (N_13456,N_12832,N_12514);
xnor U13457 (N_13457,N_12008,N_12400);
nor U13458 (N_13458,N_12634,N_12287);
nor U13459 (N_13459,N_12308,N_12873);
and U13460 (N_13460,N_12273,N_12262);
or U13461 (N_13461,N_12176,N_12451);
xor U13462 (N_13462,N_12607,N_12938);
or U13463 (N_13463,N_12864,N_12124);
and U13464 (N_13464,N_12074,N_12921);
and U13465 (N_13465,N_12948,N_12614);
nor U13466 (N_13466,N_12523,N_12321);
or U13467 (N_13467,N_12577,N_12816);
nor U13468 (N_13468,N_12080,N_12513);
nand U13469 (N_13469,N_12453,N_12359);
xor U13470 (N_13470,N_12530,N_12452);
xnor U13471 (N_13471,N_12525,N_12588);
and U13472 (N_13472,N_12448,N_12932);
xor U13473 (N_13473,N_12978,N_12172);
and U13474 (N_13474,N_12393,N_12855);
or U13475 (N_13475,N_12403,N_12013);
and U13476 (N_13476,N_12198,N_12646);
xor U13477 (N_13477,N_12300,N_12673);
nand U13478 (N_13478,N_12966,N_12035);
and U13479 (N_13479,N_12916,N_12692);
and U13480 (N_13480,N_12381,N_12348);
and U13481 (N_13481,N_12475,N_12792);
nand U13482 (N_13482,N_12501,N_12295);
xnor U13483 (N_13483,N_12350,N_12680);
nand U13484 (N_13484,N_12791,N_12764);
xnor U13485 (N_13485,N_12115,N_12710);
and U13486 (N_13486,N_12009,N_12675);
nand U13487 (N_13487,N_12886,N_12690);
nand U13488 (N_13488,N_12446,N_12162);
xnor U13489 (N_13489,N_12040,N_12552);
or U13490 (N_13490,N_12085,N_12934);
xor U13491 (N_13491,N_12048,N_12187);
and U13492 (N_13492,N_12661,N_12319);
xor U13493 (N_13493,N_12955,N_12800);
nand U13494 (N_13494,N_12790,N_12876);
nor U13495 (N_13495,N_12379,N_12072);
nor U13496 (N_13496,N_12070,N_12107);
nor U13497 (N_13497,N_12761,N_12497);
and U13498 (N_13498,N_12069,N_12711);
xor U13499 (N_13499,N_12421,N_12352);
or U13500 (N_13500,N_12387,N_12901);
and U13501 (N_13501,N_12122,N_12609);
and U13502 (N_13502,N_12684,N_12743);
and U13503 (N_13503,N_12014,N_12932);
and U13504 (N_13504,N_12472,N_12192);
nand U13505 (N_13505,N_12265,N_12099);
nand U13506 (N_13506,N_12873,N_12589);
or U13507 (N_13507,N_12573,N_12588);
nand U13508 (N_13508,N_12477,N_12499);
xnor U13509 (N_13509,N_12232,N_12405);
nand U13510 (N_13510,N_12195,N_12255);
nor U13511 (N_13511,N_12428,N_12819);
or U13512 (N_13512,N_12065,N_12311);
and U13513 (N_13513,N_12265,N_12595);
xnor U13514 (N_13514,N_12117,N_12113);
xnor U13515 (N_13515,N_12619,N_12893);
or U13516 (N_13516,N_12590,N_12319);
nor U13517 (N_13517,N_12526,N_12392);
nand U13518 (N_13518,N_12651,N_12467);
nand U13519 (N_13519,N_12318,N_12845);
or U13520 (N_13520,N_12589,N_12737);
or U13521 (N_13521,N_12482,N_12101);
nand U13522 (N_13522,N_12724,N_12715);
and U13523 (N_13523,N_12772,N_12968);
nor U13524 (N_13524,N_12742,N_12333);
nand U13525 (N_13525,N_12712,N_12982);
or U13526 (N_13526,N_12912,N_12968);
nor U13527 (N_13527,N_12694,N_12516);
nor U13528 (N_13528,N_12104,N_12878);
nand U13529 (N_13529,N_12517,N_12158);
nor U13530 (N_13530,N_12821,N_12856);
nor U13531 (N_13531,N_12355,N_12278);
xor U13532 (N_13532,N_12583,N_12197);
and U13533 (N_13533,N_12172,N_12420);
and U13534 (N_13534,N_12215,N_12782);
xor U13535 (N_13535,N_12877,N_12627);
or U13536 (N_13536,N_12748,N_12269);
xor U13537 (N_13537,N_12895,N_12851);
nand U13538 (N_13538,N_12435,N_12504);
xor U13539 (N_13539,N_12583,N_12615);
and U13540 (N_13540,N_12627,N_12211);
and U13541 (N_13541,N_12645,N_12826);
nor U13542 (N_13542,N_12122,N_12026);
nor U13543 (N_13543,N_12101,N_12447);
and U13544 (N_13544,N_12776,N_12774);
nor U13545 (N_13545,N_12673,N_12428);
and U13546 (N_13546,N_12842,N_12477);
xnor U13547 (N_13547,N_12124,N_12644);
and U13548 (N_13548,N_12375,N_12932);
and U13549 (N_13549,N_12366,N_12757);
and U13550 (N_13550,N_12846,N_12719);
and U13551 (N_13551,N_12174,N_12558);
xor U13552 (N_13552,N_12168,N_12760);
or U13553 (N_13553,N_12915,N_12576);
xnor U13554 (N_13554,N_12873,N_12560);
or U13555 (N_13555,N_12918,N_12993);
xor U13556 (N_13556,N_12966,N_12080);
or U13557 (N_13557,N_12066,N_12372);
and U13558 (N_13558,N_12503,N_12854);
xnor U13559 (N_13559,N_12438,N_12876);
and U13560 (N_13560,N_12009,N_12726);
nor U13561 (N_13561,N_12232,N_12651);
and U13562 (N_13562,N_12162,N_12851);
nor U13563 (N_13563,N_12089,N_12920);
nor U13564 (N_13564,N_12718,N_12934);
xor U13565 (N_13565,N_12971,N_12758);
nor U13566 (N_13566,N_12982,N_12848);
or U13567 (N_13567,N_12012,N_12826);
or U13568 (N_13568,N_12031,N_12941);
nor U13569 (N_13569,N_12593,N_12868);
nor U13570 (N_13570,N_12172,N_12008);
nand U13571 (N_13571,N_12885,N_12562);
nor U13572 (N_13572,N_12260,N_12810);
nor U13573 (N_13573,N_12107,N_12770);
or U13574 (N_13574,N_12549,N_12212);
and U13575 (N_13575,N_12212,N_12503);
or U13576 (N_13576,N_12505,N_12577);
or U13577 (N_13577,N_12875,N_12805);
or U13578 (N_13578,N_12974,N_12418);
xor U13579 (N_13579,N_12291,N_12331);
and U13580 (N_13580,N_12333,N_12793);
or U13581 (N_13581,N_12441,N_12981);
nand U13582 (N_13582,N_12202,N_12806);
nand U13583 (N_13583,N_12136,N_12202);
nand U13584 (N_13584,N_12121,N_12510);
nand U13585 (N_13585,N_12109,N_12893);
xor U13586 (N_13586,N_12459,N_12894);
and U13587 (N_13587,N_12641,N_12324);
and U13588 (N_13588,N_12973,N_12747);
and U13589 (N_13589,N_12152,N_12303);
nor U13590 (N_13590,N_12052,N_12878);
nand U13591 (N_13591,N_12437,N_12319);
and U13592 (N_13592,N_12150,N_12560);
nor U13593 (N_13593,N_12399,N_12125);
and U13594 (N_13594,N_12564,N_12903);
nand U13595 (N_13595,N_12340,N_12584);
nand U13596 (N_13596,N_12437,N_12817);
nor U13597 (N_13597,N_12791,N_12890);
nand U13598 (N_13598,N_12952,N_12212);
and U13599 (N_13599,N_12178,N_12013);
nand U13600 (N_13600,N_12934,N_12801);
xnor U13601 (N_13601,N_12456,N_12262);
xnor U13602 (N_13602,N_12499,N_12960);
nand U13603 (N_13603,N_12619,N_12975);
nor U13604 (N_13604,N_12044,N_12658);
xnor U13605 (N_13605,N_12963,N_12016);
xor U13606 (N_13606,N_12985,N_12931);
nand U13607 (N_13607,N_12451,N_12481);
and U13608 (N_13608,N_12247,N_12801);
nand U13609 (N_13609,N_12892,N_12019);
nor U13610 (N_13610,N_12273,N_12086);
nor U13611 (N_13611,N_12457,N_12785);
nor U13612 (N_13612,N_12396,N_12324);
and U13613 (N_13613,N_12021,N_12056);
nor U13614 (N_13614,N_12522,N_12553);
and U13615 (N_13615,N_12613,N_12247);
nor U13616 (N_13616,N_12205,N_12534);
nor U13617 (N_13617,N_12154,N_12536);
nor U13618 (N_13618,N_12880,N_12836);
and U13619 (N_13619,N_12415,N_12849);
or U13620 (N_13620,N_12984,N_12219);
nor U13621 (N_13621,N_12964,N_12174);
or U13622 (N_13622,N_12386,N_12144);
nand U13623 (N_13623,N_12872,N_12346);
nor U13624 (N_13624,N_12165,N_12294);
xnor U13625 (N_13625,N_12319,N_12024);
xor U13626 (N_13626,N_12212,N_12685);
xor U13627 (N_13627,N_12636,N_12200);
nor U13628 (N_13628,N_12437,N_12447);
and U13629 (N_13629,N_12656,N_12824);
or U13630 (N_13630,N_12601,N_12329);
nand U13631 (N_13631,N_12986,N_12565);
xnor U13632 (N_13632,N_12679,N_12537);
or U13633 (N_13633,N_12193,N_12591);
or U13634 (N_13634,N_12085,N_12049);
or U13635 (N_13635,N_12532,N_12861);
or U13636 (N_13636,N_12700,N_12047);
and U13637 (N_13637,N_12929,N_12036);
nor U13638 (N_13638,N_12051,N_12112);
nor U13639 (N_13639,N_12463,N_12641);
nor U13640 (N_13640,N_12464,N_12761);
or U13641 (N_13641,N_12894,N_12575);
or U13642 (N_13642,N_12918,N_12064);
or U13643 (N_13643,N_12490,N_12921);
nand U13644 (N_13644,N_12791,N_12199);
nor U13645 (N_13645,N_12587,N_12860);
xnor U13646 (N_13646,N_12767,N_12077);
nand U13647 (N_13647,N_12668,N_12093);
or U13648 (N_13648,N_12868,N_12718);
and U13649 (N_13649,N_12499,N_12402);
and U13650 (N_13650,N_12498,N_12138);
nor U13651 (N_13651,N_12599,N_12255);
nand U13652 (N_13652,N_12199,N_12079);
nand U13653 (N_13653,N_12380,N_12459);
or U13654 (N_13654,N_12506,N_12369);
nand U13655 (N_13655,N_12659,N_12241);
nor U13656 (N_13656,N_12125,N_12599);
nor U13657 (N_13657,N_12840,N_12211);
or U13658 (N_13658,N_12058,N_12472);
and U13659 (N_13659,N_12406,N_12924);
or U13660 (N_13660,N_12328,N_12205);
nor U13661 (N_13661,N_12584,N_12223);
or U13662 (N_13662,N_12478,N_12613);
and U13663 (N_13663,N_12353,N_12933);
nand U13664 (N_13664,N_12274,N_12575);
or U13665 (N_13665,N_12998,N_12605);
and U13666 (N_13666,N_12171,N_12804);
and U13667 (N_13667,N_12592,N_12381);
and U13668 (N_13668,N_12478,N_12903);
or U13669 (N_13669,N_12876,N_12033);
and U13670 (N_13670,N_12472,N_12153);
and U13671 (N_13671,N_12710,N_12633);
nor U13672 (N_13672,N_12142,N_12343);
nor U13673 (N_13673,N_12993,N_12499);
xor U13674 (N_13674,N_12688,N_12091);
xor U13675 (N_13675,N_12721,N_12468);
nor U13676 (N_13676,N_12886,N_12145);
and U13677 (N_13677,N_12224,N_12541);
or U13678 (N_13678,N_12566,N_12723);
and U13679 (N_13679,N_12528,N_12503);
or U13680 (N_13680,N_12106,N_12945);
nand U13681 (N_13681,N_12485,N_12604);
nor U13682 (N_13682,N_12698,N_12621);
or U13683 (N_13683,N_12017,N_12137);
nand U13684 (N_13684,N_12697,N_12760);
or U13685 (N_13685,N_12243,N_12218);
nor U13686 (N_13686,N_12738,N_12861);
and U13687 (N_13687,N_12204,N_12413);
and U13688 (N_13688,N_12440,N_12368);
nand U13689 (N_13689,N_12735,N_12728);
and U13690 (N_13690,N_12778,N_12014);
nor U13691 (N_13691,N_12524,N_12853);
nor U13692 (N_13692,N_12947,N_12903);
xor U13693 (N_13693,N_12835,N_12265);
nor U13694 (N_13694,N_12348,N_12493);
and U13695 (N_13695,N_12606,N_12354);
nor U13696 (N_13696,N_12899,N_12698);
and U13697 (N_13697,N_12467,N_12222);
xnor U13698 (N_13698,N_12171,N_12410);
nor U13699 (N_13699,N_12959,N_12851);
or U13700 (N_13700,N_12540,N_12348);
nand U13701 (N_13701,N_12784,N_12419);
xnor U13702 (N_13702,N_12742,N_12492);
xnor U13703 (N_13703,N_12209,N_12170);
and U13704 (N_13704,N_12119,N_12098);
or U13705 (N_13705,N_12371,N_12914);
and U13706 (N_13706,N_12839,N_12871);
or U13707 (N_13707,N_12224,N_12815);
xor U13708 (N_13708,N_12078,N_12509);
nand U13709 (N_13709,N_12586,N_12316);
nor U13710 (N_13710,N_12733,N_12891);
or U13711 (N_13711,N_12215,N_12220);
xor U13712 (N_13712,N_12340,N_12140);
nor U13713 (N_13713,N_12019,N_12510);
and U13714 (N_13714,N_12104,N_12704);
xnor U13715 (N_13715,N_12911,N_12920);
or U13716 (N_13716,N_12186,N_12948);
nand U13717 (N_13717,N_12074,N_12460);
or U13718 (N_13718,N_12395,N_12350);
nor U13719 (N_13719,N_12266,N_12159);
or U13720 (N_13720,N_12601,N_12444);
nor U13721 (N_13721,N_12290,N_12491);
or U13722 (N_13722,N_12685,N_12055);
and U13723 (N_13723,N_12495,N_12637);
nor U13724 (N_13724,N_12489,N_12711);
xor U13725 (N_13725,N_12696,N_12215);
and U13726 (N_13726,N_12710,N_12187);
xnor U13727 (N_13727,N_12963,N_12864);
or U13728 (N_13728,N_12072,N_12368);
xor U13729 (N_13729,N_12916,N_12820);
nand U13730 (N_13730,N_12035,N_12536);
nor U13731 (N_13731,N_12284,N_12016);
or U13732 (N_13732,N_12330,N_12585);
nor U13733 (N_13733,N_12927,N_12351);
or U13734 (N_13734,N_12567,N_12862);
and U13735 (N_13735,N_12682,N_12677);
or U13736 (N_13736,N_12766,N_12757);
xnor U13737 (N_13737,N_12140,N_12912);
nor U13738 (N_13738,N_12828,N_12695);
nand U13739 (N_13739,N_12494,N_12615);
and U13740 (N_13740,N_12968,N_12986);
xor U13741 (N_13741,N_12455,N_12712);
nand U13742 (N_13742,N_12209,N_12103);
nor U13743 (N_13743,N_12709,N_12449);
nand U13744 (N_13744,N_12706,N_12687);
and U13745 (N_13745,N_12637,N_12408);
nand U13746 (N_13746,N_12865,N_12883);
or U13747 (N_13747,N_12932,N_12091);
nor U13748 (N_13748,N_12611,N_12878);
and U13749 (N_13749,N_12646,N_12033);
and U13750 (N_13750,N_12869,N_12032);
nor U13751 (N_13751,N_12923,N_12886);
and U13752 (N_13752,N_12906,N_12510);
nand U13753 (N_13753,N_12125,N_12716);
nor U13754 (N_13754,N_12723,N_12351);
or U13755 (N_13755,N_12310,N_12709);
xnor U13756 (N_13756,N_12707,N_12672);
nand U13757 (N_13757,N_12408,N_12098);
and U13758 (N_13758,N_12619,N_12018);
nor U13759 (N_13759,N_12570,N_12476);
xnor U13760 (N_13760,N_12017,N_12766);
xnor U13761 (N_13761,N_12378,N_12321);
xor U13762 (N_13762,N_12053,N_12093);
nor U13763 (N_13763,N_12156,N_12812);
or U13764 (N_13764,N_12293,N_12956);
and U13765 (N_13765,N_12379,N_12532);
and U13766 (N_13766,N_12719,N_12036);
xor U13767 (N_13767,N_12531,N_12239);
or U13768 (N_13768,N_12791,N_12504);
nand U13769 (N_13769,N_12553,N_12667);
or U13770 (N_13770,N_12726,N_12506);
xor U13771 (N_13771,N_12026,N_12912);
nand U13772 (N_13772,N_12232,N_12977);
xnor U13773 (N_13773,N_12490,N_12405);
nand U13774 (N_13774,N_12703,N_12383);
or U13775 (N_13775,N_12014,N_12189);
xor U13776 (N_13776,N_12726,N_12863);
and U13777 (N_13777,N_12120,N_12854);
or U13778 (N_13778,N_12776,N_12899);
nand U13779 (N_13779,N_12012,N_12951);
nand U13780 (N_13780,N_12745,N_12317);
xor U13781 (N_13781,N_12172,N_12914);
nand U13782 (N_13782,N_12481,N_12919);
and U13783 (N_13783,N_12907,N_12060);
xnor U13784 (N_13784,N_12873,N_12915);
and U13785 (N_13785,N_12155,N_12115);
xnor U13786 (N_13786,N_12164,N_12751);
nand U13787 (N_13787,N_12368,N_12223);
nand U13788 (N_13788,N_12007,N_12803);
xor U13789 (N_13789,N_12690,N_12007);
nand U13790 (N_13790,N_12508,N_12971);
and U13791 (N_13791,N_12089,N_12608);
nor U13792 (N_13792,N_12169,N_12263);
or U13793 (N_13793,N_12086,N_12670);
nand U13794 (N_13794,N_12257,N_12058);
or U13795 (N_13795,N_12234,N_12932);
nand U13796 (N_13796,N_12903,N_12425);
xnor U13797 (N_13797,N_12395,N_12185);
and U13798 (N_13798,N_12112,N_12768);
xor U13799 (N_13799,N_12321,N_12670);
xor U13800 (N_13800,N_12480,N_12165);
xnor U13801 (N_13801,N_12432,N_12103);
xor U13802 (N_13802,N_12423,N_12412);
nor U13803 (N_13803,N_12929,N_12824);
nand U13804 (N_13804,N_12907,N_12652);
nor U13805 (N_13805,N_12622,N_12787);
nor U13806 (N_13806,N_12554,N_12904);
nand U13807 (N_13807,N_12151,N_12506);
xnor U13808 (N_13808,N_12372,N_12562);
and U13809 (N_13809,N_12812,N_12818);
and U13810 (N_13810,N_12290,N_12108);
nand U13811 (N_13811,N_12910,N_12077);
nor U13812 (N_13812,N_12231,N_12013);
and U13813 (N_13813,N_12705,N_12601);
and U13814 (N_13814,N_12646,N_12042);
xor U13815 (N_13815,N_12108,N_12249);
and U13816 (N_13816,N_12347,N_12195);
xnor U13817 (N_13817,N_12816,N_12662);
and U13818 (N_13818,N_12931,N_12456);
and U13819 (N_13819,N_12479,N_12176);
xor U13820 (N_13820,N_12515,N_12652);
xnor U13821 (N_13821,N_12724,N_12708);
or U13822 (N_13822,N_12883,N_12700);
nor U13823 (N_13823,N_12190,N_12704);
and U13824 (N_13824,N_12340,N_12763);
or U13825 (N_13825,N_12806,N_12951);
nand U13826 (N_13826,N_12891,N_12156);
nand U13827 (N_13827,N_12940,N_12415);
xnor U13828 (N_13828,N_12078,N_12018);
xnor U13829 (N_13829,N_12935,N_12276);
xnor U13830 (N_13830,N_12405,N_12149);
nand U13831 (N_13831,N_12195,N_12520);
nand U13832 (N_13832,N_12947,N_12626);
nor U13833 (N_13833,N_12438,N_12138);
xnor U13834 (N_13834,N_12965,N_12590);
or U13835 (N_13835,N_12132,N_12369);
or U13836 (N_13836,N_12598,N_12122);
and U13837 (N_13837,N_12519,N_12056);
or U13838 (N_13838,N_12999,N_12567);
nor U13839 (N_13839,N_12388,N_12562);
nor U13840 (N_13840,N_12175,N_12686);
or U13841 (N_13841,N_12098,N_12711);
nand U13842 (N_13842,N_12936,N_12486);
nand U13843 (N_13843,N_12275,N_12730);
and U13844 (N_13844,N_12087,N_12892);
or U13845 (N_13845,N_12652,N_12789);
and U13846 (N_13846,N_12450,N_12697);
or U13847 (N_13847,N_12707,N_12912);
or U13848 (N_13848,N_12010,N_12887);
and U13849 (N_13849,N_12211,N_12122);
nand U13850 (N_13850,N_12007,N_12384);
xnor U13851 (N_13851,N_12320,N_12812);
xor U13852 (N_13852,N_12234,N_12860);
or U13853 (N_13853,N_12098,N_12028);
nor U13854 (N_13854,N_12625,N_12574);
nor U13855 (N_13855,N_12159,N_12891);
or U13856 (N_13856,N_12386,N_12984);
and U13857 (N_13857,N_12454,N_12255);
nor U13858 (N_13858,N_12009,N_12925);
nand U13859 (N_13859,N_12302,N_12756);
and U13860 (N_13860,N_12416,N_12667);
and U13861 (N_13861,N_12327,N_12165);
or U13862 (N_13862,N_12403,N_12944);
xnor U13863 (N_13863,N_12111,N_12747);
nand U13864 (N_13864,N_12146,N_12819);
nor U13865 (N_13865,N_12887,N_12992);
nand U13866 (N_13866,N_12776,N_12539);
xnor U13867 (N_13867,N_12620,N_12670);
nand U13868 (N_13868,N_12191,N_12503);
xnor U13869 (N_13869,N_12749,N_12714);
nand U13870 (N_13870,N_12431,N_12785);
xnor U13871 (N_13871,N_12922,N_12970);
nor U13872 (N_13872,N_12262,N_12521);
nor U13873 (N_13873,N_12494,N_12481);
nand U13874 (N_13874,N_12086,N_12240);
nor U13875 (N_13875,N_12367,N_12445);
xnor U13876 (N_13876,N_12802,N_12873);
or U13877 (N_13877,N_12707,N_12304);
nand U13878 (N_13878,N_12377,N_12197);
xnor U13879 (N_13879,N_12237,N_12523);
or U13880 (N_13880,N_12305,N_12724);
and U13881 (N_13881,N_12415,N_12572);
or U13882 (N_13882,N_12585,N_12785);
nor U13883 (N_13883,N_12429,N_12106);
nand U13884 (N_13884,N_12834,N_12967);
nand U13885 (N_13885,N_12237,N_12776);
or U13886 (N_13886,N_12568,N_12031);
or U13887 (N_13887,N_12377,N_12450);
or U13888 (N_13888,N_12697,N_12981);
and U13889 (N_13889,N_12590,N_12450);
xnor U13890 (N_13890,N_12994,N_12150);
or U13891 (N_13891,N_12015,N_12577);
nor U13892 (N_13892,N_12220,N_12080);
xor U13893 (N_13893,N_12337,N_12776);
xor U13894 (N_13894,N_12770,N_12781);
xnor U13895 (N_13895,N_12818,N_12617);
or U13896 (N_13896,N_12894,N_12131);
nor U13897 (N_13897,N_12831,N_12379);
and U13898 (N_13898,N_12681,N_12743);
and U13899 (N_13899,N_12357,N_12075);
and U13900 (N_13900,N_12689,N_12788);
xor U13901 (N_13901,N_12910,N_12888);
and U13902 (N_13902,N_12147,N_12691);
and U13903 (N_13903,N_12089,N_12579);
nor U13904 (N_13904,N_12877,N_12946);
nor U13905 (N_13905,N_12277,N_12315);
and U13906 (N_13906,N_12730,N_12596);
xor U13907 (N_13907,N_12046,N_12791);
or U13908 (N_13908,N_12063,N_12159);
nand U13909 (N_13909,N_12534,N_12215);
or U13910 (N_13910,N_12700,N_12289);
and U13911 (N_13911,N_12552,N_12611);
nand U13912 (N_13912,N_12275,N_12709);
nor U13913 (N_13913,N_12293,N_12352);
and U13914 (N_13914,N_12532,N_12430);
nand U13915 (N_13915,N_12116,N_12349);
nand U13916 (N_13916,N_12564,N_12862);
or U13917 (N_13917,N_12094,N_12617);
nand U13918 (N_13918,N_12136,N_12923);
nor U13919 (N_13919,N_12296,N_12862);
or U13920 (N_13920,N_12552,N_12198);
and U13921 (N_13921,N_12793,N_12461);
nand U13922 (N_13922,N_12167,N_12174);
and U13923 (N_13923,N_12174,N_12388);
and U13924 (N_13924,N_12976,N_12395);
nand U13925 (N_13925,N_12677,N_12508);
nand U13926 (N_13926,N_12092,N_12080);
or U13927 (N_13927,N_12902,N_12052);
or U13928 (N_13928,N_12630,N_12500);
and U13929 (N_13929,N_12034,N_12675);
nand U13930 (N_13930,N_12045,N_12675);
nor U13931 (N_13931,N_12505,N_12869);
and U13932 (N_13932,N_12087,N_12263);
or U13933 (N_13933,N_12144,N_12648);
and U13934 (N_13934,N_12677,N_12641);
nor U13935 (N_13935,N_12245,N_12256);
nor U13936 (N_13936,N_12005,N_12465);
or U13937 (N_13937,N_12781,N_12246);
nand U13938 (N_13938,N_12171,N_12550);
nor U13939 (N_13939,N_12520,N_12770);
nor U13940 (N_13940,N_12273,N_12333);
nor U13941 (N_13941,N_12255,N_12137);
and U13942 (N_13942,N_12769,N_12998);
nor U13943 (N_13943,N_12113,N_12873);
nand U13944 (N_13944,N_12462,N_12583);
and U13945 (N_13945,N_12035,N_12527);
nand U13946 (N_13946,N_12903,N_12716);
nor U13947 (N_13947,N_12297,N_12107);
and U13948 (N_13948,N_12737,N_12788);
or U13949 (N_13949,N_12087,N_12221);
nand U13950 (N_13950,N_12742,N_12975);
or U13951 (N_13951,N_12553,N_12024);
or U13952 (N_13952,N_12426,N_12875);
and U13953 (N_13953,N_12632,N_12820);
or U13954 (N_13954,N_12986,N_12907);
nand U13955 (N_13955,N_12777,N_12107);
nand U13956 (N_13956,N_12434,N_12751);
nor U13957 (N_13957,N_12968,N_12083);
xnor U13958 (N_13958,N_12788,N_12639);
nand U13959 (N_13959,N_12398,N_12861);
and U13960 (N_13960,N_12254,N_12984);
and U13961 (N_13961,N_12827,N_12749);
and U13962 (N_13962,N_12158,N_12027);
and U13963 (N_13963,N_12987,N_12629);
and U13964 (N_13964,N_12662,N_12903);
nand U13965 (N_13965,N_12295,N_12118);
and U13966 (N_13966,N_12926,N_12564);
and U13967 (N_13967,N_12958,N_12845);
xnor U13968 (N_13968,N_12836,N_12632);
nand U13969 (N_13969,N_12337,N_12593);
nand U13970 (N_13970,N_12521,N_12938);
xor U13971 (N_13971,N_12154,N_12618);
xor U13972 (N_13972,N_12418,N_12310);
xnor U13973 (N_13973,N_12641,N_12678);
xnor U13974 (N_13974,N_12504,N_12541);
and U13975 (N_13975,N_12770,N_12654);
xnor U13976 (N_13976,N_12254,N_12337);
xnor U13977 (N_13977,N_12317,N_12401);
nor U13978 (N_13978,N_12290,N_12198);
nor U13979 (N_13979,N_12027,N_12532);
and U13980 (N_13980,N_12393,N_12849);
xor U13981 (N_13981,N_12271,N_12894);
xor U13982 (N_13982,N_12747,N_12750);
xor U13983 (N_13983,N_12705,N_12883);
nor U13984 (N_13984,N_12663,N_12915);
nand U13985 (N_13985,N_12410,N_12796);
nand U13986 (N_13986,N_12046,N_12152);
or U13987 (N_13987,N_12123,N_12533);
nand U13988 (N_13988,N_12794,N_12437);
or U13989 (N_13989,N_12233,N_12503);
and U13990 (N_13990,N_12455,N_12403);
xor U13991 (N_13991,N_12825,N_12698);
xor U13992 (N_13992,N_12460,N_12593);
nor U13993 (N_13993,N_12102,N_12392);
nand U13994 (N_13994,N_12026,N_12001);
xnor U13995 (N_13995,N_12501,N_12185);
and U13996 (N_13996,N_12536,N_12444);
and U13997 (N_13997,N_12656,N_12366);
and U13998 (N_13998,N_12945,N_12066);
nor U13999 (N_13999,N_12329,N_12768);
or U14000 (N_14000,N_13360,N_13670);
nor U14001 (N_14001,N_13059,N_13462);
and U14002 (N_14002,N_13148,N_13025);
or U14003 (N_14003,N_13395,N_13169);
nor U14004 (N_14004,N_13663,N_13932);
nor U14005 (N_14005,N_13149,N_13470);
and U14006 (N_14006,N_13558,N_13328);
xnor U14007 (N_14007,N_13875,N_13235);
nand U14008 (N_14008,N_13352,N_13814);
and U14009 (N_14009,N_13614,N_13623);
nor U14010 (N_14010,N_13868,N_13442);
or U14011 (N_14011,N_13505,N_13234);
or U14012 (N_14012,N_13602,N_13630);
or U14013 (N_14013,N_13575,N_13696);
xnor U14014 (N_14014,N_13774,N_13295);
nand U14015 (N_14015,N_13960,N_13044);
or U14016 (N_14016,N_13695,N_13921);
and U14017 (N_14017,N_13068,N_13162);
nand U14018 (N_14018,N_13142,N_13514);
xor U14019 (N_14019,N_13997,N_13970);
nand U14020 (N_14020,N_13474,N_13631);
xor U14021 (N_14021,N_13646,N_13222);
nor U14022 (N_14022,N_13746,N_13440);
and U14023 (N_14023,N_13698,N_13892);
nand U14024 (N_14024,N_13513,N_13512);
xor U14025 (N_14025,N_13040,N_13680);
and U14026 (N_14026,N_13750,N_13396);
and U14027 (N_14027,N_13361,N_13160);
nor U14028 (N_14028,N_13483,N_13290);
xnor U14029 (N_14029,N_13706,N_13246);
xnor U14030 (N_14030,N_13000,N_13096);
nor U14031 (N_14031,N_13278,N_13381);
nand U14032 (N_14032,N_13658,N_13419);
nand U14033 (N_14033,N_13820,N_13786);
or U14034 (N_14034,N_13065,N_13760);
xnor U14035 (N_14035,N_13403,N_13035);
nor U14036 (N_14036,N_13883,N_13161);
nor U14037 (N_14037,N_13109,N_13332);
nand U14038 (N_14038,N_13240,N_13218);
or U14039 (N_14039,N_13342,N_13701);
or U14040 (N_14040,N_13775,N_13668);
xor U14041 (N_14041,N_13231,N_13560);
and U14042 (N_14042,N_13117,N_13902);
and U14043 (N_14043,N_13446,N_13028);
and U14044 (N_14044,N_13020,N_13275);
xor U14045 (N_14045,N_13433,N_13432);
xnor U14046 (N_14046,N_13016,N_13785);
or U14047 (N_14047,N_13128,N_13792);
or U14048 (N_14048,N_13227,N_13485);
nand U14049 (N_14049,N_13158,N_13642);
nor U14050 (N_14050,N_13046,N_13077);
xnor U14051 (N_14051,N_13959,N_13539);
or U14052 (N_14052,N_13652,N_13681);
nand U14053 (N_14053,N_13624,N_13833);
or U14054 (N_14054,N_13209,N_13811);
nor U14055 (N_14055,N_13369,N_13769);
xnor U14056 (N_14056,N_13723,N_13302);
nor U14057 (N_14057,N_13274,N_13978);
nand U14058 (N_14058,N_13541,N_13612);
or U14059 (N_14059,N_13210,N_13859);
nand U14060 (N_14060,N_13364,N_13173);
xor U14061 (N_14061,N_13828,N_13581);
or U14062 (N_14062,N_13954,N_13186);
xor U14063 (N_14063,N_13074,N_13124);
or U14064 (N_14064,N_13480,N_13172);
nor U14065 (N_14065,N_13836,N_13365);
nor U14066 (N_14066,N_13277,N_13041);
or U14067 (N_14067,N_13490,N_13386);
nor U14068 (N_14068,N_13577,N_13551);
nand U14069 (N_14069,N_13644,N_13821);
nor U14070 (N_14070,N_13861,N_13250);
nor U14071 (N_14071,N_13003,N_13983);
nand U14072 (N_14072,N_13457,N_13191);
and U14073 (N_14073,N_13152,N_13322);
nand U14074 (N_14074,N_13633,N_13837);
or U14075 (N_14075,N_13181,N_13380);
and U14076 (N_14076,N_13586,N_13141);
nand U14077 (N_14077,N_13176,N_13076);
and U14078 (N_14078,N_13579,N_13957);
xnor U14079 (N_14079,N_13886,N_13156);
nor U14080 (N_14080,N_13654,N_13582);
nor U14081 (N_14081,N_13776,N_13098);
or U14082 (N_14082,N_13693,N_13043);
or U14083 (N_14083,N_13980,N_13420);
or U14084 (N_14084,N_13982,N_13439);
and U14085 (N_14085,N_13678,N_13280);
nor U14086 (N_14086,N_13761,N_13253);
xor U14087 (N_14087,N_13387,N_13058);
or U14088 (N_14088,N_13466,N_13832);
or U14089 (N_14089,N_13337,N_13468);
nor U14090 (N_14090,N_13784,N_13615);
and U14091 (N_14091,N_13409,N_13852);
and U14092 (N_14092,N_13824,N_13477);
xor U14093 (N_14093,N_13700,N_13800);
xnor U14094 (N_14094,N_13931,N_13516);
and U14095 (N_14095,N_13893,N_13952);
nor U14096 (N_14096,N_13896,N_13956);
xor U14097 (N_14097,N_13827,N_13242);
nor U14098 (N_14098,N_13587,N_13005);
nand U14099 (N_14099,N_13948,N_13780);
xor U14100 (N_14100,N_13282,N_13969);
or U14101 (N_14101,N_13145,N_13968);
nor U14102 (N_14102,N_13323,N_13255);
or U14103 (N_14103,N_13961,N_13618);
nor U14104 (N_14104,N_13782,N_13885);
nor U14105 (N_14105,N_13223,N_13851);
xnor U14106 (N_14106,N_13267,N_13019);
or U14107 (N_14107,N_13427,N_13854);
or U14108 (N_14108,N_13572,N_13042);
or U14109 (N_14109,N_13316,N_13350);
nand U14110 (N_14110,N_13802,N_13762);
xnor U14111 (N_14111,N_13953,N_13412);
and U14112 (N_14112,N_13989,N_13617);
and U14113 (N_14113,N_13174,N_13715);
nor U14114 (N_14114,N_13086,N_13532);
or U14115 (N_14115,N_13294,N_13378);
or U14116 (N_14116,N_13819,N_13682);
or U14117 (N_14117,N_13733,N_13276);
and U14118 (N_14118,N_13333,N_13704);
nor U14119 (N_14119,N_13125,N_13595);
nor U14120 (N_14120,N_13325,N_13258);
nor U14121 (N_14121,N_13348,N_13436);
nor U14122 (N_14122,N_13795,N_13708);
or U14123 (N_14123,N_13425,N_13745);
nor U14124 (N_14124,N_13536,N_13731);
or U14125 (N_14125,N_13229,N_13492);
and U14126 (N_14126,N_13722,N_13528);
nor U14127 (N_14127,N_13345,N_13321);
nand U14128 (N_14128,N_13026,N_13689);
xnor U14129 (N_14129,N_13180,N_13054);
xnor U14130 (N_14130,N_13224,N_13544);
xor U14131 (N_14131,N_13881,N_13647);
and U14132 (N_14132,N_13500,N_13744);
and U14133 (N_14133,N_13183,N_13263);
xor U14134 (N_14134,N_13573,N_13525);
nand U14135 (N_14135,N_13840,N_13203);
xnor U14136 (N_14136,N_13766,N_13127);
nand U14137 (N_14137,N_13106,N_13876);
nor U14138 (N_14138,N_13576,N_13661);
xor U14139 (N_14139,N_13081,N_13139);
xnor U14140 (N_14140,N_13632,N_13107);
nor U14141 (N_14141,N_13664,N_13542);
nor U14142 (N_14142,N_13371,N_13464);
xnor U14143 (N_14143,N_13199,N_13697);
or U14144 (N_14144,N_13699,N_13320);
and U14145 (N_14145,N_13600,N_13688);
nand U14146 (N_14146,N_13206,N_13606);
nor U14147 (N_14147,N_13767,N_13335);
xnor U14148 (N_14148,N_13013,N_13554);
nor U14149 (N_14149,N_13574,N_13066);
or U14150 (N_14150,N_13011,N_13626);
nor U14151 (N_14151,N_13829,N_13374);
nor U14152 (N_14152,N_13835,N_13933);
xnor U14153 (N_14153,N_13495,N_13950);
or U14154 (N_14154,N_13339,N_13373);
or U14155 (N_14155,N_13445,N_13146);
xor U14156 (N_14156,N_13928,N_13478);
xor U14157 (N_14157,N_13537,N_13341);
and U14158 (N_14158,N_13270,N_13848);
nor U14159 (N_14159,N_13356,N_13287);
and U14160 (N_14160,N_13872,N_13324);
and U14161 (N_14161,N_13069,N_13738);
xor U14162 (N_14162,N_13488,N_13676);
and U14163 (N_14163,N_13032,N_13313);
xor U14164 (N_14164,N_13591,N_13392);
or U14165 (N_14165,N_13545,N_13252);
nand U14166 (N_14166,N_13717,N_13207);
nor U14167 (N_14167,N_13414,N_13904);
and U14168 (N_14168,N_13809,N_13794);
xor U14169 (N_14169,N_13557,N_13482);
nor U14170 (N_14170,N_13400,N_13448);
nor U14171 (N_14171,N_13131,N_13383);
and U14172 (N_14172,N_13055,N_13526);
xor U14173 (N_14173,N_13362,N_13211);
and U14174 (N_14174,N_13251,N_13232);
xor U14175 (N_14175,N_13583,N_13562);
nand U14176 (N_14176,N_13165,N_13944);
nand U14177 (N_14177,N_13111,N_13771);
xor U14178 (N_14178,N_13281,N_13805);
xor U14179 (N_14179,N_13105,N_13147);
xnor U14180 (N_14180,N_13268,N_13538);
nor U14181 (N_14181,N_13164,N_13834);
or U14182 (N_14182,N_13453,N_13846);
nor U14183 (N_14183,N_13197,N_13925);
or U14184 (N_14184,N_13724,N_13552);
xnor U14185 (N_14185,N_13755,N_13079);
nor U14186 (N_14186,N_13764,N_13641);
nor U14187 (N_14187,N_13039,N_13976);
nor U14188 (N_14188,N_13789,N_13129);
nand U14189 (N_14189,N_13934,N_13728);
nand U14190 (N_14190,N_13547,N_13841);
xnor U14191 (N_14191,N_13118,N_13447);
and U14192 (N_14192,N_13057,N_13874);
and U14193 (N_14193,N_13384,N_13064);
xor U14194 (N_14194,N_13895,N_13300);
nor U14195 (N_14195,N_13645,N_13914);
nor U14196 (N_14196,N_13659,N_13807);
or U14197 (N_14197,N_13297,N_13894);
and U14198 (N_14198,N_13126,N_13977);
nand U14199 (N_14199,N_13465,N_13765);
or U14200 (N_14200,N_13912,N_13053);
nor U14201 (N_14201,N_13084,N_13006);
or U14202 (N_14202,N_13556,N_13228);
or U14203 (N_14203,N_13757,N_13790);
xnor U14204 (N_14204,N_13908,N_13882);
or U14205 (N_14205,N_13990,N_13085);
nand U14206 (N_14206,N_13429,N_13196);
nand U14207 (N_14207,N_13101,N_13018);
nor U14208 (N_14208,N_13310,N_13402);
nor U14209 (N_14209,N_13730,N_13718);
and U14210 (N_14210,N_13103,N_13877);
and U14211 (N_14211,N_13075,N_13190);
or U14212 (N_14212,N_13924,N_13571);
and U14213 (N_14213,N_13563,N_13091);
xor U14214 (N_14214,N_13388,N_13866);
and U14215 (N_14215,N_13372,N_13498);
xor U14216 (N_14216,N_13001,N_13357);
nor U14217 (N_14217,N_13692,N_13566);
xor U14218 (N_14218,N_13015,N_13946);
and U14219 (N_14219,N_13561,N_13408);
xnor U14220 (N_14220,N_13114,N_13651);
nand U14221 (N_14221,N_13534,N_13119);
or U14222 (N_14222,N_13285,N_13452);
or U14223 (N_14223,N_13411,N_13671);
or U14224 (N_14224,N_13441,N_13343);
nor U14225 (N_14225,N_13878,N_13097);
nor U14226 (N_14226,N_13201,N_13476);
xor U14227 (N_14227,N_13523,N_13330);
nor U14228 (N_14228,N_13088,N_13455);
nand U14229 (N_14229,N_13907,N_13120);
nand U14230 (N_14230,N_13812,N_13022);
nand U14231 (N_14231,N_13949,N_13753);
and U14232 (N_14232,N_13639,N_13565);
nor U14233 (N_14233,N_13208,N_13407);
and U14234 (N_14234,N_13230,N_13247);
xnor U14235 (N_14235,N_13502,N_13927);
xor U14236 (N_14236,N_13233,N_13522);
or U14237 (N_14237,N_13454,N_13175);
and U14238 (N_14238,N_13923,N_13071);
or U14239 (N_14239,N_13694,N_13569);
nor U14240 (N_14240,N_13418,N_13916);
nand U14241 (N_14241,N_13241,N_13024);
and U14242 (N_14242,N_13517,N_13986);
nor U14243 (N_14243,N_13501,N_13036);
and U14244 (N_14244,N_13340,N_13962);
xnor U14245 (N_14245,N_13375,N_13987);
nor U14246 (N_14246,N_13604,N_13917);
or U14247 (N_14247,N_13260,N_13955);
or U14248 (N_14248,N_13214,N_13702);
and U14249 (N_14249,N_13404,N_13867);
nand U14250 (N_14250,N_13014,N_13008);
xnor U14251 (N_14251,N_13354,N_13919);
or U14252 (N_14252,N_13616,N_13168);
nand U14253 (N_14253,N_13305,N_13672);
xor U14254 (N_14254,N_13423,N_13212);
nor U14255 (N_14255,N_13564,N_13416);
and U14256 (N_14256,N_13319,N_13472);
or U14257 (N_14257,N_13603,N_13585);
nand U14258 (N_14258,N_13179,N_13047);
and U14259 (N_14259,N_13810,N_13685);
xor U14260 (N_14260,N_13506,N_13435);
and U14261 (N_14261,N_13239,N_13653);
nand U14262 (N_14262,N_13338,N_13622);
nor U14263 (N_14263,N_13494,N_13100);
xnor U14264 (N_14264,N_13625,N_13479);
and U14265 (N_14265,N_13817,N_13519);
xnor U14266 (N_14266,N_13673,N_13437);
or U14267 (N_14267,N_13958,N_13690);
xnor U14268 (N_14268,N_13216,N_13655);
nand U14269 (N_14269,N_13930,N_13463);
xor U14270 (N_14270,N_13748,N_13911);
nand U14271 (N_14271,N_13507,N_13449);
or U14272 (N_14272,N_13844,N_13598);
or U14273 (N_14273,N_13888,N_13903);
xnor U14274 (N_14274,N_13326,N_13570);
xor U14275 (N_14275,N_13467,N_13002);
nand U14276 (N_14276,N_13543,N_13823);
nand U14277 (N_14277,N_13284,N_13359);
nor U14278 (N_14278,N_13660,N_13808);
and U14279 (N_14279,N_13458,N_13797);
or U14280 (N_14280,N_13461,N_13918);
nand U14281 (N_14281,N_13306,N_13004);
nor U14282 (N_14282,N_13596,N_13862);
or U14283 (N_14283,N_13801,N_13635);
nand U14284 (N_14284,N_13499,N_13845);
and U14285 (N_14285,N_13864,N_13311);
or U14286 (N_14286,N_13988,N_13189);
nand U14287 (N_14287,N_13758,N_13010);
xor U14288 (N_14288,N_13971,N_13677);
and U14289 (N_14289,N_13226,N_13609);
nand U14290 (N_14290,N_13742,N_13707);
nand U14291 (N_14291,N_13714,N_13225);
and U14292 (N_14292,N_13346,N_13589);
xor U14293 (N_14293,N_13051,N_13727);
and U14294 (N_14294,N_13890,N_13353);
or U14295 (N_14295,N_13607,N_13710);
nor U14296 (N_14296,N_13734,N_13122);
and U14297 (N_14297,N_13301,N_13390);
xor U14298 (N_14298,N_13291,N_13999);
and U14299 (N_14299,N_13264,N_13567);
nor U14300 (N_14300,N_13703,N_13711);
nor U14301 (N_14301,N_13674,N_13666);
nor U14302 (N_14302,N_13743,N_13087);
nand U14303 (N_14303,N_13497,N_13627);
nor U14304 (N_14304,N_13972,N_13398);
nand U14305 (N_14305,N_13597,N_13308);
nor U14306 (N_14306,N_13279,N_13740);
nor U14307 (N_14307,N_13130,N_13818);
or U14308 (N_14308,N_13336,N_13344);
nor U14309 (N_14309,N_13965,N_13858);
and U14310 (N_14310,N_13092,N_13768);
or U14311 (N_14311,N_13050,N_13082);
nand U14312 (N_14312,N_13116,N_13590);
nand U14313 (N_14313,N_13729,N_13102);
xnor U14314 (N_14314,N_13177,N_13108);
or U14315 (N_14315,N_13679,N_13192);
and U14316 (N_14316,N_13049,N_13150);
xnor U14317 (N_14317,N_13033,N_13273);
nor U14318 (N_14318,N_13038,N_13220);
nand U14319 (N_14319,N_13620,N_13842);
nor U14320 (N_14320,N_13481,N_13611);
xnor U14321 (N_14321,N_13629,N_13580);
and U14322 (N_14322,N_13721,N_13136);
and U14323 (N_14323,N_13428,N_13099);
nand U14324 (N_14324,N_13469,N_13331);
and U14325 (N_14325,N_13601,N_13796);
xor U14326 (N_14326,N_13613,N_13593);
or U14327 (N_14327,N_13656,N_13843);
and U14328 (N_14328,N_13104,N_13363);
and U14329 (N_14329,N_13935,N_13559);
and U14330 (N_14330,N_13838,N_13110);
and U14331 (N_14331,N_13521,N_13393);
xor U14332 (N_14332,N_13546,N_13473);
xnor U14333 (N_14333,N_13610,N_13397);
or U14334 (N_14334,N_13889,N_13998);
nor U14335 (N_14335,N_13315,N_13993);
nor U14336 (N_14336,N_13286,N_13424);
xor U14337 (N_14337,N_13184,N_13863);
xnor U14338 (N_14338,N_13687,N_13080);
xnor U14339 (N_14339,N_13157,N_13806);
and U14340 (N_14340,N_13256,N_13456);
xnor U14341 (N_14341,N_13984,N_13996);
or U14342 (N_14342,N_13317,N_13493);
or U14343 (N_14343,N_13849,N_13078);
nand U14344 (N_14344,N_13856,N_13860);
xor U14345 (N_14345,N_13045,N_13029);
xnor U14346 (N_14346,N_13739,N_13410);
nand U14347 (N_14347,N_13847,N_13549);
and U14348 (N_14348,N_13072,N_13134);
or U14349 (N_14349,N_13265,N_13347);
nor U14350 (N_14350,N_13178,N_13995);
nand U14351 (N_14351,N_13822,N_13599);
and U14352 (N_14352,N_13634,N_13204);
nand U14353 (N_14353,N_13777,N_13638);
nor U14354 (N_14354,N_13531,N_13471);
nand U14355 (N_14355,N_13853,N_13816);
nor U14356 (N_14356,N_13073,N_13399);
nor U14357 (N_14357,N_13027,N_13568);
nor U14358 (N_14358,N_13636,N_13171);
nand U14359 (N_14359,N_13056,N_13299);
xor U14360 (N_14360,N_13803,N_13459);
and U14361 (N_14361,N_13870,N_13289);
xnor U14362 (N_14362,N_13248,N_13669);
xnor U14363 (N_14363,N_13030,N_13370);
nor U14364 (N_14364,N_13747,N_13377);
or U14365 (N_14365,N_13787,N_13113);
xnor U14366 (N_14366,N_13391,N_13530);
nand U14367 (N_14367,N_13401,N_13063);
xor U14368 (N_14368,N_13304,N_13608);
xor U14369 (N_14369,N_13675,N_13548);
nand U14370 (N_14370,N_13713,N_13358);
nand U14371 (N_14371,N_13185,N_13198);
nand U14372 (N_14372,N_13550,N_13298);
or U14373 (N_14373,N_13637,N_13182);
nand U14374 (N_14374,N_13154,N_13737);
nor U14375 (N_14375,N_13444,N_13756);
xor U14376 (N_14376,N_13272,N_13155);
nor U14377 (N_14377,N_13665,N_13389);
nor U14378 (N_14378,N_13245,N_13773);
xor U14379 (N_14379,N_13520,N_13947);
nand U14380 (N_14380,N_13657,N_13060);
or U14381 (N_14381,N_13244,N_13451);
nand U14382 (N_14382,N_13791,N_13249);
nand U14383 (N_14383,N_13804,N_13385);
nand U14384 (N_14384,N_13938,N_13307);
or U14385 (N_14385,N_13799,N_13132);
or U14386 (N_14386,N_13187,N_13712);
xor U14387 (N_14387,N_13188,N_13351);
nand U14388 (N_14388,N_13865,N_13779);
xnor U14389 (N_14389,N_13112,N_13553);
or U14390 (N_14390,N_13269,N_13318);
and U14391 (N_14391,N_13394,N_13138);
and U14392 (N_14392,N_13735,N_13292);
nand U14393 (N_14393,N_13850,N_13508);
nand U14394 (N_14394,N_13535,N_13144);
xnor U14395 (N_14395,N_13070,N_13509);
nor U14396 (N_14396,N_13605,N_13941);
nand U14397 (N_14397,N_13426,N_13009);
and U14398 (N_14398,N_13510,N_13720);
nor U14399 (N_14399,N_13621,N_13966);
nand U14400 (N_14400,N_13592,N_13588);
xor U14401 (N_14401,N_13376,N_13314);
xnor U14402 (N_14402,N_13662,N_13221);
and U14403 (N_14403,N_13417,N_13936);
and U14404 (N_14404,N_13140,N_13151);
nor U14405 (N_14405,N_13891,N_13012);
or U14406 (N_14406,N_13257,N_13855);
nor U14407 (N_14407,N_13871,N_13413);
xor U14408 (N_14408,N_13684,N_13309);
nand U14409 (N_14409,N_13193,N_13533);
nor U14410 (N_14410,N_13839,N_13783);
xor U14411 (N_14411,N_13052,N_13994);
and U14412 (N_14412,N_13926,N_13382);
and U14413 (N_14413,N_13741,N_13491);
nand U14414 (N_14414,N_13899,N_13649);
and U14415 (N_14415,N_13238,N_13167);
nand U14416 (N_14416,N_13975,N_13643);
nand U14417 (N_14417,N_13686,N_13061);
nand U14418 (N_14418,N_13213,N_13974);
xor U14419 (N_14419,N_13062,N_13985);
and U14420 (N_14420,N_13137,N_13754);
and U14421 (N_14421,N_13202,N_13725);
or U14422 (N_14422,N_13143,N_13450);
nor U14423 (N_14423,N_13798,N_13489);
nor U14424 (N_14424,N_13529,N_13123);
nand U14425 (N_14425,N_13527,N_13170);
nand U14426 (N_14426,N_13288,N_13312);
xor U14427 (N_14427,N_13778,N_13431);
xnor U14428 (N_14428,N_13628,N_13496);
nor U14429 (N_14429,N_13475,N_13825);
or U14430 (N_14430,N_13619,N_13772);
and U14431 (N_14431,N_13254,N_13940);
or U14432 (N_14432,N_13486,N_13716);
xor U14433 (N_14433,N_13815,N_13094);
nor U14434 (N_14434,N_13992,N_13217);
xnor U14435 (N_14435,N_13034,N_13135);
and U14436 (N_14436,N_13909,N_13751);
nand U14437 (N_14437,N_13963,N_13503);
xnor U14438 (N_14438,N_13913,N_13945);
nand U14439 (N_14439,N_13887,N_13266);
or U14440 (N_14440,N_13705,N_13089);
nand U14441 (N_14441,N_13973,N_13195);
and U14442 (N_14442,N_13283,N_13857);
nand U14443 (N_14443,N_13200,N_13083);
nor U14444 (N_14444,N_13732,N_13991);
nand U14445 (N_14445,N_13271,N_13910);
and U14446 (N_14446,N_13578,N_13379);
and U14447 (N_14447,N_13243,N_13021);
nor U14448 (N_14448,N_13367,N_13540);
nor U14449 (N_14449,N_13770,N_13906);
and U14450 (N_14450,N_13095,N_13219);
or U14451 (N_14451,N_13942,N_13115);
and U14452 (N_14452,N_13900,N_13434);
xor U14453 (N_14453,N_13979,N_13293);
nor U14454 (N_14454,N_13422,N_13133);
xor U14455 (N_14455,N_13460,N_13366);
xnor U14456 (N_14456,N_13236,N_13967);
and U14457 (N_14457,N_13901,N_13421);
xnor U14458 (N_14458,N_13943,N_13939);
and U14459 (N_14459,N_13726,N_13898);
nor U14460 (N_14460,N_13905,N_13261);
nor U14461 (N_14461,N_13262,N_13159);
xor U14462 (N_14462,N_13487,N_13484);
xnor U14463 (N_14463,N_13869,N_13884);
nor U14464 (N_14464,N_13915,N_13215);
nor U14465 (N_14465,N_13736,N_13719);
nor U14466 (N_14466,N_13880,N_13920);
xor U14467 (N_14467,N_13121,N_13438);
xnor U14468 (N_14468,N_13831,N_13524);
nor U14469 (N_14469,N_13048,N_13406);
nor U14470 (N_14470,N_13007,N_13709);
and U14471 (N_14471,N_13415,N_13518);
or U14472 (N_14472,N_13922,N_13329);
nand U14473 (N_14473,N_13826,N_13093);
nor U14474 (N_14474,N_13511,N_13683);
xnor U14475 (N_14475,N_13752,N_13640);
and U14476 (N_14476,N_13349,N_13023);
and U14477 (N_14477,N_13691,N_13237);
nor U14478 (N_14478,N_13296,N_13937);
xor U14479 (N_14479,N_13334,N_13153);
xnor U14480 (N_14480,N_13759,N_13443);
and U14481 (N_14481,N_13430,N_13327);
and U14482 (N_14482,N_13031,N_13981);
nand U14483 (N_14483,N_13594,N_13667);
nor U14484 (N_14484,N_13897,N_13163);
xnor U14485 (N_14485,N_13405,N_13355);
nand U14486 (N_14486,N_13205,N_13648);
and U14487 (N_14487,N_13555,N_13515);
nor U14488 (N_14488,N_13368,N_13650);
nor U14489 (N_14489,N_13749,N_13813);
nor U14490 (N_14490,N_13879,N_13303);
nor U14491 (N_14491,N_13166,N_13090);
or U14492 (N_14492,N_13017,N_13788);
or U14493 (N_14493,N_13194,N_13504);
and U14494 (N_14494,N_13951,N_13584);
xnor U14495 (N_14495,N_13929,N_13793);
xnor U14496 (N_14496,N_13037,N_13259);
nand U14497 (N_14497,N_13830,N_13067);
or U14498 (N_14498,N_13964,N_13873);
xnor U14499 (N_14499,N_13781,N_13763);
xor U14500 (N_14500,N_13861,N_13559);
nor U14501 (N_14501,N_13621,N_13169);
nor U14502 (N_14502,N_13106,N_13681);
and U14503 (N_14503,N_13209,N_13020);
and U14504 (N_14504,N_13238,N_13518);
nand U14505 (N_14505,N_13020,N_13232);
nand U14506 (N_14506,N_13875,N_13935);
nand U14507 (N_14507,N_13101,N_13411);
or U14508 (N_14508,N_13642,N_13187);
or U14509 (N_14509,N_13393,N_13626);
nor U14510 (N_14510,N_13796,N_13711);
nor U14511 (N_14511,N_13864,N_13705);
nor U14512 (N_14512,N_13460,N_13059);
and U14513 (N_14513,N_13124,N_13433);
and U14514 (N_14514,N_13926,N_13170);
or U14515 (N_14515,N_13704,N_13875);
nand U14516 (N_14516,N_13357,N_13233);
and U14517 (N_14517,N_13880,N_13277);
nand U14518 (N_14518,N_13852,N_13102);
xnor U14519 (N_14519,N_13558,N_13887);
and U14520 (N_14520,N_13873,N_13445);
nand U14521 (N_14521,N_13619,N_13902);
or U14522 (N_14522,N_13433,N_13285);
xnor U14523 (N_14523,N_13985,N_13933);
or U14524 (N_14524,N_13204,N_13933);
xor U14525 (N_14525,N_13226,N_13334);
xor U14526 (N_14526,N_13221,N_13816);
xor U14527 (N_14527,N_13323,N_13954);
or U14528 (N_14528,N_13827,N_13445);
and U14529 (N_14529,N_13395,N_13398);
nor U14530 (N_14530,N_13213,N_13900);
nand U14531 (N_14531,N_13150,N_13641);
or U14532 (N_14532,N_13522,N_13784);
and U14533 (N_14533,N_13201,N_13899);
nand U14534 (N_14534,N_13217,N_13043);
or U14535 (N_14535,N_13872,N_13380);
nand U14536 (N_14536,N_13027,N_13855);
nand U14537 (N_14537,N_13159,N_13858);
nor U14538 (N_14538,N_13308,N_13846);
or U14539 (N_14539,N_13572,N_13649);
nand U14540 (N_14540,N_13727,N_13610);
and U14541 (N_14541,N_13015,N_13393);
nor U14542 (N_14542,N_13002,N_13846);
xnor U14543 (N_14543,N_13944,N_13455);
or U14544 (N_14544,N_13472,N_13786);
nor U14545 (N_14545,N_13092,N_13639);
xor U14546 (N_14546,N_13912,N_13454);
and U14547 (N_14547,N_13707,N_13255);
or U14548 (N_14548,N_13328,N_13072);
nand U14549 (N_14549,N_13765,N_13518);
and U14550 (N_14550,N_13594,N_13766);
and U14551 (N_14551,N_13547,N_13903);
or U14552 (N_14552,N_13343,N_13088);
nand U14553 (N_14553,N_13046,N_13348);
nand U14554 (N_14554,N_13901,N_13819);
nand U14555 (N_14555,N_13821,N_13342);
xor U14556 (N_14556,N_13685,N_13584);
nor U14557 (N_14557,N_13880,N_13232);
or U14558 (N_14558,N_13185,N_13249);
nand U14559 (N_14559,N_13552,N_13284);
nand U14560 (N_14560,N_13771,N_13207);
xor U14561 (N_14561,N_13047,N_13990);
nor U14562 (N_14562,N_13688,N_13552);
or U14563 (N_14563,N_13110,N_13460);
nor U14564 (N_14564,N_13359,N_13819);
nand U14565 (N_14565,N_13245,N_13173);
and U14566 (N_14566,N_13038,N_13851);
xnor U14567 (N_14567,N_13105,N_13437);
xor U14568 (N_14568,N_13721,N_13550);
and U14569 (N_14569,N_13289,N_13821);
nor U14570 (N_14570,N_13202,N_13210);
nand U14571 (N_14571,N_13148,N_13494);
xnor U14572 (N_14572,N_13280,N_13534);
or U14573 (N_14573,N_13594,N_13017);
nand U14574 (N_14574,N_13988,N_13206);
nand U14575 (N_14575,N_13518,N_13298);
nor U14576 (N_14576,N_13277,N_13487);
and U14577 (N_14577,N_13094,N_13680);
and U14578 (N_14578,N_13998,N_13659);
nand U14579 (N_14579,N_13199,N_13299);
nand U14580 (N_14580,N_13436,N_13705);
and U14581 (N_14581,N_13322,N_13719);
or U14582 (N_14582,N_13784,N_13827);
xnor U14583 (N_14583,N_13485,N_13835);
or U14584 (N_14584,N_13849,N_13386);
or U14585 (N_14585,N_13761,N_13497);
xor U14586 (N_14586,N_13868,N_13365);
xnor U14587 (N_14587,N_13329,N_13512);
and U14588 (N_14588,N_13777,N_13741);
nor U14589 (N_14589,N_13117,N_13434);
or U14590 (N_14590,N_13061,N_13715);
nor U14591 (N_14591,N_13736,N_13201);
nand U14592 (N_14592,N_13385,N_13664);
and U14593 (N_14593,N_13043,N_13416);
or U14594 (N_14594,N_13575,N_13785);
or U14595 (N_14595,N_13532,N_13440);
and U14596 (N_14596,N_13324,N_13089);
or U14597 (N_14597,N_13021,N_13049);
xnor U14598 (N_14598,N_13723,N_13343);
or U14599 (N_14599,N_13033,N_13350);
or U14600 (N_14600,N_13401,N_13079);
or U14601 (N_14601,N_13786,N_13031);
nand U14602 (N_14602,N_13119,N_13797);
or U14603 (N_14603,N_13347,N_13522);
nand U14604 (N_14604,N_13548,N_13493);
xnor U14605 (N_14605,N_13154,N_13779);
nand U14606 (N_14606,N_13023,N_13462);
or U14607 (N_14607,N_13038,N_13294);
nor U14608 (N_14608,N_13248,N_13832);
nor U14609 (N_14609,N_13250,N_13991);
and U14610 (N_14610,N_13454,N_13326);
and U14611 (N_14611,N_13793,N_13676);
xnor U14612 (N_14612,N_13623,N_13504);
and U14613 (N_14613,N_13932,N_13310);
and U14614 (N_14614,N_13860,N_13155);
nor U14615 (N_14615,N_13538,N_13807);
xnor U14616 (N_14616,N_13545,N_13400);
nor U14617 (N_14617,N_13215,N_13236);
or U14618 (N_14618,N_13396,N_13065);
nor U14619 (N_14619,N_13034,N_13543);
xnor U14620 (N_14620,N_13836,N_13733);
and U14621 (N_14621,N_13063,N_13810);
xnor U14622 (N_14622,N_13964,N_13593);
nor U14623 (N_14623,N_13054,N_13936);
nor U14624 (N_14624,N_13472,N_13588);
nor U14625 (N_14625,N_13662,N_13401);
or U14626 (N_14626,N_13329,N_13041);
nand U14627 (N_14627,N_13619,N_13294);
and U14628 (N_14628,N_13643,N_13572);
xor U14629 (N_14629,N_13084,N_13302);
and U14630 (N_14630,N_13996,N_13315);
nor U14631 (N_14631,N_13560,N_13770);
nand U14632 (N_14632,N_13877,N_13778);
and U14633 (N_14633,N_13879,N_13019);
and U14634 (N_14634,N_13320,N_13710);
and U14635 (N_14635,N_13541,N_13443);
nor U14636 (N_14636,N_13785,N_13204);
nor U14637 (N_14637,N_13095,N_13854);
nand U14638 (N_14638,N_13701,N_13560);
or U14639 (N_14639,N_13657,N_13095);
and U14640 (N_14640,N_13410,N_13829);
nor U14641 (N_14641,N_13553,N_13627);
and U14642 (N_14642,N_13676,N_13375);
nor U14643 (N_14643,N_13852,N_13331);
xor U14644 (N_14644,N_13039,N_13179);
nor U14645 (N_14645,N_13120,N_13284);
or U14646 (N_14646,N_13190,N_13076);
nor U14647 (N_14647,N_13365,N_13338);
nor U14648 (N_14648,N_13909,N_13685);
or U14649 (N_14649,N_13520,N_13223);
xnor U14650 (N_14650,N_13935,N_13402);
xor U14651 (N_14651,N_13886,N_13033);
or U14652 (N_14652,N_13159,N_13041);
nor U14653 (N_14653,N_13947,N_13210);
nor U14654 (N_14654,N_13203,N_13100);
and U14655 (N_14655,N_13079,N_13509);
nor U14656 (N_14656,N_13210,N_13224);
nor U14657 (N_14657,N_13513,N_13661);
nor U14658 (N_14658,N_13556,N_13270);
nand U14659 (N_14659,N_13279,N_13080);
xnor U14660 (N_14660,N_13587,N_13323);
nand U14661 (N_14661,N_13843,N_13760);
nor U14662 (N_14662,N_13812,N_13773);
nand U14663 (N_14663,N_13540,N_13229);
or U14664 (N_14664,N_13257,N_13908);
nor U14665 (N_14665,N_13716,N_13984);
nor U14666 (N_14666,N_13613,N_13958);
nor U14667 (N_14667,N_13432,N_13054);
and U14668 (N_14668,N_13322,N_13147);
and U14669 (N_14669,N_13192,N_13950);
nor U14670 (N_14670,N_13231,N_13859);
or U14671 (N_14671,N_13279,N_13287);
nand U14672 (N_14672,N_13168,N_13782);
or U14673 (N_14673,N_13841,N_13534);
xor U14674 (N_14674,N_13446,N_13305);
nand U14675 (N_14675,N_13949,N_13790);
nand U14676 (N_14676,N_13875,N_13700);
or U14677 (N_14677,N_13272,N_13474);
xor U14678 (N_14678,N_13589,N_13649);
and U14679 (N_14679,N_13264,N_13854);
or U14680 (N_14680,N_13618,N_13016);
or U14681 (N_14681,N_13189,N_13758);
nand U14682 (N_14682,N_13721,N_13602);
xor U14683 (N_14683,N_13857,N_13194);
and U14684 (N_14684,N_13444,N_13990);
and U14685 (N_14685,N_13308,N_13490);
nor U14686 (N_14686,N_13945,N_13820);
and U14687 (N_14687,N_13067,N_13475);
nand U14688 (N_14688,N_13661,N_13385);
nor U14689 (N_14689,N_13561,N_13655);
and U14690 (N_14690,N_13244,N_13418);
and U14691 (N_14691,N_13897,N_13936);
xor U14692 (N_14692,N_13672,N_13207);
or U14693 (N_14693,N_13569,N_13510);
nor U14694 (N_14694,N_13849,N_13006);
nand U14695 (N_14695,N_13121,N_13277);
nand U14696 (N_14696,N_13904,N_13542);
nor U14697 (N_14697,N_13998,N_13932);
xor U14698 (N_14698,N_13878,N_13972);
and U14699 (N_14699,N_13513,N_13108);
nand U14700 (N_14700,N_13308,N_13722);
or U14701 (N_14701,N_13667,N_13644);
xor U14702 (N_14702,N_13614,N_13681);
xnor U14703 (N_14703,N_13113,N_13729);
or U14704 (N_14704,N_13731,N_13107);
and U14705 (N_14705,N_13975,N_13394);
xnor U14706 (N_14706,N_13064,N_13518);
and U14707 (N_14707,N_13327,N_13207);
and U14708 (N_14708,N_13008,N_13749);
xor U14709 (N_14709,N_13581,N_13831);
nor U14710 (N_14710,N_13251,N_13235);
nor U14711 (N_14711,N_13738,N_13199);
or U14712 (N_14712,N_13768,N_13941);
xor U14713 (N_14713,N_13969,N_13996);
nor U14714 (N_14714,N_13427,N_13286);
nor U14715 (N_14715,N_13437,N_13148);
nand U14716 (N_14716,N_13476,N_13081);
or U14717 (N_14717,N_13468,N_13893);
nor U14718 (N_14718,N_13609,N_13705);
xnor U14719 (N_14719,N_13967,N_13008);
nand U14720 (N_14720,N_13383,N_13804);
nand U14721 (N_14721,N_13209,N_13480);
xor U14722 (N_14722,N_13733,N_13970);
or U14723 (N_14723,N_13776,N_13531);
nand U14724 (N_14724,N_13224,N_13829);
nand U14725 (N_14725,N_13792,N_13156);
nand U14726 (N_14726,N_13849,N_13122);
nand U14727 (N_14727,N_13708,N_13398);
or U14728 (N_14728,N_13134,N_13654);
and U14729 (N_14729,N_13443,N_13582);
and U14730 (N_14730,N_13265,N_13928);
xnor U14731 (N_14731,N_13720,N_13880);
and U14732 (N_14732,N_13839,N_13280);
or U14733 (N_14733,N_13338,N_13876);
or U14734 (N_14734,N_13924,N_13373);
nand U14735 (N_14735,N_13347,N_13780);
and U14736 (N_14736,N_13406,N_13373);
xnor U14737 (N_14737,N_13113,N_13070);
nor U14738 (N_14738,N_13929,N_13825);
nor U14739 (N_14739,N_13239,N_13306);
or U14740 (N_14740,N_13839,N_13232);
nand U14741 (N_14741,N_13229,N_13623);
nor U14742 (N_14742,N_13509,N_13835);
nand U14743 (N_14743,N_13838,N_13237);
and U14744 (N_14744,N_13176,N_13348);
nor U14745 (N_14745,N_13276,N_13041);
nor U14746 (N_14746,N_13477,N_13128);
or U14747 (N_14747,N_13126,N_13849);
and U14748 (N_14748,N_13856,N_13976);
or U14749 (N_14749,N_13840,N_13990);
or U14750 (N_14750,N_13173,N_13598);
xnor U14751 (N_14751,N_13383,N_13743);
or U14752 (N_14752,N_13890,N_13720);
and U14753 (N_14753,N_13121,N_13989);
xnor U14754 (N_14754,N_13866,N_13223);
nor U14755 (N_14755,N_13384,N_13477);
or U14756 (N_14756,N_13217,N_13662);
nor U14757 (N_14757,N_13021,N_13998);
nor U14758 (N_14758,N_13482,N_13148);
and U14759 (N_14759,N_13958,N_13665);
and U14760 (N_14760,N_13123,N_13252);
nor U14761 (N_14761,N_13342,N_13925);
xor U14762 (N_14762,N_13687,N_13219);
nand U14763 (N_14763,N_13753,N_13328);
nand U14764 (N_14764,N_13041,N_13929);
and U14765 (N_14765,N_13216,N_13858);
and U14766 (N_14766,N_13851,N_13594);
nor U14767 (N_14767,N_13444,N_13025);
xor U14768 (N_14768,N_13130,N_13052);
or U14769 (N_14769,N_13300,N_13015);
and U14770 (N_14770,N_13706,N_13492);
nor U14771 (N_14771,N_13971,N_13065);
and U14772 (N_14772,N_13418,N_13334);
xor U14773 (N_14773,N_13920,N_13949);
nand U14774 (N_14774,N_13614,N_13413);
nand U14775 (N_14775,N_13269,N_13691);
and U14776 (N_14776,N_13419,N_13535);
xnor U14777 (N_14777,N_13820,N_13589);
and U14778 (N_14778,N_13441,N_13149);
nor U14779 (N_14779,N_13393,N_13602);
xor U14780 (N_14780,N_13486,N_13345);
or U14781 (N_14781,N_13315,N_13496);
and U14782 (N_14782,N_13040,N_13876);
nor U14783 (N_14783,N_13334,N_13922);
nor U14784 (N_14784,N_13852,N_13013);
and U14785 (N_14785,N_13796,N_13393);
or U14786 (N_14786,N_13514,N_13284);
nand U14787 (N_14787,N_13477,N_13867);
nor U14788 (N_14788,N_13789,N_13656);
xor U14789 (N_14789,N_13635,N_13841);
and U14790 (N_14790,N_13529,N_13518);
nor U14791 (N_14791,N_13726,N_13164);
nor U14792 (N_14792,N_13513,N_13352);
or U14793 (N_14793,N_13159,N_13811);
nor U14794 (N_14794,N_13457,N_13741);
nand U14795 (N_14795,N_13580,N_13584);
or U14796 (N_14796,N_13644,N_13783);
or U14797 (N_14797,N_13152,N_13757);
and U14798 (N_14798,N_13100,N_13514);
nor U14799 (N_14799,N_13011,N_13180);
xnor U14800 (N_14800,N_13206,N_13945);
xnor U14801 (N_14801,N_13504,N_13248);
xor U14802 (N_14802,N_13508,N_13812);
nand U14803 (N_14803,N_13159,N_13562);
and U14804 (N_14804,N_13713,N_13961);
and U14805 (N_14805,N_13548,N_13680);
nand U14806 (N_14806,N_13542,N_13145);
and U14807 (N_14807,N_13788,N_13162);
xnor U14808 (N_14808,N_13694,N_13053);
and U14809 (N_14809,N_13051,N_13111);
nand U14810 (N_14810,N_13421,N_13964);
and U14811 (N_14811,N_13593,N_13320);
nor U14812 (N_14812,N_13646,N_13339);
nor U14813 (N_14813,N_13260,N_13111);
or U14814 (N_14814,N_13863,N_13550);
or U14815 (N_14815,N_13607,N_13769);
or U14816 (N_14816,N_13022,N_13310);
or U14817 (N_14817,N_13764,N_13117);
and U14818 (N_14818,N_13777,N_13625);
and U14819 (N_14819,N_13445,N_13440);
nor U14820 (N_14820,N_13821,N_13129);
nand U14821 (N_14821,N_13562,N_13473);
xor U14822 (N_14822,N_13506,N_13885);
nor U14823 (N_14823,N_13968,N_13608);
or U14824 (N_14824,N_13675,N_13683);
and U14825 (N_14825,N_13441,N_13017);
and U14826 (N_14826,N_13951,N_13825);
nor U14827 (N_14827,N_13269,N_13188);
or U14828 (N_14828,N_13124,N_13827);
xnor U14829 (N_14829,N_13755,N_13153);
xnor U14830 (N_14830,N_13525,N_13132);
xor U14831 (N_14831,N_13640,N_13731);
nand U14832 (N_14832,N_13417,N_13361);
or U14833 (N_14833,N_13155,N_13645);
nor U14834 (N_14834,N_13765,N_13495);
xor U14835 (N_14835,N_13928,N_13804);
and U14836 (N_14836,N_13147,N_13283);
nand U14837 (N_14837,N_13553,N_13615);
and U14838 (N_14838,N_13414,N_13310);
or U14839 (N_14839,N_13290,N_13535);
nor U14840 (N_14840,N_13920,N_13600);
xnor U14841 (N_14841,N_13332,N_13690);
and U14842 (N_14842,N_13964,N_13971);
or U14843 (N_14843,N_13811,N_13124);
nor U14844 (N_14844,N_13286,N_13673);
nor U14845 (N_14845,N_13502,N_13115);
nor U14846 (N_14846,N_13546,N_13489);
xnor U14847 (N_14847,N_13500,N_13617);
xor U14848 (N_14848,N_13974,N_13980);
nand U14849 (N_14849,N_13777,N_13681);
nand U14850 (N_14850,N_13656,N_13376);
nand U14851 (N_14851,N_13062,N_13341);
nand U14852 (N_14852,N_13994,N_13017);
and U14853 (N_14853,N_13549,N_13607);
or U14854 (N_14854,N_13710,N_13916);
nor U14855 (N_14855,N_13816,N_13383);
nor U14856 (N_14856,N_13719,N_13151);
nand U14857 (N_14857,N_13241,N_13360);
and U14858 (N_14858,N_13484,N_13486);
nand U14859 (N_14859,N_13088,N_13479);
and U14860 (N_14860,N_13007,N_13689);
xor U14861 (N_14861,N_13666,N_13702);
xnor U14862 (N_14862,N_13798,N_13378);
nand U14863 (N_14863,N_13430,N_13406);
xor U14864 (N_14864,N_13008,N_13908);
and U14865 (N_14865,N_13706,N_13043);
and U14866 (N_14866,N_13389,N_13639);
nor U14867 (N_14867,N_13127,N_13698);
and U14868 (N_14868,N_13811,N_13568);
xnor U14869 (N_14869,N_13174,N_13777);
nor U14870 (N_14870,N_13997,N_13602);
xor U14871 (N_14871,N_13106,N_13630);
nand U14872 (N_14872,N_13228,N_13361);
xor U14873 (N_14873,N_13967,N_13316);
xnor U14874 (N_14874,N_13094,N_13981);
xnor U14875 (N_14875,N_13797,N_13230);
nand U14876 (N_14876,N_13694,N_13317);
and U14877 (N_14877,N_13528,N_13213);
and U14878 (N_14878,N_13345,N_13260);
or U14879 (N_14879,N_13577,N_13122);
nor U14880 (N_14880,N_13461,N_13257);
nor U14881 (N_14881,N_13205,N_13813);
or U14882 (N_14882,N_13017,N_13857);
nor U14883 (N_14883,N_13645,N_13898);
xor U14884 (N_14884,N_13981,N_13326);
or U14885 (N_14885,N_13844,N_13147);
xor U14886 (N_14886,N_13433,N_13816);
xnor U14887 (N_14887,N_13051,N_13297);
nand U14888 (N_14888,N_13339,N_13329);
nor U14889 (N_14889,N_13496,N_13073);
nand U14890 (N_14890,N_13631,N_13129);
nand U14891 (N_14891,N_13769,N_13034);
or U14892 (N_14892,N_13837,N_13372);
and U14893 (N_14893,N_13510,N_13567);
xnor U14894 (N_14894,N_13511,N_13857);
or U14895 (N_14895,N_13127,N_13401);
and U14896 (N_14896,N_13060,N_13363);
nand U14897 (N_14897,N_13826,N_13773);
nand U14898 (N_14898,N_13624,N_13537);
xnor U14899 (N_14899,N_13668,N_13135);
or U14900 (N_14900,N_13419,N_13092);
nor U14901 (N_14901,N_13071,N_13723);
and U14902 (N_14902,N_13724,N_13924);
and U14903 (N_14903,N_13154,N_13386);
nor U14904 (N_14904,N_13408,N_13194);
and U14905 (N_14905,N_13101,N_13463);
nor U14906 (N_14906,N_13980,N_13474);
xnor U14907 (N_14907,N_13678,N_13035);
and U14908 (N_14908,N_13961,N_13168);
nor U14909 (N_14909,N_13784,N_13760);
and U14910 (N_14910,N_13496,N_13204);
nor U14911 (N_14911,N_13005,N_13337);
or U14912 (N_14912,N_13178,N_13608);
nand U14913 (N_14913,N_13905,N_13224);
or U14914 (N_14914,N_13595,N_13068);
and U14915 (N_14915,N_13727,N_13615);
xor U14916 (N_14916,N_13988,N_13170);
nor U14917 (N_14917,N_13947,N_13761);
or U14918 (N_14918,N_13093,N_13858);
nand U14919 (N_14919,N_13244,N_13934);
or U14920 (N_14920,N_13589,N_13282);
nor U14921 (N_14921,N_13093,N_13085);
nand U14922 (N_14922,N_13139,N_13312);
or U14923 (N_14923,N_13441,N_13278);
nand U14924 (N_14924,N_13696,N_13915);
or U14925 (N_14925,N_13835,N_13823);
or U14926 (N_14926,N_13397,N_13066);
and U14927 (N_14927,N_13130,N_13600);
xor U14928 (N_14928,N_13305,N_13977);
and U14929 (N_14929,N_13806,N_13011);
nor U14930 (N_14930,N_13963,N_13036);
and U14931 (N_14931,N_13185,N_13159);
nand U14932 (N_14932,N_13485,N_13202);
xnor U14933 (N_14933,N_13179,N_13144);
or U14934 (N_14934,N_13146,N_13556);
nor U14935 (N_14935,N_13488,N_13077);
nand U14936 (N_14936,N_13973,N_13344);
xor U14937 (N_14937,N_13880,N_13784);
xor U14938 (N_14938,N_13054,N_13002);
or U14939 (N_14939,N_13923,N_13661);
or U14940 (N_14940,N_13101,N_13867);
nand U14941 (N_14941,N_13080,N_13511);
xnor U14942 (N_14942,N_13187,N_13665);
nand U14943 (N_14943,N_13065,N_13578);
and U14944 (N_14944,N_13485,N_13744);
nor U14945 (N_14945,N_13915,N_13023);
and U14946 (N_14946,N_13493,N_13183);
or U14947 (N_14947,N_13576,N_13287);
xnor U14948 (N_14948,N_13930,N_13095);
nor U14949 (N_14949,N_13257,N_13710);
nor U14950 (N_14950,N_13906,N_13957);
nand U14951 (N_14951,N_13597,N_13673);
xnor U14952 (N_14952,N_13111,N_13665);
xnor U14953 (N_14953,N_13534,N_13633);
nor U14954 (N_14954,N_13944,N_13461);
or U14955 (N_14955,N_13365,N_13486);
xnor U14956 (N_14956,N_13059,N_13804);
and U14957 (N_14957,N_13915,N_13232);
and U14958 (N_14958,N_13245,N_13521);
xnor U14959 (N_14959,N_13965,N_13288);
xnor U14960 (N_14960,N_13361,N_13531);
nor U14961 (N_14961,N_13783,N_13395);
nand U14962 (N_14962,N_13388,N_13441);
nor U14963 (N_14963,N_13061,N_13106);
xnor U14964 (N_14964,N_13212,N_13216);
nor U14965 (N_14965,N_13270,N_13614);
and U14966 (N_14966,N_13294,N_13715);
and U14967 (N_14967,N_13330,N_13981);
xnor U14968 (N_14968,N_13936,N_13952);
and U14969 (N_14969,N_13547,N_13159);
or U14970 (N_14970,N_13910,N_13053);
and U14971 (N_14971,N_13189,N_13747);
and U14972 (N_14972,N_13544,N_13104);
xnor U14973 (N_14973,N_13097,N_13243);
nand U14974 (N_14974,N_13726,N_13531);
nor U14975 (N_14975,N_13944,N_13099);
and U14976 (N_14976,N_13859,N_13880);
and U14977 (N_14977,N_13558,N_13030);
nand U14978 (N_14978,N_13708,N_13657);
and U14979 (N_14979,N_13722,N_13520);
nor U14980 (N_14980,N_13605,N_13894);
xor U14981 (N_14981,N_13332,N_13365);
nor U14982 (N_14982,N_13955,N_13947);
and U14983 (N_14983,N_13858,N_13049);
or U14984 (N_14984,N_13654,N_13694);
nor U14985 (N_14985,N_13164,N_13442);
xor U14986 (N_14986,N_13848,N_13855);
nand U14987 (N_14987,N_13849,N_13564);
nor U14988 (N_14988,N_13189,N_13711);
xor U14989 (N_14989,N_13261,N_13680);
xnor U14990 (N_14990,N_13025,N_13584);
and U14991 (N_14991,N_13271,N_13501);
nor U14992 (N_14992,N_13908,N_13904);
nand U14993 (N_14993,N_13919,N_13774);
nand U14994 (N_14994,N_13625,N_13334);
and U14995 (N_14995,N_13315,N_13310);
and U14996 (N_14996,N_13993,N_13913);
xor U14997 (N_14997,N_13557,N_13523);
nand U14998 (N_14998,N_13960,N_13765);
or U14999 (N_14999,N_13763,N_13981);
and U15000 (N_15000,N_14633,N_14727);
xnor U15001 (N_15001,N_14610,N_14855);
and U15002 (N_15002,N_14442,N_14611);
and U15003 (N_15003,N_14078,N_14620);
xnor U15004 (N_15004,N_14344,N_14183);
nor U15005 (N_15005,N_14098,N_14250);
or U15006 (N_15006,N_14042,N_14103);
or U15007 (N_15007,N_14313,N_14529);
or U15008 (N_15008,N_14389,N_14733);
nand U15009 (N_15009,N_14572,N_14152);
xnor U15010 (N_15010,N_14781,N_14840);
nor U15011 (N_15011,N_14866,N_14374);
xor U15012 (N_15012,N_14211,N_14566);
xnor U15013 (N_15013,N_14940,N_14767);
and U15014 (N_15014,N_14047,N_14385);
nand U15015 (N_15015,N_14519,N_14160);
xnor U15016 (N_15016,N_14808,N_14467);
xor U15017 (N_15017,N_14458,N_14701);
nor U15018 (N_15018,N_14127,N_14999);
nor U15019 (N_15019,N_14897,N_14121);
nor U15020 (N_15020,N_14925,N_14687);
nor U15021 (N_15021,N_14594,N_14192);
xor U15022 (N_15022,N_14386,N_14278);
nand U15023 (N_15023,N_14315,N_14931);
nor U15024 (N_15024,N_14626,N_14492);
xnor U15025 (N_15025,N_14031,N_14876);
nor U15026 (N_15026,N_14268,N_14388);
nand U15027 (N_15027,N_14728,N_14437);
xnor U15028 (N_15028,N_14994,N_14692);
or U15029 (N_15029,N_14478,N_14394);
nand U15030 (N_15030,N_14026,N_14327);
nand U15031 (N_15031,N_14011,N_14396);
and U15032 (N_15032,N_14469,N_14254);
or U15033 (N_15033,N_14191,N_14898);
xnor U15034 (N_15034,N_14227,N_14669);
or U15035 (N_15035,N_14190,N_14653);
and U15036 (N_15036,N_14498,N_14907);
or U15037 (N_15037,N_14844,N_14271);
nand U15038 (N_15038,N_14277,N_14102);
and U15039 (N_15039,N_14032,N_14184);
nor U15040 (N_15040,N_14599,N_14223);
or U15041 (N_15041,N_14361,N_14380);
xor U15042 (N_15042,N_14915,N_14238);
xnor U15043 (N_15043,N_14731,N_14048);
nand U15044 (N_15044,N_14601,N_14944);
nand U15045 (N_15045,N_14792,N_14966);
xor U15046 (N_15046,N_14038,N_14283);
or U15047 (N_15047,N_14305,N_14249);
or U15048 (N_15048,N_14001,N_14597);
nand U15049 (N_15049,N_14137,N_14883);
and U15050 (N_15050,N_14723,N_14295);
nand U15051 (N_15051,N_14387,N_14646);
xor U15052 (N_15052,N_14563,N_14892);
nor U15053 (N_15053,N_14658,N_14642);
or U15054 (N_15054,N_14612,N_14555);
and U15055 (N_15055,N_14124,N_14065);
nand U15056 (N_15056,N_14694,N_14319);
or U15057 (N_15057,N_14096,N_14707);
and U15058 (N_15058,N_14012,N_14756);
xor U15059 (N_15059,N_14325,N_14774);
nand U15060 (N_15060,N_14814,N_14422);
nand U15061 (N_15061,N_14076,N_14812);
nand U15062 (N_15062,N_14314,N_14104);
and U15063 (N_15063,N_14435,N_14013);
xor U15064 (N_15064,N_14644,N_14182);
or U15065 (N_15065,N_14963,N_14595);
or U15066 (N_15066,N_14805,N_14430);
nor U15067 (N_15067,N_14588,N_14662);
nand U15068 (N_15068,N_14894,N_14819);
xnor U15069 (N_15069,N_14933,N_14260);
and U15070 (N_15070,N_14000,N_14901);
nor U15071 (N_15071,N_14400,N_14123);
and U15072 (N_15072,N_14280,N_14275);
nor U15073 (N_15073,N_14266,N_14220);
or U15074 (N_15074,N_14230,N_14831);
and U15075 (N_15075,N_14711,N_14861);
nor U15076 (N_15076,N_14348,N_14288);
xnor U15077 (N_15077,N_14432,N_14824);
xnor U15078 (N_15078,N_14689,N_14281);
or U15079 (N_15079,N_14961,N_14217);
nand U15080 (N_15080,N_14444,N_14638);
and U15081 (N_15081,N_14450,N_14110);
or U15082 (N_15082,N_14058,N_14600);
nor U15083 (N_15083,N_14213,N_14801);
or U15084 (N_15084,N_14057,N_14856);
and U15085 (N_15085,N_14815,N_14089);
nand U15086 (N_15086,N_14232,N_14079);
xor U15087 (N_15087,N_14481,N_14429);
or U15088 (N_15088,N_14797,N_14670);
and U15089 (N_15089,N_14234,N_14914);
nor U15090 (N_15090,N_14331,N_14616);
or U15091 (N_15091,N_14393,N_14377);
nor U15092 (N_15092,N_14911,N_14068);
xor U15093 (N_15093,N_14535,N_14991);
nor U15094 (N_15094,N_14782,N_14099);
and U15095 (N_15095,N_14335,N_14912);
and U15096 (N_15096,N_14242,N_14164);
nor U15097 (N_15097,N_14645,N_14857);
and U15098 (N_15098,N_14292,N_14142);
and U15099 (N_15099,N_14251,N_14061);
or U15100 (N_15100,N_14603,N_14128);
and U15101 (N_15101,N_14997,N_14412);
or U15102 (N_15102,N_14904,N_14527);
xor U15103 (N_15103,N_14204,N_14162);
nor U15104 (N_15104,N_14365,N_14029);
nor U15105 (N_15105,N_14246,N_14093);
nor U15106 (N_15106,N_14918,N_14871);
or U15107 (N_15107,N_14346,N_14482);
xor U15108 (N_15108,N_14417,N_14425);
nand U15109 (N_15109,N_14177,N_14917);
nand U15110 (N_15110,N_14008,N_14896);
xnor U15111 (N_15111,N_14686,N_14452);
or U15112 (N_15112,N_14743,N_14524);
or U15113 (N_15113,N_14475,N_14521);
nand U15114 (N_15114,N_14114,N_14285);
nand U15115 (N_15115,N_14221,N_14958);
and U15116 (N_15116,N_14874,N_14431);
xor U15117 (N_15117,N_14328,N_14980);
nor U15118 (N_15118,N_14556,N_14965);
or U15119 (N_15119,N_14153,N_14456);
and U15120 (N_15120,N_14567,N_14820);
and U15121 (N_15121,N_14559,N_14274);
nor U15122 (N_15122,N_14919,N_14439);
nand U15123 (N_15123,N_14582,N_14647);
nand U15124 (N_15124,N_14257,N_14621);
and U15125 (N_15125,N_14130,N_14256);
nand U15126 (N_15126,N_14222,N_14451);
nor U15127 (N_15127,N_14859,N_14712);
nand U15128 (N_15128,N_14290,N_14839);
nor U15129 (N_15129,N_14636,N_14625);
or U15130 (N_15130,N_14462,N_14675);
and U15131 (N_15131,N_14214,N_14705);
and U15132 (N_15132,N_14847,N_14846);
and U15133 (N_15133,N_14643,N_14156);
nor U15134 (N_15134,N_14334,N_14818);
xor U15135 (N_15135,N_14040,N_14542);
xnor U15136 (N_15136,N_14323,N_14485);
nor U15137 (N_15137,N_14690,N_14070);
nor U15138 (N_15138,N_14447,N_14071);
nor U15139 (N_15139,N_14186,N_14009);
xor U15140 (N_15140,N_14592,N_14623);
xor U15141 (N_15141,N_14209,N_14970);
nand U15142 (N_15142,N_14253,N_14024);
nand U15143 (N_15143,N_14373,N_14858);
xor U15144 (N_15144,N_14516,N_14522);
and U15145 (N_15145,N_14660,N_14165);
nor U15146 (N_15146,N_14459,N_14472);
or U15147 (N_15147,N_14320,N_14979);
nor U15148 (N_15148,N_14715,N_14391);
nor U15149 (N_15149,N_14986,N_14004);
nor U15150 (N_15150,N_14838,N_14816);
and U15151 (N_15151,N_14695,N_14877);
nand U15152 (N_15152,N_14585,N_14548);
nand U15153 (N_15153,N_14166,N_14113);
or U15154 (N_15154,N_14730,N_14515);
xor U15155 (N_15155,N_14457,N_14414);
xor U15156 (N_15156,N_14025,N_14353);
nand U15157 (N_15157,N_14552,N_14806);
nor U15158 (N_15158,N_14413,N_14960);
or U15159 (N_15159,N_14484,N_14860);
nor U15160 (N_15160,N_14580,N_14329);
or U15161 (N_15161,N_14893,N_14651);
and U15162 (N_15162,N_14202,N_14746);
and U15163 (N_15163,N_14398,N_14569);
xnor U15164 (N_15164,N_14879,N_14330);
or U15165 (N_15165,N_14590,N_14537);
xnor U15166 (N_15166,N_14419,N_14203);
xor U15167 (N_15167,N_14796,N_14787);
nand U15168 (N_15168,N_14639,N_14115);
nor U15169 (N_15169,N_14433,N_14120);
nand U15170 (N_15170,N_14971,N_14678);
or U15171 (N_15171,N_14117,N_14577);
or U15172 (N_15172,N_14721,N_14265);
xnor U15173 (N_15173,N_14005,N_14108);
xor U15174 (N_15174,N_14229,N_14403);
xor U15175 (N_15175,N_14967,N_14667);
and U15176 (N_15176,N_14423,N_14943);
or U15177 (N_15177,N_14946,N_14528);
or U15178 (N_15178,N_14852,N_14188);
or U15179 (N_15179,N_14648,N_14195);
and U15180 (N_15180,N_14789,N_14404);
and U15181 (N_15181,N_14872,N_14929);
or U15182 (N_15182,N_14509,N_14953);
xor U15183 (N_15183,N_14363,N_14118);
xor U15184 (N_15184,N_14978,N_14228);
and U15185 (N_15185,N_14354,N_14109);
and U15186 (N_15186,N_14685,N_14410);
or U15187 (N_15187,N_14794,N_14030);
nand U15188 (N_15188,N_14084,N_14366);
and U15189 (N_15189,N_14095,N_14225);
or U15190 (N_15190,N_14698,N_14074);
and U15191 (N_15191,N_14749,N_14307);
or U15192 (N_15192,N_14710,N_14501);
xnor U15193 (N_15193,N_14027,N_14573);
and U15194 (N_15194,N_14504,N_14411);
nor U15195 (N_15195,N_14306,N_14825);
and U15196 (N_15196,N_14742,N_14196);
nor U15197 (N_15197,N_14359,N_14656);
nand U15198 (N_15198,N_14575,N_14201);
nand U15199 (N_15199,N_14461,N_14773);
or U15200 (N_15200,N_14218,N_14163);
nand U15201 (N_15201,N_14215,N_14833);
nand U15202 (N_15202,N_14378,N_14021);
xor U15203 (N_15203,N_14640,N_14972);
and U15204 (N_15204,N_14069,N_14783);
nor U15205 (N_15205,N_14887,N_14672);
or U15206 (N_15206,N_14854,N_14652);
or U15207 (N_15207,N_14637,N_14902);
xor U15208 (N_15208,N_14134,N_14959);
xnor U15209 (N_15209,N_14576,N_14405);
xor U15210 (N_15210,N_14176,N_14035);
and U15211 (N_15211,N_14748,N_14937);
nand U15212 (N_15212,N_14468,N_14523);
nor U15213 (N_15213,N_14751,N_14453);
xor U15214 (N_15214,N_14677,N_14718);
nand U15215 (N_15215,N_14141,N_14438);
xor U15216 (N_15216,N_14992,N_14862);
and U15217 (N_15217,N_14136,N_14090);
xnor U15218 (N_15218,N_14039,N_14022);
nor U15219 (N_15219,N_14550,N_14880);
xor U15220 (N_15220,N_14514,N_14878);
or U15221 (N_15221,N_14370,N_14360);
and U15222 (N_15222,N_14362,N_14493);
nand U15223 (N_15223,N_14416,N_14622);
xor U15224 (N_15224,N_14488,N_14807);
and U15225 (N_15225,N_14499,N_14395);
xnor U15226 (N_15226,N_14836,N_14780);
nand U15227 (N_15227,N_14697,N_14664);
nand U15228 (N_15228,N_14544,N_14744);
xnor U15229 (N_15229,N_14083,N_14635);
or U15230 (N_15230,N_14799,N_14784);
and U15231 (N_15231,N_14541,N_14741);
xnor U15232 (N_15232,N_14041,N_14954);
or U15233 (N_15233,N_14684,N_14270);
xnor U15234 (N_15234,N_14064,N_14267);
nand U15235 (N_15235,N_14018,N_14899);
and U15236 (N_15236,N_14464,N_14171);
nor U15237 (N_15237,N_14298,N_14489);
and U15238 (N_15238,N_14154,N_14473);
or U15239 (N_15239,N_14553,N_14116);
and U15240 (N_15240,N_14460,N_14341);
nand U15241 (N_15241,N_14140,N_14198);
nor U15242 (N_15242,N_14668,N_14843);
and U15243 (N_15243,N_14261,N_14988);
and U15244 (N_15244,N_14778,N_14945);
nand U15245 (N_15245,N_14490,N_14886);
and U15246 (N_15246,N_14981,N_14180);
xor U15247 (N_15247,N_14149,N_14036);
xor U15248 (N_15248,N_14200,N_14920);
or U15249 (N_15249,N_14736,N_14755);
nand U15250 (N_15250,N_14659,N_14976);
xnor U15251 (N_15251,N_14532,N_14665);
xor U15252 (N_15252,N_14949,N_14881);
xor U15253 (N_15253,N_14564,N_14562);
or U15254 (N_15254,N_14734,N_14157);
xor U15255 (N_15255,N_14206,N_14427);
or U15256 (N_15256,N_14724,N_14615);
nand U15257 (N_15257,N_14845,N_14345);
and U15258 (N_15258,N_14173,N_14131);
nor U15259 (N_15259,N_14921,N_14798);
and U15260 (N_15260,N_14571,N_14072);
xor U15261 (N_15261,N_14947,N_14052);
xor U15262 (N_15262,N_14511,N_14606);
and U15263 (N_15263,N_14471,N_14974);
nand U15264 (N_15264,N_14530,N_14604);
nand U15265 (N_15265,N_14494,N_14605);
xnor U15266 (N_15266,N_14015,N_14301);
and U15267 (N_15267,N_14702,N_14474);
nor U15268 (N_15268,N_14826,N_14983);
nor U15269 (N_15269,N_14936,N_14044);
or U15270 (N_15270,N_14415,N_14382);
and U15271 (N_15271,N_14324,N_14602);
nand U15272 (N_15272,N_14147,N_14252);
or U15273 (N_15273,N_14312,N_14409);
nand U15274 (N_15274,N_14863,N_14465);
nand U15275 (N_15275,N_14884,N_14517);
nor U15276 (N_15276,N_14477,N_14709);
nand U15277 (N_15277,N_14169,N_14739);
or U15278 (N_15278,N_14758,N_14407);
xor U15279 (N_15279,N_14151,N_14769);
xnor U15280 (N_15280,N_14060,N_14406);
nor U15281 (N_15281,N_14053,N_14627);
and U15282 (N_15282,N_14584,N_14062);
nand U15283 (N_15283,N_14682,N_14436);
xor U15284 (N_15284,N_14139,N_14063);
nand U15285 (N_15285,N_14939,N_14168);
nor U15286 (N_15286,N_14033,N_14159);
or U15287 (N_15287,N_14932,N_14003);
and U15288 (N_15288,N_14598,N_14355);
or U15289 (N_15289,N_14289,N_14297);
xor U15290 (N_15290,N_14938,N_14143);
nor U15291 (N_15291,N_14086,N_14888);
xor U15292 (N_15292,N_14207,N_14367);
nor U15293 (N_15293,N_14683,N_14119);
and U15294 (N_15294,N_14513,N_14955);
and U15295 (N_15295,N_14837,N_14813);
xor U15296 (N_15296,N_14657,N_14082);
nor U15297 (N_15297,N_14596,N_14512);
xor U15298 (N_15298,N_14122,N_14302);
nand U15299 (N_15299,N_14236,N_14608);
and U15300 (N_15300,N_14628,N_14969);
and U15301 (N_15301,N_14757,N_14817);
nand U15302 (N_15302,N_14158,N_14379);
nand U15303 (N_15303,N_14941,N_14303);
xnor U15304 (N_15304,N_14273,N_14194);
nor U15305 (N_15305,N_14985,N_14922);
xnor U15306 (N_15306,N_14421,N_14631);
nand U15307 (N_15307,N_14101,N_14020);
nor U15308 (N_15308,N_14371,N_14219);
nor U15309 (N_15309,N_14614,N_14752);
nand U15310 (N_15310,N_14506,N_14002);
nand U15311 (N_15311,N_14593,N_14226);
xor U15312 (N_15312,N_14491,N_14750);
nand U15313 (N_15313,N_14729,N_14558);
or U15314 (N_15314,N_14014,N_14336);
xor U15315 (N_15315,N_14241,N_14446);
nor U15316 (N_15316,N_14508,N_14247);
nor U15317 (N_15317,N_14497,N_14231);
or U15318 (N_15318,N_14834,N_14017);
and U15319 (N_15319,N_14426,N_14714);
and U15320 (N_15320,N_14067,N_14924);
or U15321 (N_15321,N_14531,N_14720);
or U15322 (N_15322,N_14129,N_14822);
nor U15323 (N_15323,N_14870,N_14263);
or U15324 (N_15324,N_14187,N_14835);
xor U15325 (N_15325,N_14455,N_14364);
xnor U15326 (N_15326,N_14007,N_14760);
and U15327 (N_15327,N_14913,N_14989);
and U15328 (N_15328,N_14868,N_14765);
nand U15329 (N_15329,N_14926,N_14332);
xnor U15330 (N_15330,N_14565,N_14586);
and U15331 (N_15331,N_14258,N_14560);
xor U15332 (N_15332,N_14486,N_14487);
or U15333 (N_15333,N_14545,N_14111);
xnor U15334 (N_15334,N_14466,N_14347);
xor U15335 (N_15335,N_14869,N_14356);
and U15336 (N_15336,N_14617,N_14269);
nor U15337 (N_15337,N_14144,N_14753);
or U15338 (N_15338,N_14952,N_14264);
nor U15339 (N_15339,N_14525,N_14185);
nand U15340 (N_15340,N_14105,N_14629);
nand U15341 (N_15341,N_14443,N_14681);
and U15342 (N_15342,N_14763,N_14287);
xor U15343 (N_15343,N_14085,N_14713);
nand U15344 (N_15344,N_14338,N_14693);
nand U15345 (N_15345,N_14761,N_14050);
nor U15346 (N_15346,N_14540,N_14240);
nor U15347 (N_15347,N_14823,N_14181);
nor U15348 (N_15348,N_14827,N_14316);
or U15349 (N_15349,N_14674,N_14996);
nand U15350 (N_15350,N_14726,N_14066);
nor U15351 (N_15351,N_14351,N_14088);
nand U15352 (N_15352,N_14759,N_14568);
and U15353 (N_15353,N_14865,N_14679);
nand U15354 (N_15354,N_14770,N_14853);
nor U15355 (N_15355,N_14340,N_14526);
nand U15356 (N_15356,N_14279,N_14830);
and U15357 (N_15357,N_14654,N_14766);
and U15358 (N_15358,N_14737,N_14293);
or U15359 (N_15359,N_14700,N_14538);
nand U15360 (N_15360,N_14133,N_14777);
and U15361 (N_15361,N_14906,N_14779);
and U15362 (N_15362,N_14311,N_14276);
or U15363 (N_15363,N_14634,N_14549);
nor U15364 (N_15364,N_14383,N_14851);
and U15365 (N_15365,N_14245,N_14543);
nor U15366 (N_15366,N_14381,N_14581);
nor U15367 (N_15367,N_14178,N_14080);
or U15368 (N_15368,N_14375,N_14463);
xor U15369 (N_15369,N_14091,N_14804);
xnor U15370 (N_15370,N_14957,N_14318);
and U15371 (N_15371,N_14304,N_14950);
xnor U15372 (N_15372,N_14449,N_14891);
xnor U15373 (N_15373,N_14776,N_14772);
nand U15374 (N_15374,N_14775,N_14500);
nor U15375 (N_15375,N_14977,N_14930);
and U15376 (N_15376,N_14696,N_14503);
and U15377 (N_15377,N_14092,N_14810);
nand U15378 (N_15378,N_14732,N_14272);
and U15379 (N_15379,N_14350,N_14326);
xnor U15380 (N_15380,N_14189,N_14045);
nand U15381 (N_15381,N_14155,N_14179);
and U15382 (N_15382,N_14800,N_14125);
or U15383 (N_15383,N_14424,N_14591);
or U15384 (N_15384,N_14975,N_14867);
nor U15385 (N_15385,N_14802,N_14754);
or U15386 (N_15386,N_14583,N_14745);
and U15387 (N_15387,N_14821,N_14942);
xnor U15388 (N_15388,N_14402,N_14905);
and U15389 (N_15389,N_14300,N_14903);
or U15390 (N_15390,N_14212,N_14510);
nand U15391 (N_15391,N_14671,N_14357);
xnor U15392 (N_15392,N_14547,N_14408);
xnor U15393 (N_15393,N_14909,N_14587);
nor U15394 (N_15394,N_14536,N_14418);
nand U15395 (N_15395,N_14081,N_14243);
and U15396 (N_15396,N_14112,N_14010);
nand U15397 (N_15397,N_14619,N_14502);
and U15398 (N_15398,N_14055,N_14372);
nor U15399 (N_15399,N_14900,N_14019);
or U15400 (N_15400,N_14771,N_14339);
and U15401 (N_15401,N_14376,N_14661);
xnor U15402 (N_15402,N_14135,N_14795);
nand U15403 (N_15403,N_14401,N_14023);
and U15404 (N_15404,N_14570,N_14688);
or U15405 (N_15405,N_14193,N_14308);
and U15406 (N_15406,N_14358,N_14719);
or U15407 (N_15407,N_14259,N_14850);
xor U15408 (N_15408,N_14928,N_14885);
xnor U15409 (N_15409,N_14262,N_14392);
and U15410 (N_15410,N_14397,N_14927);
nor U15411 (N_15411,N_14454,N_14641);
nor U15412 (N_15412,N_14244,N_14968);
nand U15413 (N_15413,N_14995,N_14016);
nand U15414 (N_15414,N_14740,N_14294);
or U15415 (N_15415,N_14321,N_14786);
nor U15416 (N_15416,N_14964,N_14650);
and U15417 (N_15417,N_14768,N_14889);
nor U15418 (N_15418,N_14046,N_14107);
nand U15419 (N_15419,N_14704,N_14717);
xor U15420 (N_15420,N_14809,N_14145);
nor U15421 (N_15421,N_14337,N_14059);
and U15422 (N_15422,N_14174,N_14811);
nand U15423 (N_15423,N_14873,N_14910);
or U15424 (N_15424,N_14791,N_14284);
xnor U15425 (N_15425,N_14051,N_14399);
xor U15426 (N_15426,N_14496,N_14895);
and U15427 (N_15427,N_14935,N_14097);
nand U15428 (N_15428,N_14148,N_14578);
xor U15429 (N_15429,N_14998,N_14237);
and U15430 (N_15430,N_14589,N_14546);
nand U15431 (N_15431,N_14150,N_14309);
nand U15432 (N_15432,N_14073,N_14982);
nand U15433 (N_15433,N_14205,N_14882);
or U15434 (N_15434,N_14934,N_14673);
and U15435 (N_15435,N_14613,N_14434);
xnor U15436 (N_15436,N_14908,N_14483);
nor U15437 (N_15437,N_14956,N_14352);
and U15438 (N_15438,N_14923,N_14170);
nand U15439 (N_15439,N_14832,N_14445);
xnor U15440 (N_15440,N_14077,N_14703);
xnor U15441 (N_15441,N_14428,N_14716);
nand U15442 (N_15442,N_14987,N_14507);
xor U15443 (N_15443,N_14708,N_14842);
nand U15444 (N_15444,N_14172,N_14663);
or U15445 (N_15445,N_14138,N_14006);
and U15446 (N_15446,N_14049,N_14666);
nand U15447 (N_15447,N_14448,N_14216);
xor U15448 (N_15448,N_14793,N_14233);
nand U15449 (N_15449,N_14785,N_14722);
or U15450 (N_15450,N_14551,N_14890);
or U15451 (N_15451,N_14094,N_14291);
or U15452 (N_15452,N_14951,N_14607);
nor U15453 (N_15453,N_14557,N_14480);
nor U15454 (N_15454,N_14175,N_14476);
nor U15455 (N_15455,N_14132,N_14075);
nand U15456 (N_15456,N_14609,N_14829);
nand U15457 (N_15457,N_14146,N_14699);
nor U15458 (N_15458,N_14199,N_14649);
xnor U15459 (N_15459,N_14803,N_14579);
nor U15460 (N_15460,N_14235,N_14790);
or U15461 (N_15461,N_14864,N_14479);
xnor U15462 (N_15462,N_14747,N_14632);
nand U15463 (N_15463,N_14440,N_14948);
or U15464 (N_15464,N_14343,N_14691);
nor U15465 (N_15465,N_14197,N_14384);
nor U15466 (N_15466,N_14764,N_14962);
or U15467 (N_15467,N_14762,N_14210);
xor U15468 (N_15468,N_14849,N_14239);
and U15469 (N_15469,N_14990,N_14706);
and U15470 (N_15470,N_14848,N_14618);
or U15471 (N_15471,N_14333,N_14034);
and U15472 (N_15472,N_14322,N_14161);
or U15473 (N_15473,N_14630,N_14561);
xnor U15474 (N_15474,N_14282,N_14973);
xor U15475 (N_15475,N_14828,N_14495);
nand U15476 (N_15476,N_14680,N_14299);
nor U15477 (N_15477,N_14054,N_14310);
nand U15478 (N_15478,N_14574,N_14100);
nor U15479 (N_15479,N_14368,N_14296);
nor U15480 (N_15480,N_14106,N_14655);
and U15481 (N_15481,N_14248,N_14520);
nand U15482 (N_15482,N_14916,N_14534);
nand U15483 (N_15483,N_14028,N_14554);
xor U15484 (N_15484,N_14369,N_14841);
nor U15485 (N_15485,N_14788,N_14993);
nand U15486 (N_15486,N_14420,N_14208);
xor U15487 (N_15487,N_14349,N_14738);
nor U15488 (N_15488,N_14875,N_14505);
xor U15489 (N_15489,N_14725,N_14286);
or U15490 (N_15490,N_14441,N_14056);
nor U15491 (N_15491,N_14087,N_14255);
xnor U15492 (N_15492,N_14043,N_14224);
and U15493 (N_15493,N_14317,N_14518);
xnor U15494 (N_15494,N_14676,N_14984);
xor U15495 (N_15495,N_14390,N_14167);
and U15496 (N_15496,N_14533,N_14735);
and U15497 (N_15497,N_14126,N_14624);
nand U15498 (N_15498,N_14470,N_14539);
or U15499 (N_15499,N_14037,N_14342);
and U15500 (N_15500,N_14994,N_14063);
or U15501 (N_15501,N_14472,N_14806);
and U15502 (N_15502,N_14628,N_14104);
xor U15503 (N_15503,N_14469,N_14707);
xor U15504 (N_15504,N_14113,N_14106);
nor U15505 (N_15505,N_14816,N_14377);
nand U15506 (N_15506,N_14099,N_14820);
nor U15507 (N_15507,N_14031,N_14783);
nor U15508 (N_15508,N_14428,N_14326);
nand U15509 (N_15509,N_14548,N_14846);
and U15510 (N_15510,N_14872,N_14185);
nor U15511 (N_15511,N_14316,N_14442);
nand U15512 (N_15512,N_14027,N_14575);
nor U15513 (N_15513,N_14665,N_14016);
nand U15514 (N_15514,N_14034,N_14723);
xnor U15515 (N_15515,N_14410,N_14821);
nand U15516 (N_15516,N_14333,N_14513);
and U15517 (N_15517,N_14909,N_14601);
nor U15518 (N_15518,N_14738,N_14739);
nor U15519 (N_15519,N_14306,N_14424);
and U15520 (N_15520,N_14469,N_14743);
and U15521 (N_15521,N_14559,N_14811);
nor U15522 (N_15522,N_14550,N_14213);
xor U15523 (N_15523,N_14726,N_14985);
nor U15524 (N_15524,N_14873,N_14699);
or U15525 (N_15525,N_14326,N_14123);
nand U15526 (N_15526,N_14749,N_14588);
and U15527 (N_15527,N_14429,N_14012);
nand U15528 (N_15528,N_14238,N_14465);
xnor U15529 (N_15529,N_14899,N_14561);
nor U15530 (N_15530,N_14748,N_14691);
xor U15531 (N_15531,N_14203,N_14611);
or U15532 (N_15532,N_14171,N_14169);
xor U15533 (N_15533,N_14986,N_14977);
nand U15534 (N_15534,N_14305,N_14399);
and U15535 (N_15535,N_14680,N_14619);
or U15536 (N_15536,N_14194,N_14855);
xor U15537 (N_15537,N_14976,N_14564);
and U15538 (N_15538,N_14309,N_14560);
nor U15539 (N_15539,N_14027,N_14140);
xor U15540 (N_15540,N_14208,N_14083);
or U15541 (N_15541,N_14115,N_14476);
nor U15542 (N_15542,N_14456,N_14109);
or U15543 (N_15543,N_14434,N_14853);
xnor U15544 (N_15544,N_14363,N_14197);
or U15545 (N_15545,N_14435,N_14174);
or U15546 (N_15546,N_14367,N_14575);
or U15547 (N_15547,N_14593,N_14885);
nor U15548 (N_15548,N_14165,N_14391);
or U15549 (N_15549,N_14333,N_14471);
nor U15550 (N_15550,N_14155,N_14366);
nor U15551 (N_15551,N_14131,N_14548);
nand U15552 (N_15552,N_14271,N_14000);
xor U15553 (N_15553,N_14171,N_14001);
xnor U15554 (N_15554,N_14407,N_14657);
or U15555 (N_15555,N_14928,N_14445);
nor U15556 (N_15556,N_14386,N_14586);
or U15557 (N_15557,N_14037,N_14528);
nand U15558 (N_15558,N_14353,N_14774);
nand U15559 (N_15559,N_14530,N_14111);
nor U15560 (N_15560,N_14854,N_14848);
and U15561 (N_15561,N_14050,N_14195);
and U15562 (N_15562,N_14731,N_14091);
nand U15563 (N_15563,N_14168,N_14700);
or U15564 (N_15564,N_14399,N_14796);
and U15565 (N_15565,N_14408,N_14180);
xor U15566 (N_15566,N_14631,N_14881);
and U15567 (N_15567,N_14641,N_14285);
xor U15568 (N_15568,N_14405,N_14090);
xnor U15569 (N_15569,N_14111,N_14488);
xnor U15570 (N_15570,N_14467,N_14549);
xor U15571 (N_15571,N_14885,N_14874);
or U15572 (N_15572,N_14709,N_14190);
xnor U15573 (N_15573,N_14081,N_14750);
nand U15574 (N_15574,N_14593,N_14635);
nor U15575 (N_15575,N_14029,N_14209);
and U15576 (N_15576,N_14426,N_14677);
xnor U15577 (N_15577,N_14863,N_14284);
or U15578 (N_15578,N_14007,N_14364);
xor U15579 (N_15579,N_14862,N_14749);
nor U15580 (N_15580,N_14081,N_14148);
nand U15581 (N_15581,N_14682,N_14024);
nand U15582 (N_15582,N_14808,N_14425);
xor U15583 (N_15583,N_14436,N_14700);
nand U15584 (N_15584,N_14811,N_14760);
or U15585 (N_15585,N_14723,N_14445);
and U15586 (N_15586,N_14208,N_14419);
nand U15587 (N_15587,N_14255,N_14723);
nand U15588 (N_15588,N_14172,N_14447);
xor U15589 (N_15589,N_14404,N_14811);
xnor U15590 (N_15590,N_14116,N_14697);
xor U15591 (N_15591,N_14883,N_14810);
nor U15592 (N_15592,N_14648,N_14975);
or U15593 (N_15593,N_14062,N_14310);
xnor U15594 (N_15594,N_14936,N_14481);
nor U15595 (N_15595,N_14758,N_14330);
xnor U15596 (N_15596,N_14280,N_14692);
nand U15597 (N_15597,N_14847,N_14388);
or U15598 (N_15598,N_14431,N_14087);
nand U15599 (N_15599,N_14869,N_14785);
or U15600 (N_15600,N_14418,N_14577);
and U15601 (N_15601,N_14200,N_14340);
nor U15602 (N_15602,N_14845,N_14028);
nand U15603 (N_15603,N_14625,N_14518);
nor U15604 (N_15604,N_14463,N_14187);
xor U15605 (N_15605,N_14700,N_14549);
nor U15606 (N_15606,N_14005,N_14794);
nand U15607 (N_15607,N_14540,N_14083);
nor U15608 (N_15608,N_14015,N_14283);
xor U15609 (N_15609,N_14980,N_14368);
and U15610 (N_15610,N_14403,N_14625);
or U15611 (N_15611,N_14443,N_14125);
and U15612 (N_15612,N_14137,N_14838);
and U15613 (N_15613,N_14228,N_14332);
nand U15614 (N_15614,N_14453,N_14345);
xnor U15615 (N_15615,N_14012,N_14109);
nand U15616 (N_15616,N_14429,N_14274);
nor U15617 (N_15617,N_14941,N_14085);
or U15618 (N_15618,N_14501,N_14159);
nor U15619 (N_15619,N_14535,N_14016);
and U15620 (N_15620,N_14277,N_14238);
nor U15621 (N_15621,N_14471,N_14343);
nand U15622 (N_15622,N_14116,N_14467);
xor U15623 (N_15623,N_14521,N_14350);
nor U15624 (N_15624,N_14202,N_14799);
xor U15625 (N_15625,N_14059,N_14759);
or U15626 (N_15626,N_14367,N_14415);
and U15627 (N_15627,N_14866,N_14442);
or U15628 (N_15628,N_14713,N_14381);
nand U15629 (N_15629,N_14818,N_14930);
or U15630 (N_15630,N_14756,N_14278);
and U15631 (N_15631,N_14961,N_14502);
and U15632 (N_15632,N_14591,N_14058);
or U15633 (N_15633,N_14954,N_14637);
xor U15634 (N_15634,N_14764,N_14287);
nand U15635 (N_15635,N_14467,N_14928);
or U15636 (N_15636,N_14360,N_14078);
nand U15637 (N_15637,N_14164,N_14927);
nor U15638 (N_15638,N_14071,N_14366);
xnor U15639 (N_15639,N_14494,N_14076);
or U15640 (N_15640,N_14714,N_14217);
nor U15641 (N_15641,N_14748,N_14012);
nor U15642 (N_15642,N_14894,N_14839);
nand U15643 (N_15643,N_14539,N_14441);
nor U15644 (N_15644,N_14490,N_14342);
or U15645 (N_15645,N_14885,N_14526);
and U15646 (N_15646,N_14956,N_14678);
or U15647 (N_15647,N_14533,N_14236);
nor U15648 (N_15648,N_14295,N_14573);
nand U15649 (N_15649,N_14433,N_14361);
xor U15650 (N_15650,N_14690,N_14726);
and U15651 (N_15651,N_14562,N_14274);
and U15652 (N_15652,N_14089,N_14603);
and U15653 (N_15653,N_14551,N_14405);
nor U15654 (N_15654,N_14030,N_14928);
or U15655 (N_15655,N_14968,N_14020);
and U15656 (N_15656,N_14278,N_14822);
and U15657 (N_15657,N_14691,N_14517);
and U15658 (N_15658,N_14374,N_14412);
or U15659 (N_15659,N_14748,N_14622);
or U15660 (N_15660,N_14715,N_14614);
and U15661 (N_15661,N_14698,N_14614);
xor U15662 (N_15662,N_14132,N_14276);
xnor U15663 (N_15663,N_14866,N_14249);
xor U15664 (N_15664,N_14491,N_14023);
xor U15665 (N_15665,N_14586,N_14681);
or U15666 (N_15666,N_14190,N_14275);
nor U15667 (N_15667,N_14155,N_14298);
and U15668 (N_15668,N_14549,N_14715);
nand U15669 (N_15669,N_14402,N_14355);
and U15670 (N_15670,N_14607,N_14134);
or U15671 (N_15671,N_14799,N_14300);
nand U15672 (N_15672,N_14042,N_14196);
xor U15673 (N_15673,N_14021,N_14123);
and U15674 (N_15674,N_14660,N_14694);
and U15675 (N_15675,N_14801,N_14853);
nand U15676 (N_15676,N_14446,N_14047);
and U15677 (N_15677,N_14911,N_14710);
nor U15678 (N_15678,N_14682,N_14737);
nand U15679 (N_15679,N_14376,N_14105);
nand U15680 (N_15680,N_14380,N_14370);
nand U15681 (N_15681,N_14162,N_14879);
nor U15682 (N_15682,N_14325,N_14139);
nand U15683 (N_15683,N_14127,N_14500);
and U15684 (N_15684,N_14734,N_14488);
or U15685 (N_15685,N_14902,N_14700);
nor U15686 (N_15686,N_14310,N_14504);
nor U15687 (N_15687,N_14015,N_14629);
nand U15688 (N_15688,N_14285,N_14394);
and U15689 (N_15689,N_14774,N_14226);
nand U15690 (N_15690,N_14452,N_14966);
nor U15691 (N_15691,N_14678,N_14510);
or U15692 (N_15692,N_14284,N_14015);
nor U15693 (N_15693,N_14955,N_14808);
nand U15694 (N_15694,N_14582,N_14999);
nand U15695 (N_15695,N_14912,N_14776);
and U15696 (N_15696,N_14244,N_14236);
xnor U15697 (N_15697,N_14006,N_14709);
nor U15698 (N_15698,N_14232,N_14991);
nand U15699 (N_15699,N_14776,N_14165);
or U15700 (N_15700,N_14575,N_14769);
nand U15701 (N_15701,N_14341,N_14303);
nand U15702 (N_15702,N_14107,N_14238);
and U15703 (N_15703,N_14494,N_14735);
and U15704 (N_15704,N_14638,N_14577);
and U15705 (N_15705,N_14128,N_14450);
or U15706 (N_15706,N_14466,N_14565);
and U15707 (N_15707,N_14717,N_14207);
and U15708 (N_15708,N_14638,N_14779);
xnor U15709 (N_15709,N_14514,N_14182);
or U15710 (N_15710,N_14200,N_14348);
and U15711 (N_15711,N_14457,N_14906);
or U15712 (N_15712,N_14488,N_14633);
or U15713 (N_15713,N_14759,N_14966);
or U15714 (N_15714,N_14727,N_14907);
nand U15715 (N_15715,N_14332,N_14532);
or U15716 (N_15716,N_14398,N_14816);
and U15717 (N_15717,N_14222,N_14025);
nor U15718 (N_15718,N_14196,N_14300);
or U15719 (N_15719,N_14863,N_14555);
xor U15720 (N_15720,N_14303,N_14058);
nand U15721 (N_15721,N_14348,N_14469);
and U15722 (N_15722,N_14623,N_14274);
or U15723 (N_15723,N_14552,N_14051);
nor U15724 (N_15724,N_14275,N_14979);
and U15725 (N_15725,N_14019,N_14113);
nor U15726 (N_15726,N_14336,N_14708);
nand U15727 (N_15727,N_14823,N_14168);
nand U15728 (N_15728,N_14385,N_14489);
nor U15729 (N_15729,N_14182,N_14165);
nor U15730 (N_15730,N_14444,N_14801);
or U15731 (N_15731,N_14234,N_14607);
or U15732 (N_15732,N_14988,N_14564);
and U15733 (N_15733,N_14118,N_14819);
xnor U15734 (N_15734,N_14243,N_14770);
and U15735 (N_15735,N_14410,N_14048);
xnor U15736 (N_15736,N_14429,N_14103);
nor U15737 (N_15737,N_14621,N_14473);
nand U15738 (N_15738,N_14678,N_14490);
or U15739 (N_15739,N_14802,N_14706);
nand U15740 (N_15740,N_14627,N_14389);
xor U15741 (N_15741,N_14210,N_14302);
or U15742 (N_15742,N_14758,N_14792);
or U15743 (N_15743,N_14264,N_14622);
or U15744 (N_15744,N_14507,N_14342);
and U15745 (N_15745,N_14776,N_14004);
nor U15746 (N_15746,N_14699,N_14461);
and U15747 (N_15747,N_14906,N_14999);
xor U15748 (N_15748,N_14037,N_14899);
xor U15749 (N_15749,N_14157,N_14115);
nand U15750 (N_15750,N_14814,N_14369);
or U15751 (N_15751,N_14846,N_14608);
and U15752 (N_15752,N_14165,N_14256);
nor U15753 (N_15753,N_14469,N_14443);
and U15754 (N_15754,N_14502,N_14988);
and U15755 (N_15755,N_14962,N_14088);
nor U15756 (N_15756,N_14609,N_14495);
xnor U15757 (N_15757,N_14437,N_14848);
nor U15758 (N_15758,N_14729,N_14324);
nor U15759 (N_15759,N_14920,N_14159);
nand U15760 (N_15760,N_14183,N_14105);
nor U15761 (N_15761,N_14812,N_14208);
nor U15762 (N_15762,N_14916,N_14764);
nor U15763 (N_15763,N_14675,N_14069);
or U15764 (N_15764,N_14478,N_14821);
nand U15765 (N_15765,N_14600,N_14224);
nor U15766 (N_15766,N_14829,N_14886);
and U15767 (N_15767,N_14587,N_14546);
nor U15768 (N_15768,N_14037,N_14373);
nand U15769 (N_15769,N_14452,N_14041);
xor U15770 (N_15770,N_14831,N_14300);
and U15771 (N_15771,N_14039,N_14721);
nand U15772 (N_15772,N_14386,N_14338);
or U15773 (N_15773,N_14794,N_14928);
nor U15774 (N_15774,N_14194,N_14264);
or U15775 (N_15775,N_14328,N_14782);
nand U15776 (N_15776,N_14878,N_14677);
and U15777 (N_15777,N_14803,N_14485);
xor U15778 (N_15778,N_14007,N_14051);
nor U15779 (N_15779,N_14983,N_14665);
nor U15780 (N_15780,N_14044,N_14410);
and U15781 (N_15781,N_14765,N_14364);
nand U15782 (N_15782,N_14586,N_14106);
and U15783 (N_15783,N_14379,N_14466);
xnor U15784 (N_15784,N_14146,N_14258);
and U15785 (N_15785,N_14146,N_14627);
or U15786 (N_15786,N_14095,N_14836);
or U15787 (N_15787,N_14424,N_14696);
nand U15788 (N_15788,N_14928,N_14135);
xnor U15789 (N_15789,N_14360,N_14826);
nor U15790 (N_15790,N_14997,N_14314);
xnor U15791 (N_15791,N_14118,N_14700);
nand U15792 (N_15792,N_14786,N_14357);
nor U15793 (N_15793,N_14465,N_14933);
or U15794 (N_15794,N_14676,N_14040);
nor U15795 (N_15795,N_14160,N_14027);
or U15796 (N_15796,N_14858,N_14512);
nor U15797 (N_15797,N_14622,N_14380);
nand U15798 (N_15798,N_14977,N_14837);
xnor U15799 (N_15799,N_14744,N_14806);
or U15800 (N_15800,N_14775,N_14298);
nor U15801 (N_15801,N_14244,N_14436);
nand U15802 (N_15802,N_14862,N_14670);
nor U15803 (N_15803,N_14750,N_14043);
and U15804 (N_15804,N_14397,N_14755);
and U15805 (N_15805,N_14147,N_14205);
and U15806 (N_15806,N_14597,N_14518);
nand U15807 (N_15807,N_14176,N_14399);
or U15808 (N_15808,N_14532,N_14231);
xnor U15809 (N_15809,N_14043,N_14946);
nand U15810 (N_15810,N_14808,N_14335);
and U15811 (N_15811,N_14014,N_14234);
xor U15812 (N_15812,N_14838,N_14023);
or U15813 (N_15813,N_14460,N_14838);
and U15814 (N_15814,N_14588,N_14932);
nor U15815 (N_15815,N_14551,N_14646);
and U15816 (N_15816,N_14925,N_14701);
nand U15817 (N_15817,N_14157,N_14204);
nor U15818 (N_15818,N_14661,N_14776);
or U15819 (N_15819,N_14132,N_14571);
nand U15820 (N_15820,N_14686,N_14551);
and U15821 (N_15821,N_14788,N_14078);
nor U15822 (N_15822,N_14525,N_14537);
and U15823 (N_15823,N_14518,N_14404);
nor U15824 (N_15824,N_14513,N_14769);
or U15825 (N_15825,N_14639,N_14371);
and U15826 (N_15826,N_14294,N_14819);
nand U15827 (N_15827,N_14022,N_14583);
and U15828 (N_15828,N_14386,N_14100);
and U15829 (N_15829,N_14457,N_14898);
xor U15830 (N_15830,N_14152,N_14049);
nand U15831 (N_15831,N_14542,N_14650);
xor U15832 (N_15832,N_14010,N_14630);
nor U15833 (N_15833,N_14335,N_14236);
xor U15834 (N_15834,N_14332,N_14741);
and U15835 (N_15835,N_14085,N_14154);
and U15836 (N_15836,N_14526,N_14640);
nor U15837 (N_15837,N_14814,N_14681);
nand U15838 (N_15838,N_14295,N_14398);
xnor U15839 (N_15839,N_14747,N_14892);
or U15840 (N_15840,N_14594,N_14476);
and U15841 (N_15841,N_14197,N_14927);
nand U15842 (N_15842,N_14819,N_14845);
xor U15843 (N_15843,N_14055,N_14405);
and U15844 (N_15844,N_14598,N_14208);
xor U15845 (N_15845,N_14676,N_14214);
or U15846 (N_15846,N_14679,N_14010);
nor U15847 (N_15847,N_14150,N_14192);
nor U15848 (N_15848,N_14466,N_14723);
nor U15849 (N_15849,N_14776,N_14869);
nand U15850 (N_15850,N_14222,N_14715);
xor U15851 (N_15851,N_14163,N_14395);
and U15852 (N_15852,N_14207,N_14235);
xor U15853 (N_15853,N_14562,N_14829);
or U15854 (N_15854,N_14605,N_14488);
or U15855 (N_15855,N_14847,N_14479);
xor U15856 (N_15856,N_14244,N_14945);
nor U15857 (N_15857,N_14151,N_14955);
nand U15858 (N_15858,N_14376,N_14536);
nor U15859 (N_15859,N_14290,N_14585);
and U15860 (N_15860,N_14104,N_14867);
xor U15861 (N_15861,N_14052,N_14530);
xnor U15862 (N_15862,N_14316,N_14462);
nand U15863 (N_15863,N_14190,N_14409);
nor U15864 (N_15864,N_14844,N_14865);
or U15865 (N_15865,N_14188,N_14088);
and U15866 (N_15866,N_14531,N_14450);
xnor U15867 (N_15867,N_14643,N_14565);
or U15868 (N_15868,N_14368,N_14349);
and U15869 (N_15869,N_14587,N_14916);
and U15870 (N_15870,N_14463,N_14689);
xor U15871 (N_15871,N_14413,N_14795);
nor U15872 (N_15872,N_14271,N_14668);
or U15873 (N_15873,N_14485,N_14480);
xnor U15874 (N_15874,N_14379,N_14478);
or U15875 (N_15875,N_14950,N_14021);
xnor U15876 (N_15876,N_14252,N_14621);
nor U15877 (N_15877,N_14049,N_14195);
or U15878 (N_15878,N_14654,N_14590);
and U15879 (N_15879,N_14491,N_14578);
nor U15880 (N_15880,N_14747,N_14021);
xnor U15881 (N_15881,N_14879,N_14502);
and U15882 (N_15882,N_14020,N_14592);
and U15883 (N_15883,N_14418,N_14744);
nor U15884 (N_15884,N_14889,N_14755);
or U15885 (N_15885,N_14902,N_14557);
and U15886 (N_15886,N_14259,N_14202);
and U15887 (N_15887,N_14007,N_14151);
nand U15888 (N_15888,N_14096,N_14504);
and U15889 (N_15889,N_14582,N_14297);
nand U15890 (N_15890,N_14823,N_14633);
xnor U15891 (N_15891,N_14412,N_14493);
or U15892 (N_15892,N_14431,N_14939);
and U15893 (N_15893,N_14253,N_14747);
and U15894 (N_15894,N_14875,N_14158);
or U15895 (N_15895,N_14496,N_14382);
xor U15896 (N_15896,N_14864,N_14186);
nand U15897 (N_15897,N_14334,N_14432);
nand U15898 (N_15898,N_14918,N_14587);
nand U15899 (N_15899,N_14661,N_14889);
nor U15900 (N_15900,N_14649,N_14865);
xor U15901 (N_15901,N_14143,N_14079);
nor U15902 (N_15902,N_14390,N_14242);
nor U15903 (N_15903,N_14721,N_14187);
nor U15904 (N_15904,N_14323,N_14429);
and U15905 (N_15905,N_14350,N_14600);
and U15906 (N_15906,N_14397,N_14840);
and U15907 (N_15907,N_14283,N_14625);
and U15908 (N_15908,N_14707,N_14357);
and U15909 (N_15909,N_14606,N_14834);
and U15910 (N_15910,N_14874,N_14756);
and U15911 (N_15911,N_14289,N_14078);
or U15912 (N_15912,N_14221,N_14587);
and U15913 (N_15913,N_14383,N_14209);
xor U15914 (N_15914,N_14649,N_14698);
xor U15915 (N_15915,N_14147,N_14095);
and U15916 (N_15916,N_14138,N_14702);
nand U15917 (N_15917,N_14313,N_14271);
xor U15918 (N_15918,N_14603,N_14035);
xor U15919 (N_15919,N_14671,N_14688);
and U15920 (N_15920,N_14255,N_14476);
nand U15921 (N_15921,N_14943,N_14946);
xnor U15922 (N_15922,N_14024,N_14380);
and U15923 (N_15923,N_14250,N_14682);
nand U15924 (N_15924,N_14008,N_14398);
or U15925 (N_15925,N_14451,N_14099);
xnor U15926 (N_15926,N_14994,N_14138);
nor U15927 (N_15927,N_14481,N_14110);
xor U15928 (N_15928,N_14687,N_14918);
nor U15929 (N_15929,N_14811,N_14788);
or U15930 (N_15930,N_14396,N_14500);
xor U15931 (N_15931,N_14086,N_14670);
or U15932 (N_15932,N_14493,N_14785);
nand U15933 (N_15933,N_14554,N_14989);
and U15934 (N_15934,N_14197,N_14815);
nand U15935 (N_15935,N_14355,N_14164);
or U15936 (N_15936,N_14416,N_14533);
and U15937 (N_15937,N_14695,N_14542);
xnor U15938 (N_15938,N_14317,N_14772);
or U15939 (N_15939,N_14820,N_14155);
or U15940 (N_15940,N_14454,N_14449);
nand U15941 (N_15941,N_14675,N_14686);
and U15942 (N_15942,N_14800,N_14888);
or U15943 (N_15943,N_14860,N_14536);
or U15944 (N_15944,N_14937,N_14381);
xnor U15945 (N_15945,N_14764,N_14137);
nor U15946 (N_15946,N_14828,N_14771);
nor U15947 (N_15947,N_14800,N_14733);
or U15948 (N_15948,N_14589,N_14620);
and U15949 (N_15949,N_14854,N_14955);
and U15950 (N_15950,N_14815,N_14253);
and U15951 (N_15951,N_14066,N_14044);
nor U15952 (N_15952,N_14853,N_14842);
or U15953 (N_15953,N_14887,N_14500);
nor U15954 (N_15954,N_14490,N_14298);
nand U15955 (N_15955,N_14641,N_14247);
xor U15956 (N_15956,N_14615,N_14381);
and U15957 (N_15957,N_14521,N_14103);
nor U15958 (N_15958,N_14596,N_14426);
nand U15959 (N_15959,N_14539,N_14835);
nand U15960 (N_15960,N_14045,N_14072);
nand U15961 (N_15961,N_14787,N_14922);
nand U15962 (N_15962,N_14488,N_14147);
nand U15963 (N_15963,N_14837,N_14024);
nor U15964 (N_15964,N_14764,N_14644);
xor U15965 (N_15965,N_14411,N_14185);
nor U15966 (N_15966,N_14747,N_14337);
or U15967 (N_15967,N_14061,N_14156);
or U15968 (N_15968,N_14212,N_14320);
and U15969 (N_15969,N_14117,N_14175);
xor U15970 (N_15970,N_14748,N_14689);
or U15971 (N_15971,N_14080,N_14308);
or U15972 (N_15972,N_14805,N_14978);
and U15973 (N_15973,N_14853,N_14597);
xnor U15974 (N_15974,N_14525,N_14209);
and U15975 (N_15975,N_14381,N_14511);
xor U15976 (N_15976,N_14837,N_14903);
nor U15977 (N_15977,N_14247,N_14466);
nor U15978 (N_15978,N_14182,N_14489);
nand U15979 (N_15979,N_14043,N_14513);
nand U15980 (N_15980,N_14706,N_14700);
xnor U15981 (N_15981,N_14208,N_14382);
nor U15982 (N_15982,N_14234,N_14401);
nor U15983 (N_15983,N_14295,N_14943);
and U15984 (N_15984,N_14530,N_14382);
nand U15985 (N_15985,N_14599,N_14292);
and U15986 (N_15986,N_14820,N_14943);
nand U15987 (N_15987,N_14770,N_14073);
nor U15988 (N_15988,N_14377,N_14846);
xor U15989 (N_15989,N_14238,N_14789);
and U15990 (N_15990,N_14344,N_14458);
xor U15991 (N_15991,N_14657,N_14034);
or U15992 (N_15992,N_14757,N_14823);
nand U15993 (N_15993,N_14430,N_14400);
xor U15994 (N_15994,N_14829,N_14791);
nand U15995 (N_15995,N_14800,N_14722);
xor U15996 (N_15996,N_14837,N_14565);
nand U15997 (N_15997,N_14084,N_14873);
xor U15998 (N_15998,N_14926,N_14532);
and U15999 (N_15999,N_14466,N_14318);
nand U16000 (N_16000,N_15267,N_15798);
or U16001 (N_16001,N_15606,N_15067);
nor U16002 (N_16002,N_15247,N_15892);
nand U16003 (N_16003,N_15757,N_15467);
or U16004 (N_16004,N_15992,N_15410);
nand U16005 (N_16005,N_15667,N_15850);
nor U16006 (N_16006,N_15005,N_15002);
nor U16007 (N_16007,N_15224,N_15732);
or U16008 (N_16008,N_15801,N_15384);
nor U16009 (N_16009,N_15649,N_15511);
nand U16010 (N_16010,N_15958,N_15065);
nor U16011 (N_16011,N_15442,N_15391);
and U16012 (N_16012,N_15050,N_15964);
or U16013 (N_16013,N_15293,N_15236);
nor U16014 (N_16014,N_15994,N_15806);
and U16015 (N_16015,N_15825,N_15284);
xnor U16016 (N_16016,N_15895,N_15403);
or U16017 (N_16017,N_15976,N_15222);
nand U16018 (N_16018,N_15154,N_15575);
xor U16019 (N_16019,N_15011,N_15281);
xnor U16020 (N_16020,N_15858,N_15180);
xnor U16021 (N_16021,N_15231,N_15074);
and U16022 (N_16022,N_15693,N_15387);
or U16023 (N_16023,N_15034,N_15450);
nor U16024 (N_16024,N_15592,N_15555);
xor U16025 (N_16025,N_15347,N_15323);
or U16026 (N_16026,N_15171,N_15163);
or U16027 (N_16027,N_15036,N_15717);
or U16028 (N_16028,N_15635,N_15708);
nor U16029 (N_16029,N_15530,N_15153);
xnor U16030 (N_16030,N_15474,N_15871);
nand U16031 (N_16031,N_15977,N_15091);
nand U16032 (N_16032,N_15255,N_15272);
and U16033 (N_16033,N_15351,N_15501);
nand U16034 (N_16034,N_15857,N_15400);
or U16035 (N_16035,N_15271,N_15630);
and U16036 (N_16036,N_15605,N_15142);
nor U16037 (N_16037,N_15202,N_15237);
and U16038 (N_16038,N_15765,N_15967);
or U16039 (N_16039,N_15041,N_15165);
nand U16040 (N_16040,N_15779,N_15356);
xnor U16041 (N_16041,N_15952,N_15793);
xor U16042 (N_16042,N_15081,N_15105);
and U16043 (N_16043,N_15565,N_15586);
nand U16044 (N_16044,N_15889,N_15077);
nand U16045 (N_16045,N_15042,N_15978);
nand U16046 (N_16046,N_15618,N_15220);
nand U16047 (N_16047,N_15006,N_15126);
nand U16048 (N_16048,N_15320,N_15223);
and U16049 (N_16049,N_15758,N_15552);
xnor U16050 (N_16050,N_15874,N_15327);
and U16051 (N_16051,N_15828,N_15848);
nor U16052 (N_16052,N_15553,N_15397);
or U16053 (N_16053,N_15083,N_15738);
and U16054 (N_16054,N_15197,N_15069);
and U16055 (N_16055,N_15880,N_15244);
xor U16056 (N_16056,N_15401,N_15125);
nand U16057 (N_16057,N_15492,N_15665);
xor U16058 (N_16058,N_15517,N_15597);
xnor U16059 (N_16059,N_15346,N_15359);
xnor U16060 (N_16060,N_15845,N_15715);
nor U16061 (N_16061,N_15633,N_15658);
nor U16062 (N_16062,N_15875,N_15532);
xor U16063 (N_16063,N_15203,N_15997);
and U16064 (N_16064,N_15268,N_15856);
or U16065 (N_16065,N_15364,N_15123);
and U16066 (N_16066,N_15479,N_15712);
or U16067 (N_16067,N_15431,N_15756);
and U16068 (N_16068,N_15319,N_15088);
nor U16069 (N_16069,N_15386,N_15701);
and U16070 (N_16070,N_15527,N_15312);
nor U16071 (N_16071,N_15937,N_15417);
xor U16072 (N_16072,N_15315,N_15440);
and U16073 (N_16073,N_15610,N_15705);
nand U16074 (N_16074,N_15189,N_15514);
and U16075 (N_16075,N_15599,N_15972);
or U16076 (N_16076,N_15071,N_15700);
nor U16077 (N_16077,N_15489,N_15852);
nand U16078 (N_16078,N_15644,N_15383);
nor U16079 (N_16079,N_15415,N_15234);
xor U16080 (N_16080,N_15464,N_15653);
xnor U16081 (N_16081,N_15004,N_15776);
xnor U16082 (N_16082,N_15660,N_15556);
xnor U16083 (N_16083,N_15016,N_15689);
and U16084 (N_16084,N_15944,N_15767);
xnor U16085 (N_16085,N_15411,N_15047);
nand U16086 (N_16086,N_15777,N_15743);
xnor U16087 (N_16087,N_15716,N_15557);
and U16088 (N_16088,N_15815,N_15007);
xnor U16089 (N_16089,N_15001,N_15576);
nand U16090 (N_16090,N_15145,N_15064);
nand U16091 (N_16091,N_15233,N_15009);
xor U16092 (N_16092,N_15646,N_15424);
nor U16093 (N_16093,N_15876,N_15294);
or U16094 (N_16094,N_15860,N_15209);
or U16095 (N_16095,N_15690,N_15340);
xor U16096 (N_16096,N_15306,N_15582);
xnor U16097 (N_16097,N_15604,N_15598);
or U16098 (N_16098,N_15138,N_15326);
nor U16099 (N_16099,N_15353,N_15711);
nand U16100 (N_16100,N_15836,N_15988);
or U16101 (N_16101,N_15245,N_15632);
nor U16102 (N_16102,N_15699,N_15648);
nand U16103 (N_16103,N_15526,N_15607);
xnor U16104 (N_16104,N_15573,N_15012);
and U16105 (N_16105,N_15457,N_15110);
nand U16106 (N_16106,N_15460,N_15300);
nor U16107 (N_16107,N_15161,N_15558);
nand U16108 (N_16108,N_15000,N_15325);
nor U16109 (N_16109,N_15038,N_15210);
nand U16110 (N_16110,N_15430,N_15162);
nand U16111 (N_16111,N_15546,N_15191);
nor U16112 (N_16112,N_15336,N_15570);
xor U16113 (N_16113,N_15185,N_15250);
nand U16114 (N_16114,N_15888,N_15748);
or U16115 (N_16115,N_15261,N_15396);
xnor U16116 (N_16116,N_15486,N_15692);
and U16117 (N_16117,N_15655,N_15572);
nor U16118 (N_16118,N_15878,N_15443);
and U16119 (N_16119,N_15803,N_15735);
or U16120 (N_16120,N_15095,N_15563);
nor U16121 (N_16121,N_15723,N_15919);
or U16122 (N_16122,N_15550,N_15774);
nor U16123 (N_16123,N_15102,N_15039);
nor U16124 (N_16124,N_15451,N_15770);
xnor U16125 (N_16125,N_15307,N_15305);
or U16126 (N_16126,N_15522,N_15761);
and U16127 (N_16127,N_15186,N_15082);
and U16128 (N_16128,N_15904,N_15051);
xnor U16129 (N_16129,N_15158,N_15429);
nand U16130 (N_16130,N_15453,N_15407);
or U16131 (N_16131,N_15024,N_15469);
nand U16132 (N_16132,N_15637,N_15683);
nand U16133 (N_16133,N_15645,N_15498);
nand U16134 (N_16134,N_15448,N_15998);
xnor U16135 (N_16135,N_15399,N_15839);
and U16136 (N_16136,N_15955,N_15003);
nand U16137 (N_16137,N_15216,N_15982);
nand U16138 (N_16138,N_15113,N_15932);
and U16139 (N_16139,N_15219,N_15275);
nand U16140 (N_16140,N_15559,N_15891);
or U16141 (N_16141,N_15434,N_15783);
or U16142 (N_16142,N_15625,N_15017);
nor U16143 (N_16143,N_15437,N_15714);
nand U16144 (N_16144,N_15694,N_15722);
and U16145 (N_16145,N_15930,N_15751);
or U16146 (N_16146,N_15178,N_15493);
nor U16147 (N_16147,N_15593,N_15273);
nand U16148 (N_16148,N_15578,N_15395);
and U16149 (N_16149,N_15833,N_15537);
and U16150 (N_16150,N_15931,N_15378);
nor U16151 (N_16151,N_15811,N_15361);
xnor U16152 (N_16152,N_15840,N_15152);
nor U16153 (N_16153,N_15502,N_15547);
xor U16154 (N_16154,N_15979,N_15179);
or U16155 (N_16155,N_15744,N_15938);
and U16156 (N_16156,N_15989,N_15554);
xnor U16157 (N_16157,N_15863,N_15100);
or U16158 (N_16158,N_15279,N_15936);
and U16159 (N_16159,N_15331,N_15781);
nor U16160 (N_16160,N_15508,N_15452);
nor U16161 (N_16161,N_15942,N_15710);
nand U16162 (N_16162,N_15441,N_15263);
or U16163 (N_16163,N_15476,N_15089);
or U16164 (N_16164,N_15949,N_15205);
nor U16165 (N_16165,N_15029,N_15917);
or U16166 (N_16166,N_15821,N_15943);
nand U16167 (N_16167,N_15373,N_15601);
and U16168 (N_16168,N_15368,N_15729);
nor U16169 (N_16169,N_15674,N_15130);
and U16170 (N_16170,N_15503,N_15996);
nor U16171 (N_16171,N_15897,N_15531);
nand U16172 (N_16172,N_15313,N_15535);
or U16173 (N_16173,N_15355,N_15046);
nand U16174 (N_16174,N_15887,N_15214);
or U16175 (N_16175,N_15536,N_15496);
nand U16176 (N_16176,N_15243,N_15831);
xnor U16177 (N_16177,N_15120,N_15687);
xnor U16178 (N_16178,N_15405,N_15631);
nor U16179 (N_16179,N_15718,N_15843);
xor U16180 (N_16180,N_15264,N_15807);
or U16181 (N_16181,N_15427,N_15829);
and U16182 (N_16182,N_15086,N_15800);
xnor U16183 (N_16183,N_15567,N_15176);
nand U16184 (N_16184,N_15772,N_15249);
and U16185 (N_16185,N_15684,N_15805);
nand U16186 (N_16186,N_15438,N_15144);
nor U16187 (N_16187,N_15851,N_15640);
nor U16188 (N_16188,N_15792,N_15137);
nand U16189 (N_16189,N_15149,N_15902);
nor U16190 (N_16190,N_15623,N_15461);
xnor U16191 (N_16191,N_15406,N_15691);
nand U16192 (N_16192,N_15169,N_15775);
nor U16193 (N_16193,N_15092,N_15339);
and U16194 (N_16194,N_15804,N_15975);
nor U16195 (N_16195,N_15893,N_15168);
or U16196 (N_16196,N_15885,N_15352);
nor U16197 (N_16197,N_15745,N_15468);
nand U16198 (N_16198,N_15033,N_15881);
xor U16199 (N_16199,N_15287,N_15369);
nor U16200 (N_16200,N_15864,N_15256);
xor U16201 (N_16201,N_15797,N_15588);
xor U16202 (N_16202,N_15232,N_15303);
or U16203 (N_16203,N_15311,N_15974);
nand U16204 (N_16204,N_15679,N_15916);
and U16205 (N_16205,N_15362,N_15600);
or U16206 (N_16206,N_15560,N_15622);
xnor U16207 (N_16207,N_15817,N_15132);
nor U16208 (N_16208,N_15960,N_15666);
nand U16209 (N_16209,N_15087,N_15986);
and U16210 (N_16210,N_15076,N_15981);
xor U16211 (N_16211,N_15737,N_15208);
xor U16212 (N_16212,N_15966,N_15616);
xnor U16213 (N_16213,N_15096,N_15070);
and U16214 (N_16214,N_15900,N_15345);
and U16215 (N_16215,N_15215,N_15780);
and U16216 (N_16216,N_15301,N_15118);
or U16217 (N_16217,N_15529,N_15810);
or U16218 (N_16218,N_15238,N_15459);
nand U16219 (N_16219,N_15869,N_15270);
and U16220 (N_16220,N_15923,N_15111);
or U16221 (N_16221,N_15827,N_15151);
nand U16222 (N_16222,N_15366,N_15146);
nand U16223 (N_16223,N_15520,N_15728);
nand U16224 (N_16224,N_15444,N_15289);
nor U16225 (N_16225,N_15905,N_15196);
or U16226 (N_16226,N_15971,N_15439);
xnor U16227 (N_16227,N_15398,N_15544);
xnor U16228 (N_16228,N_15921,N_15926);
xnor U16229 (N_16229,N_15198,N_15954);
or U16230 (N_16230,N_15435,N_15676);
nor U16231 (N_16231,N_15040,N_15870);
nand U16232 (N_16232,N_15354,N_15372);
or U16233 (N_16233,N_15032,N_15020);
or U16234 (N_16234,N_15022,N_15078);
xor U16235 (N_16235,N_15935,N_15436);
xor U16236 (N_16236,N_15659,N_15480);
xnor U16237 (N_16237,N_15119,N_15019);
or U16238 (N_16238,N_15823,N_15910);
nand U16239 (N_16239,N_15611,N_15755);
or U16240 (N_16240,N_15199,N_15494);
xnor U16241 (N_16241,N_15915,N_15172);
and U16242 (N_16242,N_15388,N_15408);
xnor U16243 (N_16243,N_15733,N_15112);
nand U16244 (N_16244,N_15835,N_15968);
or U16245 (N_16245,N_15031,N_15485);
xor U16246 (N_16246,N_15799,N_15357);
nand U16247 (N_16247,N_15995,N_15473);
nor U16248 (N_16248,N_15157,N_15795);
and U16249 (N_16249,N_15656,N_15321);
nor U16250 (N_16250,N_15939,N_15052);
or U16251 (N_16251,N_15059,N_15762);
nand U16252 (N_16252,N_15505,N_15545);
xnor U16253 (N_16253,N_15472,N_15899);
or U16254 (N_16254,N_15521,N_15073);
or U16255 (N_16255,N_15778,N_15227);
xor U16256 (N_16256,N_15912,N_15379);
or U16257 (N_16257,N_15782,N_15055);
nand U16258 (N_16258,N_15054,N_15262);
or U16259 (N_16259,N_15822,N_15808);
xnor U16260 (N_16260,N_15764,N_15277);
nor U16261 (N_16261,N_15542,N_15638);
nand U16262 (N_16262,N_15675,N_15101);
nand U16263 (N_16263,N_15619,N_15376);
or U16264 (N_16264,N_15414,N_15865);
nand U16265 (N_16265,N_15702,N_15669);
and U16266 (N_16266,N_15866,N_15204);
nor U16267 (N_16267,N_15048,N_15533);
and U16268 (N_16268,N_15564,N_15540);
nand U16269 (N_16269,N_15670,N_15957);
and U16270 (N_16270,N_15365,N_15419);
or U16271 (N_16271,N_15181,N_15927);
nand U16272 (N_16272,N_15121,N_15360);
xnor U16273 (N_16273,N_15122,N_15662);
nor U16274 (N_16274,N_15730,N_15826);
or U16275 (N_16275,N_15446,N_15491);
nor U16276 (N_16276,N_15103,N_15724);
nand U16277 (N_16277,N_15317,N_15838);
or U16278 (N_16278,N_15108,N_15626);
or U16279 (N_16279,N_15348,N_15324);
and U16280 (N_16280,N_15175,N_15235);
nand U16281 (N_16281,N_15282,N_15241);
nand U16282 (N_16282,N_15741,N_15328);
xnor U16283 (N_16283,N_15842,N_15206);
nand U16284 (N_16284,N_15886,N_15107);
and U16285 (N_16285,N_15056,N_15925);
nand U16286 (N_16286,N_15338,N_15523);
and U16287 (N_16287,N_15654,N_15615);
or U16288 (N_16288,N_15490,N_15940);
nor U16289 (N_16289,N_15258,N_15682);
xor U16290 (N_16290,N_15240,N_15385);
xnor U16291 (N_16291,N_15375,N_15297);
or U16292 (N_16292,N_15873,N_15721);
nor U16293 (N_16293,N_15574,N_15079);
xnor U16294 (N_16294,N_15285,N_15296);
nor U16295 (N_16295,N_15901,N_15725);
nand U16296 (N_16296,N_15085,N_15672);
xnor U16297 (N_16297,N_15747,N_15796);
and U16298 (N_16298,N_15420,N_15044);
and U16299 (N_16299,N_15677,N_15134);
nand U16300 (N_16300,N_15759,N_15416);
nor U16301 (N_16301,N_15504,N_15104);
nand U16302 (N_16302,N_15213,N_15335);
and U16303 (N_16303,N_15212,N_15713);
xor U16304 (N_16304,N_15855,N_15587);
nor U16305 (N_16305,N_15948,N_15025);
xnor U16306 (N_16306,N_15909,N_15045);
or U16307 (N_16307,N_15771,N_15380);
or U16308 (N_16308,N_15959,N_15456);
nand U16309 (N_16309,N_15661,N_15195);
nand U16310 (N_16310,N_15200,N_15075);
nor U16311 (N_16311,N_15187,N_15697);
or U16312 (N_16312,N_15370,N_15896);
xnor U16313 (N_16313,N_15330,N_15481);
or U16314 (N_16314,N_15478,N_15159);
or U16315 (N_16315,N_15528,N_15129);
or U16316 (N_16316,N_15663,N_15507);
and U16317 (N_16317,N_15276,N_15624);
nand U16318 (N_16318,N_15686,N_15894);
and U16319 (N_16319,N_15642,N_15298);
xor U16320 (N_16320,N_15062,N_15617);
nand U16321 (N_16321,N_15766,N_15286);
and U16322 (N_16322,N_15248,N_15274);
nor U16323 (N_16323,N_15188,N_15820);
or U16324 (N_16324,N_15174,N_15740);
nor U16325 (N_16325,N_15028,N_15841);
nand U16326 (N_16326,N_15094,N_15150);
xor U16327 (N_16327,N_15639,N_15719);
and U16328 (N_16328,N_15333,N_15133);
or U16329 (N_16329,N_15704,N_15636);
nor U16330 (N_16330,N_15602,N_15184);
and U16331 (N_16331,N_15727,N_15349);
xor U16332 (N_16332,N_15500,N_15278);
or U16333 (N_16333,N_15513,N_15525);
and U16334 (N_16334,N_15920,N_15846);
xor U16335 (N_16335,N_15155,N_15953);
nor U16336 (N_16336,N_15812,N_15515);
or U16337 (N_16337,N_15924,N_15160);
nand U16338 (N_16338,N_15116,N_15922);
and U16339 (N_16339,N_15634,N_15941);
and U16340 (N_16340,N_15608,N_15859);
xor U16341 (N_16341,N_15769,N_15066);
or U16342 (N_16342,N_15316,N_15984);
xnor U16343 (N_16343,N_15377,N_15334);
or U16344 (N_16344,N_15115,N_15962);
xnor U16345 (N_16345,N_15518,N_15329);
nand U16346 (N_16346,N_15620,N_15844);
nand U16347 (N_16347,N_15426,N_15548);
nor U16348 (N_16348,N_15265,N_15834);
nor U16349 (N_16349,N_15549,N_15678);
xor U16350 (N_16350,N_15251,N_15389);
nand U16351 (N_16351,N_15970,N_15580);
and U16352 (N_16352,N_15283,N_15135);
and U16353 (N_16353,N_15629,N_15791);
or U16354 (N_16354,N_15847,N_15650);
xnor U16355 (N_16355,N_15973,N_15463);
nand U16356 (N_16356,N_15148,N_15309);
nand U16357 (N_16357,N_15288,N_15685);
nand U16358 (N_16358,N_15412,N_15603);
nor U16359 (N_16359,N_15872,N_15680);
nor U16360 (N_16360,N_15561,N_15292);
or U16361 (N_16361,N_15890,N_15192);
xor U16362 (N_16362,N_15819,N_15318);
or U16363 (N_16363,N_15789,N_15488);
or U16364 (N_16364,N_15470,N_15963);
or U16365 (N_16365,N_15190,N_15754);
nand U16366 (N_16366,N_15097,N_15117);
or U16367 (N_16367,N_15060,N_15409);
and U16368 (N_16368,N_15314,N_15449);
and U16369 (N_16369,N_15594,N_15350);
and U16370 (N_16370,N_15688,N_15008);
or U16371 (N_16371,N_15367,N_15698);
or U16372 (N_16372,N_15832,N_15455);
nor U16373 (N_16373,N_15614,N_15595);
and U16374 (N_16374,N_15853,N_15990);
or U16375 (N_16375,N_15341,N_15736);
or U16376 (N_16376,N_15577,N_15483);
nand U16377 (N_16377,N_15706,N_15332);
and U16378 (N_16378,N_15280,N_15402);
nor U16379 (N_16379,N_15128,N_15106);
and U16380 (N_16380,N_15739,N_15731);
or U16381 (N_16381,N_15589,N_15664);
or U16382 (N_16382,N_15302,N_15788);
nor U16383 (N_16383,N_15908,N_15295);
nand U16384 (N_16384,N_15703,N_15911);
nor U16385 (N_16385,N_15239,N_15862);
xnor U16386 (N_16386,N_15985,N_15393);
and U16387 (N_16387,N_15609,N_15950);
and U16388 (N_16388,N_15173,N_15342);
nor U16389 (N_16389,N_15933,N_15510);
nand U16390 (N_16390,N_15432,N_15177);
xnor U16391 (N_16391,N_15058,N_15809);
nand U16392 (N_16392,N_15147,N_15918);
nand U16393 (N_16393,N_15023,N_15760);
nand U16394 (N_16394,N_15425,N_15534);
nor U16395 (N_16395,N_15969,N_15965);
nand U16396 (N_16396,N_15877,N_15057);
nor U16397 (N_16397,N_15254,N_15934);
or U16398 (N_16398,N_15454,N_15043);
or U16399 (N_16399,N_15021,N_15818);
nand U16400 (N_16400,N_15193,N_15668);
nand U16401 (N_16401,N_15585,N_15166);
or U16402 (N_16402,N_15566,N_15310);
nor U16403 (N_16403,N_15956,N_15230);
or U16404 (N_16404,N_15786,N_15651);
and U16405 (N_16405,N_15879,N_15471);
or U16406 (N_16406,N_15404,N_15344);
nand U16407 (N_16407,N_15499,N_15929);
and U16408 (N_16408,N_15308,N_15013);
xor U16409 (N_16409,N_15290,N_15266);
nor U16410 (N_16410,N_15773,N_15246);
nor U16411 (N_16411,N_15433,N_15337);
nand U16412 (N_16412,N_15583,N_15418);
xnor U16413 (N_16413,N_15484,N_15182);
and U16414 (N_16414,N_15524,N_15695);
xnor U16415 (N_16415,N_15136,N_15824);
xnor U16416 (N_16416,N_15201,N_15539);
nand U16417 (N_16417,N_15322,N_15709);
nor U16418 (N_16418,N_15516,N_15621);
nand U16419 (N_16419,N_15913,N_15217);
and U16420 (N_16420,N_15482,N_15026);
and U16421 (N_16421,N_15830,N_15363);
and U16422 (N_16422,N_15541,N_15093);
nand U16423 (N_16423,N_15229,N_15422);
nor U16424 (N_16424,N_15072,N_15627);
and U16425 (N_16425,N_15579,N_15221);
or U16426 (N_16426,N_15945,N_15428);
nor U16427 (N_16427,N_15225,N_15752);
nand U16428 (N_16428,N_15837,N_15156);
or U16429 (N_16429,N_15183,N_15343);
nand U16430 (N_16430,N_15671,N_15061);
or U16431 (N_16431,N_15140,N_15734);
or U16432 (N_16432,N_15014,N_15257);
nor U16433 (N_16433,N_15590,N_15951);
nor U16434 (N_16434,N_15194,N_15987);
and U16435 (N_16435,N_15720,N_15794);
or U16436 (N_16436,N_15458,N_15613);
and U16437 (N_16437,N_15445,N_15983);
nor U16438 (N_16438,N_15049,N_15269);
and U16439 (N_16439,N_15802,N_15487);
xnor U16440 (N_16440,N_15519,N_15787);
or U16441 (N_16441,N_15027,N_15749);
nor U16442 (N_16442,N_15673,N_15015);
or U16443 (N_16443,N_15164,N_15652);
nand U16444 (N_16444,N_15647,N_15068);
nand U16445 (N_16445,N_15750,N_15980);
nand U16446 (N_16446,N_15551,N_15657);
or U16447 (N_16447,N_15849,N_15681);
or U16448 (N_16448,N_15906,N_15928);
or U16449 (N_16449,N_15141,N_15569);
xor U16450 (N_16450,N_15170,N_15512);
nor U16451 (N_16451,N_15946,N_15785);
xnor U16452 (N_16452,N_15643,N_15726);
nand U16453 (N_16453,N_15947,N_15571);
nor U16454 (N_16454,N_15581,N_15131);
or U16455 (N_16455,N_15562,N_15010);
nand U16456 (N_16456,N_15696,N_15903);
nand U16457 (N_16457,N_15465,N_15228);
or U16458 (N_16458,N_15259,N_15477);
and U16459 (N_16459,N_15098,N_15030);
nand U16460 (N_16460,N_15867,N_15596);
and U16461 (N_16461,N_15790,N_15543);
xor U16462 (N_16462,N_15218,N_15382);
nand U16463 (N_16463,N_15080,N_15861);
or U16464 (N_16464,N_15814,N_15063);
nand U16465 (N_16465,N_15497,N_15763);
and U16466 (N_16466,N_15358,N_15907);
nor U16467 (N_16467,N_15584,N_15413);
nand U16468 (N_16468,N_15753,N_15139);
nand U16469 (N_16469,N_15991,N_15475);
nor U16470 (N_16470,N_15423,N_15883);
nor U16471 (N_16471,N_15914,N_15641);
nor U16472 (N_16472,N_15746,N_15253);
xnor U16473 (N_16473,N_15167,N_15768);
nor U16474 (N_16474,N_15374,N_15242);
xor U16475 (N_16475,N_15868,N_15707);
or U16476 (N_16476,N_15882,N_15421);
and U16477 (N_16477,N_15466,N_15109);
nor U16478 (N_16478,N_15742,N_15591);
xnor U16479 (N_16479,N_15035,N_15509);
nand U16480 (N_16480,N_15961,N_15784);
nand U16481 (N_16481,N_15299,N_15381);
nor U16482 (N_16482,N_15090,N_15084);
or U16483 (N_16483,N_15291,N_15394);
or U16484 (N_16484,N_15628,N_15816);
nor U16485 (N_16485,N_15099,N_15612);
or U16486 (N_16486,N_15252,N_15506);
nor U16487 (N_16487,N_15260,N_15018);
nor U16488 (N_16488,N_15053,N_15568);
xor U16489 (N_16489,N_15884,N_15447);
nand U16490 (N_16490,N_15124,N_15304);
nor U16491 (N_16491,N_15143,N_15999);
nor U16492 (N_16492,N_15127,N_15037);
or U16493 (N_16493,N_15993,N_15371);
or U16494 (N_16494,N_15226,N_15211);
nand U16495 (N_16495,N_15898,N_15495);
nand U16496 (N_16496,N_15392,N_15114);
or U16497 (N_16497,N_15390,N_15854);
or U16498 (N_16498,N_15813,N_15207);
and U16499 (N_16499,N_15462,N_15538);
or U16500 (N_16500,N_15595,N_15419);
and U16501 (N_16501,N_15758,N_15549);
xor U16502 (N_16502,N_15062,N_15338);
or U16503 (N_16503,N_15241,N_15610);
nor U16504 (N_16504,N_15142,N_15864);
nand U16505 (N_16505,N_15876,N_15970);
or U16506 (N_16506,N_15306,N_15237);
nor U16507 (N_16507,N_15959,N_15233);
xor U16508 (N_16508,N_15844,N_15866);
or U16509 (N_16509,N_15436,N_15097);
nor U16510 (N_16510,N_15526,N_15310);
nand U16511 (N_16511,N_15778,N_15551);
and U16512 (N_16512,N_15893,N_15253);
nor U16513 (N_16513,N_15189,N_15152);
nand U16514 (N_16514,N_15933,N_15418);
nor U16515 (N_16515,N_15227,N_15191);
nand U16516 (N_16516,N_15364,N_15590);
and U16517 (N_16517,N_15075,N_15860);
nand U16518 (N_16518,N_15483,N_15299);
xnor U16519 (N_16519,N_15989,N_15260);
xor U16520 (N_16520,N_15727,N_15340);
nor U16521 (N_16521,N_15771,N_15238);
or U16522 (N_16522,N_15214,N_15082);
nor U16523 (N_16523,N_15121,N_15128);
and U16524 (N_16524,N_15130,N_15987);
nor U16525 (N_16525,N_15377,N_15684);
nand U16526 (N_16526,N_15686,N_15013);
and U16527 (N_16527,N_15638,N_15227);
nand U16528 (N_16528,N_15580,N_15811);
nand U16529 (N_16529,N_15222,N_15025);
or U16530 (N_16530,N_15999,N_15772);
nand U16531 (N_16531,N_15860,N_15458);
nand U16532 (N_16532,N_15737,N_15116);
and U16533 (N_16533,N_15339,N_15470);
xor U16534 (N_16534,N_15572,N_15777);
or U16535 (N_16535,N_15935,N_15497);
and U16536 (N_16536,N_15867,N_15215);
nand U16537 (N_16537,N_15898,N_15670);
and U16538 (N_16538,N_15866,N_15671);
or U16539 (N_16539,N_15664,N_15128);
nor U16540 (N_16540,N_15299,N_15705);
xor U16541 (N_16541,N_15450,N_15493);
or U16542 (N_16542,N_15248,N_15095);
nor U16543 (N_16543,N_15141,N_15422);
nand U16544 (N_16544,N_15176,N_15963);
or U16545 (N_16545,N_15920,N_15079);
and U16546 (N_16546,N_15298,N_15216);
nor U16547 (N_16547,N_15288,N_15988);
xnor U16548 (N_16548,N_15394,N_15166);
xnor U16549 (N_16549,N_15051,N_15293);
xnor U16550 (N_16550,N_15158,N_15842);
nand U16551 (N_16551,N_15277,N_15011);
nor U16552 (N_16552,N_15313,N_15576);
nor U16553 (N_16553,N_15540,N_15129);
nor U16554 (N_16554,N_15601,N_15884);
nor U16555 (N_16555,N_15777,N_15260);
xor U16556 (N_16556,N_15348,N_15007);
nor U16557 (N_16557,N_15917,N_15389);
xor U16558 (N_16558,N_15990,N_15837);
or U16559 (N_16559,N_15574,N_15985);
nand U16560 (N_16560,N_15197,N_15020);
nor U16561 (N_16561,N_15477,N_15522);
and U16562 (N_16562,N_15580,N_15692);
and U16563 (N_16563,N_15187,N_15779);
or U16564 (N_16564,N_15903,N_15948);
and U16565 (N_16565,N_15304,N_15680);
nor U16566 (N_16566,N_15583,N_15958);
nor U16567 (N_16567,N_15864,N_15645);
xnor U16568 (N_16568,N_15388,N_15358);
and U16569 (N_16569,N_15970,N_15672);
or U16570 (N_16570,N_15947,N_15685);
xnor U16571 (N_16571,N_15102,N_15684);
nor U16572 (N_16572,N_15218,N_15174);
xnor U16573 (N_16573,N_15596,N_15420);
and U16574 (N_16574,N_15940,N_15715);
xnor U16575 (N_16575,N_15252,N_15231);
xor U16576 (N_16576,N_15254,N_15164);
nand U16577 (N_16577,N_15317,N_15571);
or U16578 (N_16578,N_15995,N_15447);
or U16579 (N_16579,N_15874,N_15174);
or U16580 (N_16580,N_15753,N_15963);
and U16581 (N_16581,N_15603,N_15281);
nor U16582 (N_16582,N_15452,N_15345);
xor U16583 (N_16583,N_15481,N_15747);
nand U16584 (N_16584,N_15350,N_15328);
nand U16585 (N_16585,N_15986,N_15381);
or U16586 (N_16586,N_15198,N_15953);
or U16587 (N_16587,N_15005,N_15249);
or U16588 (N_16588,N_15610,N_15062);
nand U16589 (N_16589,N_15420,N_15256);
xor U16590 (N_16590,N_15151,N_15375);
nor U16591 (N_16591,N_15866,N_15225);
and U16592 (N_16592,N_15115,N_15023);
nand U16593 (N_16593,N_15908,N_15155);
nor U16594 (N_16594,N_15340,N_15725);
or U16595 (N_16595,N_15968,N_15400);
nor U16596 (N_16596,N_15266,N_15031);
or U16597 (N_16597,N_15641,N_15251);
or U16598 (N_16598,N_15130,N_15386);
xor U16599 (N_16599,N_15984,N_15841);
nor U16600 (N_16600,N_15673,N_15607);
nand U16601 (N_16601,N_15085,N_15977);
nor U16602 (N_16602,N_15463,N_15432);
or U16603 (N_16603,N_15332,N_15417);
or U16604 (N_16604,N_15408,N_15462);
nand U16605 (N_16605,N_15936,N_15421);
nand U16606 (N_16606,N_15551,N_15080);
and U16607 (N_16607,N_15580,N_15924);
nand U16608 (N_16608,N_15085,N_15359);
nor U16609 (N_16609,N_15628,N_15745);
and U16610 (N_16610,N_15999,N_15268);
and U16611 (N_16611,N_15446,N_15158);
or U16612 (N_16612,N_15139,N_15510);
xor U16613 (N_16613,N_15741,N_15816);
and U16614 (N_16614,N_15446,N_15732);
nand U16615 (N_16615,N_15295,N_15208);
xnor U16616 (N_16616,N_15916,N_15307);
nand U16617 (N_16617,N_15084,N_15220);
or U16618 (N_16618,N_15649,N_15287);
xnor U16619 (N_16619,N_15050,N_15760);
and U16620 (N_16620,N_15830,N_15806);
and U16621 (N_16621,N_15772,N_15209);
nand U16622 (N_16622,N_15248,N_15600);
xor U16623 (N_16623,N_15377,N_15575);
xor U16624 (N_16624,N_15738,N_15720);
xnor U16625 (N_16625,N_15373,N_15214);
nand U16626 (N_16626,N_15034,N_15789);
nor U16627 (N_16627,N_15016,N_15191);
nor U16628 (N_16628,N_15844,N_15630);
and U16629 (N_16629,N_15249,N_15786);
xnor U16630 (N_16630,N_15864,N_15767);
or U16631 (N_16631,N_15116,N_15764);
and U16632 (N_16632,N_15463,N_15038);
nand U16633 (N_16633,N_15328,N_15600);
nand U16634 (N_16634,N_15549,N_15646);
xnor U16635 (N_16635,N_15053,N_15955);
nor U16636 (N_16636,N_15664,N_15878);
or U16637 (N_16637,N_15309,N_15429);
nor U16638 (N_16638,N_15073,N_15536);
nand U16639 (N_16639,N_15422,N_15349);
and U16640 (N_16640,N_15983,N_15663);
xor U16641 (N_16641,N_15473,N_15891);
or U16642 (N_16642,N_15217,N_15931);
nor U16643 (N_16643,N_15174,N_15815);
or U16644 (N_16644,N_15316,N_15675);
and U16645 (N_16645,N_15319,N_15598);
or U16646 (N_16646,N_15503,N_15821);
or U16647 (N_16647,N_15506,N_15572);
or U16648 (N_16648,N_15223,N_15297);
or U16649 (N_16649,N_15434,N_15342);
nor U16650 (N_16650,N_15272,N_15584);
nor U16651 (N_16651,N_15015,N_15526);
nand U16652 (N_16652,N_15314,N_15386);
or U16653 (N_16653,N_15251,N_15031);
and U16654 (N_16654,N_15320,N_15908);
or U16655 (N_16655,N_15692,N_15914);
nor U16656 (N_16656,N_15245,N_15456);
and U16657 (N_16657,N_15922,N_15768);
nor U16658 (N_16658,N_15463,N_15397);
nor U16659 (N_16659,N_15055,N_15602);
xnor U16660 (N_16660,N_15987,N_15442);
and U16661 (N_16661,N_15386,N_15644);
xnor U16662 (N_16662,N_15069,N_15570);
nor U16663 (N_16663,N_15028,N_15370);
nor U16664 (N_16664,N_15596,N_15721);
xnor U16665 (N_16665,N_15827,N_15809);
nor U16666 (N_16666,N_15178,N_15837);
nor U16667 (N_16667,N_15262,N_15071);
nand U16668 (N_16668,N_15665,N_15419);
and U16669 (N_16669,N_15137,N_15848);
xnor U16670 (N_16670,N_15765,N_15154);
or U16671 (N_16671,N_15454,N_15164);
nor U16672 (N_16672,N_15629,N_15192);
nand U16673 (N_16673,N_15290,N_15483);
nor U16674 (N_16674,N_15496,N_15326);
and U16675 (N_16675,N_15640,N_15612);
and U16676 (N_16676,N_15060,N_15399);
and U16677 (N_16677,N_15394,N_15783);
nor U16678 (N_16678,N_15787,N_15009);
and U16679 (N_16679,N_15864,N_15502);
or U16680 (N_16680,N_15029,N_15542);
xnor U16681 (N_16681,N_15037,N_15741);
xor U16682 (N_16682,N_15719,N_15406);
nand U16683 (N_16683,N_15064,N_15131);
and U16684 (N_16684,N_15151,N_15085);
nor U16685 (N_16685,N_15614,N_15054);
nor U16686 (N_16686,N_15295,N_15608);
or U16687 (N_16687,N_15060,N_15665);
xor U16688 (N_16688,N_15008,N_15907);
or U16689 (N_16689,N_15041,N_15314);
nand U16690 (N_16690,N_15579,N_15462);
nand U16691 (N_16691,N_15598,N_15736);
or U16692 (N_16692,N_15932,N_15180);
nand U16693 (N_16693,N_15713,N_15489);
nand U16694 (N_16694,N_15192,N_15757);
nor U16695 (N_16695,N_15840,N_15317);
or U16696 (N_16696,N_15910,N_15483);
and U16697 (N_16697,N_15958,N_15418);
nor U16698 (N_16698,N_15318,N_15553);
xor U16699 (N_16699,N_15488,N_15699);
xnor U16700 (N_16700,N_15543,N_15373);
nand U16701 (N_16701,N_15485,N_15653);
nor U16702 (N_16702,N_15911,N_15485);
and U16703 (N_16703,N_15588,N_15484);
nor U16704 (N_16704,N_15942,N_15453);
xor U16705 (N_16705,N_15094,N_15696);
or U16706 (N_16706,N_15361,N_15521);
nand U16707 (N_16707,N_15709,N_15160);
and U16708 (N_16708,N_15601,N_15927);
nor U16709 (N_16709,N_15340,N_15974);
nor U16710 (N_16710,N_15251,N_15437);
and U16711 (N_16711,N_15499,N_15079);
xnor U16712 (N_16712,N_15898,N_15139);
nand U16713 (N_16713,N_15340,N_15394);
xnor U16714 (N_16714,N_15831,N_15643);
nor U16715 (N_16715,N_15244,N_15995);
nor U16716 (N_16716,N_15098,N_15780);
and U16717 (N_16717,N_15385,N_15488);
and U16718 (N_16718,N_15264,N_15792);
xnor U16719 (N_16719,N_15118,N_15386);
xnor U16720 (N_16720,N_15100,N_15834);
and U16721 (N_16721,N_15899,N_15227);
or U16722 (N_16722,N_15719,N_15085);
or U16723 (N_16723,N_15986,N_15161);
nand U16724 (N_16724,N_15900,N_15661);
xnor U16725 (N_16725,N_15177,N_15851);
nor U16726 (N_16726,N_15696,N_15150);
or U16727 (N_16727,N_15029,N_15747);
and U16728 (N_16728,N_15343,N_15218);
and U16729 (N_16729,N_15916,N_15403);
nor U16730 (N_16730,N_15405,N_15393);
nand U16731 (N_16731,N_15549,N_15187);
xor U16732 (N_16732,N_15073,N_15423);
nand U16733 (N_16733,N_15371,N_15763);
xnor U16734 (N_16734,N_15089,N_15000);
xor U16735 (N_16735,N_15523,N_15620);
or U16736 (N_16736,N_15973,N_15630);
nand U16737 (N_16737,N_15512,N_15736);
and U16738 (N_16738,N_15944,N_15278);
xnor U16739 (N_16739,N_15116,N_15757);
xor U16740 (N_16740,N_15759,N_15002);
and U16741 (N_16741,N_15181,N_15670);
nand U16742 (N_16742,N_15255,N_15807);
nand U16743 (N_16743,N_15984,N_15916);
or U16744 (N_16744,N_15522,N_15399);
xnor U16745 (N_16745,N_15550,N_15223);
or U16746 (N_16746,N_15793,N_15573);
or U16747 (N_16747,N_15705,N_15450);
xnor U16748 (N_16748,N_15251,N_15093);
nor U16749 (N_16749,N_15424,N_15831);
nand U16750 (N_16750,N_15776,N_15181);
nand U16751 (N_16751,N_15078,N_15848);
xor U16752 (N_16752,N_15750,N_15114);
xnor U16753 (N_16753,N_15672,N_15920);
xor U16754 (N_16754,N_15687,N_15004);
nand U16755 (N_16755,N_15896,N_15529);
or U16756 (N_16756,N_15443,N_15957);
xor U16757 (N_16757,N_15131,N_15779);
xnor U16758 (N_16758,N_15490,N_15510);
xnor U16759 (N_16759,N_15055,N_15091);
xor U16760 (N_16760,N_15752,N_15569);
nand U16761 (N_16761,N_15100,N_15986);
and U16762 (N_16762,N_15466,N_15903);
nand U16763 (N_16763,N_15419,N_15126);
xnor U16764 (N_16764,N_15872,N_15194);
nand U16765 (N_16765,N_15171,N_15974);
and U16766 (N_16766,N_15243,N_15382);
or U16767 (N_16767,N_15283,N_15126);
and U16768 (N_16768,N_15915,N_15343);
nand U16769 (N_16769,N_15505,N_15411);
xnor U16770 (N_16770,N_15208,N_15111);
and U16771 (N_16771,N_15881,N_15790);
nor U16772 (N_16772,N_15562,N_15529);
nand U16773 (N_16773,N_15085,N_15056);
and U16774 (N_16774,N_15358,N_15886);
and U16775 (N_16775,N_15395,N_15365);
nand U16776 (N_16776,N_15930,N_15033);
and U16777 (N_16777,N_15283,N_15076);
and U16778 (N_16778,N_15565,N_15210);
nor U16779 (N_16779,N_15185,N_15838);
nand U16780 (N_16780,N_15441,N_15965);
or U16781 (N_16781,N_15573,N_15766);
and U16782 (N_16782,N_15358,N_15748);
or U16783 (N_16783,N_15625,N_15857);
nor U16784 (N_16784,N_15015,N_15012);
nor U16785 (N_16785,N_15786,N_15457);
and U16786 (N_16786,N_15607,N_15444);
and U16787 (N_16787,N_15578,N_15374);
nand U16788 (N_16788,N_15842,N_15697);
nor U16789 (N_16789,N_15782,N_15339);
and U16790 (N_16790,N_15007,N_15037);
nor U16791 (N_16791,N_15509,N_15748);
xnor U16792 (N_16792,N_15452,N_15009);
nor U16793 (N_16793,N_15534,N_15552);
xor U16794 (N_16794,N_15237,N_15765);
nor U16795 (N_16795,N_15805,N_15985);
nand U16796 (N_16796,N_15079,N_15113);
or U16797 (N_16797,N_15655,N_15421);
xnor U16798 (N_16798,N_15883,N_15240);
nor U16799 (N_16799,N_15960,N_15900);
and U16800 (N_16800,N_15461,N_15065);
or U16801 (N_16801,N_15205,N_15656);
nor U16802 (N_16802,N_15424,N_15417);
xor U16803 (N_16803,N_15024,N_15235);
nor U16804 (N_16804,N_15281,N_15154);
nor U16805 (N_16805,N_15929,N_15712);
or U16806 (N_16806,N_15828,N_15756);
and U16807 (N_16807,N_15568,N_15679);
nand U16808 (N_16808,N_15726,N_15945);
or U16809 (N_16809,N_15389,N_15524);
and U16810 (N_16810,N_15913,N_15270);
xnor U16811 (N_16811,N_15202,N_15234);
and U16812 (N_16812,N_15032,N_15750);
nand U16813 (N_16813,N_15286,N_15656);
xnor U16814 (N_16814,N_15822,N_15228);
xor U16815 (N_16815,N_15462,N_15620);
nor U16816 (N_16816,N_15713,N_15897);
nor U16817 (N_16817,N_15063,N_15025);
and U16818 (N_16818,N_15126,N_15545);
or U16819 (N_16819,N_15774,N_15058);
or U16820 (N_16820,N_15199,N_15732);
nand U16821 (N_16821,N_15796,N_15052);
nand U16822 (N_16822,N_15067,N_15717);
and U16823 (N_16823,N_15723,N_15483);
or U16824 (N_16824,N_15979,N_15910);
nand U16825 (N_16825,N_15234,N_15349);
or U16826 (N_16826,N_15307,N_15889);
nand U16827 (N_16827,N_15517,N_15160);
nand U16828 (N_16828,N_15239,N_15679);
and U16829 (N_16829,N_15588,N_15922);
nand U16830 (N_16830,N_15317,N_15537);
or U16831 (N_16831,N_15275,N_15370);
and U16832 (N_16832,N_15397,N_15985);
and U16833 (N_16833,N_15330,N_15680);
and U16834 (N_16834,N_15167,N_15304);
nor U16835 (N_16835,N_15805,N_15979);
and U16836 (N_16836,N_15109,N_15013);
or U16837 (N_16837,N_15053,N_15362);
nor U16838 (N_16838,N_15726,N_15846);
xnor U16839 (N_16839,N_15457,N_15237);
or U16840 (N_16840,N_15338,N_15585);
and U16841 (N_16841,N_15283,N_15684);
nor U16842 (N_16842,N_15951,N_15450);
nand U16843 (N_16843,N_15779,N_15501);
nand U16844 (N_16844,N_15446,N_15106);
or U16845 (N_16845,N_15076,N_15861);
and U16846 (N_16846,N_15164,N_15287);
nor U16847 (N_16847,N_15786,N_15251);
xnor U16848 (N_16848,N_15280,N_15062);
nor U16849 (N_16849,N_15223,N_15106);
nor U16850 (N_16850,N_15680,N_15763);
nor U16851 (N_16851,N_15113,N_15408);
and U16852 (N_16852,N_15141,N_15513);
nor U16853 (N_16853,N_15543,N_15033);
or U16854 (N_16854,N_15514,N_15854);
xor U16855 (N_16855,N_15978,N_15990);
xnor U16856 (N_16856,N_15130,N_15218);
xor U16857 (N_16857,N_15382,N_15981);
and U16858 (N_16858,N_15227,N_15755);
nand U16859 (N_16859,N_15884,N_15844);
nor U16860 (N_16860,N_15945,N_15027);
xor U16861 (N_16861,N_15262,N_15250);
and U16862 (N_16862,N_15941,N_15189);
or U16863 (N_16863,N_15960,N_15118);
xnor U16864 (N_16864,N_15532,N_15705);
nor U16865 (N_16865,N_15376,N_15430);
and U16866 (N_16866,N_15030,N_15488);
nor U16867 (N_16867,N_15300,N_15358);
and U16868 (N_16868,N_15578,N_15647);
xor U16869 (N_16869,N_15589,N_15360);
or U16870 (N_16870,N_15697,N_15952);
or U16871 (N_16871,N_15413,N_15532);
nor U16872 (N_16872,N_15599,N_15657);
nand U16873 (N_16873,N_15920,N_15396);
nor U16874 (N_16874,N_15347,N_15808);
xor U16875 (N_16875,N_15260,N_15262);
or U16876 (N_16876,N_15542,N_15633);
nor U16877 (N_16877,N_15053,N_15959);
or U16878 (N_16878,N_15936,N_15197);
or U16879 (N_16879,N_15545,N_15049);
or U16880 (N_16880,N_15841,N_15471);
and U16881 (N_16881,N_15481,N_15990);
nand U16882 (N_16882,N_15358,N_15727);
nor U16883 (N_16883,N_15309,N_15944);
xor U16884 (N_16884,N_15346,N_15369);
nand U16885 (N_16885,N_15942,N_15731);
xor U16886 (N_16886,N_15303,N_15201);
nand U16887 (N_16887,N_15002,N_15244);
xor U16888 (N_16888,N_15291,N_15384);
or U16889 (N_16889,N_15206,N_15066);
xor U16890 (N_16890,N_15350,N_15612);
nor U16891 (N_16891,N_15803,N_15708);
nor U16892 (N_16892,N_15617,N_15934);
nor U16893 (N_16893,N_15710,N_15089);
xor U16894 (N_16894,N_15267,N_15255);
or U16895 (N_16895,N_15164,N_15096);
nand U16896 (N_16896,N_15384,N_15134);
and U16897 (N_16897,N_15348,N_15932);
xor U16898 (N_16898,N_15868,N_15947);
xor U16899 (N_16899,N_15308,N_15526);
and U16900 (N_16900,N_15756,N_15333);
xnor U16901 (N_16901,N_15801,N_15653);
xor U16902 (N_16902,N_15043,N_15429);
nand U16903 (N_16903,N_15861,N_15707);
nor U16904 (N_16904,N_15916,N_15847);
or U16905 (N_16905,N_15633,N_15223);
nor U16906 (N_16906,N_15034,N_15223);
xor U16907 (N_16907,N_15208,N_15552);
or U16908 (N_16908,N_15247,N_15205);
xor U16909 (N_16909,N_15039,N_15203);
and U16910 (N_16910,N_15960,N_15413);
nand U16911 (N_16911,N_15405,N_15648);
or U16912 (N_16912,N_15628,N_15096);
or U16913 (N_16913,N_15416,N_15561);
xnor U16914 (N_16914,N_15658,N_15724);
or U16915 (N_16915,N_15488,N_15162);
xor U16916 (N_16916,N_15182,N_15839);
nand U16917 (N_16917,N_15888,N_15495);
or U16918 (N_16918,N_15825,N_15922);
nor U16919 (N_16919,N_15572,N_15494);
and U16920 (N_16920,N_15885,N_15664);
or U16921 (N_16921,N_15386,N_15248);
nor U16922 (N_16922,N_15869,N_15653);
and U16923 (N_16923,N_15832,N_15695);
xnor U16924 (N_16924,N_15232,N_15793);
and U16925 (N_16925,N_15642,N_15024);
nand U16926 (N_16926,N_15944,N_15665);
or U16927 (N_16927,N_15679,N_15691);
and U16928 (N_16928,N_15795,N_15361);
nand U16929 (N_16929,N_15364,N_15846);
or U16930 (N_16930,N_15882,N_15418);
and U16931 (N_16931,N_15624,N_15563);
nand U16932 (N_16932,N_15415,N_15681);
nor U16933 (N_16933,N_15661,N_15497);
or U16934 (N_16934,N_15343,N_15806);
nor U16935 (N_16935,N_15971,N_15807);
and U16936 (N_16936,N_15735,N_15593);
and U16937 (N_16937,N_15338,N_15491);
nand U16938 (N_16938,N_15692,N_15094);
nor U16939 (N_16939,N_15872,N_15444);
nand U16940 (N_16940,N_15056,N_15132);
nand U16941 (N_16941,N_15171,N_15519);
and U16942 (N_16942,N_15081,N_15788);
nor U16943 (N_16943,N_15551,N_15580);
xnor U16944 (N_16944,N_15844,N_15179);
nand U16945 (N_16945,N_15368,N_15765);
or U16946 (N_16946,N_15704,N_15080);
xor U16947 (N_16947,N_15808,N_15362);
nor U16948 (N_16948,N_15371,N_15216);
or U16949 (N_16949,N_15714,N_15088);
nand U16950 (N_16950,N_15756,N_15924);
nand U16951 (N_16951,N_15906,N_15099);
or U16952 (N_16952,N_15778,N_15649);
xor U16953 (N_16953,N_15226,N_15959);
nand U16954 (N_16954,N_15263,N_15557);
and U16955 (N_16955,N_15966,N_15879);
xor U16956 (N_16956,N_15837,N_15667);
or U16957 (N_16957,N_15069,N_15358);
nor U16958 (N_16958,N_15620,N_15107);
or U16959 (N_16959,N_15729,N_15976);
xnor U16960 (N_16960,N_15768,N_15924);
xnor U16961 (N_16961,N_15397,N_15782);
or U16962 (N_16962,N_15595,N_15734);
or U16963 (N_16963,N_15951,N_15941);
and U16964 (N_16964,N_15213,N_15013);
or U16965 (N_16965,N_15260,N_15569);
or U16966 (N_16966,N_15083,N_15498);
and U16967 (N_16967,N_15722,N_15769);
and U16968 (N_16968,N_15433,N_15693);
nand U16969 (N_16969,N_15872,N_15458);
nor U16970 (N_16970,N_15733,N_15677);
xor U16971 (N_16971,N_15049,N_15528);
nand U16972 (N_16972,N_15523,N_15763);
or U16973 (N_16973,N_15525,N_15518);
nand U16974 (N_16974,N_15966,N_15853);
or U16975 (N_16975,N_15010,N_15715);
nor U16976 (N_16976,N_15650,N_15459);
xor U16977 (N_16977,N_15446,N_15238);
nand U16978 (N_16978,N_15291,N_15252);
nand U16979 (N_16979,N_15112,N_15570);
nand U16980 (N_16980,N_15803,N_15106);
nand U16981 (N_16981,N_15585,N_15325);
xor U16982 (N_16982,N_15127,N_15101);
or U16983 (N_16983,N_15325,N_15787);
or U16984 (N_16984,N_15191,N_15047);
or U16985 (N_16985,N_15208,N_15044);
nand U16986 (N_16986,N_15032,N_15323);
nor U16987 (N_16987,N_15963,N_15706);
xor U16988 (N_16988,N_15488,N_15313);
nor U16989 (N_16989,N_15431,N_15178);
and U16990 (N_16990,N_15005,N_15671);
or U16991 (N_16991,N_15519,N_15880);
or U16992 (N_16992,N_15145,N_15048);
nand U16993 (N_16993,N_15405,N_15330);
xnor U16994 (N_16994,N_15759,N_15613);
and U16995 (N_16995,N_15320,N_15998);
xor U16996 (N_16996,N_15751,N_15986);
nor U16997 (N_16997,N_15176,N_15165);
or U16998 (N_16998,N_15322,N_15984);
nor U16999 (N_16999,N_15916,N_15965);
nand U17000 (N_17000,N_16228,N_16757);
nand U17001 (N_17001,N_16151,N_16802);
nor U17002 (N_17002,N_16898,N_16128);
nand U17003 (N_17003,N_16311,N_16369);
xnor U17004 (N_17004,N_16753,N_16696);
or U17005 (N_17005,N_16784,N_16471);
xor U17006 (N_17006,N_16506,N_16177);
or U17007 (N_17007,N_16928,N_16601);
nor U17008 (N_17008,N_16965,N_16908);
xor U17009 (N_17009,N_16521,N_16457);
and U17010 (N_17010,N_16640,N_16192);
nand U17011 (N_17011,N_16490,N_16671);
nand U17012 (N_17012,N_16948,N_16257);
xor U17013 (N_17013,N_16466,N_16312);
nor U17014 (N_17014,N_16609,N_16843);
nand U17015 (N_17015,N_16256,N_16786);
nor U17016 (N_17016,N_16858,N_16031);
nand U17017 (N_17017,N_16867,N_16193);
nor U17018 (N_17018,N_16752,N_16015);
or U17019 (N_17019,N_16452,N_16921);
and U17020 (N_17020,N_16517,N_16206);
and U17021 (N_17021,N_16902,N_16258);
and U17022 (N_17022,N_16191,N_16366);
or U17023 (N_17023,N_16040,N_16890);
nor U17024 (N_17024,N_16555,N_16404);
and U17025 (N_17025,N_16895,N_16087);
or U17026 (N_17026,N_16994,N_16028);
and U17027 (N_17027,N_16263,N_16230);
or U17028 (N_17028,N_16590,N_16959);
nand U17029 (N_17029,N_16243,N_16475);
or U17030 (N_17030,N_16787,N_16726);
and U17031 (N_17031,N_16350,N_16387);
nor U17032 (N_17032,N_16358,N_16016);
and U17033 (N_17033,N_16109,N_16134);
or U17034 (N_17034,N_16832,N_16045);
or U17035 (N_17035,N_16712,N_16096);
and U17036 (N_17036,N_16957,N_16659);
or U17037 (N_17037,N_16493,N_16770);
and U17038 (N_17038,N_16993,N_16054);
or U17039 (N_17039,N_16344,N_16660);
nor U17040 (N_17040,N_16581,N_16967);
nand U17041 (N_17041,N_16587,N_16478);
nor U17042 (N_17042,N_16981,N_16773);
or U17043 (N_17043,N_16060,N_16329);
nand U17044 (N_17044,N_16918,N_16767);
xor U17045 (N_17045,N_16069,N_16132);
and U17046 (N_17046,N_16279,N_16951);
nand U17047 (N_17047,N_16942,N_16064);
nand U17048 (N_17048,N_16322,N_16864);
nand U17049 (N_17049,N_16120,N_16670);
or U17050 (N_17050,N_16063,N_16630);
or U17051 (N_17051,N_16771,N_16719);
nor U17052 (N_17052,N_16023,N_16791);
nand U17053 (N_17053,N_16524,N_16997);
or U17054 (N_17054,N_16084,N_16025);
nor U17055 (N_17055,N_16731,N_16481);
nand U17056 (N_17056,N_16042,N_16920);
nor U17057 (N_17057,N_16463,N_16559);
or U17058 (N_17058,N_16769,N_16812);
and U17059 (N_17059,N_16224,N_16533);
xnor U17060 (N_17060,N_16716,N_16205);
or U17061 (N_17061,N_16221,N_16119);
nand U17062 (N_17062,N_16455,N_16852);
and U17063 (N_17063,N_16187,N_16778);
nor U17064 (N_17064,N_16672,N_16302);
or U17065 (N_17065,N_16354,N_16952);
xnor U17066 (N_17066,N_16090,N_16764);
and U17067 (N_17067,N_16372,N_16596);
nand U17068 (N_17068,N_16103,N_16605);
xnor U17069 (N_17069,N_16241,N_16627);
xnor U17070 (N_17070,N_16085,N_16112);
xor U17071 (N_17071,N_16698,N_16511);
or U17072 (N_17072,N_16901,N_16472);
xnor U17073 (N_17073,N_16116,N_16435);
and U17074 (N_17074,N_16557,N_16909);
and U17075 (N_17075,N_16600,N_16580);
nand U17076 (N_17076,N_16208,N_16628);
xnor U17077 (N_17077,N_16088,N_16652);
nor U17078 (N_17078,N_16343,N_16202);
nor U17079 (N_17079,N_16785,N_16926);
nand U17080 (N_17080,N_16199,N_16484);
xnor U17081 (N_17081,N_16092,N_16695);
xnor U17082 (N_17082,N_16197,N_16178);
xor U17083 (N_17083,N_16968,N_16098);
and U17084 (N_17084,N_16700,N_16138);
nand U17085 (N_17085,N_16974,N_16891);
or U17086 (N_17086,N_16247,N_16080);
and U17087 (N_17087,N_16528,N_16194);
and U17088 (N_17088,N_16516,N_16795);
and U17089 (N_17089,N_16711,N_16339);
nor U17090 (N_17090,N_16223,N_16518);
or U17091 (N_17091,N_16743,N_16548);
or U17092 (N_17092,N_16393,N_16415);
nand U17093 (N_17093,N_16888,N_16604);
xor U17094 (N_17094,N_16474,N_16978);
xnor U17095 (N_17095,N_16639,N_16992);
xnor U17096 (N_17096,N_16419,N_16094);
xor U17097 (N_17097,N_16827,N_16488);
xor U17098 (N_17098,N_16610,N_16410);
and U17099 (N_17099,N_16411,N_16447);
xor U17100 (N_17100,N_16856,N_16677);
and U17101 (N_17101,N_16765,N_16004);
or U17102 (N_17102,N_16741,N_16621);
or U17103 (N_17103,N_16229,N_16730);
xnor U17104 (N_17104,N_16385,N_16991);
xnor U17105 (N_17105,N_16577,N_16146);
nand U17106 (N_17106,N_16217,N_16725);
nor U17107 (N_17107,N_16955,N_16983);
or U17108 (N_17108,N_16445,N_16267);
and U17109 (N_17109,N_16568,N_16531);
and U17110 (N_17110,N_16878,N_16550);
and U17111 (N_17111,N_16270,N_16656);
xnor U17112 (N_17112,N_16790,N_16772);
or U17113 (N_17113,N_16136,N_16564);
or U17114 (N_17114,N_16530,N_16966);
nor U17115 (N_17115,N_16851,N_16091);
xor U17116 (N_17116,N_16995,N_16275);
nand U17117 (N_17117,N_16813,N_16546);
or U17118 (N_17118,N_16566,N_16514);
nor U17119 (N_17119,N_16391,N_16699);
nor U17120 (N_17120,N_16181,N_16917);
nand U17121 (N_17121,N_16664,N_16880);
xnor U17122 (N_17122,N_16746,N_16924);
or U17123 (N_17123,N_16265,N_16056);
nor U17124 (N_17124,N_16195,N_16417);
nor U17125 (N_17125,N_16465,N_16857);
nand U17126 (N_17126,N_16125,N_16051);
nand U17127 (N_17127,N_16383,N_16907);
nand U17128 (N_17128,N_16883,N_16847);
and U17129 (N_17129,N_16459,N_16451);
nand U17130 (N_17130,N_16936,N_16705);
nor U17131 (N_17131,N_16346,N_16406);
and U17132 (N_17132,N_16689,N_16432);
and U17133 (N_17133,N_16482,N_16496);
and U17134 (N_17134,N_16844,N_16048);
xor U17135 (N_17135,N_16853,N_16649);
nor U17136 (N_17136,N_16044,N_16029);
nand U17137 (N_17137,N_16817,N_16688);
xor U17138 (N_17138,N_16253,N_16101);
or U17139 (N_17139,N_16710,N_16958);
nand U17140 (N_17140,N_16180,N_16246);
nand U17141 (N_17141,N_16122,N_16427);
nand U17142 (N_17142,N_16848,N_16830);
nand U17143 (N_17143,N_16679,N_16295);
or U17144 (N_17144,N_16733,N_16375);
xnor U17145 (N_17145,N_16681,N_16248);
nor U17146 (N_17146,N_16473,N_16763);
nand U17147 (N_17147,N_16704,N_16495);
xnor U17148 (N_17148,N_16569,N_16519);
nand U17149 (N_17149,N_16632,N_16058);
and U17150 (N_17150,N_16131,N_16829);
xor U17151 (N_17151,N_16422,N_16439);
and U17152 (N_17152,N_16794,N_16359);
nor U17153 (N_17153,N_16776,N_16026);
nand U17154 (N_17154,N_16185,N_16617);
nand U17155 (N_17155,N_16616,N_16460);
and U17156 (N_17156,N_16803,N_16884);
xnor U17157 (N_17157,N_16624,N_16603);
xor U17158 (N_17158,N_16130,N_16446);
xor U17159 (N_17159,N_16340,N_16413);
or U17160 (N_17160,N_16214,N_16213);
and U17161 (N_17161,N_16777,N_16846);
or U17162 (N_17162,N_16875,N_16333);
nand U17163 (N_17163,N_16932,N_16424);
and U17164 (N_17164,N_16212,N_16144);
nand U17165 (N_17165,N_16738,N_16104);
nand U17166 (N_17166,N_16071,N_16887);
nor U17167 (N_17167,N_16290,N_16826);
nand U17168 (N_17168,N_16370,N_16553);
or U17169 (N_17169,N_16012,N_16618);
nor U17170 (N_17170,N_16871,N_16188);
or U17171 (N_17171,N_16287,N_16701);
nor U17172 (N_17172,N_16706,N_16161);
nor U17173 (N_17173,N_16984,N_16934);
nand U17174 (N_17174,N_16399,N_16114);
xnor U17175 (N_17175,N_16793,N_16444);
nor U17176 (N_17176,N_16798,N_16849);
nor U17177 (N_17177,N_16549,N_16274);
or U17178 (N_17178,N_16933,N_16059);
nor U17179 (N_17179,N_16877,N_16100);
xnor U17180 (N_17180,N_16434,N_16337);
nor U17181 (N_17181,N_16425,N_16373);
nand U17182 (N_17182,N_16653,N_16124);
nor U17183 (N_17183,N_16661,N_16821);
nand U17184 (N_17184,N_16072,N_16956);
or U17185 (N_17185,N_16489,N_16464);
or U17186 (N_17186,N_16486,N_16266);
nor U17187 (N_17187,N_16173,N_16565);
nor U17188 (N_17188,N_16750,N_16781);
and U17189 (N_17189,N_16374,N_16523);
or U17190 (N_17190,N_16693,N_16328);
xor U17191 (N_17191,N_16280,N_16401);
nand U17192 (N_17192,N_16234,N_16189);
or U17193 (N_17193,N_16005,N_16536);
xnor U17194 (N_17194,N_16003,N_16551);
or U17195 (N_17195,N_16236,N_16945);
nor U17196 (N_17196,N_16286,N_16986);
nand U17197 (N_17197,N_16316,N_16885);
nand U17198 (N_17198,N_16102,N_16783);
nor U17199 (N_17199,N_16662,N_16588);
or U17200 (N_17200,N_16532,N_16408);
or U17201 (N_17201,N_16911,N_16886);
and U17202 (N_17202,N_16893,N_16749);
nor U17203 (N_17203,N_16673,N_16799);
nand U17204 (N_17204,N_16050,N_16915);
xor U17205 (N_17205,N_16001,N_16779);
nor U17206 (N_17206,N_16162,N_16367);
or U17207 (N_17207,N_16201,N_16612);
or U17208 (N_17208,N_16904,N_16222);
and U17209 (N_17209,N_16756,N_16397);
or U17210 (N_17210,N_16303,N_16013);
or U17211 (N_17211,N_16708,N_16685);
xnor U17212 (N_17212,N_16646,N_16049);
nand U17213 (N_17213,N_16052,N_16082);
and U17214 (N_17214,N_16825,N_16547);
nor U17215 (N_17215,N_16625,N_16836);
nand U17216 (N_17216,N_16582,N_16310);
or U17217 (N_17217,N_16149,N_16240);
or U17218 (N_17218,N_16027,N_16567);
or U17219 (N_17219,N_16483,N_16107);
nand U17220 (N_17220,N_16468,N_16745);
nand U17221 (N_17221,N_16226,N_16635);
or U17222 (N_17222,N_16436,N_16014);
or U17223 (N_17223,N_16513,N_16309);
and U17224 (N_17224,N_16225,N_16651);
xor U17225 (N_17225,N_16259,N_16336);
and U17226 (N_17226,N_16327,N_16047);
or U17227 (N_17227,N_16019,N_16944);
xnor U17228 (N_17228,N_16563,N_16637);
xnor U17229 (N_17229,N_16633,N_16816);
or U17230 (N_17230,N_16800,N_16441);
xnor U17231 (N_17231,N_16331,N_16143);
xnor U17232 (N_17232,N_16811,N_16219);
nor U17233 (N_17233,N_16163,N_16152);
nor U17234 (N_17234,N_16873,N_16381);
or U17235 (N_17235,N_16492,N_16200);
nor U17236 (N_17236,N_16272,N_16768);
nand U17237 (N_17237,N_16641,N_16081);
nor U17238 (N_17238,N_16947,N_16634);
xor U17239 (N_17239,N_16414,N_16539);
or U17240 (N_17240,N_16389,N_16147);
nand U17241 (N_17241,N_16494,N_16395);
and U17242 (N_17242,N_16782,N_16126);
and U17243 (N_17243,N_16325,N_16076);
or U17244 (N_17244,N_16529,N_16057);
nor U17245 (N_17245,N_16655,N_16368);
nor U17246 (N_17246,N_16356,N_16931);
or U17247 (N_17247,N_16407,N_16925);
nand U17248 (N_17248,N_16674,N_16430);
nand U17249 (N_17249,N_16692,N_16043);
nor U17250 (N_17250,N_16055,N_16544);
nand U17251 (N_17251,N_16682,N_16033);
nor U17252 (N_17252,N_16378,N_16892);
or U17253 (N_17253,N_16657,N_16535);
nor U17254 (N_17254,N_16110,N_16861);
or U17255 (N_17255,N_16334,N_16801);
nand U17256 (N_17256,N_16304,N_16823);
or U17257 (N_17257,N_16894,N_16850);
nand U17258 (N_17258,N_16261,N_16251);
or U17259 (N_17259,N_16074,N_16089);
nor U17260 (N_17260,N_16810,N_16815);
or U17261 (N_17261,N_16868,N_16245);
xnor U17262 (N_17262,N_16929,N_16963);
or U17263 (N_17263,N_16807,N_16160);
nand U17264 (N_17264,N_16386,N_16355);
nand U17265 (N_17265,N_16724,N_16363);
nor U17266 (N_17266,N_16137,N_16186);
or U17267 (N_17267,N_16906,N_16900);
or U17268 (N_17268,N_16204,N_16937);
nand U17269 (N_17269,N_16075,N_16687);
nand U17270 (N_17270,N_16686,N_16876);
nor U17271 (N_17271,N_16775,N_16207);
xnor U17272 (N_17272,N_16950,N_16307);
xor U17273 (N_17273,N_16556,N_16164);
xnor U17274 (N_17274,N_16232,N_16854);
nand U17275 (N_17275,N_16797,N_16831);
xnor U17276 (N_17276,N_16169,N_16298);
or U17277 (N_17277,N_16504,N_16168);
or U17278 (N_17278,N_16273,N_16863);
xor U17279 (N_17279,N_16461,N_16808);
nand U17280 (N_17280,N_16335,N_16129);
nand U17281 (N_17281,N_16842,N_16330);
or U17282 (N_17282,N_16105,N_16319);
or U17283 (N_17283,N_16845,N_16505);
nor U17284 (N_17284,N_16118,N_16910);
and U17285 (N_17285,N_16982,N_16809);
nand U17286 (N_17286,N_16839,N_16941);
or U17287 (N_17287,N_16405,N_16613);
or U17288 (N_17288,N_16540,N_16561);
nand U17289 (N_17289,N_16061,N_16394);
nand U17290 (N_17290,N_16606,N_16713);
and U17291 (N_17291,N_16597,N_16690);
nand U17292 (N_17292,N_16766,N_16141);
or U17293 (N_17293,N_16534,N_16707);
nand U17294 (N_17294,N_16824,N_16837);
nand U17295 (N_17295,N_16216,N_16755);
and U17296 (N_17296,N_16384,N_16940);
nor U17297 (N_17297,N_16423,N_16658);
and U17298 (N_17298,N_16663,N_16297);
nand U17299 (N_17299,N_16077,N_16573);
and U17300 (N_17300,N_16636,N_16046);
nand U17301 (N_17301,N_16697,N_16715);
nand U17302 (N_17302,N_16510,N_16041);
or U17303 (N_17303,N_16039,N_16804);
or U17304 (N_17304,N_16835,N_16589);
xor U17305 (N_17305,N_16030,N_16034);
nand U17306 (N_17306,N_16338,N_16231);
nand U17307 (N_17307,N_16860,N_16006);
and U17308 (N_17308,N_16011,N_16905);
nor U17309 (N_17309,N_16281,N_16949);
nand U17310 (N_17310,N_16233,N_16780);
and U17311 (N_17311,N_16127,N_16215);
xor U17312 (N_17312,N_16897,N_16987);
nor U17313 (N_17313,N_16211,N_16739);
xnor U17314 (N_17314,N_16449,N_16067);
or U17315 (N_17315,N_16477,N_16792);
nor U17316 (N_17316,N_16392,N_16970);
nand U17317 (N_17317,N_16209,N_16734);
nor U17318 (N_17318,N_16537,N_16282);
and U17319 (N_17319,N_16068,N_16623);
nand U17320 (N_17320,N_16499,N_16916);
or U17321 (N_17321,N_16645,N_16418);
nand U17322 (N_17322,N_16454,N_16694);
xor U17323 (N_17323,N_16083,N_16456);
xnor U17324 (N_17324,N_16053,N_16560);
xnor U17325 (N_17325,N_16476,N_16292);
nor U17326 (N_17326,N_16838,N_16989);
and U17327 (N_17327,N_16421,N_16647);
xor U17328 (N_17328,N_16479,N_16239);
or U17329 (N_17329,N_16976,N_16691);
nor U17330 (N_17330,N_16935,N_16717);
nand U17331 (N_17331,N_16889,N_16183);
and U17332 (N_17332,N_16939,N_16244);
and U17333 (N_17333,N_16431,N_16242);
xor U17334 (N_17334,N_16912,N_16789);
and U17335 (N_17335,N_16165,N_16527);
or U17336 (N_17336,N_16315,N_16254);
nand U17337 (N_17337,N_16615,N_16501);
or U17338 (N_17338,N_16796,N_16667);
nand U17339 (N_17339,N_16874,N_16522);
nor U17340 (N_17340,N_16148,N_16879);
xnor U17341 (N_17341,N_16362,N_16979);
or U17342 (N_17342,N_16462,N_16353);
nor U17343 (N_17343,N_16683,N_16525);
nand U17344 (N_17344,N_16308,N_16973);
and U17345 (N_17345,N_16238,N_16620);
xnor U17346 (N_17346,N_16584,N_16095);
nor U17347 (N_17347,N_16520,N_16759);
nand U17348 (N_17348,N_16788,N_16429);
nor U17349 (N_17349,N_16313,N_16442);
and U17350 (N_17350,N_16296,N_16930);
nor U17351 (N_17351,N_16278,N_16007);
nand U17352 (N_17352,N_16602,N_16388);
and U17353 (N_17353,N_16364,N_16480);
nand U17354 (N_17354,N_16988,N_16038);
nor U17355 (N_17355,N_16545,N_16293);
nor U17356 (N_17356,N_16971,N_16881);
or U17357 (N_17357,N_16190,N_16509);
or U17358 (N_17358,N_16250,N_16182);
nor U17359 (N_17359,N_16073,N_16913);
or U17360 (N_17360,N_16748,N_16167);
or U17361 (N_17361,N_16351,N_16172);
xor U17362 (N_17362,N_16440,N_16133);
xnor U17363 (N_17363,N_16996,N_16158);
and U17364 (N_17364,N_16321,N_16576);
nand U17365 (N_17365,N_16437,N_16271);
and U17366 (N_17366,N_16721,N_16341);
xor U17367 (N_17367,N_16382,N_16252);
xnor U17368 (N_17368,N_16318,N_16171);
nor U17369 (N_17369,N_16503,N_16317);
or U17370 (N_17370,N_16668,N_16583);
nand U17371 (N_17371,N_16675,N_16269);
or U17372 (N_17372,N_16607,N_16469);
nand U17373 (N_17373,N_16666,N_16720);
or U17374 (N_17374,N_16872,N_16291);
nand U17375 (N_17375,N_16062,N_16398);
or U17376 (N_17376,N_16106,N_16543);
or U17377 (N_17377,N_16732,N_16644);
and U17378 (N_17378,N_16943,N_16320);
nor U17379 (N_17379,N_16841,N_16289);
nand U17380 (N_17380,N_16111,N_16498);
nand U17381 (N_17381,N_16412,N_16450);
nor U17382 (N_17382,N_16032,N_16323);
and U17383 (N_17383,N_16485,N_16729);
nand U17384 (N_17384,N_16703,N_16175);
or U17385 (N_17385,N_16727,N_16869);
xnor U17386 (N_17386,N_16654,N_16819);
nand U17387 (N_17387,N_16300,N_16115);
nand U17388 (N_17388,N_16249,N_16896);
and U17389 (N_17389,N_16299,N_16284);
or U17390 (N_17390,N_16962,N_16184);
and U17391 (N_17391,N_16010,N_16702);
and U17392 (N_17392,N_16453,N_16020);
and U17393 (N_17393,N_16742,N_16669);
or U17394 (N_17394,N_16598,N_16761);
xor U17395 (N_17395,N_16002,N_16762);
or U17396 (N_17396,N_16751,N_16179);
or U17397 (N_17397,N_16998,N_16870);
xor U17398 (N_17398,N_16153,N_16631);
nor U17399 (N_17399,N_16357,N_16024);
and U17400 (N_17400,N_16264,N_16348);
xor U17401 (N_17401,N_16542,N_16972);
or U17402 (N_17402,N_16740,N_16117);
xor U17403 (N_17403,N_16255,N_16360);
and U17404 (N_17404,N_16332,N_16579);
or U17405 (N_17405,N_16571,N_16737);
nand U17406 (N_17406,N_16735,N_16035);
and U17407 (N_17407,N_16145,N_16680);
nand U17408 (N_17408,N_16000,N_16574);
or U17409 (N_17409,N_16980,N_16037);
nand U17410 (N_17410,N_16416,N_16157);
xnor U17411 (N_17411,N_16097,N_16558);
xor U17412 (N_17412,N_16608,N_16828);
nor U17413 (N_17413,N_16306,N_16502);
and U17414 (N_17414,N_16237,N_16210);
nor U17415 (N_17415,N_16578,N_16396);
nor U17416 (N_17416,N_16426,N_16288);
xnor U17417 (N_17417,N_16923,N_16139);
nand U17418 (N_17418,N_16990,N_16428);
nor U17419 (N_17419,N_16500,N_16156);
and U17420 (N_17420,N_16150,N_16744);
xor U17421 (N_17421,N_16593,N_16922);
and U17422 (N_17422,N_16170,N_16283);
nand U17423 (N_17423,N_16758,N_16722);
nor U17424 (N_17424,N_16196,N_16774);
nor U17425 (N_17425,N_16326,N_16570);
nand U17426 (N_17426,N_16009,N_16552);
and U17427 (N_17427,N_16866,N_16512);
xor U17428 (N_17428,N_16638,N_16855);
and U17429 (N_17429,N_16946,N_16626);
nand U17430 (N_17430,N_16420,N_16665);
xor U17431 (N_17431,N_16642,N_16113);
nand U17432 (N_17432,N_16760,N_16723);
nand U17433 (N_17433,N_16314,N_16349);
or U17434 (N_17434,N_16123,N_16822);
nor U17435 (N_17435,N_16121,N_16220);
or U17436 (N_17436,N_16470,N_16099);
and U17437 (N_17437,N_16166,N_16285);
xor U17438 (N_17438,N_16650,N_16865);
nor U17439 (N_17439,N_16964,N_16078);
or U17440 (N_17440,N_16805,N_16592);
xnor U17441 (N_17441,N_16961,N_16806);
nand U17442 (N_17442,N_16086,N_16142);
or U17443 (N_17443,N_16575,N_16714);
and U17444 (N_17444,N_16648,N_16260);
or U17445 (N_17445,N_16718,N_16927);
nor U17446 (N_17446,N_16585,N_16008);
and U17447 (N_17447,N_16066,N_16409);
nand U17448 (N_17448,N_16365,N_16953);
or U17449 (N_17449,N_16859,N_16975);
or U17450 (N_17450,N_16159,N_16562);
xnor U17451 (N_17451,N_16611,N_16021);
or U17452 (N_17452,N_16526,N_16352);
or U17453 (N_17453,N_16277,N_16438);
or U17454 (N_17454,N_16467,N_16491);
nor U17455 (N_17455,N_16433,N_16515);
nand U17456 (N_17456,N_16305,N_16174);
or U17457 (N_17457,N_16347,N_16919);
or U17458 (N_17458,N_16914,N_16684);
nand U17459 (N_17459,N_16676,N_16629);
nand U17460 (N_17460,N_16176,N_16538);
nor U17461 (N_17461,N_16377,N_16622);
or U17462 (N_17462,N_16403,N_16262);
or U17463 (N_17463,N_16022,N_16954);
and U17464 (N_17464,N_16862,N_16614);
or U17465 (N_17465,N_16709,N_16301);
or U17466 (N_17466,N_16342,N_16345);
nand U17467 (N_17467,N_16218,N_16443);
or U17468 (N_17468,N_16093,N_16599);
xor U17469 (N_17469,N_16899,N_16135);
nand U17470 (N_17470,N_16591,N_16586);
xnor U17471 (N_17471,N_16678,N_16140);
xor U17472 (N_17472,N_16507,N_16108);
xnor U17473 (N_17473,N_16820,N_16361);
xor U17474 (N_17474,N_16736,N_16508);
xnor U17475 (N_17475,N_16814,N_16227);
nand U17476 (N_17476,N_16276,N_16402);
nor U17477 (N_17477,N_16487,N_16818);
and U17478 (N_17478,N_16882,N_16619);
xor U17479 (N_17479,N_16268,N_16999);
or U17480 (N_17480,N_16079,N_16497);
xor U17481 (N_17481,N_16595,N_16458);
nand U17482 (N_17482,N_16070,N_16541);
and U17483 (N_17483,N_16754,N_16985);
or U17484 (N_17484,N_16155,N_16036);
or U17485 (N_17485,N_16400,N_16371);
nand U17486 (N_17486,N_16572,N_16833);
or U17487 (N_17487,N_16154,N_16203);
nor U17488 (N_17488,N_16017,N_16380);
nand U17489 (N_17489,N_16390,N_16960);
nand U17490 (N_17490,N_16728,N_16379);
nand U17491 (N_17491,N_16324,N_16903);
and U17492 (N_17492,N_16834,N_16977);
nor U17493 (N_17493,N_16554,N_16448);
nor U17494 (N_17494,N_16018,N_16235);
or U17495 (N_17495,N_16065,N_16294);
or U17496 (N_17496,N_16198,N_16747);
xnor U17497 (N_17497,N_16840,N_16376);
or U17498 (N_17498,N_16594,N_16938);
nand U17499 (N_17499,N_16969,N_16643);
xor U17500 (N_17500,N_16755,N_16403);
xor U17501 (N_17501,N_16729,N_16289);
nor U17502 (N_17502,N_16265,N_16507);
xnor U17503 (N_17503,N_16296,N_16727);
or U17504 (N_17504,N_16651,N_16121);
and U17505 (N_17505,N_16492,N_16232);
nand U17506 (N_17506,N_16082,N_16302);
xnor U17507 (N_17507,N_16132,N_16265);
or U17508 (N_17508,N_16022,N_16702);
and U17509 (N_17509,N_16943,N_16526);
nand U17510 (N_17510,N_16605,N_16716);
or U17511 (N_17511,N_16015,N_16627);
nand U17512 (N_17512,N_16372,N_16828);
nor U17513 (N_17513,N_16227,N_16695);
nor U17514 (N_17514,N_16146,N_16691);
and U17515 (N_17515,N_16118,N_16214);
nor U17516 (N_17516,N_16557,N_16388);
xor U17517 (N_17517,N_16151,N_16253);
nor U17518 (N_17518,N_16092,N_16313);
or U17519 (N_17519,N_16379,N_16074);
and U17520 (N_17520,N_16920,N_16107);
nor U17521 (N_17521,N_16993,N_16920);
and U17522 (N_17522,N_16560,N_16995);
nand U17523 (N_17523,N_16112,N_16954);
nor U17524 (N_17524,N_16722,N_16408);
xnor U17525 (N_17525,N_16058,N_16231);
and U17526 (N_17526,N_16418,N_16609);
nand U17527 (N_17527,N_16574,N_16504);
nand U17528 (N_17528,N_16651,N_16924);
or U17529 (N_17529,N_16591,N_16226);
nor U17530 (N_17530,N_16174,N_16589);
or U17531 (N_17531,N_16021,N_16891);
nand U17532 (N_17532,N_16507,N_16710);
or U17533 (N_17533,N_16281,N_16035);
and U17534 (N_17534,N_16565,N_16918);
or U17535 (N_17535,N_16588,N_16577);
xor U17536 (N_17536,N_16946,N_16832);
xnor U17537 (N_17537,N_16459,N_16981);
and U17538 (N_17538,N_16387,N_16897);
nand U17539 (N_17539,N_16829,N_16248);
or U17540 (N_17540,N_16412,N_16347);
xor U17541 (N_17541,N_16117,N_16763);
nor U17542 (N_17542,N_16031,N_16527);
and U17543 (N_17543,N_16337,N_16704);
nor U17544 (N_17544,N_16786,N_16184);
and U17545 (N_17545,N_16938,N_16599);
xnor U17546 (N_17546,N_16859,N_16771);
or U17547 (N_17547,N_16487,N_16210);
and U17548 (N_17548,N_16169,N_16522);
nor U17549 (N_17549,N_16804,N_16583);
nor U17550 (N_17550,N_16188,N_16795);
nor U17551 (N_17551,N_16627,N_16114);
xnor U17552 (N_17552,N_16033,N_16714);
nor U17553 (N_17553,N_16199,N_16505);
xor U17554 (N_17554,N_16070,N_16976);
or U17555 (N_17555,N_16894,N_16012);
or U17556 (N_17556,N_16864,N_16956);
xor U17557 (N_17557,N_16347,N_16814);
or U17558 (N_17558,N_16343,N_16629);
nor U17559 (N_17559,N_16902,N_16005);
nor U17560 (N_17560,N_16391,N_16177);
and U17561 (N_17561,N_16615,N_16864);
nor U17562 (N_17562,N_16147,N_16712);
or U17563 (N_17563,N_16432,N_16803);
or U17564 (N_17564,N_16660,N_16072);
and U17565 (N_17565,N_16190,N_16923);
xnor U17566 (N_17566,N_16952,N_16840);
nand U17567 (N_17567,N_16985,N_16329);
nor U17568 (N_17568,N_16351,N_16764);
nand U17569 (N_17569,N_16804,N_16972);
or U17570 (N_17570,N_16680,N_16612);
nor U17571 (N_17571,N_16766,N_16365);
and U17572 (N_17572,N_16721,N_16615);
nand U17573 (N_17573,N_16039,N_16847);
or U17574 (N_17574,N_16920,N_16289);
nand U17575 (N_17575,N_16897,N_16747);
nor U17576 (N_17576,N_16273,N_16515);
or U17577 (N_17577,N_16704,N_16969);
nor U17578 (N_17578,N_16014,N_16491);
xnor U17579 (N_17579,N_16272,N_16403);
xnor U17580 (N_17580,N_16209,N_16531);
nor U17581 (N_17581,N_16046,N_16851);
or U17582 (N_17582,N_16243,N_16292);
xor U17583 (N_17583,N_16896,N_16248);
and U17584 (N_17584,N_16368,N_16034);
xor U17585 (N_17585,N_16912,N_16611);
xnor U17586 (N_17586,N_16289,N_16257);
or U17587 (N_17587,N_16017,N_16855);
xnor U17588 (N_17588,N_16836,N_16700);
nor U17589 (N_17589,N_16786,N_16721);
and U17590 (N_17590,N_16422,N_16434);
nand U17591 (N_17591,N_16347,N_16477);
or U17592 (N_17592,N_16252,N_16870);
nor U17593 (N_17593,N_16440,N_16827);
nor U17594 (N_17594,N_16470,N_16043);
and U17595 (N_17595,N_16608,N_16892);
nor U17596 (N_17596,N_16318,N_16553);
or U17597 (N_17597,N_16351,N_16614);
nand U17598 (N_17598,N_16038,N_16449);
xor U17599 (N_17599,N_16876,N_16650);
nor U17600 (N_17600,N_16656,N_16187);
nor U17601 (N_17601,N_16226,N_16112);
or U17602 (N_17602,N_16927,N_16261);
and U17603 (N_17603,N_16505,N_16859);
xor U17604 (N_17604,N_16669,N_16717);
xor U17605 (N_17605,N_16982,N_16566);
and U17606 (N_17606,N_16400,N_16064);
or U17607 (N_17607,N_16721,N_16491);
and U17608 (N_17608,N_16629,N_16331);
and U17609 (N_17609,N_16267,N_16325);
or U17610 (N_17610,N_16738,N_16733);
nor U17611 (N_17611,N_16082,N_16874);
or U17612 (N_17612,N_16363,N_16189);
nand U17613 (N_17613,N_16071,N_16516);
and U17614 (N_17614,N_16042,N_16382);
nand U17615 (N_17615,N_16658,N_16190);
and U17616 (N_17616,N_16963,N_16241);
nor U17617 (N_17617,N_16507,N_16432);
and U17618 (N_17618,N_16073,N_16826);
nor U17619 (N_17619,N_16303,N_16885);
nand U17620 (N_17620,N_16060,N_16811);
nor U17621 (N_17621,N_16687,N_16231);
nand U17622 (N_17622,N_16263,N_16734);
xor U17623 (N_17623,N_16796,N_16286);
or U17624 (N_17624,N_16843,N_16650);
xnor U17625 (N_17625,N_16812,N_16659);
nand U17626 (N_17626,N_16833,N_16224);
and U17627 (N_17627,N_16374,N_16285);
xnor U17628 (N_17628,N_16797,N_16209);
and U17629 (N_17629,N_16850,N_16692);
xor U17630 (N_17630,N_16707,N_16184);
or U17631 (N_17631,N_16580,N_16711);
and U17632 (N_17632,N_16690,N_16871);
and U17633 (N_17633,N_16408,N_16344);
nand U17634 (N_17634,N_16179,N_16606);
and U17635 (N_17635,N_16714,N_16664);
nand U17636 (N_17636,N_16202,N_16817);
nand U17637 (N_17637,N_16173,N_16792);
nand U17638 (N_17638,N_16556,N_16371);
xor U17639 (N_17639,N_16442,N_16546);
and U17640 (N_17640,N_16324,N_16026);
and U17641 (N_17641,N_16472,N_16527);
or U17642 (N_17642,N_16471,N_16225);
nor U17643 (N_17643,N_16369,N_16528);
nand U17644 (N_17644,N_16631,N_16805);
nor U17645 (N_17645,N_16206,N_16558);
nand U17646 (N_17646,N_16841,N_16810);
xnor U17647 (N_17647,N_16068,N_16671);
nand U17648 (N_17648,N_16076,N_16913);
xor U17649 (N_17649,N_16893,N_16062);
and U17650 (N_17650,N_16066,N_16493);
xor U17651 (N_17651,N_16256,N_16247);
or U17652 (N_17652,N_16859,N_16531);
and U17653 (N_17653,N_16736,N_16195);
nor U17654 (N_17654,N_16054,N_16394);
xnor U17655 (N_17655,N_16503,N_16252);
nand U17656 (N_17656,N_16938,N_16949);
or U17657 (N_17657,N_16954,N_16370);
or U17658 (N_17658,N_16492,N_16224);
nor U17659 (N_17659,N_16174,N_16179);
or U17660 (N_17660,N_16757,N_16628);
nand U17661 (N_17661,N_16020,N_16135);
or U17662 (N_17662,N_16224,N_16457);
or U17663 (N_17663,N_16548,N_16617);
xor U17664 (N_17664,N_16163,N_16382);
xnor U17665 (N_17665,N_16965,N_16453);
xnor U17666 (N_17666,N_16889,N_16911);
and U17667 (N_17667,N_16368,N_16962);
and U17668 (N_17668,N_16070,N_16274);
xnor U17669 (N_17669,N_16886,N_16319);
and U17670 (N_17670,N_16102,N_16909);
or U17671 (N_17671,N_16280,N_16714);
xor U17672 (N_17672,N_16671,N_16285);
nor U17673 (N_17673,N_16192,N_16769);
nand U17674 (N_17674,N_16448,N_16699);
nor U17675 (N_17675,N_16530,N_16336);
xor U17676 (N_17676,N_16033,N_16121);
nor U17677 (N_17677,N_16123,N_16209);
or U17678 (N_17678,N_16444,N_16286);
xnor U17679 (N_17679,N_16467,N_16008);
xnor U17680 (N_17680,N_16675,N_16742);
nand U17681 (N_17681,N_16519,N_16389);
or U17682 (N_17682,N_16661,N_16091);
nand U17683 (N_17683,N_16515,N_16036);
nor U17684 (N_17684,N_16791,N_16283);
and U17685 (N_17685,N_16827,N_16250);
nor U17686 (N_17686,N_16240,N_16978);
xor U17687 (N_17687,N_16346,N_16392);
and U17688 (N_17688,N_16567,N_16999);
or U17689 (N_17689,N_16046,N_16653);
xor U17690 (N_17690,N_16541,N_16301);
and U17691 (N_17691,N_16376,N_16537);
or U17692 (N_17692,N_16995,N_16975);
xor U17693 (N_17693,N_16949,N_16247);
and U17694 (N_17694,N_16353,N_16479);
nand U17695 (N_17695,N_16607,N_16285);
nand U17696 (N_17696,N_16575,N_16741);
and U17697 (N_17697,N_16199,N_16822);
nand U17698 (N_17698,N_16091,N_16447);
xor U17699 (N_17699,N_16425,N_16307);
nor U17700 (N_17700,N_16842,N_16696);
xor U17701 (N_17701,N_16992,N_16774);
nand U17702 (N_17702,N_16309,N_16053);
nor U17703 (N_17703,N_16747,N_16976);
or U17704 (N_17704,N_16894,N_16452);
nor U17705 (N_17705,N_16920,N_16579);
xor U17706 (N_17706,N_16265,N_16583);
xnor U17707 (N_17707,N_16469,N_16914);
xnor U17708 (N_17708,N_16597,N_16561);
and U17709 (N_17709,N_16901,N_16183);
and U17710 (N_17710,N_16460,N_16144);
nand U17711 (N_17711,N_16497,N_16944);
nor U17712 (N_17712,N_16310,N_16132);
xnor U17713 (N_17713,N_16455,N_16954);
or U17714 (N_17714,N_16450,N_16249);
xnor U17715 (N_17715,N_16469,N_16276);
or U17716 (N_17716,N_16884,N_16109);
xnor U17717 (N_17717,N_16342,N_16377);
and U17718 (N_17718,N_16498,N_16593);
nand U17719 (N_17719,N_16364,N_16513);
and U17720 (N_17720,N_16267,N_16059);
nor U17721 (N_17721,N_16554,N_16978);
nand U17722 (N_17722,N_16542,N_16656);
nand U17723 (N_17723,N_16966,N_16682);
or U17724 (N_17724,N_16525,N_16456);
or U17725 (N_17725,N_16681,N_16424);
nand U17726 (N_17726,N_16584,N_16593);
or U17727 (N_17727,N_16611,N_16485);
nor U17728 (N_17728,N_16190,N_16142);
nor U17729 (N_17729,N_16830,N_16030);
and U17730 (N_17730,N_16260,N_16453);
nor U17731 (N_17731,N_16515,N_16678);
and U17732 (N_17732,N_16725,N_16277);
and U17733 (N_17733,N_16809,N_16249);
nand U17734 (N_17734,N_16165,N_16061);
and U17735 (N_17735,N_16111,N_16628);
xnor U17736 (N_17736,N_16453,N_16354);
nand U17737 (N_17737,N_16432,N_16304);
nor U17738 (N_17738,N_16631,N_16039);
xor U17739 (N_17739,N_16760,N_16250);
or U17740 (N_17740,N_16017,N_16249);
and U17741 (N_17741,N_16961,N_16854);
and U17742 (N_17742,N_16851,N_16533);
xor U17743 (N_17743,N_16815,N_16896);
xor U17744 (N_17744,N_16354,N_16865);
nand U17745 (N_17745,N_16423,N_16537);
nor U17746 (N_17746,N_16721,N_16777);
or U17747 (N_17747,N_16416,N_16556);
and U17748 (N_17748,N_16601,N_16059);
nand U17749 (N_17749,N_16288,N_16123);
or U17750 (N_17750,N_16182,N_16639);
xor U17751 (N_17751,N_16915,N_16850);
nor U17752 (N_17752,N_16895,N_16131);
or U17753 (N_17753,N_16538,N_16342);
xor U17754 (N_17754,N_16573,N_16940);
or U17755 (N_17755,N_16847,N_16139);
and U17756 (N_17756,N_16480,N_16689);
xor U17757 (N_17757,N_16241,N_16813);
or U17758 (N_17758,N_16191,N_16726);
xnor U17759 (N_17759,N_16171,N_16455);
nand U17760 (N_17760,N_16161,N_16938);
nand U17761 (N_17761,N_16763,N_16622);
nor U17762 (N_17762,N_16019,N_16801);
xnor U17763 (N_17763,N_16952,N_16669);
nand U17764 (N_17764,N_16070,N_16733);
or U17765 (N_17765,N_16259,N_16237);
xor U17766 (N_17766,N_16370,N_16587);
xor U17767 (N_17767,N_16913,N_16195);
and U17768 (N_17768,N_16214,N_16523);
and U17769 (N_17769,N_16534,N_16504);
and U17770 (N_17770,N_16654,N_16264);
and U17771 (N_17771,N_16581,N_16189);
nand U17772 (N_17772,N_16480,N_16145);
nor U17773 (N_17773,N_16100,N_16738);
and U17774 (N_17774,N_16189,N_16357);
or U17775 (N_17775,N_16339,N_16516);
nand U17776 (N_17776,N_16583,N_16442);
nor U17777 (N_17777,N_16743,N_16089);
xnor U17778 (N_17778,N_16458,N_16764);
nand U17779 (N_17779,N_16663,N_16807);
or U17780 (N_17780,N_16538,N_16335);
or U17781 (N_17781,N_16357,N_16052);
nor U17782 (N_17782,N_16382,N_16968);
xnor U17783 (N_17783,N_16093,N_16890);
or U17784 (N_17784,N_16784,N_16216);
and U17785 (N_17785,N_16937,N_16233);
xor U17786 (N_17786,N_16528,N_16941);
or U17787 (N_17787,N_16861,N_16386);
or U17788 (N_17788,N_16718,N_16252);
nand U17789 (N_17789,N_16924,N_16516);
or U17790 (N_17790,N_16430,N_16502);
or U17791 (N_17791,N_16339,N_16569);
nor U17792 (N_17792,N_16365,N_16812);
nor U17793 (N_17793,N_16688,N_16352);
or U17794 (N_17794,N_16715,N_16301);
nand U17795 (N_17795,N_16432,N_16572);
nor U17796 (N_17796,N_16829,N_16750);
nand U17797 (N_17797,N_16660,N_16388);
or U17798 (N_17798,N_16166,N_16393);
and U17799 (N_17799,N_16155,N_16027);
xnor U17800 (N_17800,N_16667,N_16588);
nor U17801 (N_17801,N_16728,N_16832);
nor U17802 (N_17802,N_16537,N_16608);
nand U17803 (N_17803,N_16688,N_16648);
nand U17804 (N_17804,N_16938,N_16153);
xor U17805 (N_17805,N_16408,N_16426);
and U17806 (N_17806,N_16355,N_16139);
or U17807 (N_17807,N_16297,N_16385);
nor U17808 (N_17808,N_16466,N_16835);
nor U17809 (N_17809,N_16406,N_16779);
and U17810 (N_17810,N_16601,N_16153);
xor U17811 (N_17811,N_16799,N_16242);
or U17812 (N_17812,N_16543,N_16350);
nand U17813 (N_17813,N_16431,N_16209);
and U17814 (N_17814,N_16006,N_16423);
and U17815 (N_17815,N_16239,N_16222);
and U17816 (N_17816,N_16712,N_16742);
xnor U17817 (N_17817,N_16986,N_16098);
xor U17818 (N_17818,N_16526,N_16929);
and U17819 (N_17819,N_16300,N_16964);
and U17820 (N_17820,N_16356,N_16246);
nor U17821 (N_17821,N_16128,N_16922);
nor U17822 (N_17822,N_16479,N_16879);
nand U17823 (N_17823,N_16916,N_16134);
xnor U17824 (N_17824,N_16183,N_16713);
nand U17825 (N_17825,N_16935,N_16157);
xor U17826 (N_17826,N_16569,N_16479);
nor U17827 (N_17827,N_16444,N_16214);
nand U17828 (N_17828,N_16919,N_16664);
nor U17829 (N_17829,N_16985,N_16785);
and U17830 (N_17830,N_16347,N_16115);
nand U17831 (N_17831,N_16532,N_16674);
nor U17832 (N_17832,N_16883,N_16472);
nor U17833 (N_17833,N_16582,N_16097);
nor U17834 (N_17834,N_16262,N_16713);
nand U17835 (N_17835,N_16588,N_16075);
or U17836 (N_17836,N_16275,N_16029);
and U17837 (N_17837,N_16380,N_16983);
and U17838 (N_17838,N_16461,N_16048);
or U17839 (N_17839,N_16129,N_16384);
nand U17840 (N_17840,N_16617,N_16445);
nand U17841 (N_17841,N_16869,N_16359);
nand U17842 (N_17842,N_16445,N_16562);
or U17843 (N_17843,N_16711,N_16902);
xnor U17844 (N_17844,N_16969,N_16085);
nand U17845 (N_17845,N_16340,N_16362);
nand U17846 (N_17846,N_16179,N_16100);
nor U17847 (N_17847,N_16257,N_16809);
nand U17848 (N_17848,N_16787,N_16836);
or U17849 (N_17849,N_16684,N_16035);
nand U17850 (N_17850,N_16376,N_16315);
nand U17851 (N_17851,N_16551,N_16137);
nor U17852 (N_17852,N_16824,N_16560);
nand U17853 (N_17853,N_16163,N_16492);
nor U17854 (N_17854,N_16104,N_16352);
nand U17855 (N_17855,N_16339,N_16923);
nand U17856 (N_17856,N_16074,N_16131);
nor U17857 (N_17857,N_16471,N_16203);
xor U17858 (N_17858,N_16612,N_16299);
nor U17859 (N_17859,N_16467,N_16449);
nand U17860 (N_17860,N_16501,N_16429);
nor U17861 (N_17861,N_16961,N_16048);
nand U17862 (N_17862,N_16832,N_16119);
or U17863 (N_17863,N_16905,N_16690);
xor U17864 (N_17864,N_16172,N_16816);
xor U17865 (N_17865,N_16946,N_16494);
nor U17866 (N_17866,N_16059,N_16752);
nor U17867 (N_17867,N_16395,N_16566);
xnor U17868 (N_17868,N_16256,N_16421);
or U17869 (N_17869,N_16621,N_16650);
nand U17870 (N_17870,N_16048,N_16570);
xnor U17871 (N_17871,N_16554,N_16137);
nor U17872 (N_17872,N_16116,N_16254);
and U17873 (N_17873,N_16493,N_16359);
nor U17874 (N_17874,N_16436,N_16692);
or U17875 (N_17875,N_16020,N_16979);
nor U17876 (N_17876,N_16129,N_16089);
nand U17877 (N_17877,N_16152,N_16681);
xnor U17878 (N_17878,N_16280,N_16190);
xor U17879 (N_17879,N_16740,N_16823);
xor U17880 (N_17880,N_16118,N_16615);
nor U17881 (N_17881,N_16694,N_16678);
or U17882 (N_17882,N_16497,N_16983);
nor U17883 (N_17883,N_16345,N_16244);
and U17884 (N_17884,N_16838,N_16543);
nand U17885 (N_17885,N_16652,N_16986);
or U17886 (N_17886,N_16791,N_16300);
nand U17887 (N_17887,N_16210,N_16940);
nor U17888 (N_17888,N_16359,N_16287);
xor U17889 (N_17889,N_16359,N_16208);
xor U17890 (N_17890,N_16520,N_16772);
or U17891 (N_17891,N_16421,N_16999);
xor U17892 (N_17892,N_16432,N_16742);
xor U17893 (N_17893,N_16491,N_16199);
xnor U17894 (N_17894,N_16668,N_16174);
nor U17895 (N_17895,N_16760,N_16854);
nor U17896 (N_17896,N_16152,N_16474);
xnor U17897 (N_17897,N_16753,N_16479);
and U17898 (N_17898,N_16288,N_16385);
xnor U17899 (N_17899,N_16701,N_16371);
or U17900 (N_17900,N_16367,N_16015);
and U17901 (N_17901,N_16892,N_16235);
or U17902 (N_17902,N_16397,N_16514);
nand U17903 (N_17903,N_16413,N_16300);
nand U17904 (N_17904,N_16258,N_16761);
xor U17905 (N_17905,N_16644,N_16826);
and U17906 (N_17906,N_16695,N_16146);
xnor U17907 (N_17907,N_16124,N_16947);
nand U17908 (N_17908,N_16116,N_16990);
nand U17909 (N_17909,N_16566,N_16292);
nor U17910 (N_17910,N_16377,N_16331);
nor U17911 (N_17911,N_16515,N_16526);
and U17912 (N_17912,N_16121,N_16658);
or U17913 (N_17913,N_16652,N_16772);
or U17914 (N_17914,N_16713,N_16625);
nand U17915 (N_17915,N_16383,N_16930);
and U17916 (N_17916,N_16028,N_16977);
and U17917 (N_17917,N_16466,N_16124);
and U17918 (N_17918,N_16998,N_16099);
xnor U17919 (N_17919,N_16596,N_16733);
or U17920 (N_17920,N_16675,N_16407);
nand U17921 (N_17921,N_16733,N_16681);
xnor U17922 (N_17922,N_16786,N_16432);
xor U17923 (N_17923,N_16878,N_16557);
nand U17924 (N_17924,N_16054,N_16906);
nand U17925 (N_17925,N_16685,N_16581);
xor U17926 (N_17926,N_16335,N_16043);
xor U17927 (N_17927,N_16470,N_16150);
nor U17928 (N_17928,N_16637,N_16340);
nand U17929 (N_17929,N_16513,N_16292);
and U17930 (N_17930,N_16694,N_16257);
and U17931 (N_17931,N_16348,N_16684);
nand U17932 (N_17932,N_16490,N_16019);
xnor U17933 (N_17933,N_16851,N_16124);
nor U17934 (N_17934,N_16198,N_16256);
xnor U17935 (N_17935,N_16681,N_16705);
nor U17936 (N_17936,N_16565,N_16859);
or U17937 (N_17937,N_16471,N_16389);
nor U17938 (N_17938,N_16311,N_16679);
nor U17939 (N_17939,N_16183,N_16426);
nand U17940 (N_17940,N_16190,N_16129);
nand U17941 (N_17941,N_16647,N_16683);
or U17942 (N_17942,N_16192,N_16187);
nor U17943 (N_17943,N_16250,N_16381);
nor U17944 (N_17944,N_16943,N_16006);
xnor U17945 (N_17945,N_16468,N_16156);
or U17946 (N_17946,N_16604,N_16614);
nand U17947 (N_17947,N_16465,N_16672);
xnor U17948 (N_17948,N_16877,N_16929);
xnor U17949 (N_17949,N_16805,N_16789);
nand U17950 (N_17950,N_16599,N_16944);
or U17951 (N_17951,N_16201,N_16475);
and U17952 (N_17952,N_16163,N_16372);
xnor U17953 (N_17953,N_16770,N_16227);
nand U17954 (N_17954,N_16363,N_16351);
and U17955 (N_17955,N_16567,N_16306);
and U17956 (N_17956,N_16677,N_16683);
xnor U17957 (N_17957,N_16405,N_16712);
xnor U17958 (N_17958,N_16821,N_16933);
nand U17959 (N_17959,N_16014,N_16589);
xor U17960 (N_17960,N_16916,N_16683);
or U17961 (N_17961,N_16689,N_16861);
nand U17962 (N_17962,N_16873,N_16669);
nand U17963 (N_17963,N_16705,N_16304);
and U17964 (N_17964,N_16268,N_16939);
and U17965 (N_17965,N_16500,N_16141);
or U17966 (N_17966,N_16552,N_16894);
or U17967 (N_17967,N_16899,N_16864);
xnor U17968 (N_17968,N_16449,N_16483);
nand U17969 (N_17969,N_16772,N_16836);
and U17970 (N_17970,N_16705,N_16445);
nor U17971 (N_17971,N_16492,N_16906);
nor U17972 (N_17972,N_16985,N_16674);
and U17973 (N_17973,N_16598,N_16970);
nand U17974 (N_17974,N_16919,N_16978);
or U17975 (N_17975,N_16033,N_16500);
nor U17976 (N_17976,N_16495,N_16483);
xor U17977 (N_17977,N_16960,N_16494);
and U17978 (N_17978,N_16569,N_16277);
xnor U17979 (N_17979,N_16507,N_16767);
xnor U17980 (N_17980,N_16302,N_16280);
and U17981 (N_17981,N_16306,N_16714);
nand U17982 (N_17982,N_16917,N_16384);
xor U17983 (N_17983,N_16178,N_16839);
and U17984 (N_17984,N_16956,N_16030);
xor U17985 (N_17985,N_16816,N_16585);
or U17986 (N_17986,N_16106,N_16440);
nor U17987 (N_17987,N_16227,N_16791);
xnor U17988 (N_17988,N_16385,N_16275);
or U17989 (N_17989,N_16378,N_16534);
nor U17990 (N_17990,N_16426,N_16001);
nand U17991 (N_17991,N_16988,N_16190);
nor U17992 (N_17992,N_16889,N_16329);
nand U17993 (N_17993,N_16512,N_16266);
nand U17994 (N_17994,N_16001,N_16159);
nand U17995 (N_17995,N_16960,N_16017);
nor U17996 (N_17996,N_16076,N_16442);
or U17997 (N_17997,N_16026,N_16522);
nand U17998 (N_17998,N_16742,N_16777);
or U17999 (N_17999,N_16054,N_16142);
xnor U18000 (N_18000,N_17600,N_17327);
nor U18001 (N_18001,N_17933,N_17695);
and U18002 (N_18002,N_17035,N_17120);
nor U18003 (N_18003,N_17009,N_17438);
xnor U18004 (N_18004,N_17848,N_17267);
or U18005 (N_18005,N_17004,N_17800);
nand U18006 (N_18006,N_17949,N_17156);
nor U18007 (N_18007,N_17172,N_17819);
or U18008 (N_18008,N_17828,N_17412);
and U18009 (N_18009,N_17142,N_17101);
and U18010 (N_18010,N_17333,N_17409);
nor U18011 (N_18011,N_17166,N_17794);
xor U18012 (N_18012,N_17132,N_17261);
or U18013 (N_18013,N_17401,N_17430);
nand U18014 (N_18014,N_17399,N_17840);
and U18015 (N_18015,N_17861,N_17739);
nor U18016 (N_18016,N_17047,N_17332);
and U18017 (N_18017,N_17025,N_17415);
or U18018 (N_18018,N_17114,N_17992);
nand U18019 (N_18019,N_17658,N_17467);
nand U18020 (N_18020,N_17504,N_17281);
or U18021 (N_18021,N_17212,N_17494);
or U18022 (N_18022,N_17429,N_17975);
nor U18023 (N_18023,N_17977,N_17970);
nor U18024 (N_18024,N_17817,N_17884);
nor U18025 (N_18025,N_17956,N_17950);
xor U18026 (N_18026,N_17338,N_17485);
nor U18027 (N_18027,N_17017,N_17051);
and U18028 (N_18028,N_17974,N_17566);
or U18029 (N_18029,N_17735,N_17124);
nand U18030 (N_18030,N_17957,N_17562);
nor U18031 (N_18031,N_17366,N_17516);
xnor U18032 (N_18032,N_17618,N_17894);
xnor U18033 (N_18033,N_17592,N_17610);
nor U18034 (N_18034,N_17876,N_17134);
and U18035 (N_18035,N_17940,N_17639);
nor U18036 (N_18036,N_17147,N_17784);
or U18037 (N_18037,N_17468,N_17622);
nand U18038 (N_18038,N_17460,N_17307);
xnor U18039 (N_18039,N_17763,N_17030);
nand U18040 (N_18040,N_17837,N_17103);
nand U18041 (N_18041,N_17442,N_17295);
nand U18042 (N_18042,N_17753,N_17698);
or U18043 (N_18043,N_17274,N_17221);
xnor U18044 (N_18044,N_17663,N_17509);
nor U18045 (N_18045,N_17318,N_17407);
nand U18046 (N_18046,N_17305,N_17402);
nand U18047 (N_18047,N_17972,N_17928);
and U18048 (N_18048,N_17766,N_17629);
nand U18049 (N_18049,N_17078,N_17759);
or U18050 (N_18050,N_17608,N_17821);
xor U18051 (N_18051,N_17843,N_17079);
xnor U18052 (N_18052,N_17311,N_17667);
or U18053 (N_18053,N_17724,N_17097);
xnor U18054 (N_18054,N_17184,N_17827);
nor U18055 (N_18055,N_17590,N_17532);
nor U18056 (N_18056,N_17614,N_17576);
nand U18057 (N_18057,N_17432,N_17077);
nand U18058 (N_18058,N_17553,N_17322);
nor U18059 (N_18059,N_17162,N_17368);
or U18060 (N_18060,N_17507,N_17313);
nand U18061 (N_18061,N_17359,N_17041);
and U18062 (N_18062,N_17679,N_17067);
nand U18063 (N_18063,N_17436,N_17642);
nand U18064 (N_18064,N_17619,N_17013);
nand U18065 (N_18065,N_17584,N_17207);
or U18066 (N_18066,N_17547,N_17606);
and U18067 (N_18067,N_17541,N_17196);
xnor U18068 (N_18068,N_17841,N_17499);
or U18069 (N_18069,N_17781,N_17703);
nor U18070 (N_18070,N_17382,N_17945);
xor U18071 (N_18071,N_17088,N_17683);
and U18072 (N_18072,N_17830,N_17666);
nand U18073 (N_18073,N_17561,N_17746);
and U18074 (N_18074,N_17091,N_17820);
xor U18075 (N_18075,N_17376,N_17981);
or U18076 (N_18076,N_17498,N_17080);
nor U18077 (N_18077,N_17104,N_17413);
or U18078 (N_18078,N_17326,N_17993);
or U18079 (N_18079,N_17016,N_17689);
nand U18080 (N_18080,N_17024,N_17059);
nand U18081 (N_18081,N_17119,N_17756);
nor U18082 (N_18082,N_17270,N_17866);
or U18083 (N_18083,N_17908,N_17681);
xnor U18084 (N_18084,N_17772,N_17268);
nand U18085 (N_18085,N_17692,N_17996);
or U18086 (N_18086,N_17582,N_17265);
or U18087 (N_18087,N_17143,N_17810);
nor U18088 (N_18088,N_17994,N_17350);
or U18089 (N_18089,N_17767,N_17877);
or U18090 (N_18090,N_17251,N_17653);
and U18091 (N_18091,N_17701,N_17337);
nor U18092 (N_18092,N_17447,N_17502);
nor U18093 (N_18093,N_17090,N_17854);
nand U18094 (N_18094,N_17719,N_17976);
and U18095 (N_18095,N_17937,N_17813);
nand U18096 (N_18096,N_17577,N_17804);
nor U18097 (N_18097,N_17082,N_17217);
xnor U18098 (N_18098,N_17700,N_17792);
xnor U18099 (N_18099,N_17360,N_17954);
nand U18100 (N_18100,N_17573,N_17410);
nand U18101 (N_18101,N_17304,N_17095);
xor U18102 (N_18102,N_17284,N_17336);
xnor U18103 (N_18103,N_17129,N_17697);
xnor U18104 (N_18104,N_17631,N_17801);
or U18105 (N_18105,N_17849,N_17930);
nand U18106 (N_18106,N_17776,N_17023);
nand U18107 (N_18107,N_17086,N_17064);
nand U18108 (N_18108,N_17560,N_17643);
xor U18109 (N_18109,N_17010,N_17380);
nand U18110 (N_18110,N_17721,N_17216);
xnor U18111 (N_18111,N_17913,N_17448);
and U18112 (N_18112,N_17527,N_17427);
xor U18113 (N_18113,N_17807,N_17397);
nand U18114 (N_18114,N_17883,N_17728);
or U18115 (N_18115,N_17795,N_17676);
nor U18116 (N_18116,N_17100,N_17179);
and U18117 (N_18117,N_17144,N_17652);
and U18118 (N_18118,N_17938,N_17300);
nand U18119 (N_18119,N_17967,N_17364);
xnor U18120 (N_18120,N_17372,N_17717);
or U18121 (N_18121,N_17116,N_17985);
nor U18122 (N_18122,N_17015,N_17654);
xor U18123 (N_18123,N_17001,N_17968);
xor U18124 (N_18124,N_17459,N_17493);
nand U18125 (N_18125,N_17780,N_17672);
xnor U18126 (N_18126,N_17369,N_17315);
nand U18127 (N_18127,N_17660,N_17882);
or U18128 (N_18128,N_17685,N_17012);
nand U18129 (N_18129,N_17534,N_17236);
or U18130 (N_18130,N_17121,N_17388);
nand U18131 (N_18131,N_17462,N_17314);
nand U18132 (N_18132,N_17531,N_17483);
xor U18133 (N_18133,N_17105,N_17519);
xor U18134 (N_18134,N_17452,N_17157);
or U18135 (N_18135,N_17093,N_17109);
or U18136 (N_18136,N_17137,N_17244);
xor U18137 (N_18137,N_17623,N_17550);
and U18138 (N_18138,N_17063,N_17812);
xnor U18139 (N_18139,N_17647,N_17390);
or U18140 (N_18140,N_17141,N_17674);
nor U18141 (N_18141,N_17011,N_17000);
xor U18142 (N_18142,N_17889,N_17711);
xnor U18143 (N_18143,N_17897,N_17056);
nand U18144 (N_18144,N_17554,N_17238);
xnor U18145 (N_18145,N_17040,N_17328);
or U18146 (N_18146,N_17158,N_17099);
and U18147 (N_18147,N_17193,N_17515);
and U18148 (N_18148,N_17720,N_17526);
and U18149 (N_18149,N_17638,N_17572);
nor U18150 (N_18150,N_17456,N_17732);
and U18151 (N_18151,N_17909,N_17754);
and U18152 (N_18152,N_17260,N_17190);
and U18153 (N_18153,N_17615,N_17433);
nor U18154 (N_18154,N_17049,N_17223);
and U18155 (N_18155,N_17856,N_17558);
xnor U18156 (N_18156,N_17123,N_17487);
nor U18157 (N_18157,N_17523,N_17072);
xor U18158 (N_18158,N_17242,N_17929);
xor U18159 (N_18159,N_17014,N_17964);
nor U18160 (N_18160,N_17862,N_17916);
xnor U18161 (N_18161,N_17375,N_17549);
and U18162 (N_18162,N_17518,N_17678);
or U18163 (N_18163,N_17521,N_17525);
and U18164 (N_18164,N_17716,N_17832);
or U18165 (N_18165,N_17246,N_17387);
nor U18166 (N_18166,N_17505,N_17989);
nor U18167 (N_18167,N_17220,N_17736);
or U18168 (N_18168,N_17321,N_17478);
and U18169 (N_18169,N_17750,N_17389);
or U18170 (N_18170,N_17280,N_17888);
xnor U18171 (N_18171,N_17464,N_17965);
nor U18172 (N_18172,N_17655,N_17818);
or U18173 (N_18173,N_17871,N_17227);
nor U18174 (N_18174,N_17323,N_17651);
and U18175 (N_18175,N_17215,N_17511);
or U18176 (N_18176,N_17228,N_17210);
nand U18177 (N_18177,N_17755,N_17370);
xnor U18178 (N_18178,N_17159,N_17297);
nor U18179 (N_18179,N_17878,N_17741);
and U18180 (N_18180,N_17363,N_17037);
nor U18181 (N_18181,N_17367,N_17749);
and U18182 (N_18182,N_17708,N_17334);
nor U18183 (N_18183,N_17508,N_17834);
xnor U18184 (N_18184,N_17490,N_17596);
and U18185 (N_18185,N_17520,N_17362);
or U18186 (N_18186,N_17868,N_17312);
nand U18187 (N_18187,N_17186,N_17071);
and U18188 (N_18188,N_17115,N_17988);
nor U18189 (N_18189,N_17192,N_17910);
nand U18190 (N_18190,N_17924,N_17714);
nor U18191 (N_18191,N_17497,N_17718);
xor U18192 (N_18192,N_17420,N_17206);
nor U18193 (N_18193,N_17627,N_17935);
and U18194 (N_18194,N_17029,N_17942);
nand U18195 (N_18195,N_17453,N_17987);
nor U18196 (N_18196,N_17943,N_17038);
xor U18197 (N_18197,N_17565,N_17068);
and U18198 (N_18198,N_17850,N_17133);
xnor U18199 (N_18199,N_17302,N_17982);
and U18200 (N_18200,N_17269,N_17570);
nor U18201 (N_18201,N_17771,N_17624);
nor U18202 (N_18202,N_17744,N_17403);
xnor U18203 (N_18203,N_17858,N_17995);
and U18204 (N_18204,N_17536,N_17458);
nand U18205 (N_18205,N_17555,N_17803);
or U18206 (N_18206,N_17748,N_17997);
nand U18207 (N_18207,N_17126,N_17440);
xor U18208 (N_18208,N_17715,N_17282);
nand U18209 (N_18209,N_17348,N_17028);
nor U18210 (N_18210,N_17428,N_17587);
nor U18211 (N_18211,N_17860,N_17904);
and U18212 (N_18212,N_17501,N_17761);
and U18213 (N_18213,N_17791,N_17354);
or U18214 (N_18214,N_17229,N_17919);
and U18215 (N_18215,N_17500,N_17696);
nand U18216 (N_18216,N_17768,N_17425);
xnor U18217 (N_18217,N_17661,N_17208);
and U18218 (N_18218,N_17557,N_17903);
nor U18219 (N_18219,N_17686,N_17241);
and U18220 (N_18220,N_17342,N_17296);
and U18221 (N_18221,N_17613,N_17019);
or U18222 (N_18222,N_17778,N_17451);
or U18223 (N_18223,N_17125,N_17445);
xor U18224 (N_18224,N_17659,N_17486);
xnor U18225 (N_18225,N_17214,N_17912);
nor U18226 (N_18226,N_17953,N_17495);
and U18227 (N_18227,N_17605,N_17583);
nor U18228 (N_18228,N_17959,N_17796);
xnor U18229 (N_18229,N_17852,N_17202);
or U18230 (N_18230,N_17036,N_17797);
xnor U18231 (N_18231,N_17470,N_17838);
and U18232 (N_18232,N_17675,N_17809);
nand U18233 (N_18233,N_17303,N_17626);
and U18234 (N_18234,N_17863,N_17008);
nor U18235 (N_18235,N_17847,N_17551);
or U18236 (N_18236,N_17839,N_17075);
or U18237 (N_18237,N_17253,N_17379);
or U18238 (N_18238,N_17747,N_17385);
and U18239 (N_18239,N_17998,N_17690);
nand U18240 (N_18240,N_17680,N_17574);
nor U18241 (N_18241,N_17875,N_17374);
nand U18242 (N_18242,N_17266,N_17783);
xor U18243 (N_18243,N_17371,N_17290);
nor U18244 (N_18244,N_17154,N_17278);
nor U18245 (N_18245,N_17102,N_17469);
and U18246 (N_18246,N_17224,N_17579);
nand U18247 (N_18247,N_17693,N_17391);
and U18248 (N_18248,N_17727,N_17506);
xnor U18249 (N_18249,N_17277,N_17931);
nand U18250 (N_18250,N_17219,N_17880);
nor U18251 (N_18251,N_17779,N_17404);
nand U18252 (N_18252,N_17074,N_17252);
and U18253 (N_18253,N_17081,N_17053);
and U18254 (N_18254,N_17538,N_17317);
and U18255 (N_18255,N_17769,N_17249);
or U18256 (N_18256,N_17108,N_17405);
nand U18257 (N_18257,N_17729,N_17073);
or U18258 (N_18258,N_17823,N_17089);
nand U18259 (N_18259,N_17168,N_17640);
and U18260 (N_18260,N_17320,N_17491);
xnor U18261 (N_18261,N_17301,N_17775);
or U18262 (N_18262,N_17272,N_17512);
xnor U18263 (N_18263,N_17752,N_17816);
and U18264 (N_18264,N_17543,N_17130);
and U18265 (N_18265,N_17087,N_17588);
xor U18266 (N_18266,N_17222,N_17170);
and U18267 (N_18267,N_17477,N_17611);
nor U18268 (N_18268,N_17226,N_17594);
nor U18269 (N_18269,N_17955,N_17039);
nand U18270 (N_18270,N_17032,N_17991);
or U18271 (N_18271,N_17734,N_17177);
nand U18272 (N_18272,N_17829,N_17593);
and U18273 (N_18273,N_17707,N_17757);
xnor U18274 (N_18274,N_17595,N_17806);
xnor U18275 (N_18275,N_17127,N_17331);
nor U18276 (N_18276,N_17033,N_17330);
nor U18277 (N_18277,N_17925,N_17983);
nor U18278 (N_18278,N_17620,N_17762);
xnor U18279 (N_18279,N_17774,N_17589);
and U18280 (N_18280,N_17662,N_17522);
nor U18281 (N_18281,N_17926,N_17233);
xor U18282 (N_18282,N_17439,N_17349);
nand U18283 (N_18283,N_17112,N_17174);
nor U18284 (N_18284,N_17240,N_17182);
nand U18285 (N_18285,N_17031,N_17417);
nand U18286 (N_18286,N_17770,N_17824);
and U18287 (N_18287,N_17636,N_17891);
nor U18288 (N_18288,N_17406,N_17211);
and U18289 (N_18289,N_17645,N_17185);
nand U18290 (N_18290,N_17450,N_17670);
nor U18291 (N_18291,N_17237,N_17632);
or U18292 (N_18292,N_17649,N_17422);
and U18293 (N_18293,N_17153,N_17218);
and U18294 (N_18294,N_17225,N_17646);
and U18295 (N_18295,N_17948,N_17963);
nor U18296 (N_18296,N_17630,N_17437);
and U18297 (N_18297,N_17879,N_17058);
or U18298 (N_18298,N_17107,N_17567);
nand U18299 (N_18299,N_17984,N_17283);
nor U18300 (N_18300,N_17291,N_17263);
or U18301 (N_18301,N_17482,N_17355);
xnor U18302 (N_18302,N_17932,N_17230);
and U18303 (N_18303,N_17351,N_17421);
or U18304 (N_18304,N_17634,N_17285);
xor U18305 (N_18305,N_17786,N_17597);
and U18306 (N_18306,N_17293,N_17138);
and U18307 (N_18307,N_17052,N_17245);
xnor U18308 (N_18308,N_17050,N_17545);
xnor U18309 (N_18309,N_17329,N_17833);
nand U18310 (N_18310,N_17069,N_17286);
nand U18311 (N_18311,N_17393,N_17886);
nor U18312 (N_18312,N_17018,N_17969);
or U18313 (N_18313,N_17900,N_17258);
and U18314 (N_18314,N_17461,N_17197);
nor U18315 (N_18315,N_17822,N_17484);
nor U18316 (N_18316,N_17978,N_17952);
xor U18317 (N_18317,N_17083,N_17664);
and U18318 (N_18318,N_17423,N_17394);
and U18319 (N_18319,N_17310,N_17887);
and U18320 (N_18320,N_17481,N_17668);
or U18321 (N_18321,N_17378,N_17869);
or U18322 (N_18322,N_17292,N_17044);
or U18323 (N_18323,N_17092,N_17764);
and U18324 (N_18324,N_17872,N_17431);
or U18325 (N_18325,N_17239,N_17287);
nand U18326 (N_18326,N_17529,N_17234);
nor U18327 (N_18327,N_17256,N_17203);
nor U18328 (N_18328,N_17669,N_17835);
or U18329 (N_18329,N_17540,N_17340);
nand U18330 (N_18330,N_17022,N_17671);
nand U18331 (N_18331,N_17279,N_17826);
xor U18332 (N_18332,N_17128,N_17475);
nor U18333 (N_18333,N_17414,N_17339);
or U18334 (N_18334,N_17927,N_17146);
nor U18335 (N_18335,N_17788,N_17556);
nor U18336 (N_18336,N_17195,N_17730);
nand U18337 (N_18337,N_17737,N_17773);
nor U18338 (N_18338,N_17055,N_17895);
and U18339 (N_18339,N_17152,N_17607);
nand U18340 (N_18340,N_17936,N_17194);
nor U18341 (N_18341,N_17601,N_17548);
nor U18342 (N_18342,N_17738,N_17454);
and U18343 (N_18343,N_17633,N_17325);
nand U18344 (N_18344,N_17528,N_17061);
nand U18345 (N_18345,N_17434,N_17905);
xor U18346 (N_18346,N_17140,N_17160);
and U18347 (N_18347,N_17424,N_17787);
xor U18348 (N_18348,N_17045,N_17145);
nor U18349 (N_18349,N_17187,N_17085);
and U18350 (N_18350,N_17065,N_17966);
nor U18351 (N_18351,N_17851,N_17255);
or U18352 (N_18352,N_17918,N_17745);
xor U18353 (N_18353,N_17885,N_17042);
xor U18354 (N_18354,N_17906,N_17113);
or U18355 (N_18355,N_17694,N_17917);
nor U18356 (N_18356,N_17066,N_17899);
and U18357 (N_18357,N_17377,N_17864);
nand U18358 (N_18358,N_17625,N_17947);
nor U18359 (N_18359,N_17740,N_17874);
or U18360 (N_18360,N_17914,N_17199);
and U18361 (N_18361,N_17463,N_17398);
nor U18362 (N_18362,N_17578,N_17163);
or U18363 (N_18363,N_17855,N_17898);
or U18364 (N_18364,N_17479,N_17542);
or U18365 (N_18365,N_17136,N_17513);
nand U18366 (N_18366,N_17713,N_17922);
nand U18367 (N_18367,N_17201,N_17441);
xor U18368 (N_18368,N_17859,N_17357);
or U18369 (N_18369,N_17496,N_17361);
xnor U18370 (N_18370,N_17189,N_17564);
nor U18371 (N_18371,N_17324,N_17273);
or U18372 (N_18372,N_17699,N_17979);
or U18373 (N_18373,N_17005,N_17726);
and U18374 (N_18374,N_17621,N_17276);
nor U18375 (N_18375,N_17076,N_17760);
nand U18376 (N_18376,N_17920,N_17533);
nand U18377 (N_18377,N_17148,N_17785);
xnor U18378 (N_18378,N_17492,N_17559);
nor U18379 (N_18379,N_17373,N_17175);
xor U18380 (N_18380,N_17581,N_17893);
or U18381 (N_18381,N_17723,N_17489);
xor U18382 (N_18382,N_17790,N_17111);
nand U18383 (N_18383,N_17356,N_17198);
and U18384 (N_18384,N_17161,N_17782);
and U18385 (N_18385,N_17873,N_17743);
xor U18386 (N_18386,N_17510,N_17173);
nand U18387 (N_18387,N_17384,N_17443);
and U18388 (N_18388,N_17907,N_17980);
nor U18389 (N_18389,N_17971,N_17169);
and U18390 (N_18390,N_17825,N_17209);
nand U18391 (N_18391,N_17188,N_17973);
or U18392 (N_18392,N_17309,N_17003);
and U18393 (N_18393,N_17259,N_17831);
or U18394 (N_18394,N_17688,N_17705);
and U18395 (N_18395,N_17815,N_17167);
nor U18396 (N_18396,N_17751,N_17007);
and U18397 (N_18397,N_17006,N_17923);
xor U18398 (N_18398,N_17961,N_17789);
and U18399 (N_18399,N_17999,N_17704);
xnor U18400 (N_18400,N_17777,N_17271);
or U18401 (N_18401,N_17183,N_17386);
and U18402 (N_18402,N_17990,N_17345);
xnor U18403 (N_18403,N_17395,N_17706);
nand U18404 (N_18404,N_17546,N_17524);
and U18405 (N_18405,N_17106,N_17381);
nand U18406 (N_18406,N_17396,N_17165);
xor U18407 (N_18407,N_17656,N_17644);
or U18408 (N_18408,N_17383,N_17235);
nand U18409 (N_18409,N_17358,N_17084);
nand U18410 (N_18410,N_17846,N_17289);
and U18411 (N_18411,N_17027,N_17335);
or U18412 (N_18412,N_17231,N_17098);
xnor U18413 (N_18413,N_17094,N_17944);
nand U18414 (N_18414,N_17444,N_17476);
and U18415 (N_18415,N_17117,N_17808);
and U18416 (N_18416,N_17725,N_17793);
and U18417 (N_18417,N_17473,N_17842);
nand U18418 (N_18418,N_17575,N_17308);
nor U18419 (N_18419,N_17118,N_17805);
xnor U18420 (N_18420,N_17205,N_17845);
or U18421 (N_18421,N_17319,N_17811);
nor U18422 (N_18422,N_17934,N_17365);
nor U18423 (N_18423,N_17503,N_17537);
nand U18424 (N_18424,N_17722,N_17939);
nor U18425 (N_18425,N_17488,N_17002);
nand U18426 (N_18426,N_17465,N_17609);
nand U18427 (N_18427,N_17568,N_17164);
nand U18428 (N_18428,N_17299,N_17802);
xor U18429 (N_18429,N_17288,N_17602);
nand U18430 (N_18430,N_17257,N_17844);
nor U18431 (N_18431,N_17054,N_17446);
and U18432 (N_18432,N_17673,N_17539);
and U18433 (N_18433,N_17637,N_17650);
nand U18434 (N_18434,N_17480,N_17921);
or U18435 (N_18435,N_17691,N_17435);
nand U18436 (N_18436,N_17867,N_17986);
xor U18437 (N_18437,N_17426,N_17598);
nor U18438 (N_18438,N_17298,N_17641);
or U18439 (N_18439,N_17911,N_17896);
xnor U18440 (N_18440,N_17799,N_17677);
and U18441 (N_18441,N_17648,N_17070);
and U18442 (N_18442,N_17684,N_17254);
nor U18443 (N_18443,N_17026,N_17457);
or U18444 (N_18444,N_17343,N_17294);
and U18445 (N_18445,N_17742,N_17392);
or U18446 (N_18446,N_17710,N_17472);
xor U18447 (N_18447,N_17306,N_17344);
and U18448 (N_18448,N_17657,N_17131);
nor U18449 (N_18449,N_17046,N_17419);
or U18450 (N_18450,N_17798,N_17057);
xnor U18451 (N_18451,N_17043,N_17155);
or U18452 (N_18452,N_17599,N_17275);
nor U18453 (N_18453,N_17603,N_17178);
or U18454 (N_18454,N_17617,N_17712);
xor U18455 (N_18455,N_17408,N_17892);
or U18456 (N_18456,N_17530,N_17247);
nand U18457 (N_18457,N_17151,N_17471);
or U18458 (N_18458,N_17316,N_17865);
and U18459 (N_18459,N_17213,N_17733);
and U18460 (N_18460,N_17552,N_17449);
and U18461 (N_18461,N_17571,N_17902);
nor U18462 (N_18462,N_17890,N_17264);
nand U18463 (N_18463,N_17466,N_17758);
or U18464 (N_18464,N_17586,N_17122);
and U18465 (N_18465,N_17181,N_17418);
or U18466 (N_18466,N_17110,N_17200);
nor U18467 (N_18467,N_17702,N_17191);
nand U18468 (N_18468,N_17901,N_17021);
xnor U18469 (N_18469,N_17232,N_17946);
nor U18470 (N_18470,N_17062,N_17616);
or U18471 (N_18471,N_17150,N_17020);
nor U18472 (N_18472,N_17535,N_17604);
nand U18473 (N_18473,N_17060,N_17347);
and U18474 (N_18474,N_17591,N_17765);
xnor U18475 (N_18475,N_17682,N_17951);
or U18476 (N_18476,N_17243,N_17857);
nor U18477 (N_18477,N_17352,N_17411);
nand U18478 (N_18478,N_17585,N_17474);
xnor U18479 (N_18479,N_17870,N_17400);
and U18480 (N_18480,N_17353,N_17204);
or U18481 (N_18481,N_17048,N_17171);
nand U18482 (N_18482,N_17709,N_17853);
nand U18483 (N_18483,N_17248,N_17731);
nand U18484 (N_18484,N_17180,N_17135);
and U18485 (N_18485,N_17962,N_17569);
and U18486 (N_18486,N_17250,N_17941);
and U18487 (N_18487,N_17544,N_17960);
nor U18488 (N_18488,N_17612,N_17580);
and U18489 (N_18489,N_17687,N_17149);
nor U18490 (N_18490,N_17958,N_17514);
nand U18491 (N_18491,N_17915,N_17176);
or U18492 (N_18492,N_17836,N_17416);
nor U18493 (N_18493,N_17034,N_17262);
nor U18494 (N_18494,N_17881,N_17814);
nor U18495 (N_18495,N_17665,N_17455);
or U18496 (N_18496,N_17628,N_17341);
and U18497 (N_18497,N_17635,N_17096);
nor U18498 (N_18498,N_17139,N_17346);
or U18499 (N_18499,N_17517,N_17563);
nand U18500 (N_18500,N_17941,N_17711);
and U18501 (N_18501,N_17673,N_17970);
xnor U18502 (N_18502,N_17484,N_17456);
nor U18503 (N_18503,N_17395,N_17177);
and U18504 (N_18504,N_17463,N_17437);
or U18505 (N_18505,N_17870,N_17360);
xnor U18506 (N_18506,N_17008,N_17733);
xnor U18507 (N_18507,N_17820,N_17702);
and U18508 (N_18508,N_17028,N_17288);
or U18509 (N_18509,N_17143,N_17837);
xor U18510 (N_18510,N_17138,N_17314);
nor U18511 (N_18511,N_17875,N_17862);
nand U18512 (N_18512,N_17198,N_17765);
nor U18513 (N_18513,N_17993,N_17268);
and U18514 (N_18514,N_17091,N_17769);
xor U18515 (N_18515,N_17330,N_17154);
and U18516 (N_18516,N_17405,N_17627);
nor U18517 (N_18517,N_17189,N_17197);
xor U18518 (N_18518,N_17069,N_17806);
nand U18519 (N_18519,N_17790,N_17931);
and U18520 (N_18520,N_17903,N_17575);
or U18521 (N_18521,N_17720,N_17448);
and U18522 (N_18522,N_17059,N_17163);
xor U18523 (N_18523,N_17546,N_17830);
xor U18524 (N_18524,N_17899,N_17468);
or U18525 (N_18525,N_17204,N_17279);
xnor U18526 (N_18526,N_17483,N_17903);
and U18527 (N_18527,N_17745,N_17315);
and U18528 (N_18528,N_17060,N_17506);
nand U18529 (N_18529,N_17995,N_17912);
or U18530 (N_18530,N_17512,N_17941);
nand U18531 (N_18531,N_17079,N_17270);
xnor U18532 (N_18532,N_17792,N_17565);
nor U18533 (N_18533,N_17165,N_17868);
nand U18534 (N_18534,N_17184,N_17495);
nor U18535 (N_18535,N_17117,N_17258);
and U18536 (N_18536,N_17222,N_17907);
xor U18537 (N_18537,N_17406,N_17540);
or U18538 (N_18538,N_17211,N_17083);
and U18539 (N_18539,N_17668,N_17379);
nor U18540 (N_18540,N_17218,N_17373);
nand U18541 (N_18541,N_17467,N_17065);
or U18542 (N_18542,N_17698,N_17813);
xor U18543 (N_18543,N_17126,N_17974);
xor U18544 (N_18544,N_17045,N_17808);
nor U18545 (N_18545,N_17838,N_17905);
or U18546 (N_18546,N_17455,N_17269);
xor U18547 (N_18547,N_17156,N_17924);
xnor U18548 (N_18548,N_17836,N_17932);
and U18549 (N_18549,N_17206,N_17061);
nand U18550 (N_18550,N_17960,N_17952);
nor U18551 (N_18551,N_17083,N_17165);
or U18552 (N_18552,N_17010,N_17762);
nand U18553 (N_18553,N_17546,N_17538);
nand U18554 (N_18554,N_17005,N_17215);
and U18555 (N_18555,N_17277,N_17167);
and U18556 (N_18556,N_17812,N_17059);
nor U18557 (N_18557,N_17560,N_17042);
nand U18558 (N_18558,N_17225,N_17170);
xnor U18559 (N_18559,N_17997,N_17851);
nor U18560 (N_18560,N_17000,N_17628);
xor U18561 (N_18561,N_17606,N_17996);
and U18562 (N_18562,N_17678,N_17451);
and U18563 (N_18563,N_17082,N_17344);
nor U18564 (N_18564,N_17358,N_17519);
and U18565 (N_18565,N_17546,N_17061);
or U18566 (N_18566,N_17747,N_17759);
nand U18567 (N_18567,N_17878,N_17131);
nand U18568 (N_18568,N_17759,N_17911);
or U18569 (N_18569,N_17360,N_17208);
or U18570 (N_18570,N_17384,N_17062);
and U18571 (N_18571,N_17826,N_17116);
xnor U18572 (N_18572,N_17692,N_17536);
or U18573 (N_18573,N_17059,N_17518);
or U18574 (N_18574,N_17226,N_17360);
and U18575 (N_18575,N_17156,N_17456);
and U18576 (N_18576,N_17090,N_17332);
xor U18577 (N_18577,N_17072,N_17475);
nor U18578 (N_18578,N_17368,N_17412);
xnor U18579 (N_18579,N_17660,N_17055);
nand U18580 (N_18580,N_17602,N_17030);
xor U18581 (N_18581,N_17399,N_17147);
and U18582 (N_18582,N_17442,N_17162);
nand U18583 (N_18583,N_17155,N_17552);
nand U18584 (N_18584,N_17181,N_17690);
xor U18585 (N_18585,N_17390,N_17712);
nor U18586 (N_18586,N_17530,N_17954);
xnor U18587 (N_18587,N_17369,N_17912);
nor U18588 (N_18588,N_17295,N_17116);
nand U18589 (N_18589,N_17094,N_17166);
nand U18590 (N_18590,N_17872,N_17899);
or U18591 (N_18591,N_17684,N_17155);
and U18592 (N_18592,N_17335,N_17861);
nor U18593 (N_18593,N_17768,N_17046);
nor U18594 (N_18594,N_17839,N_17520);
or U18595 (N_18595,N_17592,N_17875);
and U18596 (N_18596,N_17700,N_17120);
or U18597 (N_18597,N_17196,N_17508);
or U18598 (N_18598,N_17772,N_17514);
nor U18599 (N_18599,N_17581,N_17843);
nand U18600 (N_18600,N_17888,N_17951);
and U18601 (N_18601,N_17680,N_17666);
nor U18602 (N_18602,N_17296,N_17963);
nand U18603 (N_18603,N_17402,N_17431);
nand U18604 (N_18604,N_17149,N_17111);
nand U18605 (N_18605,N_17213,N_17658);
nor U18606 (N_18606,N_17334,N_17943);
and U18607 (N_18607,N_17650,N_17175);
or U18608 (N_18608,N_17157,N_17638);
xnor U18609 (N_18609,N_17921,N_17577);
nand U18610 (N_18610,N_17189,N_17357);
nor U18611 (N_18611,N_17465,N_17453);
and U18612 (N_18612,N_17244,N_17834);
and U18613 (N_18613,N_17416,N_17560);
and U18614 (N_18614,N_17629,N_17806);
nor U18615 (N_18615,N_17661,N_17718);
xnor U18616 (N_18616,N_17290,N_17400);
xor U18617 (N_18617,N_17773,N_17973);
nor U18618 (N_18618,N_17065,N_17116);
nand U18619 (N_18619,N_17593,N_17181);
xor U18620 (N_18620,N_17827,N_17642);
and U18621 (N_18621,N_17073,N_17140);
xor U18622 (N_18622,N_17145,N_17826);
or U18623 (N_18623,N_17294,N_17479);
and U18624 (N_18624,N_17326,N_17772);
xor U18625 (N_18625,N_17833,N_17597);
xnor U18626 (N_18626,N_17949,N_17463);
nand U18627 (N_18627,N_17798,N_17437);
or U18628 (N_18628,N_17653,N_17853);
nor U18629 (N_18629,N_17102,N_17784);
nand U18630 (N_18630,N_17134,N_17468);
nor U18631 (N_18631,N_17604,N_17150);
and U18632 (N_18632,N_17753,N_17979);
nor U18633 (N_18633,N_17708,N_17584);
xor U18634 (N_18634,N_17604,N_17115);
nand U18635 (N_18635,N_17564,N_17743);
nor U18636 (N_18636,N_17657,N_17752);
nand U18637 (N_18637,N_17608,N_17525);
xor U18638 (N_18638,N_17249,N_17386);
nor U18639 (N_18639,N_17677,N_17950);
or U18640 (N_18640,N_17933,N_17158);
xor U18641 (N_18641,N_17812,N_17912);
xor U18642 (N_18642,N_17035,N_17208);
or U18643 (N_18643,N_17088,N_17680);
xor U18644 (N_18644,N_17895,N_17177);
or U18645 (N_18645,N_17651,N_17997);
nor U18646 (N_18646,N_17398,N_17915);
nand U18647 (N_18647,N_17833,N_17359);
nand U18648 (N_18648,N_17969,N_17663);
nor U18649 (N_18649,N_17524,N_17550);
and U18650 (N_18650,N_17775,N_17928);
nand U18651 (N_18651,N_17940,N_17514);
nor U18652 (N_18652,N_17884,N_17355);
and U18653 (N_18653,N_17559,N_17936);
xor U18654 (N_18654,N_17028,N_17684);
and U18655 (N_18655,N_17733,N_17829);
nand U18656 (N_18656,N_17270,N_17633);
nand U18657 (N_18657,N_17399,N_17876);
and U18658 (N_18658,N_17466,N_17708);
xor U18659 (N_18659,N_17462,N_17641);
nand U18660 (N_18660,N_17629,N_17080);
and U18661 (N_18661,N_17475,N_17510);
or U18662 (N_18662,N_17178,N_17077);
or U18663 (N_18663,N_17061,N_17436);
nor U18664 (N_18664,N_17875,N_17810);
nand U18665 (N_18665,N_17726,N_17414);
nand U18666 (N_18666,N_17919,N_17270);
and U18667 (N_18667,N_17584,N_17332);
or U18668 (N_18668,N_17428,N_17128);
nand U18669 (N_18669,N_17758,N_17840);
and U18670 (N_18670,N_17488,N_17354);
nor U18671 (N_18671,N_17366,N_17974);
and U18672 (N_18672,N_17523,N_17587);
nand U18673 (N_18673,N_17242,N_17941);
or U18674 (N_18674,N_17906,N_17944);
xnor U18675 (N_18675,N_17634,N_17780);
and U18676 (N_18676,N_17962,N_17119);
nand U18677 (N_18677,N_17686,N_17274);
xnor U18678 (N_18678,N_17889,N_17592);
or U18679 (N_18679,N_17666,N_17920);
or U18680 (N_18680,N_17124,N_17871);
and U18681 (N_18681,N_17512,N_17306);
or U18682 (N_18682,N_17103,N_17684);
nand U18683 (N_18683,N_17911,N_17318);
or U18684 (N_18684,N_17986,N_17929);
or U18685 (N_18685,N_17174,N_17784);
nand U18686 (N_18686,N_17255,N_17836);
nor U18687 (N_18687,N_17139,N_17028);
nor U18688 (N_18688,N_17249,N_17154);
nor U18689 (N_18689,N_17036,N_17925);
or U18690 (N_18690,N_17885,N_17456);
xor U18691 (N_18691,N_17806,N_17734);
nand U18692 (N_18692,N_17791,N_17710);
nor U18693 (N_18693,N_17102,N_17866);
nand U18694 (N_18694,N_17102,N_17672);
xor U18695 (N_18695,N_17467,N_17727);
or U18696 (N_18696,N_17562,N_17031);
or U18697 (N_18697,N_17804,N_17216);
and U18698 (N_18698,N_17947,N_17042);
xor U18699 (N_18699,N_17279,N_17683);
nand U18700 (N_18700,N_17916,N_17172);
nor U18701 (N_18701,N_17697,N_17641);
nor U18702 (N_18702,N_17081,N_17639);
or U18703 (N_18703,N_17097,N_17924);
or U18704 (N_18704,N_17944,N_17620);
nor U18705 (N_18705,N_17049,N_17230);
nor U18706 (N_18706,N_17825,N_17268);
xnor U18707 (N_18707,N_17888,N_17250);
nor U18708 (N_18708,N_17248,N_17018);
nand U18709 (N_18709,N_17013,N_17256);
and U18710 (N_18710,N_17128,N_17057);
nor U18711 (N_18711,N_17460,N_17131);
or U18712 (N_18712,N_17868,N_17599);
and U18713 (N_18713,N_17606,N_17804);
and U18714 (N_18714,N_17288,N_17120);
and U18715 (N_18715,N_17814,N_17264);
or U18716 (N_18716,N_17714,N_17781);
nor U18717 (N_18717,N_17094,N_17970);
or U18718 (N_18718,N_17881,N_17433);
and U18719 (N_18719,N_17519,N_17840);
and U18720 (N_18720,N_17367,N_17615);
nand U18721 (N_18721,N_17222,N_17557);
nand U18722 (N_18722,N_17575,N_17410);
nand U18723 (N_18723,N_17839,N_17191);
nand U18724 (N_18724,N_17100,N_17585);
and U18725 (N_18725,N_17406,N_17458);
nor U18726 (N_18726,N_17137,N_17047);
and U18727 (N_18727,N_17889,N_17300);
or U18728 (N_18728,N_17225,N_17812);
nor U18729 (N_18729,N_17344,N_17839);
xor U18730 (N_18730,N_17257,N_17086);
xor U18731 (N_18731,N_17698,N_17138);
nor U18732 (N_18732,N_17399,N_17347);
nand U18733 (N_18733,N_17607,N_17471);
nand U18734 (N_18734,N_17021,N_17298);
and U18735 (N_18735,N_17388,N_17878);
xnor U18736 (N_18736,N_17957,N_17420);
nand U18737 (N_18737,N_17385,N_17572);
nor U18738 (N_18738,N_17969,N_17447);
nor U18739 (N_18739,N_17210,N_17233);
xor U18740 (N_18740,N_17244,N_17418);
xor U18741 (N_18741,N_17047,N_17556);
nand U18742 (N_18742,N_17213,N_17999);
nor U18743 (N_18743,N_17112,N_17460);
xnor U18744 (N_18744,N_17506,N_17752);
and U18745 (N_18745,N_17759,N_17908);
nand U18746 (N_18746,N_17684,N_17287);
nor U18747 (N_18747,N_17006,N_17841);
xor U18748 (N_18748,N_17640,N_17172);
and U18749 (N_18749,N_17590,N_17956);
and U18750 (N_18750,N_17466,N_17287);
nor U18751 (N_18751,N_17791,N_17578);
xnor U18752 (N_18752,N_17435,N_17962);
nor U18753 (N_18753,N_17511,N_17437);
xor U18754 (N_18754,N_17668,N_17222);
xor U18755 (N_18755,N_17142,N_17417);
or U18756 (N_18756,N_17307,N_17871);
nor U18757 (N_18757,N_17138,N_17440);
and U18758 (N_18758,N_17222,N_17237);
or U18759 (N_18759,N_17118,N_17434);
or U18760 (N_18760,N_17521,N_17346);
xor U18761 (N_18761,N_17906,N_17885);
and U18762 (N_18762,N_17542,N_17060);
nor U18763 (N_18763,N_17754,N_17077);
or U18764 (N_18764,N_17162,N_17748);
or U18765 (N_18765,N_17358,N_17399);
xnor U18766 (N_18766,N_17128,N_17865);
nand U18767 (N_18767,N_17692,N_17273);
xor U18768 (N_18768,N_17701,N_17293);
and U18769 (N_18769,N_17414,N_17694);
nand U18770 (N_18770,N_17526,N_17927);
or U18771 (N_18771,N_17024,N_17904);
and U18772 (N_18772,N_17638,N_17859);
nand U18773 (N_18773,N_17416,N_17523);
nor U18774 (N_18774,N_17395,N_17035);
nor U18775 (N_18775,N_17510,N_17063);
xnor U18776 (N_18776,N_17540,N_17804);
and U18777 (N_18777,N_17101,N_17999);
or U18778 (N_18778,N_17979,N_17065);
nand U18779 (N_18779,N_17008,N_17040);
or U18780 (N_18780,N_17488,N_17352);
nand U18781 (N_18781,N_17742,N_17328);
or U18782 (N_18782,N_17172,N_17001);
xnor U18783 (N_18783,N_17360,N_17383);
nand U18784 (N_18784,N_17787,N_17598);
and U18785 (N_18785,N_17706,N_17103);
xnor U18786 (N_18786,N_17213,N_17489);
or U18787 (N_18787,N_17890,N_17517);
or U18788 (N_18788,N_17754,N_17662);
and U18789 (N_18789,N_17477,N_17129);
nor U18790 (N_18790,N_17263,N_17295);
and U18791 (N_18791,N_17015,N_17383);
xnor U18792 (N_18792,N_17161,N_17239);
nand U18793 (N_18793,N_17205,N_17668);
xnor U18794 (N_18794,N_17510,N_17397);
and U18795 (N_18795,N_17496,N_17516);
xnor U18796 (N_18796,N_17257,N_17902);
xor U18797 (N_18797,N_17096,N_17906);
xor U18798 (N_18798,N_17639,N_17057);
nand U18799 (N_18799,N_17406,N_17675);
xor U18800 (N_18800,N_17896,N_17602);
and U18801 (N_18801,N_17728,N_17990);
and U18802 (N_18802,N_17915,N_17200);
or U18803 (N_18803,N_17363,N_17822);
nor U18804 (N_18804,N_17063,N_17178);
or U18805 (N_18805,N_17232,N_17217);
and U18806 (N_18806,N_17106,N_17593);
or U18807 (N_18807,N_17727,N_17047);
nor U18808 (N_18808,N_17342,N_17397);
nor U18809 (N_18809,N_17053,N_17162);
nor U18810 (N_18810,N_17101,N_17475);
xnor U18811 (N_18811,N_17981,N_17580);
nor U18812 (N_18812,N_17461,N_17164);
xnor U18813 (N_18813,N_17818,N_17825);
and U18814 (N_18814,N_17594,N_17884);
xnor U18815 (N_18815,N_17681,N_17407);
and U18816 (N_18816,N_17760,N_17995);
nand U18817 (N_18817,N_17453,N_17098);
xor U18818 (N_18818,N_17681,N_17634);
and U18819 (N_18819,N_17293,N_17023);
or U18820 (N_18820,N_17137,N_17282);
xnor U18821 (N_18821,N_17499,N_17491);
nor U18822 (N_18822,N_17920,N_17537);
or U18823 (N_18823,N_17227,N_17397);
and U18824 (N_18824,N_17788,N_17644);
xnor U18825 (N_18825,N_17072,N_17163);
nor U18826 (N_18826,N_17146,N_17839);
or U18827 (N_18827,N_17532,N_17917);
nand U18828 (N_18828,N_17346,N_17167);
nand U18829 (N_18829,N_17685,N_17390);
or U18830 (N_18830,N_17305,N_17072);
xnor U18831 (N_18831,N_17274,N_17599);
nor U18832 (N_18832,N_17275,N_17058);
nor U18833 (N_18833,N_17199,N_17273);
xor U18834 (N_18834,N_17389,N_17956);
nor U18835 (N_18835,N_17546,N_17708);
nor U18836 (N_18836,N_17664,N_17903);
or U18837 (N_18837,N_17474,N_17296);
or U18838 (N_18838,N_17887,N_17132);
nor U18839 (N_18839,N_17300,N_17835);
or U18840 (N_18840,N_17222,N_17873);
xnor U18841 (N_18841,N_17590,N_17868);
nand U18842 (N_18842,N_17740,N_17803);
and U18843 (N_18843,N_17730,N_17213);
or U18844 (N_18844,N_17410,N_17283);
nand U18845 (N_18845,N_17664,N_17502);
nor U18846 (N_18846,N_17244,N_17440);
nor U18847 (N_18847,N_17563,N_17147);
nand U18848 (N_18848,N_17102,N_17295);
nand U18849 (N_18849,N_17059,N_17789);
xnor U18850 (N_18850,N_17599,N_17744);
xnor U18851 (N_18851,N_17871,N_17827);
nand U18852 (N_18852,N_17737,N_17950);
nor U18853 (N_18853,N_17990,N_17406);
and U18854 (N_18854,N_17698,N_17490);
and U18855 (N_18855,N_17818,N_17701);
or U18856 (N_18856,N_17317,N_17828);
xor U18857 (N_18857,N_17405,N_17388);
nor U18858 (N_18858,N_17421,N_17242);
or U18859 (N_18859,N_17852,N_17006);
and U18860 (N_18860,N_17493,N_17655);
or U18861 (N_18861,N_17183,N_17647);
nand U18862 (N_18862,N_17950,N_17488);
or U18863 (N_18863,N_17409,N_17396);
xnor U18864 (N_18864,N_17717,N_17492);
or U18865 (N_18865,N_17815,N_17298);
xor U18866 (N_18866,N_17762,N_17887);
or U18867 (N_18867,N_17777,N_17194);
nand U18868 (N_18868,N_17588,N_17012);
nand U18869 (N_18869,N_17760,N_17838);
xnor U18870 (N_18870,N_17150,N_17849);
or U18871 (N_18871,N_17155,N_17763);
nor U18872 (N_18872,N_17853,N_17701);
nor U18873 (N_18873,N_17543,N_17470);
or U18874 (N_18874,N_17533,N_17428);
nor U18875 (N_18875,N_17547,N_17505);
xnor U18876 (N_18876,N_17560,N_17387);
nand U18877 (N_18877,N_17649,N_17180);
nand U18878 (N_18878,N_17514,N_17086);
and U18879 (N_18879,N_17029,N_17554);
or U18880 (N_18880,N_17343,N_17354);
nor U18881 (N_18881,N_17334,N_17998);
xnor U18882 (N_18882,N_17467,N_17853);
xor U18883 (N_18883,N_17566,N_17238);
nand U18884 (N_18884,N_17944,N_17078);
nor U18885 (N_18885,N_17366,N_17219);
or U18886 (N_18886,N_17631,N_17102);
or U18887 (N_18887,N_17729,N_17118);
nand U18888 (N_18888,N_17255,N_17661);
xor U18889 (N_18889,N_17107,N_17390);
nor U18890 (N_18890,N_17257,N_17206);
nand U18891 (N_18891,N_17909,N_17945);
and U18892 (N_18892,N_17391,N_17110);
xor U18893 (N_18893,N_17275,N_17611);
nor U18894 (N_18894,N_17699,N_17383);
and U18895 (N_18895,N_17854,N_17965);
xor U18896 (N_18896,N_17478,N_17342);
nand U18897 (N_18897,N_17042,N_17049);
nand U18898 (N_18898,N_17223,N_17105);
or U18899 (N_18899,N_17184,N_17760);
xnor U18900 (N_18900,N_17340,N_17700);
nand U18901 (N_18901,N_17283,N_17736);
nand U18902 (N_18902,N_17641,N_17307);
xor U18903 (N_18903,N_17918,N_17763);
xor U18904 (N_18904,N_17605,N_17446);
and U18905 (N_18905,N_17293,N_17670);
nand U18906 (N_18906,N_17617,N_17919);
nor U18907 (N_18907,N_17810,N_17873);
nand U18908 (N_18908,N_17544,N_17614);
or U18909 (N_18909,N_17008,N_17912);
nand U18910 (N_18910,N_17265,N_17146);
and U18911 (N_18911,N_17412,N_17005);
nand U18912 (N_18912,N_17706,N_17492);
xor U18913 (N_18913,N_17220,N_17101);
or U18914 (N_18914,N_17935,N_17760);
xor U18915 (N_18915,N_17768,N_17369);
nor U18916 (N_18916,N_17251,N_17993);
xnor U18917 (N_18917,N_17247,N_17180);
nand U18918 (N_18918,N_17521,N_17190);
xor U18919 (N_18919,N_17893,N_17393);
or U18920 (N_18920,N_17356,N_17931);
nor U18921 (N_18921,N_17119,N_17689);
nor U18922 (N_18922,N_17570,N_17934);
or U18923 (N_18923,N_17879,N_17665);
and U18924 (N_18924,N_17969,N_17227);
xor U18925 (N_18925,N_17948,N_17605);
nand U18926 (N_18926,N_17350,N_17248);
and U18927 (N_18927,N_17523,N_17273);
or U18928 (N_18928,N_17664,N_17926);
nor U18929 (N_18929,N_17267,N_17699);
nand U18930 (N_18930,N_17934,N_17614);
and U18931 (N_18931,N_17194,N_17009);
nand U18932 (N_18932,N_17725,N_17396);
or U18933 (N_18933,N_17603,N_17848);
nor U18934 (N_18934,N_17283,N_17803);
or U18935 (N_18935,N_17849,N_17480);
nand U18936 (N_18936,N_17473,N_17989);
or U18937 (N_18937,N_17003,N_17946);
nor U18938 (N_18938,N_17143,N_17291);
or U18939 (N_18939,N_17618,N_17354);
or U18940 (N_18940,N_17525,N_17921);
or U18941 (N_18941,N_17859,N_17279);
nand U18942 (N_18942,N_17324,N_17381);
nand U18943 (N_18943,N_17132,N_17021);
and U18944 (N_18944,N_17246,N_17464);
or U18945 (N_18945,N_17460,N_17952);
nor U18946 (N_18946,N_17890,N_17446);
and U18947 (N_18947,N_17354,N_17505);
or U18948 (N_18948,N_17953,N_17273);
nand U18949 (N_18949,N_17466,N_17906);
nor U18950 (N_18950,N_17211,N_17892);
nand U18951 (N_18951,N_17571,N_17618);
nor U18952 (N_18952,N_17448,N_17897);
nand U18953 (N_18953,N_17783,N_17865);
or U18954 (N_18954,N_17324,N_17898);
nor U18955 (N_18955,N_17562,N_17033);
or U18956 (N_18956,N_17670,N_17116);
and U18957 (N_18957,N_17808,N_17963);
or U18958 (N_18958,N_17327,N_17935);
nor U18959 (N_18959,N_17176,N_17532);
nor U18960 (N_18960,N_17796,N_17399);
xnor U18961 (N_18961,N_17933,N_17694);
and U18962 (N_18962,N_17539,N_17985);
and U18963 (N_18963,N_17441,N_17280);
and U18964 (N_18964,N_17980,N_17172);
or U18965 (N_18965,N_17158,N_17142);
and U18966 (N_18966,N_17376,N_17459);
nand U18967 (N_18967,N_17299,N_17776);
or U18968 (N_18968,N_17912,N_17103);
and U18969 (N_18969,N_17926,N_17296);
nor U18970 (N_18970,N_17012,N_17178);
nand U18971 (N_18971,N_17559,N_17999);
xor U18972 (N_18972,N_17832,N_17681);
and U18973 (N_18973,N_17694,N_17615);
nand U18974 (N_18974,N_17186,N_17155);
nor U18975 (N_18975,N_17905,N_17160);
and U18976 (N_18976,N_17439,N_17496);
or U18977 (N_18977,N_17011,N_17059);
or U18978 (N_18978,N_17642,N_17623);
xnor U18979 (N_18979,N_17467,N_17197);
or U18980 (N_18980,N_17472,N_17059);
nand U18981 (N_18981,N_17009,N_17510);
and U18982 (N_18982,N_17513,N_17608);
nor U18983 (N_18983,N_17123,N_17075);
and U18984 (N_18984,N_17097,N_17259);
nand U18985 (N_18985,N_17583,N_17716);
or U18986 (N_18986,N_17675,N_17462);
nor U18987 (N_18987,N_17460,N_17613);
or U18988 (N_18988,N_17125,N_17009);
nand U18989 (N_18989,N_17073,N_17443);
and U18990 (N_18990,N_17241,N_17944);
xnor U18991 (N_18991,N_17358,N_17649);
and U18992 (N_18992,N_17060,N_17670);
xor U18993 (N_18993,N_17224,N_17942);
and U18994 (N_18994,N_17427,N_17524);
and U18995 (N_18995,N_17530,N_17608);
xnor U18996 (N_18996,N_17964,N_17155);
xor U18997 (N_18997,N_17780,N_17737);
or U18998 (N_18998,N_17207,N_17615);
nand U18999 (N_18999,N_17568,N_17341);
and U19000 (N_19000,N_18399,N_18672);
and U19001 (N_19001,N_18220,N_18119);
and U19002 (N_19002,N_18273,N_18713);
or U19003 (N_19003,N_18025,N_18870);
and U19004 (N_19004,N_18855,N_18152);
nor U19005 (N_19005,N_18262,N_18379);
or U19006 (N_19006,N_18709,N_18380);
xnor U19007 (N_19007,N_18969,N_18931);
and U19008 (N_19008,N_18035,N_18808);
nand U19009 (N_19009,N_18533,N_18727);
and U19010 (N_19010,N_18984,N_18677);
and U19011 (N_19011,N_18584,N_18178);
or U19012 (N_19012,N_18690,N_18587);
xor U19013 (N_19013,N_18743,N_18937);
or U19014 (N_19014,N_18358,N_18736);
nand U19015 (N_19015,N_18260,N_18346);
or U19016 (N_19016,N_18771,N_18852);
and U19017 (N_19017,N_18548,N_18619);
nor U19018 (N_19018,N_18943,N_18641);
and U19019 (N_19019,N_18885,N_18590);
nor U19020 (N_19020,N_18310,N_18518);
and U19021 (N_19021,N_18552,N_18502);
and U19022 (N_19022,N_18401,N_18429);
nor U19023 (N_19023,N_18348,N_18209);
or U19024 (N_19024,N_18109,N_18261);
nand U19025 (N_19025,N_18469,N_18047);
nor U19026 (N_19026,N_18092,N_18388);
nand U19027 (N_19027,N_18583,N_18848);
nand U19028 (N_19028,N_18711,N_18577);
xnor U19029 (N_19029,N_18072,N_18654);
nand U19030 (N_19030,N_18068,N_18942);
or U19031 (N_19031,N_18345,N_18434);
nand U19032 (N_19032,N_18881,N_18982);
and U19033 (N_19033,N_18222,N_18461);
or U19034 (N_19034,N_18567,N_18500);
xor U19035 (N_19035,N_18366,N_18298);
and U19036 (N_19036,N_18053,N_18341);
nand U19037 (N_19037,N_18048,N_18285);
and U19038 (N_19038,N_18739,N_18030);
xnor U19039 (N_19039,N_18156,N_18286);
xnor U19040 (N_19040,N_18194,N_18008);
nor U19041 (N_19041,N_18452,N_18701);
nand U19042 (N_19042,N_18451,N_18819);
and U19043 (N_19043,N_18698,N_18055);
or U19044 (N_19044,N_18205,N_18287);
xnor U19045 (N_19045,N_18783,N_18763);
nand U19046 (N_19046,N_18077,N_18418);
nor U19047 (N_19047,N_18467,N_18618);
and U19048 (N_19048,N_18844,N_18371);
nand U19049 (N_19049,N_18865,N_18566);
or U19050 (N_19050,N_18520,N_18915);
xor U19051 (N_19051,N_18210,N_18160);
nor U19052 (N_19052,N_18253,N_18793);
nor U19053 (N_19053,N_18407,N_18213);
and U19054 (N_19054,N_18738,N_18464);
nand U19055 (N_19055,N_18192,N_18324);
nand U19056 (N_19056,N_18560,N_18661);
or U19057 (N_19057,N_18015,N_18350);
nand U19058 (N_19058,N_18305,N_18666);
nor U19059 (N_19059,N_18498,N_18197);
nor U19060 (N_19060,N_18516,N_18607);
nand U19061 (N_19061,N_18921,N_18689);
and U19062 (N_19062,N_18961,N_18717);
or U19063 (N_19063,N_18532,N_18440);
and U19064 (N_19064,N_18471,N_18934);
and U19065 (N_19065,N_18188,N_18483);
or U19066 (N_19066,N_18172,N_18397);
nand U19067 (N_19067,N_18400,N_18255);
nor U19068 (N_19068,N_18311,N_18017);
nor U19069 (N_19069,N_18417,N_18144);
or U19070 (N_19070,N_18993,N_18662);
or U19071 (N_19071,N_18167,N_18880);
or U19072 (N_19072,N_18105,N_18540);
nand U19073 (N_19073,N_18510,N_18300);
and U19074 (N_19074,N_18912,N_18707);
nand U19075 (N_19075,N_18482,N_18496);
and U19076 (N_19076,N_18408,N_18538);
nor U19077 (N_19077,N_18193,N_18712);
nand U19078 (N_19078,N_18140,N_18060);
or U19079 (N_19079,N_18450,N_18497);
xor U19080 (N_19080,N_18876,N_18335);
and U19081 (N_19081,N_18040,N_18064);
or U19082 (N_19082,N_18445,N_18734);
nand U19083 (N_19083,N_18322,N_18492);
and U19084 (N_19084,N_18612,N_18766);
nand U19085 (N_19085,N_18892,N_18276);
xor U19086 (N_19086,N_18901,N_18363);
nor U19087 (N_19087,N_18703,N_18569);
nor U19088 (N_19088,N_18603,N_18221);
nand U19089 (N_19089,N_18330,N_18280);
nand U19090 (N_19090,N_18155,N_18997);
nand U19091 (N_19091,N_18826,N_18905);
or U19092 (N_19092,N_18853,N_18941);
or U19093 (N_19093,N_18874,N_18256);
xnor U19094 (N_19094,N_18393,N_18326);
or U19095 (N_19095,N_18395,N_18232);
xor U19096 (N_19096,N_18320,N_18179);
and U19097 (N_19097,N_18091,N_18438);
or U19098 (N_19098,N_18882,N_18229);
nor U19099 (N_19099,N_18034,N_18671);
or U19100 (N_19100,N_18457,N_18086);
and U19101 (N_19101,N_18331,N_18906);
xor U19102 (N_19102,N_18107,N_18480);
xnor U19103 (N_19103,N_18237,N_18202);
nor U19104 (N_19104,N_18974,N_18499);
or U19105 (N_19105,N_18267,N_18066);
nor U19106 (N_19106,N_18663,N_18889);
nor U19107 (N_19107,N_18744,N_18359);
or U19108 (N_19108,N_18725,N_18090);
and U19109 (N_19109,N_18585,N_18329);
nor U19110 (N_19110,N_18686,N_18057);
nor U19111 (N_19111,N_18594,N_18138);
or U19112 (N_19112,N_18275,N_18697);
nand U19113 (N_19113,N_18849,N_18375);
xor U19114 (N_19114,N_18867,N_18589);
nor U19115 (N_19115,N_18554,N_18123);
or U19116 (N_19116,N_18888,N_18815);
nor U19117 (N_19117,N_18441,N_18682);
and U19118 (N_19118,N_18460,N_18095);
and U19119 (N_19119,N_18730,N_18531);
or U19120 (N_19120,N_18546,N_18317);
nand U19121 (N_19121,N_18952,N_18318);
nor U19122 (N_19122,N_18243,N_18128);
and U19123 (N_19123,N_18611,N_18837);
xnor U19124 (N_19124,N_18693,N_18512);
and U19125 (N_19125,N_18652,N_18802);
xor U19126 (N_19126,N_18597,N_18547);
or U19127 (N_19127,N_18147,N_18288);
nor U19128 (N_19128,N_18543,N_18410);
nor U19129 (N_19129,N_18005,N_18196);
nand U19130 (N_19130,N_18575,N_18283);
nand U19131 (N_19131,N_18474,N_18559);
nor U19132 (N_19132,N_18838,N_18878);
or U19133 (N_19133,N_18685,N_18307);
or U19134 (N_19134,N_18922,N_18604);
nand U19135 (N_19135,N_18344,N_18930);
or U19136 (N_19136,N_18297,N_18565);
nor U19137 (N_19137,N_18443,N_18812);
nand U19138 (N_19138,N_18303,N_18938);
nor U19139 (N_19139,N_18032,N_18814);
xnor U19140 (N_19140,N_18054,N_18978);
nor U19141 (N_19141,N_18225,N_18792);
xor U19142 (N_19142,N_18405,N_18023);
nand U19143 (N_19143,N_18551,N_18487);
and U19144 (N_19144,N_18511,N_18349);
nor U19145 (N_19145,N_18608,N_18831);
xnor U19146 (N_19146,N_18673,N_18351);
or U19147 (N_19147,N_18101,N_18760);
and U19148 (N_19148,N_18126,N_18100);
xnor U19149 (N_19149,N_18694,N_18636);
and U19150 (N_19150,N_18239,N_18732);
xnor U19151 (N_19151,N_18757,N_18268);
nand U19152 (N_19152,N_18056,N_18266);
or U19153 (N_19153,N_18678,N_18890);
xor U19154 (N_19154,N_18336,N_18505);
and U19155 (N_19155,N_18011,N_18564);
nand U19156 (N_19156,N_18644,N_18807);
nand U19157 (N_19157,N_18235,N_18816);
xnor U19158 (N_19158,N_18866,N_18455);
nand U19159 (N_19159,N_18365,N_18122);
and U19160 (N_19160,N_18463,N_18115);
or U19161 (N_19161,N_18264,N_18596);
nor U19162 (N_19162,N_18384,N_18823);
or U19163 (N_19163,N_18149,N_18373);
nand U19164 (N_19164,N_18428,N_18761);
and U19165 (N_19165,N_18165,N_18572);
or U19166 (N_19166,N_18503,N_18389);
and U19167 (N_19167,N_18251,N_18019);
or U19168 (N_19168,N_18650,N_18490);
and U19169 (N_19169,N_18340,N_18754);
or U19170 (N_19170,N_18805,N_18489);
nor U19171 (N_19171,N_18333,N_18083);
nor U19172 (N_19172,N_18720,N_18453);
nand U19173 (N_19173,N_18491,N_18785);
and U19174 (N_19174,N_18269,N_18014);
nand U19175 (N_19175,N_18879,N_18245);
and U19176 (N_19176,N_18506,N_18781);
nor U19177 (N_19177,N_18247,N_18829);
xor U19178 (N_19178,N_18216,N_18075);
xnor U19179 (N_19179,N_18044,N_18708);
and U19180 (N_19180,N_18782,N_18659);
nor U19181 (N_19181,N_18378,N_18290);
and U19182 (N_19182,N_18241,N_18386);
nor U19183 (N_19183,N_18945,N_18404);
or U19184 (N_19184,N_18919,N_18555);
nor U19185 (N_19185,N_18224,N_18895);
xor U19186 (N_19186,N_18150,N_18824);
nand U19187 (N_19187,N_18817,N_18076);
or U19188 (N_19188,N_18230,N_18478);
and U19189 (N_19189,N_18797,N_18700);
nor U19190 (N_19190,N_18561,N_18877);
and U19191 (N_19191,N_18541,N_18534);
nand U19192 (N_19192,N_18563,N_18896);
and U19193 (N_19193,N_18306,N_18319);
and U19194 (N_19194,N_18680,N_18900);
nor U19195 (N_19195,N_18951,N_18841);
nand U19196 (N_19196,N_18606,N_18588);
xnor U19197 (N_19197,N_18470,N_18124);
or U19198 (N_19198,N_18142,N_18998);
nand U19199 (N_19199,N_18111,N_18139);
nor U19200 (N_19200,N_18125,N_18437);
nand U19201 (N_19201,N_18999,N_18493);
and U19202 (N_19202,N_18522,N_18535);
or U19203 (N_19203,N_18448,N_18811);
and U19204 (N_19204,N_18581,N_18414);
nand U19205 (N_19205,N_18813,N_18980);
or U19206 (N_19206,N_18010,N_18120);
or U19207 (N_19207,N_18312,N_18148);
nor U19208 (N_19208,N_18858,N_18946);
xor U19209 (N_19209,N_18121,N_18668);
or U19210 (N_19210,N_18164,N_18836);
nand U19211 (N_19211,N_18021,N_18657);
xor U19212 (N_19212,N_18893,N_18473);
and U19213 (N_19213,N_18684,N_18421);
and U19214 (N_19214,N_18332,N_18394);
nand U19215 (N_19215,N_18598,N_18809);
xnor U19216 (N_19216,N_18145,N_18871);
or U19217 (N_19217,N_18250,N_18526);
nor U19218 (N_19218,N_18923,N_18186);
nor U19219 (N_19219,N_18729,N_18114);
nand U19220 (N_19220,N_18970,N_18078);
nand U19221 (N_19221,N_18517,N_18976);
nor U19222 (N_19222,N_18718,N_18254);
and U19223 (N_19223,N_18238,N_18003);
and U19224 (N_19224,N_18313,N_18085);
xor U19225 (N_19225,N_18314,N_18353);
nor U19226 (N_19226,N_18909,N_18347);
xnor U19227 (N_19227,N_18530,N_18277);
nand U19228 (N_19228,N_18772,N_18272);
xor U19229 (N_19229,N_18681,N_18519);
xnor U19230 (N_19230,N_18759,N_18869);
xnor U19231 (N_19231,N_18016,N_18131);
xnor U19232 (N_19232,N_18012,N_18265);
nor U19233 (N_19233,N_18454,N_18664);
nand U19234 (N_19234,N_18356,N_18102);
nand U19235 (N_19235,N_18529,N_18284);
xor U19236 (N_19236,N_18898,N_18579);
or U19237 (N_19237,N_18791,N_18752);
xnor U19238 (N_19238,N_18843,N_18001);
nand U19239 (N_19239,N_18136,N_18721);
xor U19240 (N_19240,N_18660,N_18556);
nand U19241 (N_19241,N_18550,N_18964);
or U19242 (N_19242,N_18986,N_18328);
xor U19243 (N_19243,N_18586,N_18971);
xnor U19244 (N_19244,N_18651,N_18479);
xor U19245 (N_19245,N_18431,N_18605);
nor U19246 (N_19246,N_18316,N_18468);
xnor U19247 (N_19247,N_18582,N_18279);
or U19248 (N_19248,N_18638,N_18198);
nand U19249 (N_19249,N_18884,N_18323);
xnor U19250 (N_19250,N_18631,N_18762);
nor U19251 (N_19251,N_18907,N_18402);
and U19252 (N_19252,N_18413,N_18965);
nand U19253 (N_19253,N_18617,N_18459);
nand U19254 (N_19254,N_18616,N_18226);
xor U19255 (N_19255,N_18742,N_18180);
xnor U19256 (N_19256,N_18472,N_18475);
and U19257 (N_19257,N_18857,N_18248);
nand U19258 (N_19258,N_18977,N_18006);
xor U19259 (N_19259,N_18427,N_18177);
xor U19260 (N_19260,N_18850,N_18501);
or U19261 (N_19261,N_18485,N_18170);
xnor U19262 (N_19262,N_18737,N_18846);
or U19263 (N_19263,N_18749,N_18702);
and U19264 (N_19264,N_18840,N_18181);
xor U19265 (N_19265,N_18920,N_18342);
xnor U19266 (N_19266,N_18691,N_18667);
xnor U19267 (N_19267,N_18724,N_18296);
nand U19268 (N_19268,N_18822,N_18623);
and U19269 (N_19269,N_18308,N_18542);
nor U19270 (N_19270,N_18106,N_18525);
nor U19271 (N_19271,N_18028,N_18218);
and U19272 (N_19272,N_18495,N_18796);
nor U19273 (N_19273,N_18458,N_18183);
or U19274 (N_19274,N_18887,N_18804);
nand U19275 (N_19275,N_18787,N_18292);
nor U19276 (N_19276,N_18444,N_18046);
xor U19277 (N_19277,N_18995,N_18203);
and U19278 (N_19278,N_18281,N_18642);
and U19279 (N_19279,N_18204,N_18031);
or U19280 (N_19280,N_18465,N_18439);
xnor U19281 (N_19281,N_18169,N_18185);
or U19282 (N_19282,N_18835,N_18908);
or U19283 (N_19283,N_18062,N_18143);
nor U19284 (N_19284,N_18132,N_18765);
nor U19285 (N_19285,N_18476,N_18190);
and U19286 (N_19286,N_18630,N_18416);
or U19287 (N_19287,N_18058,N_18979);
nor U19288 (N_19288,N_18168,N_18112);
and U19289 (N_19289,N_18362,N_18430);
or U19290 (N_19290,N_18928,N_18988);
xnor U19291 (N_19291,N_18462,N_18571);
or U19292 (N_19292,N_18656,N_18904);
nand U19293 (N_19293,N_18045,N_18041);
xor U19294 (N_19294,N_18270,N_18377);
nor U19295 (N_19295,N_18856,N_18806);
or U19296 (N_19296,N_18514,N_18918);
xnor U19297 (N_19297,N_18756,N_18159);
nor U19298 (N_19298,N_18774,N_18081);
nor U19299 (N_19299,N_18679,N_18304);
and U19300 (N_19300,N_18873,N_18067);
or U19301 (N_19301,N_18233,N_18875);
or U19302 (N_19302,N_18842,N_18549);
nor U19303 (N_19303,N_18820,N_18917);
nand U19304 (N_19304,N_18675,N_18236);
xor U19305 (N_19305,N_18282,N_18925);
nand U19306 (N_19306,N_18624,N_18302);
and U19307 (N_19307,N_18504,N_18257);
and U19308 (N_19308,N_18412,N_18271);
nand U19309 (N_19309,N_18246,N_18669);
nor U19310 (N_19310,N_18484,N_18983);
or U19311 (N_19311,N_18049,N_18352);
and U19312 (N_19312,N_18601,N_18424);
xnor U19313 (N_19313,N_18643,N_18768);
nand U19314 (N_19314,N_18770,N_18595);
xor U19315 (N_19315,N_18217,N_18162);
or U19316 (N_19316,N_18291,N_18116);
and U19317 (N_19317,N_18939,N_18574);
nand U19318 (N_19318,N_18171,N_18859);
and U19319 (N_19319,N_18828,N_18208);
or U19320 (N_19320,N_18442,N_18903);
nand U19321 (N_19321,N_18206,N_18295);
or U19322 (N_19322,N_18433,N_18073);
or U19323 (N_19323,N_18798,N_18803);
or U19324 (N_19324,N_18151,N_18403);
nand U19325 (N_19325,N_18810,N_18655);
nor U19326 (N_19326,N_18883,N_18728);
and U19327 (N_19327,N_18789,N_18665);
nor U19328 (N_19328,N_18769,N_18710);
xnor U19329 (N_19329,N_18715,N_18639);
nor U19330 (N_19330,N_18343,N_18524);
or U19331 (N_19331,N_18117,N_18851);
nand U19332 (N_19332,N_18227,N_18374);
or U19333 (N_19333,N_18419,N_18080);
nor U19334 (N_19334,N_18981,N_18024);
xor U19335 (N_19335,N_18627,N_18199);
xnor U19336 (N_19336,N_18456,N_18558);
and U19337 (N_19337,N_18944,N_18130);
or U19338 (N_19338,N_18207,N_18423);
xnor U19339 (N_19339,N_18750,N_18042);
nor U19340 (N_19340,N_18714,N_18966);
nor U19341 (N_19341,N_18381,N_18845);
nor U19342 (N_19342,N_18098,N_18794);
nor U19343 (N_19343,N_18626,N_18364);
or U19344 (N_19344,N_18422,N_18648);
nor U19345 (N_19345,N_18383,N_18447);
nor U19346 (N_19346,N_18360,N_18370);
or U19347 (N_19347,N_18731,N_18093);
or U19348 (N_19348,N_18411,N_18544);
or U19349 (N_19349,N_18065,N_18020);
xnor U19350 (N_19350,N_18299,N_18758);
and U19351 (N_19351,N_18773,N_18449);
nor U19352 (N_19352,N_18830,N_18187);
or U19353 (N_19353,N_18426,N_18082);
nor U19354 (N_19354,N_18097,N_18420);
or U19355 (N_19355,N_18634,N_18784);
and U19356 (N_19356,N_18670,N_18258);
xnor U19357 (N_19357,N_18954,N_18334);
nand U19358 (N_19358,N_18367,N_18398);
nor U19359 (N_19359,N_18932,N_18609);
or U19360 (N_19360,N_18050,N_18406);
and U19361 (N_19361,N_18635,N_18392);
nor U19362 (N_19362,N_18989,N_18897);
or U19363 (N_19363,N_18704,N_18527);
nand U19364 (N_19364,N_18933,N_18950);
and U19365 (N_19365,N_18074,N_18600);
or U19366 (N_19366,N_18593,N_18294);
and U19367 (N_19367,N_18800,N_18972);
and U19368 (N_19368,N_18234,N_18914);
nand U19369 (N_19369,N_18834,N_18839);
and U19370 (N_19370,N_18521,N_18973);
xor U19371 (N_19371,N_18211,N_18947);
nor U19372 (N_19372,N_18613,N_18240);
nor U19373 (N_19373,N_18985,N_18103);
xnor U19374 (N_19374,N_18104,N_18553);
and U19375 (N_19375,N_18396,N_18215);
nor U19376 (N_19376,N_18968,N_18301);
xor U19377 (N_19377,N_18432,N_18274);
nand U19378 (N_19378,N_18926,N_18687);
xnor U19379 (N_19379,N_18182,N_18037);
or U19380 (N_19380,N_18975,N_18633);
nor U19381 (N_19381,N_18523,N_18992);
nor U19382 (N_19382,N_18753,N_18385);
nand U19383 (N_19383,N_18929,N_18191);
xor U19384 (N_19384,N_18927,N_18825);
and U19385 (N_19385,N_18509,N_18629);
nand U19386 (N_19386,N_18436,N_18735);
nor U19387 (N_19387,N_18860,N_18786);
and U19388 (N_19388,N_18955,N_18004);
nor U19389 (N_19389,N_18747,N_18002);
or U19390 (N_19390,N_18991,N_18173);
nand U19391 (N_19391,N_18508,N_18212);
nor U19392 (N_19392,N_18146,N_18309);
nor U19393 (N_19393,N_18936,N_18799);
nor U19394 (N_19394,N_18862,N_18621);
nand U19395 (N_19395,N_18899,N_18369);
nand U19396 (N_19396,N_18894,N_18244);
and U19397 (N_19397,N_18528,N_18137);
nand U19398 (N_19398,N_18872,N_18357);
or U19399 (N_19399,N_18924,N_18231);
nor U19400 (N_19400,N_18368,N_18647);
nand U19401 (N_19401,N_18949,N_18637);
and U19402 (N_19402,N_18013,N_18599);
or U19403 (N_19403,N_18706,N_18916);
and U19404 (N_19404,N_18646,N_18719);
nand U19405 (N_19405,N_18692,N_18415);
xnor U19406 (N_19406,N_18958,N_18321);
and U19407 (N_19407,N_18610,N_18486);
and U19408 (N_19408,N_18361,N_18052);
and U19409 (N_19409,N_18507,N_18391);
and U19410 (N_19410,N_18339,N_18026);
xnor U19411 (N_19411,N_18163,N_18818);
xor U19412 (N_19412,N_18801,N_18223);
and U19413 (N_19413,N_18069,N_18674);
or U19414 (N_19414,N_18158,N_18488);
or U19415 (N_19415,N_18088,N_18960);
nand U19416 (N_19416,N_18990,N_18748);
and U19417 (N_19417,N_18161,N_18956);
and U19418 (N_19418,N_18864,N_18832);
nor U19419 (N_19419,N_18745,N_18355);
xor U19420 (N_19420,N_18539,N_18602);
or U19421 (N_19421,N_18133,N_18953);
and U19422 (N_19422,N_18084,N_18699);
or U19423 (N_19423,N_18537,N_18070);
nand U19424 (N_19424,N_18578,N_18716);
or U19425 (N_19425,N_18778,N_18863);
nor U19426 (N_19426,N_18278,N_18622);
nand U19427 (N_19427,N_18263,N_18777);
or U19428 (N_19428,N_18536,N_18705);
xnor U19429 (N_19429,N_18576,N_18166);
and U19430 (N_19430,N_18446,N_18570);
nand U19431 (N_19431,N_18515,N_18252);
or U19432 (N_19432,N_18726,N_18134);
xor U19433 (N_19433,N_18741,N_18861);
or U19434 (N_19434,N_18201,N_18967);
xnor U19435 (N_19435,N_18249,N_18039);
nand U19436 (N_19436,N_18940,N_18390);
or U19437 (N_19437,N_18755,N_18127);
or U19438 (N_19438,N_18000,N_18683);
nand U19439 (N_19439,N_18029,N_18591);
xnor U19440 (N_19440,N_18723,N_18481);
xor U19441 (N_19441,N_18994,N_18315);
nor U19442 (N_19442,N_18141,N_18079);
or U19443 (N_19443,N_18653,N_18387);
and U19444 (N_19444,N_18910,N_18195);
and U19445 (N_19445,N_18722,N_18788);
or U19446 (N_19446,N_18821,N_18625);
and U19447 (N_19447,N_18614,N_18094);
nand U19448 (N_19448,N_18573,N_18963);
xnor U19449 (N_19449,N_18327,N_18996);
nor U19450 (N_19450,N_18854,N_18409);
xor U19451 (N_19451,N_18113,N_18764);
nand U19452 (N_19452,N_18289,N_18033);
or U19453 (N_19453,N_18780,N_18027);
nor U19454 (N_19454,N_18036,N_18695);
xor U19455 (N_19455,N_18051,N_18628);
and U19456 (N_19456,N_18174,N_18891);
xor U19457 (N_19457,N_18827,N_18200);
or U19458 (N_19458,N_18688,N_18435);
and U19459 (N_19459,N_18337,N_18513);
xor U19460 (N_19460,N_18733,N_18494);
nor U19461 (N_19461,N_18135,N_18776);
nand U19462 (N_19462,N_18382,N_18425);
nand U19463 (N_19463,N_18059,N_18833);
or U19464 (N_19464,N_18096,N_18018);
xnor U19465 (N_19465,N_18354,N_18562);
xnor U19466 (N_19466,N_18376,N_18795);
and U19467 (N_19467,N_18009,N_18157);
or U19468 (N_19468,N_18259,N_18118);
nor U19469 (N_19469,N_18767,N_18219);
xnor U19470 (N_19470,N_18746,N_18228);
and U19471 (N_19471,N_18022,N_18154);
nor U19472 (N_19472,N_18775,N_18580);
and U19473 (N_19473,N_18214,N_18338);
xnor U19474 (N_19474,N_18696,N_18913);
and U19475 (N_19475,N_18293,N_18615);
nor U19476 (N_19476,N_18176,N_18959);
nand U19477 (N_19477,N_18592,N_18847);
nand U19478 (N_19478,N_18129,N_18620);
nand U19479 (N_19479,N_18911,N_18751);
and U19480 (N_19480,N_18189,N_18545);
xnor U19481 (N_19481,N_18325,N_18676);
nor U19482 (N_19482,N_18184,N_18987);
xnor U19483 (N_19483,N_18645,N_18740);
or U19484 (N_19484,N_18007,N_18071);
xnor U19485 (N_19485,N_18372,N_18962);
and U19486 (N_19486,N_18242,N_18948);
xnor U19487 (N_19487,N_18779,N_18099);
nor U19488 (N_19488,N_18957,N_18087);
and U19489 (N_19489,N_18063,N_18790);
nand U19490 (N_19490,N_18935,N_18089);
nor U19491 (N_19491,N_18110,N_18043);
nor U19492 (N_19492,N_18886,N_18632);
xnor U19493 (N_19493,N_18466,N_18557);
or U19494 (N_19494,N_18640,N_18568);
nor U19495 (N_19495,N_18649,N_18868);
nor U19496 (N_19496,N_18061,N_18038);
xor U19497 (N_19497,N_18108,N_18175);
nor U19498 (N_19498,N_18477,N_18902);
xor U19499 (N_19499,N_18153,N_18658);
and U19500 (N_19500,N_18369,N_18592);
and U19501 (N_19501,N_18074,N_18809);
nand U19502 (N_19502,N_18749,N_18794);
or U19503 (N_19503,N_18238,N_18769);
and U19504 (N_19504,N_18126,N_18640);
or U19505 (N_19505,N_18655,N_18758);
or U19506 (N_19506,N_18226,N_18166);
nand U19507 (N_19507,N_18379,N_18900);
or U19508 (N_19508,N_18648,N_18128);
nor U19509 (N_19509,N_18630,N_18403);
nand U19510 (N_19510,N_18291,N_18874);
or U19511 (N_19511,N_18902,N_18685);
xor U19512 (N_19512,N_18747,N_18340);
xor U19513 (N_19513,N_18373,N_18529);
or U19514 (N_19514,N_18971,N_18600);
nor U19515 (N_19515,N_18181,N_18176);
or U19516 (N_19516,N_18614,N_18105);
or U19517 (N_19517,N_18630,N_18057);
nor U19518 (N_19518,N_18286,N_18891);
or U19519 (N_19519,N_18700,N_18495);
or U19520 (N_19520,N_18551,N_18620);
nor U19521 (N_19521,N_18526,N_18814);
nand U19522 (N_19522,N_18312,N_18799);
xnor U19523 (N_19523,N_18362,N_18915);
xor U19524 (N_19524,N_18378,N_18828);
nand U19525 (N_19525,N_18154,N_18779);
xnor U19526 (N_19526,N_18781,N_18690);
and U19527 (N_19527,N_18349,N_18340);
and U19528 (N_19528,N_18107,N_18704);
xor U19529 (N_19529,N_18083,N_18951);
or U19530 (N_19530,N_18158,N_18436);
nor U19531 (N_19531,N_18573,N_18255);
xnor U19532 (N_19532,N_18564,N_18654);
xor U19533 (N_19533,N_18881,N_18985);
or U19534 (N_19534,N_18987,N_18702);
and U19535 (N_19535,N_18979,N_18758);
and U19536 (N_19536,N_18494,N_18371);
or U19537 (N_19537,N_18128,N_18193);
and U19538 (N_19538,N_18268,N_18745);
or U19539 (N_19539,N_18673,N_18185);
and U19540 (N_19540,N_18380,N_18076);
nand U19541 (N_19541,N_18678,N_18120);
nand U19542 (N_19542,N_18774,N_18236);
or U19543 (N_19543,N_18638,N_18460);
or U19544 (N_19544,N_18684,N_18213);
and U19545 (N_19545,N_18361,N_18538);
or U19546 (N_19546,N_18645,N_18230);
and U19547 (N_19547,N_18923,N_18974);
xnor U19548 (N_19548,N_18050,N_18845);
nand U19549 (N_19549,N_18366,N_18976);
and U19550 (N_19550,N_18468,N_18262);
and U19551 (N_19551,N_18436,N_18912);
xnor U19552 (N_19552,N_18016,N_18678);
xor U19553 (N_19553,N_18992,N_18147);
nor U19554 (N_19554,N_18668,N_18927);
nand U19555 (N_19555,N_18679,N_18113);
nor U19556 (N_19556,N_18067,N_18878);
nand U19557 (N_19557,N_18278,N_18322);
nor U19558 (N_19558,N_18047,N_18161);
nor U19559 (N_19559,N_18396,N_18811);
nand U19560 (N_19560,N_18185,N_18081);
xor U19561 (N_19561,N_18092,N_18626);
or U19562 (N_19562,N_18548,N_18177);
xnor U19563 (N_19563,N_18983,N_18587);
and U19564 (N_19564,N_18141,N_18685);
nor U19565 (N_19565,N_18340,N_18447);
and U19566 (N_19566,N_18988,N_18520);
and U19567 (N_19567,N_18349,N_18788);
nand U19568 (N_19568,N_18780,N_18207);
or U19569 (N_19569,N_18444,N_18998);
xnor U19570 (N_19570,N_18761,N_18317);
xnor U19571 (N_19571,N_18176,N_18359);
xnor U19572 (N_19572,N_18188,N_18696);
nor U19573 (N_19573,N_18892,N_18373);
and U19574 (N_19574,N_18739,N_18423);
and U19575 (N_19575,N_18089,N_18021);
and U19576 (N_19576,N_18241,N_18934);
and U19577 (N_19577,N_18534,N_18088);
nand U19578 (N_19578,N_18419,N_18390);
and U19579 (N_19579,N_18720,N_18037);
and U19580 (N_19580,N_18342,N_18471);
or U19581 (N_19581,N_18226,N_18458);
xor U19582 (N_19582,N_18030,N_18065);
and U19583 (N_19583,N_18607,N_18436);
xor U19584 (N_19584,N_18344,N_18859);
and U19585 (N_19585,N_18620,N_18425);
nor U19586 (N_19586,N_18863,N_18994);
xor U19587 (N_19587,N_18537,N_18269);
or U19588 (N_19588,N_18232,N_18431);
nand U19589 (N_19589,N_18442,N_18600);
and U19590 (N_19590,N_18305,N_18636);
and U19591 (N_19591,N_18775,N_18475);
nor U19592 (N_19592,N_18620,N_18804);
xnor U19593 (N_19593,N_18084,N_18333);
nand U19594 (N_19594,N_18019,N_18324);
nand U19595 (N_19595,N_18775,N_18118);
nand U19596 (N_19596,N_18323,N_18841);
nor U19597 (N_19597,N_18598,N_18715);
xor U19598 (N_19598,N_18761,N_18440);
xnor U19599 (N_19599,N_18906,N_18919);
nor U19600 (N_19600,N_18386,N_18804);
nand U19601 (N_19601,N_18230,N_18075);
or U19602 (N_19602,N_18183,N_18583);
xor U19603 (N_19603,N_18302,N_18108);
and U19604 (N_19604,N_18095,N_18547);
or U19605 (N_19605,N_18021,N_18205);
nand U19606 (N_19606,N_18272,N_18335);
or U19607 (N_19607,N_18020,N_18399);
nor U19608 (N_19608,N_18429,N_18763);
nor U19609 (N_19609,N_18495,N_18907);
nor U19610 (N_19610,N_18028,N_18373);
xnor U19611 (N_19611,N_18343,N_18258);
or U19612 (N_19612,N_18413,N_18453);
and U19613 (N_19613,N_18794,N_18114);
and U19614 (N_19614,N_18116,N_18069);
or U19615 (N_19615,N_18185,N_18920);
nand U19616 (N_19616,N_18491,N_18488);
nor U19617 (N_19617,N_18016,N_18525);
xnor U19618 (N_19618,N_18917,N_18120);
xor U19619 (N_19619,N_18220,N_18174);
or U19620 (N_19620,N_18276,N_18899);
xnor U19621 (N_19621,N_18692,N_18238);
nand U19622 (N_19622,N_18559,N_18410);
and U19623 (N_19623,N_18606,N_18489);
nor U19624 (N_19624,N_18057,N_18379);
nand U19625 (N_19625,N_18157,N_18415);
nand U19626 (N_19626,N_18698,N_18905);
nand U19627 (N_19627,N_18125,N_18492);
xor U19628 (N_19628,N_18336,N_18842);
nand U19629 (N_19629,N_18124,N_18342);
xnor U19630 (N_19630,N_18359,N_18123);
nor U19631 (N_19631,N_18324,N_18330);
xnor U19632 (N_19632,N_18319,N_18925);
nand U19633 (N_19633,N_18834,N_18661);
nor U19634 (N_19634,N_18974,N_18451);
and U19635 (N_19635,N_18040,N_18466);
nand U19636 (N_19636,N_18212,N_18715);
xor U19637 (N_19637,N_18045,N_18375);
xnor U19638 (N_19638,N_18099,N_18821);
or U19639 (N_19639,N_18108,N_18344);
xor U19640 (N_19640,N_18544,N_18909);
nor U19641 (N_19641,N_18538,N_18444);
and U19642 (N_19642,N_18855,N_18321);
or U19643 (N_19643,N_18738,N_18018);
xnor U19644 (N_19644,N_18613,N_18126);
and U19645 (N_19645,N_18278,N_18408);
nor U19646 (N_19646,N_18669,N_18966);
nand U19647 (N_19647,N_18070,N_18667);
xnor U19648 (N_19648,N_18009,N_18077);
nand U19649 (N_19649,N_18926,N_18650);
nor U19650 (N_19650,N_18634,N_18242);
nor U19651 (N_19651,N_18068,N_18276);
nand U19652 (N_19652,N_18588,N_18354);
and U19653 (N_19653,N_18733,N_18808);
nor U19654 (N_19654,N_18828,N_18730);
nor U19655 (N_19655,N_18533,N_18354);
and U19656 (N_19656,N_18758,N_18646);
or U19657 (N_19657,N_18287,N_18886);
and U19658 (N_19658,N_18710,N_18131);
and U19659 (N_19659,N_18097,N_18311);
nand U19660 (N_19660,N_18623,N_18713);
or U19661 (N_19661,N_18355,N_18207);
xnor U19662 (N_19662,N_18630,N_18926);
or U19663 (N_19663,N_18394,N_18824);
nor U19664 (N_19664,N_18006,N_18272);
and U19665 (N_19665,N_18132,N_18832);
nor U19666 (N_19666,N_18700,N_18667);
nand U19667 (N_19667,N_18307,N_18494);
nand U19668 (N_19668,N_18871,N_18276);
nor U19669 (N_19669,N_18333,N_18180);
nand U19670 (N_19670,N_18972,N_18237);
xor U19671 (N_19671,N_18203,N_18194);
nor U19672 (N_19672,N_18034,N_18037);
xor U19673 (N_19673,N_18826,N_18113);
and U19674 (N_19674,N_18908,N_18563);
xor U19675 (N_19675,N_18968,N_18488);
or U19676 (N_19676,N_18791,N_18156);
xor U19677 (N_19677,N_18385,N_18448);
xnor U19678 (N_19678,N_18252,N_18489);
and U19679 (N_19679,N_18361,N_18623);
or U19680 (N_19680,N_18601,N_18258);
nor U19681 (N_19681,N_18609,N_18951);
and U19682 (N_19682,N_18955,N_18823);
xnor U19683 (N_19683,N_18703,N_18802);
nor U19684 (N_19684,N_18286,N_18682);
nand U19685 (N_19685,N_18298,N_18934);
and U19686 (N_19686,N_18369,N_18963);
nor U19687 (N_19687,N_18451,N_18469);
or U19688 (N_19688,N_18271,N_18586);
or U19689 (N_19689,N_18306,N_18283);
xor U19690 (N_19690,N_18324,N_18798);
xnor U19691 (N_19691,N_18528,N_18293);
xnor U19692 (N_19692,N_18771,N_18383);
and U19693 (N_19693,N_18971,N_18995);
and U19694 (N_19694,N_18257,N_18447);
or U19695 (N_19695,N_18663,N_18948);
xor U19696 (N_19696,N_18909,N_18057);
nand U19697 (N_19697,N_18313,N_18470);
and U19698 (N_19698,N_18569,N_18128);
or U19699 (N_19699,N_18717,N_18066);
and U19700 (N_19700,N_18497,N_18460);
and U19701 (N_19701,N_18014,N_18177);
nor U19702 (N_19702,N_18111,N_18712);
nand U19703 (N_19703,N_18511,N_18314);
xor U19704 (N_19704,N_18827,N_18247);
nand U19705 (N_19705,N_18820,N_18815);
xor U19706 (N_19706,N_18328,N_18829);
xnor U19707 (N_19707,N_18105,N_18200);
xnor U19708 (N_19708,N_18320,N_18645);
xnor U19709 (N_19709,N_18765,N_18900);
xnor U19710 (N_19710,N_18760,N_18090);
or U19711 (N_19711,N_18321,N_18325);
xor U19712 (N_19712,N_18964,N_18605);
nor U19713 (N_19713,N_18031,N_18913);
xnor U19714 (N_19714,N_18417,N_18708);
xor U19715 (N_19715,N_18796,N_18328);
and U19716 (N_19716,N_18295,N_18641);
and U19717 (N_19717,N_18384,N_18952);
and U19718 (N_19718,N_18470,N_18210);
xor U19719 (N_19719,N_18539,N_18593);
and U19720 (N_19720,N_18293,N_18816);
nand U19721 (N_19721,N_18193,N_18884);
nor U19722 (N_19722,N_18728,N_18477);
xnor U19723 (N_19723,N_18834,N_18869);
nor U19724 (N_19724,N_18725,N_18408);
and U19725 (N_19725,N_18868,N_18946);
and U19726 (N_19726,N_18765,N_18982);
xnor U19727 (N_19727,N_18568,N_18643);
nor U19728 (N_19728,N_18321,N_18521);
and U19729 (N_19729,N_18384,N_18473);
nor U19730 (N_19730,N_18757,N_18055);
xor U19731 (N_19731,N_18732,N_18814);
xor U19732 (N_19732,N_18789,N_18995);
or U19733 (N_19733,N_18787,N_18843);
nor U19734 (N_19734,N_18807,N_18482);
nand U19735 (N_19735,N_18949,N_18600);
or U19736 (N_19736,N_18783,N_18092);
xor U19737 (N_19737,N_18909,N_18935);
or U19738 (N_19738,N_18466,N_18856);
nand U19739 (N_19739,N_18823,N_18285);
and U19740 (N_19740,N_18546,N_18977);
or U19741 (N_19741,N_18576,N_18939);
or U19742 (N_19742,N_18830,N_18123);
nand U19743 (N_19743,N_18157,N_18626);
nor U19744 (N_19744,N_18480,N_18673);
or U19745 (N_19745,N_18507,N_18291);
and U19746 (N_19746,N_18279,N_18584);
xor U19747 (N_19747,N_18811,N_18092);
or U19748 (N_19748,N_18709,N_18613);
and U19749 (N_19749,N_18631,N_18104);
nand U19750 (N_19750,N_18847,N_18988);
nor U19751 (N_19751,N_18888,N_18168);
or U19752 (N_19752,N_18790,N_18650);
and U19753 (N_19753,N_18151,N_18058);
nand U19754 (N_19754,N_18419,N_18255);
nand U19755 (N_19755,N_18203,N_18243);
nor U19756 (N_19756,N_18498,N_18404);
and U19757 (N_19757,N_18502,N_18146);
nor U19758 (N_19758,N_18728,N_18802);
nand U19759 (N_19759,N_18825,N_18710);
or U19760 (N_19760,N_18673,N_18942);
nor U19761 (N_19761,N_18109,N_18132);
xor U19762 (N_19762,N_18049,N_18584);
nand U19763 (N_19763,N_18948,N_18272);
and U19764 (N_19764,N_18096,N_18935);
xor U19765 (N_19765,N_18816,N_18182);
nand U19766 (N_19766,N_18090,N_18503);
xnor U19767 (N_19767,N_18664,N_18048);
xnor U19768 (N_19768,N_18863,N_18110);
or U19769 (N_19769,N_18596,N_18850);
xor U19770 (N_19770,N_18722,N_18245);
nand U19771 (N_19771,N_18137,N_18926);
xor U19772 (N_19772,N_18431,N_18745);
xnor U19773 (N_19773,N_18784,N_18611);
nor U19774 (N_19774,N_18016,N_18177);
and U19775 (N_19775,N_18892,N_18694);
nor U19776 (N_19776,N_18060,N_18947);
xnor U19777 (N_19777,N_18642,N_18821);
nand U19778 (N_19778,N_18747,N_18056);
nor U19779 (N_19779,N_18615,N_18094);
nand U19780 (N_19780,N_18085,N_18053);
nor U19781 (N_19781,N_18345,N_18567);
and U19782 (N_19782,N_18193,N_18405);
nor U19783 (N_19783,N_18778,N_18204);
xnor U19784 (N_19784,N_18634,N_18165);
nor U19785 (N_19785,N_18179,N_18514);
or U19786 (N_19786,N_18310,N_18796);
nor U19787 (N_19787,N_18526,N_18198);
or U19788 (N_19788,N_18714,N_18200);
nor U19789 (N_19789,N_18963,N_18415);
nand U19790 (N_19790,N_18384,N_18796);
and U19791 (N_19791,N_18204,N_18585);
or U19792 (N_19792,N_18773,N_18605);
and U19793 (N_19793,N_18659,N_18701);
and U19794 (N_19794,N_18095,N_18199);
nand U19795 (N_19795,N_18494,N_18938);
and U19796 (N_19796,N_18630,N_18267);
nand U19797 (N_19797,N_18756,N_18190);
xnor U19798 (N_19798,N_18787,N_18553);
and U19799 (N_19799,N_18166,N_18097);
and U19800 (N_19800,N_18932,N_18885);
nor U19801 (N_19801,N_18569,N_18814);
xor U19802 (N_19802,N_18258,N_18528);
xor U19803 (N_19803,N_18233,N_18171);
nor U19804 (N_19804,N_18709,N_18184);
and U19805 (N_19805,N_18330,N_18915);
xnor U19806 (N_19806,N_18778,N_18482);
and U19807 (N_19807,N_18456,N_18716);
xnor U19808 (N_19808,N_18988,N_18169);
and U19809 (N_19809,N_18383,N_18320);
or U19810 (N_19810,N_18171,N_18526);
nand U19811 (N_19811,N_18992,N_18182);
xnor U19812 (N_19812,N_18086,N_18962);
or U19813 (N_19813,N_18534,N_18784);
or U19814 (N_19814,N_18391,N_18518);
nand U19815 (N_19815,N_18102,N_18981);
nor U19816 (N_19816,N_18084,N_18964);
and U19817 (N_19817,N_18157,N_18303);
xor U19818 (N_19818,N_18599,N_18430);
and U19819 (N_19819,N_18005,N_18490);
nand U19820 (N_19820,N_18572,N_18407);
xor U19821 (N_19821,N_18059,N_18566);
or U19822 (N_19822,N_18898,N_18650);
nand U19823 (N_19823,N_18744,N_18529);
nor U19824 (N_19824,N_18470,N_18501);
nand U19825 (N_19825,N_18380,N_18729);
nand U19826 (N_19826,N_18220,N_18057);
or U19827 (N_19827,N_18187,N_18010);
nor U19828 (N_19828,N_18261,N_18961);
nand U19829 (N_19829,N_18871,N_18183);
or U19830 (N_19830,N_18182,N_18225);
or U19831 (N_19831,N_18193,N_18835);
nand U19832 (N_19832,N_18856,N_18927);
nand U19833 (N_19833,N_18057,N_18139);
nor U19834 (N_19834,N_18347,N_18034);
nor U19835 (N_19835,N_18561,N_18088);
xnor U19836 (N_19836,N_18569,N_18664);
or U19837 (N_19837,N_18629,N_18367);
nand U19838 (N_19838,N_18631,N_18034);
or U19839 (N_19839,N_18972,N_18616);
nor U19840 (N_19840,N_18211,N_18331);
xor U19841 (N_19841,N_18308,N_18544);
xor U19842 (N_19842,N_18958,N_18221);
xnor U19843 (N_19843,N_18266,N_18402);
or U19844 (N_19844,N_18515,N_18147);
nand U19845 (N_19845,N_18452,N_18414);
xor U19846 (N_19846,N_18363,N_18631);
and U19847 (N_19847,N_18097,N_18708);
or U19848 (N_19848,N_18276,N_18192);
xnor U19849 (N_19849,N_18214,N_18618);
xor U19850 (N_19850,N_18998,N_18915);
and U19851 (N_19851,N_18553,N_18914);
nand U19852 (N_19852,N_18576,N_18548);
nand U19853 (N_19853,N_18638,N_18818);
or U19854 (N_19854,N_18954,N_18033);
nand U19855 (N_19855,N_18873,N_18787);
nand U19856 (N_19856,N_18085,N_18396);
xnor U19857 (N_19857,N_18674,N_18734);
or U19858 (N_19858,N_18664,N_18553);
and U19859 (N_19859,N_18437,N_18243);
and U19860 (N_19860,N_18136,N_18567);
or U19861 (N_19861,N_18670,N_18020);
nand U19862 (N_19862,N_18455,N_18233);
and U19863 (N_19863,N_18143,N_18977);
and U19864 (N_19864,N_18710,N_18783);
or U19865 (N_19865,N_18463,N_18707);
or U19866 (N_19866,N_18005,N_18855);
or U19867 (N_19867,N_18235,N_18884);
or U19868 (N_19868,N_18696,N_18829);
xnor U19869 (N_19869,N_18205,N_18077);
xor U19870 (N_19870,N_18290,N_18347);
and U19871 (N_19871,N_18525,N_18430);
and U19872 (N_19872,N_18548,N_18874);
nor U19873 (N_19873,N_18778,N_18217);
and U19874 (N_19874,N_18319,N_18549);
or U19875 (N_19875,N_18419,N_18105);
xor U19876 (N_19876,N_18353,N_18626);
xor U19877 (N_19877,N_18299,N_18857);
or U19878 (N_19878,N_18363,N_18876);
or U19879 (N_19879,N_18385,N_18539);
nor U19880 (N_19880,N_18853,N_18590);
nand U19881 (N_19881,N_18809,N_18026);
and U19882 (N_19882,N_18760,N_18612);
nand U19883 (N_19883,N_18602,N_18095);
xnor U19884 (N_19884,N_18214,N_18273);
nand U19885 (N_19885,N_18119,N_18860);
xor U19886 (N_19886,N_18552,N_18231);
nor U19887 (N_19887,N_18398,N_18194);
xnor U19888 (N_19888,N_18943,N_18670);
nor U19889 (N_19889,N_18004,N_18780);
nor U19890 (N_19890,N_18576,N_18762);
nor U19891 (N_19891,N_18911,N_18055);
or U19892 (N_19892,N_18444,N_18539);
nand U19893 (N_19893,N_18628,N_18843);
nor U19894 (N_19894,N_18948,N_18796);
nand U19895 (N_19895,N_18273,N_18618);
nor U19896 (N_19896,N_18050,N_18495);
or U19897 (N_19897,N_18225,N_18723);
nor U19898 (N_19898,N_18742,N_18046);
nand U19899 (N_19899,N_18810,N_18308);
or U19900 (N_19900,N_18017,N_18405);
xor U19901 (N_19901,N_18249,N_18376);
nand U19902 (N_19902,N_18438,N_18596);
xnor U19903 (N_19903,N_18484,N_18887);
or U19904 (N_19904,N_18588,N_18090);
nor U19905 (N_19905,N_18737,N_18464);
nor U19906 (N_19906,N_18897,N_18420);
and U19907 (N_19907,N_18856,N_18547);
xor U19908 (N_19908,N_18673,N_18222);
nor U19909 (N_19909,N_18127,N_18178);
nand U19910 (N_19910,N_18806,N_18217);
nand U19911 (N_19911,N_18193,N_18868);
and U19912 (N_19912,N_18391,N_18754);
and U19913 (N_19913,N_18158,N_18903);
nor U19914 (N_19914,N_18763,N_18479);
nand U19915 (N_19915,N_18807,N_18271);
nand U19916 (N_19916,N_18619,N_18371);
nand U19917 (N_19917,N_18205,N_18552);
nor U19918 (N_19918,N_18169,N_18494);
nand U19919 (N_19919,N_18954,N_18686);
nand U19920 (N_19920,N_18248,N_18837);
nor U19921 (N_19921,N_18767,N_18500);
nor U19922 (N_19922,N_18463,N_18594);
nand U19923 (N_19923,N_18021,N_18752);
or U19924 (N_19924,N_18391,N_18222);
and U19925 (N_19925,N_18177,N_18105);
xor U19926 (N_19926,N_18997,N_18773);
xnor U19927 (N_19927,N_18477,N_18472);
nand U19928 (N_19928,N_18491,N_18347);
nor U19929 (N_19929,N_18017,N_18433);
nor U19930 (N_19930,N_18789,N_18786);
and U19931 (N_19931,N_18135,N_18414);
nand U19932 (N_19932,N_18205,N_18942);
and U19933 (N_19933,N_18242,N_18575);
nor U19934 (N_19934,N_18388,N_18666);
nor U19935 (N_19935,N_18864,N_18661);
xnor U19936 (N_19936,N_18371,N_18763);
nand U19937 (N_19937,N_18695,N_18356);
or U19938 (N_19938,N_18217,N_18059);
and U19939 (N_19939,N_18604,N_18329);
xor U19940 (N_19940,N_18127,N_18919);
or U19941 (N_19941,N_18343,N_18207);
nor U19942 (N_19942,N_18410,N_18969);
or U19943 (N_19943,N_18288,N_18646);
xor U19944 (N_19944,N_18522,N_18073);
and U19945 (N_19945,N_18788,N_18662);
nor U19946 (N_19946,N_18888,N_18514);
and U19947 (N_19947,N_18781,N_18481);
nor U19948 (N_19948,N_18461,N_18894);
nor U19949 (N_19949,N_18916,N_18457);
nand U19950 (N_19950,N_18885,N_18253);
or U19951 (N_19951,N_18951,N_18196);
and U19952 (N_19952,N_18405,N_18565);
nand U19953 (N_19953,N_18481,N_18687);
nor U19954 (N_19954,N_18149,N_18817);
nor U19955 (N_19955,N_18626,N_18845);
and U19956 (N_19956,N_18878,N_18700);
nor U19957 (N_19957,N_18551,N_18577);
xor U19958 (N_19958,N_18319,N_18514);
nand U19959 (N_19959,N_18450,N_18462);
xnor U19960 (N_19960,N_18971,N_18067);
nand U19961 (N_19961,N_18312,N_18973);
and U19962 (N_19962,N_18499,N_18380);
xnor U19963 (N_19963,N_18797,N_18137);
nor U19964 (N_19964,N_18510,N_18015);
xnor U19965 (N_19965,N_18174,N_18419);
nor U19966 (N_19966,N_18697,N_18266);
nor U19967 (N_19967,N_18411,N_18163);
xor U19968 (N_19968,N_18543,N_18883);
xor U19969 (N_19969,N_18364,N_18577);
or U19970 (N_19970,N_18574,N_18271);
and U19971 (N_19971,N_18784,N_18670);
and U19972 (N_19972,N_18627,N_18807);
xor U19973 (N_19973,N_18395,N_18397);
nand U19974 (N_19974,N_18538,N_18238);
or U19975 (N_19975,N_18861,N_18843);
nor U19976 (N_19976,N_18441,N_18676);
nand U19977 (N_19977,N_18088,N_18922);
xnor U19978 (N_19978,N_18352,N_18431);
or U19979 (N_19979,N_18713,N_18358);
nand U19980 (N_19980,N_18592,N_18924);
nand U19981 (N_19981,N_18905,N_18789);
xor U19982 (N_19982,N_18133,N_18453);
and U19983 (N_19983,N_18749,N_18399);
xnor U19984 (N_19984,N_18115,N_18501);
xnor U19985 (N_19985,N_18724,N_18329);
xor U19986 (N_19986,N_18625,N_18329);
or U19987 (N_19987,N_18389,N_18066);
and U19988 (N_19988,N_18339,N_18171);
xor U19989 (N_19989,N_18218,N_18565);
and U19990 (N_19990,N_18451,N_18668);
and U19991 (N_19991,N_18263,N_18136);
nor U19992 (N_19992,N_18637,N_18852);
and U19993 (N_19993,N_18647,N_18427);
nor U19994 (N_19994,N_18277,N_18889);
nor U19995 (N_19995,N_18648,N_18624);
nor U19996 (N_19996,N_18071,N_18469);
and U19997 (N_19997,N_18539,N_18711);
and U19998 (N_19998,N_18264,N_18129);
nand U19999 (N_19999,N_18461,N_18791);
xor UO_0 (O_0,N_19389,N_19375);
nor UO_1 (O_1,N_19795,N_19861);
or UO_2 (O_2,N_19292,N_19628);
or UO_3 (O_3,N_19981,N_19313);
and UO_4 (O_4,N_19223,N_19338);
or UO_5 (O_5,N_19351,N_19521);
nor UO_6 (O_6,N_19060,N_19399);
nand UO_7 (O_7,N_19465,N_19341);
xnor UO_8 (O_8,N_19850,N_19691);
nor UO_9 (O_9,N_19961,N_19989);
xor UO_10 (O_10,N_19063,N_19584);
or UO_11 (O_11,N_19992,N_19664);
and UO_12 (O_12,N_19764,N_19071);
and UO_13 (O_13,N_19830,N_19903);
nor UO_14 (O_14,N_19839,N_19394);
nand UO_15 (O_15,N_19626,N_19242);
and UO_16 (O_16,N_19315,N_19878);
nand UO_17 (O_17,N_19382,N_19478);
nand UO_18 (O_18,N_19600,N_19115);
nor UO_19 (O_19,N_19845,N_19704);
nand UO_20 (O_20,N_19350,N_19675);
xor UO_21 (O_21,N_19009,N_19834);
nand UO_22 (O_22,N_19390,N_19291);
or UO_23 (O_23,N_19948,N_19793);
and UO_24 (O_24,N_19235,N_19352);
nor UO_25 (O_25,N_19774,N_19707);
nor UO_26 (O_26,N_19792,N_19544);
xnor UO_27 (O_27,N_19897,N_19416);
or UO_28 (O_28,N_19448,N_19752);
and UO_29 (O_29,N_19611,N_19592);
and UO_30 (O_30,N_19567,N_19965);
or UO_31 (O_31,N_19682,N_19739);
or UO_32 (O_32,N_19210,N_19196);
nor UO_33 (O_33,N_19936,N_19493);
or UO_34 (O_34,N_19028,N_19773);
nor UO_35 (O_35,N_19491,N_19954);
or UO_36 (O_36,N_19634,N_19983);
and UO_37 (O_37,N_19877,N_19179);
nor UO_38 (O_38,N_19650,N_19787);
nor UO_39 (O_39,N_19469,N_19947);
nor UO_40 (O_40,N_19854,N_19255);
nor UO_41 (O_41,N_19804,N_19248);
xor UO_42 (O_42,N_19636,N_19940);
nor UO_43 (O_43,N_19610,N_19320);
nand UO_44 (O_44,N_19464,N_19266);
and UO_45 (O_45,N_19213,N_19109);
or UO_46 (O_46,N_19360,N_19061);
or UO_47 (O_47,N_19186,N_19617);
nand UO_48 (O_48,N_19907,N_19660);
or UO_49 (O_49,N_19005,N_19588);
nand UO_50 (O_50,N_19837,N_19112);
or UO_51 (O_51,N_19128,N_19163);
nor UO_52 (O_52,N_19645,N_19721);
or UO_53 (O_53,N_19011,N_19153);
or UO_54 (O_54,N_19507,N_19539);
and UO_55 (O_55,N_19549,N_19003);
xor UO_56 (O_56,N_19219,N_19101);
and UO_57 (O_57,N_19695,N_19767);
or UO_58 (O_58,N_19287,N_19272);
nand UO_59 (O_59,N_19724,N_19788);
or UO_60 (O_60,N_19683,N_19879);
xnor UO_61 (O_61,N_19395,N_19342);
nand UO_62 (O_62,N_19976,N_19159);
xnor UO_63 (O_63,N_19277,N_19910);
nor UO_64 (O_64,N_19303,N_19590);
or UO_65 (O_65,N_19913,N_19890);
nor UO_66 (O_66,N_19502,N_19720);
or UO_67 (O_67,N_19917,N_19024);
xor UO_68 (O_68,N_19184,N_19236);
nor UO_69 (O_69,N_19942,N_19149);
nand UO_70 (O_70,N_19893,N_19228);
and UO_71 (O_71,N_19922,N_19385);
nor UO_72 (O_72,N_19538,N_19957);
xnor UO_73 (O_73,N_19037,N_19039);
nor UO_74 (O_74,N_19117,N_19908);
nor UO_75 (O_75,N_19169,N_19353);
nand UO_76 (O_76,N_19755,N_19311);
and UO_77 (O_77,N_19462,N_19734);
xnor UO_78 (O_78,N_19646,N_19863);
xor UO_79 (O_79,N_19882,N_19378);
nand UO_80 (O_80,N_19825,N_19512);
and UO_81 (O_81,N_19547,N_19497);
nor UO_82 (O_82,N_19031,N_19434);
nor UO_83 (O_83,N_19644,N_19397);
nand UO_84 (O_84,N_19870,N_19006);
xor UO_85 (O_85,N_19096,N_19529);
and UO_86 (O_86,N_19124,N_19077);
nand UO_87 (O_87,N_19154,N_19460);
or UO_88 (O_88,N_19806,N_19987);
or UO_89 (O_89,N_19361,N_19499);
nor UO_90 (O_90,N_19639,N_19571);
xor UO_91 (O_91,N_19820,N_19828);
nor UO_92 (O_92,N_19412,N_19677);
nand UO_93 (O_93,N_19715,N_19199);
xor UO_94 (O_94,N_19383,N_19607);
nand UO_95 (O_95,N_19405,N_19120);
or UO_96 (O_96,N_19373,N_19443);
or UO_97 (O_97,N_19629,N_19275);
and UO_98 (O_98,N_19307,N_19819);
nand UO_99 (O_99,N_19344,N_19400);
nand UO_100 (O_100,N_19862,N_19986);
and UO_101 (O_101,N_19240,N_19032);
xor UO_102 (O_102,N_19925,N_19094);
nor UO_103 (O_103,N_19132,N_19613);
and UO_104 (O_104,N_19326,N_19622);
or UO_105 (O_105,N_19216,N_19689);
xnor UO_106 (O_106,N_19065,N_19871);
and UO_107 (O_107,N_19531,N_19758);
and UO_108 (O_108,N_19211,N_19824);
or UO_109 (O_109,N_19427,N_19826);
nor UO_110 (O_110,N_19569,N_19359);
and UO_111 (O_111,N_19302,N_19178);
and UO_112 (O_112,N_19973,N_19885);
and UO_113 (O_113,N_19388,N_19367);
xor UO_114 (O_114,N_19221,N_19487);
and UO_115 (O_115,N_19763,N_19197);
or UO_116 (O_116,N_19789,N_19975);
xnor UO_117 (O_117,N_19376,N_19558);
or UO_118 (O_118,N_19935,N_19042);
and UO_119 (O_119,N_19073,N_19717);
nand UO_120 (O_120,N_19815,N_19408);
xor UO_121 (O_121,N_19494,N_19182);
or UO_122 (O_122,N_19348,N_19485);
nand UO_123 (O_123,N_19730,N_19679);
nand UO_124 (O_124,N_19699,N_19288);
nand UO_125 (O_125,N_19340,N_19933);
or UO_126 (O_126,N_19528,N_19540);
nor UO_127 (O_127,N_19778,N_19585);
nand UO_128 (O_128,N_19949,N_19504);
or UO_129 (O_129,N_19560,N_19188);
or UO_130 (O_130,N_19030,N_19035);
and UO_131 (O_131,N_19444,N_19552);
nor UO_132 (O_132,N_19786,N_19190);
and UO_133 (O_133,N_19233,N_19768);
xor UO_134 (O_134,N_19534,N_19386);
or UO_135 (O_135,N_19098,N_19777);
nand UO_136 (O_136,N_19618,N_19329);
or UO_137 (O_137,N_19895,N_19046);
xor UO_138 (O_138,N_19172,N_19511);
nor UO_139 (O_139,N_19290,N_19358);
xor UO_140 (O_140,N_19737,N_19103);
xnor UO_141 (O_141,N_19398,N_19939);
nand UO_142 (O_142,N_19483,N_19245);
nor UO_143 (O_143,N_19174,N_19356);
nand UO_144 (O_144,N_19923,N_19802);
or UO_145 (O_145,N_19924,N_19106);
nor UO_146 (O_146,N_19195,N_19155);
and UO_147 (O_147,N_19714,N_19308);
or UO_148 (O_148,N_19131,N_19581);
xor UO_149 (O_149,N_19433,N_19999);
or UO_150 (O_150,N_19086,N_19387);
or UO_151 (O_151,N_19570,N_19817);
or UO_152 (O_152,N_19294,N_19916);
nor UO_153 (O_153,N_19333,N_19851);
xor UO_154 (O_154,N_19556,N_19330);
and UO_155 (O_155,N_19800,N_19582);
xnor UO_156 (O_156,N_19310,N_19403);
or UO_157 (O_157,N_19074,N_19161);
xor UO_158 (O_158,N_19612,N_19673);
and UO_159 (O_159,N_19357,N_19979);
xor UO_160 (O_160,N_19604,N_19813);
and UO_161 (O_161,N_19193,N_19822);
xnor UO_162 (O_162,N_19316,N_19753);
and UO_163 (O_163,N_19305,N_19598);
xnor UO_164 (O_164,N_19145,N_19391);
xnor UO_165 (O_165,N_19743,N_19765);
xor UO_166 (O_166,N_19919,N_19551);
nor UO_167 (O_167,N_19215,N_19043);
or UO_168 (O_168,N_19418,N_19008);
xor UO_169 (O_169,N_19454,N_19587);
and UO_170 (O_170,N_19869,N_19708);
nand UO_171 (O_171,N_19951,N_19880);
and UO_172 (O_172,N_19067,N_19413);
or UO_173 (O_173,N_19222,N_19262);
and UO_174 (O_174,N_19718,N_19619);
and UO_175 (O_175,N_19889,N_19536);
nand UO_176 (O_176,N_19282,N_19921);
or UO_177 (O_177,N_19790,N_19865);
and UO_178 (O_178,N_19858,N_19142);
and UO_179 (O_179,N_19119,N_19323);
and UO_180 (O_180,N_19393,N_19415);
xor UO_181 (O_181,N_19713,N_19796);
xor UO_182 (O_182,N_19762,N_19772);
xnor UO_183 (O_183,N_19187,N_19722);
or UO_184 (O_184,N_19295,N_19991);
and UO_185 (O_185,N_19165,N_19506);
and UO_186 (O_186,N_19264,N_19500);
nor UO_187 (O_187,N_19621,N_19371);
nor UO_188 (O_188,N_19943,N_19568);
nor UO_189 (O_189,N_19816,N_19445);
nand UO_190 (O_190,N_19230,N_19859);
nand UO_191 (O_191,N_19509,N_19299);
nand UO_192 (O_192,N_19105,N_19204);
nor UO_193 (O_193,N_19967,N_19779);
xnor UO_194 (O_194,N_19104,N_19955);
nand UO_195 (O_195,N_19684,N_19363);
and UO_196 (O_196,N_19602,N_19702);
xor UO_197 (O_197,N_19127,N_19705);
or UO_198 (O_198,N_19244,N_19580);
nand UO_199 (O_199,N_19997,N_19548);
xor UO_200 (O_200,N_19212,N_19953);
xnor UO_201 (O_201,N_19475,N_19798);
nor UO_202 (O_202,N_19080,N_19489);
or UO_203 (O_203,N_19285,N_19420);
nor UO_204 (O_204,N_19108,N_19446);
and UO_205 (O_205,N_19181,N_19896);
or UO_206 (O_206,N_19331,N_19892);
nand UO_207 (O_207,N_19474,N_19505);
and UO_208 (O_208,N_19881,N_19959);
nand UO_209 (O_209,N_19530,N_19467);
xnor UO_210 (O_210,N_19681,N_19716);
xnor UO_211 (O_211,N_19492,N_19998);
nor UO_212 (O_212,N_19234,N_19392);
and UO_213 (O_213,N_19561,N_19107);
nor UO_214 (O_214,N_19081,N_19423);
or UO_215 (O_215,N_19846,N_19891);
xor UO_216 (O_216,N_19557,N_19956);
or UO_217 (O_217,N_19263,N_19832);
xor UO_218 (O_218,N_19599,N_19458);
and UO_219 (O_219,N_19318,N_19033);
xnor UO_220 (O_220,N_19055,N_19872);
xor UO_221 (O_221,N_19225,N_19808);
nor UO_222 (O_222,N_19332,N_19988);
or UO_223 (O_223,N_19665,N_19449);
or UO_224 (O_224,N_19814,N_19572);
and UO_225 (O_225,N_19022,N_19852);
or UO_226 (O_226,N_19671,N_19630);
xnor UO_227 (O_227,N_19384,N_19267);
nand UO_228 (O_228,N_19346,N_19336);
xor UO_229 (O_229,N_19680,N_19615);
nand UO_230 (O_230,N_19928,N_19945);
and UO_231 (O_231,N_19740,N_19821);
nand UO_232 (O_232,N_19775,N_19731);
or UO_233 (O_233,N_19152,N_19586);
nand UO_234 (O_234,N_19206,N_19058);
nand UO_235 (O_235,N_19335,N_19253);
and UO_236 (O_236,N_19709,N_19428);
nand UO_237 (O_237,N_19100,N_19960);
nor UO_238 (O_238,N_19237,N_19805);
xor UO_239 (O_239,N_19057,N_19044);
and UO_240 (O_240,N_19426,N_19324);
and UO_241 (O_241,N_19062,N_19453);
and UO_242 (O_242,N_19214,N_19651);
or UO_243 (O_243,N_19593,N_19457);
xnor UO_244 (O_244,N_19963,N_19001);
xor UO_245 (O_245,N_19517,N_19564);
or UO_246 (O_246,N_19741,N_19934);
xnor UO_247 (O_247,N_19855,N_19799);
nor UO_248 (O_248,N_19915,N_19286);
xnor UO_249 (O_249,N_19579,N_19461);
or UO_250 (O_250,N_19810,N_19856);
and UO_251 (O_251,N_19726,N_19952);
xor UO_252 (O_252,N_19273,N_19012);
and UO_253 (O_253,N_19513,N_19669);
xor UO_254 (O_254,N_19728,N_19970);
nor UO_255 (O_255,N_19902,N_19546);
nor UO_256 (O_256,N_19662,N_19054);
and UO_257 (O_257,N_19250,N_19269);
xnor UO_258 (O_258,N_19047,N_19972);
xnor UO_259 (O_259,N_19173,N_19655);
nor UO_260 (O_260,N_19971,N_19995);
nor UO_261 (O_261,N_19591,N_19706);
and UO_262 (O_262,N_19377,N_19676);
and UO_263 (O_263,N_19157,N_19914);
nor UO_264 (O_264,N_19719,N_19435);
nand UO_265 (O_265,N_19514,N_19803);
nand UO_266 (O_266,N_19906,N_19092);
nand UO_267 (O_267,N_19140,N_19090);
xnor UO_268 (O_268,N_19625,N_19135);
nand UO_269 (O_269,N_19209,N_19113);
nand UO_270 (O_270,N_19577,N_19756);
or UO_271 (O_271,N_19553,N_19455);
or UO_272 (O_272,N_19354,N_19409);
and UO_273 (O_273,N_19381,N_19984);
or UO_274 (O_274,N_19900,N_19725);
and UO_275 (O_275,N_19470,N_19537);
nand UO_276 (O_276,N_19041,N_19432);
nand UO_277 (O_277,N_19627,N_19343);
xor UO_278 (O_278,N_19148,N_19437);
xnor UO_279 (O_279,N_19289,N_19198);
or UO_280 (O_280,N_19147,N_19450);
nor UO_281 (O_281,N_19898,N_19162);
nand UO_282 (O_282,N_19093,N_19831);
xor UO_283 (O_283,N_19766,N_19258);
or UO_284 (O_284,N_19853,N_19251);
nor UO_285 (O_285,N_19017,N_19185);
nor UO_286 (O_286,N_19609,N_19424);
or UO_287 (O_287,N_19224,N_19328);
or UO_288 (O_288,N_19946,N_19659);
or UO_289 (O_289,N_19379,N_19068);
nand UO_290 (O_290,N_19532,N_19501);
nand UO_291 (O_291,N_19056,N_19129);
nand UO_292 (O_292,N_19439,N_19738);
nand UO_293 (O_293,N_19620,N_19770);
nor UO_294 (O_294,N_19518,N_19314);
or UO_295 (O_295,N_19334,N_19578);
nand UO_296 (O_296,N_19747,N_19150);
and UO_297 (O_297,N_19040,N_19369);
nand UO_298 (O_298,N_19927,N_19782);
and UO_299 (O_299,N_19541,N_19141);
nor UO_300 (O_300,N_19301,N_19254);
or UO_301 (O_301,N_19138,N_19797);
xnor UO_302 (O_302,N_19297,N_19566);
or UO_303 (O_303,N_19596,N_19711);
or UO_304 (O_304,N_19259,N_19312);
xnor UO_305 (O_305,N_19648,N_19362);
xor UO_306 (O_306,N_19686,N_19685);
nand UO_307 (O_307,N_19298,N_19126);
xnor UO_308 (O_308,N_19985,N_19887);
and UO_309 (O_309,N_19515,N_19158);
and UO_310 (O_310,N_19075,N_19666);
or UO_311 (O_311,N_19189,N_19525);
or UO_312 (O_312,N_19281,N_19430);
nor UO_313 (O_313,N_19052,N_19868);
nor UO_314 (O_314,N_19735,N_19873);
nand UO_315 (O_315,N_19490,N_19631);
nand UO_316 (O_316,N_19911,N_19495);
xnor UO_317 (O_317,N_19652,N_19079);
xnor UO_318 (O_318,N_19888,N_19769);
or UO_319 (O_319,N_19252,N_19633);
xor UO_320 (O_320,N_19217,N_19441);
or UO_321 (O_321,N_19524,N_19573);
and UO_322 (O_322,N_19347,N_19143);
nor UO_323 (O_323,N_19516,N_19904);
nand UO_324 (O_324,N_19700,N_19232);
nand UO_325 (O_325,N_19678,N_19051);
nor UO_326 (O_326,N_19635,N_19300);
and UO_327 (O_327,N_19761,N_19306);
nand UO_328 (O_328,N_19076,N_19482);
xor UO_329 (O_329,N_19647,N_19151);
nand UO_330 (O_330,N_19208,N_19085);
nand UO_331 (O_331,N_19000,N_19406);
and UO_332 (O_332,N_19018,N_19614);
nor UO_333 (O_333,N_19941,N_19144);
xnor UO_334 (O_334,N_19156,N_19070);
xor UO_335 (O_335,N_19095,N_19729);
xnor UO_336 (O_336,N_19750,N_19429);
and UO_337 (O_337,N_19674,N_19279);
nand UO_338 (O_338,N_19038,N_19550);
or UO_339 (O_339,N_19014,N_19227);
or UO_340 (O_340,N_19239,N_19034);
and UO_341 (O_341,N_19710,N_19349);
nand UO_342 (O_342,N_19603,N_19595);
nand UO_343 (O_343,N_19472,N_19164);
and UO_344 (O_344,N_19050,N_19136);
or UO_345 (O_345,N_19533,N_19059);
and UO_346 (O_346,N_19002,N_19121);
nand UO_347 (O_347,N_19200,N_19833);
nand UO_348 (O_348,N_19261,N_19543);
or UO_349 (O_349,N_19909,N_19304);
or UO_350 (O_350,N_19442,N_19139);
nor UO_351 (O_351,N_19701,N_19624);
or UO_352 (O_352,N_19886,N_19257);
nor UO_353 (O_353,N_19431,N_19372);
and UO_354 (O_354,N_19527,N_19407);
or UO_355 (O_355,N_19565,N_19843);
xor UO_356 (O_356,N_19175,N_19226);
and UO_357 (O_357,N_19545,N_19088);
xnor UO_358 (O_358,N_19045,N_19876);
xnor UO_359 (O_359,N_19791,N_19759);
or UO_360 (O_360,N_19220,N_19690);
and UO_361 (O_361,N_19694,N_19703);
nand UO_362 (O_362,N_19559,N_19594);
xnor UO_363 (O_363,N_19848,N_19823);
or UO_364 (O_364,N_19177,N_19661);
or UO_365 (O_365,N_19576,N_19122);
nand UO_366 (O_366,N_19337,N_19696);
or UO_367 (O_367,N_19962,N_19510);
xor UO_368 (O_368,N_19801,N_19486);
nand UO_369 (O_369,N_19268,N_19994);
or UO_370 (O_370,N_19072,N_19938);
nor UO_371 (O_371,N_19421,N_19542);
nor UO_372 (O_372,N_19688,N_19597);
or UO_373 (O_373,N_19194,N_19663);
and UO_374 (O_374,N_19180,N_19114);
nand UO_375 (O_375,N_19087,N_19355);
nand UO_376 (O_376,N_19732,N_19535);
and UO_377 (O_377,N_19083,N_19950);
xnor UO_378 (O_378,N_19498,N_19698);
nor UO_379 (O_379,N_19751,N_19968);
nor UO_380 (O_380,N_19066,N_19857);
nor UO_381 (O_381,N_19969,N_19471);
nand UO_382 (O_382,N_19125,N_19283);
xnor UO_383 (O_383,N_19176,N_19748);
or UO_384 (O_384,N_19010,N_19866);
or UO_385 (O_385,N_19964,N_19274);
and UO_386 (O_386,N_19744,N_19742);
or UO_387 (O_387,N_19401,N_19327);
xor UO_388 (O_388,N_19091,N_19563);
nor UO_389 (O_389,N_19667,N_19672);
and UO_390 (O_390,N_19656,N_19452);
xor UO_391 (O_391,N_19463,N_19201);
and UO_392 (O_392,N_19654,N_19937);
xor UO_393 (O_393,N_19918,N_19013);
nor UO_394 (O_394,N_19203,N_19642);
or UO_395 (O_395,N_19958,N_19668);
or UO_396 (O_396,N_19807,N_19606);
or UO_397 (O_397,N_19670,N_19118);
nor UO_398 (O_398,N_19520,N_19912);
nand UO_399 (O_399,N_19456,N_19345);
or UO_400 (O_400,N_19278,N_19477);
nor UO_401 (O_401,N_19110,N_19171);
and UO_402 (O_402,N_19476,N_19523);
or UO_403 (O_403,N_19322,N_19374);
nand UO_404 (O_404,N_19980,N_19867);
and UO_405 (O_405,N_19754,N_19990);
nor UO_406 (O_406,N_19522,N_19026);
or UO_407 (O_407,N_19926,N_19812);
and UO_408 (O_408,N_19589,N_19894);
or UO_409 (O_409,N_19425,N_19692);
xnor UO_410 (O_410,N_19601,N_19265);
and UO_411 (O_411,N_19339,N_19168);
and UO_412 (O_412,N_19844,N_19309);
xnor UO_413 (O_413,N_19982,N_19745);
nor UO_414 (O_414,N_19794,N_19218);
xnor UO_415 (O_415,N_19811,N_19827);
or UO_416 (O_416,N_19658,N_19899);
nor UO_417 (O_417,N_19183,N_19712);
and UO_418 (O_418,N_19167,N_19883);
nor UO_419 (O_419,N_19864,N_19840);
and UO_420 (O_420,N_19978,N_19023);
nor UO_421 (O_421,N_19519,N_19293);
or UO_422 (O_422,N_19929,N_19757);
nor UO_423 (O_423,N_19649,N_19160);
and UO_424 (O_424,N_19451,N_19238);
xor UO_425 (O_425,N_19640,N_19019);
nand UO_426 (O_426,N_19246,N_19207);
nand UO_427 (O_427,N_19260,N_19901);
or UO_428 (O_428,N_19526,N_19249);
and UO_429 (O_429,N_19321,N_19130);
nand UO_430 (O_430,N_19025,N_19473);
xnor UO_431 (O_431,N_19166,N_19776);
nand UO_432 (O_432,N_19317,N_19370);
nor UO_433 (O_433,N_19480,N_19111);
or UO_434 (O_434,N_19760,N_19027);
and UO_435 (O_435,N_19785,N_19693);
nand UO_436 (O_436,N_19366,N_19396);
and UO_437 (O_437,N_19723,N_19605);
or UO_438 (O_438,N_19687,N_19727);
or UO_439 (O_439,N_19319,N_19229);
or UO_440 (O_440,N_19781,N_19069);
or UO_441 (O_441,N_19653,N_19481);
and UO_442 (O_442,N_19977,N_19410);
or UO_443 (O_443,N_19733,N_19368);
xor UO_444 (O_444,N_19422,N_19641);
and UO_445 (O_445,N_19296,N_19746);
xor UO_446 (O_446,N_19170,N_19944);
and UO_447 (O_447,N_19116,N_19884);
nor UO_448 (O_448,N_19503,N_19459);
xor UO_449 (O_449,N_19847,N_19053);
or UO_450 (O_450,N_19829,N_19736);
and UO_451 (O_451,N_19479,N_19841);
nand UO_452 (O_452,N_19325,N_19049);
nand UO_453 (O_453,N_19276,N_19256);
xor UO_454 (O_454,N_19484,N_19616);
or UO_455 (O_455,N_19191,N_19436);
xor UO_456 (O_456,N_19202,N_19466);
and UO_457 (O_457,N_19875,N_19993);
and UO_458 (O_458,N_19099,N_19657);
and UO_459 (O_459,N_19440,N_19608);
and UO_460 (O_460,N_19780,N_19123);
and UO_461 (O_461,N_19562,N_19016);
nor UO_462 (O_462,N_19932,N_19247);
nor UO_463 (O_463,N_19133,N_19205);
nor UO_464 (O_464,N_19447,N_19048);
nand UO_465 (O_465,N_19931,N_19749);
nand UO_466 (O_466,N_19496,N_19842);
and UO_467 (O_467,N_19583,N_19271);
or UO_468 (O_468,N_19137,N_19231);
nand UO_469 (O_469,N_19007,N_19554);
xor UO_470 (O_470,N_19417,N_19102);
and UO_471 (O_471,N_19488,N_19241);
or UO_472 (O_472,N_19468,N_19380);
or UO_473 (O_473,N_19835,N_19818);
and UO_474 (O_474,N_19637,N_19134);
nand UO_475 (O_475,N_19004,N_19836);
nor UO_476 (O_476,N_19280,N_19783);
and UO_477 (O_477,N_19036,N_19078);
nor UO_478 (O_478,N_19874,N_19097);
nand UO_479 (O_479,N_19089,N_19021);
nor UO_480 (O_480,N_19084,N_19438);
nand UO_481 (O_481,N_19192,N_19771);
xor UO_482 (O_482,N_19029,N_19809);
xor UO_483 (O_483,N_19623,N_19920);
or UO_484 (O_484,N_19574,N_19411);
xnor UO_485 (O_485,N_19555,N_19860);
or UO_486 (O_486,N_19966,N_19905);
or UO_487 (O_487,N_19146,N_19404);
nor UO_488 (O_488,N_19414,N_19930);
or UO_489 (O_489,N_19575,N_19015);
nand UO_490 (O_490,N_19284,N_19064);
xor UO_491 (O_491,N_19243,N_19365);
xor UO_492 (O_492,N_19364,N_19508);
xnor UO_493 (O_493,N_19419,N_19849);
nor UO_494 (O_494,N_19020,N_19974);
xor UO_495 (O_495,N_19082,N_19270);
and UO_496 (O_496,N_19632,N_19638);
nand UO_497 (O_497,N_19643,N_19784);
and UO_498 (O_498,N_19402,N_19697);
or UO_499 (O_499,N_19838,N_19996);
and UO_500 (O_500,N_19318,N_19960);
xor UO_501 (O_501,N_19294,N_19361);
nand UO_502 (O_502,N_19760,N_19997);
nor UO_503 (O_503,N_19529,N_19179);
xnor UO_504 (O_504,N_19774,N_19497);
and UO_505 (O_505,N_19048,N_19562);
nand UO_506 (O_506,N_19761,N_19236);
nand UO_507 (O_507,N_19853,N_19922);
xnor UO_508 (O_508,N_19261,N_19041);
nor UO_509 (O_509,N_19069,N_19578);
or UO_510 (O_510,N_19985,N_19067);
and UO_511 (O_511,N_19646,N_19120);
nor UO_512 (O_512,N_19168,N_19312);
xnor UO_513 (O_513,N_19417,N_19032);
xnor UO_514 (O_514,N_19542,N_19056);
nand UO_515 (O_515,N_19550,N_19492);
or UO_516 (O_516,N_19973,N_19745);
nand UO_517 (O_517,N_19109,N_19608);
nor UO_518 (O_518,N_19599,N_19766);
and UO_519 (O_519,N_19793,N_19904);
nor UO_520 (O_520,N_19477,N_19205);
nand UO_521 (O_521,N_19183,N_19224);
xnor UO_522 (O_522,N_19221,N_19007);
nand UO_523 (O_523,N_19448,N_19339);
nand UO_524 (O_524,N_19793,N_19526);
xor UO_525 (O_525,N_19830,N_19147);
xnor UO_526 (O_526,N_19837,N_19209);
and UO_527 (O_527,N_19534,N_19265);
and UO_528 (O_528,N_19027,N_19211);
and UO_529 (O_529,N_19623,N_19726);
nand UO_530 (O_530,N_19945,N_19245);
nand UO_531 (O_531,N_19960,N_19273);
and UO_532 (O_532,N_19447,N_19257);
xnor UO_533 (O_533,N_19077,N_19751);
nor UO_534 (O_534,N_19469,N_19286);
nor UO_535 (O_535,N_19997,N_19288);
nand UO_536 (O_536,N_19427,N_19499);
xnor UO_537 (O_537,N_19746,N_19220);
nor UO_538 (O_538,N_19194,N_19304);
and UO_539 (O_539,N_19171,N_19147);
or UO_540 (O_540,N_19898,N_19682);
nor UO_541 (O_541,N_19764,N_19650);
or UO_542 (O_542,N_19155,N_19747);
nand UO_543 (O_543,N_19271,N_19407);
nand UO_544 (O_544,N_19677,N_19328);
nand UO_545 (O_545,N_19166,N_19079);
nand UO_546 (O_546,N_19943,N_19165);
or UO_547 (O_547,N_19410,N_19020);
nand UO_548 (O_548,N_19474,N_19889);
and UO_549 (O_549,N_19982,N_19552);
nand UO_550 (O_550,N_19533,N_19080);
or UO_551 (O_551,N_19080,N_19571);
nor UO_552 (O_552,N_19650,N_19200);
and UO_553 (O_553,N_19149,N_19422);
and UO_554 (O_554,N_19706,N_19758);
nor UO_555 (O_555,N_19488,N_19244);
nand UO_556 (O_556,N_19985,N_19597);
or UO_557 (O_557,N_19855,N_19615);
nor UO_558 (O_558,N_19114,N_19727);
and UO_559 (O_559,N_19653,N_19622);
nor UO_560 (O_560,N_19439,N_19052);
or UO_561 (O_561,N_19667,N_19968);
nand UO_562 (O_562,N_19141,N_19319);
nor UO_563 (O_563,N_19016,N_19170);
and UO_564 (O_564,N_19908,N_19842);
nor UO_565 (O_565,N_19843,N_19194);
xor UO_566 (O_566,N_19839,N_19093);
nor UO_567 (O_567,N_19239,N_19662);
nand UO_568 (O_568,N_19291,N_19610);
and UO_569 (O_569,N_19106,N_19657);
xor UO_570 (O_570,N_19821,N_19157);
nand UO_571 (O_571,N_19317,N_19668);
nand UO_572 (O_572,N_19609,N_19245);
nor UO_573 (O_573,N_19339,N_19184);
nor UO_574 (O_574,N_19287,N_19292);
nand UO_575 (O_575,N_19309,N_19653);
xnor UO_576 (O_576,N_19067,N_19507);
xnor UO_577 (O_577,N_19255,N_19412);
or UO_578 (O_578,N_19096,N_19213);
nor UO_579 (O_579,N_19076,N_19605);
nor UO_580 (O_580,N_19264,N_19584);
xnor UO_581 (O_581,N_19329,N_19085);
xor UO_582 (O_582,N_19296,N_19859);
or UO_583 (O_583,N_19238,N_19336);
or UO_584 (O_584,N_19064,N_19594);
nor UO_585 (O_585,N_19748,N_19895);
and UO_586 (O_586,N_19063,N_19010);
nand UO_587 (O_587,N_19765,N_19320);
nand UO_588 (O_588,N_19421,N_19019);
and UO_589 (O_589,N_19250,N_19272);
or UO_590 (O_590,N_19511,N_19685);
or UO_591 (O_591,N_19326,N_19747);
and UO_592 (O_592,N_19265,N_19033);
or UO_593 (O_593,N_19740,N_19015);
and UO_594 (O_594,N_19516,N_19641);
or UO_595 (O_595,N_19012,N_19053);
or UO_596 (O_596,N_19765,N_19051);
and UO_597 (O_597,N_19262,N_19116);
nor UO_598 (O_598,N_19438,N_19582);
or UO_599 (O_599,N_19956,N_19031);
and UO_600 (O_600,N_19774,N_19071);
nand UO_601 (O_601,N_19109,N_19367);
nand UO_602 (O_602,N_19242,N_19881);
nand UO_603 (O_603,N_19283,N_19102);
nor UO_604 (O_604,N_19204,N_19669);
and UO_605 (O_605,N_19963,N_19800);
or UO_606 (O_606,N_19988,N_19697);
and UO_607 (O_607,N_19148,N_19215);
xor UO_608 (O_608,N_19836,N_19192);
or UO_609 (O_609,N_19653,N_19820);
nand UO_610 (O_610,N_19786,N_19573);
nor UO_611 (O_611,N_19532,N_19485);
xor UO_612 (O_612,N_19558,N_19345);
xnor UO_613 (O_613,N_19617,N_19978);
nor UO_614 (O_614,N_19581,N_19510);
and UO_615 (O_615,N_19323,N_19684);
or UO_616 (O_616,N_19464,N_19193);
nor UO_617 (O_617,N_19488,N_19534);
xnor UO_618 (O_618,N_19262,N_19134);
nor UO_619 (O_619,N_19212,N_19640);
or UO_620 (O_620,N_19051,N_19719);
or UO_621 (O_621,N_19013,N_19255);
or UO_622 (O_622,N_19108,N_19293);
xor UO_623 (O_623,N_19952,N_19614);
or UO_624 (O_624,N_19465,N_19642);
nor UO_625 (O_625,N_19717,N_19838);
xnor UO_626 (O_626,N_19965,N_19566);
or UO_627 (O_627,N_19152,N_19992);
nor UO_628 (O_628,N_19679,N_19368);
and UO_629 (O_629,N_19584,N_19259);
and UO_630 (O_630,N_19557,N_19766);
and UO_631 (O_631,N_19425,N_19637);
and UO_632 (O_632,N_19223,N_19406);
nand UO_633 (O_633,N_19166,N_19467);
nor UO_634 (O_634,N_19434,N_19390);
xnor UO_635 (O_635,N_19115,N_19952);
nand UO_636 (O_636,N_19394,N_19542);
xnor UO_637 (O_637,N_19830,N_19242);
xnor UO_638 (O_638,N_19245,N_19824);
and UO_639 (O_639,N_19190,N_19747);
and UO_640 (O_640,N_19146,N_19871);
xor UO_641 (O_641,N_19638,N_19125);
or UO_642 (O_642,N_19352,N_19427);
and UO_643 (O_643,N_19256,N_19746);
and UO_644 (O_644,N_19080,N_19274);
nand UO_645 (O_645,N_19575,N_19475);
nor UO_646 (O_646,N_19546,N_19269);
xnor UO_647 (O_647,N_19755,N_19176);
nor UO_648 (O_648,N_19028,N_19146);
nand UO_649 (O_649,N_19742,N_19392);
xnor UO_650 (O_650,N_19365,N_19457);
nand UO_651 (O_651,N_19766,N_19804);
nor UO_652 (O_652,N_19241,N_19922);
or UO_653 (O_653,N_19341,N_19236);
nor UO_654 (O_654,N_19347,N_19536);
xnor UO_655 (O_655,N_19374,N_19201);
nand UO_656 (O_656,N_19378,N_19500);
nor UO_657 (O_657,N_19128,N_19229);
or UO_658 (O_658,N_19228,N_19216);
or UO_659 (O_659,N_19567,N_19231);
nand UO_660 (O_660,N_19469,N_19148);
nand UO_661 (O_661,N_19377,N_19168);
or UO_662 (O_662,N_19951,N_19080);
nor UO_663 (O_663,N_19371,N_19519);
and UO_664 (O_664,N_19874,N_19064);
and UO_665 (O_665,N_19537,N_19987);
nand UO_666 (O_666,N_19603,N_19888);
nand UO_667 (O_667,N_19388,N_19121);
nor UO_668 (O_668,N_19365,N_19054);
nor UO_669 (O_669,N_19138,N_19839);
nor UO_670 (O_670,N_19595,N_19648);
nand UO_671 (O_671,N_19586,N_19657);
and UO_672 (O_672,N_19576,N_19526);
and UO_673 (O_673,N_19909,N_19067);
and UO_674 (O_674,N_19315,N_19711);
or UO_675 (O_675,N_19658,N_19247);
nand UO_676 (O_676,N_19039,N_19626);
and UO_677 (O_677,N_19686,N_19103);
nand UO_678 (O_678,N_19424,N_19721);
and UO_679 (O_679,N_19178,N_19843);
xor UO_680 (O_680,N_19175,N_19506);
or UO_681 (O_681,N_19219,N_19806);
and UO_682 (O_682,N_19087,N_19648);
and UO_683 (O_683,N_19662,N_19670);
nand UO_684 (O_684,N_19653,N_19114);
xnor UO_685 (O_685,N_19243,N_19466);
nor UO_686 (O_686,N_19654,N_19341);
nor UO_687 (O_687,N_19969,N_19754);
or UO_688 (O_688,N_19596,N_19193);
xnor UO_689 (O_689,N_19635,N_19773);
nor UO_690 (O_690,N_19061,N_19722);
or UO_691 (O_691,N_19324,N_19658);
and UO_692 (O_692,N_19480,N_19627);
nand UO_693 (O_693,N_19336,N_19504);
xnor UO_694 (O_694,N_19802,N_19591);
nor UO_695 (O_695,N_19536,N_19734);
xnor UO_696 (O_696,N_19046,N_19901);
or UO_697 (O_697,N_19200,N_19749);
or UO_698 (O_698,N_19023,N_19555);
nor UO_699 (O_699,N_19472,N_19911);
nand UO_700 (O_700,N_19791,N_19062);
nor UO_701 (O_701,N_19629,N_19099);
nor UO_702 (O_702,N_19233,N_19517);
xor UO_703 (O_703,N_19211,N_19790);
nand UO_704 (O_704,N_19545,N_19252);
nor UO_705 (O_705,N_19397,N_19595);
or UO_706 (O_706,N_19057,N_19622);
nand UO_707 (O_707,N_19709,N_19770);
and UO_708 (O_708,N_19849,N_19123);
nor UO_709 (O_709,N_19144,N_19603);
xor UO_710 (O_710,N_19528,N_19925);
nand UO_711 (O_711,N_19799,N_19808);
and UO_712 (O_712,N_19255,N_19669);
or UO_713 (O_713,N_19610,N_19214);
nand UO_714 (O_714,N_19928,N_19176);
nand UO_715 (O_715,N_19223,N_19001);
nor UO_716 (O_716,N_19716,N_19139);
or UO_717 (O_717,N_19195,N_19609);
nand UO_718 (O_718,N_19590,N_19308);
or UO_719 (O_719,N_19169,N_19438);
nand UO_720 (O_720,N_19258,N_19423);
xnor UO_721 (O_721,N_19647,N_19535);
or UO_722 (O_722,N_19938,N_19376);
nand UO_723 (O_723,N_19901,N_19209);
nor UO_724 (O_724,N_19920,N_19816);
xnor UO_725 (O_725,N_19717,N_19152);
nand UO_726 (O_726,N_19841,N_19051);
xnor UO_727 (O_727,N_19496,N_19646);
nor UO_728 (O_728,N_19705,N_19559);
xnor UO_729 (O_729,N_19420,N_19990);
or UO_730 (O_730,N_19917,N_19452);
nand UO_731 (O_731,N_19624,N_19748);
xnor UO_732 (O_732,N_19343,N_19300);
and UO_733 (O_733,N_19956,N_19508);
nor UO_734 (O_734,N_19338,N_19818);
xor UO_735 (O_735,N_19840,N_19297);
and UO_736 (O_736,N_19372,N_19877);
or UO_737 (O_737,N_19755,N_19518);
nor UO_738 (O_738,N_19584,N_19738);
and UO_739 (O_739,N_19709,N_19324);
or UO_740 (O_740,N_19162,N_19358);
xor UO_741 (O_741,N_19974,N_19154);
or UO_742 (O_742,N_19329,N_19128);
nand UO_743 (O_743,N_19505,N_19160);
xor UO_744 (O_744,N_19518,N_19156);
or UO_745 (O_745,N_19754,N_19109);
and UO_746 (O_746,N_19797,N_19358);
nand UO_747 (O_747,N_19370,N_19820);
xor UO_748 (O_748,N_19326,N_19062);
or UO_749 (O_749,N_19612,N_19254);
nand UO_750 (O_750,N_19690,N_19039);
nor UO_751 (O_751,N_19701,N_19241);
xnor UO_752 (O_752,N_19637,N_19837);
nor UO_753 (O_753,N_19195,N_19153);
or UO_754 (O_754,N_19957,N_19143);
nor UO_755 (O_755,N_19031,N_19675);
nand UO_756 (O_756,N_19269,N_19761);
xor UO_757 (O_757,N_19822,N_19511);
or UO_758 (O_758,N_19373,N_19608);
xnor UO_759 (O_759,N_19291,N_19176);
nor UO_760 (O_760,N_19231,N_19685);
or UO_761 (O_761,N_19582,N_19556);
or UO_762 (O_762,N_19953,N_19121);
nand UO_763 (O_763,N_19863,N_19629);
or UO_764 (O_764,N_19274,N_19810);
and UO_765 (O_765,N_19904,N_19827);
and UO_766 (O_766,N_19471,N_19178);
nor UO_767 (O_767,N_19174,N_19344);
or UO_768 (O_768,N_19136,N_19283);
or UO_769 (O_769,N_19861,N_19262);
and UO_770 (O_770,N_19348,N_19268);
or UO_771 (O_771,N_19884,N_19861);
nand UO_772 (O_772,N_19414,N_19030);
and UO_773 (O_773,N_19278,N_19168);
nand UO_774 (O_774,N_19605,N_19130);
and UO_775 (O_775,N_19788,N_19174);
xor UO_776 (O_776,N_19272,N_19305);
and UO_777 (O_777,N_19592,N_19349);
and UO_778 (O_778,N_19993,N_19975);
nand UO_779 (O_779,N_19761,N_19686);
or UO_780 (O_780,N_19018,N_19392);
nand UO_781 (O_781,N_19903,N_19026);
nor UO_782 (O_782,N_19748,N_19884);
xnor UO_783 (O_783,N_19121,N_19484);
or UO_784 (O_784,N_19192,N_19991);
xor UO_785 (O_785,N_19456,N_19750);
or UO_786 (O_786,N_19172,N_19845);
and UO_787 (O_787,N_19167,N_19607);
nor UO_788 (O_788,N_19027,N_19615);
or UO_789 (O_789,N_19995,N_19117);
and UO_790 (O_790,N_19700,N_19246);
nand UO_791 (O_791,N_19296,N_19562);
and UO_792 (O_792,N_19181,N_19704);
xor UO_793 (O_793,N_19364,N_19525);
xor UO_794 (O_794,N_19194,N_19594);
and UO_795 (O_795,N_19589,N_19372);
xor UO_796 (O_796,N_19899,N_19342);
nand UO_797 (O_797,N_19746,N_19684);
xor UO_798 (O_798,N_19809,N_19749);
and UO_799 (O_799,N_19061,N_19519);
and UO_800 (O_800,N_19323,N_19108);
nand UO_801 (O_801,N_19589,N_19242);
nor UO_802 (O_802,N_19969,N_19323);
nor UO_803 (O_803,N_19235,N_19184);
xnor UO_804 (O_804,N_19157,N_19751);
nor UO_805 (O_805,N_19875,N_19497);
nand UO_806 (O_806,N_19776,N_19035);
or UO_807 (O_807,N_19740,N_19911);
and UO_808 (O_808,N_19603,N_19953);
and UO_809 (O_809,N_19748,N_19892);
nand UO_810 (O_810,N_19412,N_19596);
or UO_811 (O_811,N_19067,N_19351);
nand UO_812 (O_812,N_19482,N_19293);
nand UO_813 (O_813,N_19885,N_19704);
nor UO_814 (O_814,N_19025,N_19095);
and UO_815 (O_815,N_19198,N_19321);
and UO_816 (O_816,N_19420,N_19421);
or UO_817 (O_817,N_19747,N_19096);
or UO_818 (O_818,N_19323,N_19345);
nor UO_819 (O_819,N_19733,N_19110);
xor UO_820 (O_820,N_19021,N_19065);
or UO_821 (O_821,N_19228,N_19284);
nor UO_822 (O_822,N_19112,N_19309);
nor UO_823 (O_823,N_19088,N_19175);
or UO_824 (O_824,N_19778,N_19244);
nand UO_825 (O_825,N_19775,N_19800);
xor UO_826 (O_826,N_19336,N_19965);
or UO_827 (O_827,N_19236,N_19855);
or UO_828 (O_828,N_19672,N_19253);
or UO_829 (O_829,N_19340,N_19846);
nor UO_830 (O_830,N_19455,N_19040);
nand UO_831 (O_831,N_19827,N_19791);
nor UO_832 (O_832,N_19276,N_19832);
nor UO_833 (O_833,N_19564,N_19401);
and UO_834 (O_834,N_19692,N_19725);
xnor UO_835 (O_835,N_19008,N_19798);
or UO_836 (O_836,N_19626,N_19593);
and UO_837 (O_837,N_19624,N_19725);
nand UO_838 (O_838,N_19677,N_19712);
or UO_839 (O_839,N_19576,N_19278);
or UO_840 (O_840,N_19124,N_19868);
nand UO_841 (O_841,N_19453,N_19905);
and UO_842 (O_842,N_19963,N_19873);
nand UO_843 (O_843,N_19590,N_19989);
nand UO_844 (O_844,N_19326,N_19577);
and UO_845 (O_845,N_19181,N_19691);
or UO_846 (O_846,N_19531,N_19558);
or UO_847 (O_847,N_19414,N_19671);
nand UO_848 (O_848,N_19421,N_19135);
or UO_849 (O_849,N_19948,N_19557);
nor UO_850 (O_850,N_19486,N_19595);
nor UO_851 (O_851,N_19743,N_19938);
nor UO_852 (O_852,N_19358,N_19932);
or UO_853 (O_853,N_19254,N_19074);
or UO_854 (O_854,N_19192,N_19731);
or UO_855 (O_855,N_19606,N_19861);
nor UO_856 (O_856,N_19605,N_19814);
xor UO_857 (O_857,N_19999,N_19373);
nand UO_858 (O_858,N_19189,N_19721);
nor UO_859 (O_859,N_19421,N_19313);
xnor UO_860 (O_860,N_19253,N_19759);
or UO_861 (O_861,N_19199,N_19003);
or UO_862 (O_862,N_19741,N_19254);
nand UO_863 (O_863,N_19492,N_19425);
or UO_864 (O_864,N_19319,N_19323);
xnor UO_865 (O_865,N_19752,N_19821);
or UO_866 (O_866,N_19562,N_19675);
xnor UO_867 (O_867,N_19068,N_19512);
nor UO_868 (O_868,N_19703,N_19409);
and UO_869 (O_869,N_19826,N_19515);
or UO_870 (O_870,N_19143,N_19377);
and UO_871 (O_871,N_19597,N_19418);
or UO_872 (O_872,N_19080,N_19733);
or UO_873 (O_873,N_19807,N_19785);
xor UO_874 (O_874,N_19178,N_19152);
nor UO_875 (O_875,N_19274,N_19429);
and UO_876 (O_876,N_19760,N_19455);
nor UO_877 (O_877,N_19556,N_19376);
or UO_878 (O_878,N_19685,N_19727);
xnor UO_879 (O_879,N_19234,N_19748);
or UO_880 (O_880,N_19778,N_19735);
nand UO_881 (O_881,N_19841,N_19862);
xor UO_882 (O_882,N_19346,N_19253);
nor UO_883 (O_883,N_19577,N_19054);
nor UO_884 (O_884,N_19962,N_19379);
nand UO_885 (O_885,N_19608,N_19691);
and UO_886 (O_886,N_19452,N_19727);
or UO_887 (O_887,N_19343,N_19050);
and UO_888 (O_888,N_19324,N_19106);
xor UO_889 (O_889,N_19489,N_19862);
nand UO_890 (O_890,N_19904,N_19881);
xnor UO_891 (O_891,N_19302,N_19806);
nand UO_892 (O_892,N_19245,N_19369);
nand UO_893 (O_893,N_19678,N_19273);
or UO_894 (O_894,N_19674,N_19986);
xor UO_895 (O_895,N_19722,N_19341);
nand UO_896 (O_896,N_19282,N_19995);
nand UO_897 (O_897,N_19519,N_19978);
or UO_898 (O_898,N_19243,N_19359);
nor UO_899 (O_899,N_19856,N_19013);
xnor UO_900 (O_900,N_19373,N_19929);
nand UO_901 (O_901,N_19075,N_19620);
or UO_902 (O_902,N_19595,N_19107);
and UO_903 (O_903,N_19953,N_19660);
nand UO_904 (O_904,N_19359,N_19539);
nand UO_905 (O_905,N_19651,N_19955);
nor UO_906 (O_906,N_19395,N_19603);
nand UO_907 (O_907,N_19944,N_19540);
nand UO_908 (O_908,N_19836,N_19403);
or UO_909 (O_909,N_19065,N_19414);
nand UO_910 (O_910,N_19918,N_19246);
or UO_911 (O_911,N_19325,N_19623);
and UO_912 (O_912,N_19255,N_19672);
or UO_913 (O_913,N_19675,N_19278);
and UO_914 (O_914,N_19062,N_19999);
and UO_915 (O_915,N_19574,N_19168);
xnor UO_916 (O_916,N_19970,N_19232);
or UO_917 (O_917,N_19279,N_19478);
nor UO_918 (O_918,N_19189,N_19002);
xor UO_919 (O_919,N_19100,N_19039);
and UO_920 (O_920,N_19591,N_19007);
nor UO_921 (O_921,N_19749,N_19170);
or UO_922 (O_922,N_19610,N_19222);
or UO_923 (O_923,N_19743,N_19533);
or UO_924 (O_924,N_19420,N_19401);
nor UO_925 (O_925,N_19960,N_19478);
or UO_926 (O_926,N_19478,N_19401);
and UO_927 (O_927,N_19345,N_19980);
nor UO_928 (O_928,N_19375,N_19021);
nor UO_929 (O_929,N_19415,N_19352);
xor UO_930 (O_930,N_19686,N_19428);
and UO_931 (O_931,N_19975,N_19871);
or UO_932 (O_932,N_19100,N_19105);
nand UO_933 (O_933,N_19906,N_19596);
or UO_934 (O_934,N_19448,N_19516);
nand UO_935 (O_935,N_19282,N_19360);
nand UO_936 (O_936,N_19900,N_19586);
xnor UO_937 (O_937,N_19855,N_19569);
and UO_938 (O_938,N_19351,N_19429);
nor UO_939 (O_939,N_19021,N_19976);
xor UO_940 (O_940,N_19375,N_19942);
and UO_941 (O_941,N_19992,N_19702);
nor UO_942 (O_942,N_19477,N_19755);
nand UO_943 (O_943,N_19146,N_19055);
nand UO_944 (O_944,N_19414,N_19800);
nand UO_945 (O_945,N_19654,N_19886);
xor UO_946 (O_946,N_19002,N_19386);
nor UO_947 (O_947,N_19328,N_19201);
nand UO_948 (O_948,N_19372,N_19709);
or UO_949 (O_949,N_19148,N_19514);
nand UO_950 (O_950,N_19424,N_19493);
nor UO_951 (O_951,N_19811,N_19209);
nand UO_952 (O_952,N_19542,N_19575);
nand UO_953 (O_953,N_19329,N_19523);
and UO_954 (O_954,N_19894,N_19612);
or UO_955 (O_955,N_19988,N_19018);
and UO_956 (O_956,N_19064,N_19516);
nand UO_957 (O_957,N_19711,N_19926);
nor UO_958 (O_958,N_19197,N_19395);
xor UO_959 (O_959,N_19447,N_19410);
nand UO_960 (O_960,N_19117,N_19716);
or UO_961 (O_961,N_19695,N_19570);
and UO_962 (O_962,N_19865,N_19397);
nand UO_963 (O_963,N_19556,N_19149);
nand UO_964 (O_964,N_19807,N_19690);
nand UO_965 (O_965,N_19299,N_19843);
xnor UO_966 (O_966,N_19882,N_19202);
or UO_967 (O_967,N_19687,N_19203);
xor UO_968 (O_968,N_19280,N_19126);
nand UO_969 (O_969,N_19352,N_19542);
and UO_970 (O_970,N_19350,N_19156);
nor UO_971 (O_971,N_19999,N_19882);
nor UO_972 (O_972,N_19765,N_19340);
nand UO_973 (O_973,N_19279,N_19460);
or UO_974 (O_974,N_19814,N_19201);
nor UO_975 (O_975,N_19504,N_19071);
nand UO_976 (O_976,N_19945,N_19544);
or UO_977 (O_977,N_19176,N_19219);
nand UO_978 (O_978,N_19337,N_19898);
and UO_979 (O_979,N_19032,N_19179);
nand UO_980 (O_980,N_19337,N_19042);
nor UO_981 (O_981,N_19539,N_19969);
and UO_982 (O_982,N_19782,N_19017);
nor UO_983 (O_983,N_19997,N_19903);
nor UO_984 (O_984,N_19202,N_19400);
and UO_985 (O_985,N_19848,N_19078);
and UO_986 (O_986,N_19291,N_19923);
or UO_987 (O_987,N_19096,N_19404);
nor UO_988 (O_988,N_19645,N_19221);
and UO_989 (O_989,N_19197,N_19496);
and UO_990 (O_990,N_19871,N_19286);
nor UO_991 (O_991,N_19426,N_19842);
and UO_992 (O_992,N_19763,N_19683);
and UO_993 (O_993,N_19020,N_19879);
xnor UO_994 (O_994,N_19845,N_19400);
xor UO_995 (O_995,N_19044,N_19720);
or UO_996 (O_996,N_19785,N_19774);
xnor UO_997 (O_997,N_19510,N_19842);
xnor UO_998 (O_998,N_19886,N_19214);
or UO_999 (O_999,N_19937,N_19724);
nand UO_1000 (O_1000,N_19488,N_19669);
nand UO_1001 (O_1001,N_19192,N_19354);
and UO_1002 (O_1002,N_19203,N_19916);
xnor UO_1003 (O_1003,N_19192,N_19120);
and UO_1004 (O_1004,N_19705,N_19966);
xor UO_1005 (O_1005,N_19288,N_19073);
nor UO_1006 (O_1006,N_19969,N_19948);
or UO_1007 (O_1007,N_19399,N_19418);
nand UO_1008 (O_1008,N_19342,N_19627);
nor UO_1009 (O_1009,N_19991,N_19833);
and UO_1010 (O_1010,N_19643,N_19564);
nor UO_1011 (O_1011,N_19067,N_19344);
or UO_1012 (O_1012,N_19190,N_19722);
and UO_1013 (O_1013,N_19489,N_19821);
and UO_1014 (O_1014,N_19115,N_19718);
nand UO_1015 (O_1015,N_19685,N_19471);
or UO_1016 (O_1016,N_19479,N_19728);
or UO_1017 (O_1017,N_19332,N_19220);
or UO_1018 (O_1018,N_19358,N_19040);
or UO_1019 (O_1019,N_19604,N_19038);
xnor UO_1020 (O_1020,N_19467,N_19067);
nor UO_1021 (O_1021,N_19298,N_19270);
or UO_1022 (O_1022,N_19098,N_19794);
nand UO_1023 (O_1023,N_19537,N_19701);
nor UO_1024 (O_1024,N_19897,N_19344);
nor UO_1025 (O_1025,N_19468,N_19115);
or UO_1026 (O_1026,N_19209,N_19728);
or UO_1027 (O_1027,N_19938,N_19564);
xor UO_1028 (O_1028,N_19659,N_19626);
xnor UO_1029 (O_1029,N_19234,N_19322);
xor UO_1030 (O_1030,N_19550,N_19995);
or UO_1031 (O_1031,N_19940,N_19895);
nand UO_1032 (O_1032,N_19104,N_19279);
and UO_1033 (O_1033,N_19953,N_19949);
nand UO_1034 (O_1034,N_19445,N_19015);
or UO_1035 (O_1035,N_19158,N_19795);
nand UO_1036 (O_1036,N_19625,N_19171);
and UO_1037 (O_1037,N_19528,N_19256);
and UO_1038 (O_1038,N_19178,N_19845);
or UO_1039 (O_1039,N_19889,N_19366);
and UO_1040 (O_1040,N_19931,N_19255);
xnor UO_1041 (O_1041,N_19585,N_19896);
and UO_1042 (O_1042,N_19504,N_19273);
and UO_1043 (O_1043,N_19203,N_19292);
or UO_1044 (O_1044,N_19269,N_19780);
nand UO_1045 (O_1045,N_19293,N_19992);
nor UO_1046 (O_1046,N_19326,N_19296);
xnor UO_1047 (O_1047,N_19042,N_19032);
or UO_1048 (O_1048,N_19456,N_19288);
and UO_1049 (O_1049,N_19381,N_19181);
nand UO_1050 (O_1050,N_19736,N_19600);
nand UO_1051 (O_1051,N_19519,N_19762);
xnor UO_1052 (O_1052,N_19505,N_19281);
nand UO_1053 (O_1053,N_19610,N_19916);
xnor UO_1054 (O_1054,N_19885,N_19503);
xor UO_1055 (O_1055,N_19364,N_19943);
or UO_1056 (O_1056,N_19003,N_19194);
and UO_1057 (O_1057,N_19814,N_19490);
xnor UO_1058 (O_1058,N_19269,N_19140);
and UO_1059 (O_1059,N_19085,N_19909);
nand UO_1060 (O_1060,N_19403,N_19708);
xor UO_1061 (O_1061,N_19689,N_19092);
xnor UO_1062 (O_1062,N_19446,N_19918);
or UO_1063 (O_1063,N_19328,N_19426);
nor UO_1064 (O_1064,N_19617,N_19912);
nor UO_1065 (O_1065,N_19576,N_19405);
xor UO_1066 (O_1066,N_19283,N_19788);
and UO_1067 (O_1067,N_19135,N_19295);
and UO_1068 (O_1068,N_19903,N_19628);
and UO_1069 (O_1069,N_19426,N_19436);
xnor UO_1070 (O_1070,N_19570,N_19430);
xor UO_1071 (O_1071,N_19405,N_19729);
and UO_1072 (O_1072,N_19510,N_19361);
xor UO_1073 (O_1073,N_19405,N_19933);
nand UO_1074 (O_1074,N_19332,N_19768);
nand UO_1075 (O_1075,N_19676,N_19921);
nor UO_1076 (O_1076,N_19928,N_19034);
or UO_1077 (O_1077,N_19721,N_19262);
or UO_1078 (O_1078,N_19307,N_19998);
nor UO_1079 (O_1079,N_19018,N_19203);
or UO_1080 (O_1080,N_19338,N_19812);
nand UO_1081 (O_1081,N_19461,N_19388);
nand UO_1082 (O_1082,N_19814,N_19549);
xnor UO_1083 (O_1083,N_19471,N_19630);
nand UO_1084 (O_1084,N_19467,N_19958);
nor UO_1085 (O_1085,N_19490,N_19606);
xor UO_1086 (O_1086,N_19809,N_19958);
xor UO_1087 (O_1087,N_19589,N_19422);
and UO_1088 (O_1088,N_19795,N_19863);
or UO_1089 (O_1089,N_19428,N_19501);
and UO_1090 (O_1090,N_19026,N_19385);
and UO_1091 (O_1091,N_19342,N_19099);
nor UO_1092 (O_1092,N_19317,N_19519);
or UO_1093 (O_1093,N_19966,N_19965);
or UO_1094 (O_1094,N_19640,N_19843);
and UO_1095 (O_1095,N_19329,N_19142);
xor UO_1096 (O_1096,N_19264,N_19677);
nor UO_1097 (O_1097,N_19701,N_19579);
nor UO_1098 (O_1098,N_19671,N_19232);
or UO_1099 (O_1099,N_19932,N_19752);
or UO_1100 (O_1100,N_19648,N_19348);
nor UO_1101 (O_1101,N_19284,N_19149);
xnor UO_1102 (O_1102,N_19348,N_19183);
or UO_1103 (O_1103,N_19796,N_19819);
xor UO_1104 (O_1104,N_19834,N_19121);
and UO_1105 (O_1105,N_19086,N_19123);
or UO_1106 (O_1106,N_19132,N_19994);
or UO_1107 (O_1107,N_19281,N_19931);
nor UO_1108 (O_1108,N_19462,N_19958);
xnor UO_1109 (O_1109,N_19371,N_19999);
and UO_1110 (O_1110,N_19107,N_19600);
nor UO_1111 (O_1111,N_19292,N_19294);
and UO_1112 (O_1112,N_19423,N_19163);
or UO_1113 (O_1113,N_19311,N_19798);
nand UO_1114 (O_1114,N_19372,N_19255);
or UO_1115 (O_1115,N_19730,N_19587);
nor UO_1116 (O_1116,N_19289,N_19154);
nor UO_1117 (O_1117,N_19770,N_19977);
nor UO_1118 (O_1118,N_19446,N_19590);
nor UO_1119 (O_1119,N_19727,N_19304);
xor UO_1120 (O_1120,N_19876,N_19555);
and UO_1121 (O_1121,N_19439,N_19635);
xor UO_1122 (O_1122,N_19394,N_19214);
nand UO_1123 (O_1123,N_19992,N_19978);
and UO_1124 (O_1124,N_19277,N_19698);
and UO_1125 (O_1125,N_19853,N_19969);
nor UO_1126 (O_1126,N_19512,N_19959);
xnor UO_1127 (O_1127,N_19360,N_19564);
and UO_1128 (O_1128,N_19026,N_19807);
and UO_1129 (O_1129,N_19927,N_19598);
xor UO_1130 (O_1130,N_19847,N_19461);
or UO_1131 (O_1131,N_19316,N_19806);
or UO_1132 (O_1132,N_19009,N_19849);
or UO_1133 (O_1133,N_19187,N_19330);
or UO_1134 (O_1134,N_19851,N_19666);
xnor UO_1135 (O_1135,N_19063,N_19522);
nand UO_1136 (O_1136,N_19470,N_19309);
xnor UO_1137 (O_1137,N_19730,N_19420);
and UO_1138 (O_1138,N_19861,N_19512);
and UO_1139 (O_1139,N_19739,N_19059);
xor UO_1140 (O_1140,N_19440,N_19556);
xor UO_1141 (O_1141,N_19859,N_19020);
xnor UO_1142 (O_1142,N_19050,N_19382);
or UO_1143 (O_1143,N_19594,N_19413);
nor UO_1144 (O_1144,N_19470,N_19869);
nand UO_1145 (O_1145,N_19216,N_19253);
and UO_1146 (O_1146,N_19625,N_19689);
xnor UO_1147 (O_1147,N_19303,N_19670);
nor UO_1148 (O_1148,N_19736,N_19718);
and UO_1149 (O_1149,N_19361,N_19359);
and UO_1150 (O_1150,N_19184,N_19671);
xnor UO_1151 (O_1151,N_19212,N_19405);
nor UO_1152 (O_1152,N_19167,N_19335);
and UO_1153 (O_1153,N_19460,N_19667);
nand UO_1154 (O_1154,N_19106,N_19917);
and UO_1155 (O_1155,N_19968,N_19837);
nor UO_1156 (O_1156,N_19287,N_19081);
nand UO_1157 (O_1157,N_19087,N_19284);
or UO_1158 (O_1158,N_19661,N_19116);
xnor UO_1159 (O_1159,N_19179,N_19350);
xnor UO_1160 (O_1160,N_19694,N_19457);
and UO_1161 (O_1161,N_19538,N_19759);
and UO_1162 (O_1162,N_19179,N_19020);
nor UO_1163 (O_1163,N_19203,N_19732);
nor UO_1164 (O_1164,N_19261,N_19916);
or UO_1165 (O_1165,N_19813,N_19732);
nand UO_1166 (O_1166,N_19441,N_19588);
and UO_1167 (O_1167,N_19569,N_19046);
or UO_1168 (O_1168,N_19364,N_19778);
and UO_1169 (O_1169,N_19134,N_19912);
nor UO_1170 (O_1170,N_19720,N_19653);
nand UO_1171 (O_1171,N_19334,N_19720);
nand UO_1172 (O_1172,N_19584,N_19768);
and UO_1173 (O_1173,N_19622,N_19075);
and UO_1174 (O_1174,N_19977,N_19361);
nor UO_1175 (O_1175,N_19343,N_19305);
or UO_1176 (O_1176,N_19896,N_19171);
xnor UO_1177 (O_1177,N_19070,N_19412);
xor UO_1178 (O_1178,N_19430,N_19917);
or UO_1179 (O_1179,N_19294,N_19170);
nand UO_1180 (O_1180,N_19526,N_19797);
and UO_1181 (O_1181,N_19926,N_19835);
and UO_1182 (O_1182,N_19043,N_19954);
and UO_1183 (O_1183,N_19640,N_19868);
xor UO_1184 (O_1184,N_19221,N_19949);
or UO_1185 (O_1185,N_19421,N_19670);
or UO_1186 (O_1186,N_19821,N_19966);
or UO_1187 (O_1187,N_19284,N_19123);
and UO_1188 (O_1188,N_19553,N_19464);
nand UO_1189 (O_1189,N_19849,N_19540);
nand UO_1190 (O_1190,N_19106,N_19446);
and UO_1191 (O_1191,N_19934,N_19776);
xor UO_1192 (O_1192,N_19171,N_19030);
nand UO_1193 (O_1193,N_19781,N_19915);
nand UO_1194 (O_1194,N_19943,N_19255);
and UO_1195 (O_1195,N_19534,N_19402);
or UO_1196 (O_1196,N_19777,N_19127);
or UO_1197 (O_1197,N_19880,N_19574);
or UO_1198 (O_1198,N_19498,N_19994);
nand UO_1199 (O_1199,N_19201,N_19265);
xnor UO_1200 (O_1200,N_19391,N_19505);
and UO_1201 (O_1201,N_19107,N_19767);
nand UO_1202 (O_1202,N_19645,N_19160);
nor UO_1203 (O_1203,N_19098,N_19324);
and UO_1204 (O_1204,N_19379,N_19690);
xnor UO_1205 (O_1205,N_19344,N_19784);
xnor UO_1206 (O_1206,N_19597,N_19830);
nor UO_1207 (O_1207,N_19144,N_19418);
xnor UO_1208 (O_1208,N_19425,N_19232);
and UO_1209 (O_1209,N_19386,N_19892);
or UO_1210 (O_1210,N_19699,N_19931);
and UO_1211 (O_1211,N_19746,N_19872);
xnor UO_1212 (O_1212,N_19302,N_19415);
xnor UO_1213 (O_1213,N_19510,N_19003);
xnor UO_1214 (O_1214,N_19704,N_19605);
nand UO_1215 (O_1215,N_19258,N_19059);
or UO_1216 (O_1216,N_19669,N_19227);
nor UO_1217 (O_1217,N_19073,N_19546);
nor UO_1218 (O_1218,N_19544,N_19028);
and UO_1219 (O_1219,N_19339,N_19175);
nor UO_1220 (O_1220,N_19729,N_19609);
nor UO_1221 (O_1221,N_19774,N_19770);
nand UO_1222 (O_1222,N_19019,N_19775);
nor UO_1223 (O_1223,N_19913,N_19180);
nor UO_1224 (O_1224,N_19483,N_19403);
and UO_1225 (O_1225,N_19774,N_19089);
nand UO_1226 (O_1226,N_19184,N_19919);
nand UO_1227 (O_1227,N_19079,N_19154);
nand UO_1228 (O_1228,N_19809,N_19632);
and UO_1229 (O_1229,N_19717,N_19904);
or UO_1230 (O_1230,N_19703,N_19155);
nor UO_1231 (O_1231,N_19839,N_19531);
and UO_1232 (O_1232,N_19517,N_19583);
nor UO_1233 (O_1233,N_19707,N_19868);
or UO_1234 (O_1234,N_19113,N_19632);
nand UO_1235 (O_1235,N_19605,N_19665);
xnor UO_1236 (O_1236,N_19505,N_19739);
or UO_1237 (O_1237,N_19098,N_19038);
nand UO_1238 (O_1238,N_19714,N_19705);
xor UO_1239 (O_1239,N_19549,N_19172);
and UO_1240 (O_1240,N_19389,N_19975);
nand UO_1241 (O_1241,N_19478,N_19215);
nand UO_1242 (O_1242,N_19882,N_19298);
and UO_1243 (O_1243,N_19064,N_19728);
nand UO_1244 (O_1244,N_19618,N_19008);
nor UO_1245 (O_1245,N_19673,N_19575);
nand UO_1246 (O_1246,N_19562,N_19558);
nand UO_1247 (O_1247,N_19250,N_19764);
xor UO_1248 (O_1248,N_19541,N_19863);
nand UO_1249 (O_1249,N_19615,N_19617);
or UO_1250 (O_1250,N_19945,N_19362);
and UO_1251 (O_1251,N_19401,N_19669);
and UO_1252 (O_1252,N_19455,N_19601);
nand UO_1253 (O_1253,N_19346,N_19102);
and UO_1254 (O_1254,N_19572,N_19348);
nand UO_1255 (O_1255,N_19482,N_19047);
nor UO_1256 (O_1256,N_19026,N_19959);
or UO_1257 (O_1257,N_19789,N_19176);
and UO_1258 (O_1258,N_19014,N_19850);
and UO_1259 (O_1259,N_19606,N_19873);
nand UO_1260 (O_1260,N_19401,N_19227);
or UO_1261 (O_1261,N_19837,N_19133);
nand UO_1262 (O_1262,N_19522,N_19457);
nor UO_1263 (O_1263,N_19943,N_19482);
xor UO_1264 (O_1264,N_19280,N_19467);
nor UO_1265 (O_1265,N_19375,N_19885);
nand UO_1266 (O_1266,N_19088,N_19227);
or UO_1267 (O_1267,N_19626,N_19056);
xnor UO_1268 (O_1268,N_19639,N_19142);
or UO_1269 (O_1269,N_19198,N_19619);
or UO_1270 (O_1270,N_19165,N_19333);
nand UO_1271 (O_1271,N_19886,N_19719);
and UO_1272 (O_1272,N_19120,N_19468);
nor UO_1273 (O_1273,N_19570,N_19927);
nor UO_1274 (O_1274,N_19640,N_19790);
nor UO_1275 (O_1275,N_19191,N_19424);
nor UO_1276 (O_1276,N_19643,N_19091);
or UO_1277 (O_1277,N_19996,N_19385);
or UO_1278 (O_1278,N_19846,N_19277);
nand UO_1279 (O_1279,N_19312,N_19824);
and UO_1280 (O_1280,N_19854,N_19519);
and UO_1281 (O_1281,N_19565,N_19446);
nor UO_1282 (O_1282,N_19949,N_19771);
or UO_1283 (O_1283,N_19887,N_19734);
and UO_1284 (O_1284,N_19194,N_19731);
nor UO_1285 (O_1285,N_19314,N_19138);
nand UO_1286 (O_1286,N_19404,N_19264);
nor UO_1287 (O_1287,N_19069,N_19764);
nor UO_1288 (O_1288,N_19732,N_19621);
nand UO_1289 (O_1289,N_19536,N_19009);
and UO_1290 (O_1290,N_19083,N_19150);
nor UO_1291 (O_1291,N_19720,N_19200);
nand UO_1292 (O_1292,N_19019,N_19246);
nor UO_1293 (O_1293,N_19206,N_19702);
nor UO_1294 (O_1294,N_19513,N_19632);
nor UO_1295 (O_1295,N_19848,N_19328);
xnor UO_1296 (O_1296,N_19863,N_19656);
nand UO_1297 (O_1297,N_19591,N_19930);
and UO_1298 (O_1298,N_19068,N_19870);
xnor UO_1299 (O_1299,N_19507,N_19875);
xor UO_1300 (O_1300,N_19472,N_19763);
nor UO_1301 (O_1301,N_19450,N_19754);
xnor UO_1302 (O_1302,N_19345,N_19265);
or UO_1303 (O_1303,N_19810,N_19003);
nand UO_1304 (O_1304,N_19173,N_19229);
or UO_1305 (O_1305,N_19967,N_19387);
or UO_1306 (O_1306,N_19596,N_19222);
nand UO_1307 (O_1307,N_19940,N_19968);
xnor UO_1308 (O_1308,N_19457,N_19578);
and UO_1309 (O_1309,N_19114,N_19286);
and UO_1310 (O_1310,N_19695,N_19979);
xnor UO_1311 (O_1311,N_19507,N_19128);
nand UO_1312 (O_1312,N_19084,N_19838);
nor UO_1313 (O_1313,N_19526,N_19128);
nor UO_1314 (O_1314,N_19973,N_19479);
nor UO_1315 (O_1315,N_19349,N_19105);
and UO_1316 (O_1316,N_19525,N_19216);
and UO_1317 (O_1317,N_19249,N_19862);
xor UO_1318 (O_1318,N_19119,N_19104);
and UO_1319 (O_1319,N_19079,N_19984);
nor UO_1320 (O_1320,N_19396,N_19407);
nand UO_1321 (O_1321,N_19659,N_19986);
and UO_1322 (O_1322,N_19572,N_19238);
nand UO_1323 (O_1323,N_19047,N_19790);
nand UO_1324 (O_1324,N_19008,N_19300);
or UO_1325 (O_1325,N_19975,N_19598);
and UO_1326 (O_1326,N_19927,N_19078);
xnor UO_1327 (O_1327,N_19083,N_19124);
nor UO_1328 (O_1328,N_19746,N_19322);
xor UO_1329 (O_1329,N_19304,N_19016);
xnor UO_1330 (O_1330,N_19002,N_19731);
nor UO_1331 (O_1331,N_19220,N_19323);
nand UO_1332 (O_1332,N_19407,N_19642);
or UO_1333 (O_1333,N_19410,N_19511);
xnor UO_1334 (O_1334,N_19773,N_19731);
and UO_1335 (O_1335,N_19267,N_19650);
or UO_1336 (O_1336,N_19472,N_19414);
xnor UO_1337 (O_1337,N_19263,N_19605);
nor UO_1338 (O_1338,N_19312,N_19478);
or UO_1339 (O_1339,N_19219,N_19837);
nor UO_1340 (O_1340,N_19161,N_19483);
nand UO_1341 (O_1341,N_19979,N_19906);
xnor UO_1342 (O_1342,N_19839,N_19863);
xnor UO_1343 (O_1343,N_19462,N_19380);
and UO_1344 (O_1344,N_19212,N_19618);
nand UO_1345 (O_1345,N_19620,N_19605);
nand UO_1346 (O_1346,N_19889,N_19277);
and UO_1347 (O_1347,N_19550,N_19540);
or UO_1348 (O_1348,N_19806,N_19779);
or UO_1349 (O_1349,N_19491,N_19888);
and UO_1350 (O_1350,N_19493,N_19654);
nand UO_1351 (O_1351,N_19692,N_19015);
or UO_1352 (O_1352,N_19327,N_19260);
nor UO_1353 (O_1353,N_19400,N_19201);
nand UO_1354 (O_1354,N_19675,N_19785);
nand UO_1355 (O_1355,N_19588,N_19718);
or UO_1356 (O_1356,N_19928,N_19081);
xnor UO_1357 (O_1357,N_19525,N_19981);
nand UO_1358 (O_1358,N_19303,N_19442);
or UO_1359 (O_1359,N_19729,N_19237);
nand UO_1360 (O_1360,N_19943,N_19295);
or UO_1361 (O_1361,N_19165,N_19975);
or UO_1362 (O_1362,N_19005,N_19993);
or UO_1363 (O_1363,N_19440,N_19371);
and UO_1364 (O_1364,N_19616,N_19019);
or UO_1365 (O_1365,N_19251,N_19864);
and UO_1366 (O_1366,N_19235,N_19830);
or UO_1367 (O_1367,N_19406,N_19073);
and UO_1368 (O_1368,N_19221,N_19844);
nand UO_1369 (O_1369,N_19845,N_19552);
or UO_1370 (O_1370,N_19086,N_19480);
nor UO_1371 (O_1371,N_19342,N_19346);
nand UO_1372 (O_1372,N_19269,N_19447);
nand UO_1373 (O_1373,N_19231,N_19079);
xor UO_1374 (O_1374,N_19552,N_19835);
xor UO_1375 (O_1375,N_19368,N_19023);
nand UO_1376 (O_1376,N_19935,N_19764);
nand UO_1377 (O_1377,N_19822,N_19907);
or UO_1378 (O_1378,N_19067,N_19108);
or UO_1379 (O_1379,N_19218,N_19527);
xnor UO_1380 (O_1380,N_19564,N_19455);
xor UO_1381 (O_1381,N_19645,N_19175);
or UO_1382 (O_1382,N_19065,N_19985);
nor UO_1383 (O_1383,N_19497,N_19420);
or UO_1384 (O_1384,N_19569,N_19961);
xnor UO_1385 (O_1385,N_19581,N_19801);
xnor UO_1386 (O_1386,N_19203,N_19820);
or UO_1387 (O_1387,N_19557,N_19890);
xnor UO_1388 (O_1388,N_19904,N_19768);
and UO_1389 (O_1389,N_19086,N_19065);
or UO_1390 (O_1390,N_19782,N_19327);
or UO_1391 (O_1391,N_19675,N_19626);
nor UO_1392 (O_1392,N_19881,N_19124);
nand UO_1393 (O_1393,N_19756,N_19441);
or UO_1394 (O_1394,N_19272,N_19808);
nand UO_1395 (O_1395,N_19042,N_19727);
or UO_1396 (O_1396,N_19831,N_19526);
nand UO_1397 (O_1397,N_19869,N_19372);
xnor UO_1398 (O_1398,N_19872,N_19945);
nand UO_1399 (O_1399,N_19062,N_19529);
nand UO_1400 (O_1400,N_19729,N_19493);
nand UO_1401 (O_1401,N_19798,N_19318);
or UO_1402 (O_1402,N_19692,N_19628);
xnor UO_1403 (O_1403,N_19145,N_19247);
nand UO_1404 (O_1404,N_19470,N_19046);
and UO_1405 (O_1405,N_19831,N_19308);
nor UO_1406 (O_1406,N_19335,N_19967);
and UO_1407 (O_1407,N_19842,N_19077);
and UO_1408 (O_1408,N_19345,N_19999);
or UO_1409 (O_1409,N_19974,N_19220);
or UO_1410 (O_1410,N_19475,N_19437);
nor UO_1411 (O_1411,N_19407,N_19110);
nand UO_1412 (O_1412,N_19254,N_19492);
nand UO_1413 (O_1413,N_19651,N_19307);
nand UO_1414 (O_1414,N_19197,N_19171);
xnor UO_1415 (O_1415,N_19581,N_19139);
or UO_1416 (O_1416,N_19175,N_19712);
nor UO_1417 (O_1417,N_19244,N_19245);
nand UO_1418 (O_1418,N_19470,N_19439);
nor UO_1419 (O_1419,N_19287,N_19100);
and UO_1420 (O_1420,N_19445,N_19958);
nand UO_1421 (O_1421,N_19843,N_19385);
xnor UO_1422 (O_1422,N_19232,N_19109);
or UO_1423 (O_1423,N_19963,N_19342);
xnor UO_1424 (O_1424,N_19181,N_19574);
xor UO_1425 (O_1425,N_19588,N_19276);
or UO_1426 (O_1426,N_19735,N_19678);
and UO_1427 (O_1427,N_19040,N_19031);
nand UO_1428 (O_1428,N_19968,N_19440);
nand UO_1429 (O_1429,N_19868,N_19001);
or UO_1430 (O_1430,N_19489,N_19297);
xor UO_1431 (O_1431,N_19778,N_19087);
and UO_1432 (O_1432,N_19272,N_19074);
nand UO_1433 (O_1433,N_19610,N_19689);
nand UO_1434 (O_1434,N_19434,N_19955);
nor UO_1435 (O_1435,N_19624,N_19367);
xnor UO_1436 (O_1436,N_19882,N_19979);
and UO_1437 (O_1437,N_19830,N_19344);
and UO_1438 (O_1438,N_19258,N_19745);
xor UO_1439 (O_1439,N_19548,N_19474);
nor UO_1440 (O_1440,N_19917,N_19187);
nand UO_1441 (O_1441,N_19939,N_19166);
or UO_1442 (O_1442,N_19881,N_19635);
and UO_1443 (O_1443,N_19838,N_19925);
nor UO_1444 (O_1444,N_19706,N_19295);
or UO_1445 (O_1445,N_19871,N_19522);
nor UO_1446 (O_1446,N_19543,N_19748);
and UO_1447 (O_1447,N_19736,N_19789);
xor UO_1448 (O_1448,N_19463,N_19244);
nand UO_1449 (O_1449,N_19360,N_19066);
nor UO_1450 (O_1450,N_19615,N_19771);
nand UO_1451 (O_1451,N_19539,N_19140);
nor UO_1452 (O_1452,N_19340,N_19697);
nor UO_1453 (O_1453,N_19482,N_19561);
nor UO_1454 (O_1454,N_19339,N_19858);
and UO_1455 (O_1455,N_19933,N_19875);
or UO_1456 (O_1456,N_19449,N_19690);
and UO_1457 (O_1457,N_19595,N_19618);
xnor UO_1458 (O_1458,N_19257,N_19452);
and UO_1459 (O_1459,N_19007,N_19190);
and UO_1460 (O_1460,N_19352,N_19848);
nor UO_1461 (O_1461,N_19729,N_19040);
xor UO_1462 (O_1462,N_19763,N_19951);
nor UO_1463 (O_1463,N_19914,N_19744);
nor UO_1464 (O_1464,N_19686,N_19824);
and UO_1465 (O_1465,N_19187,N_19370);
nor UO_1466 (O_1466,N_19492,N_19641);
or UO_1467 (O_1467,N_19658,N_19450);
nor UO_1468 (O_1468,N_19754,N_19323);
xnor UO_1469 (O_1469,N_19981,N_19467);
xor UO_1470 (O_1470,N_19240,N_19630);
and UO_1471 (O_1471,N_19565,N_19152);
nand UO_1472 (O_1472,N_19354,N_19515);
nand UO_1473 (O_1473,N_19907,N_19053);
or UO_1474 (O_1474,N_19081,N_19428);
or UO_1475 (O_1475,N_19200,N_19756);
xor UO_1476 (O_1476,N_19929,N_19866);
and UO_1477 (O_1477,N_19092,N_19655);
or UO_1478 (O_1478,N_19410,N_19822);
and UO_1479 (O_1479,N_19123,N_19548);
nor UO_1480 (O_1480,N_19922,N_19911);
and UO_1481 (O_1481,N_19440,N_19819);
nand UO_1482 (O_1482,N_19117,N_19850);
nor UO_1483 (O_1483,N_19076,N_19157);
nor UO_1484 (O_1484,N_19095,N_19156);
nor UO_1485 (O_1485,N_19058,N_19965);
and UO_1486 (O_1486,N_19576,N_19115);
and UO_1487 (O_1487,N_19193,N_19235);
xor UO_1488 (O_1488,N_19215,N_19924);
and UO_1489 (O_1489,N_19713,N_19822);
and UO_1490 (O_1490,N_19372,N_19725);
nor UO_1491 (O_1491,N_19614,N_19711);
and UO_1492 (O_1492,N_19404,N_19435);
xor UO_1493 (O_1493,N_19543,N_19411);
nand UO_1494 (O_1494,N_19282,N_19934);
and UO_1495 (O_1495,N_19982,N_19844);
nor UO_1496 (O_1496,N_19792,N_19446);
xor UO_1497 (O_1497,N_19141,N_19481);
nor UO_1498 (O_1498,N_19346,N_19444);
and UO_1499 (O_1499,N_19871,N_19067);
nor UO_1500 (O_1500,N_19132,N_19119);
and UO_1501 (O_1501,N_19821,N_19324);
nand UO_1502 (O_1502,N_19503,N_19911);
nand UO_1503 (O_1503,N_19084,N_19346);
nand UO_1504 (O_1504,N_19374,N_19586);
xnor UO_1505 (O_1505,N_19241,N_19313);
nand UO_1506 (O_1506,N_19474,N_19779);
or UO_1507 (O_1507,N_19001,N_19790);
nand UO_1508 (O_1508,N_19249,N_19792);
nand UO_1509 (O_1509,N_19892,N_19221);
nand UO_1510 (O_1510,N_19402,N_19083);
and UO_1511 (O_1511,N_19232,N_19522);
nand UO_1512 (O_1512,N_19034,N_19160);
or UO_1513 (O_1513,N_19870,N_19949);
xor UO_1514 (O_1514,N_19731,N_19865);
or UO_1515 (O_1515,N_19622,N_19010);
nor UO_1516 (O_1516,N_19337,N_19510);
nand UO_1517 (O_1517,N_19131,N_19026);
nor UO_1518 (O_1518,N_19032,N_19896);
nor UO_1519 (O_1519,N_19774,N_19060);
or UO_1520 (O_1520,N_19346,N_19688);
xnor UO_1521 (O_1521,N_19867,N_19737);
or UO_1522 (O_1522,N_19652,N_19984);
nand UO_1523 (O_1523,N_19831,N_19978);
nor UO_1524 (O_1524,N_19442,N_19466);
xor UO_1525 (O_1525,N_19041,N_19868);
or UO_1526 (O_1526,N_19475,N_19164);
or UO_1527 (O_1527,N_19503,N_19112);
or UO_1528 (O_1528,N_19040,N_19161);
or UO_1529 (O_1529,N_19437,N_19057);
or UO_1530 (O_1530,N_19547,N_19211);
and UO_1531 (O_1531,N_19192,N_19189);
xor UO_1532 (O_1532,N_19165,N_19438);
and UO_1533 (O_1533,N_19317,N_19348);
xor UO_1534 (O_1534,N_19460,N_19040);
and UO_1535 (O_1535,N_19114,N_19975);
or UO_1536 (O_1536,N_19440,N_19710);
nor UO_1537 (O_1537,N_19762,N_19197);
nand UO_1538 (O_1538,N_19810,N_19665);
or UO_1539 (O_1539,N_19979,N_19409);
nor UO_1540 (O_1540,N_19024,N_19479);
nand UO_1541 (O_1541,N_19324,N_19031);
or UO_1542 (O_1542,N_19159,N_19334);
xnor UO_1543 (O_1543,N_19713,N_19439);
or UO_1544 (O_1544,N_19504,N_19511);
xor UO_1545 (O_1545,N_19707,N_19210);
nand UO_1546 (O_1546,N_19906,N_19117);
xor UO_1547 (O_1547,N_19461,N_19173);
nand UO_1548 (O_1548,N_19515,N_19645);
nor UO_1549 (O_1549,N_19568,N_19346);
or UO_1550 (O_1550,N_19122,N_19219);
or UO_1551 (O_1551,N_19923,N_19089);
or UO_1552 (O_1552,N_19944,N_19636);
or UO_1553 (O_1553,N_19419,N_19166);
xor UO_1554 (O_1554,N_19078,N_19571);
xnor UO_1555 (O_1555,N_19637,N_19843);
nand UO_1556 (O_1556,N_19292,N_19942);
xnor UO_1557 (O_1557,N_19326,N_19915);
nand UO_1558 (O_1558,N_19977,N_19138);
nor UO_1559 (O_1559,N_19204,N_19966);
xnor UO_1560 (O_1560,N_19952,N_19628);
or UO_1561 (O_1561,N_19714,N_19444);
nand UO_1562 (O_1562,N_19463,N_19888);
nand UO_1563 (O_1563,N_19950,N_19888);
xnor UO_1564 (O_1564,N_19573,N_19834);
nand UO_1565 (O_1565,N_19072,N_19202);
nand UO_1566 (O_1566,N_19956,N_19958);
or UO_1567 (O_1567,N_19142,N_19555);
and UO_1568 (O_1568,N_19511,N_19985);
xor UO_1569 (O_1569,N_19511,N_19185);
and UO_1570 (O_1570,N_19829,N_19354);
xor UO_1571 (O_1571,N_19292,N_19413);
nor UO_1572 (O_1572,N_19576,N_19030);
xor UO_1573 (O_1573,N_19729,N_19635);
or UO_1574 (O_1574,N_19201,N_19533);
or UO_1575 (O_1575,N_19055,N_19765);
xnor UO_1576 (O_1576,N_19499,N_19110);
and UO_1577 (O_1577,N_19512,N_19910);
nand UO_1578 (O_1578,N_19138,N_19448);
nand UO_1579 (O_1579,N_19384,N_19094);
or UO_1580 (O_1580,N_19389,N_19220);
nor UO_1581 (O_1581,N_19140,N_19216);
nor UO_1582 (O_1582,N_19664,N_19529);
nand UO_1583 (O_1583,N_19464,N_19273);
nand UO_1584 (O_1584,N_19819,N_19882);
xor UO_1585 (O_1585,N_19140,N_19313);
or UO_1586 (O_1586,N_19144,N_19168);
or UO_1587 (O_1587,N_19526,N_19599);
nor UO_1588 (O_1588,N_19579,N_19315);
nand UO_1589 (O_1589,N_19830,N_19664);
nor UO_1590 (O_1590,N_19954,N_19049);
nand UO_1591 (O_1591,N_19300,N_19174);
nand UO_1592 (O_1592,N_19017,N_19805);
nand UO_1593 (O_1593,N_19321,N_19195);
nand UO_1594 (O_1594,N_19918,N_19126);
xnor UO_1595 (O_1595,N_19739,N_19573);
and UO_1596 (O_1596,N_19592,N_19449);
nand UO_1597 (O_1597,N_19226,N_19007);
xnor UO_1598 (O_1598,N_19790,N_19150);
xor UO_1599 (O_1599,N_19452,N_19547);
nor UO_1600 (O_1600,N_19146,N_19503);
and UO_1601 (O_1601,N_19562,N_19154);
or UO_1602 (O_1602,N_19712,N_19810);
or UO_1603 (O_1603,N_19497,N_19610);
xnor UO_1604 (O_1604,N_19154,N_19786);
xnor UO_1605 (O_1605,N_19040,N_19870);
or UO_1606 (O_1606,N_19339,N_19973);
nand UO_1607 (O_1607,N_19386,N_19977);
nand UO_1608 (O_1608,N_19797,N_19528);
xnor UO_1609 (O_1609,N_19317,N_19404);
or UO_1610 (O_1610,N_19429,N_19952);
nand UO_1611 (O_1611,N_19670,N_19849);
nor UO_1612 (O_1612,N_19235,N_19554);
nand UO_1613 (O_1613,N_19476,N_19765);
xnor UO_1614 (O_1614,N_19158,N_19901);
nor UO_1615 (O_1615,N_19531,N_19170);
nor UO_1616 (O_1616,N_19125,N_19709);
and UO_1617 (O_1617,N_19262,N_19703);
nand UO_1618 (O_1618,N_19803,N_19452);
nor UO_1619 (O_1619,N_19959,N_19177);
or UO_1620 (O_1620,N_19626,N_19955);
or UO_1621 (O_1621,N_19772,N_19123);
xnor UO_1622 (O_1622,N_19044,N_19181);
or UO_1623 (O_1623,N_19747,N_19223);
and UO_1624 (O_1624,N_19593,N_19495);
xnor UO_1625 (O_1625,N_19123,N_19239);
xnor UO_1626 (O_1626,N_19652,N_19135);
or UO_1627 (O_1627,N_19177,N_19489);
nand UO_1628 (O_1628,N_19015,N_19541);
or UO_1629 (O_1629,N_19783,N_19159);
nor UO_1630 (O_1630,N_19315,N_19927);
nand UO_1631 (O_1631,N_19992,N_19323);
or UO_1632 (O_1632,N_19853,N_19473);
xor UO_1633 (O_1633,N_19108,N_19205);
or UO_1634 (O_1634,N_19108,N_19062);
xor UO_1635 (O_1635,N_19575,N_19374);
nand UO_1636 (O_1636,N_19348,N_19928);
xnor UO_1637 (O_1637,N_19433,N_19619);
nand UO_1638 (O_1638,N_19363,N_19406);
nand UO_1639 (O_1639,N_19221,N_19555);
nor UO_1640 (O_1640,N_19780,N_19647);
and UO_1641 (O_1641,N_19228,N_19535);
and UO_1642 (O_1642,N_19533,N_19648);
and UO_1643 (O_1643,N_19990,N_19149);
or UO_1644 (O_1644,N_19724,N_19203);
xor UO_1645 (O_1645,N_19088,N_19124);
or UO_1646 (O_1646,N_19490,N_19615);
nor UO_1647 (O_1647,N_19119,N_19729);
or UO_1648 (O_1648,N_19205,N_19925);
or UO_1649 (O_1649,N_19723,N_19536);
nor UO_1650 (O_1650,N_19300,N_19274);
or UO_1651 (O_1651,N_19730,N_19989);
or UO_1652 (O_1652,N_19427,N_19453);
nand UO_1653 (O_1653,N_19231,N_19562);
or UO_1654 (O_1654,N_19878,N_19709);
or UO_1655 (O_1655,N_19778,N_19159);
or UO_1656 (O_1656,N_19438,N_19949);
nor UO_1657 (O_1657,N_19498,N_19346);
or UO_1658 (O_1658,N_19170,N_19209);
or UO_1659 (O_1659,N_19062,N_19538);
nand UO_1660 (O_1660,N_19455,N_19998);
nand UO_1661 (O_1661,N_19704,N_19889);
nand UO_1662 (O_1662,N_19344,N_19083);
nor UO_1663 (O_1663,N_19673,N_19360);
and UO_1664 (O_1664,N_19012,N_19090);
xor UO_1665 (O_1665,N_19621,N_19327);
nand UO_1666 (O_1666,N_19420,N_19556);
xnor UO_1667 (O_1667,N_19807,N_19426);
nand UO_1668 (O_1668,N_19319,N_19960);
or UO_1669 (O_1669,N_19590,N_19335);
xor UO_1670 (O_1670,N_19598,N_19529);
nor UO_1671 (O_1671,N_19458,N_19816);
or UO_1672 (O_1672,N_19368,N_19383);
xnor UO_1673 (O_1673,N_19337,N_19974);
xnor UO_1674 (O_1674,N_19959,N_19712);
or UO_1675 (O_1675,N_19666,N_19328);
xor UO_1676 (O_1676,N_19496,N_19109);
and UO_1677 (O_1677,N_19761,N_19614);
or UO_1678 (O_1678,N_19373,N_19593);
nand UO_1679 (O_1679,N_19126,N_19848);
or UO_1680 (O_1680,N_19089,N_19331);
xnor UO_1681 (O_1681,N_19732,N_19510);
xor UO_1682 (O_1682,N_19659,N_19003);
nand UO_1683 (O_1683,N_19295,N_19872);
nor UO_1684 (O_1684,N_19000,N_19250);
or UO_1685 (O_1685,N_19968,N_19022);
nand UO_1686 (O_1686,N_19867,N_19064);
nor UO_1687 (O_1687,N_19747,N_19380);
or UO_1688 (O_1688,N_19848,N_19712);
nand UO_1689 (O_1689,N_19249,N_19096);
and UO_1690 (O_1690,N_19263,N_19688);
xor UO_1691 (O_1691,N_19788,N_19708);
xnor UO_1692 (O_1692,N_19408,N_19473);
xor UO_1693 (O_1693,N_19142,N_19964);
nand UO_1694 (O_1694,N_19181,N_19933);
and UO_1695 (O_1695,N_19161,N_19270);
nor UO_1696 (O_1696,N_19214,N_19624);
nor UO_1697 (O_1697,N_19145,N_19222);
nor UO_1698 (O_1698,N_19892,N_19550);
xnor UO_1699 (O_1699,N_19816,N_19925);
and UO_1700 (O_1700,N_19743,N_19766);
xor UO_1701 (O_1701,N_19893,N_19428);
nand UO_1702 (O_1702,N_19662,N_19303);
and UO_1703 (O_1703,N_19807,N_19751);
xnor UO_1704 (O_1704,N_19155,N_19403);
nand UO_1705 (O_1705,N_19282,N_19507);
or UO_1706 (O_1706,N_19728,N_19192);
and UO_1707 (O_1707,N_19608,N_19164);
and UO_1708 (O_1708,N_19122,N_19164);
or UO_1709 (O_1709,N_19461,N_19398);
and UO_1710 (O_1710,N_19332,N_19436);
nor UO_1711 (O_1711,N_19627,N_19849);
nand UO_1712 (O_1712,N_19760,N_19600);
and UO_1713 (O_1713,N_19459,N_19927);
nand UO_1714 (O_1714,N_19588,N_19332);
and UO_1715 (O_1715,N_19531,N_19557);
nor UO_1716 (O_1716,N_19518,N_19870);
or UO_1717 (O_1717,N_19959,N_19784);
or UO_1718 (O_1718,N_19106,N_19379);
or UO_1719 (O_1719,N_19998,N_19510);
and UO_1720 (O_1720,N_19735,N_19787);
nor UO_1721 (O_1721,N_19483,N_19924);
nand UO_1722 (O_1722,N_19965,N_19757);
or UO_1723 (O_1723,N_19391,N_19667);
or UO_1724 (O_1724,N_19777,N_19568);
and UO_1725 (O_1725,N_19374,N_19247);
xor UO_1726 (O_1726,N_19521,N_19694);
or UO_1727 (O_1727,N_19449,N_19297);
and UO_1728 (O_1728,N_19025,N_19183);
and UO_1729 (O_1729,N_19259,N_19783);
nor UO_1730 (O_1730,N_19628,N_19814);
nand UO_1731 (O_1731,N_19643,N_19884);
nand UO_1732 (O_1732,N_19761,N_19758);
nand UO_1733 (O_1733,N_19667,N_19669);
nand UO_1734 (O_1734,N_19837,N_19232);
or UO_1735 (O_1735,N_19960,N_19128);
and UO_1736 (O_1736,N_19846,N_19957);
nor UO_1737 (O_1737,N_19129,N_19199);
or UO_1738 (O_1738,N_19532,N_19078);
xor UO_1739 (O_1739,N_19623,N_19987);
nand UO_1740 (O_1740,N_19028,N_19025);
xor UO_1741 (O_1741,N_19337,N_19388);
nand UO_1742 (O_1742,N_19649,N_19702);
xnor UO_1743 (O_1743,N_19368,N_19462);
xnor UO_1744 (O_1744,N_19050,N_19673);
or UO_1745 (O_1745,N_19703,N_19891);
xnor UO_1746 (O_1746,N_19560,N_19328);
or UO_1747 (O_1747,N_19881,N_19487);
nand UO_1748 (O_1748,N_19024,N_19346);
xor UO_1749 (O_1749,N_19223,N_19387);
nor UO_1750 (O_1750,N_19048,N_19415);
or UO_1751 (O_1751,N_19504,N_19579);
and UO_1752 (O_1752,N_19410,N_19504);
xor UO_1753 (O_1753,N_19571,N_19342);
and UO_1754 (O_1754,N_19046,N_19908);
nor UO_1755 (O_1755,N_19221,N_19273);
nand UO_1756 (O_1756,N_19458,N_19071);
xnor UO_1757 (O_1757,N_19268,N_19979);
nand UO_1758 (O_1758,N_19219,N_19597);
nand UO_1759 (O_1759,N_19122,N_19564);
nor UO_1760 (O_1760,N_19790,N_19765);
and UO_1761 (O_1761,N_19862,N_19663);
nor UO_1762 (O_1762,N_19900,N_19653);
xnor UO_1763 (O_1763,N_19952,N_19525);
nand UO_1764 (O_1764,N_19923,N_19143);
or UO_1765 (O_1765,N_19816,N_19198);
or UO_1766 (O_1766,N_19967,N_19476);
xnor UO_1767 (O_1767,N_19792,N_19922);
xor UO_1768 (O_1768,N_19960,N_19238);
nor UO_1769 (O_1769,N_19991,N_19892);
xor UO_1770 (O_1770,N_19094,N_19097);
and UO_1771 (O_1771,N_19223,N_19776);
xor UO_1772 (O_1772,N_19356,N_19604);
nand UO_1773 (O_1773,N_19324,N_19818);
nor UO_1774 (O_1774,N_19510,N_19329);
xnor UO_1775 (O_1775,N_19008,N_19601);
or UO_1776 (O_1776,N_19353,N_19589);
or UO_1777 (O_1777,N_19446,N_19394);
nand UO_1778 (O_1778,N_19926,N_19502);
nand UO_1779 (O_1779,N_19904,N_19223);
and UO_1780 (O_1780,N_19898,N_19215);
or UO_1781 (O_1781,N_19926,N_19393);
and UO_1782 (O_1782,N_19968,N_19707);
nand UO_1783 (O_1783,N_19490,N_19867);
nor UO_1784 (O_1784,N_19463,N_19535);
or UO_1785 (O_1785,N_19042,N_19930);
or UO_1786 (O_1786,N_19652,N_19020);
xnor UO_1787 (O_1787,N_19232,N_19806);
xor UO_1788 (O_1788,N_19374,N_19395);
nand UO_1789 (O_1789,N_19150,N_19363);
nor UO_1790 (O_1790,N_19878,N_19482);
and UO_1791 (O_1791,N_19679,N_19978);
or UO_1792 (O_1792,N_19055,N_19370);
and UO_1793 (O_1793,N_19579,N_19676);
xor UO_1794 (O_1794,N_19947,N_19418);
nor UO_1795 (O_1795,N_19077,N_19635);
or UO_1796 (O_1796,N_19225,N_19049);
xnor UO_1797 (O_1797,N_19021,N_19328);
or UO_1798 (O_1798,N_19110,N_19932);
nor UO_1799 (O_1799,N_19946,N_19106);
nor UO_1800 (O_1800,N_19086,N_19393);
nand UO_1801 (O_1801,N_19579,N_19604);
nor UO_1802 (O_1802,N_19443,N_19501);
or UO_1803 (O_1803,N_19839,N_19782);
xnor UO_1804 (O_1804,N_19084,N_19471);
nor UO_1805 (O_1805,N_19937,N_19995);
nor UO_1806 (O_1806,N_19936,N_19997);
and UO_1807 (O_1807,N_19261,N_19191);
nor UO_1808 (O_1808,N_19006,N_19719);
or UO_1809 (O_1809,N_19107,N_19121);
nand UO_1810 (O_1810,N_19191,N_19213);
xor UO_1811 (O_1811,N_19564,N_19054);
and UO_1812 (O_1812,N_19437,N_19604);
or UO_1813 (O_1813,N_19089,N_19747);
or UO_1814 (O_1814,N_19092,N_19427);
or UO_1815 (O_1815,N_19118,N_19285);
nand UO_1816 (O_1816,N_19182,N_19526);
or UO_1817 (O_1817,N_19338,N_19176);
nand UO_1818 (O_1818,N_19358,N_19333);
xor UO_1819 (O_1819,N_19420,N_19930);
and UO_1820 (O_1820,N_19231,N_19584);
and UO_1821 (O_1821,N_19331,N_19475);
and UO_1822 (O_1822,N_19605,N_19671);
or UO_1823 (O_1823,N_19052,N_19711);
or UO_1824 (O_1824,N_19958,N_19170);
nand UO_1825 (O_1825,N_19399,N_19424);
and UO_1826 (O_1826,N_19557,N_19898);
and UO_1827 (O_1827,N_19939,N_19782);
nor UO_1828 (O_1828,N_19840,N_19762);
nor UO_1829 (O_1829,N_19438,N_19190);
nor UO_1830 (O_1830,N_19274,N_19191);
or UO_1831 (O_1831,N_19079,N_19813);
xor UO_1832 (O_1832,N_19439,N_19185);
and UO_1833 (O_1833,N_19031,N_19611);
nand UO_1834 (O_1834,N_19893,N_19388);
nand UO_1835 (O_1835,N_19313,N_19202);
or UO_1836 (O_1836,N_19318,N_19832);
xnor UO_1837 (O_1837,N_19725,N_19360);
and UO_1838 (O_1838,N_19880,N_19756);
nand UO_1839 (O_1839,N_19881,N_19589);
and UO_1840 (O_1840,N_19710,N_19203);
xor UO_1841 (O_1841,N_19466,N_19782);
nand UO_1842 (O_1842,N_19195,N_19277);
nor UO_1843 (O_1843,N_19568,N_19292);
xor UO_1844 (O_1844,N_19818,N_19950);
nand UO_1845 (O_1845,N_19059,N_19589);
and UO_1846 (O_1846,N_19290,N_19538);
and UO_1847 (O_1847,N_19105,N_19432);
or UO_1848 (O_1848,N_19243,N_19027);
nor UO_1849 (O_1849,N_19775,N_19023);
nor UO_1850 (O_1850,N_19524,N_19203);
nand UO_1851 (O_1851,N_19117,N_19884);
and UO_1852 (O_1852,N_19982,N_19673);
xor UO_1853 (O_1853,N_19745,N_19947);
nor UO_1854 (O_1854,N_19768,N_19588);
or UO_1855 (O_1855,N_19227,N_19678);
and UO_1856 (O_1856,N_19129,N_19892);
or UO_1857 (O_1857,N_19421,N_19827);
xor UO_1858 (O_1858,N_19296,N_19223);
nand UO_1859 (O_1859,N_19926,N_19610);
nor UO_1860 (O_1860,N_19941,N_19716);
and UO_1861 (O_1861,N_19296,N_19712);
or UO_1862 (O_1862,N_19748,N_19622);
or UO_1863 (O_1863,N_19207,N_19690);
and UO_1864 (O_1864,N_19797,N_19162);
xor UO_1865 (O_1865,N_19249,N_19927);
nor UO_1866 (O_1866,N_19379,N_19882);
or UO_1867 (O_1867,N_19885,N_19935);
or UO_1868 (O_1868,N_19345,N_19150);
xor UO_1869 (O_1869,N_19395,N_19644);
nand UO_1870 (O_1870,N_19380,N_19836);
xor UO_1871 (O_1871,N_19096,N_19677);
xnor UO_1872 (O_1872,N_19935,N_19365);
nand UO_1873 (O_1873,N_19319,N_19649);
or UO_1874 (O_1874,N_19324,N_19638);
nand UO_1875 (O_1875,N_19308,N_19119);
and UO_1876 (O_1876,N_19458,N_19667);
nor UO_1877 (O_1877,N_19510,N_19044);
or UO_1878 (O_1878,N_19980,N_19145);
and UO_1879 (O_1879,N_19238,N_19755);
xnor UO_1880 (O_1880,N_19958,N_19804);
and UO_1881 (O_1881,N_19509,N_19340);
and UO_1882 (O_1882,N_19356,N_19202);
nand UO_1883 (O_1883,N_19319,N_19941);
xor UO_1884 (O_1884,N_19114,N_19845);
and UO_1885 (O_1885,N_19802,N_19919);
and UO_1886 (O_1886,N_19057,N_19819);
xor UO_1887 (O_1887,N_19175,N_19875);
nand UO_1888 (O_1888,N_19893,N_19954);
and UO_1889 (O_1889,N_19572,N_19850);
nand UO_1890 (O_1890,N_19220,N_19689);
nand UO_1891 (O_1891,N_19799,N_19393);
and UO_1892 (O_1892,N_19828,N_19417);
nand UO_1893 (O_1893,N_19575,N_19819);
nor UO_1894 (O_1894,N_19413,N_19655);
and UO_1895 (O_1895,N_19303,N_19966);
nor UO_1896 (O_1896,N_19043,N_19713);
xnor UO_1897 (O_1897,N_19312,N_19777);
nor UO_1898 (O_1898,N_19254,N_19560);
xnor UO_1899 (O_1899,N_19999,N_19842);
and UO_1900 (O_1900,N_19154,N_19514);
nand UO_1901 (O_1901,N_19597,N_19145);
xnor UO_1902 (O_1902,N_19542,N_19471);
xnor UO_1903 (O_1903,N_19399,N_19626);
or UO_1904 (O_1904,N_19268,N_19154);
xor UO_1905 (O_1905,N_19805,N_19015);
nand UO_1906 (O_1906,N_19915,N_19661);
or UO_1907 (O_1907,N_19162,N_19011);
or UO_1908 (O_1908,N_19615,N_19185);
xnor UO_1909 (O_1909,N_19833,N_19505);
and UO_1910 (O_1910,N_19960,N_19050);
or UO_1911 (O_1911,N_19066,N_19934);
and UO_1912 (O_1912,N_19851,N_19226);
nand UO_1913 (O_1913,N_19302,N_19253);
nor UO_1914 (O_1914,N_19029,N_19701);
xnor UO_1915 (O_1915,N_19446,N_19257);
and UO_1916 (O_1916,N_19181,N_19429);
nand UO_1917 (O_1917,N_19102,N_19667);
nor UO_1918 (O_1918,N_19101,N_19290);
and UO_1919 (O_1919,N_19876,N_19465);
and UO_1920 (O_1920,N_19464,N_19417);
nor UO_1921 (O_1921,N_19390,N_19693);
nand UO_1922 (O_1922,N_19909,N_19589);
nand UO_1923 (O_1923,N_19291,N_19684);
and UO_1924 (O_1924,N_19001,N_19168);
or UO_1925 (O_1925,N_19274,N_19542);
or UO_1926 (O_1926,N_19793,N_19521);
nor UO_1927 (O_1927,N_19299,N_19256);
or UO_1928 (O_1928,N_19429,N_19348);
nand UO_1929 (O_1929,N_19400,N_19811);
or UO_1930 (O_1930,N_19648,N_19718);
xor UO_1931 (O_1931,N_19838,N_19236);
xnor UO_1932 (O_1932,N_19316,N_19072);
nand UO_1933 (O_1933,N_19169,N_19868);
and UO_1934 (O_1934,N_19411,N_19650);
and UO_1935 (O_1935,N_19205,N_19062);
and UO_1936 (O_1936,N_19132,N_19577);
xnor UO_1937 (O_1937,N_19385,N_19908);
nor UO_1938 (O_1938,N_19499,N_19957);
nor UO_1939 (O_1939,N_19492,N_19918);
nor UO_1940 (O_1940,N_19474,N_19049);
or UO_1941 (O_1941,N_19539,N_19786);
nor UO_1942 (O_1942,N_19347,N_19670);
xnor UO_1943 (O_1943,N_19100,N_19860);
or UO_1944 (O_1944,N_19611,N_19951);
xor UO_1945 (O_1945,N_19978,N_19098);
nor UO_1946 (O_1946,N_19350,N_19046);
and UO_1947 (O_1947,N_19170,N_19245);
nand UO_1948 (O_1948,N_19823,N_19493);
nand UO_1949 (O_1949,N_19151,N_19560);
nand UO_1950 (O_1950,N_19567,N_19901);
nand UO_1951 (O_1951,N_19448,N_19217);
or UO_1952 (O_1952,N_19846,N_19350);
nand UO_1953 (O_1953,N_19201,N_19818);
xnor UO_1954 (O_1954,N_19278,N_19427);
or UO_1955 (O_1955,N_19354,N_19748);
xor UO_1956 (O_1956,N_19658,N_19545);
nand UO_1957 (O_1957,N_19058,N_19200);
nand UO_1958 (O_1958,N_19951,N_19333);
xor UO_1959 (O_1959,N_19360,N_19215);
nand UO_1960 (O_1960,N_19495,N_19723);
xnor UO_1961 (O_1961,N_19392,N_19063);
or UO_1962 (O_1962,N_19742,N_19065);
and UO_1963 (O_1963,N_19354,N_19898);
and UO_1964 (O_1964,N_19012,N_19586);
and UO_1965 (O_1965,N_19829,N_19278);
nor UO_1966 (O_1966,N_19366,N_19296);
and UO_1967 (O_1967,N_19403,N_19080);
xor UO_1968 (O_1968,N_19494,N_19455);
nor UO_1969 (O_1969,N_19120,N_19489);
nand UO_1970 (O_1970,N_19849,N_19614);
and UO_1971 (O_1971,N_19582,N_19022);
nand UO_1972 (O_1972,N_19017,N_19019);
nor UO_1973 (O_1973,N_19303,N_19812);
nand UO_1974 (O_1974,N_19579,N_19382);
nor UO_1975 (O_1975,N_19116,N_19378);
nor UO_1976 (O_1976,N_19775,N_19048);
and UO_1977 (O_1977,N_19230,N_19799);
xor UO_1978 (O_1978,N_19590,N_19487);
nand UO_1979 (O_1979,N_19940,N_19396);
and UO_1980 (O_1980,N_19069,N_19216);
and UO_1981 (O_1981,N_19068,N_19048);
nor UO_1982 (O_1982,N_19197,N_19280);
and UO_1983 (O_1983,N_19107,N_19342);
or UO_1984 (O_1984,N_19352,N_19711);
or UO_1985 (O_1985,N_19266,N_19750);
and UO_1986 (O_1986,N_19641,N_19826);
xnor UO_1987 (O_1987,N_19937,N_19355);
and UO_1988 (O_1988,N_19615,N_19986);
nor UO_1989 (O_1989,N_19080,N_19711);
and UO_1990 (O_1990,N_19174,N_19831);
and UO_1991 (O_1991,N_19106,N_19990);
or UO_1992 (O_1992,N_19488,N_19348);
xor UO_1993 (O_1993,N_19710,N_19721);
or UO_1994 (O_1994,N_19174,N_19244);
xor UO_1995 (O_1995,N_19063,N_19638);
nand UO_1996 (O_1996,N_19175,N_19340);
xor UO_1997 (O_1997,N_19867,N_19243);
and UO_1998 (O_1998,N_19651,N_19218);
nor UO_1999 (O_1999,N_19015,N_19128);
nor UO_2000 (O_2000,N_19624,N_19721);
nor UO_2001 (O_2001,N_19893,N_19858);
and UO_2002 (O_2002,N_19208,N_19494);
nor UO_2003 (O_2003,N_19675,N_19566);
or UO_2004 (O_2004,N_19333,N_19809);
nand UO_2005 (O_2005,N_19061,N_19391);
nand UO_2006 (O_2006,N_19718,N_19803);
nand UO_2007 (O_2007,N_19250,N_19742);
and UO_2008 (O_2008,N_19245,N_19327);
xor UO_2009 (O_2009,N_19460,N_19969);
and UO_2010 (O_2010,N_19892,N_19672);
nand UO_2011 (O_2011,N_19080,N_19035);
and UO_2012 (O_2012,N_19460,N_19256);
nand UO_2013 (O_2013,N_19291,N_19479);
nand UO_2014 (O_2014,N_19983,N_19507);
and UO_2015 (O_2015,N_19539,N_19820);
and UO_2016 (O_2016,N_19355,N_19459);
xor UO_2017 (O_2017,N_19564,N_19608);
nor UO_2018 (O_2018,N_19236,N_19508);
xor UO_2019 (O_2019,N_19192,N_19090);
nand UO_2020 (O_2020,N_19638,N_19983);
or UO_2021 (O_2021,N_19218,N_19742);
nor UO_2022 (O_2022,N_19257,N_19358);
and UO_2023 (O_2023,N_19491,N_19168);
and UO_2024 (O_2024,N_19324,N_19693);
or UO_2025 (O_2025,N_19411,N_19460);
nor UO_2026 (O_2026,N_19106,N_19090);
nand UO_2027 (O_2027,N_19272,N_19208);
or UO_2028 (O_2028,N_19265,N_19569);
nand UO_2029 (O_2029,N_19677,N_19095);
or UO_2030 (O_2030,N_19878,N_19133);
and UO_2031 (O_2031,N_19194,N_19376);
xor UO_2032 (O_2032,N_19042,N_19982);
xnor UO_2033 (O_2033,N_19625,N_19062);
nor UO_2034 (O_2034,N_19638,N_19824);
xor UO_2035 (O_2035,N_19844,N_19396);
and UO_2036 (O_2036,N_19001,N_19301);
or UO_2037 (O_2037,N_19130,N_19940);
and UO_2038 (O_2038,N_19069,N_19997);
xor UO_2039 (O_2039,N_19524,N_19830);
or UO_2040 (O_2040,N_19342,N_19489);
nor UO_2041 (O_2041,N_19201,N_19330);
or UO_2042 (O_2042,N_19894,N_19606);
xor UO_2043 (O_2043,N_19377,N_19426);
nor UO_2044 (O_2044,N_19984,N_19422);
nor UO_2045 (O_2045,N_19886,N_19073);
and UO_2046 (O_2046,N_19591,N_19788);
nor UO_2047 (O_2047,N_19483,N_19966);
xor UO_2048 (O_2048,N_19933,N_19294);
nor UO_2049 (O_2049,N_19137,N_19176);
xor UO_2050 (O_2050,N_19662,N_19700);
nand UO_2051 (O_2051,N_19706,N_19026);
and UO_2052 (O_2052,N_19162,N_19584);
xnor UO_2053 (O_2053,N_19583,N_19795);
nor UO_2054 (O_2054,N_19761,N_19846);
nand UO_2055 (O_2055,N_19960,N_19418);
and UO_2056 (O_2056,N_19537,N_19543);
or UO_2057 (O_2057,N_19342,N_19801);
xor UO_2058 (O_2058,N_19733,N_19919);
and UO_2059 (O_2059,N_19003,N_19377);
xor UO_2060 (O_2060,N_19762,N_19863);
or UO_2061 (O_2061,N_19348,N_19342);
nor UO_2062 (O_2062,N_19787,N_19533);
or UO_2063 (O_2063,N_19894,N_19903);
or UO_2064 (O_2064,N_19647,N_19186);
nor UO_2065 (O_2065,N_19573,N_19093);
and UO_2066 (O_2066,N_19851,N_19388);
and UO_2067 (O_2067,N_19289,N_19776);
or UO_2068 (O_2068,N_19207,N_19706);
or UO_2069 (O_2069,N_19459,N_19032);
nor UO_2070 (O_2070,N_19409,N_19989);
xnor UO_2071 (O_2071,N_19359,N_19100);
and UO_2072 (O_2072,N_19598,N_19030);
xnor UO_2073 (O_2073,N_19259,N_19725);
or UO_2074 (O_2074,N_19143,N_19763);
and UO_2075 (O_2075,N_19363,N_19865);
or UO_2076 (O_2076,N_19425,N_19110);
nand UO_2077 (O_2077,N_19842,N_19190);
nand UO_2078 (O_2078,N_19384,N_19253);
xor UO_2079 (O_2079,N_19430,N_19641);
and UO_2080 (O_2080,N_19613,N_19951);
nor UO_2081 (O_2081,N_19935,N_19314);
and UO_2082 (O_2082,N_19261,N_19169);
xor UO_2083 (O_2083,N_19235,N_19362);
xor UO_2084 (O_2084,N_19039,N_19146);
and UO_2085 (O_2085,N_19695,N_19965);
or UO_2086 (O_2086,N_19142,N_19981);
xnor UO_2087 (O_2087,N_19043,N_19331);
and UO_2088 (O_2088,N_19296,N_19132);
and UO_2089 (O_2089,N_19889,N_19699);
and UO_2090 (O_2090,N_19347,N_19009);
or UO_2091 (O_2091,N_19289,N_19097);
or UO_2092 (O_2092,N_19567,N_19924);
or UO_2093 (O_2093,N_19576,N_19314);
and UO_2094 (O_2094,N_19599,N_19169);
or UO_2095 (O_2095,N_19737,N_19118);
nor UO_2096 (O_2096,N_19936,N_19002);
xnor UO_2097 (O_2097,N_19599,N_19342);
and UO_2098 (O_2098,N_19697,N_19199);
xor UO_2099 (O_2099,N_19826,N_19727);
nand UO_2100 (O_2100,N_19552,N_19478);
nand UO_2101 (O_2101,N_19895,N_19713);
and UO_2102 (O_2102,N_19013,N_19439);
nor UO_2103 (O_2103,N_19111,N_19831);
or UO_2104 (O_2104,N_19832,N_19121);
nor UO_2105 (O_2105,N_19451,N_19036);
and UO_2106 (O_2106,N_19298,N_19528);
xor UO_2107 (O_2107,N_19360,N_19212);
nor UO_2108 (O_2108,N_19955,N_19653);
nor UO_2109 (O_2109,N_19982,N_19861);
nand UO_2110 (O_2110,N_19420,N_19870);
or UO_2111 (O_2111,N_19418,N_19451);
or UO_2112 (O_2112,N_19475,N_19939);
and UO_2113 (O_2113,N_19378,N_19379);
or UO_2114 (O_2114,N_19595,N_19778);
nor UO_2115 (O_2115,N_19083,N_19153);
xnor UO_2116 (O_2116,N_19496,N_19636);
xor UO_2117 (O_2117,N_19204,N_19977);
or UO_2118 (O_2118,N_19555,N_19533);
xnor UO_2119 (O_2119,N_19154,N_19954);
or UO_2120 (O_2120,N_19174,N_19183);
nand UO_2121 (O_2121,N_19566,N_19903);
and UO_2122 (O_2122,N_19477,N_19201);
nand UO_2123 (O_2123,N_19050,N_19715);
xor UO_2124 (O_2124,N_19591,N_19493);
nor UO_2125 (O_2125,N_19463,N_19399);
nor UO_2126 (O_2126,N_19441,N_19404);
nand UO_2127 (O_2127,N_19637,N_19483);
or UO_2128 (O_2128,N_19435,N_19421);
xor UO_2129 (O_2129,N_19091,N_19104);
or UO_2130 (O_2130,N_19158,N_19438);
and UO_2131 (O_2131,N_19987,N_19596);
nand UO_2132 (O_2132,N_19845,N_19670);
nand UO_2133 (O_2133,N_19250,N_19556);
nand UO_2134 (O_2134,N_19638,N_19952);
nand UO_2135 (O_2135,N_19826,N_19534);
and UO_2136 (O_2136,N_19996,N_19703);
nand UO_2137 (O_2137,N_19514,N_19878);
or UO_2138 (O_2138,N_19834,N_19928);
or UO_2139 (O_2139,N_19511,N_19460);
and UO_2140 (O_2140,N_19207,N_19868);
nand UO_2141 (O_2141,N_19668,N_19293);
or UO_2142 (O_2142,N_19637,N_19236);
nor UO_2143 (O_2143,N_19717,N_19802);
or UO_2144 (O_2144,N_19893,N_19969);
or UO_2145 (O_2145,N_19371,N_19687);
and UO_2146 (O_2146,N_19596,N_19283);
and UO_2147 (O_2147,N_19407,N_19779);
nor UO_2148 (O_2148,N_19786,N_19958);
or UO_2149 (O_2149,N_19333,N_19948);
and UO_2150 (O_2150,N_19395,N_19517);
nor UO_2151 (O_2151,N_19895,N_19770);
and UO_2152 (O_2152,N_19952,N_19996);
and UO_2153 (O_2153,N_19128,N_19601);
xor UO_2154 (O_2154,N_19113,N_19366);
and UO_2155 (O_2155,N_19616,N_19869);
and UO_2156 (O_2156,N_19130,N_19994);
or UO_2157 (O_2157,N_19908,N_19368);
xor UO_2158 (O_2158,N_19196,N_19775);
xor UO_2159 (O_2159,N_19931,N_19193);
or UO_2160 (O_2160,N_19147,N_19076);
nor UO_2161 (O_2161,N_19936,N_19712);
and UO_2162 (O_2162,N_19856,N_19085);
or UO_2163 (O_2163,N_19587,N_19684);
and UO_2164 (O_2164,N_19835,N_19262);
xnor UO_2165 (O_2165,N_19442,N_19401);
or UO_2166 (O_2166,N_19541,N_19025);
xor UO_2167 (O_2167,N_19268,N_19401);
and UO_2168 (O_2168,N_19033,N_19675);
nand UO_2169 (O_2169,N_19517,N_19455);
and UO_2170 (O_2170,N_19751,N_19434);
or UO_2171 (O_2171,N_19944,N_19333);
and UO_2172 (O_2172,N_19066,N_19359);
nand UO_2173 (O_2173,N_19049,N_19250);
nor UO_2174 (O_2174,N_19146,N_19112);
or UO_2175 (O_2175,N_19486,N_19781);
nor UO_2176 (O_2176,N_19686,N_19877);
nor UO_2177 (O_2177,N_19726,N_19226);
nand UO_2178 (O_2178,N_19627,N_19350);
or UO_2179 (O_2179,N_19460,N_19158);
xnor UO_2180 (O_2180,N_19732,N_19288);
nand UO_2181 (O_2181,N_19819,N_19862);
xor UO_2182 (O_2182,N_19223,N_19966);
and UO_2183 (O_2183,N_19013,N_19339);
nand UO_2184 (O_2184,N_19071,N_19792);
nand UO_2185 (O_2185,N_19853,N_19953);
xor UO_2186 (O_2186,N_19990,N_19931);
xnor UO_2187 (O_2187,N_19089,N_19738);
nand UO_2188 (O_2188,N_19512,N_19615);
and UO_2189 (O_2189,N_19215,N_19997);
or UO_2190 (O_2190,N_19990,N_19972);
nor UO_2191 (O_2191,N_19060,N_19226);
nand UO_2192 (O_2192,N_19136,N_19083);
and UO_2193 (O_2193,N_19833,N_19873);
and UO_2194 (O_2194,N_19068,N_19615);
nor UO_2195 (O_2195,N_19209,N_19410);
or UO_2196 (O_2196,N_19087,N_19240);
nor UO_2197 (O_2197,N_19481,N_19906);
or UO_2198 (O_2198,N_19905,N_19328);
or UO_2199 (O_2199,N_19186,N_19439);
xnor UO_2200 (O_2200,N_19746,N_19989);
xnor UO_2201 (O_2201,N_19018,N_19282);
and UO_2202 (O_2202,N_19584,N_19949);
xor UO_2203 (O_2203,N_19231,N_19284);
nand UO_2204 (O_2204,N_19762,N_19072);
xor UO_2205 (O_2205,N_19422,N_19194);
or UO_2206 (O_2206,N_19251,N_19271);
or UO_2207 (O_2207,N_19429,N_19840);
and UO_2208 (O_2208,N_19527,N_19222);
and UO_2209 (O_2209,N_19298,N_19200);
nor UO_2210 (O_2210,N_19716,N_19577);
and UO_2211 (O_2211,N_19961,N_19093);
xnor UO_2212 (O_2212,N_19014,N_19241);
nand UO_2213 (O_2213,N_19521,N_19587);
or UO_2214 (O_2214,N_19472,N_19400);
xor UO_2215 (O_2215,N_19355,N_19215);
and UO_2216 (O_2216,N_19625,N_19967);
xnor UO_2217 (O_2217,N_19507,N_19248);
or UO_2218 (O_2218,N_19948,N_19710);
nor UO_2219 (O_2219,N_19561,N_19642);
nand UO_2220 (O_2220,N_19654,N_19038);
nor UO_2221 (O_2221,N_19827,N_19534);
and UO_2222 (O_2222,N_19068,N_19167);
nor UO_2223 (O_2223,N_19434,N_19557);
xor UO_2224 (O_2224,N_19503,N_19350);
and UO_2225 (O_2225,N_19397,N_19888);
nand UO_2226 (O_2226,N_19494,N_19959);
and UO_2227 (O_2227,N_19499,N_19287);
nand UO_2228 (O_2228,N_19731,N_19441);
or UO_2229 (O_2229,N_19172,N_19595);
xor UO_2230 (O_2230,N_19787,N_19922);
and UO_2231 (O_2231,N_19912,N_19444);
nor UO_2232 (O_2232,N_19746,N_19779);
or UO_2233 (O_2233,N_19981,N_19827);
nand UO_2234 (O_2234,N_19945,N_19818);
nand UO_2235 (O_2235,N_19934,N_19366);
nor UO_2236 (O_2236,N_19914,N_19982);
and UO_2237 (O_2237,N_19617,N_19793);
xnor UO_2238 (O_2238,N_19747,N_19244);
nor UO_2239 (O_2239,N_19631,N_19385);
xor UO_2240 (O_2240,N_19704,N_19097);
and UO_2241 (O_2241,N_19385,N_19812);
xnor UO_2242 (O_2242,N_19439,N_19782);
nand UO_2243 (O_2243,N_19481,N_19246);
nand UO_2244 (O_2244,N_19486,N_19886);
nand UO_2245 (O_2245,N_19857,N_19077);
and UO_2246 (O_2246,N_19843,N_19341);
or UO_2247 (O_2247,N_19604,N_19373);
xor UO_2248 (O_2248,N_19331,N_19849);
nor UO_2249 (O_2249,N_19862,N_19094);
nor UO_2250 (O_2250,N_19043,N_19699);
nor UO_2251 (O_2251,N_19241,N_19438);
and UO_2252 (O_2252,N_19902,N_19178);
nor UO_2253 (O_2253,N_19307,N_19953);
and UO_2254 (O_2254,N_19544,N_19952);
xnor UO_2255 (O_2255,N_19851,N_19569);
xor UO_2256 (O_2256,N_19582,N_19658);
and UO_2257 (O_2257,N_19951,N_19053);
and UO_2258 (O_2258,N_19776,N_19343);
or UO_2259 (O_2259,N_19698,N_19293);
or UO_2260 (O_2260,N_19119,N_19694);
xor UO_2261 (O_2261,N_19805,N_19824);
or UO_2262 (O_2262,N_19223,N_19209);
and UO_2263 (O_2263,N_19227,N_19036);
and UO_2264 (O_2264,N_19230,N_19875);
nor UO_2265 (O_2265,N_19852,N_19864);
nor UO_2266 (O_2266,N_19938,N_19808);
nand UO_2267 (O_2267,N_19094,N_19440);
xnor UO_2268 (O_2268,N_19276,N_19466);
and UO_2269 (O_2269,N_19365,N_19698);
or UO_2270 (O_2270,N_19428,N_19093);
and UO_2271 (O_2271,N_19600,N_19591);
and UO_2272 (O_2272,N_19201,N_19091);
and UO_2273 (O_2273,N_19520,N_19657);
xnor UO_2274 (O_2274,N_19658,N_19538);
xor UO_2275 (O_2275,N_19268,N_19706);
xor UO_2276 (O_2276,N_19711,N_19913);
nor UO_2277 (O_2277,N_19890,N_19183);
or UO_2278 (O_2278,N_19030,N_19997);
nor UO_2279 (O_2279,N_19929,N_19505);
xor UO_2280 (O_2280,N_19777,N_19561);
or UO_2281 (O_2281,N_19425,N_19457);
nor UO_2282 (O_2282,N_19847,N_19330);
nor UO_2283 (O_2283,N_19385,N_19057);
xnor UO_2284 (O_2284,N_19833,N_19588);
nor UO_2285 (O_2285,N_19362,N_19466);
nor UO_2286 (O_2286,N_19031,N_19512);
xor UO_2287 (O_2287,N_19757,N_19751);
or UO_2288 (O_2288,N_19085,N_19712);
xor UO_2289 (O_2289,N_19134,N_19061);
or UO_2290 (O_2290,N_19845,N_19874);
xnor UO_2291 (O_2291,N_19872,N_19167);
or UO_2292 (O_2292,N_19860,N_19394);
and UO_2293 (O_2293,N_19238,N_19803);
or UO_2294 (O_2294,N_19982,N_19543);
and UO_2295 (O_2295,N_19137,N_19941);
xor UO_2296 (O_2296,N_19551,N_19454);
nor UO_2297 (O_2297,N_19159,N_19219);
xnor UO_2298 (O_2298,N_19252,N_19356);
nand UO_2299 (O_2299,N_19775,N_19405);
nor UO_2300 (O_2300,N_19271,N_19593);
or UO_2301 (O_2301,N_19716,N_19684);
xor UO_2302 (O_2302,N_19113,N_19835);
nor UO_2303 (O_2303,N_19470,N_19029);
nand UO_2304 (O_2304,N_19833,N_19679);
nand UO_2305 (O_2305,N_19669,N_19308);
or UO_2306 (O_2306,N_19634,N_19607);
xor UO_2307 (O_2307,N_19517,N_19664);
nor UO_2308 (O_2308,N_19146,N_19014);
nor UO_2309 (O_2309,N_19138,N_19463);
or UO_2310 (O_2310,N_19456,N_19931);
nand UO_2311 (O_2311,N_19928,N_19663);
xnor UO_2312 (O_2312,N_19085,N_19544);
and UO_2313 (O_2313,N_19313,N_19830);
or UO_2314 (O_2314,N_19127,N_19704);
nand UO_2315 (O_2315,N_19617,N_19221);
and UO_2316 (O_2316,N_19586,N_19580);
xor UO_2317 (O_2317,N_19322,N_19255);
xnor UO_2318 (O_2318,N_19175,N_19835);
nand UO_2319 (O_2319,N_19553,N_19205);
nor UO_2320 (O_2320,N_19873,N_19840);
or UO_2321 (O_2321,N_19462,N_19509);
and UO_2322 (O_2322,N_19318,N_19810);
and UO_2323 (O_2323,N_19877,N_19599);
nor UO_2324 (O_2324,N_19652,N_19668);
xnor UO_2325 (O_2325,N_19747,N_19105);
or UO_2326 (O_2326,N_19893,N_19091);
or UO_2327 (O_2327,N_19936,N_19869);
xnor UO_2328 (O_2328,N_19923,N_19864);
and UO_2329 (O_2329,N_19263,N_19764);
and UO_2330 (O_2330,N_19483,N_19923);
xor UO_2331 (O_2331,N_19875,N_19683);
nor UO_2332 (O_2332,N_19424,N_19994);
and UO_2333 (O_2333,N_19313,N_19095);
nand UO_2334 (O_2334,N_19616,N_19747);
or UO_2335 (O_2335,N_19092,N_19994);
nor UO_2336 (O_2336,N_19301,N_19760);
nand UO_2337 (O_2337,N_19211,N_19984);
nor UO_2338 (O_2338,N_19090,N_19552);
xnor UO_2339 (O_2339,N_19298,N_19020);
nand UO_2340 (O_2340,N_19960,N_19537);
nand UO_2341 (O_2341,N_19942,N_19964);
nor UO_2342 (O_2342,N_19170,N_19213);
nand UO_2343 (O_2343,N_19184,N_19757);
xor UO_2344 (O_2344,N_19456,N_19638);
nor UO_2345 (O_2345,N_19817,N_19340);
nand UO_2346 (O_2346,N_19714,N_19718);
nor UO_2347 (O_2347,N_19487,N_19170);
or UO_2348 (O_2348,N_19677,N_19643);
and UO_2349 (O_2349,N_19432,N_19830);
and UO_2350 (O_2350,N_19664,N_19106);
or UO_2351 (O_2351,N_19057,N_19555);
or UO_2352 (O_2352,N_19216,N_19674);
and UO_2353 (O_2353,N_19256,N_19599);
xnor UO_2354 (O_2354,N_19148,N_19971);
nand UO_2355 (O_2355,N_19007,N_19553);
nand UO_2356 (O_2356,N_19523,N_19691);
or UO_2357 (O_2357,N_19150,N_19038);
nor UO_2358 (O_2358,N_19334,N_19741);
nand UO_2359 (O_2359,N_19679,N_19358);
and UO_2360 (O_2360,N_19277,N_19885);
and UO_2361 (O_2361,N_19575,N_19081);
and UO_2362 (O_2362,N_19527,N_19364);
nor UO_2363 (O_2363,N_19091,N_19012);
and UO_2364 (O_2364,N_19248,N_19568);
and UO_2365 (O_2365,N_19259,N_19854);
nand UO_2366 (O_2366,N_19731,N_19364);
xnor UO_2367 (O_2367,N_19901,N_19272);
and UO_2368 (O_2368,N_19069,N_19805);
or UO_2369 (O_2369,N_19339,N_19732);
nor UO_2370 (O_2370,N_19416,N_19932);
nor UO_2371 (O_2371,N_19462,N_19007);
nand UO_2372 (O_2372,N_19974,N_19375);
or UO_2373 (O_2373,N_19420,N_19595);
and UO_2374 (O_2374,N_19577,N_19524);
and UO_2375 (O_2375,N_19887,N_19784);
nand UO_2376 (O_2376,N_19705,N_19576);
and UO_2377 (O_2377,N_19910,N_19155);
and UO_2378 (O_2378,N_19019,N_19818);
nor UO_2379 (O_2379,N_19840,N_19304);
nand UO_2380 (O_2380,N_19499,N_19182);
or UO_2381 (O_2381,N_19699,N_19696);
xor UO_2382 (O_2382,N_19801,N_19044);
nor UO_2383 (O_2383,N_19912,N_19774);
or UO_2384 (O_2384,N_19942,N_19035);
nand UO_2385 (O_2385,N_19342,N_19814);
nor UO_2386 (O_2386,N_19376,N_19543);
xnor UO_2387 (O_2387,N_19608,N_19392);
and UO_2388 (O_2388,N_19917,N_19297);
xnor UO_2389 (O_2389,N_19931,N_19750);
nor UO_2390 (O_2390,N_19441,N_19949);
nor UO_2391 (O_2391,N_19520,N_19142);
or UO_2392 (O_2392,N_19057,N_19651);
xor UO_2393 (O_2393,N_19887,N_19501);
xor UO_2394 (O_2394,N_19038,N_19169);
nor UO_2395 (O_2395,N_19620,N_19249);
nand UO_2396 (O_2396,N_19315,N_19235);
xnor UO_2397 (O_2397,N_19220,N_19534);
nand UO_2398 (O_2398,N_19405,N_19324);
xor UO_2399 (O_2399,N_19234,N_19003);
xnor UO_2400 (O_2400,N_19955,N_19183);
and UO_2401 (O_2401,N_19001,N_19077);
or UO_2402 (O_2402,N_19550,N_19577);
and UO_2403 (O_2403,N_19432,N_19814);
nor UO_2404 (O_2404,N_19071,N_19472);
and UO_2405 (O_2405,N_19894,N_19656);
or UO_2406 (O_2406,N_19724,N_19501);
nor UO_2407 (O_2407,N_19457,N_19460);
and UO_2408 (O_2408,N_19876,N_19662);
xnor UO_2409 (O_2409,N_19048,N_19783);
and UO_2410 (O_2410,N_19852,N_19758);
xor UO_2411 (O_2411,N_19466,N_19779);
or UO_2412 (O_2412,N_19649,N_19530);
or UO_2413 (O_2413,N_19708,N_19837);
xnor UO_2414 (O_2414,N_19138,N_19889);
nand UO_2415 (O_2415,N_19151,N_19047);
xnor UO_2416 (O_2416,N_19786,N_19739);
or UO_2417 (O_2417,N_19113,N_19326);
xor UO_2418 (O_2418,N_19907,N_19308);
xnor UO_2419 (O_2419,N_19610,N_19063);
nand UO_2420 (O_2420,N_19526,N_19915);
nor UO_2421 (O_2421,N_19039,N_19221);
nand UO_2422 (O_2422,N_19562,N_19423);
or UO_2423 (O_2423,N_19995,N_19004);
and UO_2424 (O_2424,N_19680,N_19676);
and UO_2425 (O_2425,N_19151,N_19165);
nor UO_2426 (O_2426,N_19097,N_19791);
and UO_2427 (O_2427,N_19652,N_19573);
or UO_2428 (O_2428,N_19546,N_19053);
and UO_2429 (O_2429,N_19206,N_19762);
nand UO_2430 (O_2430,N_19425,N_19396);
nand UO_2431 (O_2431,N_19043,N_19469);
nand UO_2432 (O_2432,N_19547,N_19722);
xnor UO_2433 (O_2433,N_19961,N_19142);
nor UO_2434 (O_2434,N_19888,N_19552);
and UO_2435 (O_2435,N_19677,N_19124);
and UO_2436 (O_2436,N_19074,N_19262);
and UO_2437 (O_2437,N_19060,N_19888);
or UO_2438 (O_2438,N_19903,N_19351);
nand UO_2439 (O_2439,N_19615,N_19416);
nor UO_2440 (O_2440,N_19983,N_19980);
nor UO_2441 (O_2441,N_19824,N_19533);
xnor UO_2442 (O_2442,N_19197,N_19729);
and UO_2443 (O_2443,N_19023,N_19323);
nand UO_2444 (O_2444,N_19549,N_19930);
nand UO_2445 (O_2445,N_19788,N_19592);
or UO_2446 (O_2446,N_19288,N_19757);
or UO_2447 (O_2447,N_19377,N_19334);
nor UO_2448 (O_2448,N_19282,N_19876);
nand UO_2449 (O_2449,N_19779,N_19324);
or UO_2450 (O_2450,N_19650,N_19284);
or UO_2451 (O_2451,N_19402,N_19926);
and UO_2452 (O_2452,N_19443,N_19512);
nor UO_2453 (O_2453,N_19707,N_19659);
or UO_2454 (O_2454,N_19322,N_19917);
nor UO_2455 (O_2455,N_19039,N_19458);
xor UO_2456 (O_2456,N_19718,N_19003);
xor UO_2457 (O_2457,N_19692,N_19808);
nand UO_2458 (O_2458,N_19012,N_19487);
or UO_2459 (O_2459,N_19416,N_19610);
xor UO_2460 (O_2460,N_19569,N_19695);
nand UO_2461 (O_2461,N_19729,N_19898);
and UO_2462 (O_2462,N_19303,N_19400);
nand UO_2463 (O_2463,N_19412,N_19906);
nand UO_2464 (O_2464,N_19966,N_19406);
and UO_2465 (O_2465,N_19038,N_19219);
nand UO_2466 (O_2466,N_19704,N_19219);
or UO_2467 (O_2467,N_19779,N_19575);
xor UO_2468 (O_2468,N_19887,N_19557);
xnor UO_2469 (O_2469,N_19364,N_19048);
nor UO_2470 (O_2470,N_19816,N_19645);
or UO_2471 (O_2471,N_19340,N_19149);
or UO_2472 (O_2472,N_19624,N_19093);
and UO_2473 (O_2473,N_19360,N_19794);
nand UO_2474 (O_2474,N_19226,N_19826);
nor UO_2475 (O_2475,N_19368,N_19491);
nor UO_2476 (O_2476,N_19290,N_19209);
and UO_2477 (O_2477,N_19024,N_19481);
nand UO_2478 (O_2478,N_19860,N_19500);
nand UO_2479 (O_2479,N_19159,N_19777);
nor UO_2480 (O_2480,N_19806,N_19860);
or UO_2481 (O_2481,N_19302,N_19947);
nor UO_2482 (O_2482,N_19640,N_19838);
and UO_2483 (O_2483,N_19814,N_19288);
nand UO_2484 (O_2484,N_19703,N_19060);
nand UO_2485 (O_2485,N_19560,N_19488);
nand UO_2486 (O_2486,N_19814,N_19347);
or UO_2487 (O_2487,N_19151,N_19366);
nand UO_2488 (O_2488,N_19679,N_19123);
xor UO_2489 (O_2489,N_19032,N_19607);
and UO_2490 (O_2490,N_19948,N_19832);
xor UO_2491 (O_2491,N_19637,N_19008);
nor UO_2492 (O_2492,N_19117,N_19006);
nor UO_2493 (O_2493,N_19338,N_19146);
and UO_2494 (O_2494,N_19080,N_19981);
nor UO_2495 (O_2495,N_19064,N_19832);
nor UO_2496 (O_2496,N_19427,N_19022);
xor UO_2497 (O_2497,N_19961,N_19898);
and UO_2498 (O_2498,N_19245,N_19701);
and UO_2499 (O_2499,N_19982,N_19360);
endmodule