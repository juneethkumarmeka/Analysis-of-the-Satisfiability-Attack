module basic_1500_15000_2000_15_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_1083,In_171);
nand U1 (N_1,In_815,In_1317);
xnor U2 (N_2,In_1047,In_1475);
or U3 (N_3,In_796,In_872);
and U4 (N_4,In_315,In_264);
and U5 (N_5,In_172,In_323);
or U6 (N_6,In_1232,In_333);
nor U7 (N_7,In_1128,In_1145);
nor U8 (N_8,In_257,In_554);
and U9 (N_9,In_318,In_115);
nand U10 (N_10,In_392,In_447);
xnor U11 (N_11,In_1339,In_1235);
nor U12 (N_12,In_837,In_929);
xnor U13 (N_13,In_375,In_520);
and U14 (N_14,In_1064,In_1291);
or U15 (N_15,In_1476,In_985);
and U16 (N_16,In_640,In_1039);
xor U17 (N_17,In_1237,In_618);
or U18 (N_18,In_442,In_561);
nor U19 (N_19,In_1321,In_1377);
xor U20 (N_20,In_641,In_453);
nor U21 (N_21,In_804,In_384);
and U22 (N_22,In_55,In_776);
and U23 (N_23,In_125,In_998);
xnor U24 (N_24,In_911,In_105);
nor U25 (N_25,In_1286,In_200);
nand U26 (N_26,In_69,In_1497);
nor U27 (N_27,In_1161,In_143);
and U28 (N_28,In_361,In_879);
nor U29 (N_29,In_1385,In_622);
xnor U30 (N_30,In_819,In_619);
nor U31 (N_31,In_512,In_1263);
nor U32 (N_32,In_459,In_1439);
xor U33 (N_33,In_445,In_136);
nand U34 (N_34,In_247,In_405);
nand U35 (N_35,In_1487,In_614);
nor U36 (N_36,In_1103,In_224);
nand U37 (N_37,In_1437,In_100);
nor U38 (N_38,In_962,In_1372);
xor U39 (N_39,In_1243,In_83);
and U40 (N_40,In_904,In_1096);
and U41 (N_41,In_1347,In_436);
nand U42 (N_42,In_893,In_1044);
and U43 (N_43,In_133,In_429);
or U44 (N_44,In_861,In_1416);
and U45 (N_45,In_811,In_1203);
or U46 (N_46,In_424,In_580);
and U47 (N_47,In_1113,In_1087);
nor U48 (N_48,In_944,In_1197);
or U49 (N_49,In_282,In_868);
nor U50 (N_50,In_1228,In_1020);
or U51 (N_51,In_949,In_1117);
nor U52 (N_52,In_588,In_1373);
xor U53 (N_53,In_1125,In_1015);
xnor U54 (N_54,In_150,In_1411);
xnor U55 (N_55,In_87,In_1054);
xnor U56 (N_56,In_832,In_945);
nand U57 (N_57,In_1436,In_1010);
xnor U58 (N_58,In_543,In_1362);
and U59 (N_59,In_1366,In_1075);
and U60 (N_60,In_369,In_702);
nor U61 (N_61,In_704,In_5);
nand U62 (N_62,In_178,In_1495);
nand U63 (N_63,In_542,In_1481);
xor U64 (N_64,In_1443,In_1383);
and U65 (N_65,In_102,In_1360);
nor U66 (N_66,In_1223,In_350);
or U67 (N_67,In_517,In_711);
nor U68 (N_68,In_1494,In_1143);
or U69 (N_69,In_357,In_1297);
or U70 (N_70,In_1406,In_1488);
or U71 (N_71,In_97,In_1204);
nand U72 (N_72,In_1049,In_1420);
or U73 (N_73,In_283,In_823);
nor U74 (N_74,In_808,In_791);
or U75 (N_75,In_27,In_403);
and U76 (N_76,In_267,In_1472);
xor U77 (N_77,In_1303,In_840);
nand U78 (N_78,In_714,In_336);
nand U79 (N_79,In_570,In_431);
xnor U80 (N_80,In_862,In_662);
or U81 (N_81,In_980,In_84);
nand U82 (N_82,In_498,In_466);
nand U83 (N_83,In_1335,In_1169);
and U84 (N_84,In_216,In_1449);
or U85 (N_85,In_807,In_434);
nor U86 (N_86,In_1340,In_1478);
xor U87 (N_87,In_1455,In_635);
nand U88 (N_88,In_907,In_217);
xnor U89 (N_89,In_733,In_1329);
nor U90 (N_90,In_644,In_1273);
xnor U91 (N_91,In_93,In_1060);
or U92 (N_92,In_365,In_667);
and U93 (N_93,In_1392,In_956);
nand U94 (N_94,In_1191,In_1283);
or U95 (N_95,In_1162,In_404);
and U96 (N_96,In_1133,In_1301);
or U97 (N_97,In_731,In_65);
nor U98 (N_98,In_457,In_249);
nand U99 (N_99,In_600,In_1230);
nand U100 (N_100,In_1208,In_1043);
and U101 (N_101,In_555,In_737);
and U102 (N_102,In_747,In_1042);
and U103 (N_103,In_510,In_423);
or U104 (N_104,In_1390,In_825);
nor U105 (N_105,In_1142,In_699);
and U106 (N_106,In_829,In_210);
nand U107 (N_107,In_1129,In_1241);
or U108 (N_108,In_661,In_793);
nand U109 (N_109,In_158,In_354);
xnor U110 (N_110,In_279,In_854);
nand U111 (N_111,In_1287,In_687);
nor U112 (N_112,In_877,In_259);
nor U113 (N_113,In_697,In_340);
nand U114 (N_114,In_508,In_1171);
nand U115 (N_115,In_846,In_1355);
and U116 (N_116,In_500,In_1393);
nand U117 (N_117,In_1192,In_986);
nor U118 (N_118,In_1052,In_203);
or U119 (N_119,In_1121,In_666);
nor U120 (N_120,In_652,In_408);
nor U121 (N_121,In_1423,In_473);
or U122 (N_122,In_1115,In_1483);
nor U123 (N_123,In_491,In_1177);
or U124 (N_124,In_1207,In_299);
or U125 (N_125,In_1091,In_214);
xor U126 (N_126,In_251,In_947);
nand U127 (N_127,In_397,In_430);
xor U128 (N_128,In_530,In_1220);
or U129 (N_129,In_677,In_1082);
nand U130 (N_130,In_694,In_566);
xnor U131 (N_131,In_1299,In_730);
nor U132 (N_132,In_1012,In_1030);
nand U133 (N_133,In_858,In_799);
and U134 (N_134,In_161,In_1343);
or U135 (N_135,In_1410,In_191);
nor U136 (N_136,In_876,In_1247);
or U137 (N_137,In_114,In_1099);
nor U138 (N_138,In_1338,In_806);
and U139 (N_139,In_253,In_1092);
and U140 (N_140,In_831,In_1007);
or U141 (N_141,In_673,In_426);
and U142 (N_142,In_1137,In_464);
nor U143 (N_143,In_1023,In_612);
xor U144 (N_144,In_1489,In_707);
xor U145 (N_145,In_513,In_295);
nand U146 (N_146,In_1306,In_1492);
and U147 (N_147,In_1069,In_935);
nand U148 (N_148,In_304,In_1305);
nor U149 (N_149,In_889,In_668);
xor U150 (N_150,In_581,In_376);
xnor U151 (N_151,In_1394,In_212);
xor U152 (N_152,In_1370,In_119);
xnor U153 (N_153,In_1460,In_723);
xor U154 (N_154,In_435,In_422);
nand U155 (N_155,In_589,In_310);
and U156 (N_156,In_79,In_1289);
and U157 (N_157,In_263,In_71);
or U158 (N_158,In_1031,In_772);
nand U159 (N_159,In_739,In_111);
xor U160 (N_160,In_122,In_803);
and U161 (N_161,In_1359,In_497);
and U162 (N_162,In_242,In_965);
and U163 (N_163,In_785,In_594);
and U164 (N_164,In_1149,In_738);
and U165 (N_165,In_269,In_1139);
nor U166 (N_166,In_932,In_951);
xor U167 (N_167,In_1018,In_1);
nor U168 (N_168,In_607,In_827);
xor U169 (N_169,In_1496,In_875);
nand U170 (N_170,In_625,In_1326);
and U171 (N_171,In_678,In_533);
and U172 (N_172,In_1259,In_950);
xor U173 (N_173,In_712,In_1063);
and U174 (N_174,In_1098,In_1395);
nor U175 (N_175,In_693,In_1413);
xnor U176 (N_176,In_1477,In_984);
nand U177 (N_177,In_1210,In_1490);
or U178 (N_178,In_628,In_782);
and U179 (N_179,In_1140,In_33);
or U180 (N_180,In_227,In_732);
xor U181 (N_181,In_1308,In_123);
nand U182 (N_182,In_639,In_703);
xor U183 (N_183,In_49,In_196);
nand U184 (N_184,In_1111,In_812);
nor U185 (N_185,In_176,In_281);
nor U186 (N_186,In_1053,In_1095);
and U187 (N_187,In_1222,In_349);
or U188 (N_188,In_623,In_1256);
xnor U189 (N_189,In_331,In_1364);
nand U190 (N_190,In_124,In_1186);
nand U191 (N_191,In_983,In_1499);
or U192 (N_192,In_298,In_483);
and U193 (N_193,In_1467,In_82);
nand U194 (N_194,In_94,In_1403);
and U195 (N_195,In_103,In_725);
and U196 (N_196,In_213,In_1310);
nand U197 (N_197,In_547,In_348);
nand U198 (N_198,In_1456,In_710);
and U199 (N_199,In_1267,In_132);
xnor U200 (N_200,In_1131,In_345);
and U201 (N_201,In_407,In_314);
nand U202 (N_202,In_1132,In_1365);
nand U203 (N_203,In_149,In_767);
xor U204 (N_204,In_917,In_624);
and U205 (N_205,In_891,In_1036);
nand U206 (N_206,In_140,In_1397);
nor U207 (N_207,In_833,In_1122);
nand U208 (N_208,In_326,In_335);
xnor U209 (N_209,In_910,In_768);
nor U210 (N_210,In_748,In_494);
xor U211 (N_211,In_964,In_866);
xor U212 (N_212,In_1073,In_1251);
nand U213 (N_213,In_599,In_409);
nor U214 (N_214,In_1320,In_47);
or U215 (N_215,In_1022,In_481);
nor U216 (N_216,In_1454,In_1041);
xor U217 (N_217,In_617,In_557);
nand U218 (N_218,In_1334,In_39);
xor U219 (N_219,In_851,In_38);
or U220 (N_220,In_895,In_52);
nor U221 (N_221,In_1302,In_110);
and U222 (N_222,In_709,In_615);
or U223 (N_223,In_156,In_1175);
nand U224 (N_224,In_1120,In_1071);
or U225 (N_225,In_523,In_745);
nor U226 (N_226,In_129,In_208);
xor U227 (N_227,In_443,In_465);
nand U228 (N_228,In_237,In_1101);
and U229 (N_229,In_234,In_1061);
nor U230 (N_230,In_387,In_1389);
xnor U231 (N_231,In_118,In_1024);
xor U232 (N_232,In_954,In_669);
nor U233 (N_233,In_476,In_1382);
nor U234 (N_234,In_108,In_230);
xnor U235 (N_235,In_1470,In_1005);
or U236 (N_236,In_721,In_922);
and U237 (N_237,In_1166,In_585);
nand U238 (N_238,In_1266,In_353);
nor U239 (N_239,In_413,In_1038);
or U240 (N_240,In_660,In_941);
xnor U241 (N_241,In_255,In_386);
xnor U242 (N_242,In_696,In_924);
xnor U243 (N_243,In_1376,In_301);
nor U244 (N_244,In_968,In_814);
xor U245 (N_245,In_990,In_981);
and U246 (N_246,In_682,In_1248);
or U247 (N_247,In_629,In_309);
xnor U248 (N_248,In_416,In_1438);
xnor U249 (N_249,In_1182,In_943);
or U250 (N_250,In_1067,In_1179);
and U251 (N_251,In_648,In_1013);
or U252 (N_252,In_1086,In_233);
nor U253 (N_253,In_290,In_254);
xor U254 (N_254,In_193,In_953);
nand U255 (N_255,In_421,In_395);
xor U256 (N_256,In_1311,In_653);
or U257 (N_257,In_797,In_1379);
or U258 (N_258,In_313,In_1414);
nor U259 (N_259,In_1001,In_1158);
nand U260 (N_260,In_32,In_72);
xor U261 (N_261,In_439,In_926);
nand U262 (N_262,In_189,In_463);
nor U263 (N_263,In_1292,In_571);
xnor U264 (N_264,In_1484,In_544);
and U265 (N_265,In_1019,In_284);
or U266 (N_266,In_724,In_142);
nor U267 (N_267,In_1336,In_1211);
or U268 (N_268,In_920,In_502);
nor U269 (N_269,In_425,In_857);
nand U270 (N_270,In_1349,In_1037);
xor U271 (N_271,In_906,In_1107);
or U272 (N_272,In_14,In_278);
nor U273 (N_273,In_1108,In_402);
and U274 (N_274,In_1380,In_801);
nor U275 (N_275,In_444,In_974);
nor U276 (N_276,In_346,In_1350);
nand U277 (N_277,In_221,In_1065);
or U278 (N_278,In_1363,In_437);
nor U279 (N_279,In_592,In_275);
xnor U280 (N_280,In_378,In_680);
xnor U281 (N_281,In_865,In_1000);
and U282 (N_282,In_265,In_1090);
or U283 (N_283,In_164,In_1188);
and U284 (N_284,In_1459,In_238);
nand U285 (N_285,In_51,In_1109);
xor U286 (N_286,In_287,In_764);
or U287 (N_287,In_244,In_1400);
and U288 (N_288,In_1447,In_1035);
nor U289 (N_289,In_1221,In_205);
xnor U290 (N_290,In_900,In_993);
nand U291 (N_291,In_1268,In_449);
and U292 (N_292,In_976,In_537);
or U293 (N_293,In_1205,In_43);
nor U294 (N_294,In_828,In_139);
nor U295 (N_295,In_564,In_12);
and U296 (N_296,In_185,In_899);
or U297 (N_297,In_236,In_1144);
nand U298 (N_298,In_163,In_415);
or U299 (N_299,In_360,In_1167);
nand U300 (N_300,In_104,In_428);
or U301 (N_301,In_740,In_228);
nor U302 (N_302,In_198,In_96);
xor U303 (N_303,In_177,In_367);
xor U304 (N_304,In_1159,In_1183);
nor U305 (N_305,In_760,In_190);
nor U306 (N_306,In_207,In_595);
nand U307 (N_307,In_705,In_506);
nand U308 (N_308,In_1319,In_881);
xor U309 (N_309,In_509,In_266);
nand U310 (N_310,In_209,In_1401);
nor U311 (N_311,In_305,In_1451);
or U312 (N_312,In_23,In_64);
or U313 (N_313,In_897,In_490);
and U314 (N_314,In_252,In_487);
xnor U315 (N_315,In_596,In_1441);
nor U316 (N_316,In_560,In_713);
or U317 (N_317,In_591,In_590);
nor U318 (N_318,In_182,In_141);
nand U319 (N_319,In_432,In_671);
nand U320 (N_320,In_1025,In_778);
or U321 (N_321,In_843,In_1050);
nor U322 (N_322,In_321,In_276);
nand U323 (N_323,In_1076,In_1016);
nand U324 (N_324,In_95,In_180);
nor U325 (N_325,In_1316,In_1246);
or U326 (N_326,In_874,In_729);
xor U327 (N_327,In_59,In_853);
nand U328 (N_328,In_126,In_1402);
nand U329 (N_329,In_414,In_138);
xnor U330 (N_330,In_1262,In_885);
and U331 (N_331,In_572,In_1146);
nand U332 (N_332,In_960,In_836);
nor U333 (N_333,In_1242,In_385);
xor U334 (N_334,In_446,In_145);
or U335 (N_335,In_1479,In_90);
xnor U336 (N_336,In_1432,In_363);
nor U337 (N_337,In_685,In_440);
xor U338 (N_338,In_10,In_582);
or U339 (N_339,In_1165,In_1045);
nor U340 (N_340,In_1127,In_219);
and U341 (N_341,In_206,In_277);
or U342 (N_342,In_1173,In_174);
nor U343 (N_343,In_720,In_849);
nand U344 (N_344,In_1431,In_1130);
and U345 (N_345,In_54,In_153);
nand U346 (N_346,In_789,In_522);
nand U347 (N_347,In_374,In_29);
xnor U348 (N_348,In_46,In_1274);
nor U349 (N_349,In_679,In_690);
nor U350 (N_350,In_1255,In_1187);
nand U351 (N_351,In_824,In_6);
and U352 (N_352,In_1427,In_741);
xnor U353 (N_353,In_1461,In_942);
nor U354 (N_354,In_137,In_1399);
nand U355 (N_355,In_400,In_1196);
nand U356 (N_356,In_996,In_536);
nand U357 (N_357,In_1253,In_1231);
nand U358 (N_358,In_1358,In_1072);
xor U359 (N_359,In_130,In_1464);
nand U360 (N_360,In_1147,In_896);
nor U361 (N_361,In_239,In_235);
xor U362 (N_362,In_525,In_790);
nor U363 (N_363,In_674,In_1298);
xnor U364 (N_364,In_1124,In_856);
xor U365 (N_365,In_651,In_553);
or U366 (N_366,In_184,In_864);
or U367 (N_367,In_240,In_609);
and U368 (N_368,In_1014,In_1004);
nand U369 (N_369,In_584,In_352);
and U370 (N_370,In_700,In_1160);
and U371 (N_371,In_496,In_1446);
nor U372 (N_372,In_1415,In_810);
nor U373 (N_373,In_1463,In_603);
or U374 (N_374,In_1276,In_394);
or U375 (N_375,In_9,In_1341);
xor U376 (N_376,In_398,In_220);
or U377 (N_377,In_98,In_1026);
xnor U378 (N_378,In_794,In_451);
xnor U379 (N_379,In_1094,In_468);
nor U380 (N_380,In_577,In_1258);
nor U381 (N_381,In_1239,In_579);
nor U382 (N_382,In_933,In_608);
xnor U383 (N_383,In_602,In_1445);
xor U384 (N_384,In_777,In_780);
nand U385 (N_385,In_692,In_759);
xor U386 (N_386,In_1138,In_746);
xnor U387 (N_387,In_977,In_68);
xor U388 (N_388,In_1354,In_638);
xor U389 (N_389,In_1429,In_955);
xnor U390 (N_390,In_531,In_1055);
xor U391 (N_391,In_527,In_519);
nand U392 (N_392,In_19,In_199);
nor U393 (N_393,In_1155,In_486);
nand U394 (N_394,In_308,In_1405);
or U395 (N_395,In_839,In_1046);
nor U396 (N_396,In_192,In_620);
nor U397 (N_397,In_576,In_616);
and U398 (N_398,In_850,In_894);
nand U399 (N_399,In_322,In_225);
xor U400 (N_400,In_967,In_860);
and U401 (N_401,In_946,In_1048);
and U402 (N_402,In_475,In_1240);
xnor U403 (N_403,In_356,In_60);
nand U404 (N_404,In_166,In_1105);
nor U405 (N_405,In_418,In_388);
nand U406 (N_406,In_146,In_514);
nand U407 (N_407,In_175,In_148);
nand U408 (N_408,In_1051,In_813);
nor U409 (N_409,In_959,In_293);
nor U410 (N_410,In_30,In_505);
nor U411 (N_411,In_1224,In_834);
nand U412 (N_412,In_67,In_1398);
nor U413 (N_413,In_358,In_871);
nand U414 (N_414,In_939,In_873);
xnor U415 (N_415,In_963,In_727);
nor U416 (N_416,In_1353,In_726);
nor U417 (N_417,In_878,In_223);
and U418 (N_418,In_545,In_1371);
xor U419 (N_419,In_307,In_7);
nor U420 (N_420,In_120,In_1056);
nor U421 (N_421,In_887,In_890);
and U422 (N_422,In_18,In_1330);
or U423 (N_423,In_1294,In_320);
nor U424 (N_424,In_155,In_1219);
nand U425 (N_425,In_1491,In_1152);
nand U426 (N_426,In_1104,In_1151);
or U427 (N_427,In_22,In_366);
or U428 (N_428,In_1245,In_1206);
nand U429 (N_429,In_11,In_165);
and U430 (N_430,In_1418,In_89);
nand U431 (N_431,In_1386,In_676);
xnor U432 (N_432,In_755,In_48);
nor U433 (N_433,In_1422,In_1327);
nor U434 (N_434,In_1284,In_50);
or U435 (N_435,In_170,In_556);
and U436 (N_436,In_324,In_948);
xnor U437 (N_437,In_1021,In_835);
and U438 (N_438,In_34,In_1227);
or U439 (N_439,In_918,In_994);
or U440 (N_440,In_672,In_681);
nor U441 (N_441,In_1011,In_575);
nand U442 (N_442,In_770,In_1028);
nor U443 (N_443,In_1323,In_135);
xor U444 (N_444,In_550,In_952);
or U445 (N_445,In_197,In_245);
nor U446 (N_446,In_45,In_495);
nand U447 (N_447,In_1332,In_325);
xnor U448 (N_448,In_1261,In_1080);
or U449 (N_449,In_1361,In_75);
and U450 (N_450,In_880,In_371);
nand U451 (N_451,In_1170,In_85);
or U452 (N_452,In_419,In_80);
nand U453 (N_453,In_21,In_1384);
nor U454 (N_454,In_817,In_913);
xnor U455 (N_455,In_567,In_106);
nand U456 (N_456,In_999,In_1199);
or U457 (N_457,In_1296,In_1181);
or U458 (N_458,In_286,In_218);
nand U459 (N_459,In_1369,In_1378);
or U460 (N_460,In_892,In_1066);
nand U461 (N_461,In_665,In_73);
xor U462 (N_462,In_92,In_1190);
or U463 (N_463,In_66,In_1184);
and U464 (N_464,In_53,In_1408);
or U465 (N_465,In_1254,In_1034);
and U466 (N_466,In_898,In_633);
nor U467 (N_467,In_152,In_455);
nor U468 (N_468,In_417,In_1176);
and U469 (N_469,In_1008,In_563);
nand U470 (N_470,In_1295,In_1412);
nand U471 (N_471,In_1313,In_396);
and U472 (N_472,In_742,In_229);
nor U473 (N_473,In_1209,In_107);
xor U474 (N_474,In_930,In_701);
nand U475 (N_475,In_1126,In_187);
xor U476 (N_476,In_698,In_663);
xnor U477 (N_477,In_593,In_383);
xor U478 (N_478,In_154,In_775);
xnor U479 (N_479,In_1356,In_1345);
xor U480 (N_480,In_695,In_774);
nor U481 (N_481,In_1387,In_478);
nor U482 (N_482,In_743,In_1304);
xor U483 (N_483,In_292,In_1156);
or U484 (N_484,In_319,In_147);
xor U485 (N_485,In_1424,In_971);
or U486 (N_486,In_691,In_606);
nand U487 (N_487,In_433,In_8);
and U488 (N_488,In_1368,In_144);
nor U489 (N_489,In_1214,In_1027);
and U490 (N_490,In_1078,In_243);
nor U491 (N_491,In_469,In_1419);
or U492 (N_492,In_40,In_393);
nand U493 (N_493,In_845,In_630);
nand U494 (N_494,In_1084,In_786);
xor U495 (N_495,In_128,In_1351);
nand U496 (N_496,In_1281,In_706);
or U497 (N_497,In_380,In_821);
xor U498 (N_498,In_484,In_485);
xor U499 (N_499,In_61,In_1217);
nor U500 (N_500,In_1265,In_1017);
nand U501 (N_501,In_1457,In_1193);
nand U502 (N_502,In_1325,In_1425);
nor U503 (N_503,In_1236,In_334);
or U504 (N_504,In_1216,In_1346);
nor U505 (N_505,In_1453,In_1277);
nand U506 (N_506,In_632,In_1272);
xor U507 (N_507,In_169,In_342);
nand U508 (N_508,In_246,In_1250);
xnor U509 (N_509,In_870,In_204);
nor U510 (N_510,In_232,In_1331);
nand U511 (N_511,In_489,In_1102);
or U512 (N_512,In_1134,In_1498);
and U513 (N_513,In_982,In_186);
and U514 (N_514,In_756,In_634);
or U515 (N_515,In_450,In_936);
xnor U516 (N_516,In_969,In_769);
and U517 (N_517,In_56,In_1079);
or U518 (N_518,In_479,In_852);
nand U519 (N_519,In_1150,In_882);
and U520 (N_520,In_461,In_830);
and U521 (N_521,In_765,In_1033);
or U522 (N_522,In_1278,In_285);
nor U523 (N_523,In_558,In_1417);
or U524 (N_524,In_1333,In_76);
xnor U525 (N_525,In_524,In_781);
nand U526 (N_526,In_645,In_1275);
nor U527 (N_527,In_1428,In_1213);
xnor U528 (N_528,In_302,In_1002);
and U529 (N_529,In_1375,In_162);
and U530 (N_530,In_250,In_1229);
and U531 (N_531,In_1433,In_751);
nand U532 (N_532,In_1391,In_816);
xnor U533 (N_533,In_534,In_1458);
or U534 (N_534,In_1081,In_241);
and U535 (N_535,In_792,In_1450);
and U536 (N_536,In_1352,In_642);
xor U537 (N_537,In_613,In_841);
and U538 (N_538,In_1348,In_116);
xnor U539 (N_539,In_1452,In_541);
nor U540 (N_540,In_659,In_631);
or U541 (N_541,In_1404,In_1480);
nand U542 (N_542,In_1314,In_1300);
nand U543 (N_543,In_1029,In_903);
nand U544 (N_544,In_372,In_159);
nor U545 (N_545,In_735,In_601);
nor U546 (N_546,In_805,In_121);
nor U547 (N_547,In_788,In_16);
and U548 (N_548,In_270,In_44);
and U549 (N_549,In_329,In_362);
and U550 (N_550,In_1136,In_1148);
and U551 (N_551,In_306,In_991);
or U552 (N_552,In_1324,In_957);
nor U553 (N_553,In_504,In_610);
or U554 (N_554,In_989,In_438);
nor U555 (N_555,In_773,In_377);
nand U556 (N_556,In_359,In_70);
and U557 (N_557,In_296,In_1178);
nand U558 (N_558,In_1116,In_1465);
nor U559 (N_559,In_1106,In_127);
nand U560 (N_560,In_1270,In_637);
xnor U561 (N_561,In_516,In_294);
and U562 (N_562,In_1466,In_507);
or U563 (N_563,In_655,In_1174);
nand U564 (N_564,In_752,In_274);
or U565 (N_565,In_1077,In_202);
and U566 (N_566,In_389,In_1068);
nor U567 (N_567,In_689,In_1238);
nand U568 (N_568,In_291,In_753);
nand U569 (N_569,In_1264,In_565);
and U570 (N_570,In_722,In_26);
xnor U571 (N_571,In_884,In_410);
xnor U572 (N_572,In_460,In_573);
and U573 (N_573,In_482,In_272);
nand U574 (N_574,In_1493,In_37);
xor U575 (N_575,In_1448,In_35);
nand U576 (N_576,In_1444,In_649);
or U577 (N_577,In_57,In_1164);
nand U578 (N_578,In_650,In_1442);
xnor U579 (N_579,In_787,In_715);
nand U580 (N_580,In_728,In_518);
or U581 (N_581,In_647,In_1468);
and U582 (N_582,In_848,In_1257);
or U583 (N_583,In_859,In_1157);
or U584 (N_584,In_1110,In_112);
nor U585 (N_585,In_62,In_343);
xnor U586 (N_586,In_919,In_934);
nor U587 (N_587,In_467,In_1342);
nor U588 (N_588,In_569,In_915);
nor U589 (N_589,In_401,In_261);
or U590 (N_590,In_195,In_493);
nand U591 (N_591,In_1234,In_717);
or U592 (N_592,In_1293,In_36);
xor U593 (N_593,In_1100,In_248);
or U594 (N_594,In_1252,In_1430);
or U595 (N_595,In_838,In_188);
xor U596 (N_596,In_355,In_1058);
and U597 (N_597,In_540,In_316);
or U598 (N_598,In_1434,In_636);
xnor U599 (N_599,In_488,In_842);
and U600 (N_600,In_1195,In_501);
xor U601 (N_601,In_975,In_312);
or U602 (N_602,In_273,In_758);
and U603 (N_603,In_179,In_961);
or U604 (N_604,In_338,In_766);
xor U605 (N_605,In_626,In_927);
xor U606 (N_606,In_916,In_88);
nand U607 (N_607,In_262,In_503);
nor U608 (N_608,In_1180,In_42);
nand U609 (N_609,In_1118,In_940);
nand U610 (N_610,In_462,In_1282);
and U611 (N_611,In_1374,In_1093);
nand U612 (N_612,In_1218,In_675);
nand U613 (N_613,In_480,In_420);
and U614 (N_614,In_587,In_1322);
nor U615 (N_615,In_1290,In_379);
or U616 (N_616,In_515,In_173);
and U617 (N_617,In_784,In_1307);
nor U618 (N_618,In_1244,In_373);
and U619 (N_619,In_351,In_1194);
nand U620 (N_620,In_972,In_1089);
nand U621 (N_621,In_492,In_1168);
and U622 (N_622,In_855,In_966);
nor U623 (N_623,In_381,In_330);
and U624 (N_624,In_1185,In_337);
or U625 (N_625,In_905,In_719);
nand U626 (N_626,In_458,In_526);
nor U627 (N_627,In_1388,In_113);
nor U628 (N_628,In_1469,In_99);
xor U629 (N_629,In_231,In_822);
and U630 (N_630,In_74,In_1440);
or U631 (N_631,In_1074,In_332);
nand U632 (N_632,In_211,In_657);
and U633 (N_633,In_260,In_1215);
nor U634 (N_634,In_280,In_686);
and U635 (N_635,In_970,In_937);
and U636 (N_636,In_406,In_474);
nand U637 (N_637,In_1153,In_901);
xor U638 (N_638,In_598,In_1271);
and U639 (N_639,In_1233,In_716);
xor U640 (N_640,In_347,In_783);
or U641 (N_641,In_448,In_1396);
nor U642 (N_642,In_1309,In_471);
nor U643 (N_643,In_194,In_988);
or U644 (N_644,In_958,In_1070);
xor U645 (N_645,In_226,In_914);
xnor U646 (N_646,In_1426,In_167);
nand U647 (N_647,In_1485,In_736);
xnor U648 (N_648,In_923,In_317);
or U649 (N_649,In_844,In_168);
or U650 (N_650,In_863,In_1226);
nor U651 (N_651,In_928,In_24);
nor U652 (N_652,In_28,In_1337);
and U653 (N_653,In_902,In_1482);
nand U654 (N_654,In_368,In_1357);
xor U655 (N_655,In_1032,In_364);
nor U656 (N_656,In_708,In_271);
xnor U657 (N_657,In_456,In_818);
xnor U658 (N_658,In_311,In_91);
nand U659 (N_659,In_546,In_222);
and U660 (N_660,In_744,In_761);
nor U661 (N_661,In_683,In_908);
nand U662 (N_662,In_763,In_552);
xor U663 (N_663,In_303,In_912);
nand U664 (N_664,In_562,In_869);
or U665 (N_665,In_798,In_1367);
nand U666 (N_666,In_268,In_1285);
nand U667 (N_667,In_151,In_973);
and U668 (N_668,In_586,In_521);
nor U669 (N_669,In_1280,In_1279);
nand U670 (N_670,In_131,In_718);
and U671 (N_671,In_604,In_1003);
and U672 (N_672,In_101,In_909);
nor U673 (N_673,In_734,In_256);
xor U674 (N_674,In_1189,In_528);
xor U675 (N_675,In_551,In_134);
nor U676 (N_676,In_1202,In_1407);
nor U677 (N_677,In_1119,In_1085);
or U678 (N_678,In_13,In_297);
xor U679 (N_679,In_992,In_802);
or U680 (N_680,In_2,In_1344);
xnor U681 (N_681,In_382,In_800);
nand U682 (N_682,In_339,In_399);
xor U683 (N_683,In_809,In_627);
nand U684 (N_684,In_995,In_1114);
xor U685 (N_685,In_883,In_654);
or U686 (N_686,In_1288,In_886);
or U687 (N_687,In_921,In_341);
nand U688 (N_688,In_643,In_1088);
and U689 (N_689,In_1315,In_559);
nor U690 (N_690,In_86,In_117);
or U691 (N_691,In_472,In_548);
and U692 (N_692,In_867,In_0);
or U693 (N_693,In_452,In_3);
xnor U694 (N_694,In_17,In_670);
or U695 (N_695,In_762,In_529);
or U696 (N_696,In_1486,In_757);
xor U697 (N_697,In_1471,In_1006);
nand U698 (N_698,In_539,In_1009);
xnor U699 (N_699,In_183,In_1201);
nor U700 (N_700,In_412,In_31);
nand U701 (N_701,In_81,In_499);
or U702 (N_702,In_201,In_344);
xor U703 (N_703,In_289,In_454);
nand U704 (N_704,In_578,In_771);
nand U705 (N_705,In_684,In_931);
or U706 (N_706,In_1135,In_795);
and U707 (N_707,In_1328,In_925);
and U708 (N_708,In_1212,In_370);
or U709 (N_709,In_754,In_1163);
and U710 (N_710,In_820,In_656);
nor U711 (N_711,In_605,In_1057);
nand U712 (N_712,In_664,In_1462);
nor U713 (N_713,In_58,In_181);
nand U714 (N_714,In_583,In_1062);
nand U715 (N_715,In_411,In_1123);
nor U716 (N_716,In_1154,In_41);
xor U717 (N_717,In_1040,In_477);
or U718 (N_718,In_750,In_78);
nand U719 (N_719,In_1198,In_288);
or U720 (N_720,In_470,In_1112);
nand U721 (N_721,In_1059,In_1474);
nand U722 (N_722,In_511,In_888);
nand U723 (N_723,In_688,In_1473);
xnor U724 (N_724,In_1200,In_826);
and U725 (N_725,In_1318,In_25);
nor U726 (N_726,In_1097,In_1269);
nand U727 (N_727,In_77,In_532);
xnor U728 (N_728,In_109,In_847);
nand U729 (N_729,In_441,In_979);
or U730 (N_730,In_20,In_327);
xnor U731 (N_731,In_1249,In_779);
and U732 (N_732,In_427,In_574);
nor U733 (N_733,In_987,In_549);
xnor U734 (N_734,In_658,In_300);
nand U735 (N_735,In_1409,In_535);
nor U736 (N_736,In_157,In_611);
or U737 (N_737,In_997,In_15);
and U738 (N_738,In_1421,In_1312);
nor U739 (N_739,In_258,In_1260);
or U740 (N_740,In_328,In_749);
or U741 (N_741,In_621,In_1435);
nor U742 (N_742,In_4,In_1141);
nand U743 (N_743,In_160,In_538);
nand U744 (N_744,In_597,In_63);
or U745 (N_745,In_1172,In_215);
nand U746 (N_746,In_391,In_978);
and U747 (N_747,In_1225,In_390);
and U748 (N_748,In_1381,In_938);
xor U749 (N_749,In_646,In_568);
and U750 (N_750,In_224,In_395);
nand U751 (N_751,In_717,In_510);
xnor U752 (N_752,In_622,In_857);
nor U753 (N_753,In_581,In_38);
or U754 (N_754,In_1023,In_1094);
nor U755 (N_755,In_937,In_1158);
xnor U756 (N_756,In_536,In_832);
nand U757 (N_757,In_1232,In_960);
and U758 (N_758,In_11,In_1203);
xor U759 (N_759,In_71,In_128);
and U760 (N_760,In_605,In_920);
and U761 (N_761,In_548,In_673);
nand U762 (N_762,In_580,In_686);
nor U763 (N_763,In_1080,In_1087);
nor U764 (N_764,In_130,In_728);
or U765 (N_765,In_1094,In_1058);
and U766 (N_766,In_990,In_1158);
nand U767 (N_767,In_1465,In_448);
nor U768 (N_768,In_853,In_167);
xor U769 (N_769,In_531,In_284);
and U770 (N_770,In_1384,In_1451);
or U771 (N_771,In_562,In_1483);
or U772 (N_772,In_815,In_568);
xor U773 (N_773,In_14,In_624);
xor U774 (N_774,In_697,In_403);
nand U775 (N_775,In_1215,In_1185);
xor U776 (N_776,In_93,In_767);
nor U777 (N_777,In_777,In_481);
or U778 (N_778,In_559,In_1301);
xnor U779 (N_779,In_960,In_489);
xor U780 (N_780,In_557,In_1317);
nand U781 (N_781,In_753,In_1216);
nor U782 (N_782,In_1319,In_117);
xor U783 (N_783,In_872,In_1286);
nand U784 (N_784,In_150,In_1183);
or U785 (N_785,In_680,In_164);
nor U786 (N_786,In_245,In_1184);
and U787 (N_787,In_587,In_1068);
xor U788 (N_788,In_608,In_361);
nand U789 (N_789,In_10,In_292);
and U790 (N_790,In_1225,In_586);
or U791 (N_791,In_1016,In_1326);
or U792 (N_792,In_673,In_1064);
nand U793 (N_793,In_304,In_91);
xnor U794 (N_794,In_374,In_1024);
and U795 (N_795,In_507,In_88);
and U796 (N_796,In_5,In_1409);
xor U797 (N_797,In_1341,In_527);
xor U798 (N_798,In_1443,In_177);
nor U799 (N_799,In_327,In_23);
or U800 (N_800,In_1088,In_270);
nor U801 (N_801,In_248,In_418);
nand U802 (N_802,In_1087,In_1392);
nand U803 (N_803,In_709,In_600);
nor U804 (N_804,In_903,In_1336);
nor U805 (N_805,In_368,In_62);
and U806 (N_806,In_560,In_75);
xor U807 (N_807,In_539,In_28);
xor U808 (N_808,In_342,In_503);
nand U809 (N_809,In_745,In_1225);
xor U810 (N_810,In_590,In_750);
or U811 (N_811,In_517,In_1084);
nand U812 (N_812,In_416,In_1254);
nand U813 (N_813,In_81,In_1475);
nand U814 (N_814,In_638,In_1108);
or U815 (N_815,In_983,In_784);
nor U816 (N_816,In_591,In_11);
nor U817 (N_817,In_26,In_175);
or U818 (N_818,In_1232,In_610);
nor U819 (N_819,In_560,In_1461);
nor U820 (N_820,In_1475,In_1444);
and U821 (N_821,In_720,In_142);
nor U822 (N_822,In_1482,In_1322);
nand U823 (N_823,In_550,In_719);
nand U824 (N_824,In_1247,In_1349);
nor U825 (N_825,In_1498,In_52);
xnor U826 (N_826,In_453,In_317);
xnor U827 (N_827,In_247,In_662);
or U828 (N_828,In_140,In_12);
and U829 (N_829,In_1471,In_829);
nor U830 (N_830,In_1276,In_1142);
nor U831 (N_831,In_759,In_138);
nand U832 (N_832,In_289,In_828);
or U833 (N_833,In_1395,In_116);
nand U834 (N_834,In_582,In_229);
or U835 (N_835,In_1205,In_1006);
and U836 (N_836,In_28,In_1209);
and U837 (N_837,In_781,In_1265);
nand U838 (N_838,In_904,In_1429);
nand U839 (N_839,In_329,In_1341);
and U840 (N_840,In_402,In_658);
or U841 (N_841,In_77,In_1301);
nand U842 (N_842,In_235,In_72);
nand U843 (N_843,In_1238,In_0);
and U844 (N_844,In_164,In_804);
or U845 (N_845,In_1423,In_971);
nand U846 (N_846,In_222,In_6);
xnor U847 (N_847,In_88,In_1311);
or U848 (N_848,In_744,In_342);
or U849 (N_849,In_265,In_1022);
and U850 (N_850,In_702,In_1116);
nand U851 (N_851,In_553,In_755);
and U852 (N_852,In_646,In_207);
nor U853 (N_853,In_65,In_1260);
xnor U854 (N_854,In_20,In_1376);
xor U855 (N_855,In_300,In_1144);
nand U856 (N_856,In_1111,In_1043);
and U857 (N_857,In_1420,In_84);
or U858 (N_858,In_836,In_746);
nand U859 (N_859,In_827,In_794);
and U860 (N_860,In_1317,In_1202);
nor U861 (N_861,In_972,In_865);
nor U862 (N_862,In_22,In_759);
and U863 (N_863,In_875,In_422);
and U864 (N_864,In_1076,In_1039);
xor U865 (N_865,In_334,In_513);
xnor U866 (N_866,In_17,In_295);
nand U867 (N_867,In_12,In_368);
and U868 (N_868,In_16,In_451);
xnor U869 (N_869,In_937,In_59);
xor U870 (N_870,In_650,In_596);
nand U871 (N_871,In_3,In_101);
xor U872 (N_872,In_238,In_1043);
nor U873 (N_873,In_990,In_19);
and U874 (N_874,In_1124,In_573);
nor U875 (N_875,In_1463,In_1257);
xor U876 (N_876,In_781,In_446);
nor U877 (N_877,In_1377,In_535);
xnor U878 (N_878,In_758,In_1487);
xor U879 (N_879,In_584,In_563);
and U880 (N_880,In_674,In_740);
and U881 (N_881,In_1087,In_636);
nand U882 (N_882,In_78,In_1283);
and U883 (N_883,In_688,In_908);
or U884 (N_884,In_771,In_1232);
nor U885 (N_885,In_679,In_194);
and U886 (N_886,In_893,In_70);
nand U887 (N_887,In_168,In_498);
and U888 (N_888,In_1149,In_122);
nor U889 (N_889,In_597,In_857);
xnor U890 (N_890,In_572,In_576);
nand U891 (N_891,In_455,In_1284);
or U892 (N_892,In_1443,In_985);
and U893 (N_893,In_1240,In_1044);
nor U894 (N_894,In_133,In_775);
or U895 (N_895,In_411,In_166);
nor U896 (N_896,In_58,In_663);
nor U897 (N_897,In_763,In_1003);
nor U898 (N_898,In_307,In_964);
and U899 (N_899,In_271,In_580);
nand U900 (N_900,In_1111,In_232);
nand U901 (N_901,In_1171,In_1178);
nor U902 (N_902,In_1190,In_1222);
xor U903 (N_903,In_338,In_894);
or U904 (N_904,In_790,In_913);
and U905 (N_905,In_450,In_192);
nor U906 (N_906,In_423,In_207);
nor U907 (N_907,In_791,In_80);
or U908 (N_908,In_1192,In_333);
and U909 (N_909,In_1331,In_1253);
or U910 (N_910,In_1455,In_24);
nand U911 (N_911,In_646,In_1449);
xor U912 (N_912,In_269,In_1402);
or U913 (N_913,In_784,In_371);
xor U914 (N_914,In_1464,In_1007);
nand U915 (N_915,In_770,In_1044);
nor U916 (N_916,In_831,In_433);
nor U917 (N_917,In_1320,In_691);
and U918 (N_918,In_1337,In_1289);
nand U919 (N_919,In_114,In_224);
xor U920 (N_920,In_755,In_349);
nor U921 (N_921,In_477,In_377);
nor U922 (N_922,In_679,In_360);
and U923 (N_923,In_234,In_1267);
xor U924 (N_924,In_950,In_37);
or U925 (N_925,In_290,In_56);
nor U926 (N_926,In_829,In_97);
and U927 (N_927,In_824,In_1207);
or U928 (N_928,In_612,In_958);
nor U929 (N_929,In_1081,In_1252);
xor U930 (N_930,In_154,In_1488);
or U931 (N_931,In_582,In_137);
and U932 (N_932,In_606,In_565);
nand U933 (N_933,In_25,In_1338);
nand U934 (N_934,In_1172,In_1324);
xnor U935 (N_935,In_456,In_710);
nand U936 (N_936,In_702,In_782);
or U937 (N_937,In_881,In_280);
nand U938 (N_938,In_1121,In_514);
xor U939 (N_939,In_818,In_1131);
or U940 (N_940,In_1246,In_1099);
nand U941 (N_941,In_581,In_750);
xor U942 (N_942,In_398,In_980);
and U943 (N_943,In_1256,In_930);
nor U944 (N_944,In_799,In_1250);
nor U945 (N_945,In_1260,In_642);
nand U946 (N_946,In_1176,In_1356);
nor U947 (N_947,In_69,In_474);
or U948 (N_948,In_157,In_1077);
xnor U949 (N_949,In_335,In_1401);
nand U950 (N_950,In_1110,In_79);
or U951 (N_951,In_266,In_155);
nand U952 (N_952,In_1147,In_1288);
and U953 (N_953,In_1077,In_877);
nand U954 (N_954,In_1208,In_1448);
and U955 (N_955,In_1090,In_749);
or U956 (N_956,In_1442,In_1157);
nor U957 (N_957,In_147,In_158);
nand U958 (N_958,In_1119,In_130);
nand U959 (N_959,In_1340,In_1416);
nand U960 (N_960,In_1184,In_528);
and U961 (N_961,In_849,In_510);
nor U962 (N_962,In_1458,In_214);
or U963 (N_963,In_822,In_769);
nor U964 (N_964,In_249,In_836);
xnor U965 (N_965,In_687,In_274);
xor U966 (N_966,In_1163,In_1430);
nand U967 (N_967,In_1097,In_1186);
and U968 (N_968,In_999,In_617);
or U969 (N_969,In_630,In_1439);
nand U970 (N_970,In_643,In_760);
and U971 (N_971,In_795,In_986);
and U972 (N_972,In_300,In_722);
nor U973 (N_973,In_1010,In_1289);
or U974 (N_974,In_809,In_933);
nand U975 (N_975,In_283,In_1233);
xnor U976 (N_976,In_414,In_3);
nand U977 (N_977,In_999,In_365);
nor U978 (N_978,In_1415,In_1430);
xor U979 (N_979,In_676,In_76);
nor U980 (N_980,In_1160,In_1202);
nor U981 (N_981,In_1337,In_1417);
xnor U982 (N_982,In_104,In_214);
or U983 (N_983,In_577,In_1301);
xnor U984 (N_984,In_1201,In_194);
nand U985 (N_985,In_1397,In_1050);
nand U986 (N_986,In_384,In_1485);
nand U987 (N_987,In_304,In_172);
nand U988 (N_988,In_1123,In_364);
xor U989 (N_989,In_1114,In_1105);
and U990 (N_990,In_194,In_744);
and U991 (N_991,In_83,In_1441);
and U992 (N_992,In_644,In_1188);
xnor U993 (N_993,In_1340,In_82);
xnor U994 (N_994,In_461,In_1389);
nor U995 (N_995,In_833,In_820);
nand U996 (N_996,In_190,In_521);
nand U997 (N_997,In_213,In_1174);
xor U998 (N_998,In_88,In_273);
xnor U999 (N_999,In_76,In_408);
and U1000 (N_1000,N_415,N_943);
or U1001 (N_1001,N_750,N_511);
nand U1002 (N_1002,N_563,N_488);
xor U1003 (N_1003,N_895,N_594);
and U1004 (N_1004,N_773,N_208);
or U1005 (N_1005,N_637,N_199);
and U1006 (N_1006,N_356,N_619);
and U1007 (N_1007,N_880,N_770);
or U1008 (N_1008,N_794,N_400);
nand U1009 (N_1009,N_19,N_187);
and U1010 (N_1010,N_504,N_654);
and U1011 (N_1011,N_303,N_788);
nor U1012 (N_1012,N_996,N_477);
nand U1013 (N_1013,N_168,N_211);
or U1014 (N_1014,N_836,N_431);
and U1015 (N_1015,N_696,N_178);
nor U1016 (N_1016,N_159,N_130);
nor U1017 (N_1017,N_925,N_30);
xnor U1018 (N_1018,N_582,N_702);
or U1019 (N_1019,N_67,N_122);
nand U1020 (N_1020,N_737,N_331);
nand U1021 (N_1021,N_534,N_601);
and U1022 (N_1022,N_983,N_722);
nor U1023 (N_1023,N_884,N_471);
or U1024 (N_1024,N_146,N_580);
and U1025 (N_1025,N_965,N_283);
or U1026 (N_1026,N_756,N_599);
xor U1027 (N_1027,N_946,N_189);
nand U1028 (N_1028,N_430,N_721);
nand U1029 (N_1029,N_265,N_913);
and U1030 (N_1030,N_995,N_197);
or U1031 (N_1031,N_768,N_23);
or U1032 (N_1032,N_450,N_801);
nor U1033 (N_1033,N_171,N_157);
nor U1034 (N_1034,N_20,N_759);
or U1035 (N_1035,N_394,N_52);
nor U1036 (N_1036,N_490,N_334);
or U1037 (N_1037,N_395,N_120);
and U1038 (N_1038,N_893,N_495);
nor U1039 (N_1039,N_101,N_68);
xnor U1040 (N_1040,N_507,N_964);
nand U1041 (N_1041,N_418,N_644);
or U1042 (N_1042,N_41,N_290);
and U1043 (N_1043,N_322,N_5);
xnor U1044 (N_1044,N_414,N_686);
or U1045 (N_1045,N_660,N_738);
or U1046 (N_1046,N_358,N_703);
or U1047 (N_1047,N_554,N_131);
or U1048 (N_1048,N_989,N_911);
and U1049 (N_1049,N_851,N_314);
nand U1050 (N_1050,N_53,N_274);
xor U1051 (N_1051,N_466,N_917);
or U1052 (N_1052,N_147,N_976);
nor U1053 (N_1053,N_27,N_932);
nor U1054 (N_1054,N_907,N_225);
and U1055 (N_1055,N_36,N_399);
xor U1056 (N_1056,N_304,N_835);
and U1057 (N_1057,N_92,N_906);
and U1058 (N_1058,N_43,N_396);
or U1059 (N_1059,N_61,N_833);
nand U1060 (N_1060,N_695,N_849);
or U1061 (N_1061,N_842,N_612);
nor U1062 (N_1062,N_669,N_106);
nand U1063 (N_1063,N_433,N_521);
nand U1064 (N_1064,N_538,N_897);
and U1065 (N_1065,N_832,N_776);
xor U1066 (N_1066,N_295,N_866);
nor U1067 (N_1067,N_542,N_524);
or U1068 (N_1068,N_624,N_903);
nand U1069 (N_1069,N_104,N_319);
xor U1070 (N_1070,N_748,N_991);
nor U1071 (N_1071,N_997,N_522);
nand U1072 (N_1072,N_847,N_180);
nor U1073 (N_1073,N_80,N_479);
or U1074 (N_1074,N_839,N_803);
nand U1075 (N_1075,N_465,N_480);
and U1076 (N_1076,N_209,N_64);
or U1077 (N_1077,N_714,N_88);
or U1078 (N_1078,N_456,N_564);
nor U1079 (N_1079,N_69,N_55);
nor U1080 (N_1080,N_129,N_775);
nand U1081 (N_1081,N_17,N_867);
nor U1082 (N_1082,N_629,N_685);
xor U1083 (N_1083,N_39,N_975);
and U1084 (N_1084,N_8,N_416);
nand U1085 (N_1085,N_713,N_525);
or U1086 (N_1086,N_77,N_827);
or U1087 (N_1087,N_231,N_93);
or U1088 (N_1088,N_467,N_586);
nand U1089 (N_1089,N_203,N_840);
and U1090 (N_1090,N_362,N_162);
nor U1091 (N_1091,N_59,N_323);
nor U1092 (N_1092,N_992,N_901);
nor U1093 (N_1093,N_643,N_742);
nor U1094 (N_1094,N_270,N_709);
xnor U1095 (N_1095,N_710,N_165);
xnor U1096 (N_1096,N_959,N_892);
or U1097 (N_1097,N_166,N_514);
xnor U1098 (N_1098,N_60,N_325);
xor U1099 (N_1099,N_112,N_74);
nor U1100 (N_1100,N_558,N_778);
xnor U1101 (N_1101,N_54,N_349);
nand U1102 (N_1102,N_355,N_927);
or U1103 (N_1103,N_711,N_291);
and U1104 (N_1104,N_248,N_447);
xnor U1105 (N_1105,N_734,N_151);
xnor U1106 (N_1106,N_752,N_767);
or U1107 (N_1107,N_741,N_556);
nand U1108 (N_1108,N_58,N_857);
nor U1109 (N_1109,N_18,N_732);
and U1110 (N_1110,N_947,N_70);
or U1111 (N_1111,N_384,N_21);
nor U1112 (N_1112,N_366,N_571);
or U1113 (N_1113,N_215,N_13);
xor U1114 (N_1114,N_649,N_406);
xnor U1115 (N_1115,N_682,N_766);
xnor U1116 (N_1116,N_618,N_56);
nor U1117 (N_1117,N_500,N_177);
nor U1118 (N_1118,N_44,N_11);
nand U1119 (N_1119,N_754,N_850);
xor U1120 (N_1120,N_278,N_547);
and U1121 (N_1121,N_760,N_296);
or U1122 (N_1122,N_4,N_535);
or U1123 (N_1123,N_133,N_970);
nand U1124 (N_1124,N_391,N_105);
and U1125 (N_1125,N_668,N_672);
and U1126 (N_1126,N_779,N_555);
nand U1127 (N_1127,N_135,N_289);
xnor U1128 (N_1128,N_977,N_720);
nor U1129 (N_1129,N_95,N_864);
or U1130 (N_1130,N_12,N_592);
nor U1131 (N_1131,N_606,N_182);
or U1132 (N_1132,N_510,N_340);
nand U1133 (N_1133,N_985,N_883);
nor U1134 (N_1134,N_417,N_268);
xor U1135 (N_1135,N_875,N_824);
or U1136 (N_1136,N_676,N_724);
nor U1137 (N_1137,N_663,N_132);
nand U1138 (N_1138,N_730,N_320);
or U1139 (N_1139,N_587,N_518);
xor U1140 (N_1140,N_424,N_483);
nor U1141 (N_1141,N_569,N_935);
nor U1142 (N_1142,N_755,N_622);
xor U1143 (N_1143,N_276,N_853);
or U1144 (N_1144,N_621,N_223);
nand U1145 (N_1145,N_999,N_717);
xnor U1146 (N_1146,N_163,N_693);
xor U1147 (N_1147,N_715,N_308);
and U1148 (N_1148,N_256,N_688);
and U1149 (N_1149,N_46,N_214);
nor U1150 (N_1150,N_733,N_86);
and U1151 (N_1151,N_912,N_623);
xor U1152 (N_1152,N_350,N_380);
and U1153 (N_1153,N_980,N_566);
xnor U1154 (N_1154,N_607,N_657);
nor U1155 (N_1155,N_261,N_800);
nand U1156 (N_1156,N_952,N_729);
xnor U1157 (N_1157,N_786,N_889);
and U1158 (N_1158,N_899,N_352);
or U1159 (N_1159,N_597,N_367);
xnor U1160 (N_1160,N_916,N_705);
nor U1161 (N_1161,N_749,N_718);
or U1162 (N_1162,N_790,N_285);
nand U1163 (N_1163,N_813,N_793);
or U1164 (N_1164,N_653,N_236);
nand U1165 (N_1165,N_342,N_751);
nand U1166 (N_1166,N_302,N_631);
nor U1167 (N_1167,N_854,N_922);
or U1168 (N_1168,N_967,N_888);
and U1169 (N_1169,N_99,N_258);
xnor U1170 (N_1170,N_953,N_108);
or U1171 (N_1171,N_700,N_119);
nand U1172 (N_1172,N_33,N_411);
and U1173 (N_1173,N_224,N_890);
or U1174 (N_1174,N_675,N_408);
nand U1175 (N_1175,N_140,N_658);
and U1176 (N_1176,N_740,N_628);
nor U1177 (N_1177,N_89,N_255);
or U1178 (N_1178,N_206,N_110);
and U1179 (N_1179,N_817,N_924);
nand U1180 (N_1180,N_559,N_613);
xor U1181 (N_1181,N_492,N_427);
nand U1182 (N_1182,N_868,N_962);
or U1183 (N_1183,N_124,N_680);
or U1184 (N_1184,N_968,N_526);
or U1185 (N_1185,N_647,N_543);
nor U1186 (N_1186,N_532,N_611);
nor U1187 (N_1187,N_42,N_451);
nor U1188 (N_1188,N_879,N_841);
or U1189 (N_1189,N_727,N_91);
xor U1190 (N_1190,N_780,N_886);
nand U1191 (N_1191,N_377,N_15);
or U1192 (N_1192,N_26,N_200);
and U1193 (N_1193,N_550,N_527);
or U1194 (N_1194,N_798,N_869);
nor U1195 (N_1195,N_708,N_3);
nor U1196 (N_1196,N_993,N_292);
nand U1197 (N_1197,N_299,N_179);
nor U1198 (N_1198,N_218,N_50);
nand U1199 (N_1199,N_938,N_670);
or U1200 (N_1200,N_264,N_860);
xnor U1201 (N_1201,N_990,N_633);
nor U1202 (N_1202,N_142,N_681);
xnor U1203 (N_1203,N_359,N_988);
and U1204 (N_1204,N_781,N_123);
or U1205 (N_1205,N_409,N_118);
nor U1206 (N_1206,N_332,N_307);
nor U1207 (N_1207,N_245,N_808);
or U1208 (N_1208,N_152,N_82);
and U1209 (N_1209,N_160,N_29);
xor U1210 (N_1210,N_503,N_858);
or U1211 (N_1211,N_2,N_944);
and U1212 (N_1212,N_615,N_398);
nor U1213 (N_1213,N_636,N_969);
xnor U1214 (N_1214,N_329,N_448);
xor U1215 (N_1215,N_324,N_844);
and U1216 (N_1216,N_412,N_181);
or U1217 (N_1217,N_634,N_222);
xor U1218 (N_1218,N_574,N_508);
nand U1219 (N_1219,N_862,N_785);
and U1220 (N_1220,N_515,N_62);
nand U1221 (N_1221,N_470,N_317);
xnor U1222 (N_1222,N_513,N_347);
xnor U1223 (N_1223,N_247,N_48);
and U1224 (N_1224,N_425,N_143);
or U1225 (N_1225,N_812,N_297);
nand U1226 (N_1226,N_787,N_478);
nor U1227 (N_1227,N_934,N_294);
xor U1228 (N_1228,N_158,N_379);
and U1229 (N_1229,N_175,N_260);
nand U1230 (N_1230,N_589,N_83);
xnor U1231 (N_1231,N_413,N_987);
nor U1232 (N_1232,N_830,N_739);
nand U1233 (N_1233,N_281,N_172);
xor U1234 (N_1234,N_173,N_232);
nand U1235 (N_1235,N_905,N_455);
xnor U1236 (N_1236,N_777,N_441);
nor U1237 (N_1237,N_948,N_529);
nor U1238 (N_1238,N_828,N_421);
xor U1239 (N_1239,N_701,N_584);
nand U1240 (N_1240,N_114,N_116);
nand U1241 (N_1241,N_257,N_536);
and U1242 (N_1242,N_743,N_769);
nand U1243 (N_1243,N_961,N_139);
nor U1244 (N_1244,N_570,N_505);
nor U1245 (N_1245,N_7,N_63);
xor U1246 (N_1246,N_789,N_848);
nand U1247 (N_1247,N_799,N_614);
nor U1248 (N_1248,N_174,N_193);
nor U1249 (N_1249,N_354,N_533);
nor U1250 (N_1250,N_902,N_345);
nor U1251 (N_1251,N_677,N_982);
nor U1252 (N_1252,N_422,N_551);
and U1253 (N_1253,N_298,N_782);
nor U1254 (N_1254,N_665,N_90);
or U1255 (N_1255,N_545,N_861);
and U1256 (N_1256,N_994,N_809);
xnor U1257 (N_1257,N_918,N_852);
and U1258 (N_1258,N_47,N_578);
nor U1259 (N_1259,N_57,N_144);
and U1260 (N_1260,N_169,N_138);
or U1261 (N_1261,N_369,N_326);
nor U1262 (N_1262,N_954,N_188);
or U1263 (N_1263,N_929,N_242);
and U1264 (N_1264,N_195,N_98);
nor U1265 (N_1265,N_402,N_16);
and U1266 (N_1266,N_397,N_509);
or U1267 (N_1267,N_616,N_246);
nor U1268 (N_1268,N_468,N_419);
xor U1269 (N_1269,N_443,N_435);
or U1270 (N_1270,N_667,N_335);
or U1271 (N_1271,N_951,N_458);
or U1272 (N_1272,N_269,N_309);
nor U1273 (N_1273,N_609,N_339);
xor U1274 (N_1274,N_482,N_35);
and U1275 (N_1275,N_972,N_544);
and U1276 (N_1276,N_216,N_882);
or U1277 (N_1277,N_694,N_221);
and U1278 (N_1278,N_572,N_617);
nor U1279 (N_1279,N_318,N_263);
and U1280 (N_1280,N_491,N_34);
xnor U1281 (N_1281,N_440,N_386);
xor U1282 (N_1282,N_71,N_293);
nor U1283 (N_1283,N_552,N_390);
and U1284 (N_1284,N_645,N_272);
nor U1285 (N_1285,N_382,N_437);
xor U1286 (N_1286,N_337,N_473);
and U1287 (N_1287,N_300,N_568);
nand U1288 (N_1288,N_671,N_600);
or U1289 (N_1289,N_141,N_423);
and U1290 (N_1290,N_499,N_316);
nor U1291 (N_1291,N_485,N_815);
and U1292 (N_1292,N_149,N_531);
and U1293 (N_1293,N_931,N_373);
or U1294 (N_1294,N_457,N_585);
and U1295 (N_1295,N_10,N_712);
nor U1296 (N_1296,N_904,N_72);
xnor U1297 (N_1297,N_745,N_85);
nand U1298 (N_1298,N_184,N_134);
nand U1299 (N_1299,N_392,N_288);
nor U1300 (N_1300,N_1,N_333);
nand U1301 (N_1301,N_679,N_148);
nor U1302 (N_1302,N_966,N_338);
xor U1303 (N_1303,N_6,N_960);
xnor U1304 (N_1304,N_530,N_204);
and U1305 (N_1305,N_389,N_267);
nand U1306 (N_1306,N_638,N_881);
and U1307 (N_1307,N_874,N_438);
nor U1308 (N_1308,N_364,N_341);
or U1309 (N_1309,N_420,N_939);
nor U1310 (N_1310,N_220,N_872);
nor U1311 (N_1311,N_641,N_385);
and U1312 (N_1312,N_674,N_113);
nor U1313 (N_1313,N_212,N_706);
and U1314 (N_1314,N_243,N_561);
nor U1315 (N_1315,N_933,N_540);
xor U1316 (N_1316,N_845,N_576);
or U1317 (N_1317,N_176,N_648);
and U1318 (N_1318,N_0,N_981);
nor U1319 (N_1319,N_125,N_791);
nand U1320 (N_1320,N_191,N_249);
nor U1321 (N_1321,N_97,N_115);
and U1322 (N_1322,N_519,N_923);
nand U1323 (N_1323,N_460,N_481);
xor U1324 (N_1324,N_735,N_546);
xor U1325 (N_1325,N_873,N_928);
or U1326 (N_1326,N_651,N_494);
xor U1327 (N_1327,N_65,N_31);
or U1328 (N_1328,N_646,N_84);
xor U1329 (N_1329,N_446,N_956);
nor U1330 (N_1330,N_838,N_383);
nor U1331 (N_1331,N_957,N_639);
nand U1332 (N_1332,N_254,N_805);
nor U1333 (N_1333,N_426,N_940);
or U1334 (N_1334,N_971,N_156);
or U1335 (N_1335,N_161,N_25);
nand U1336 (N_1336,N_627,N_14);
nand U1337 (N_1337,N_583,N_401);
xnor U1338 (N_1338,N_719,N_823);
xnor U1339 (N_1339,N_262,N_819);
and U1340 (N_1340,N_910,N_201);
xnor U1341 (N_1341,N_567,N_445);
and U1342 (N_1342,N_153,N_774);
or U1343 (N_1343,N_655,N_235);
nand U1344 (N_1344,N_51,N_493);
or U1345 (N_1345,N_603,N_489);
or U1346 (N_1346,N_45,N_652);
nor U1347 (N_1347,N_286,N_228);
and U1348 (N_1348,N_949,N_626);
or U1349 (N_1349,N_915,N_66);
xor U1350 (N_1350,N_442,N_541);
xor U1351 (N_1351,N_94,N_136);
or U1352 (N_1352,N_363,N_170);
xnor U1353 (N_1353,N_312,N_747);
nor U1354 (N_1354,N_941,N_908);
nand U1355 (N_1355,N_829,N_871);
xor U1356 (N_1356,N_404,N_516);
xor U1357 (N_1357,N_549,N_226);
nor U1358 (N_1358,N_986,N_539);
nor U1359 (N_1359,N_818,N_374);
and U1360 (N_1360,N_461,N_353);
nor U1361 (N_1361,N_802,N_661);
or U1362 (N_1362,N_444,N_429);
xnor U1363 (N_1363,N_807,N_877);
nor U1364 (N_1364,N_311,N_327);
or U1365 (N_1365,N_496,N_371);
and U1366 (N_1366,N_79,N_831);
nor U1367 (N_1367,N_591,N_687);
nor U1368 (N_1368,N_210,N_520);
and U1369 (N_1369,N_75,N_678);
xnor U1370 (N_1370,N_692,N_32);
nand U1371 (N_1371,N_577,N_239);
nand U1372 (N_1372,N_921,N_81);
and U1373 (N_1373,N_605,N_562);
and U1374 (N_1374,N_804,N_475);
nor U1375 (N_1375,N_484,N_78);
nand U1376 (N_1376,N_487,N_764);
nor U1377 (N_1377,N_428,N_190);
nand U1378 (N_1378,N_217,N_310);
and U1379 (N_1379,N_579,N_252);
nor U1380 (N_1380,N_328,N_183);
xor U1381 (N_1381,N_771,N_234);
xor U1382 (N_1382,N_914,N_588);
and U1383 (N_1383,N_315,N_816);
xnor U1384 (N_1384,N_207,N_357);
and U1385 (N_1385,N_523,N_375);
or U1386 (N_1386,N_449,N_909);
nand U1387 (N_1387,N_313,N_103);
or U1388 (N_1388,N_271,N_744);
xor U1389 (N_1389,N_9,N_107);
or U1390 (N_1390,N_859,N_573);
nor U1391 (N_1391,N_820,N_978);
and U1392 (N_1392,N_761,N_942);
nand U1393 (N_1393,N_656,N_662);
xor U1394 (N_1394,N_673,N_900);
nor U1395 (N_1395,N_266,N_287);
and U1396 (N_1396,N_659,N_305);
nand U1397 (N_1397,N_683,N_604);
nor U1398 (N_1398,N_843,N_919);
nand U1399 (N_1399,N_878,N_233);
and U1400 (N_1400,N_301,N_891);
nand U1401 (N_1401,N_387,N_728);
nor U1402 (N_1402,N_463,N_111);
or U1403 (N_1403,N_109,N_497);
nand U1404 (N_1404,N_560,N_469);
nand U1405 (N_1405,N_811,N_725);
xor U1406 (N_1406,N_691,N_762);
nor U1407 (N_1407,N_608,N_963);
and U1408 (N_1408,N_595,N_593);
or U1409 (N_1409,N_432,N_979);
nand U1410 (N_1410,N_698,N_517);
and U1411 (N_1411,N_284,N_100);
nand U1412 (N_1412,N_229,N_640);
nor U1413 (N_1413,N_279,N_155);
and U1414 (N_1414,N_486,N_219);
and U1415 (N_1415,N_610,N_548);
and U1416 (N_1416,N_894,N_837);
nand U1417 (N_1417,N_462,N_306);
nor U1418 (N_1418,N_945,N_365);
xnor U1419 (N_1419,N_241,N_145);
nand U1420 (N_1420,N_635,N_783);
nor U1421 (N_1421,N_958,N_821);
nand U1422 (N_1422,N_277,N_506);
xnor U1423 (N_1423,N_253,N_453);
nand U1424 (N_1424,N_650,N_664);
nor U1425 (N_1425,N_117,N_336);
or U1426 (N_1426,N_378,N_575);
xor U1427 (N_1427,N_185,N_796);
nand U1428 (N_1428,N_73,N_826);
or U1429 (N_1429,N_454,N_863);
nand U1430 (N_1430,N_590,N_330);
and U1431 (N_1431,N_96,N_403);
or U1432 (N_1432,N_49,N_726);
nand U1433 (N_1433,N_393,N_855);
nor U1434 (N_1434,N_846,N_885);
or U1435 (N_1435,N_361,N_689);
or U1436 (N_1436,N_128,N_360);
and U1437 (N_1437,N_707,N_273);
xnor U1438 (N_1438,N_666,N_464);
and U1439 (N_1439,N_684,N_557);
xnor U1440 (N_1440,N_930,N_474);
nor U1441 (N_1441,N_596,N_126);
nor U1442 (N_1442,N_731,N_434);
nand U1443 (N_1443,N_955,N_876);
nand U1444 (N_1444,N_410,N_280);
nor U1445 (N_1445,N_772,N_810);
xor U1446 (N_1446,N_381,N_736);
nor U1447 (N_1447,N_723,N_870);
xor U1448 (N_1448,N_512,N_87);
and U1449 (N_1449,N_194,N_28);
and U1450 (N_1450,N_984,N_690);
xnor U1451 (N_1451,N_202,N_537);
nor U1452 (N_1452,N_763,N_405);
nor U1453 (N_1453,N_38,N_472);
xor U1454 (N_1454,N_630,N_372);
or U1455 (N_1455,N_244,N_602);
and U1456 (N_1456,N_37,N_150);
xor U1457 (N_1457,N_825,N_237);
nor U1458 (N_1458,N_76,N_40);
xor U1459 (N_1459,N_822,N_344);
nor U1460 (N_1460,N_565,N_502);
and U1461 (N_1461,N_973,N_581);
xnor U1462 (N_1462,N_898,N_407);
or U1463 (N_1463,N_758,N_368);
nand U1464 (N_1464,N_321,N_998);
nand U1465 (N_1465,N_282,N_24);
and U1466 (N_1466,N_501,N_797);
xnor U1467 (N_1467,N_834,N_167);
or U1468 (N_1468,N_865,N_137);
nor U1469 (N_1469,N_498,N_598);
nand U1470 (N_1470,N_896,N_926);
and U1471 (N_1471,N_784,N_459);
nor U1472 (N_1472,N_227,N_251);
nand U1473 (N_1473,N_238,N_121);
and U1474 (N_1474,N_950,N_164);
or U1475 (N_1475,N_436,N_351);
nor U1476 (N_1476,N_452,N_814);
and U1477 (N_1477,N_697,N_528);
nand U1478 (N_1478,N_699,N_746);
xnor U1479 (N_1479,N_376,N_625);
or U1480 (N_1480,N_920,N_936);
xor U1481 (N_1481,N_186,N_620);
nand U1482 (N_1482,N_198,N_213);
or U1483 (N_1483,N_765,N_154);
and U1484 (N_1484,N_343,N_250);
or U1485 (N_1485,N_792,N_370);
and U1486 (N_1486,N_22,N_553);
and U1487 (N_1487,N_795,N_196);
or U1488 (N_1488,N_856,N_439);
xnor U1489 (N_1489,N_716,N_240);
nor U1490 (N_1490,N_205,N_346);
xnor U1491 (N_1491,N_753,N_348);
or U1492 (N_1492,N_632,N_102);
nor U1493 (N_1493,N_275,N_974);
nor U1494 (N_1494,N_937,N_757);
or U1495 (N_1495,N_259,N_192);
nor U1496 (N_1496,N_476,N_127);
or U1497 (N_1497,N_230,N_388);
or U1498 (N_1498,N_642,N_704);
or U1499 (N_1499,N_887,N_806);
or U1500 (N_1500,N_1,N_297);
and U1501 (N_1501,N_539,N_907);
or U1502 (N_1502,N_630,N_531);
or U1503 (N_1503,N_112,N_329);
or U1504 (N_1504,N_427,N_467);
and U1505 (N_1505,N_547,N_560);
and U1506 (N_1506,N_606,N_259);
xor U1507 (N_1507,N_816,N_875);
and U1508 (N_1508,N_591,N_759);
or U1509 (N_1509,N_854,N_321);
and U1510 (N_1510,N_358,N_842);
nand U1511 (N_1511,N_400,N_435);
or U1512 (N_1512,N_439,N_488);
or U1513 (N_1513,N_564,N_694);
or U1514 (N_1514,N_980,N_779);
nand U1515 (N_1515,N_932,N_719);
nor U1516 (N_1516,N_331,N_827);
nand U1517 (N_1517,N_103,N_326);
xor U1518 (N_1518,N_402,N_616);
nor U1519 (N_1519,N_134,N_439);
or U1520 (N_1520,N_439,N_780);
and U1521 (N_1521,N_620,N_153);
nor U1522 (N_1522,N_895,N_878);
and U1523 (N_1523,N_740,N_694);
nor U1524 (N_1524,N_844,N_783);
and U1525 (N_1525,N_763,N_691);
nor U1526 (N_1526,N_802,N_390);
nand U1527 (N_1527,N_609,N_294);
or U1528 (N_1528,N_726,N_755);
nand U1529 (N_1529,N_564,N_746);
nand U1530 (N_1530,N_417,N_406);
nor U1531 (N_1531,N_497,N_507);
xor U1532 (N_1532,N_897,N_595);
nor U1533 (N_1533,N_802,N_373);
nor U1534 (N_1534,N_135,N_659);
or U1535 (N_1535,N_109,N_144);
and U1536 (N_1536,N_786,N_111);
and U1537 (N_1537,N_412,N_494);
xnor U1538 (N_1538,N_697,N_801);
nand U1539 (N_1539,N_615,N_31);
xor U1540 (N_1540,N_55,N_591);
nand U1541 (N_1541,N_989,N_40);
xor U1542 (N_1542,N_432,N_447);
or U1543 (N_1543,N_89,N_439);
and U1544 (N_1544,N_153,N_806);
nand U1545 (N_1545,N_457,N_332);
xnor U1546 (N_1546,N_616,N_652);
xor U1547 (N_1547,N_307,N_645);
xor U1548 (N_1548,N_94,N_768);
nand U1549 (N_1549,N_77,N_959);
nand U1550 (N_1550,N_883,N_453);
xnor U1551 (N_1551,N_360,N_203);
xor U1552 (N_1552,N_138,N_211);
and U1553 (N_1553,N_220,N_531);
or U1554 (N_1554,N_757,N_959);
nand U1555 (N_1555,N_185,N_471);
xor U1556 (N_1556,N_678,N_728);
or U1557 (N_1557,N_666,N_540);
nor U1558 (N_1558,N_945,N_968);
nor U1559 (N_1559,N_979,N_298);
or U1560 (N_1560,N_748,N_948);
or U1561 (N_1561,N_269,N_159);
and U1562 (N_1562,N_774,N_667);
nand U1563 (N_1563,N_891,N_675);
nor U1564 (N_1564,N_193,N_779);
or U1565 (N_1565,N_637,N_911);
and U1566 (N_1566,N_729,N_825);
nor U1567 (N_1567,N_351,N_101);
xor U1568 (N_1568,N_826,N_300);
nor U1569 (N_1569,N_641,N_77);
xor U1570 (N_1570,N_673,N_825);
nand U1571 (N_1571,N_688,N_45);
nor U1572 (N_1572,N_238,N_289);
and U1573 (N_1573,N_497,N_140);
or U1574 (N_1574,N_572,N_304);
nor U1575 (N_1575,N_450,N_59);
or U1576 (N_1576,N_262,N_961);
nor U1577 (N_1577,N_679,N_353);
or U1578 (N_1578,N_13,N_683);
and U1579 (N_1579,N_607,N_369);
or U1580 (N_1580,N_877,N_867);
or U1581 (N_1581,N_435,N_760);
or U1582 (N_1582,N_758,N_593);
or U1583 (N_1583,N_761,N_894);
nand U1584 (N_1584,N_979,N_587);
nor U1585 (N_1585,N_12,N_825);
xnor U1586 (N_1586,N_281,N_711);
nand U1587 (N_1587,N_75,N_318);
and U1588 (N_1588,N_381,N_258);
xnor U1589 (N_1589,N_530,N_441);
nor U1590 (N_1590,N_629,N_889);
xor U1591 (N_1591,N_998,N_320);
and U1592 (N_1592,N_961,N_164);
nand U1593 (N_1593,N_625,N_903);
or U1594 (N_1594,N_534,N_426);
and U1595 (N_1595,N_773,N_623);
nand U1596 (N_1596,N_332,N_539);
nand U1597 (N_1597,N_538,N_103);
or U1598 (N_1598,N_961,N_128);
and U1599 (N_1599,N_707,N_166);
nand U1600 (N_1600,N_987,N_109);
and U1601 (N_1601,N_259,N_80);
nand U1602 (N_1602,N_479,N_184);
nand U1603 (N_1603,N_890,N_369);
and U1604 (N_1604,N_15,N_591);
xor U1605 (N_1605,N_874,N_92);
nand U1606 (N_1606,N_352,N_13);
and U1607 (N_1607,N_40,N_864);
and U1608 (N_1608,N_912,N_336);
nand U1609 (N_1609,N_941,N_54);
or U1610 (N_1610,N_375,N_403);
xor U1611 (N_1611,N_860,N_936);
nand U1612 (N_1612,N_3,N_172);
nand U1613 (N_1613,N_301,N_392);
nand U1614 (N_1614,N_495,N_572);
nor U1615 (N_1615,N_444,N_602);
and U1616 (N_1616,N_389,N_355);
or U1617 (N_1617,N_144,N_118);
nor U1618 (N_1618,N_475,N_920);
nand U1619 (N_1619,N_650,N_95);
or U1620 (N_1620,N_909,N_559);
and U1621 (N_1621,N_57,N_66);
or U1622 (N_1622,N_122,N_674);
nand U1623 (N_1623,N_909,N_997);
or U1624 (N_1624,N_812,N_431);
or U1625 (N_1625,N_167,N_994);
and U1626 (N_1626,N_153,N_60);
and U1627 (N_1627,N_467,N_537);
and U1628 (N_1628,N_633,N_124);
nor U1629 (N_1629,N_766,N_559);
and U1630 (N_1630,N_555,N_386);
xnor U1631 (N_1631,N_370,N_356);
nand U1632 (N_1632,N_947,N_245);
nand U1633 (N_1633,N_284,N_8);
or U1634 (N_1634,N_649,N_174);
nor U1635 (N_1635,N_749,N_796);
and U1636 (N_1636,N_310,N_616);
nand U1637 (N_1637,N_940,N_280);
nand U1638 (N_1638,N_644,N_703);
xor U1639 (N_1639,N_195,N_527);
xor U1640 (N_1640,N_923,N_736);
nor U1641 (N_1641,N_377,N_948);
or U1642 (N_1642,N_842,N_463);
or U1643 (N_1643,N_461,N_399);
and U1644 (N_1644,N_644,N_660);
nand U1645 (N_1645,N_981,N_670);
nor U1646 (N_1646,N_85,N_398);
nand U1647 (N_1647,N_96,N_182);
xnor U1648 (N_1648,N_209,N_921);
nor U1649 (N_1649,N_175,N_637);
or U1650 (N_1650,N_619,N_274);
xor U1651 (N_1651,N_683,N_288);
nor U1652 (N_1652,N_187,N_728);
nand U1653 (N_1653,N_939,N_6);
nand U1654 (N_1654,N_671,N_747);
nor U1655 (N_1655,N_624,N_356);
nor U1656 (N_1656,N_133,N_116);
nand U1657 (N_1657,N_705,N_181);
nor U1658 (N_1658,N_267,N_495);
or U1659 (N_1659,N_43,N_378);
and U1660 (N_1660,N_190,N_636);
or U1661 (N_1661,N_370,N_591);
or U1662 (N_1662,N_859,N_172);
or U1663 (N_1663,N_459,N_762);
xnor U1664 (N_1664,N_618,N_422);
and U1665 (N_1665,N_502,N_751);
nor U1666 (N_1666,N_35,N_91);
and U1667 (N_1667,N_333,N_434);
or U1668 (N_1668,N_523,N_509);
or U1669 (N_1669,N_425,N_554);
or U1670 (N_1670,N_632,N_427);
or U1671 (N_1671,N_254,N_994);
and U1672 (N_1672,N_508,N_770);
or U1673 (N_1673,N_457,N_57);
xnor U1674 (N_1674,N_560,N_129);
and U1675 (N_1675,N_140,N_750);
nor U1676 (N_1676,N_334,N_808);
and U1677 (N_1677,N_850,N_765);
and U1678 (N_1678,N_184,N_581);
xnor U1679 (N_1679,N_852,N_814);
and U1680 (N_1680,N_791,N_392);
nor U1681 (N_1681,N_702,N_822);
nand U1682 (N_1682,N_321,N_627);
nand U1683 (N_1683,N_157,N_356);
or U1684 (N_1684,N_954,N_252);
xnor U1685 (N_1685,N_161,N_136);
and U1686 (N_1686,N_980,N_867);
nor U1687 (N_1687,N_246,N_311);
nand U1688 (N_1688,N_118,N_428);
nand U1689 (N_1689,N_312,N_718);
or U1690 (N_1690,N_56,N_565);
or U1691 (N_1691,N_691,N_742);
nand U1692 (N_1692,N_942,N_968);
nor U1693 (N_1693,N_464,N_147);
xnor U1694 (N_1694,N_580,N_33);
xnor U1695 (N_1695,N_656,N_212);
and U1696 (N_1696,N_956,N_949);
or U1697 (N_1697,N_888,N_559);
nor U1698 (N_1698,N_466,N_342);
nor U1699 (N_1699,N_877,N_131);
xnor U1700 (N_1700,N_97,N_121);
or U1701 (N_1701,N_644,N_247);
xor U1702 (N_1702,N_307,N_578);
or U1703 (N_1703,N_813,N_439);
or U1704 (N_1704,N_18,N_547);
or U1705 (N_1705,N_463,N_685);
xor U1706 (N_1706,N_552,N_695);
nor U1707 (N_1707,N_468,N_623);
xor U1708 (N_1708,N_819,N_800);
xor U1709 (N_1709,N_121,N_38);
or U1710 (N_1710,N_213,N_894);
nor U1711 (N_1711,N_707,N_578);
or U1712 (N_1712,N_467,N_617);
or U1713 (N_1713,N_788,N_579);
and U1714 (N_1714,N_208,N_709);
and U1715 (N_1715,N_241,N_434);
nand U1716 (N_1716,N_986,N_861);
and U1717 (N_1717,N_669,N_42);
and U1718 (N_1718,N_606,N_192);
nor U1719 (N_1719,N_422,N_731);
nand U1720 (N_1720,N_865,N_517);
nor U1721 (N_1721,N_839,N_269);
nor U1722 (N_1722,N_159,N_732);
xor U1723 (N_1723,N_392,N_628);
nand U1724 (N_1724,N_760,N_336);
nor U1725 (N_1725,N_777,N_566);
nand U1726 (N_1726,N_659,N_986);
and U1727 (N_1727,N_545,N_211);
xor U1728 (N_1728,N_318,N_430);
or U1729 (N_1729,N_756,N_697);
nand U1730 (N_1730,N_610,N_14);
or U1731 (N_1731,N_588,N_229);
nor U1732 (N_1732,N_864,N_169);
and U1733 (N_1733,N_299,N_822);
xor U1734 (N_1734,N_100,N_888);
and U1735 (N_1735,N_501,N_457);
nand U1736 (N_1736,N_133,N_100);
and U1737 (N_1737,N_948,N_671);
or U1738 (N_1738,N_388,N_207);
and U1739 (N_1739,N_360,N_401);
xor U1740 (N_1740,N_887,N_525);
and U1741 (N_1741,N_608,N_135);
nand U1742 (N_1742,N_217,N_30);
xor U1743 (N_1743,N_58,N_603);
nor U1744 (N_1744,N_776,N_949);
nor U1745 (N_1745,N_784,N_344);
xnor U1746 (N_1746,N_342,N_581);
nor U1747 (N_1747,N_181,N_15);
and U1748 (N_1748,N_94,N_448);
or U1749 (N_1749,N_205,N_468);
nand U1750 (N_1750,N_106,N_125);
nor U1751 (N_1751,N_238,N_277);
xnor U1752 (N_1752,N_220,N_476);
xnor U1753 (N_1753,N_764,N_937);
nor U1754 (N_1754,N_852,N_481);
and U1755 (N_1755,N_301,N_271);
nand U1756 (N_1756,N_329,N_259);
or U1757 (N_1757,N_759,N_28);
or U1758 (N_1758,N_500,N_50);
nor U1759 (N_1759,N_542,N_752);
or U1760 (N_1760,N_499,N_90);
or U1761 (N_1761,N_799,N_906);
nand U1762 (N_1762,N_114,N_581);
nor U1763 (N_1763,N_453,N_601);
xor U1764 (N_1764,N_300,N_444);
and U1765 (N_1765,N_194,N_163);
or U1766 (N_1766,N_917,N_939);
nand U1767 (N_1767,N_980,N_482);
nor U1768 (N_1768,N_445,N_117);
xor U1769 (N_1769,N_281,N_272);
nor U1770 (N_1770,N_227,N_337);
and U1771 (N_1771,N_946,N_240);
or U1772 (N_1772,N_570,N_473);
nor U1773 (N_1773,N_577,N_268);
nor U1774 (N_1774,N_587,N_47);
nor U1775 (N_1775,N_534,N_756);
xnor U1776 (N_1776,N_814,N_412);
or U1777 (N_1777,N_89,N_288);
nand U1778 (N_1778,N_86,N_143);
and U1779 (N_1779,N_792,N_798);
xor U1780 (N_1780,N_68,N_692);
xor U1781 (N_1781,N_64,N_800);
nor U1782 (N_1782,N_181,N_176);
nor U1783 (N_1783,N_892,N_490);
xnor U1784 (N_1784,N_512,N_904);
xnor U1785 (N_1785,N_282,N_623);
and U1786 (N_1786,N_217,N_138);
xnor U1787 (N_1787,N_825,N_328);
nor U1788 (N_1788,N_262,N_470);
nor U1789 (N_1789,N_414,N_186);
nand U1790 (N_1790,N_481,N_446);
or U1791 (N_1791,N_94,N_705);
nor U1792 (N_1792,N_355,N_85);
nor U1793 (N_1793,N_410,N_934);
and U1794 (N_1794,N_257,N_856);
nor U1795 (N_1795,N_529,N_353);
nand U1796 (N_1796,N_739,N_569);
xnor U1797 (N_1797,N_525,N_267);
nor U1798 (N_1798,N_983,N_450);
nor U1799 (N_1799,N_465,N_354);
and U1800 (N_1800,N_16,N_212);
nor U1801 (N_1801,N_869,N_887);
and U1802 (N_1802,N_143,N_205);
nor U1803 (N_1803,N_233,N_698);
nand U1804 (N_1804,N_278,N_218);
nor U1805 (N_1805,N_689,N_5);
nor U1806 (N_1806,N_706,N_996);
nand U1807 (N_1807,N_872,N_821);
and U1808 (N_1808,N_997,N_779);
nand U1809 (N_1809,N_38,N_708);
nand U1810 (N_1810,N_353,N_384);
nand U1811 (N_1811,N_493,N_883);
nand U1812 (N_1812,N_748,N_299);
nor U1813 (N_1813,N_985,N_403);
xnor U1814 (N_1814,N_900,N_705);
and U1815 (N_1815,N_331,N_721);
and U1816 (N_1816,N_741,N_775);
xor U1817 (N_1817,N_792,N_830);
xnor U1818 (N_1818,N_744,N_824);
or U1819 (N_1819,N_283,N_226);
nor U1820 (N_1820,N_234,N_832);
xnor U1821 (N_1821,N_88,N_102);
and U1822 (N_1822,N_373,N_997);
or U1823 (N_1823,N_797,N_108);
xor U1824 (N_1824,N_93,N_199);
nand U1825 (N_1825,N_622,N_279);
nor U1826 (N_1826,N_856,N_545);
or U1827 (N_1827,N_403,N_859);
and U1828 (N_1828,N_810,N_708);
nand U1829 (N_1829,N_522,N_40);
nand U1830 (N_1830,N_197,N_876);
xnor U1831 (N_1831,N_132,N_254);
xnor U1832 (N_1832,N_84,N_599);
or U1833 (N_1833,N_525,N_139);
or U1834 (N_1834,N_774,N_978);
xnor U1835 (N_1835,N_20,N_241);
nand U1836 (N_1836,N_657,N_814);
or U1837 (N_1837,N_290,N_18);
nor U1838 (N_1838,N_727,N_506);
nor U1839 (N_1839,N_760,N_570);
and U1840 (N_1840,N_4,N_105);
and U1841 (N_1841,N_193,N_248);
xor U1842 (N_1842,N_702,N_237);
and U1843 (N_1843,N_490,N_476);
nor U1844 (N_1844,N_471,N_318);
xor U1845 (N_1845,N_101,N_440);
and U1846 (N_1846,N_391,N_876);
or U1847 (N_1847,N_620,N_986);
or U1848 (N_1848,N_424,N_499);
nor U1849 (N_1849,N_752,N_314);
and U1850 (N_1850,N_368,N_650);
nand U1851 (N_1851,N_492,N_87);
and U1852 (N_1852,N_453,N_51);
or U1853 (N_1853,N_771,N_543);
nand U1854 (N_1854,N_913,N_908);
nor U1855 (N_1855,N_832,N_915);
or U1856 (N_1856,N_688,N_891);
and U1857 (N_1857,N_569,N_663);
and U1858 (N_1858,N_881,N_380);
nand U1859 (N_1859,N_164,N_101);
nor U1860 (N_1860,N_502,N_345);
nand U1861 (N_1861,N_904,N_151);
xnor U1862 (N_1862,N_615,N_277);
xnor U1863 (N_1863,N_979,N_242);
or U1864 (N_1864,N_464,N_553);
xor U1865 (N_1865,N_974,N_74);
xor U1866 (N_1866,N_286,N_650);
and U1867 (N_1867,N_391,N_726);
or U1868 (N_1868,N_61,N_326);
and U1869 (N_1869,N_85,N_118);
and U1870 (N_1870,N_494,N_530);
nor U1871 (N_1871,N_574,N_961);
and U1872 (N_1872,N_493,N_74);
or U1873 (N_1873,N_443,N_234);
and U1874 (N_1874,N_165,N_923);
and U1875 (N_1875,N_73,N_185);
nor U1876 (N_1876,N_99,N_978);
xor U1877 (N_1877,N_458,N_664);
and U1878 (N_1878,N_832,N_416);
and U1879 (N_1879,N_96,N_657);
and U1880 (N_1880,N_241,N_562);
and U1881 (N_1881,N_655,N_11);
xnor U1882 (N_1882,N_342,N_959);
or U1883 (N_1883,N_508,N_293);
nor U1884 (N_1884,N_404,N_511);
and U1885 (N_1885,N_152,N_884);
or U1886 (N_1886,N_797,N_531);
and U1887 (N_1887,N_611,N_206);
nand U1888 (N_1888,N_658,N_354);
nand U1889 (N_1889,N_100,N_338);
xnor U1890 (N_1890,N_645,N_740);
xor U1891 (N_1891,N_567,N_252);
and U1892 (N_1892,N_962,N_404);
or U1893 (N_1893,N_27,N_584);
nand U1894 (N_1894,N_609,N_966);
nor U1895 (N_1895,N_630,N_947);
nand U1896 (N_1896,N_889,N_323);
nor U1897 (N_1897,N_91,N_558);
nand U1898 (N_1898,N_419,N_910);
or U1899 (N_1899,N_451,N_339);
or U1900 (N_1900,N_797,N_696);
nand U1901 (N_1901,N_555,N_335);
and U1902 (N_1902,N_816,N_95);
and U1903 (N_1903,N_944,N_54);
and U1904 (N_1904,N_265,N_299);
nor U1905 (N_1905,N_463,N_28);
nand U1906 (N_1906,N_643,N_525);
or U1907 (N_1907,N_380,N_220);
nand U1908 (N_1908,N_214,N_276);
xor U1909 (N_1909,N_626,N_96);
nor U1910 (N_1910,N_39,N_688);
and U1911 (N_1911,N_612,N_816);
or U1912 (N_1912,N_445,N_679);
xnor U1913 (N_1913,N_525,N_422);
and U1914 (N_1914,N_749,N_577);
nand U1915 (N_1915,N_104,N_680);
or U1916 (N_1916,N_793,N_881);
nor U1917 (N_1917,N_506,N_621);
nor U1918 (N_1918,N_26,N_568);
or U1919 (N_1919,N_931,N_348);
nand U1920 (N_1920,N_192,N_680);
nor U1921 (N_1921,N_134,N_759);
nor U1922 (N_1922,N_503,N_953);
and U1923 (N_1923,N_606,N_169);
nor U1924 (N_1924,N_49,N_171);
or U1925 (N_1925,N_137,N_218);
xnor U1926 (N_1926,N_162,N_122);
nor U1927 (N_1927,N_393,N_967);
nand U1928 (N_1928,N_348,N_820);
or U1929 (N_1929,N_753,N_411);
xnor U1930 (N_1930,N_657,N_160);
and U1931 (N_1931,N_316,N_444);
or U1932 (N_1932,N_441,N_430);
or U1933 (N_1933,N_218,N_652);
and U1934 (N_1934,N_38,N_860);
or U1935 (N_1935,N_387,N_865);
nor U1936 (N_1936,N_257,N_432);
and U1937 (N_1937,N_954,N_190);
nor U1938 (N_1938,N_595,N_836);
or U1939 (N_1939,N_682,N_739);
nand U1940 (N_1940,N_345,N_349);
nor U1941 (N_1941,N_56,N_831);
xnor U1942 (N_1942,N_253,N_385);
xor U1943 (N_1943,N_986,N_603);
and U1944 (N_1944,N_209,N_349);
and U1945 (N_1945,N_545,N_43);
xor U1946 (N_1946,N_552,N_126);
xor U1947 (N_1947,N_339,N_180);
or U1948 (N_1948,N_677,N_157);
nor U1949 (N_1949,N_299,N_459);
and U1950 (N_1950,N_759,N_478);
nand U1951 (N_1951,N_525,N_393);
xor U1952 (N_1952,N_832,N_391);
and U1953 (N_1953,N_411,N_478);
and U1954 (N_1954,N_712,N_891);
nand U1955 (N_1955,N_874,N_504);
nand U1956 (N_1956,N_560,N_478);
nand U1957 (N_1957,N_51,N_557);
or U1958 (N_1958,N_214,N_978);
nor U1959 (N_1959,N_811,N_427);
and U1960 (N_1960,N_308,N_411);
or U1961 (N_1961,N_928,N_674);
nor U1962 (N_1962,N_123,N_823);
nor U1963 (N_1963,N_615,N_143);
and U1964 (N_1964,N_54,N_450);
and U1965 (N_1965,N_825,N_502);
nand U1966 (N_1966,N_492,N_955);
nor U1967 (N_1967,N_306,N_521);
nand U1968 (N_1968,N_513,N_207);
and U1969 (N_1969,N_622,N_111);
xor U1970 (N_1970,N_25,N_885);
or U1971 (N_1971,N_823,N_548);
or U1972 (N_1972,N_16,N_478);
and U1973 (N_1973,N_583,N_148);
nand U1974 (N_1974,N_964,N_347);
nand U1975 (N_1975,N_847,N_130);
and U1976 (N_1976,N_711,N_990);
and U1977 (N_1977,N_696,N_11);
nand U1978 (N_1978,N_534,N_816);
nor U1979 (N_1979,N_680,N_789);
and U1980 (N_1980,N_963,N_425);
and U1981 (N_1981,N_756,N_673);
xnor U1982 (N_1982,N_259,N_245);
nand U1983 (N_1983,N_96,N_827);
or U1984 (N_1984,N_112,N_672);
and U1985 (N_1985,N_584,N_921);
nor U1986 (N_1986,N_759,N_530);
xor U1987 (N_1987,N_523,N_395);
or U1988 (N_1988,N_682,N_538);
or U1989 (N_1989,N_444,N_269);
and U1990 (N_1990,N_772,N_938);
and U1991 (N_1991,N_711,N_366);
nand U1992 (N_1992,N_121,N_913);
and U1993 (N_1993,N_204,N_680);
xor U1994 (N_1994,N_977,N_837);
nand U1995 (N_1995,N_414,N_892);
xnor U1996 (N_1996,N_478,N_311);
xnor U1997 (N_1997,N_878,N_41);
and U1998 (N_1998,N_196,N_838);
xor U1999 (N_1999,N_333,N_790);
and U2000 (N_2000,N_1988,N_1796);
xor U2001 (N_2001,N_1685,N_1901);
nand U2002 (N_2002,N_1217,N_1229);
nand U2003 (N_2003,N_1463,N_1477);
and U2004 (N_2004,N_1992,N_1505);
or U2005 (N_2005,N_1414,N_1244);
nor U2006 (N_2006,N_1693,N_1629);
or U2007 (N_2007,N_1269,N_1516);
and U2008 (N_2008,N_1432,N_1977);
nand U2009 (N_2009,N_1096,N_1068);
nor U2010 (N_2010,N_1262,N_1117);
or U2011 (N_2011,N_1311,N_1519);
xor U2012 (N_2012,N_1819,N_1597);
and U2013 (N_2013,N_1923,N_1409);
xnor U2014 (N_2014,N_1765,N_1037);
nor U2015 (N_2015,N_1954,N_1042);
and U2016 (N_2016,N_1856,N_1888);
nor U2017 (N_2017,N_1001,N_1695);
and U2018 (N_2018,N_1958,N_1836);
nor U2019 (N_2019,N_1300,N_1258);
nand U2020 (N_2020,N_1509,N_1458);
nor U2021 (N_2021,N_1489,N_1305);
xnor U2022 (N_2022,N_1083,N_1593);
nand U2023 (N_2023,N_1683,N_1193);
xnor U2024 (N_2024,N_1080,N_1082);
nor U2025 (N_2025,N_1885,N_1199);
and U2026 (N_2026,N_1767,N_1890);
xor U2027 (N_2027,N_1708,N_1338);
and U2028 (N_2028,N_1580,N_1047);
xor U2029 (N_2029,N_1592,N_1802);
nor U2030 (N_2030,N_1315,N_1946);
xor U2031 (N_2031,N_1492,N_1542);
or U2032 (N_2032,N_1773,N_1833);
or U2033 (N_2033,N_1549,N_1438);
or U2034 (N_2034,N_1655,N_1533);
nor U2035 (N_2035,N_1378,N_1099);
nand U2036 (N_2036,N_1002,N_1886);
nand U2037 (N_2037,N_1652,N_1972);
and U2038 (N_2038,N_1361,N_1405);
nor U2039 (N_2039,N_1600,N_1084);
xor U2040 (N_2040,N_1844,N_1555);
nand U2041 (N_2041,N_1271,N_1337);
or U2042 (N_2042,N_1771,N_1702);
nand U2043 (N_2043,N_1110,N_1257);
nand U2044 (N_2044,N_1237,N_1241);
and U2045 (N_2045,N_1916,N_1172);
or U2046 (N_2046,N_1399,N_1014);
or U2047 (N_2047,N_1725,N_1766);
nor U2048 (N_2048,N_1232,N_1926);
and U2049 (N_2049,N_1433,N_1673);
and U2050 (N_2050,N_1528,N_1670);
or U2051 (N_2051,N_1609,N_1859);
nor U2052 (N_2052,N_1281,N_1675);
or U2053 (N_2053,N_1276,N_1248);
xor U2054 (N_2054,N_1090,N_1897);
and U2055 (N_2055,N_1895,N_1967);
nand U2056 (N_2056,N_1633,N_1191);
and U2057 (N_2057,N_1547,N_1335);
xnor U2058 (N_2058,N_1436,N_1575);
or U2059 (N_2059,N_1267,N_1349);
and U2060 (N_2060,N_1862,N_1346);
or U2061 (N_2061,N_1488,N_1131);
nand U2062 (N_2062,N_1651,N_1716);
or U2063 (N_2063,N_1826,N_1984);
nor U2064 (N_2064,N_1423,N_1273);
xnor U2065 (N_2065,N_1297,N_1175);
xnor U2066 (N_2066,N_1919,N_1818);
or U2067 (N_2067,N_1918,N_1931);
nor U2068 (N_2068,N_1539,N_1166);
and U2069 (N_2069,N_1266,N_1159);
nand U2070 (N_2070,N_1548,N_1161);
nor U2071 (N_2071,N_1251,N_1933);
and U2072 (N_2072,N_1843,N_1393);
and U2073 (N_2073,N_1362,N_1447);
nor U2074 (N_2074,N_1989,N_1216);
and U2075 (N_2075,N_1665,N_1720);
and U2076 (N_2076,N_1801,N_1385);
and U2077 (N_2077,N_1207,N_1390);
nor U2078 (N_2078,N_1482,N_1824);
or U2079 (N_2079,N_1736,N_1303);
or U2080 (N_2080,N_1376,N_1927);
nor U2081 (N_2081,N_1408,N_1957);
nor U2082 (N_2082,N_1640,N_1682);
nor U2083 (N_2083,N_1004,N_1581);
or U2084 (N_2084,N_1025,N_1807);
xor U2085 (N_2085,N_1781,N_1061);
or U2086 (N_2086,N_1316,N_1636);
or U2087 (N_2087,N_1871,N_1270);
nor U2088 (N_2088,N_1914,N_1878);
and U2089 (N_2089,N_1421,N_1317);
or U2090 (N_2090,N_1615,N_1688);
xor U2091 (N_2091,N_1956,N_1472);
nand U2092 (N_2092,N_1288,N_1321);
or U2093 (N_2093,N_1469,N_1788);
xnor U2094 (N_2094,N_1278,N_1461);
nor U2095 (N_2095,N_1457,N_1471);
or U2096 (N_2096,N_1664,N_1176);
nor U2097 (N_2097,N_1272,N_1095);
or U2098 (N_2098,N_1427,N_1106);
and U2099 (N_2099,N_1586,N_1787);
nor U2100 (N_2100,N_1920,N_1026);
and U2101 (N_2101,N_1975,N_1546);
or U2102 (N_2102,N_1779,N_1732);
and U2103 (N_2103,N_1997,N_1980);
nand U2104 (N_2104,N_1413,N_1504);
xnor U2105 (N_2105,N_1033,N_1121);
nand U2106 (N_2106,N_1299,N_1704);
nor U2107 (N_2107,N_1120,N_1738);
and U2108 (N_2108,N_1127,N_1345);
or U2109 (N_2109,N_1326,N_1480);
nor U2110 (N_2110,N_1085,N_1924);
nand U2111 (N_2111,N_1769,N_1048);
xor U2112 (N_2112,N_1981,N_1202);
nor U2113 (N_2113,N_1745,N_1728);
or U2114 (N_2114,N_1727,N_1333);
nor U2115 (N_2115,N_1611,N_1006);
xor U2116 (N_2116,N_1356,N_1647);
and U2117 (N_2117,N_1696,N_1793);
and U2118 (N_2118,N_1309,N_1701);
nor U2119 (N_2119,N_1604,N_1874);
or U2120 (N_2120,N_1778,N_1606);
nor U2121 (N_2121,N_1577,N_1298);
xnor U2122 (N_2122,N_1301,N_1541);
and U2123 (N_2123,N_1021,N_1177);
xor U2124 (N_2124,N_1860,N_1621);
nand U2125 (N_2125,N_1674,N_1135);
nand U2126 (N_2126,N_1970,N_1236);
and U2127 (N_2127,N_1884,N_1784);
or U2128 (N_2128,N_1576,N_1858);
or U2129 (N_2129,N_1731,N_1396);
nor U2130 (N_2130,N_1147,N_1103);
xor U2131 (N_2131,N_1097,N_1797);
or U2132 (N_2132,N_1540,N_1848);
and U2133 (N_2133,N_1864,N_1173);
nor U2134 (N_2134,N_1192,N_1060);
or U2135 (N_2135,N_1518,N_1973);
or U2136 (N_2136,N_1478,N_1368);
nand U2137 (N_2137,N_1840,N_1046);
nor U2138 (N_2138,N_1941,N_1906);
nand U2139 (N_2139,N_1086,N_1650);
nor U2140 (N_2140,N_1929,N_1454);
nor U2141 (N_2141,N_1557,N_1442);
or U2142 (N_2142,N_1998,N_1292);
nor U2143 (N_2143,N_1059,N_1877);
nor U2144 (N_2144,N_1772,N_1870);
xor U2145 (N_2145,N_1689,N_1510);
nand U2146 (N_2146,N_1990,N_1608);
or U2147 (N_2147,N_1210,N_1717);
and U2148 (N_2148,N_1464,N_1063);
nand U2149 (N_2149,N_1323,N_1680);
and U2150 (N_2150,N_1669,N_1032);
xnor U2151 (N_2151,N_1829,N_1486);
or U2152 (N_2152,N_1206,N_1122);
xor U2153 (N_2153,N_1003,N_1625);
xnor U2154 (N_2154,N_1805,N_1714);
or U2155 (N_2155,N_1286,N_1056);
nand U2156 (N_2156,N_1287,N_1863);
or U2157 (N_2157,N_1430,N_1839);
nand U2158 (N_2158,N_1841,N_1564);
or U2159 (N_2159,N_1184,N_1164);
xor U2160 (N_2160,N_1743,N_1699);
or U2161 (N_2161,N_1293,N_1630);
nand U2162 (N_2162,N_1452,N_1986);
xor U2163 (N_2163,N_1587,N_1729);
and U2164 (N_2164,N_1439,N_1538);
and U2165 (N_2165,N_1995,N_1320);
and U2166 (N_2166,N_1149,N_1676);
or U2167 (N_2167,N_1294,N_1648);
xor U2168 (N_2168,N_1188,N_1571);
and U2169 (N_2169,N_1764,N_1443);
xor U2170 (N_2170,N_1394,N_1775);
or U2171 (N_2171,N_1698,N_1656);
nand U2172 (N_2172,N_1429,N_1107);
or U2173 (N_2173,N_1198,N_1196);
and U2174 (N_2174,N_1734,N_1041);
or U2175 (N_2175,N_1247,N_1614);
nand U2176 (N_2176,N_1075,N_1749);
or U2177 (N_2177,N_1327,N_1307);
and U2178 (N_2178,N_1126,N_1343);
nand U2179 (N_2179,N_1602,N_1579);
or U2180 (N_2180,N_1130,N_1373);
or U2181 (N_2181,N_1976,N_1289);
and U2182 (N_2182,N_1619,N_1588);
or U2183 (N_2183,N_1465,N_1827);
nor U2184 (N_2184,N_1092,N_1360);
or U2185 (N_2185,N_1948,N_1102);
and U2186 (N_2186,N_1435,N_1357);
xor U2187 (N_2187,N_1978,N_1391);
nand U2188 (N_2188,N_1366,N_1653);
nand U2189 (N_2189,N_1453,N_1211);
or U2190 (N_2190,N_1560,N_1044);
and U2191 (N_2191,N_1200,N_1329);
nand U2192 (N_2192,N_1077,N_1017);
nor U2193 (N_2193,N_1881,N_1562);
or U2194 (N_2194,N_1785,N_1585);
nand U2195 (N_2195,N_1055,N_1529);
nor U2196 (N_2196,N_1649,N_1851);
and U2197 (N_2197,N_1777,N_1114);
xor U2198 (N_2198,N_1145,N_1567);
or U2199 (N_2199,N_1726,N_1383);
nand U2200 (N_2200,N_1238,N_1181);
and U2201 (N_2201,N_1506,N_1468);
and U2202 (N_2202,N_1559,N_1328);
and U2203 (N_2203,N_1950,N_1554);
nor U2204 (N_2204,N_1961,N_1312);
nand U2205 (N_2205,N_1220,N_1049);
nor U2206 (N_2206,N_1907,N_1475);
xor U2207 (N_2207,N_1310,N_1431);
xor U2208 (N_2208,N_1719,N_1138);
or U2209 (N_2209,N_1628,N_1991);
nor U2210 (N_2210,N_1476,N_1228);
nor U2211 (N_2211,N_1511,N_1353);
or U2212 (N_2212,N_1804,N_1324);
and U2213 (N_2213,N_1525,N_1341);
nand U2214 (N_2214,N_1253,N_1190);
or U2215 (N_2215,N_1005,N_1474);
nor U2216 (N_2216,N_1180,N_1865);
xnor U2217 (N_2217,N_1620,N_1798);
and U2218 (N_2218,N_1178,N_1484);
and U2219 (N_2219,N_1544,N_1815);
nand U2220 (N_2220,N_1142,N_1275);
xnor U2221 (N_2221,N_1873,N_1896);
nand U2222 (N_2222,N_1296,N_1274);
and U2223 (N_2223,N_1389,N_1583);
nor U2224 (N_2224,N_1700,N_1634);
or U2225 (N_2225,N_1768,N_1134);
and U2226 (N_2226,N_1022,N_1174);
xor U2227 (N_2227,N_1645,N_1119);
xor U2228 (N_2228,N_1817,N_1456);
nand U2229 (N_2229,N_1459,N_1867);
or U2230 (N_2230,N_1894,N_1491);
xor U2231 (N_2231,N_1355,N_1759);
xor U2232 (N_2232,N_1868,N_1069);
or U2233 (N_2233,N_1012,N_1460);
or U2234 (N_2234,N_1502,N_1939);
nand U2235 (N_2235,N_1291,N_1955);
xnor U2236 (N_2236,N_1064,N_1481);
nor U2237 (N_2237,N_1748,N_1382);
and U2238 (N_2238,N_1898,N_1799);
nor U2239 (N_2239,N_1569,N_1842);
nand U2240 (N_2240,N_1832,N_1325);
or U2241 (N_2241,N_1395,N_1747);
nor U2242 (N_2242,N_1233,N_1483);
nand U2243 (N_2243,N_1155,N_1524);
xor U2244 (N_2244,N_1133,N_1637);
and U2245 (N_2245,N_1574,N_1850);
nand U2246 (N_2246,N_1411,N_1831);
or U2247 (N_2247,N_1657,N_1902);
xnor U2248 (N_2248,N_1009,N_1887);
xnor U2249 (N_2249,N_1031,N_1835);
nand U2250 (N_2250,N_1514,N_1959);
nor U2251 (N_2251,N_1953,N_1380);
or U2252 (N_2252,N_1040,N_1783);
xor U2253 (N_2253,N_1162,N_1372);
nand U2254 (N_2254,N_1662,N_1553);
or U2255 (N_2255,N_1111,N_1790);
nand U2256 (N_2256,N_1379,N_1617);
nor U2257 (N_2257,N_1952,N_1537);
and U2258 (N_2258,N_1942,N_1422);
xor U2259 (N_2259,N_1183,N_1935);
nand U2260 (N_2260,N_1712,N_1883);
and U2261 (N_2261,N_1915,N_1322);
nand U2262 (N_2262,N_1485,N_1760);
nor U2263 (N_2263,N_1479,N_1171);
nand U2264 (N_2264,N_1691,N_1302);
xor U2265 (N_2265,N_1370,N_1150);
nand U2266 (N_2266,N_1869,N_1146);
or U2267 (N_2267,N_1644,N_1028);
and U2268 (N_2268,N_1219,N_1104);
or U2269 (N_2269,N_1962,N_1215);
xnor U2270 (N_2270,N_1521,N_1853);
nor U2271 (N_2271,N_1501,N_1234);
or U2272 (N_2272,N_1034,N_1710);
nor U2273 (N_2273,N_1761,N_1347);
or U2274 (N_2274,N_1638,N_1938);
xor U2275 (N_2275,N_1550,N_1814);
and U2276 (N_2276,N_1904,N_1803);
and U2277 (N_2277,N_1187,N_1318);
or U2278 (N_2278,N_1365,N_1227);
nand U2279 (N_2279,N_1222,N_1757);
nand U2280 (N_2280,N_1808,N_1124);
nor U2281 (N_2281,N_1330,N_1879);
xnor U2282 (N_2282,N_1816,N_1515);
nand U2283 (N_2283,N_1319,N_1721);
and U2284 (N_2284,N_1074,N_1256);
xor U2285 (N_2285,N_1601,N_1358);
nand U2286 (N_2286,N_1596,N_1201);
xnor U2287 (N_2287,N_1532,N_1160);
xnor U2288 (N_2288,N_1987,N_1921);
xor U2289 (N_2289,N_1951,N_1444);
nand U2290 (N_2290,N_1925,N_1561);
nand U2291 (N_2291,N_1910,N_1038);
nor U2292 (N_2292,N_1045,N_1071);
and U2293 (N_2293,N_1285,N_1945);
xnor U2294 (N_2294,N_1030,N_1163);
or U2295 (N_2295,N_1051,N_1354);
nand U2296 (N_2296,N_1616,N_1572);
and U2297 (N_2297,N_1066,N_1806);
nand U2298 (N_2298,N_1966,N_1654);
or U2299 (N_2299,N_1861,N_1448);
and U2300 (N_2300,N_1526,N_1535);
nand U2301 (N_2301,N_1566,N_1093);
and U2302 (N_2302,N_1407,N_1369);
nand U2303 (N_2303,N_1057,N_1733);
xor U2304 (N_2304,N_1306,N_1899);
nor U2305 (N_2305,N_1158,N_1756);
nand U2306 (N_2306,N_1866,N_1240);
nand U2307 (N_2307,N_1893,N_1404);
and U2308 (N_2308,N_1203,N_1812);
or U2309 (N_2309,N_1058,N_1010);
or U2310 (N_2310,N_1857,N_1632);
nand U2311 (N_2311,N_1744,N_1118);
and U2312 (N_2312,N_1612,N_1008);
nand U2313 (N_2313,N_1445,N_1239);
xnor U2314 (N_2314,N_1882,N_1208);
nor U2315 (N_2315,N_1344,N_1410);
and U2316 (N_2316,N_1993,N_1681);
nand U2317 (N_2317,N_1179,N_1255);
and U2318 (N_2318,N_1892,N_1496);
nor U2319 (N_2319,N_1499,N_1949);
or U2320 (N_2320,N_1838,N_1168);
and U2321 (N_2321,N_1594,N_1451);
and U2322 (N_2322,N_1283,N_1723);
and U2323 (N_2323,N_1377,N_1350);
nor U2324 (N_2324,N_1641,N_1054);
nand U2325 (N_2325,N_1195,N_1610);
nand U2326 (N_2326,N_1936,N_1658);
and U2327 (N_2327,N_1416,N_1212);
nor U2328 (N_2328,N_1011,N_1437);
xnor U2329 (N_2329,N_1268,N_1245);
nor U2330 (N_2330,N_1050,N_1367);
nand U2331 (N_2331,N_1500,N_1157);
nor U2332 (N_2332,N_1282,N_1406);
nor U2333 (N_2333,N_1613,N_1144);
xor U2334 (N_2334,N_1023,N_1622);
nor U2335 (N_2335,N_1332,N_1128);
nand U2336 (N_2336,N_1226,N_1739);
nand U2337 (N_2337,N_1223,N_1875);
and U2338 (N_2338,N_1340,N_1308);
nand U2339 (N_2339,N_1678,N_1170);
nor U2340 (N_2340,N_1348,N_1758);
or U2341 (N_2341,N_1419,N_1243);
nand U2342 (N_2342,N_1754,N_1339);
xnor U2343 (N_2343,N_1624,N_1230);
nor U2344 (N_2344,N_1584,N_1094);
and U2345 (N_2345,N_1917,N_1737);
xnor U2346 (N_2346,N_1552,N_1908);
nor U2347 (N_2347,N_1473,N_1375);
or U2348 (N_2348,N_1570,N_1224);
nand U2349 (N_2349,N_1813,N_1746);
xnor U2350 (N_2350,N_1847,N_1928);
xnor U2351 (N_2351,N_1167,N_1755);
and U2352 (N_2352,N_1697,N_1690);
nand U2353 (N_2353,N_1999,N_1663);
nor U2354 (N_2354,N_1763,N_1139);
xor U2355 (N_2355,N_1522,N_1589);
nand U2356 (N_2356,N_1715,N_1013);
xor U2357 (N_2357,N_1284,N_1374);
nor U2358 (N_2358,N_1052,N_1742);
nor U2359 (N_2359,N_1551,N_1252);
and U2360 (N_2360,N_1112,N_1132);
and U2361 (N_2361,N_1101,N_1852);
nor U2362 (N_2362,N_1627,N_1667);
and U2363 (N_2363,N_1930,N_1225);
nor U2364 (N_2364,N_1590,N_1249);
and U2365 (N_2365,N_1591,N_1115);
or U2366 (N_2366,N_1677,N_1810);
or U2367 (N_2367,N_1467,N_1724);
and U2368 (N_2368,N_1019,N_1334);
nand U2369 (N_2369,N_1455,N_1635);
xor U2370 (N_2370,N_1671,N_1072);
or U2371 (N_2371,N_1290,N_1730);
nor U2372 (N_2372,N_1098,N_1845);
or U2373 (N_2373,N_1398,N_1076);
nor U2374 (N_2374,N_1666,N_1336);
nor U2375 (N_2375,N_1036,N_1425);
nor U2376 (N_2376,N_1053,N_1364);
and U2377 (N_2377,N_1381,N_1789);
and U2378 (N_2378,N_1070,N_1351);
nor U2379 (N_2379,N_1631,N_1568);
nor U2380 (N_2380,N_1194,N_1872);
xnor U2381 (N_2381,N_1821,N_1235);
nor U2382 (N_2382,N_1039,N_1470);
xor U2383 (N_2383,N_1711,N_1129);
nand U2384 (N_2384,N_1903,N_1125);
and U2385 (N_2385,N_1441,N_1259);
nand U2386 (N_2386,N_1169,N_1913);
or U2387 (N_2387,N_1782,N_1507);
and U2388 (N_2388,N_1982,N_1646);
or U2389 (N_2389,N_1363,N_1822);
xor U2390 (N_2390,N_1709,N_1141);
nor U2391 (N_2391,N_1944,N_1545);
xnor U2392 (N_2392,N_1932,N_1820);
or U2393 (N_2393,N_1417,N_1794);
or U2394 (N_2394,N_1420,N_1397);
or U2395 (N_2395,N_1151,N_1752);
or U2396 (N_2396,N_1722,N_1679);
xor U2397 (N_2397,N_1791,N_1912);
nor U2398 (N_2398,N_1035,N_1081);
xor U2399 (N_2399,N_1969,N_1979);
nor U2400 (N_2400,N_1762,N_1062);
and U2401 (N_2401,N_1020,N_1000);
xnor U2402 (N_2402,N_1684,N_1260);
and U2403 (N_2403,N_1154,N_1740);
nor U2404 (N_2404,N_1934,N_1512);
or U2405 (N_2405,N_1985,N_1828);
xnor U2406 (N_2406,N_1313,N_1527);
xor U2407 (N_2407,N_1067,N_1314);
nor U2408 (N_2408,N_1264,N_1205);
or U2409 (N_2409,N_1943,N_1209);
nor U2410 (N_2410,N_1186,N_1520);
and U2411 (N_2411,N_1493,N_1900);
and U2412 (N_2412,N_1153,N_1971);
nor U2413 (N_2413,N_1446,N_1741);
xnor U2414 (N_2414,N_1091,N_1922);
and U2415 (N_2415,N_1400,N_1466);
nand U2416 (N_2416,N_1494,N_1123);
and U2417 (N_2417,N_1672,N_1450);
and U2418 (N_2418,N_1668,N_1974);
and U2419 (N_2419,N_1359,N_1774);
nand U2420 (N_2420,N_1497,N_1603);
nor U2421 (N_2421,N_1079,N_1029);
and U2422 (N_2422,N_1462,N_1531);
nand U2423 (N_2423,N_1434,N_1792);
nand U2424 (N_2424,N_1043,N_1089);
xor U2425 (N_2425,N_1280,N_1854);
nor U2426 (N_2426,N_1643,N_1795);
or U2427 (N_2427,N_1607,N_1498);
or U2428 (N_2428,N_1983,N_1116);
or U2429 (N_2429,N_1265,N_1136);
or U2430 (N_2430,N_1024,N_1964);
and U2431 (N_2431,N_1880,N_1642);
nor U2432 (N_2432,N_1213,N_1889);
and U2433 (N_2433,N_1189,N_1108);
xor U2434 (N_2434,N_1261,N_1113);
xor U2435 (N_2435,N_1837,N_1578);
or U2436 (N_2436,N_1384,N_1786);
nand U2437 (N_2437,N_1751,N_1148);
nand U2438 (N_2438,N_1304,N_1718);
xnor U2439 (N_2439,N_1523,N_1246);
and U2440 (N_2440,N_1937,N_1140);
nor U2441 (N_2441,N_1996,N_1440);
nor U2442 (N_2442,N_1088,N_1753);
xor U2443 (N_2443,N_1558,N_1846);
nand U2444 (N_2444,N_1027,N_1109);
and U2445 (N_2445,N_1418,N_1618);
xnor U2446 (N_2446,N_1428,N_1947);
or U2447 (N_2447,N_1735,N_1536);
xnor U2448 (N_2448,N_1279,N_1968);
and U2449 (N_2449,N_1849,N_1543);
xor U2450 (N_2450,N_1007,N_1563);
and U2451 (N_2451,N_1403,N_1940);
or U2452 (N_2452,N_1660,N_1078);
nor U2453 (N_2453,N_1073,N_1143);
and U2454 (N_2454,N_1556,N_1426);
nand U2455 (N_2455,N_1855,N_1963);
nor U2456 (N_2456,N_1692,N_1214);
nor U2457 (N_2457,N_1776,N_1595);
or U2458 (N_2458,N_1331,N_1834);
xor U2459 (N_2459,N_1825,N_1197);
or U2460 (N_2460,N_1706,N_1534);
or U2461 (N_2461,N_1295,N_1830);
and U2462 (N_2462,N_1242,N_1876);
or U2463 (N_2463,N_1909,N_1960);
xor U2464 (N_2464,N_1352,N_1016);
and U2465 (N_2465,N_1254,N_1424);
nand U2466 (N_2466,N_1687,N_1263);
nor U2467 (N_2467,N_1449,N_1487);
xor U2468 (N_2468,N_1694,N_1573);
nor U2469 (N_2469,N_1401,N_1770);
or U2470 (N_2470,N_1250,N_1015);
or U2471 (N_2471,N_1087,N_1105);
xor U2472 (N_2472,N_1623,N_1371);
or U2473 (N_2473,N_1750,N_1412);
and U2474 (N_2474,N_1402,N_1599);
nand U2475 (N_2475,N_1415,N_1182);
and U2476 (N_2476,N_1165,N_1152);
xor U2477 (N_2477,N_1705,N_1905);
nand U2478 (N_2478,N_1530,N_1800);
xor U2479 (N_2479,N_1218,N_1156);
xnor U2480 (N_2480,N_1707,N_1811);
xor U2481 (N_2481,N_1713,N_1686);
and U2482 (N_2482,N_1231,N_1598);
nor U2483 (N_2483,N_1639,N_1386);
nand U2484 (N_2484,N_1809,N_1204);
nor U2485 (N_2485,N_1392,N_1626);
xor U2486 (N_2486,N_1490,N_1994);
or U2487 (N_2487,N_1503,N_1517);
xor U2488 (N_2488,N_1342,N_1387);
xor U2489 (N_2489,N_1780,N_1018);
and U2490 (N_2490,N_1137,N_1565);
and U2491 (N_2491,N_1582,N_1388);
and U2492 (N_2492,N_1891,N_1508);
or U2493 (N_2493,N_1965,N_1823);
nor U2494 (N_2494,N_1659,N_1065);
nor U2495 (N_2495,N_1185,N_1221);
xnor U2496 (N_2496,N_1911,N_1513);
nor U2497 (N_2497,N_1605,N_1100);
or U2498 (N_2498,N_1703,N_1495);
nor U2499 (N_2499,N_1661,N_1277);
xnor U2500 (N_2500,N_1960,N_1820);
or U2501 (N_2501,N_1722,N_1934);
and U2502 (N_2502,N_1721,N_1921);
and U2503 (N_2503,N_1936,N_1135);
nor U2504 (N_2504,N_1721,N_1380);
or U2505 (N_2505,N_1929,N_1824);
nand U2506 (N_2506,N_1799,N_1410);
or U2507 (N_2507,N_1606,N_1996);
nor U2508 (N_2508,N_1784,N_1254);
or U2509 (N_2509,N_1279,N_1792);
nand U2510 (N_2510,N_1555,N_1564);
nor U2511 (N_2511,N_1529,N_1776);
nand U2512 (N_2512,N_1387,N_1925);
nand U2513 (N_2513,N_1567,N_1161);
or U2514 (N_2514,N_1830,N_1124);
xor U2515 (N_2515,N_1702,N_1410);
or U2516 (N_2516,N_1253,N_1159);
nand U2517 (N_2517,N_1591,N_1263);
nor U2518 (N_2518,N_1468,N_1374);
nor U2519 (N_2519,N_1850,N_1340);
nor U2520 (N_2520,N_1529,N_1646);
xnor U2521 (N_2521,N_1390,N_1841);
and U2522 (N_2522,N_1137,N_1338);
nor U2523 (N_2523,N_1177,N_1014);
and U2524 (N_2524,N_1073,N_1145);
and U2525 (N_2525,N_1950,N_1036);
or U2526 (N_2526,N_1437,N_1496);
and U2527 (N_2527,N_1540,N_1461);
and U2528 (N_2528,N_1674,N_1758);
or U2529 (N_2529,N_1773,N_1408);
and U2530 (N_2530,N_1339,N_1726);
nand U2531 (N_2531,N_1340,N_1364);
xor U2532 (N_2532,N_1403,N_1256);
and U2533 (N_2533,N_1233,N_1486);
nor U2534 (N_2534,N_1505,N_1117);
nor U2535 (N_2535,N_1222,N_1692);
and U2536 (N_2536,N_1633,N_1330);
or U2537 (N_2537,N_1731,N_1504);
and U2538 (N_2538,N_1623,N_1071);
and U2539 (N_2539,N_1492,N_1538);
nand U2540 (N_2540,N_1760,N_1204);
nor U2541 (N_2541,N_1911,N_1025);
xnor U2542 (N_2542,N_1478,N_1786);
nand U2543 (N_2543,N_1245,N_1940);
nand U2544 (N_2544,N_1279,N_1767);
or U2545 (N_2545,N_1794,N_1640);
nand U2546 (N_2546,N_1418,N_1916);
xnor U2547 (N_2547,N_1788,N_1133);
nand U2548 (N_2548,N_1603,N_1867);
or U2549 (N_2549,N_1372,N_1142);
xor U2550 (N_2550,N_1464,N_1741);
nand U2551 (N_2551,N_1072,N_1635);
nand U2552 (N_2552,N_1911,N_1523);
nand U2553 (N_2553,N_1170,N_1533);
nor U2554 (N_2554,N_1225,N_1942);
or U2555 (N_2555,N_1936,N_1431);
nor U2556 (N_2556,N_1823,N_1639);
or U2557 (N_2557,N_1770,N_1758);
nand U2558 (N_2558,N_1965,N_1244);
and U2559 (N_2559,N_1524,N_1592);
and U2560 (N_2560,N_1680,N_1558);
nor U2561 (N_2561,N_1905,N_1094);
or U2562 (N_2562,N_1486,N_1476);
or U2563 (N_2563,N_1187,N_1138);
or U2564 (N_2564,N_1006,N_1042);
and U2565 (N_2565,N_1152,N_1836);
and U2566 (N_2566,N_1347,N_1461);
nand U2567 (N_2567,N_1847,N_1279);
xor U2568 (N_2568,N_1463,N_1701);
nand U2569 (N_2569,N_1856,N_1605);
or U2570 (N_2570,N_1847,N_1580);
or U2571 (N_2571,N_1721,N_1075);
and U2572 (N_2572,N_1556,N_1964);
nand U2573 (N_2573,N_1013,N_1951);
nand U2574 (N_2574,N_1229,N_1093);
or U2575 (N_2575,N_1000,N_1545);
nor U2576 (N_2576,N_1253,N_1081);
or U2577 (N_2577,N_1303,N_1972);
nor U2578 (N_2578,N_1130,N_1523);
xor U2579 (N_2579,N_1489,N_1996);
nand U2580 (N_2580,N_1685,N_1152);
nor U2581 (N_2581,N_1547,N_1823);
nor U2582 (N_2582,N_1240,N_1530);
nand U2583 (N_2583,N_1832,N_1435);
or U2584 (N_2584,N_1020,N_1650);
or U2585 (N_2585,N_1136,N_1036);
nor U2586 (N_2586,N_1203,N_1810);
or U2587 (N_2587,N_1809,N_1226);
xor U2588 (N_2588,N_1104,N_1497);
or U2589 (N_2589,N_1018,N_1217);
and U2590 (N_2590,N_1353,N_1234);
or U2591 (N_2591,N_1587,N_1718);
or U2592 (N_2592,N_1319,N_1618);
and U2593 (N_2593,N_1770,N_1465);
nand U2594 (N_2594,N_1482,N_1168);
xnor U2595 (N_2595,N_1627,N_1559);
or U2596 (N_2596,N_1949,N_1129);
nor U2597 (N_2597,N_1811,N_1300);
nand U2598 (N_2598,N_1881,N_1772);
nor U2599 (N_2599,N_1300,N_1378);
and U2600 (N_2600,N_1823,N_1141);
and U2601 (N_2601,N_1706,N_1484);
and U2602 (N_2602,N_1559,N_1634);
or U2603 (N_2603,N_1468,N_1701);
and U2604 (N_2604,N_1667,N_1416);
nor U2605 (N_2605,N_1850,N_1985);
nand U2606 (N_2606,N_1102,N_1044);
and U2607 (N_2607,N_1981,N_1203);
xor U2608 (N_2608,N_1068,N_1246);
nor U2609 (N_2609,N_1329,N_1020);
and U2610 (N_2610,N_1599,N_1452);
xor U2611 (N_2611,N_1954,N_1795);
and U2612 (N_2612,N_1934,N_1614);
or U2613 (N_2613,N_1744,N_1815);
nand U2614 (N_2614,N_1784,N_1367);
xor U2615 (N_2615,N_1666,N_1101);
and U2616 (N_2616,N_1606,N_1637);
xnor U2617 (N_2617,N_1249,N_1492);
nor U2618 (N_2618,N_1731,N_1536);
xnor U2619 (N_2619,N_1575,N_1445);
nand U2620 (N_2620,N_1268,N_1587);
xor U2621 (N_2621,N_1429,N_1915);
nor U2622 (N_2622,N_1149,N_1658);
xnor U2623 (N_2623,N_1646,N_1129);
and U2624 (N_2624,N_1202,N_1824);
or U2625 (N_2625,N_1109,N_1789);
xor U2626 (N_2626,N_1732,N_1805);
and U2627 (N_2627,N_1421,N_1556);
or U2628 (N_2628,N_1037,N_1630);
xnor U2629 (N_2629,N_1689,N_1095);
and U2630 (N_2630,N_1552,N_1032);
and U2631 (N_2631,N_1870,N_1564);
or U2632 (N_2632,N_1442,N_1956);
or U2633 (N_2633,N_1090,N_1202);
and U2634 (N_2634,N_1172,N_1573);
xnor U2635 (N_2635,N_1223,N_1191);
nand U2636 (N_2636,N_1170,N_1405);
nor U2637 (N_2637,N_1615,N_1112);
nor U2638 (N_2638,N_1456,N_1512);
nand U2639 (N_2639,N_1001,N_1412);
nor U2640 (N_2640,N_1084,N_1783);
or U2641 (N_2641,N_1966,N_1710);
nor U2642 (N_2642,N_1958,N_1718);
or U2643 (N_2643,N_1197,N_1199);
nor U2644 (N_2644,N_1118,N_1907);
xor U2645 (N_2645,N_1066,N_1893);
xnor U2646 (N_2646,N_1180,N_1744);
and U2647 (N_2647,N_1362,N_1277);
or U2648 (N_2648,N_1044,N_1003);
and U2649 (N_2649,N_1801,N_1147);
nand U2650 (N_2650,N_1911,N_1739);
nand U2651 (N_2651,N_1479,N_1950);
nand U2652 (N_2652,N_1203,N_1379);
nand U2653 (N_2653,N_1067,N_1493);
xnor U2654 (N_2654,N_1577,N_1709);
nor U2655 (N_2655,N_1037,N_1355);
and U2656 (N_2656,N_1384,N_1341);
nor U2657 (N_2657,N_1404,N_1915);
nor U2658 (N_2658,N_1824,N_1463);
or U2659 (N_2659,N_1541,N_1041);
or U2660 (N_2660,N_1074,N_1117);
nand U2661 (N_2661,N_1633,N_1193);
nand U2662 (N_2662,N_1236,N_1683);
xor U2663 (N_2663,N_1041,N_1810);
nand U2664 (N_2664,N_1909,N_1484);
and U2665 (N_2665,N_1489,N_1002);
and U2666 (N_2666,N_1313,N_1685);
or U2667 (N_2667,N_1229,N_1798);
xnor U2668 (N_2668,N_1583,N_1154);
nor U2669 (N_2669,N_1707,N_1222);
xnor U2670 (N_2670,N_1954,N_1146);
xor U2671 (N_2671,N_1811,N_1113);
or U2672 (N_2672,N_1441,N_1794);
nor U2673 (N_2673,N_1151,N_1869);
nor U2674 (N_2674,N_1966,N_1944);
nor U2675 (N_2675,N_1894,N_1410);
nor U2676 (N_2676,N_1625,N_1033);
or U2677 (N_2677,N_1092,N_1337);
nand U2678 (N_2678,N_1165,N_1392);
xor U2679 (N_2679,N_1015,N_1092);
nor U2680 (N_2680,N_1937,N_1527);
and U2681 (N_2681,N_1990,N_1698);
or U2682 (N_2682,N_1425,N_1820);
nand U2683 (N_2683,N_1773,N_1268);
or U2684 (N_2684,N_1727,N_1814);
and U2685 (N_2685,N_1396,N_1697);
or U2686 (N_2686,N_1582,N_1053);
nand U2687 (N_2687,N_1778,N_1112);
nand U2688 (N_2688,N_1289,N_1980);
nor U2689 (N_2689,N_1593,N_1391);
nand U2690 (N_2690,N_1820,N_1189);
xor U2691 (N_2691,N_1285,N_1975);
nand U2692 (N_2692,N_1114,N_1687);
nor U2693 (N_2693,N_1069,N_1126);
and U2694 (N_2694,N_1578,N_1785);
nand U2695 (N_2695,N_1359,N_1200);
xor U2696 (N_2696,N_1503,N_1237);
nor U2697 (N_2697,N_1110,N_1856);
nand U2698 (N_2698,N_1005,N_1639);
nand U2699 (N_2699,N_1459,N_1112);
or U2700 (N_2700,N_1547,N_1399);
nor U2701 (N_2701,N_1556,N_1889);
nor U2702 (N_2702,N_1573,N_1123);
nand U2703 (N_2703,N_1769,N_1989);
or U2704 (N_2704,N_1379,N_1913);
or U2705 (N_2705,N_1567,N_1587);
or U2706 (N_2706,N_1862,N_1032);
and U2707 (N_2707,N_1410,N_1406);
or U2708 (N_2708,N_1123,N_1600);
nand U2709 (N_2709,N_1798,N_1952);
or U2710 (N_2710,N_1930,N_1224);
or U2711 (N_2711,N_1747,N_1881);
or U2712 (N_2712,N_1443,N_1324);
nor U2713 (N_2713,N_1192,N_1201);
xor U2714 (N_2714,N_1906,N_1374);
or U2715 (N_2715,N_1991,N_1181);
or U2716 (N_2716,N_1485,N_1076);
or U2717 (N_2717,N_1102,N_1084);
or U2718 (N_2718,N_1651,N_1245);
or U2719 (N_2719,N_1266,N_1484);
xnor U2720 (N_2720,N_1958,N_1464);
xor U2721 (N_2721,N_1726,N_1028);
xnor U2722 (N_2722,N_1923,N_1854);
or U2723 (N_2723,N_1874,N_1241);
nor U2724 (N_2724,N_1293,N_1542);
and U2725 (N_2725,N_1235,N_1153);
nand U2726 (N_2726,N_1786,N_1801);
or U2727 (N_2727,N_1448,N_1648);
or U2728 (N_2728,N_1611,N_1249);
nand U2729 (N_2729,N_1891,N_1667);
nand U2730 (N_2730,N_1502,N_1356);
xor U2731 (N_2731,N_1845,N_1617);
nand U2732 (N_2732,N_1510,N_1684);
nand U2733 (N_2733,N_1269,N_1620);
and U2734 (N_2734,N_1232,N_1233);
xor U2735 (N_2735,N_1041,N_1288);
nor U2736 (N_2736,N_1027,N_1135);
or U2737 (N_2737,N_1278,N_1636);
nand U2738 (N_2738,N_1055,N_1236);
nand U2739 (N_2739,N_1043,N_1452);
xnor U2740 (N_2740,N_1874,N_1550);
xor U2741 (N_2741,N_1875,N_1032);
nand U2742 (N_2742,N_1573,N_1897);
or U2743 (N_2743,N_1984,N_1114);
or U2744 (N_2744,N_1823,N_1179);
and U2745 (N_2745,N_1310,N_1490);
xnor U2746 (N_2746,N_1845,N_1530);
nand U2747 (N_2747,N_1463,N_1765);
xor U2748 (N_2748,N_1850,N_1642);
and U2749 (N_2749,N_1724,N_1447);
xnor U2750 (N_2750,N_1931,N_1294);
or U2751 (N_2751,N_1756,N_1698);
and U2752 (N_2752,N_1516,N_1520);
xor U2753 (N_2753,N_1842,N_1771);
xnor U2754 (N_2754,N_1302,N_1288);
nand U2755 (N_2755,N_1941,N_1177);
and U2756 (N_2756,N_1490,N_1450);
and U2757 (N_2757,N_1542,N_1283);
nor U2758 (N_2758,N_1663,N_1834);
nand U2759 (N_2759,N_1587,N_1823);
nor U2760 (N_2760,N_1885,N_1413);
xor U2761 (N_2761,N_1246,N_1508);
or U2762 (N_2762,N_1134,N_1648);
and U2763 (N_2763,N_1196,N_1226);
xor U2764 (N_2764,N_1981,N_1345);
nor U2765 (N_2765,N_1038,N_1493);
or U2766 (N_2766,N_1573,N_1900);
nor U2767 (N_2767,N_1527,N_1452);
or U2768 (N_2768,N_1216,N_1251);
and U2769 (N_2769,N_1108,N_1217);
nor U2770 (N_2770,N_1764,N_1760);
xor U2771 (N_2771,N_1016,N_1669);
and U2772 (N_2772,N_1533,N_1483);
or U2773 (N_2773,N_1525,N_1779);
or U2774 (N_2774,N_1919,N_1763);
nor U2775 (N_2775,N_1609,N_1903);
or U2776 (N_2776,N_1623,N_1830);
and U2777 (N_2777,N_1456,N_1461);
nand U2778 (N_2778,N_1943,N_1437);
xor U2779 (N_2779,N_1686,N_1770);
or U2780 (N_2780,N_1325,N_1644);
xnor U2781 (N_2781,N_1303,N_1888);
nand U2782 (N_2782,N_1757,N_1974);
xor U2783 (N_2783,N_1910,N_1617);
and U2784 (N_2784,N_1718,N_1960);
nor U2785 (N_2785,N_1605,N_1962);
nor U2786 (N_2786,N_1755,N_1946);
xor U2787 (N_2787,N_1614,N_1224);
nand U2788 (N_2788,N_1346,N_1699);
or U2789 (N_2789,N_1363,N_1662);
xnor U2790 (N_2790,N_1867,N_1820);
nor U2791 (N_2791,N_1538,N_1502);
nor U2792 (N_2792,N_1777,N_1081);
or U2793 (N_2793,N_1291,N_1515);
and U2794 (N_2794,N_1704,N_1125);
xor U2795 (N_2795,N_1645,N_1722);
or U2796 (N_2796,N_1099,N_1509);
nand U2797 (N_2797,N_1282,N_1123);
xnor U2798 (N_2798,N_1300,N_1931);
nor U2799 (N_2799,N_1087,N_1065);
nand U2800 (N_2800,N_1344,N_1075);
or U2801 (N_2801,N_1807,N_1696);
or U2802 (N_2802,N_1283,N_1238);
xor U2803 (N_2803,N_1157,N_1063);
and U2804 (N_2804,N_1358,N_1201);
and U2805 (N_2805,N_1911,N_1268);
xor U2806 (N_2806,N_1463,N_1200);
and U2807 (N_2807,N_1098,N_1489);
and U2808 (N_2808,N_1579,N_1425);
xnor U2809 (N_2809,N_1429,N_1918);
or U2810 (N_2810,N_1615,N_1489);
nor U2811 (N_2811,N_1074,N_1600);
nand U2812 (N_2812,N_1227,N_1200);
xor U2813 (N_2813,N_1296,N_1281);
nand U2814 (N_2814,N_1897,N_1595);
xor U2815 (N_2815,N_1525,N_1216);
or U2816 (N_2816,N_1703,N_1040);
and U2817 (N_2817,N_1536,N_1192);
nand U2818 (N_2818,N_1274,N_1198);
nor U2819 (N_2819,N_1397,N_1445);
nand U2820 (N_2820,N_1720,N_1303);
nor U2821 (N_2821,N_1533,N_1766);
nand U2822 (N_2822,N_1951,N_1593);
and U2823 (N_2823,N_1423,N_1100);
nor U2824 (N_2824,N_1033,N_1574);
xor U2825 (N_2825,N_1602,N_1012);
or U2826 (N_2826,N_1509,N_1239);
and U2827 (N_2827,N_1539,N_1638);
or U2828 (N_2828,N_1711,N_1143);
and U2829 (N_2829,N_1052,N_1576);
nor U2830 (N_2830,N_1171,N_1515);
nor U2831 (N_2831,N_1808,N_1971);
and U2832 (N_2832,N_1638,N_1385);
nand U2833 (N_2833,N_1613,N_1014);
nand U2834 (N_2834,N_1014,N_1842);
nand U2835 (N_2835,N_1583,N_1771);
xnor U2836 (N_2836,N_1083,N_1828);
and U2837 (N_2837,N_1807,N_1108);
xor U2838 (N_2838,N_1671,N_1638);
nand U2839 (N_2839,N_1456,N_1197);
or U2840 (N_2840,N_1076,N_1124);
nor U2841 (N_2841,N_1210,N_1437);
xnor U2842 (N_2842,N_1367,N_1597);
or U2843 (N_2843,N_1354,N_1175);
or U2844 (N_2844,N_1193,N_1125);
or U2845 (N_2845,N_1993,N_1327);
and U2846 (N_2846,N_1606,N_1010);
nand U2847 (N_2847,N_1844,N_1841);
or U2848 (N_2848,N_1447,N_1709);
xnor U2849 (N_2849,N_1882,N_1512);
xor U2850 (N_2850,N_1087,N_1554);
xnor U2851 (N_2851,N_1234,N_1605);
nand U2852 (N_2852,N_1442,N_1169);
or U2853 (N_2853,N_1489,N_1928);
xnor U2854 (N_2854,N_1604,N_1600);
xnor U2855 (N_2855,N_1780,N_1592);
and U2856 (N_2856,N_1298,N_1618);
nand U2857 (N_2857,N_1764,N_1985);
nor U2858 (N_2858,N_1135,N_1000);
nand U2859 (N_2859,N_1571,N_1902);
nand U2860 (N_2860,N_1105,N_1913);
xnor U2861 (N_2861,N_1085,N_1193);
nor U2862 (N_2862,N_1107,N_1242);
nand U2863 (N_2863,N_1706,N_1667);
or U2864 (N_2864,N_1518,N_1931);
nand U2865 (N_2865,N_1444,N_1577);
nand U2866 (N_2866,N_1519,N_1013);
nor U2867 (N_2867,N_1883,N_1295);
nor U2868 (N_2868,N_1980,N_1100);
and U2869 (N_2869,N_1748,N_1148);
or U2870 (N_2870,N_1019,N_1225);
or U2871 (N_2871,N_1907,N_1049);
nand U2872 (N_2872,N_1972,N_1238);
nor U2873 (N_2873,N_1313,N_1142);
or U2874 (N_2874,N_1955,N_1583);
or U2875 (N_2875,N_1889,N_1658);
xor U2876 (N_2876,N_1653,N_1015);
and U2877 (N_2877,N_1283,N_1474);
xnor U2878 (N_2878,N_1449,N_1190);
nor U2879 (N_2879,N_1518,N_1361);
nor U2880 (N_2880,N_1118,N_1496);
nand U2881 (N_2881,N_1477,N_1900);
nor U2882 (N_2882,N_1820,N_1180);
nand U2883 (N_2883,N_1634,N_1151);
and U2884 (N_2884,N_1186,N_1837);
nor U2885 (N_2885,N_1882,N_1127);
and U2886 (N_2886,N_1956,N_1185);
nor U2887 (N_2887,N_1476,N_1652);
nand U2888 (N_2888,N_1779,N_1699);
xor U2889 (N_2889,N_1838,N_1304);
or U2890 (N_2890,N_1258,N_1150);
and U2891 (N_2891,N_1091,N_1396);
nand U2892 (N_2892,N_1948,N_1840);
or U2893 (N_2893,N_1237,N_1311);
nand U2894 (N_2894,N_1258,N_1891);
or U2895 (N_2895,N_1367,N_1652);
and U2896 (N_2896,N_1246,N_1755);
nand U2897 (N_2897,N_1396,N_1711);
nand U2898 (N_2898,N_1428,N_1446);
nor U2899 (N_2899,N_1921,N_1159);
xor U2900 (N_2900,N_1186,N_1305);
nand U2901 (N_2901,N_1859,N_1733);
nor U2902 (N_2902,N_1519,N_1313);
nor U2903 (N_2903,N_1374,N_1234);
or U2904 (N_2904,N_1279,N_1103);
and U2905 (N_2905,N_1674,N_1114);
and U2906 (N_2906,N_1534,N_1075);
and U2907 (N_2907,N_1816,N_1055);
nor U2908 (N_2908,N_1219,N_1489);
and U2909 (N_2909,N_1326,N_1570);
and U2910 (N_2910,N_1237,N_1813);
and U2911 (N_2911,N_1274,N_1084);
xor U2912 (N_2912,N_1754,N_1443);
or U2913 (N_2913,N_1568,N_1363);
or U2914 (N_2914,N_1218,N_1630);
and U2915 (N_2915,N_1068,N_1542);
xor U2916 (N_2916,N_1498,N_1315);
nor U2917 (N_2917,N_1649,N_1186);
or U2918 (N_2918,N_1843,N_1639);
nand U2919 (N_2919,N_1538,N_1721);
xor U2920 (N_2920,N_1049,N_1776);
nor U2921 (N_2921,N_1274,N_1897);
nand U2922 (N_2922,N_1684,N_1851);
and U2923 (N_2923,N_1386,N_1231);
or U2924 (N_2924,N_1572,N_1150);
nor U2925 (N_2925,N_1042,N_1416);
nand U2926 (N_2926,N_1749,N_1274);
and U2927 (N_2927,N_1775,N_1196);
or U2928 (N_2928,N_1747,N_1306);
and U2929 (N_2929,N_1921,N_1929);
nor U2930 (N_2930,N_1124,N_1601);
nor U2931 (N_2931,N_1206,N_1104);
and U2932 (N_2932,N_1365,N_1552);
xnor U2933 (N_2933,N_1968,N_1112);
and U2934 (N_2934,N_1643,N_1561);
and U2935 (N_2935,N_1821,N_1329);
nand U2936 (N_2936,N_1579,N_1408);
and U2937 (N_2937,N_1396,N_1282);
nor U2938 (N_2938,N_1440,N_1525);
nor U2939 (N_2939,N_1046,N_1614);
nor U2940 (N_2940,N_1120,N_1076);
nand U2941 (N_2941,N_1591,N_1649);
xor U2942 (N_2942,N_1186,N_1078);
nand U2943 (N_2943,N_1793,N_1415);
and U2944 (N_2944,N_1496,N_1311);
and U2945 (N_2945,N_1708,N_1764);
nor U2946 (N_2946,N_1215,N_1581);
xnor U2947 (N_2947,N_1211,N_1031);
or U2948 (N_2948,N_1446,N_1852);
and U2949 (N_2949,N_1999,N_1992);
xor U2950 (N_2950,N_1971,N_1677);
and U2951 (N_2951,N_1150,N_1610);
and U2952 (N_2952,N_1095,N_1895);
xnor U2953 (N_2953,N_1922,N_1502);
xor U2954 (N_2954,N_1757,N_1079);
or U2955 (N_2955,N_1166,N_1987);
or U2956 (N_2956,N_1278,N_1761);
and U2957 (N_2957,N_1141,N_1742);
nand U2958 (N_2958,N_1659,N_1935);
nand U2959 (N_2959,N_1591,N_1853);
or U2960 (N_2960,N_1743,N_1385);
and U2961 (N_2961,N_1793,N_1722);
xnor U2962 (N_2962,N_1730,N_1069);
xnor U2963 (N_2963,N_1202,N_1540);
nand U2964 (N_2964,N_1580,N_1027);
xor U2965 (N_2965,N_1841,N_1432);
nand U2966 (N_2966,N_1017,N_1862);
and U2967 (N_2967,N_1892,N_1311);
or U2968 (N_2968,N_1482,N_1828);
nor U2969 (N_2969,N_1881,N_1146);
and U2970 (N_2970,N_1149,N_1566);
xnor U2971 (N_2971,N_1089,N_1656);
nor U2972 (N_2972,N_1225,N_1857);
nor U2973 (N_2973,N_1955,N_1867);
nand U2974 (N_2974,N_1096,N_1315);
xor U2975 (N_2975,N_1527,N_1041);
nand U2976 (N_2976,N_1726,N_1997);
nor U2977 (N_2977,N_1281,N_1664);
or U2978 (N_2978,N_1782,N_1547);
and U2979 (N_2979,N_1669,N_1454);
or U2980 (N_2980,N_1189,N_1371);
or U2981 (N_2981,N_1988,N_1752);
or U2982 (N_2982,N_1390,N_1325);
and U2983 (N_2983,N_1160,N_1962);
xor U2984 (N_2984,N_1135,N_1096);
xnor U2985 (N_2985,N_1906,N_1821);
and U2986 (N_2986,N_1237,N_1111);
or U2987 (N_2987,N_1448,N_1968);
xnor U2988 (N_2988,N_1931,N_1330);
or U2989 (N_2989,N_1192,N_1922);
or U2990 (N_2990,N_1512,N_1982);
and U2991 (N_2991,N_1084,N_1050);
and U2992 (N_2992,N_1165,N_1847);
xnor U2993 (N_2993,N_1551,N_1863);
nand U2994 (N_2994,N_1667,N_1099);
nor U2995 (N_2995,N_1305,N_1991);
or U2996 (N_2996,N_1902,N_1592);
and U2997 (N_2997,N_1570,N_1633);
or U2998 (N_2998,N_1211,N_1897);
nand U2999 (N_2999,N_1980,N_1123);
nand U3000 (N_3000,N_2457,N_2834);
and U3001 (N_3001,N_2073,N_2609);
nor U3002 (N_3002,N_2520,N_2975);
nand U3003 (N_3003,N_2058,N_2121);
or U3004 (N_3004,N_2014,N_2514);
nand U3005 (N_3005,N_2883,N_2044);
nand U3006 (N_3006,N_2783,N_2533);
and U3007 (N_3007,N_2633,N_2133);
xor U3008 (N_3008,N_2964,N_2510);
and U3009 (N_3009,N_2188,N_2995);
and U3010 (N_3010,N_2280,N_2199);
nor U3011 (N_3011,N_2852,N_2315);
nand U3012 (N_3012,N_2996,N_2301);
and U3013 (N_3013,N_2036,N_2412);
or U3014 (N_3014,N_2773,N_2334);
nand U3015 (N_3015,N_2085,N_2824);
or U3016 (N_3016,N_2562,N_2988);
xor U3017 (N_3017,N_2637,N_2639);
nand U3018 (N_3018,N_2160,N_2837);
and U3019 (N_3019,N_2276,N_2971);
and U3020 (N_3020,N_2980,N_2254);
xor U3021 (N_3021,N_2331,N_2484);
or U3022 (N_3022,N_2542,N_2210);
xnor U3023 (N_3023,N_2653,N_2908);
xor U3024 (N_3024,N_2183,N_2829);
nor U3025 (N_3025,N_2107,N_2569);
xnor U3026 (N_3026,N_2587,N_2367);
nand U3027 (N_3027,N_2129,N_2373);
nor U3028 (N_3028,N_2157,N_2174);
or U3029 (N_3029,N_2558,N_2238);
xor U3030 (N_3030,N_2064,N_2035);
xor U3031 (N_3031,N_2365,N_2407);
and U3032 (N_3032,N_2590,N_2416);
nand U3033 (N_3033,N_2458,N_2962);
xnor U3034 (N_3034,N_2705,N_2127);
nor U3035 (N_3035,N_2319,N_2158);
nor U3036 (N_3036,N_2729,N_2218);
xor U3037 (N_3037,N_2414,N_2302);
and U3038 (N_3038,N_2349,N_2028);
xnor U3039 (N_3039,N_2152,N_2755);
nand U3040 (N_3040,N_2436,N_2310);
or U3041 (N_3041,N_2312,N_2222);
and U3042 (N_3042,N_2815,N_2667);
and U3043 (N_3043,N_2016,N_2998);
or U3044 (N_3044,N_2911,N_2846);
or U3045 (N_3045,N_2034,N_2622);
or U3046 (N_3046,N_2504,N_2206);
nor U3047 (N_3047,N_2659,N_2411);
and U3048 (N_3048,N_2330,N_2362);
xor U3049 (N_3049,N_2584,N_2765);
and U3050 (N_3050,N_2308,N_2781);
nor U3051 (N_3051,N_2958,N_2800);
xor U3052 (N_3052,N_2006,N_2855);
xor U3053 (N_3053,N_2722,N_2517);
xor U3054 (N_3054,N_2076,N_2051);
xnor U3055 (N_3055,N_2931,N_2526);
and U3056 (N_3056,N_2615,N_2828);
xor U3057 (N_3057,N_2770,N_2586);
and U3058 (N_3058,N_2271,N_2432);
and U3059 (N_3059,N_2888,N_2492);
xnor U3060 (N_3060,N_2066,N_2681);
xnor U3061 (N_3061,N_2554,N_2863);
nand U3062 (N_3062,N_2347,N_2135);
xor U3063 (N_3063,N_2187,N_2617);
or U3064 (N_3064,N_2671,N_2418);
and U3065 (N_3065,N_2697,N_2899);
or U3066 (N_3066,N_2951,N_2124);
nor U3067 (N_3067,N_2389,N_2664);
and U3068 (N_3068,N_2876,N_2730);
or U3069 (N_3069,N_2771,N_2581);
nor U3070 (N_3070,N_2428,N_2388);
and U3071 (N_3071,N_2039,N_2390);
and U3072 (N_3072,N_2241,N_2266);
nor U3073 (N_3073,N_2636,N_2348);
nor U3074 (N_3074,N_2948,N_2889);
nor U3075 (N_3075,N_2648,N_2720);
nand U3076 (N_3076,N_2508,N_2143);
and U3077 (N_3077,N_2378,N_2645);
xnor U3078 (N_3078,N_2038,N_2112);
nor U3079 (N_3079,N_2552,N_2716);
xor U3080 (N_3080,N_2052,N_2442);
xor U3081 (N_3081,N_2629,N_2983);
and U3082 (N_3082,N_2485,N_2712);
or U3083 (N_3083,N_2691,N_2043);
nor U3084 (N_3084,N_2233,N_2866);
nand U3085 (N_3085,N_2322,N_2283);
or U3086 (N_3086,N_2131,N_2742);
and U3087 (N_3087,N_2002,N_2912);
or U3088 (N_3088,N_2634,N_2200);
xor U3089 (N_3089,N_2725,N_2372);
or U3090 (N_3090,N_2156,N_2405);
xnor U3091 (N_3091,N_2326,N_2884);
and U3092 (N_3092,N_2605,N_2369);
xnor U3093 (N_3093,N_2787,N_2009);
nor U3094 (N_3094,N_2079,N_2292);
or U3095 (N_3095,N_2718,N_2259);
xnor U3096 (N_3096,N_2661,N_2102);
nor U3097 (N_3097,N_2491,N_2050);
xor U3098 (N_3098,N_2660,N_2231);
or U3099 (N_3099,N_2843,N_2343);
nand U3100 (N_3100,N_2930,N_2286);
nand U3101 (N_3101,N_2287,N_2630);
xor U3102 (N_3102,N_2454,N_2546);
nor U3103 (N_3103,N_2974,N_2366);
nand U3104 (N_3104,N_2841,N_2456);
xnor U3105 (N_3105,N_2679,N_2248);
xor U3106 (N_3106,N_2392,N_2472);
nand U3107 (N_3107,N_2677,N_2602);
or U3108 (N_3108,N_2874,N_2665);
nor U3109 (N_3109,N_2449,N_2926);
xor U3110 (N_3110,N_2225,N_2642);
nor U3111 (N_3111,N_2890,N_2196);
and U3112 (N_3112,N_2060,N_2500);
or U3113 (N_3113,N_2488,N_2556);
nor U3114 (N_3114,N_2025,N_2583);
or U3115 (N_3115,N_2342,N_2669);
nor U3116 (N_3116,N_2170,N_2136);
nor U3117 (N_3117,N_2325,N_2024);
or U3118 (N_3118,N_2450,N_2055);
or U3119 (N_3119,N_2859,N_2900);
nand U3120 (N_3120,N_2544,N_2003);
xor U3121 (N_3121,N_2059,N_2296);
nand U3122 (N_3122,N_2848,N_2563);
nor U3123 (N_3123,N_2710,N_2111);
and U3124 (N_3124,N_2668,N_2746);
xnor U3125 (N_3125,N_2421,N_2182);
nand U3126 (N_3126,N_2501,N_2784);
and U3127 (N_3127,N_2981,N_2067);
xnor U3128 (N_3128,N_2999,N_2550);
and U3129 (N_3129,N_2042,N_2105);
and U3130 (N_3130,N_2332,N_2140);
or U3131 (N_3131,N_2018,N_2460);
nor U3132 (N_3132,N_2875,N_2738);
xnor U3133 (N_3133,N_2640,N_2803);
and U3134 (N_3134,N_2870,N_2397);
xnor U3135 (N_3135,N_2600,N_2793);
or U3136 (N_3136,N_2905,N_2741);
nor U3137 (N_3137,N_2545,N_2597);
xor U3138 (N_3138,N_2949,N_2088);
and U3139 (N_3139,N_2524,N_2763);
or U3140 (N_3140,N_2108,N_2359);
and U3141 (N_3141,N_2915,N_2047);
or U3142 (N_3142,N_2574,N_2618);
xor U3143 (N_3143,N_2576,N_2408);
nand U3144 (N_3144,N_2809,N_2001);
nand U3145 (N_3145,N_2175,N_2236);
and U3146 (N_3146,N_2046,N_2540);
nor U3147 (N_3147,N_2082,N_2317);
and U3148 (N_3148,N_2095,N_2732);
nand U3149 (N_3149,N_2165,N_2277);
nor U3150 (N_3150,N_2598,N_2445);
nor U3151 (N_3151,N_2529,N_2619);
and U3152 (N_3152,N_2098,N_2811);
nor U3153 (N_3153,N_2898,N_2186);
xor U3154 (N_3154,N_2153,N_2228);
xnor U3155 (N_3155,N_2093,N_2263);
nand U3156 (N_3156,N_2758,N_2495);
nor U3157 (N_3157,N_2353,N_2178);
xnor U3158 (N_3158,N_2623,N_2877);
nand U3159 (N_3159,N_2713,N_2663);
nand U3160 (N_3160,N_2902,N_2641);
and U3161 (N_3161,N_2991,N_2764);
and U3162 (N_3162,N_2860,N_2928);
nand U3163 (N_3163,N_2417,N_2288);
and U3164 (N_3164,N_2490,N_2807);
nand U3165 (N_3165,N_2512,N_2269);
nand U3166 (N_3166,N_2409,N_2247);
nand U3167 (N_3167,N_2693,N_2478);
or U3168 (N_3168,N_2161,N_2080);
nand U3169 (N_3169,N_2092,N_2031);
nor U3170 (N_3170,N_2462,N_2522);
xnor U3171 (N_3171,N_2227,N_2149);
nand U3172 (N_3172,N_2239,N_2154);
xnor U3173 (N_3173,N_2480,N_2439);
nor U3174 (N_3174,N_2992,N_2291);
or U3175 (N_3175,N_2221,N_2446);
or U3176 (N_3176,N_2358,N_2997);
or U3177 (N_3177,N_2904,N_2850);
nor U3178 (N_3178,N_2530,N_2062);
nand U3179 (N_3179,N_2245,N_2191);
or U3180 (N_3180,N_2290,N_2965);
xor U3181 (N_3181,N_2614,N_2424);
and U3182 (N_3182,N_2589,N_2198);
or U3183 (N_3183,N_2110,N_2163);
nor U3184 (N_3184,N_2074,N_2371);
nor U3185 (N_3185,N_2425,N_2467);
or U3186 (N_3186,N_2386,N_2818);
or U3187 (N_3187,N_2728,N_2736);
or U3188 (N_3188,N_2977,N_2872);
xnor U3189 (N_3189,N_2830,N_2970);
nor U3190 (N_3190,N_2250,N_2268);
nor U3191 (N_3191,N_2822,N_2429);
and U3192 (N_3192,N_2960,N_2497);
nor U3193 (N_3193,N_2433,N_2635);
nor U3194 (N_3194,N_2171,N_2114);
xor U3195 (N_3195,N_2827,N_2721);
and U3196 (N_3196,N_2945,N_2953);
or U3197 (N_3197,N_2021,N_2923);
and U3198 (N_3198,N_2887,N_2447);
and U3199 (N_3199,N_2734,N_2063);
nand U3200 (N_3200,N_2894,N_2474);
xor U3201 (N_3201,N_2952,N_2982);
and U3202 (N_3202,N_2913,N_2935);
and U3203 (N_3203,N_2032,N_2806);
or U3204 (N_3204,N_2045,N_2090);
or U3205 (N_3205,N_2385,N_2297);
nand U3206 (N_3206,N_2747,N_2706);
or U3207 (N_3207,N_2604,N_2733);
nand U3208 (N_3208,N_2307,N_2832);
nand U3209 (N_3209,N_2232,N_2682);
xor U3210 (N_3210,N_2896,N_2189);
xor U3211 (N_3211,N_2620,N_2444);
nand U3212 (N_3212,N_2985,N_2507);
nor U3213 (N_3213,N_2836,N_2230);
nor U3214 (N_3214,N_2027,N_2201);
or U3215 (N_3215,N_2756,N_2934);
nor U3216 (N_3216,N_2061,N_2166);
or U3217 (N_3217,N_2625,N_2261);
or U3218 (N_3218,N_2769,N_2895);
or U3219 (N_3219,N_2125,N_2422);
nand U3220 (N_3220,N_2229,N_2656);
and U3221 (N_3221,N_2745,N_2528);
and U3222 (N_3222,N_2766,N_2919);
xor U3223 (N_3223,N_2845,N_2162);
nand U3224 (N_3224,N_2242,N_2657);
and U3225 (N_3225,N_2295,N_2961);
and U3226 (N_3226,N_2335,N_2826);
nand U3227 (N_3227,N_2857,N_2986);
or U3228 (N_3228,N_2094,N_2918);
nor U3229 (N_3229,N_2033,N_2134);
nor U3230 (N_3230,N_2089,N_2298);
nand U3231 (N_3231,N_2049,N_2892);
xor U3232 (N_3232,N_2476,N_2567);
or U3233 (N_3233,N_2337,N_2929);
and U3234 (N_3234,N_2410,N_2666);
xor U3235 (N_3235,N_2814,N_2258);
nor U3236 (N_3236,N_2939,N_2008);
or U3237 (N_3237,N_2083,N_2754);
and U3238 (N_3238,N_2532,N_2475);
nor U3239 (N_3239,N_2377,N_2282);
and U3240 (N_3240,N_2768,N_2413);
nand U3241 (N_3241,N_2582,N_2267);
and U3242 (N_3242,N_2548,N_2580);
xnor U3243 (N_3243,N_2113,N_2197);
xnor U3244 (N_3244,N_2571,N_2352);
nand U3245 (N_3245,N_2987,N_2654);
xor U3246 (N_3246,N_2655,N_2724);
and U3247 (N_3247,N_2118,N_2880);
xor U3248 (N_3248,N_2840,N_2438);
xnor U3249 (N_3249,N_2979,N_2179);
xnor U3250 (N_3250,N_2471,N_2211);
nor U3251 (N_3251,N_2194,N_2662);
xnor U3252 (N_3252,N_2026,N_2774);
nor U3253 (N_3253,N_2000,N_2398);
xnor U3254 (N_3254,N_2802,N_2180);
nand U3255 (N_3255,N_2394,N_2181);
or U3256 (N_3256,N_2256,N_2393);
nor U3257 (N_3257,N_2708,N_2355);
and U3258 (N_3258,N_2272,N_2916);
or U3259 (N_3259,N_2631,N_2363);
and U3260 (N_3260,N_2167,N_2675);
or U3261 (N_3261,N_2208,N_2801);
nor U3262 (N_3262,N_2954,N_2482);
nor U3263 (N_3263,N_2274,N_2012);
nor U3264 (N_3264,N_2539,N_2406);
nor U3265 (N_3265,N_2871,N_2399);
xor U3266 (N_3266,N_2573,N_2145);
or U3267 (N_3267,N_2040,N_2300);
xnor U3268 (N_3268,N_2777,N_2555);
and U3269 (N_3269,N_2727,N_2443);
and U3270 (N_3270,N_2680,N_2601);
and U3271 (N_3271,N_2316,N_2963);
nand U3272 (N_3272,N_2376,N_2862);
nand U3273 (N_3273,N_2328,N_2990);
nand U3274 (N_3274,N_2132,N_2967);
and U3275 (N_3275,N_2626,N_2150);
and U3276 (N_3276,N_2346,N_2947);
or U3277 (N_3277,N_2022,N_2202);
nand U3278 (N_3278,N_2797,N_2821);
nor U3279 (N_3279,N_2205,N_2015);
xnor U3280 (N_3280,N_2978,N_2561);
xor U3281 (N_3281,N_2023,N_2559);
xor U3282 (N_3282,N_2744,N_2213);
xor U3283 (N_3283,N_2936,N_2686);
nand U3284 (N_3284,N_2585,N_2148);
nor U3285 (N_3285,N_2466,N_2252);
nor U3286 (N_3286,N_2053,N_2069);
nand U3287 (N_3287,N_2285,N_2782);
or U3288 (N_3288,N_2791,N_2356);
and U3289 (N_3289,N_2473,N_2932);
xor U3290 (N_3290,N_2920,N_2324);
and U3291 (N_3291,N_2689,N_2382);
and U3292 (N_3292,N_2643,N_2270);
nor U3293 (N_3293,N_2515,N_2081);
nand U3294 (N_3294,N_2168,N_2177);
nand U3295 (N_3295,N_2909,N_2329);
nand U3296 (N_3296,N_2690,N_2886);
or U3297 (N_3297,N_2914,N_2103);
xnor U3298 (N_3298,N_2338,N_2214);
xnor U3299 (N_3299,N_2726,N_2608);
and U3300 (N_3300,N_2564,N_2340);
nor U3301 (N_3301,N_2086,N_2461);
xor U3302 (N_3302,N_2336,N_2715);
xor U3303 (N_3303,N_2942,N_2215);
xnor U3304 (N_3304,N_2257,N_2535);
nor U3305 (N_3305,N_2278,N_2101);
xor U3306 (N_3306,N_2683,N_2751);
and U3307 (N_3307,N_2511,N_2881);
and U3308 (N_3308,N_2479,N_2854);
nand U3309 (N_3309,N_2116,N_2516);
and U3310 (N_3310,N_2327,N_2577);
nor U3311 (N_3311,N_2709,N_2673);
nor U3312 (N_3312,N_2759,N_2844);
nand U3313 (N_3313,N_2864,N_2882);
nor U3314 (N_3314,N_2304,N_2048);
or U3315 (N_3315,N_2711,N_2610);
or U3316 (N_3316,N_2448,N_2255);
and U3317 (N_3317,N_2628,N_2427);
or U3318 (N_3318,N_2453,N_2538);
nand U3319 (N_3319,N_2139,N_2749);
xor U3320 (N_3320,N_2115,N_2305);
xor U3321 (N_3321,N_2994,N_2489);
nor U3322 (N_3322,N_2603,N_2676);
nor U3323 (N_3323,N_2703,N_2798);
and U3324 (N_3324,N_2907,N_2380);
xor U3325 (N_3325,N_2234,N_2387);
nor U3326 (N_3326,N_2944,N_2813);
nor U3327 (N_3327,N_2509,N_2265);
or U3328 (N_3328,N_2865,N_2849);
nand U3329 (N_3329,N_2071,N_2465);
or U3330 (N_3330,N_2357,N_2719);
nand U3331 (N_3331,N_2810,N_2249);
or U3332 (N_3332,N_2383,N_2212);
or U3333 (N_3333,N_2968,N_2119);
nor U3334 (N_3334,N_2565,N_2632);
and U3335 (N_3335,N_2494,N_2748);
nor U3336 (N_3336,N_2464,N_2714);
xor U3337 (N_3337,N_2606,N_2468);
or U3338 (N_3338,N_2885,N_2973);
or U3339 (N_3339,N_2289,N_2097);
nand U3340 (N_3340,N_2933,N_2123);
nor U3341 (N_3341,N_2144,N_2694);
and U3342 (N_3342,N_2940,N_2842);
or U3343 (N_3343,N_2595,N_2776);
nand U3344 (N_3344,N_2927,N_2757);
or U3345 (N_3345,N_2572,N_2243);
or U3346 (N_3346,N_2856,N_2224);
xor U3347 (N_3347,N_2503,N_2339);
or U3348 (N_3348,N_2440,N_2195);
and U3349 (N_3349,N_2649,N_2470);
nand U3350 (N_3350,N_2011,N_2607);
nor U3351 (N_3351,N_2260,N_2794);
and U3352 (N_3352,N_2638,N_2420);
and U3353 (N_3353,N_2621,N_2521);
xor U3354 (N_3354,N_2426,N_2244);
nand U3355 (N_3355,N_2379,N_2879);
and U3356 (N_3356,N_2303,N_2578);
or U3357 (N_3357,N_2068,N_2891);
and U3358 (N_3358,N_2487,N_2477);
and U3359 (N_3359,N_2838,N_2078);
nor U3360 (N_3360,N_2096,N_2344);
or U3361 (N_3361,N_2203,N_2106);
nor U3362 (N_3362,N_2650,N_2275);
nand U3363 (N_3363,N_2743,N_2019);
nand U3364 (N_3364,N_2486,N_2360);
xor U3365 (N_3365,N_2109,N_2893);
or U3366 (N_3366,N_2251,N_2543);
nor U3367 (N_3367,N_2435,N_2381);
xnor U3368 (N_3368,N_2647,N_2959);
or U3369 (N_3369,N_2396,N_2575);
nor U3370 (N_3370,N_2527,N_2700);
or U3371 (N_3371,N_2812,N_2284);
nor U3372 (N_3372,N_2553,N_2901);
and U3373 (N_3373,N_2688,N_2541);
and U3374 (N_3374,N_2753,N_2226);
nor U3375 (N_3375,N_2483,N_2796);
nand U3376 (N_3376,N_2146,N_2264);
xnor U3377 (N_3377,N_2695,N_2616);
nor U3378 (N_3378,N_2976,N_2735);
and U3379 (N_3379,N_2128,N_2851);
nor U3380 (N_3380,N_2937,N_2788);
nand U3381 (N_3381,N_2299,N_2354);
nor U3382 (N_3382,N_2141,N_2169);
nand U3383 (N_3383,N_2799,N_2104);
and U3384 (N_3384,N_2273,N_2775);
or U3385 (N_3385,N_2320,N_2184);
and U3386 (N_3386,N_2924,N_2005);
and U3387 (N_3387,N_2701,N_2126);
nand U3388 (N_3388,N_2795,N_2699);
and U3389 (N_3389,N_2917,N_2384);
nor U3390 (N_3390,N_2817,N_2767);
and U3391 (N_3391,N_2281,N_2056);
and U3392 (N_3392,N_2030,N_2219);
and U3393 (N_3393,N_2084,N_2341);
nor U3394 (N_3394,N_2395,N_2568);
or U3395 (N_3395,N_2216,N_2374);
or U3396 (N_3396,N_2816,N_2969);
nor U3397 (N_3397,N_2029,N_2858);
xnor U3398 (N_3398,N_2345,N_2792);
xnor U3399 (N_3399,N_2151,N_2192);
or U3400 (N_3400,N_2099,N_2652);
nand U3401 (N_3401,N_2557,N_2518);
or U3402 (N_3402,N_2253,N_2404);
nor U3403 (N_3403,N_2993,N_2065);
or U3404 (N_3404,N_2400,N_2938);
and U3405 (N_3405,N_2611,N_2955);
and U3406 (N_3406,N_2130,N_2313);
or U3407 (N_3407,N_2566,N_2847);
nand U3408 (N_3408,N_2309,N_2704);
and U3409 (N_3409,N_2455,N_2117);
nor U3410 (N_3410,N_2752,N_2190);
nor U3411 (N_3411,N_2306,N_2867);
nor U3412 (N_3412,N_2451,N_2138);
nor U3413 (N_3413,N_2087,N_2391);
or U3414 (N_3414,N_2020,N_2437);
nor U3415 (N_3415,N_2207,N_2246);
and U3416 (N_3416,N_2434,N_2835);
xnor U3417 (N_3417,N_2176,N_2685);
and U3418 (N_3418,N_2839,N_2070);
and U3419 (N_3419,N_2037,N_2240);
or U3420 (N_3420,N_2903,N_2966);
nand U3421 (N_3421,N_2717,N_2370);
nor U3422 (N_3422,N_2672,N_2921);
nand U3423 (N_3423,N_2702,N_2790);
or U3424 (N_3424,N_2204,N_2989);
nor U3425 (N_3425,N_2739,N_2419);
or U3426 (N_3426,N_2627,N_2159);
nand U3427 (N_3427,N_2670,N_2173);
nand U3428 (N_3428,N_2950,N_2547);
xnor U3429 (N_3429,N_2294,N_2403);
nor U3430 (N_3430,N_2142,N_2946);
nand U3431 (N_3431,N_2311,N_2823);
nor U3432 (N_3432,N_2333,N_2549);
nor U3433 (N_3433,N_2825,N_2696);
nand U3434 (N_3434,N_2692,N_2220);
xnor U3435 (N_3435,N_2122,N_2401);
or U3436 (N_3436,N_2925,N_2760);
xor U3437 (N_3437,N_2235,N_2262);
nand U3438 (N_3438,N_2646,N_2596);
xor U3439 (N_3439,N_2592,N_2209);
xnor U3440 (N_3440,N_2723,N_2513);
or U3441 (N_3441,N_2644,N_2943);
xor U3442 (N_3442,N_2525,N_2493);
nand U3443 (N_3443,N_2761,N_2853);
nor U3444 (N_3444,N_2570,N_2868);
or U3445 (N_3445,N_2613,N_2804);
nor U3446 (N_3446,N_2505,N_2599);
xnor U3447 (N_3447,N_2375,N_2415);
nand U3448 (N_3448,N_2740,N_2350);
xnor U3449 (N_3449,N_2873,N_2579);
nor U3450 (N_3450,N_2364,N_2869);
nor U3451 (N_3451,N_2057,N_2077);
nand U3452 (N_3452,N_2588,N_2013);
or U3453 (N_3453,N_2941,N_2004);
and U3454 (N_3454,N_2368,N_2041);
nor U3455 (N_3455,N_2155,N_2463);
nor U3456 (N_3456,N_2897,N_2910);
or U3457 (N_3457,N_2687,N_2172);
nor U3458 (N_3458,N_2147,N_2698);
nand U3459 (N_3459,N_2612,N_2361);
xor U3460 (N_3460,N_2789,N_2560);
nand U3461 (N_3461,N_2984,N_2531);
nand U3462 (N_3462,N_2193,N_2593);
xnor U3463 (N_3463,N_2651,N_2499);
and U3464 (N_3464,N_2861,N_2551);
xor U3465 (N_3465,N_2750,N_2594);
nor U3466 (N_3466,N_2351,N_2054);
nand U3467 (N_3467,N_2010,N_2137);
xnor U3468 (N_3468,N_2831,N_2072);
or U3469 (N_3469,N_2537,N_2502);
or U3470 (N_3470,N_2737,N_2780);
xnor U3471 (N_3471,N_2878,N_2007);
and U3472 (N_3472,N_2430,N_2100);
nor U3473 (N_3473,N_2534,N_2321);
xor U3474 (N_3474,N_2164,N_2498);
nand U3475 (N_3475,N_2684,N_2017);
nor U3476 (N_3476,N_2217,N_2185);
or U3477 (N_3477,N_2423,N_2805);
nand U3478 (N_3478,N_2293,N_2956);
or U3479 (N_3479,N_2624,N_2431);
and U3480 (N_3480,N_2469,N_2314);
nor U3481 (N_3481,N_2523,N_2820);
or U3482 (N_3482,N_2674,N_2785);
nand U3483 (N_3483,N_2452,N_2323);
xor U3484 (N_3484,N_2762,N_2120);
nor U3485 (N_3485,N_2536,N_2678);
and U3486 (N_3486,N_2833,N_2819);
or U3487 (N_3487,N_2237,N_2279);
xnor U3488 (N_3488,N_2957,N_2441);
nor U3489 (N_3489,N_2778,N_2519);
xnor U3490 (N_3490,N_2972,N_2223);
and U3491 (N_3491,N_2786,N_2808);
and U3492 (N_3492,N_2402,N_2658);
or U3493 (N_3493,N_2496,N_2591);
nor U3494 (N_3494,N_2779,N_2707);
nand U3495 (N_3495,N_2459,N_2506);
nor U3496 (N_3496,N_2091,N_2318);
nor U3497 (N_3497,N_2481,N_2906);
nand U3498 (N_3498,N_2075,N_2772);
nor U3499 (N_3499,N_2731,N_2922);
xnor U3500 (N_3500,N_2424,N_2509);
nand U3501 (N_3501,N_2255,N_2358);
or U3502 (N_3502,N_2074,N_2206);
xnor U3503 (N_3503,N_2576,N_2925);
and U3504 (N_3504,N_2135,N_2110);
nand U3505 (N_3505,N_2188,N_2719);
and U3506 (N_3506,N_2722,N_2649);
nand U3507 (N_3507,N_2349,N_2522);
nand U3508 (N_3508,N_2846,N_2126);
nor U3509 (N_3509,N_2574,N_2533);
or U3510 (N_3510,N_2681,N_2754);
nor U3511 (N_3511,N_2746,N_2361);
or U3512 (N_3512,N_2112,N_2250);
nand U3513 (N_3513,N_2293,N_2938);
xnor U3514 (N_3514,N_2005,N_2573);
xor U3515 (N_3515,N_2565,N_2659);
or U3516 (N_3516,N_2154,N_2736);
nand U3517 (N_3517,N_2160,N_2372);
nor U3518 (N_3518,N_2258,N_2163);
nor U3519 (N_3519,N_2734,N_2532);
xnor U3520 (N_3520,N_2492,N_2677);
xnor U3521 (N_3521,N_2334,N_2828);
and U3522 (N_3522,N_2916,N_2145);
nand U3523 (N_3523,N_2528,N_2100);
and U3524 (N_3524,N_2438,N_2728);
nor U3525 (N_3525,N_2855,N_2688);
or U3526 (N_3526,N_2363,N_2362);
nor U3527 (N_3527,N_2842,N_2232);
or U3528 (N_3528,N_2592,N_2571);
nand U3529 (N_3529,N_2317,N_2791);
and U3530 (N_3530,N_2182,N_2093);
nand U3531 (N_3531,N_2500,N_2216);
or U3532 (N_3532,N_2108,N_2389);
and U3533 (N_3533,N_2024,N_2869);
xor U3534 (N_3534,N_2471,N_2723);
or U3535 (N_3535,N_2533,N_2027);
and U3536 (N_3536,N_2255,N_2041);
or U3537 (N_3537,N_2461,N_2725);
nand U3538 (N_3538,N_2556,N_2867);
or U3539 (N_3539,N_2152,N_2143);
and U3540 (N_3540,N_2074,N_2597);
or U3541 (N_3541,N_2090,N_2770);
xnor U3542 (N_3542,N_2888,N_2372);
xnor U3543 (N_3543,N_2830,N_2072);
nor U3544 (N_3544,N_2294,N_2378);
or U3545 (N_3545,N_2826,N_2258);
and U3546 (N_3546,N_2194,N_2102);
or U3547 (N_3547,N_2750,N_2297);
or U3548 (N_3548,N_2387,N_2330);
nand U3549 (N_3549,N_2067,N_2463);
nand U3550 (N_3550,N_2695,N_2345);
and U3551 (N_3551,N_2759,N_2647);
and U3552 (N_3552,N_2326,N_2111);
nor U3553 (N_3553,N_2292,N_2980);
xnor U3554 (N_3554,N_2981,N_2028);
nor U3555 (N_3555,N_2465,N_2697);
or U3556 (N_3556,N_2544,N_2589);
or U3557 (N_3557,N_2686,N_2646);
xnor U3558 (N_3558,N_2011,N_2068);
nand U3559 (N_3559,N_2425,N_2166);
nor U3560 (N_3560,N_2120,N_2793);
and U3561 (N_3561,N_2148,N_2179);
and U3562 (N_3562,N_2488,N_2974);
nand U3563 (N_3563,N_2899,N_2362);
nor U3564 (N_3564,N_2170,N_2319);
nand U3565 (N_3565,N_2232,N_2060);
xnor U3566 (N_3566,N_2424,N_2915);
or U3567 (N_3567,N_2886,N_2650);
nand U3568 (N_3568,N_2874,N_2115);
nor U3569 (N_3569,N_2803,N_2496);
nor U3570 (N_3570,N_2197,N_2226);
nor U3571 (N_3571,N_2629,N_2723);
xor U3572 (N_3572,N_2077,N_2257);
nor U3573 (N_3573,N_2183,N_2809);
nor U3574 (N_3574,N_2720,N_2613);
or U3575 (N_3575,N_2682,N_2417);
and U3576 (N_3576,N_2502,N_2047);
nand U3577 (N_3577,N_2256,N_2556);
nand U3578 (N_3578,N_2652,N_2995);
or U3579 (N_3579,N_2697,N_2933);
nand U3580 (N_3580,N_2486,N_2165);
nor U3581 (N_3581,N_2324,N_2806);
or U3582 (N_3582,N_2673,N_2490);
nor U3583 (N_3583,N_2586,N_2089);
nor U3584 (N_3584,N_2491,N_2042);
nor U3585 (N_3585,N_2146,N_2459);
nor U3586 (N_3586,N_2861,N_2391);
nor U3587 (N_3587,N_2652,N_2145);
nand U3588 (N_3588,N_2910,N_2619);
and U3589 (N_3589,N_2645,N_2176);
xnor U3590 (N_3590,N_2428,N_2075);
and U3591 (N_3591,N_2802,N_2192);
and U3592 (N_3592,N_2790,N_2236);
or U3593 (N_3593,N_2967,N_2865);
nor U3594 (N_3594,N_2540,N_2862);
xor U3595 (N_3595,N_2755,N_2550);
xor U3596 (N_3596,N_2862,N_2231);
nor U3597 (N_3597,N_2640,N_2813);
or U3598 (N_3598,N_2988,N_2320);
nand U3599 (N_3599,N_2678,N_2609);
xnor U3600 (N_3600,N_2462,N_2451);
nor U3601 (N_3601,N_2146,N_2059);
or U3602 (N_3602,N_2124,N_2532);
or U3603 (N_3603,N_2815,N_2982);
xnor U3604 (N_3604,N_2185,N_2444);
xnor U3605 (N_3605,N_2071,N_2984);
nand U3606 (N_3606,N_2447,N_2249);
or U3607 (N_3607,N_2023,N_2921);
xnor U3608 (N_3608,N_2531,N_2831);
nor U3609 (N_3609,N_2870,N_2954);
xor U3610 (N_3610,N_2364,N_2455);
or U3611 (N_3611,N_2128,N_2251);
xor U3612 (N_3612,N_2369,N_2138);
nand U3613 (N_3613,N_2732,N_2822);
xnor U3614 (N_3614,N_2157,N_2936);
nand U3615 (N_3615,N_2860,N_2179);
nor U3616 (N_3616,N_2161,N_2074);
and U3617 (N_3617,N_2519,N_2483);
and U3618 (N_3618,N_2615,N_2899);
nand U3619 (N_3619,N_2865,N_2643);
and U3620 (N_3620,N_2133,N_2776);
nand U3621 (N_3621,N_2665,N_2070);
xnor U3622 (N_3622,N_2114,N_2931);
xor U3623 (N_3623,N_2643,N_2653);
xnor U3624 (N_3624,N_2732,N_2695);
or U3625 (N_3625,N_2910,N_2231);
xor U3626 (N_3626,N_2338,N_2473);
or U3627 (N_3627,N_2922,N_2164);
nand U3628 (N_3628,N_2440,N_2818);
or U3629 (N_3629,N_2115,N_2821);
nand U3630 (N_3630,N_2941,N_2513);
nand U3631 (N_3631,N_2598,N_2781);
xor U3632 (N_3632,N_2483,N_2335);
xor U3633 (N_3633,N_2389,N_2556);
or U3634 (N_3634,N_2248,N_2662);
nand U3635 (N_3635,N_2249,N_2242);
nand U3636 (N_3636,N_2360,N_2898);
nor U3637 (N_3637,N_2504,N_2692);
and U3638 (N_3638,N_2509,N_2698);
or U3639 (N_3639,N_2789,N_2620);
xnor U3640 (N_3640,N_2247,N_2386);
nor U3641 (N_3641,N_2212,N_2214);
nor U3642 (N_3642,N_2487,N_2251);
nand U3643 (N_3643,N_2825,N_2843);
and U3644 (N_3644,N_2157,N_2123);
and U3645 (N_3645,N_2425,N_2495);
or U3646 (N_3646,N_2407,N_2694);
and U3647 (N_3647,N_2755,N_2534);
nor U3648 (N_3648,N_2927,N_2070);
and U3649 (N_3649,N_2787,N_2769);
or U3650 (N_3650,N_2819,N_2996);
nand U3651 (N_3651,N_2073,N_2071);
xnor U3652 (N_3652,N_2780,N_2175);
or U3653 (N_3653,N_2384,N_2987);
and U3654 (N_3654,N_2855,N_2144);
xnor U3655 (N_3655,N_2751,N_2458);
or U3656 (N_3656,N_2818,N_2510);
nor U3657 (N_3657,N_2977,N_2928);
xnor U3658 (N_3658,N_2857,N_2609);
nand U3659 (N_3659,N_2557,N_2445);
nor U3660 (N_3660,N_2787,N_2598);
nand U3661 (N_3661,N_2117,N_2021);
nor U3662 (N_3662,N_2140,N_2402);
nand U3663 (N_3663,N_2401,N_2701);
or U3664 (N_3664,N_2058,N_2064);
xor U3665 (N_3665,N_2112,N_2684);
and U3666 (N_3666,N_2251,N_2672);
nor U3667 (N_3667,N_2557,N_2639);
and U3668 (N_3668,N_2369,N_2377);
xnor U3669 (N_3669,N_2089,N_2883);
nor U3670 (N_3670,N_2278,N_2610);
nand U3671 (N_3671,N_2421,N_2278);
and U3672 (N_3672,N_2929,N_2067);
xnor U3673 (N_3673,N_2095,N_2003);
and U3674 (N_3674,N_2272,N_2506);
xor U3675 (N_3675,N_2080,N_2827);
and U3676 (N_3676,N_2538,N_2306);
nand U3677 (N_3677,N_2131,N_2067);
or U3678 (N_3678,N_2137,N_2128);
or U3679 (N_3679,N_2641,N_2687);
or U3680 (N_3680,N_2850,N_2765);
nor U3681 (N_3681,N_2427,N_2954);
nor U3682 (N_3682,N_2994,N_2701);
or U3683 (N_3683,N_2733,N_2878);
nor U3684 (N_3684,N_2277,N_2583);
xor U3685 (N_3685,N_2911,N_2517);
or U3686 (N_3686,N_2942,N_2547);
and U3687 (N_3687,N_2728,N_2138);
or U3688 (N_3688,N_2300,N_2239);
and U3689 (N_3689,N_2397,N_2741);
and U3690 (N_3690,N_2436,N_2639);
xnor U3691 (N_3691,N_2909,N_2021);
and U3692 (N_3692,N_2118,N_2367);
nor U3693 (N_3693,N_2461,N_2212);
xnor U3694 (N_3694,N_2144,N_2189);
nand U3695 (N_3695,N_2856,N_2468);
nor U3696 (N_3696,N_2448,N_2890);
nor U3697 (N_3697,N_2880,N_2576);
or U3698 (N_3698,N_2242,N_2998);
nand U3699 (N_3699,N_2569,N_2899);
nor U3700 (N_3700,N_2461,N_2113);
xnor U3701 (N_3701,N_2626,N_2326);
nor U3702 (N_3702,N_2574,N_2767);
and U3703 (N_3703,N_2051,N_2571);
nor U3704 (N_3704,N_2467,N_2001);
and U3705 (N_3705,N_2881,N_2264);
xnor U3706 (N_3706,N_2281,N_2087);
nor U3707 (N_3707,N_2649,N_2749);
or U3708 (N_3708,N_2588,N_2165);
and U3709 (N_3709,N_2176,N_2903);
and U3710 (N_3710,N_2352,N_2354);
and U3711 (N_3711,N_2606,N_2012);
and U3712 (N_3712,N_2351,N_2857);
and U3713 (N_3713,N_2480,N_2188);
nor U3714 (N_3714,N_2285,N_2904);
xnor U3715 (N_3715,N_2646,N_2592);
nor U3716 (N_3716,N_2191,N_2705);
xnor U3717 (N_3717,N_2601,N_2866);
nor U3718 (N_3718,N_2131,N_2265);
nand U3719 (N_3719,N_2332,N_2999);
xor U3720 (N_3720,N_2586,N_2130);
nor U3721 (N_3721,N_2122,N_2263);
or U3722 (N_3722,N_2104,N_2415);
nand U3723 (N_3723,N_2584,N_2945);
nand U3724 (N_3724,N_2013,N_2615);
xnor U3725 (N_3725,N_2156,N_2783);
xor U3726 (N_3726,N_2256,N_2047);
nor U3727 (N_3727,N_2327,N_2698);
nor U3728 (N_3728,N_2157,N_2309);
and U3729 (N_3729,N_2842,N_2667);
and U3730 (N_3730,N_2536,N_2377);
xor U3731 (N_3731,N_2215,N_2342);
xor U3732 (N_3732,N_2288,N_2875);
nand U3733 (N_3733,N_2416,N_2729);
nand U3734 (N_3734,N_2477,N_2914);
and U3735 (N_3735,N_2281,N_2511);
xnor U3736 (N_3736,N_2138,N_2051);
nor U3737 (N_3737,N_2533,N_2435);
xor U3738 (N_3738,N_2291,N_2110);
nor U3739 (N_3739,N_2470,N_2960);
or U3740 (N_3740,N_2686,N_2973);
or U3741 (N_3741,N_2504,N_2680);
xor U3742 (N_3742,N_2408,N_2934);
or U3743 (N_3743,N_2473,N_2365);
or U3744 (N_3744,N_2731,N_2408);
nand U3745 (N_3745,N_2994,N_2674);
or U3746 (N_3746,N_2853,N_2564);
nand U3747 (N_3747,N_2741,N_2830);
or U3748 (N_3748,N_2054,N_2677);
or U3749 (N_3749,N_2113,N_2492);
nand U3750 (N_3750,N_2210,N_2198);
and U3751 (N_3751,N_2476,N_2418);
or U3752 (N_3752,N_2074,N_2573);
and U3753 (N_3753,N_2071,N_2077);
nand U3754 (N_3754,N_2144,N_2403);
or U3755 (N_3755,N_2771,N_2012);
xnor U3756 (N_3756,N_2845,N_2588);
xor U3757 (N_3757,N_2105,N_2739);
and U3758 (N_3758,N_2786,N_2601);
and U3759 (N_3759,N_2312,N_2850);
nor U3760 (N_3760,N_2130,N_2159);
or U3761 (N_3761,N_2219,N_2817);
xnor U3762 (N_3762,N_2634,N_2175);
nor U3763 (N_3763,N_2108,N_2128);
and U3764 (N_3764,N_2497,N_2189);
and U3765 (N_3765,N_2337,N_2409);
and U3766 (N_3766,N_2107,N_2526);
and U3767 (N_3767,N_2563,N_2520);
xnor U3768 (N_3768,N_2988,N_2589);
nor U3769 (N_3769,N_2404,N_2730);
nand U3770 (N_3770,N_2947,N_2584);
xnor U3771 (N_3771,N_2459,N_2047);
xnor U3772 (N_3772,N_2204,N_2804);
and U3773 (N_3773,N_2109,N_2879);
or U3774 (N_3774,N_2745,N_2809);
and U3775 (N_3775,N_2578,N_2196);
or U3776 (N_3776,N_2883,N_2985);
or U3777 (N_3777,N_2389,N_2524);
or U3778 (N_3778,N_2087,N_2266);
or U3779 (N_3779,N_2691,N_2557);
nand U3780 (N_3780,N_2292,N_2510);
and U3781 (N_3781,N_2394,N_2682);
and U3782 (N_3782,N_2935,N_2675);
and U3783 (N_3783,N_2695,N_2625);
and U3784 (N_3784,N_2585,N_2314);
xnor U3785 (N_3785,N_2789,N_2493);
xor U3786 (N_3786,N_2430,N_2343);
nand U3787 (N_3787,N_2670,N_2750);
xnor U3788 (N_3788,N_2848,N_2772);
or U3789 (N_3789,N_2728,N_2661);
or U3790 (N_3790,N_2427,N_2038);
nor U3791 (N_3791,N_2768,N_2204);
or U3792 (N_3792,N_2414,N_2342);
and U3793 (N_3793,N_2968,N_2607);
and U3794 (N_3794,N_2558,N_2743);
nand U3795 (N_3795,N_2729,N_2839);
and U3796 (N_3796,N_2230,N_2144);
and U3797 (N_3797,N_2208,N_2599);
nand U3798 (N_3798,N_2266,N_2471);
xor U3799 (N_3799,N_2835,N_2487);
and U3800 (N_3800,N_2898,N_2027);
or U3801 (N_3801,N_2008,N_2762);
nor U3802 (N_3802,N_2633,N_2596);
nand U3803 (N_3803,N_2034,N_2496);
nor U3804 (N_3804,N_2384,N_2507);
and U3805 (N_3805,N_2126,N_2867);
and U3806 (N_3806,N_2929,N_2833);
nor U3807 (N_3807,N_2190,N_2949);
and U3808 (N_3808,N_2434,N_2588);
or U3809 (N_3809,N_2978,N_2887);
or U3810 (N_3810,N_2792,N_2829);
or U3811 (N_3811,N_2325,N_2453);
xnor U3812 (N_3812,N_2512,N_2102);
or U3813 (N_3813,N_2393,N_2043);
or U3814 (N_3814,N_2068,N_2925);
nand U3815 (N_3815,N_2861,N_2129);
or U3816 (N_3816,N_2808,N_2146);
nand U3817 (N_3817,N_2890,N_2603);
xor U3818 (N_3818,N_2021,N_2635);
xnor U3819 (N_3819,N_2657,N_2108);
and U3820 (N_3820,N_2907,N_2122);
nor U3821 (N_3821,N_2651,N_2245);
nor U3822 (N_3822,N_2092,N_2111);
nor U3823 (N_3823,N_2663,N_2671);
xnor U3824 (N_3824,N_2291,N_2826);
xnor U3825 (N_3825,N_2188,N_2256);
xor U3826 (N_3826,N_2431,N_2261);
or U3827 (N_3827,N_2776,N_2574);
nand U3828 (N_3828,N_2193,N_2372);
xnor U3829 (N_3829,N_2418,N_2957);
nor U3830 (N_3830,N_2649,N_2192);
nand U3831 (N_3831,N_2087,N_2890);
or U3832 (N_3832,N_2814,N_2558);
nor U3833 (N_3833,N_2028,N_2000);
xor U3834 (N_3834,N_2948,N_2039);
xnor U3835 (N_3835,N_2853,N_2652);
xor U3836 (N_3836,N_2051,N_2813);
nand U3837 (N_3837,N_2112,N_2730);
and U3838 (N_3838,N_2506,N_2178);
and U3839 (N_3839,N_2222,N_2888);
or U3840 (N_3840,N_2934,N_2596);
or U3841 (N_3841,N_2743,N_2099);
or U3842 (N_3842,N_2829,N_2141);
nand U3843 (N_3843,N_2292,N_2924);
xor U3844 (N_3844,N_2605,N_2283);
nand U3845 (N_3845,N_2025,N_2443);
nand U3846 (N_3846,N_2233,N_2024);
or U3847 (N_3847,N_2982,N_2885);
and U3848 (N_3848,N_2262,N_2667);
or U3849 (N_3849,N_2561,N_2492);
or U3850 (N_3850,N_2425,N_2701);
nor U3851 (N_3851,N_2631,N_2572);
and U3852 (N_3852,N_2190,N_2698);
nor U3853 (N_3853,N_2637,N_2727);
or U3854 (N_3854,N_2171,N_2285);
and U3855 (N_3855,N_2789,N_2184);
and U3856 (N_3856,N_2027,N_2330);
and U3857 (N_3857,N_2817,N_2552);
xnor U3858 (N_3858,N_2928,N_2960);
and U3859 (N_3859,N_2964,N_2364);
xor U3860 (N_3860,N_2150,N_2047);
xor U3861 (N_3861,N_2620,N_2844);
and U3862 (N_3862,N_2399,N_2964);
nand U3863 (N_3863,N_2788,N_2022);
xnor U3864 (N_3864,N_2313,N_2569);
and U3865 (N_3865,N_2865,N_2820);
xor U3866 (N_3866,N_2277,N_2032);
xor U3867 (N_3867,N_2548,N_2067);
and U3868 (N_3868,N_2932,N_2460);
and U3869 (N_3869,N_2516,N_2709);
or U3870 (N_3870,N_2272,N_2492);
xnor U3871 (N_3871,N_2784,N_2542);
and U3872 (N_3872,N_2689,N_2869);
and U3873 (N_3873,N_2048,N_2261);
nand U3874 (N_3874,N_2722,N_2272);
xnor U3875 (N_3875,N_2757,N_2366);
nor U3876 (N_3876,N_2707,N_2432);
nor U3877 (N_3877,N_2634,N_2104);
nor U3878 (N_3878,N_2663,N_2523);
nand U3879 (N_3879,N_2578,N_2277);
nor U3880 (N_3880,N_2936,N_2236);
or U3881 (N_3881,N_2027,N_2711);
or U3882 (N_3882,N_2414,N_2103);
nand U3883 (N_3883,N_2307,N_2961);
xor U3884 (N_3884,N_2503,N_2294);
or U3885 (N_3885,N_2939,N_2202);
or U3886 (N_3886,N_2552,N_2934);
xnor U3887 (N_3887,N_2050,N_2794);
xor U3888 (N_3888,N_2596,N_2353);
and U3889 (N_3889,N_2544,N_2563);
nand U3890 (N_3890,N_2157,N_2812);
or U3891 (N_3891,N_2548,N_2453);
xnor U3892 (N_3892,N_2279,N_2158);
xor U3893 (N_3893,N_2229,N_2906);
nor U3894 (N_3894,N_2922,N_2399);
and U3895 (N_3895,N_2035,N_2942);
and U3896 (N_3896,N_2644,N_2650);
and U3897 (N_3897,N_2756,N_2944);
nand U3898 (N_3898,N_2770,N_2915);
and U3899 (N_3899,N_2228,N_2915);
or U3900 (N_3900,N_2730,N_2465);
or U3901 (N_3901,N_2789,N_2563);
nand U3902 (N_3902,N_2781,N_2251);
or U3903 (N_3903,N_2596,N_2470);
xor U3904 (N_3904,N_2317,N_2754);
and U3905 (N_3905,N_2747,N_2169);
xnor U3906 (N_3906,N_2071,N_2493);
nor U3907 (N_3907,N_2515,N_2444);
or U3908 (N_3908,N_2865,N_2590);
or U3909 (N_3909,N_2087,N_2902);
or U3910 (N_3910,N_2799,N_2524);
and U3911 (N_3911,N_2419,N_2764);
nand U3912 (N_3912,N_2929,N_2951);
or U3913 (N_3913,N_2216,N_2392);
xor U3914 (N_3914,N_2536,N_2909);
and U3915 (N_3915,N_2786,N_2815);
or U3916 (N_3916,N_2087,N_2212);
nand U3917 (N_3917,N_2076,N_2379);
and U3918 (N_3918,N_2464,N_2103);
or U3919 (N_3919,N_2915,N_2064);
or U3920 (N_3920,N_2511,N_2433);
or U3921 (N_3921,N_2619,N_2725);
or U3922 (N_3922,N_2034,N_2321);
or U3923 (N_3923,N_2171,N_2978);
xnor U3924 (N_3924,N_2044,N_2346);
nand U3925 (N_3925,N_2772,N_2345);
nand U3926 (N_3926,N_2391,N_2116);
xnor U3927 (N_3927,N_2031,N_2216);
nor U3928 (N_3928,N_2621,N_2756);
nor U3929 (N_3929,N_2310,N_2350);
xor U3930 (N_3930,N_2415,N_2605);
xnor U3931 (N_3931,N_2349,N_2989);
or U3932 (N_3932,N_2069,N_2259);
xor U3933 (N_3933,N_2977,N_2509);
or U3934 (N_3934,N_2566,N_2191);
nand U3935 (N_3935,N_2407,N_2114);
xor U3936 (N_3936,N_2054,N_2420);
nand U3937 (N_3937,N_2429,N_2889);
or U3938 (N_3938,N_2215,N_2768);
or U3939 (N_3939,N_2443,N_2192);
nand U3940 (N_3940,N_2875,N_2795);
or U3941 (N_3941,N_2321,N_2634);
nor U3942 (N_3942,N_2141,N_2313);
nor U3943 (N_3943,N_2946,N_2083);
nor U3944 (N_3944,N_2445,N_2435);
xnor U3945 (N_3945,N_2949,N_2622);
nand U3946 (N_3946,N_2055,N_2612);
nor U3947 (N_3947,N_2327,N_2748);
xnor U3948 (N_3948,N_2343,N_2500);
nor U3949 (N_3949,N_2310,N_2837);
or U3950 (N_3950,N_2536,N_2291);
nor U3951 (N_3951,N_2811,N_2738);
nor U3952 (N_3952,N_2198,N_2348);
xnor U3953 (N_3953,N_2497,N_2066);
or U3954 (N_3954,N_2152,N_2222);
nand U3955 (N_3955,N_2819,N_2934);
xnor U3956 (N_3956,N_2767,N_2334);
and U3957 (N_3957,N_2861,N_2672);
or U3958 (N_3958,N_2753,N_2974);
or U3959 (N_3959,N_2806,N_2197);
or U3960 (N_3960,N_2572,N_2855);
nand U3961 (N_3961,N_2016,N_2527);
and U3962 (N_3962,N_2053,N_2587);
xor U3963 (N_3963,N_2880,N_2642);
nor U3964 (N_3964,N_2238,N_2967);
and U3965 (N_3965,N_2698,N_2553);
and U3966 (N_3966,N_2962,N_2383);
and U3967 (N_3967,N_2210,N_2880);
xnor U3968 (N_3968,N_2318,N_2344);
nor U3969 (N_3969,N_2195,N_2121);
nor U3970 (N_3970,N_2497,N_2306);
xnor U3971 (N_3971,N_2617,N_2747);
nor U3972 (N_3972,N_2389,N_2617);
and U3973 (N_3973,N_2972,N_2786);
nand U3974 (N_3974,N_2425,N_2900);
nand U3975 (N_3975,N_2083,N_2642);
or U3976 (N_3976,N_2362,N_2129);
or U3977 (N_3977,N_2742,N_2984);
xnor U3978 (N_3978,N_2425,N_2865);
nand U3979 (N_3979,N_2266,N_2892);
or U3980 (N_3980,N_2828,N_2895);
and U3981 (N_3981,N_2748,N_2165);
and U3982 (N_3982,N_2259,N_2027);
nand U3983 (N_3983,N_2120,N_2783);
xor U3984 (N_3984,N_2087,N_2010);
nor U3985 (N_3985,N_2072,N_2892);
or U3986 (N_3986,N_2853,N_2914);
or U3987 (N_3987,N_2503,N_2965);
xnor U3988 (N_3988,N_2787,N_2003);
nor U3989 (N_3989,N_2407,N_2075);
or U3990 (N_3990,N_2754,N_2496);
xnor U3991 (N_3991,N_2221,N_2526);
nor U3992 (N_3992,N_2259,N_2801);
nand U3993 (N_3993,N_2747,N_2150);
or U3994 (N_3994,N_2570,N_2460);
and U3995 (N_3995,N_2015,N_2771);
or U3996 (N_3996,N_2565,N_2530);
nor U3997 (N_3997,N_2601,N_2332);
nor U3998 (N_3998,N_2532,N_2045);
xor U3999 (N_3999,N_2337,N_2999);
xor U4000 (N_4000,N_3613,N_3716);
nor U4001 (N_4001,N_3990,N_3538);
or U4002 (N_4002,N_3147,N_3643);
and U4003 (N_4003,N_3675,N_3073);
nor U4004 (N_4004,N_3580,N_3033);
nor U4005 (N_4005,N_3660,N_3857);
nand U4006 (N_4006,N_3091,N_3721);
nor U4007 (N_4007,N_3676,N_3395);
nand U4008 (N_4008,N_3875,N_3911);
nand U4009 (N_4009,N_3898,N_3552);
or U4010 (N_4010,N_3274,N_3119);
nor U4011 (N_4011,N_3399,N_3539);
nand U4012 (N_4012,N_3049,N_3589);
and U4013 (N_4013,N_3601,N_3175);
and U4014 (N_4014,N_3217,N_3176);
xor U4015 (N_4015,N_3725,N_3663);
xor U4016 (N_4016,N_3062,N_3684);
and U4017 (N_4017,N_3201,N_3326);
xnor U4018 (N_4018,N_3645,N_3310);
or U4019 (N_4019,N_3529,N_3603);
nor U4020 (N_4020,N_3377,N_3807);
nand U4021 (N_4021,N_3456,N_3311);
and U4022 (N_4022,N_3523,N_3141);
nand U4023 (N_4023,N_3697,N_3789);
nand U4024 (N_4024,N_3639,N_3629);
or U4025 (N_4025,N_3045,N_3080);
xnor U4026 (N_4026,N_3396,N_3886);
xnor U4027 (N_4027,N_3671,N_3350);
or U4028 (N_4028,N_3787,N_3473);
or U4029 (N_4029,N_3705,N_3347);
and U4030 (N_4030,N_3468,N_3731);
and U4031 (N_4031,N_3734,N_3284);
and U4032 (N_4032,N_3451,N_3851);
and U4033 (N_4033,N_3095,N_3391);
or U4034 (N_4034,N_3830,N_3803);
and U4035 (N_4035,N_3914,N_3328);
or U4036 (N_4036,N_3124,N_3942);
nand U4037 (N_4037,N_3460,N_3046);
xor U4038 (N_4038,N_3016,N_3753);
nor U4039 (N_4039,N_3402,N_3113);
and U4040 (N_4040,N_3883,N_3504);
nand U4041 (N_4041,N_3598,N_3491);
nor U4042 (N_4042,N_3024,N_3506);
nand U4043 (N_4043,N_3836,N_3574);
nand U4044 (N_4044,N_3696,N_3588);
or U4045 (N_4045,N_3145,N_3405);
nor U4046 (N_4046,N_3439,N_3184);
xor U4047 (N_4047,N_3779,N_3322);
nand U4048 (N_4048,N_3748,N_3125);
nand U4049 (N_4049,N_3250,N_3723);
xor U4050 (N_4050,N_3567,N_3011);
nor U4051 (N_4051,N_3679,N_3832);
nor U4052 (N_4052,N_3148,N_3013);
or U4053 (N_4053,N_3724,N_3693);
nor U4054 (N_4054,N_3888,N_3963);
xor U4055 (N_4055,N_3711,N_3253);
xnor U4056 (N_4056,N_3861,N_3076);
and U4057 (N_4057,N_3241,N_3082);
and U4058 (N_4058,N_3561,N_3925);
and U4059 (N_4059,N_3882,N_3582);
nand U4060 (N_4060,N_3710,N_3386);
nand U4061 (N_4061,N_3433,N_3918);
nand U4062 (N_4062,N_3324,N_3901);
nor U4063 (N_4063,N_3564,N_3780);
or U4064 (N_4064,N_3251,N_3577);
and U4065 (N_4065,N_3797,N_3237);
nand U4066 (N_4066,N_3855,N_3784);
or U4067 (N_4067,N_3166,N_3672);
nor U4068 (N_4068,N_3014,N_3945);
or U4069 (N_4069,N_3902,N_3246);
and U4070 (N_4070,N_3955,N_3407);
or U4071 (N_4071,N_3820,N_3615);
nand U4072 (N_4072,N_3298,N_3531);
xnor U4073 (N_4073,N_3265,N_3150);
and U4074 (N_4074,N_3075,N_3680);
or U4075 (N_4075,N_3490,N_3171);
or U4076 (N_4076,N_3065,N_3088);
xnor U4077 (N_4077,N_3694,N_3651);
or U4078 (N_4078,N_3112,N_3231);
xor U4079 (N_4079,N_3656,N_3794);
nor U4080 (N_4080,N_3876,N_3922);
nand U4081 (N_4081,N_3801,N_3604);
nor U4082 (N_4082,N_3722,N_3750);
or U4083 (N_4083,N_3267,N_3781);
and U4084 (N_4084,N_3181,N_3293);
or U4085 (N_4085,N_3444,N_3833);
nand U4086 (N_4086,N_3525,N_3636);
xnor U4087 (N_4087,N_3652,N_3870);
nor U4088 (N_4088,N_3866,N_3685);
xnor U4089 (N_4089,N_3069,N_3039);
nor U4090 (N_4090,N_3488,N_3501);
or U4091 (N_4091,N_3101,N_3634);
or U4092 (N_4092,N_3965,N_3631);
or U4093 (N_4093,N_3064,N_3387);
xor U4094 (N_4094,N_3332,N_3223);
xnor U4095 (N_4095,N_3834,N_3686);
and U4096 (N_4096,N_3149,N_3212);
nor U4097 (N_4097,N_3244,N_3996);
nand U4098 (N_4098,N_3924,N_3550);
xor U4099 (N_4099,N_3143,N_3079);
and U4100 (N_4100,N_3873,N_3971);
nor U4101 (N_4101,N_3524,N_3568);
nor U4102 (N_4102,N_3819,N_3969);
and U4103 (N_4103,N_3053,N_3499);
nor U4104 (N_4104,N_3445,N_3817);
and U4105 (N_4105,N_3454,N_3678);
nand U4106 (N_4106,N_3313,N_3554);
and U4107 (N_4107,N_3983,N_3160);
nand U4108 (N_4108,N_3247,N_3520);
or U4109 (N_4109,N_3584,N_3626);
nor U4110 (N_4110,N_3430,N_3667);
nand U4111 (N_4111,N_3742,N_3893);
or U4112 (N_4112,N_3459,N_3607);
and U4113 (N_4113,N_3170,N_3382);
xor U4114 (N_4114,N_3348,N_3361);
or U4115 (N_4115,N_3031,N_3349);
nand U4116 (N_4116,N_3597,N_3342);
and U4117 (N_4117,N_3432,N_3106);
and U4118 (N_4118,N_3336,N_3188);
and U4119 (N_4119,N_3135,N_3010);
xor U4120 (N_4120,N_3744,N_3687);
nand U4121 (N_4121,N_3042,N_3923);
xnor U4122 (N_4122,N_3989,N_3300);
and U4123 (N_4123,N_3828,N_3885);
or U4124 (N_4124,N_3436,N_3102);
and U4125 (N_4125,N_3573,N_3758);
nor U4126 (N_4126,N_3540,N_3920);
nor U4127 (N_4127,N_3163,N_3221);
and U4128 (N_4128,N_3280,N_3400);
nor U4129 (N_4129,N_3899,N_3533);
nand U4130 (N_4130,N_3610,N_3715);
or U4131 (N_4131,N_3470,N_3627);
nor U4132 (N_4132,N_3835,N_3358);
nor U4133 (N_4133,N_3822,N_3999);
nor U4134 (N_4134,N_3994,N_3172);
nand U4135 (N_4135,N_3966,N_3174);
or U4136 (N_4136,N_3976,N_3926);
nor U4137 (N_4137,N_3662,N_3500);
nor U4138 (N_4138,N_3292,N_3986);
or U4139 (N_4139,N_3952,N_3435);
and U4140 (N_4140,N_3559,N_3738);
xnor U4141 (N_4141,N_3853,N_3973);
or U4142 (N_4142,N_3850,N_3058);
nor U4143 (N_4143,N_3425,N_3424);
or U4144 (N_4144,N_3892,N_3354);
or U4145 (N_4145,N_3616,N_3000);
or U4146 (N_4146,N_3213,N_3205);
nand U4147 (N_4147,N_3369,N_3890);
nand U4148 (N_4148,N_3908,N_3129);
nand U4149 (N_4149,N_3475,N_3256);
nor U4150 (N_4150,N_3630,N_3957);
or U4151 (N_4151,N_3263,N_3620);
nand U4152 (N_4152,N_3811,N_3545);
xnor U4153 (N_4153,N_3829,N_3798);
nor U4154 (N_4154,N_3547,N_3944);
nor U4155 (N_4155,N_3617,N_3094);
xor U4156 (N_4156,N_3123,N_3596);
nor U4157 (N_4157,N_3465,N_3809);
xnor U4158 (N_4158,N_3390,N_3437);
or U4159 (N_4159,N_3704,N_3192);
xor U4160 (N_4160,N_3216,N_3299);
nand U4161 (N_4161,N_3489,N_3345);
xnor U4162 (N_4162,N_3412,N_3070);
or U4163 (N_4163,N_3974,N_3814);
xor U4164 (N_4164,N_3442,N_3578);
and U4165 (N_4165,N_3288,N_3305);
nor U4166 (N_4166,N_3674,N_3002);
or U4167 (N_4167,N_3270,N_3153);
nand U4168 (N_4168,N_3553,N_3230);
nor U4169 (N_4169,N_3340,N_3831);
xnor U4170 (N_4170,N_3019,N_3417);
or U4171 (N_4171,N_3747,N_3493);
and U4172 (N_4172,N_3931,N_3796);
nor U4173 (N_4173,N_3077,N_3770);
and U4174 (N_4174,N_3638,N_3977);
and U4175 (N_4175,N_3546,N_3248);
xnor U4176 (N_4176,N_3043,N_3838);
xor U4177 (N_4177,N_3709,N_3078);
nand U4178 (N_4178,N_3281,N_3503);
nand U4179 (N_4179,N_3338,N_3356);
or U4180 (N_4180,N_3535,N_3664);
xnor U4181 (N_4181,N_3605,N_3839);
xor U4182 (N_4182,N_3378,N_3788);
nand U4183 (N_4183,N_3793,N_3037);
and U4184 (N_4184,N_3297,N_3571);
or U4185 (N_4185,N_3012,N_3398);
nand U4186 (N_4186,N_3648,N_3273);
or U4187 (N_4187,N_3772,N_3521);
nand U4188 (N_4188,N_3707,N_3144);
nand U4189 (N_4189,N_3508,N_3654);
xnor U4190 (N_4190,N_3514,N_3915);
or U4191 (N_4191,N_3084,N_3659);
xor U4192 (N_4192,N_3257,N_3821);
and U4193 (N_4193,N_3903,N_3479);
xor U4194 (N_4194,N_3717,N_3208);
or U4195 (N_4195,N_3325,N_3894);
nand U4196 (N_4196,N_3455,N_3517);
xnor U4197 (N_4197,N_3624,N_3359);
nand U4198 (N_4198,N_3259,N_3827);
xnor U4199 (N_4199,N_3411,N_3413);
nand U4200 (N_4200,N_3602,N_3682);
xor U4201 (N_4201,N_3752,N_3757);
nor U4202 (N_4202,N_3083,N_3374);
nor U4203 (N_4203,N_3761,N_3981);
xor U4204 (N_4204,N_3528,N_3512);
or U4205 (N_4205,N_3067,N_3906);
and U4206 (N_4206,N_3728,N_3778);
nand U4207 (N_4207,N_3653,N_3351);
nand U4208 (N_4208,N_3558,N_3544);
nand U4209 (N_4209,N_3585,N_3650);
or U4210 (N_4210,N_3090,N_3428);
and U4211 (N_4211,N_3015,N_3168);
nand U4212 (N_4212,N_3337,N_3448);
nor U4213 (N_4213,N_3863,N_3766);
xnor U4214 (N_4214,N_3282,N_3303);
nor U4215 (N_4215,N_3157,N_3815);
nor U4216 (N_4216,N_3335,N_3461);
nand U4217 (N_4217,N_3532,N_3426);
nand U4218 (N_4218,N_3327,N_3127);
nor U4219 (N_4219,N_3978,N_3776);
and U4220 (N_4220,N_3673,N_3562);
and U4221 (N_4221,N_3097,N_3649);
xnor U4222 (N_4222,N_3810,N_3860);
xnor U4223 (N_4223,N_3110,N_3896);
nor U4224 (N_4224,N_3193,N_3480);
nor U4225 (N_4225,N_3258,N_3706);
or U4226 (N_4226,N_3868,N_3566);
and U4227 (N_4227,N_3118,N_3804);
and U4228 (N_4228,N_3536,N_3964);
or U4229 (N_4229,N_3249,N_3754);
nor U4230 (N_4230,N_3872,N_3495);
nor U4231 (N_4231,N_3856,N_3214);
nor U4232 (N_4232,N_3642,N_3264);
nor U4233 (N_4233,N_3916,N_3555);
nand U4234 (N_4234,N_3005,N_3290);
nand U4235 (N_4235,N_3666,N_3755);
or U4236 (N_4236,N_3462,N_3373);
nand U4237 (N_4237,N_3575,N_3291);
or U4238 (N_4238,N_3304,N_3843);
and U4239 (N_4239,N_3035,N_3365);
xor U4240 (N_4240,N_3513,N_3840);
and U4241 (N_4241,N_3569,N_3515);
xnor U4242 (N_4242,N_3262,N_3869);
nand U4243 (N_4243,N_3845,N_3104);
nor U4244 (N_4244,N_3841,N_3419);
and U4245 (N_4245,N_3484,N_3085);
nand U4246 (N_4246,N_3579,N_3404);
or U4247 (N_4247,N_3871,N_3403);
and U4248 (N_4248,N_3997,N_3469);
xnor U4249 (N_4249,N_3474,N_3414);
or U4250 (N_4250,N_3542,N_3138);
and U4251 (N_4251,N_3511,N_3092);
nor U4252 (N_4252,N_3646,N_3001);
nor U4253 (N_4253,N_3959,N_3668);
and U4254 (N_4254,N_3283,N_3478);
or U4255 (N_4255,N_3763,N_3368);
nor U4256 (N_4256,N_3186,N_3209);
xor U4257 (N_4257,N_3637,N_3623);
nand U4258 (N_4258,N_3941,N_3736);
and U4259 (N_4259,N_3929,N_3055);
and U4260 (N_4260,N_3537,N_3958);
nor U4261 (N_4261,N_3238,N_3783);
and U4262 (N_4262,N_3655,N_3583);
or U4263 (N_4263,N_3178,N_3472);
nand U4264 (N_4264,N_3530,N_3593);
and U4265 (N_4265,N_3608,N_3370);
nand U4266 (N_4266,N_3352,N_3276);
nand U4267 (N_4267,N_3441,N_3912);
or U4268 (N_4268,N_3940,N_3269);
and U4269 (N_4269,N_3140,N_3982);
xor U4270 (N_4270,N_3375,N_3917);
and U4271 (N_4271,N_3606,N_3700);
and U4272 (N_4272,N_3961,N_3393);
nand U4273 (N_4273,N_3600,N_3910);
nand U4274 (N_4274,N_3254,N_3156);
nor U4275 (N_4275,N_3086,N_3563);
or U4276 (N_4276,N_3384,N_3032);
or U4277 (N_4277,N_3587,N_3314);
xnor U4278 (N_4278,N_3765,N_3155);
and U4279 (N_4279,N_3452,N_3956);
nor U4280 (N_4280,N_3496,N_3380);
nor U4281 (N_4281,N_3355,N_3826);
and U4282 (N_4282,N_3025,N_3632);
nor U4283 (N_4283,N_3732,N_3572);
xor U4284 (N_4284,N_3089,N_3131);
nand U4285 (N_4285,N_3236,N_3132);
nor U4286 (N_4286,N_3333,N_3825);
nand U4287 (N_4287,N_3036,N_3301);
and U4288 (N_4288,N_3423,N_3346);
xor U4289 (N_4289,N_3937,N_3427);
nand U4290 (N_4290,N_3658,N_3087);
nor U4291 (N_4291,N_3560,N_3239);
and U4292 (N_4292,N_3900,N_3762);
xor U4293 (N_4293,N_3486,N_3453);
and U4294 (N_4294,N_3519,N_3027);
nor U4295 (N_4295,N_3852,N_3609);
or U4296 (N_4296,N_3570,N_3471);
xnor U4297 (N_4297,N_3897,N_3240);
nand U4298 (N_4298,N_3218,N_3726);
nor U4299 (N_4299,N_3071,N_3848);
xor U4300 (N_4300,N_3383,N_3740);
xnor U4301 (N_4301,N_3360,N_3619);
xor U4302 (N_4302,N_3099,N_3865);
nor U4303 (N_4303,N_3799,N_3858);
nand U4304 (N_4304,N_3111,N_3702);
xor U4305 (N_4305,N_3255,N_3116);
and U4306 (N_4306,N_3818,N_3341);
nand U4307 (N_4307,N_3954,N_3215);
xor U4308 (N_4308,N_3594,N_3960);
nor U4309 (N_4309,N_3953,N_3285);
nand U4310 (N_4310,N_3980,N_3447);
and U4311 (N_4311,N_3422,N_3235);
and U4312 (N_4312,N_3800,N_3034);
and U4313 (N_4313,N_3271,N_3934);
nand U4314 (N_4314,N_3041,N_3151);
nor U4315 (N_4315,N_3808,N_3907);
and U4316 (N_4316,N_3507,N_3261);
nand U4317 (N_4317,N_3159,N_3698);
xnor U4318 (N_4318,N_3446,N_3689);
and U4319 (N_4319,N_3207,N_3294);
and U4320 (N_4320,N_3203,N_3948);
or U4321 (N_4321,N_3785,N_3782);
nor U4322 (N_4322,N_3984,N_3057);
xor U4323 (N_4323,N_3316,N_3727);
and U4324 (N_4324,N_3498,N_3056);
nor U4325 (N_4325,N_3066,N_3139);
and U4326 (N_4326,N_3483,N_3120);
nor U4327 (N_4327,N_3306,N_3641);
nand U4328 (N_4328,N_3397,N_3122);
and U4329 (N_4329,N_3477,N_3194);
xnor U4330 (N_4330,N_3109,N_3366);
or U4331 (N_4331,N_3268,N_3919);
nor U4332 (N_4332,N_3518,N_3074);
nor U4333 (N_4333,N_3054,N_3379);
and U4334 (N_4334,N_3191,N_3494);
nand U4335 (N_4335,N_3887,N_3320);
nand U4336 (N_4336,N_3541,N_3182);
nand U4337 (N_4337,N_3394,N_3943);
or U4338 (N_4338,N_3434,N_3321);
xnor U4339 (N_4339,N_3197,N_3975);
xor U4340 (N_4340,N_3950,N_3362);
and U4341 (N_4341,N_3962,N_3992);
or U4342 (N_4342,N_3105,N_3344);
nand U4343 (N_4343,N_3121,N_3881);
or U4344 (N_4344,N_3421,N_3252);
nand U4345 (N_4345,N_3928,N_3098);
and U4346 (N_4346,N_3371,N_3874);
nor U4347 (N_4347,N_3993,N_3266);
or U4348 (N_4348,N_3590,N_3210);
or U4349 (N_4349,N_3988,N_3003);
or U4350 (N_4350,N_3837,N_3142);
xor U4351 (N_4351,N_3224,N_3633);
or U4352 (N_4352,N_3040,N_3749);
xnor U4353 (N_4353,N_3296,N_3846);
nand U4354 (N_4354,N_3760,N_3154);
or U4355 (N_4355,N_3998,N_3308);
xnor U4356 (N_4356,N_3879,N_3107);
nor U4357 (N_4357,N_3729,N_3720);
or U4358 (N_4358,N_3234,N_3408);
nand U4359 (N_4359,N_3245,N_3389);
and U4360 (N_4360,N_3708,N_3714);
nand U4361 (N_4361,N_3979,N_3816);
or U4362 (N_4362,N_3243,N_3510);
nand U4363 (N_4363,N_3522,N_3334);
and U4364 (N_4364,N_3242,N_3286);
nand U4365 (N_4365,N_3774,N_3777);
nor U4366 (N_4366,N_3946,N_3949);
nand U4367 (N_4367,N_3644,N_3029);
nand U4368 (N_4368,N_3677,N_3527);
or U4369 (N_4369,N_3904,N_3913);
nand U4370 (N_4370,N_3775,N_3927);
nor U4371 (N_4371,N_3161,N_3364);
or U4372 (N_4372,N_3204,N_3222);
nor U4373 (N_4373,N_3196,N_3690);
nand U4374 (N_4374,N_3392,N_3030);
xnor U4375 (N_4375,N_3185,N_3719);
xnor U4376 (N_4376,N_3739,N_3968);
and U4377 (N_4377,N_3909,N_3363);
xnor U4378 (N_4378,N_3028,N_3712);
and U4379 (N_4379,N_3891,N_3202);
nand U4380 (N_4380,N_3543,N_3628);
nor U4381 (N_4381,N_3621,N_3768);
nor U4382 (N_4382,N_3206,N_3126);
and U4383 (N_4383,N_3420,N_3795);
or U4384 (N_4384,N_3692,N_3319);
xor U4385 (N_4385,N_3061,N_3485);
xnor U4386 (N_4386,N_3930,N_3867);
and U4387 (N_4387,N_3323,N_3936);
or U4388 (N_4388,N_3093,N_3318);
and U4389 (N_4389,N_3735,N_3051);
and U4390 (N_4390,N_3023,N_3130);
xor U4391 (N_4391,N_3549,N_3859);
xnor U4392 (N_4392,N_3751,N_3289);
and U4393 (N_4393,N_3802,N_3790);
nor U4394 (N_4394,N_3625,N_3134);
or U4395 (N_4395,N_3769,N_3367);
or U4396 (N_4396,N_3232,N_3022);
xor U4397 (N_4397,N_3353,N_3226);
or U4398 (N_4398,N_3063,N_3295);
nand U4399 (N_4399,N_3683,N_3406);
nand U4400 (N_4400,N_3756,N_3277);
or U4401 (N_4401,N_3169,N_3592);
or U4402 (N_4402,N_3463,N_3180);
nor U4403 (N_4403,N_3416,N_3108);
and U4404 (N_4404,N_3786,N_3548);
nand U4405 (N_4405,N_3059,N_3877);
nand U4406 (N_4406,N_3481,N_3307);
nor U4407 (N_4407,N_3052,N_3343);
xnor U4408 (N_4408,N_3612,N_3009);
nor U4409 (N_4409,N_3179,N_3275);
and U4410 (N_4410,N_3409,N_3938);
or U4411 (N_4411,N_3450,N_3746);
xnor U4412 (N_4412,N_3339,N_3806);
xor U4413 (N_4413,N_3128,N_3038);
and U4414 (N_4414,N_3847,N_3699);
xnor U4415 (N_4415,N_3072,N_3640);
nand U4416 (N_4416,N_3759,N_3482);
and U4417 (N_4417,N_3165,N_3189);
and U4418 (N_4418,N_3773,N_3017);
xor U4419 (N_4419,N_3691,N_3136);
xor U4420 (N_4420,N_3457,N_3167);
nand U4421 (N_4421,N_3502,N_3743);
nand U4422 (N_4422,N_3467,N_3278);
and U4423 (N_4423,N_3187,N_3889);
nand U4424 (N_4424,N_3018,N_3618);
nor U4425 (N_4425,N_3260,N_3146);
xnor U4426 (N_4426,N_3190,N_3622);
nor U4427 (N_4427,N_3792,N_3440);
nand U4428 (N_4428,N_3805,N_3317);
nor U4429 (N_4429,N_3177,N_3133);
or U4430 (N_4430,N_3864,N_3703);
and U4431 (N_4431,N_3733,N_3713);
nand U4432 (N_4432,N_3985,N_3933);
or U4433 (N_4433,N_3737,N_3526);
xnor U4434 (N_4434,N_3595,N_3199);
or U4435 (N_4435,N_3044,N_3287);
nor U4436 (N_4436,N_3695,N_3935);
nor U4437 (N_4437,N_3162,N_3381);
or U4438 (N_4438,N_3464,N_3438);
nand U4439 (N_4439,N_3410,N_3591);
nand U4440 (N_4440,N_3068,N_3878);
or U4441 (N_4441,N_3991,N_3557);
or U4442 (N_4442,N_3741,N_3813);
and U4443 (N_4443,N_3932,N_3312);
nor U4444 (N_4444,N_3586,N_3458);
nand U4445 (N_4445,N_3117,N_3497);
xor U4446 (N_4446,N_3021,N_3688);
nor U4447 (N_4447,N_3158,N_3556);
xor U4448 (N_4448,N_3635,N_3100);
nand U4449 (N_4449,N_3137,N_3970);
or U4450 (N_4450,N_3152,N_3219);
xor U4451 (N_4451,N_3947,N_3844);
nand U4452 (N_4452,N_3581,N_3330);
nand U4453 (N_4453,N_3939,N_3967);
and U4454 (N_4454,N_3006,N_3730);
nand U4455 (N_4455,N_3401,N_3048);
xor U4456 (N_4456,N_3599,N_3745);
and U4457 (N_4457,N_3951,N_3164);
xor U4458 (N_4458,N_3657,N_3200);
nand U4459 (N_4459,N_3718,N_3895);
xor U4460 (N_4460,N_3449,N_3007);
and U4461 (N_4461,N_3228,N_3227);
xor U4462 (N_4462,N_3004,N_3516);
and U4463 (N_4463,N_3670,N_3509);
nor U4464 (N_4464,N_3220,N_3764);
xnor U4465 (N_4465,N_3823,N_3331);
nand U4466 (N_4466,N_3505,N_3431);
or U4467 (N_4467,N_3476,N_3225);
or U4468 (N_4468,N_3824,N_3880);
xor U4469 (N_4469,N_3429,N_3771);
or U4470 (N_4470,N_3862,N_3229);
nor U4471 (N_4471,N_3611,N_3661);
and U4472 (N_4472,N_3812,N_3103);
or U4473 (N_4473,N_3614,N_3669);
nand U4474 (N_4474,N_3415,N_3565);
nand U4475 (N_4475,N_3849,N_3173);
and U4476 (N_4476,N_3272,N_3551);
and U4477 (N_4477,N_3665,N_3647);
or U4478 (N_4478,N_3008,N_3905);
or U4479 (N_4479,N_3388,N_3576);
nor U4480 (N_4480,N_3309,N_3115);
or U4481 (N_4481,N_3842,N_3060);
nor U4482 (N_4482,N_3302,N_3183);
and U4483 (N_4483,N_3466,N_3198);
nand U4484 (N_4484,N_3385,N_3972);
nor U4485 (N_4485,N_3233,N_3195);
xnor U4486 (N_4486,N_3026,N_3443);
nor U4487 (N_4487,N_3372,N_3050);
nor U4488 (N_4488,N_3357,N_3884);
xor U4489 (N_4489,N_3047,N_3921);
nand U4490 (N_4490,N_3315,N_3995);
xor U4491 (N_4491,N_3791,N_3114);
nor U4492 (N_4492,N_3329,N_3211);
and U4493 (N_4493,N_3418,N_3534);
nand U4494 (N_4494,N_3487,N_3081);
nor U4495 (N_4495,N_3492,N_3096);
nand U4496 (N_4496,N_3681,N_3987);
nor U4497 (N_4497,N_3854,N_3767);
xnor U4498 (N_4498,N_3376,N_3020);
nor U4499 (N_4499,N_3279,N_3701);
xnor U4500 (N_4500,N_3475,N_3195);
xnor U4501 (N_4501,N_3662,N_3739);
nand U4502 (N_4502,N_3098,N_3438);
and U4503 (N_4503,N_3921,N_3196);
or U4504 (N_4504,N_3663,N_3128);
nor U4505 (N_4505,N_3562,N_3001);
nand U4506 (N_4506,N_3314,N_3464);
nand U4507 (N_4507,N_3539,N_3054);
xnor U4508 (N_4508,N_3484,N_3975);
nor U4509 (N_4509,N_3665,N_3007);
nand U4510 (N_4510,N_3179,N_3943);
and U4511 (N_4511,N_3158,N_3922);
and U4512 (N_4512,N_3943,N_3830);
nor U4513 (N_4513,N_3683,N_3916);
xnor U4514 (N_4514,N_3892,N_3719);
nor U4515 (N_4515,N_3137,N_3941);
or U4516 (N_4516,N_3432,N_3633);
or U4517 (N_4517,N_3761,N_3618);
and U4518 (N_4518,N_3492,N_3904);
xor U4519 (N_4519,N_3794,N_3621);
or U4520 (N_4520,N_3796,N_3313);
xnor U4521 (N_4521,N_3276,N_3295);
nand U4522 (N_4522,N_3187,N_3219);
nor U4523 (N_4523,N_3875,N_3131);
nand U4524 (N_4524,N_3148,N_3879);
nand U4525 (N_4525,N_3237,N_3966);
or U4526 (N_4526,N_3232,N_3237);
nand U4527 (N_4527,N_3474,N_3444);
nor U4528 (N_4528,N_3713,N_3460);
xor U4529 (N_4529,N_3820,N_3766);
or U4530 (N_4530,N_3564,N_3868);
and U4531 (N_4531,N_3930,N_3929);
nand U4532 (N_4532,N_3457,N_3220);
xnor U4533 (N_4533,N_3536,N_3338);
or U4534 (N_4534,N_3577,N_3278);
nor U4535 (N_4535,N_3265,N_3866);
nor U4536 (N_4536,N_3502,N_3080);
nand U4537 (N_4537,N_3399,N_3955);
or U4538 (N_4538,N_3693,N_3150);
nand U4539 (N_4539,N_3516,N_3304);
xor U4540 (N_4540,N_3119,N_3134);
or U4541 (N_4541,N_3340,N_3533);
xor U4542 (N_4542,N_3458,N_3456);
nand U4543 (N_4543,N_3589,N_3009);
and U4544 (N_4544,N_3251,N_3053);
nor U4545 (N_4545,N_3631,N_3231);
nor U4546 (N_4546,N_3854,N_3415);
nor U4547 (N_4547,N_3077,N_3886);
nor U4548 (N_4548,N_3499,N_3420);
xnor U4549 (N_4549,N_3158,N_3776);
xor U4550 (N_4550,N_3659,N_3316);
nand U4551 (N_4551,N_3239,N_3162);
nor U4552 (N_4552,N_3489,N_3578);
nor U4553 (N_4553,N_3276,N_3470);
nor U4554 (N_4554,N_3051,N_3688);
or U4555 (N_4555,N_3457,N_3137);
xnor U4556 (N_4556,N_3899,N_3850);
and U4557 (N_4557,N_3326,N_3125);
nor U4558 (N_4558,N_3225,N_3506);
and U4559 (N_4559,N_3851,N_3602);
or U4560 (N_4560,N_3197,N_3239);
or U4561 (N_4561,N_3348,N_3657);
nor U4562 (N_4562,N_3077,N_3490);
nand U4563 (N_4563,N_3114,N_3377);
or U4564 (N_4564,N_3045,N_3889);
or U4565 (N_4565,N_3478,N_3398);
or U4566 (N_4566,N_3959,N_3680);
or U4567 (N_4567,N_3148,N_3254);
nor U4568 (N_4568,N_3036,N_3440);
nand U4569 (N_4569,N_3557,N_3967);
nor U4570 (N_4570,N_3396,N_3604);
nor U4571 (N_4571,N_3209,N_3749);
or U4572 (N_4572,N_3872,N_3224);
or U4573 (N_4573,N_3588,N_3048);
and U4574 (N_4574,N_3189,N_3898);
nor U4575 (N_4575,N_3915,N_3893);
and U4576 (N_4576,N_3724,N_3857);
nor U4577 (N_4577,N_3450,N_3669);
nand U4578 (N_4578,N_3821,N_3355);
or U4579 (N_4579,N_3857,N_3166);
nand U4580 (N_4580,N_3723,N_3749);
or U4581 (N_4581,N_3277,N_3465);
xnor U4582 (N_4582,N_3151,N_3822);
or U4583 (N_4583,N_3636,N_3449);
or U4584 (N_4584,N_3070,N_3306);
nand U4585 (N_4585,N_3758,N_3202);
nand U4586 (N_4586,N_3454,N_3978);
nor U4587 (N_4587,N_3238,N_3002);
or U4588 (N_4588,N_3278,N_3625);
and U4589 (N_4589,N_3320,N_3118);
nand U4590 (N_4590,N_3221,N_3585);
or U4591 (N_4591,N_3897,N_3086);
nor U4592 (N_4592,N_3444,N_3302);
and U4593 (N_4593,N_3513,N_3306);
and U4594 (N_4594,N_3792,N_3057);
nand U4595 (N_4595,N_3836,N_3013);
xnor U4596 (N_4596,N_3162,N_3573);
nand U4597 (N_4597,N_3075,N_3969);
xor U4598 (N_4598,N_3190,N_3848);
or U4599 (N_4599,N_3655,N_3664);
nand U4600 (N_4600,N_3496,N_3560);
xnor U4601 (N_4601,N_3557,N_3834);
or U4602 (N_4602,N_3407,N_3467);
nor U4603 (N_4603,N_3883,N_3122);
xnor U4604 (N_4604,N_3043,N_3634);
xnor U4605 (N_4605,N_3505,N_3131);
nand U4606 (N_4606,N_3660,N_3257);
nor U4607 (N_4607,N_3780,N_3642);
nor U4608 (N_4608,N_3350,N_3693);
and U4609 (N_4609,N_3600,N_3066);
or U4610 (N_4610,N_3564,N_3297);
xnor U4611 (N_4611,N_3082,N_3615);
or U4612 (N_4612,N_3685,N_3143);
and U4613 (N_4613,N_3928,N_3560);
or U4614 (N_4614,N_3268,N_3988);
or U4615 (N_4615,N_3998,N_3676);
nor U4616 (N_4616,N_3125,N_3691);
and U4617 (N_4617,N_3334,N_3616);
nor U4618 (N_4618,N_3209,N_3666);
or U4619 (N_4619,N_3935,N_3093);
and U4620 (N_4620,N_3093,N_3374);
nand U4621 (N_4621,N_3188,N_3089);
and U4622 (N_4622,N_3579,N_3725);
or U4623 (N_4623,N_3936,N_3162);
nand U4624 (N_4624,N_3077,N_3357);
nand U4625 (N_4625,N_3942,N_3994);
or U4626 (N_4626,N_3825,N_3628);
xor U4627 (N_4627,N_3916,N_3273);
xor U4628 (N_4628,N_3402,N_3611);
or U4629 (N_4629,N_3045,N_3136);
and U4630 (N_4630,N_3612,N_3957);
or U4631 (N_4631,N_3828,N_3207);
or U4632 (N_4632,N_3470,N_3567);
nand U4633 (N_4633,N_3430,N_3928);
or U4634 (N_4634,N_3528,N_3025);
or U4635 (N_4635,N_3235,N_3433);
or U4636 (N_4636,N_3141,N_3012);
nor U4637 (N_4637,N_3267,N_3254);
nand U4638 (N_4638,N_3430,N_3124);
and U4639 (N_4639,N_3464,N_3061);
xor U4640 (N_4640,N_3191,N_3333);
nor U4641 (N_4641,N_3430,N_3337);
nor U4642 (N_4642,N_3546,N_3485);
nor U4643 (N_4643,N_3964,N_3324);
and U4644 (N_4644,N_3501,N_3149);
and U4645 (N_4645,N_3731,N_3519);
or U4646 (N_4646,N_3990,N_3629);
and U4647 (N_4647,N_3381,N_3031);
nor U4648 (N_4648,N_3998,N_3184);
nor U4649 (N_4649,N_3013,N_3290);
xor U4650 (N_4650,N_3982,N_3337);
or U4651 (N_4651,N_3290,N_3289);
nand U4652 (N_4652,N_3536,N_3424);
nor U4653 (N_4653,N_3037,N_3103);
and U4654 (N_4654,N_3621,N_3579);
or U4655 (N_4655,N_3476,N_3131);
nor U4656 (N_4656,N_3507,N_3407);
nor U4657 (N_4657,N_3255,N_3108);
xnor U4658 (N_4658,N_3373,N_3766);
or U4659 (N_4659,N_3638,N_3958);
and U4660 (N_4660,N_3173,N_3031);
nand U4661 (N_4661,N_3157,N_3576);
nand U4662 (N_4662,N_3622,N_3482);
or U4663 (N_4663,N_3402,N_3079);
or U4664 (N_4664,N_3702,N_3131);
xnor U4665 (N_4665,N_3968,N_3716);
and U4666 (N_4666,N_3418,N_3412);
or U4667 (N_4667,N_3744,N_3383);
or U4668 (N_4668,N_3226,N_3765);
xor U4669 (N_4669,N_3227,N_3987);
nor U4670 (N_4670,N_3161,N_3344);
or U4671 (N_4671,N_3541,N_3872);
and U4672 (N_4672,N_3010,N_3394);
xnor U4673 (N_4673,N_3708,N_3105);
and U4674 (N_4674,N_3127,N_3027);
nand U4675 (N_4675,N_3253,N_3576);
nor U4676 (N_4676,N_3880,N_3227);
and U4677 (N_4677,N_3019,N_3469);
or U4678 (N_4678,N_3462,N_3547);
xor U4679 (N_4679,N_3833,N_3519);
or U4680 (N_4680,N_3624,N_3357);
nand U4681 (N_4681,N_3265,N_3130);
xnor U4682 (N_4682,N_3296,N_3318);
nor U4683 (N_4683,N_3161,N_3004);
and U4684 (N_4684,N_3545,N_3484);
xnor U4685 (N_4685,N_3932,N_3885);
nand U4686 (N_4686,N_3133,N_3501);
or U4687 (N_4687,N_3580,N_3013);
or U4688 (N_4688,N_3032,N_3962);
xor U4689 (N_4689,N_3411,N_3375);
nand U4690 (N_4690,N_3696,N_3594);
or U4691 (N_4691,N_3442,N_3954);
nand U4692 (N_4692,N_3272,N_3503);
or U4693 (N_4693,N_3160,N_3582);
nor U4694 (N_4694,N_3554,N_3589);
nor U4695 (N_4695,N_3630,N_3667);
and U4696 (N_4696,N_3505,N_3404);
nor U4697 (N_4697,N_3644,N_3992);
nor U4698 (N_4698,N_3752,N_3906);
and U4699 (N_4699,N_3204,N_3918);
nor U4700 (N_4700,N_3975,N_3148);
xor U4701 (N_4701,N_3430,N_3644);
or U4702 (N_4702,N_3555,N_3056);
and U4703 (N_4703,N_3898,N_3344);
nor U4704 (N_4704,N_3248,N_3990);
and U4705 (N_4705,N_3982,N_3935);
or U4706 (N_4706,N_3017,N_3858);
nand U4707 (N_4707,N_3351,N_3798);
xor U4708 (N_4708,N_3097,N_3572);
xnor U4709 (N_4709,N_3324,N_3894);
nand U4710 (N_4710,N_3487,N_3636);
nand U4711 (N_4711,N_3689,N_3667);
xor U4712 (N_4712,N_3706,N_3107);
and U4713 (N_4713,N_3675,N_3659);
nand U4714 (N_4714,N_3455,N_3385);
nor U4715 (N_4715,N_3132,N_3563);
or U4716 (N_4716,N_3507,N_3276);
and U4717 (N_4717,N_3076,N_3875);
xnor U4718 (N_4718,N_3360,N_3705);
and U4719 (N_4719,N_3118,N_3075);
or U4720 (N_4720,N_3369,N_3415);
and U4721 (N_4721,N_3894,N_3009);
nor U4722 (N_4722,N_3622,N_3911);
xnor U4723 (N_4723,N_3106,N_3165);
or U4724 (N_4724,N_3973,N_3185);
xor U4725 (N_4725,N_3882,N_3760);
and U4726 (N_4726,N_3893,N_3788);
or U4727 (N_4727,N_3325,N_3626);
xnor U4728 (N_4728,N_3546,N_3413);
nand U4729 (N_4729,N_3871,N_3414);
xnor U4730 (N_4730,N_3395,N_3332);
or U4731 (N_4731,N_3989,N_3893);
nand U4732 (N_4732,N_3617,N_3908);
and U4733 (N_4733,N_3396,N_3330);
nor U4734 (N_4734,N_3558,N_3534);
nor U4735 (N_4735,N_3732,N_3382);
nor U4736 (N_4736,N_3679,N_3996);
nor U4737 (N_4737,N_3267,N_3624);
nor U4738 (N_4738,N_3573,N_3694);
nor U4739 (N_4739,N_3751,N_3852);
or U4740 (N_4740,N_3296,N_3015);
or U4741 (N_4741,N_3560,N_3743);
nor U4742 (N_4742,N_3341,N_3709);
nor U4743 (N_4743,N_3073,N_3621);
and U4744 (N_4744,N_3671,N_3447);
and U4745 (N_4745,N_3764,N_3842);
xnor U4746 (N_4746,N_3500,N_3245);
xor U4747 (N_4747,N_3317,N_3343);
nand U4748 (N_4748,N_3040,N_3912);
xor U4749 (N_4749,N_3020,N_3962);
nor U4750 (N_4750,N_3284,N_3832);
xnor U4751 (N_4751,N_3093,N_3412);
xnor U4752 (N_4752,N_3165,N_3003);
xor U4753 (N_4753,N_3942,N_3618);
xnor U4754 (N_4754,N_3010,N_3736);
and U4755 (N_4755,N_3602,N_3873);
or U4756 (N_4756,N_3744,N_3096);
or U4757 (N_4757,N_3487,N_3438);
xor U4758 (N_4758,N_3182,N_3342);
and U4759 (N_4759,N_3667,N_3733);
or U4760 (N_4760,N_3670,N_3629);
xor U4761 (N_4761,N_3811,N_3258);
nor U4762 (N_4762,N_3528,N_3506);
and U4763 (N_4763,N_3979,N_3308);
xor U4764 (N_4764,N_3398,N_3511);
nor U4765 (N_4765,N_3785,N_3425);
nand U4766 (N_4766,N_3783,N_3618);
nand U4767 (N_4767,N_3570,N_3775);
xnor U4768 (N_4768,N_3857,N_3438);
or U4769 (N_4769,N_3311,N_3107);
nand U4770 (N_4770,N_3717,N_3078);
nand U4771 (N_4771,N_3145,N_3809);
xor U4772 (N_4772,N_3471,N_3772);
and U4773 (N_4773,N_3603,N_3156);
nor U4774 (N_4774,N_3722,N_3463);
nand U4775 (N_4775,N_3675,N_3160);
xor U4776 (N_4776,N_3026,N_3411);
or U4777 (N_4777,N_3146,N_3979);
nand U4778 (N_4778,N_3743,N_3097);
and U4779 (N_4779,N_3406,N_3761);
and U4780 (N_4780,N_3301,N_3236);
nand U4781 (N_4781,N_3651,N_3110);
nor U4782 (N_4782,N_3717,N_3061);
or U4783 (N_4783,N_3006,N_3418);
or U4784 (N_4784,N_3166,N_3879);
xnor U4785 (N_4785,N_3861,N_3277);
and U4786 (N_4786,N_3174,N_3834);
and U4787 (N_4787,N_3331,N_3008);
or U4788 (N_4788,N_3672,N_3406);
xnor U4789 (N_4789,N_3673,N_3074);
and U4790 (N_4790,N_3096,N_3882);
nand U4791 (N_4791,N_3405,N_3144);
nand U4792 (N_4792,N_3077,N_3106);
or U4793 (N_4793,N_3572,N_3896);
and U4794 (N_4794,N_3719,N_3684);
nor U4795 (N_4795,N_3863,N_3075);
xor U4796 (N_4796,N_3330,N_3225);
nor U4797 (N_4797,N_3964,N_3957);
xnor U4798 (N_4798,N_3683,N_3115);
or U4799 (N_4799,N_3498,N_3273);
nor U4800 (N_4800,N_3923,N_3382);
xnor U4801 (N_4801,N_3588,N_3445);
nand U4802 (N_4802,N_3904,N_3366);
nor U4803 (N_4803,N_3918,N_3850);
nor U4804 (N_4804,N_3553,N_3895);
nand U4805 (N_4805,N_3272,N_3813);
or U4806 (N_4806,N_3342,N_3188);
xnor U4807 (N_4807,N_3800,N_3138);
xor U4808 (N_4808,N_3540,N_3392);
xor U4809 (N_4809,N_3153,N_3613);
xnor U4810 (N_4810,N_3538,N_3498);
xor U4811 (N_4811,N_3454,N_3551);
xnor U4812 (N_4812,N_3621,N_3510);
nand U4813 (N_4813,N_3426,N_3730);
or U4814 (N_4814,N_3658,N_3382);
and U4815 (N_4815,N_3163,N_3086);
xor U4816 (N_4816,N_3125,N_3527);
nor U4817 (N_4817,N_3683,N_3978);
nand U4818 (N_4818,N_3981,N_3059);
nand U4819 (N_4819,N_3095,N_3337);
and U4820 (N_4820,N_3124,N_3546);
nor U4821 (N_4821,N_3411,N_3157);
and U4822 (N_4822,N_3435,N_3692);
nand U4823 (N_4823,N_3067,N_3853);
nand U4824 (N_4824,N_3118,N_3605);
or U4825 (N_4825,N_3996,N_3202);
xor U4826 (N_4826,N_3857,N_3412);
or U4827 (N_4827,N_3057,N_3771);
nand U4828 (N_4828,N_3672,N_3011);
nand U4829 (N_4829,N_3992,N_3090);
nor U4830 (N_4830,N_3024,N_3152);
nor U4831 (N_4831,N_3807,N_3185);
or U4832 (N_4832,N_3615,N_3217);
xor U4833 (N_4833,N_3670,N_3838);
and U4834 (N_4834,N_3078,N_3872);
nand U4835 (N_4835,N_3951,N_3107);
and U4836 (N_4836,N_3822,N_3414);
nand U4837 (N_4837,N_3562,N_3353);
and U4838 (N_4838,N_3683,N_3464);
nor U4839 (N_4839,N_3713,N_3559);
xor U4840 (N_4840,N_3973,N_3139);
nor U4841 (N_4841,N_3318,N_3446);
nand U4842 (N_4842,N_3082,N_3980);
nor U4843 (N_4843,N_3798,N_3623);
nor U4844 (N_4844,N_3606,N_3899);
nand U4845 (N_4845,N_3360,N_3048);
nor U4846 (N_4846,N_3152,N_3331);
and U4847 (N_4847,N_3436,N_3461);
nand U4848 (N_4848,N_3379,N_3028);
and U4849 (N_4849,N_3701,N_3419);
and U4850 (N_4850,N_3669,N_3618);
nand U4851 (N_4851,N_3773,N_3688);
and U4852 (N_4852,N_3817,N_3439);
or U4853 (N_4853,N_3304,N_3976);
and U4854 (N_4854,N_3094,N_3338);
xnor U4855 (N_4855,N_3254,N_3166);
and U4856 (N_4856,N_3606,N_3761);
and U4857 (N_4857,N_3782,N_3096);
nand U4858 (N_4858,N_3024,N_3674);
and U4859 (N_4859,N_3986,N_3716);
nor U4860 (N_4860,N_3177,N_3490);
nor U4861 (N_4861,N_3833,N_3888);
or U4862 (N_4862,N_3305,N_3322);
nor U4863 (N_4863,N_3860,N_3836);
xor U4864 (N_4864,N_3719,N_3703);
or U4865 (N_4865,N_3760,N_3911);
nand U4866 (N_4866,N_3142,N_3757);
nor U4867 (N_4867,N_3217,N_3765);
nand U4868 (N_4868,N_3287,N_3155);
xnor U4869 (N_4869,N_3669,N_3506);
xnor U4870 (N_4870,N_3931,N_3590);
and U4871 (N_4871,N_3853,N_3464);
or U4872 (N_4872,N_3730,N_3181);
and U4873 (N_4873,N_3020,N_3428);
or U4874 (N_4874,N_3765,N_3112);
or U4875 (N_4875,N_3116,N_3873);
xnor U4876 (N_4876,N_3715,N_3679);
and U4877 (N_4877,N_3285,N_3775);
nor U4878 (N_4878,N_3049,N_3624);
and U4879 (N_4879,N_3470,N_3349);
or U4880 (N_4880,N_3836,N_3692);
xor U4881 (N_4881,N_3863,N_3073);
nor U4882 (N_4882,N_3057,N_3365);
nor U4883 (N_4883,N_3757,N_3196);
nor U4884 (N_4884,N_3615,N_3833);
or U4885 (N_4885,N_3529,N_3379);
nand U4886 (N_4886,N_3042,N_3974);
nand U4887 (N_4887,N_3214,N_3045);
nand U4888 (N_4888,N_3179,N_3280);
and U4889 (N_4889,N_3651,N_3729);
nand U4890 (N_4890,N_3508,N_3349);
nand U4891 (N_4891,N_3058,N_3696);
and U4892 (N_4892,N_3088,N_3078);
nor U4893 (N_4893,N_3572,N_3141);
xor U4894 (N_4894,N_3913,N_3407);
nand U4895 (N_4895,N_3535,N_3558);
or U4896 (N_4896,N_3260,N_3570);
nand U4897 (N_4897,N_3042,N_3004);
or U4898 (N_4898,N_3056,N_3340);
or U4899 (N_4899,N_3097,N_3436);
nor U4900 (N_4900,N_3840,N_3441);
nand U4901 (N_4901,N_3357,N_3003);
and U4902 (N_4902,N_3905,N_3112);
nor U4903 (N_4903,N_3383,N_3400);
xor U4904 (N_4904,N_3985,N_3795);
nor U4905 (N_4905,N_3260,N_3023);
nor U4906 (N_4906,N_3484,N_3381);
and U4907 (N_4907,N_3434,N_3408);
nor U4908 (N_4908,N_3918,N_3436);
xor U4909 (N_4909,N_3150,N_3482);
nor U4910 (N_4910,N_3253,N_3872);
and U4911 (N_4911,N_3253,N_3288);
or U4912 (N_4912,N_3601,N_3716);
xor U4913 (N_4913,N_3639,N_3699);
and U4914 (N_4914,N_3587,N_3442);
and U4915 (N_4915,N_3708,N_3867);
nand U4916 (N_4916,N_3855,N_3994);
nor U4917 (N_4917,N_3919,N_3620);
or U4918 (N_4918,N_3832,N_3443);
or U4919 (N_4919,N_3362,N_3253);
nor U4920 (N_4920,N_3281,N_3472);
and U4921 (N_4921,N_3917,N_3073);
nand U4922 (N_4922,N_3509,N_3320);
or U4923 (N_4923,N_3434,N_3922);
and U4924 (N_4924,N_3787,N_3326);
xnor U4925 (N_4925,N_3112,N_3662);
and U4926 (N_4926,N_3442,N_3605);
nor U4927 (N_4927,N_3757,N_3368);
nor U4928 (N_4928,N_3493,N_3412);
and U4929 (N_4929,N_3219,N_3345);
nand U4930 (N_4930,N_3311,N_3630);
and U4931 (N_4931,N_3396,N_3874);
or U4932 (N_4932,N_3218,N_3185);
or U4933 (N_4933,N_3531,N_3082);
nand U4934 (N_4934,N_3438,N_3596);
and U4935 (N_4935,N_3127,N_3392);
nor U4936 (N_4936,N_3118,N_3936);
nor U4937 (N_4937,N_3503,N_3596);
nand U4938 (N_4938,N_3945,N_3213);
nand U4939 (N_4939,N_3342,N_3471);
nor U4940 (N_4940,N_3443,N_3045);
and U4941 (N_4941,N_3802,N_3130);
nand U4942 (N_4942,N_3933,N_3249);
and U4943 (N_4943,N_3807,N_3552);
nor U4944 (N_4944,N_3259,N_3545);
or U4945 (N_4945,N_3089,N_3029);
xor U4946 (N_4946,N_3473,N_3679);
nand U4947 (N_4947,N_3053,N_3776);
nand U4948 (N_4948,N_3574,N_3154);
nand U4949 (N_4949,N_3057,N_3811);
or U4950 (N_4950,N_3608,N_3797);
xnor U4951 (N_4951,N_3345,N_3982);
nor U4952 (N_4952,N_3121,N_3985);
or U4953 (N_4953,N_3883,N_3072);
or U4954 (N_4954,N_3422,N_3610);
nand U4955 (N_4955,N_3587,N_3130);
or U4956 (N_4956,N_3691,N_3237);
xnor U4957 (N_4957,N_3558,N_3806);
and U4958 (N_4958,N_3881,N_3738);
or U4959 (N_4959,N_3554,N_3873);
or U4960 (N_4960,N_3247,N_3455);
or U4961 (N_4961,N_3284,N_3479);
xnor U4962 (N_4962,N_3734,N_3504);
nand U4963 (N_4963,N_3248,N_3867);
nand U4964 (N_4964,N_3196,N_3807);
nand U4965 (N_4965,N_3727,N_3884);
or U4966 (N_4966,N_3457,N_3112);
and U4967 (N_4967,N_3632,N_3657);
nor U4968 (N_4968,N_3856,N_3580);
nand U4969 (N_4969,N_3371,N_3211);
xnor U4970 (N_4970,N_3149,N_3440);
xnor U4971 (N_4971,N_3023,N_3728);
nor U4972 (N_4972,N_3423,N_3834);
or U4973 (N_4973,N_3834,N_3288);
and U4974 (N_4974,N_3548,N_3700);
xor U4975 (N_4975,N_3988,N_3555);
and U4976 (N_4976,N_3930,N_3998);
nand U4977 (N_4977,N_3643,N_3070);
xor U4978 (N_4978,N_3351,N_3145);
and U4979 (N_4979,N_3519,N_3588);
or U4980 (N_4980,N_3847,N_3143);
xnor U4981 (N_4981,N_3102,N_3677);
or U4982 (N_4982,N_3983,N_3058);
xnor U4983 (N_4983,N_3574,N_3364);
and U4984 (N_4984,N_3830,N_3884);
nor U4985 (N_4985,N_3688,N_3855);
nand U4986 (N_4986,N_3129,N_3715);
xor U4987 (N_4987,N_3982,N_3565);
and U4988 (N_4988,N_3788,N_3608);
nor U4989 (N_4989,N_3006,N_3545);
nor U4990 (N_4990,N_3539,N_3200);
or U4991 (N_4991,N_3658,N_3170);
nand U4992 (N_4992,N_3155,N_3575);
and U4993 (N_4993,N_3788,N_3249);
xnor U4994 (N_4994,N_3835,N_3489);
xor U4995 (N_4995,N_3379,N_3393);
xnor U4996 (N_4996,N_3257,N_3629);
and U4997 (N_4997,N_3367,N_3457);
and U4998 (N_4998,N_3066,N_3774);
nor U4999 (N_4999,N_3698,N_3213);
or U5000 (N_5000,N_4812,N_4533);
nor U5001 (N_5001,N_4587,N_4323);
or U5002 (N_5002,N_4976,N_4597);
nand U5003 (N_5003,N_4528,N_4128);
nand U5004 (N_5004,N_4398,N_4354);
nor U5005 (N_5005,N_4382,N_4129);
and U5006 (N_5006,N_4755,N_4737);
and U5007 (N_5007,N_4853,N_4068);
nor U5008 (N_5008,N_4941,N_4772);
nor U5009 (N_5009,N_4649,N_4286);
nor U5010 (N_5010,N_4685,N_4273);
xnor U5011 (N_5011,N_4485,N_4534);
or U5012 (N_5012,N_4960,N_4102);
nand U5013 (N_5013,N_4702,N_4059);
and U5014 (N_5014,N_4308,N_4002);
nand U5015 (N_5015,N_4787,N_4612);
and U5016 (N_5016,N_4590,N_4616);
xor U5017 (N_5017,N_4746,N_4611);
nor U5018 (N_5018,N_4520,N_4602);
nor U5019 (N_5019,N_4221,N_4939);
nor U5020 (N_5020,N_4120,N_4161);
or U5021 (N_5021,N_4364,N_4727);
xor U5022 (N_5022,N_4095,N_4598);
nand U5023 (N_5023,N_4441,N_4368);
and U5024 (N_5024,N_4314,N_4252);
and U5025 (N_5025,N_4337,N_4654);
and U5026 (N_5026,N_4034,N_4225);
nor U5027 (N_5027,N_4815,N_4464);
nand U5028 (N_5028,N_4497,N_4257);
xnor U5029 (N_5029,N_4246,N_4355);
or U5030 (N_5030,N_4300,N_4176);
or U5031 (N_5031,N_4463,N_4197);
nand U5032 (N_5032,N_4537,N_4844);
xor U5033 (N_5033,N_4829,N_4046);
and U5034 (N_5034,N_4047,N_4847);
or U5035 (N_5035,N_4322,N_4025);
or U5036 (N_5036,N_4559,N_4642);
and U5037 (N_5037,N_4747,N_4925);
nand U5038 (N_5038,N_4431,N_4868);
nor U5039 (N_5039,N_4798,N_4019);
xor U5040 (N_5040,N_4106,N_4779);
and U5041 (N_5041,N_4507,N_4065);
or U5042 (N_5042,N_4061,N_4662);
and U5043 (N_5043,N_4443,N_4233);
or U5044 (N_5044,N_4644,N_4571);
and U5045 (N_5045,N_4543,N_4473);
nand U5046 (N_5046,N_4499,N_4601);
or U5047 (N_5047,N_4591,N_4969);
nand U5048 (N_5048,N_4773,N_4149);
xor U5049 (N_5049,N_4152,N_4080);
and U5050 (N_5050,N_4752,N_4990);
xnor U5051 (N_5051,N_4998,N_4381);
nand U5052 (N_5052,N_4724,N_4881);
xnor U5053 (N_5053,N_4184,N_4613);
nand U5054 (N_5054,N_4967,N_4971);
nand U5055 (N_5055,N_4632,N_4677);
or U5056 (N_5056,N_4830,N_4171);
and U5057 (N_5057,N_4326,N_4586);
nor U5058 (N_5058,N_4387,N_4883);
nand U5059 (N_5059,N_4097,N_4493);
nand U5060 (N_5060,N_4736,N_4217);
xor U5061 (N_5061,N_4179,N_4029);
xor U5062 (N_5062,N_4470,N_4044);
and U5063 (N_5063,N_4347,N_4202);
nand U5064 (N_5064,N_4521,N_4524);
xor U5065 (N_5065,N_4251,N_4583);
nand U5066 (N_5066,N_4890,N_4385);
nand U5067 (N_5067,N_4140,N_4926);
and U5068 (N_5068,N_4523,N_4655);
nand U5069 (N_5069,N_4639,N_4449);
nand U5070 (N_5070,N_4804,N_4442);
or U5071 (N_5071,N_4942,N_4551);
and U5072 (N_5072,N_4134,N_4440);
xor U5073 (N_5073,N_4500,N_4336);
nand U5074 (N_5074,N_4640,N_4697);
or U5075 (N_5075,N_4570,N_4852);
nor U5076 (N_5076,N_4058,N_4832);
nor U5077 (N_5077,N_4077,N_4796);
and U5078 (N_5078,N_4966,N_4414);
nand U5079 (N_5079,N_4653,N_4137);
xnor U5080 (N_5080,N_4043,N_4460);
xor U5081 (N_5081,N_4838,N_4795);
nand U5082 (N_5082,N_4857,N_4010);
and U5083 (N_5083,N_4483,N_4855);
or U5084 (N_5084,N_4287,N_4413);
xor U5085 (N_5085,N_4656,N_4291);
nand U5086 (N_5086,N_4880,N_4782);
and U5087 (N_5087,N_4053,N_4907);
xnor U5088 (N_5088,N_4317,N_4643);
xnor U5089 (N_5089,N_4160,N_4879);
nand U5090 (N_5090,N_4725,N_4452);
nand U5091 (N_5091,N_4113,N_4258);
nand U5092 (N_5092,N_4709,N_4681);
nor U5093 (N_5093,N_4935,N_4556);
nand U5094 (N_5094,N_4215,N_4103);
or U5095 (N_5095,N_4581,N_4522);
nor U5096 (N_5096,N_4917,N_4631);
or U5097 (N_5097,N_4343,N_4259);
and U5098 (N_5098,N_4888,N_4970);
nand U5099 (N_5099,N_4313,N_4513);
nor U5100 (N_5100,N_4014,N_4525);
nand U5101 (N_5101,N_4800,N_4190);
and U5102 (N_5102,N_4728,N_4021);
or U5103 (N_5103,N_4188,N_4435);
and U5104 (N_5104,N_4684,N_4101);
and U5105 (N_5105,N_4318,N_4396);
nand U5106 (N_5106,N_4680,N_4212);
xor U5107 (N_5107,N_4647,N_4512);
or U5108 (N_5108,N_4474,N_4254);
and U5109 (N_5109,N_4105,N_4180);
nand U5110 (N_5110,N_4306,N_4818);
nand U5111 (N_5111,N_4913,N_4823);
xnor U5112 (N_5112,N_4519,N_4289);
and U5113 (N_5113,N_4430,N_4713);
xor U5114 (N_5114,N_4278,N_4749);
and U5115 (N_5115,N_4446,N_4905);
nand U5116 (N_5116,N_4548,N_4806);
and U5117 (N_5117,N_4220,N_4921);
and U5118 (N_5118,N_4411,N_4022);
xor U5119 (N_5119,N_4009,N_4087);
nor U5120 (N_5120,N_4841,N_4253);
and U5121 (N_5121,N_4247,N_4767);
or U5122 (N_5122,N_4480,N_4028);
nor U5123 (N_5123,N_4648,N_4734);
or U5124 (N_5124,N_4859,N_4775);
xnor U5125 (N_5125,N_4124,N_4408);
and U5126 (N_5126,N_4223,N_4987);
nor U5127 (N_5127,N_4471,N_4265);
and U5128 (N_5128,N_4371,N_4948);
or U5129 (N_5129,N_4266,N_4127);
nor U5130 (N_5130,N_4927,N_4074);
nand U5131 (N_5131,N_4788,N_4922);
nor U5132 (N_5132,N_4198,N_4887);
and U5133 (N_5133,N_4952,N_4506);
xor U5134 (N_5134,N_4017,N_4805);
nor U5135 (N_5135,N_4154,N_4013);
or U5136 (N_5136,N_4110,N_4495);
nand U5137 (N_5137,N_4748,N_4564);
nor U5138 (N_5138,N_4407,N_4981);
nand U5139 (N_5139,N_4610,N_4693);
or U5140 (N_5140,N_4863,N_4676);
nor U5141 (N_5141,N_4356,N_4900);
xor U5142 (N_5142,N_4270,N_4819);
xnor U5143 (N_5143,N_4547,N_4405);
nand U5144 (N_5144,N_4807,N_4955);
xor U5145 (N_5145,N_4057,N_4432);
and U5146 (N_5146,N_4003,N_4490);
or U5147 (N_5147,N_4542,N_4207);
or U5148 (N_5148,N_4923,N_4627);
nand U5149 (N_5149,N_4104,N_4912);
or U5150 (N_5150,N_4585,N_4731);
nor U5151 (N_5151,N_4540,N_4541);
xnor U5152 (N_5152,N_4319,N_4817);
nand U5153 (N_5153,N_4791,N_4634);
or U5154 (N_5154,N_4380,N_4866);
xnor U5155 (N_5155,N_4607,N_4236);
nand U5156 (N_5156,N_4325,N_4088);
xnor U5157 (N_5157,N_4031,N_4439);
or U5158 (N_5158,N_4238,N_4125);
and U5159 (N_5159,N_4897,N_4438);
xor U5160 (N_5160,N_4871,N_4433);
and U5161 (N_5161,N_4771,N_4756);
or U5162 (N_5162,N_4691,N_4295);
xnor U5163 (N_5163,N_4016,N_4173);
xnor U5164 (N_5164,N_4932,N_4307);
nand U5165 (N_5165,N_4060,N_4402);
nor U5166 (N_5166,N_4641,N_4930);
nor U5167 (N_5167,N_4936,N_4885);
or U5168 (N_5168,N_4115,N_4084);
or U5169 (N_5169,N_4428,N_4884);
xnor U5170 (N_5170,N_4753,N_4455);
xnor U5171 (N_5171,N_4148,N_4784);
xor U5172 (N_5172,N_4153,N_4142);
nand U5173 (N_5173,N_4194,N_4754);
nor U5174 (N_5174,N_4605,N_4039);
or U5175 (N_5175,N_4116,N_4315);
and U5176 (N_5176,N_4268,N_4650);
xor U5177 (N_5177,N_4974,N_4906);
and U5178 (N_5178,N_4657,N_4434);
nand U5179 (N_5179,N_4872,N_4679);
and U5180 (N_5180,N_4122,N_4595);
and U5181 (N_5181,N_4892,N_4934);
or U5182 (N_5182,N_4764,N_4946);
nor U5183 (N_5183,N_4001,N_4557);
or U5184 (N_5184,N_4781,N_4940);
xor U5185 (N_5185,N_4218,N_4667);
and U5186 (N_5186,N_4945,N_4185);
and U5187 (N_5187,N_4531,N_4624);
and U5188 (N_5188,N_4683,N_4666);
xor U5189 (N_5189,N_4367,N_4860);
nand U5190 (N_5190,N_4596,N_4199);
or U5191 (N_5191,N_4669,N_4532);
and U5192 (N_5192,N_4620,N_4530);
nor U5193 (N_5193,N_4415,N_4563);
and U5194 (N_5194,N_4505,N_4592);
and U5195 (N_5195,N_4304,N_4739);
xnor U5196 (N_5196,N_4893,N_4035);
nor U5197 (N_5197,N_4608,N_4156);
xnor U5198 (N_5198,N_4024,N_4929);
nor U5199 (N_5199,N_4089,N_4370);
nand U5200 (N_5200,N_4997,N_4033);
xor U5201 (N_5201,N_4334,N_4975);
or U5202 (N_5202,N_4978,N_4580);
and U5203 (N_5203,N_4394,N_4331);
nand U5204 (N_5204,N_4659,N_4100);
or U5205 (N_5205,N_4196,N_4297);
xnor U5206 (N_5206,N_4372,N_4050);
nor U5207 (N_5207,N_4600,N_4706);
xor U5208 (N_5208,N_4342,N_4665);
or U5209 (N_5209,N_4081,N_4555);
nor U5210 (N_5210,N_4719,N_4399);
or U5211 (N_5211,N_4886,N_4539);
nand U5212 (N_5212,N_4672,N_4208);
xnor U5213 (N_5213,N_4660,N_4205);
xor U5214 (N_5214,N_4763,N_4803);
xor U5215 (N_5215,N_4589,N_4023);
xor U5216 (N_5216,N_4423,N_4155);
or U5217 (N_5217,N_4450,N_4716);
nand U5218 (N_5218,N_4783,N_4690);
and U5219 (N_5219,N_4686,N_4037);
xor U5220 (N_5220,N_4111,N_4594);
nor U5221 (N_5221,N_4768,N_4496);
or U5222 (N_5222,N_4850,N_4568);
nor U5223 (N_5223,N_4544,N_4663);
nand U5224 (N_5224,N_4789,N_4451);
and U5225 (N_5225,N_4502,N_4891);
nor U5226 (N_5226,N_4882,N_4309);
nor U5227 (N_5227,N_4042,N_4409);
nor U5228 (N_5228,N_4808,N_4214);
nor U5229 (N_5229,N_4219,N_4458);
xor U5230 (N_5230,N_4072,N_4740);
and U5231 (N_5231,N_4237,N_4558);
xnor U5232 (N_5232,N_4661,N_4244);
nor U5233 (N_5233,N_4963,N_4165);
xnor U5234 (N_5234,N_4468,N_4526);
xnor U5235 (N_5235,N_4181,N_4296);
and U5236 (N_5236,N_4527,N_4330);
nand U5237 (N_5237,N_4011,N_4986);
xor U5238 (N_5238,N_4476,N_4569);
xor U5239 (N_5239,N_4840,N_4094);
and U5240 (N_5240,N_4075,N_4333);
or U5241 (N_5241,N_4876,N_4869);
xor U5242 (N_5242,N_4484,N_4834);
and U5243 (N_5243,N_4721,N_4117);
nor U5244 (N_5244,N_4138,N_4699);
nand U5245 (N_5245,N_4901,N_4720);
or U5246 (N_5246,N_4689,N_4573);
xnor U5247 (N_5247,N_4708,N_4406);
and U5248 (N_5248,N_4983,N_4671);
and U5249 (N_5249,N_4301,N_4777);
and U5250 (N_5250,N_4324,N_4412);
nor U5251 (N_5251,N_4729,N_4403);
nand U5252 (N_5252,N_4745,N_4327);
and U5253 (N_5253,N_4429,N_4515);
xor U5254 (N_5254,N_4635,N_4228);
nor U5255 (N_5255,N_4858,N_4472);
nor U5256 (N_5256,N_4168,N_4200);
nand U5257 (N_5257,N_4395,N_4492);
xor U5258 (N_5258,N_4112,N_4083);
xnor U5259 (N_5259,N_4943,N_4831);
and U5260 (N_5260,N_4478,N_4201);
or U5261 (N_5261,N_4799,N_4119);
and U5262 (N_5262,N_4126,N_4365);
and U5263 (N_5263,N_4135,N_4593);
and U5264 (N_5264,N_4972,N_4078);
nor U5265 (N_5265,N_4674,N_4933);
or U5266 (N_5266,N_4360,N_4738);
and U5267 (N_5267,N_4169,N_4707);
nor U5268 (N_5268,N_4508,N_4007);
nor U5269 (N_5269,N_4615,N_4828);
nand U5270 (N_5270,N_4132,N_4491);
nor U5271 (N_5271,N_4392,N_4744);
or U5272 (N_5272,N_4391,N_4070);
nand U5273 (N_5273,N_4562,N_4991);
nand U5274 (N_5274,N_4700,N_4419);
or U5275 (N_5275,N_4369,N_4267);
xnor U5276 (N_5276,N_4063,N_4567);
nand U5277 (N_5277,N_4827,N_4150);
and U5278 (N_5278,N_4311,N_4977);
xnor U5279 (N_5279,N_4552,N_4993);
nor U5280 (N_5280,N_4232,N_4487);
nand U5281 (N_5281,N_4264,N_4174);
nand U5282 (N_5282,N_4529,N_4166);
nor U5283 (N_5283,N_4163,N_4950);
and U5284 (N_5284,N_4376,N_4633);
nand U5285 (N_5285,N_4277,N_4488);
nor U5286 (N_5286,N_4146,N_4144);
nor U5287 (N_5287,N_4574,N_4209);
nor U5288 (N_5288,N_4861,N_4980);
and U5289 (N_5289,N_4454,N_4809);
and U5290 (N_5290,N_4284,N_4924);
or U5291 (N_5291,N_4899,N_4822);
and U5292 (N_5292,N_4790,N_4448);
nand U5293 (N_5293,N_4345,N_4427);
nor U5294 (N_5294,N_4283,N_4637);
nor U5295 (N_5295,N_4085,N_4045);
or U5296 (N_5296,N_4444,N_4750);
nor U5297 (N_5297,N_4462,N_4005);
nand U5298 (N_5298,N_4091,N_4717);
xor U5299 (N_5299,N_4560,N_4477);
or U5300 (N_5300,N_4849,N_4303);
or U5301 (N_5301,N_4896,N_4489);
and U5302 (N_5302,N_4835,N_4758);
and U5303 (N_5303,N_4918,N_4241);
and U5304 (N_5304,N_4008,N_4321);
nor U5305 (N_5305,N_4389,N_4846);
nor U5306 (N_5306,N_4549,N_4760);
or U5307 (N_5307,N_4239,N_4316);
and U5308 (N_5308,N_4704,N_4875);
nand U5309 (N_5309,N_4210,N_4421);
or U5310 (N_5310,N_4335,N_4614);
or U5311 (N_5311,N_4572,N_4159);
or U5312 (N_5312,N_4281,N_4006);
and U5313 (N_5313,N_4810,N_4959);
and U5314 (N_5314,N_4894,N_4951);
and U5315 (N_5315,N_4766,N_4695);
nor U5316 (N_5316,N_4761,N_4999);
xnor U5317 (N_5317,N_4565,N_4517);
or U5318 (N_5318,N_4664,N_4384);
and U5319 (N_5319,N_4167,N_4479);
and U5320 (N_5320,N_4629,N_4814);
nand U5321 (N_5321,N_4864,N_4466);
or U5322 (N_5322,N_4066,N_4062);
or U5323 (N_5323,N_4617,N_4914);
or U5324 (N_5324,N_4280,N_4393);
and U5325 (N_5325,N_4903,N_4420);
and U5326 (N_5326,N_4801,N_4279);
nor U5327 (N_5327,N_4157,N_4358);
nand U5328 (N_5328,N_4436,N_4410);
nor U5329 (N_5329,N_4718,N_4762);
nor U5330 (N_5330,N_4294,N_4341);
and U5331 (N_5331,N_4235,N_4973);
xor U5332 (N_5332,N_4388,N_4012);
nor U5333 (N_5333,N_4329,N_4030);
xor U5334 (N_5334,N_4692,N_4780);
nand U5335 (N_5335,N_4874,N_4302);
or U5336 (N_5336,N_4274,N_4445);
or U5337 (N_5337,N_4130,N_4038);
xnor U5338 (N_5338,N_4052,N_4988);
nand U5339 (N_5339,N_4377,N_4698);
nor U5340 (N_5340,N_4206,N_4305);
nor U5341 (N_5341,N_4867,N_4826);
or U5342 (N_5342,N_4765,N_4938);
nand U5343 (N_5343,N_4426,N_4383);
nor U5344 (N_5344,N_4786,N_4027);
nand U5345 (N_5345,N_4425,N_4919);
nor U5346 (N_5346,N_4151,N_4162);
nand U5347 (N_5347,N_4051,N_4726);
xor U5348 (N_5348,N_4510,N_4147);
and U5349 (N_5349,N_4459,N_4509);
nand U5350 (N_5350,N_4516,N_4064);
xnor U5351 (N_5351,N_4361,N_4400);
nor U5352 (N_5352,N_4743,N_4964);
nor U5353 (N_5353,N_4349,N_4645);
and U5354 (N_5354,N_4108,N_4588);
xnor U5355 (N_5355,N_4995,N_4920);
nor U5356 (N_5356,N_4131,N_4417);
or U5357 (N_5357,N_4862,N_4243);
or U5358 (N_5358,N_4953,N_4224);
or U5359 (N_5359,N_4275,N_4272);
xnor U5360 (N_5360,N_4979,N_4909);
xor U5361 (N_5361,N_4344,N_4465);
or U5362 (N_5362,N_4340,N_4514);
or U5363 (N_5363,N_4187,N_4957);
or U5364 (N_5364,N_4824,N_4067);
nand U5365 (N_5365,N_4216,N_4778);
nand U5366 (N_5366,N_4359,N_4504);
xor U5367 (N_5367,N_4298,N_4870);
xor U5368 (N_5368,N_4191,N_4949);
nor U5369 (N_5369,N_4628,N_4204);
xnor U5370 (N_5370,N_4183,N_4248);
nor U5371 (N_5371,N_4256,N_4584);
or U5372 (N_5372,N_4701,N_4833);
nor U5373 (N_5373,N_4961,N_4910);
or U5374 (N_5374,N_4651,N_4255);
xnor U5375 (N_5375,N_4742,N_4694);
nand U5376 (N_5376,N_4310,N_4164);
or U5377 (N_5377,N_4816,N_4904);
and U5378 (N_5378,N_4636,N_4386);
nor U5379 (N_5379,N_4546,N_4687);
and U5380 (N_5380,N_4056,N_4877);
xnor U5381 (N_5381,N_4582,N_4536);
nand U5382 (N_5382,N_4878,N_4982);
xnor U5383 (N_5383,N_4293,N_4213);
nand U5384 (N_5384,N_4069,N_4898);
xnor U5385 (N_5385,N_4350,N_4865);
nor U5386 (N_5386,N_4231,N_4732);
or U5387 (N_5387,N_4646,N_4312);
nand U5388 (N_5388,N_4366,N_4757);
nand U5389 (N_5389,N_4968,N_4242);
xnor U5390 (N_5390,N_4136,N_4511);
nand U5391 (N_5391,N_4328,N_4915);
nor U5392 (N_5392,N_4911,N_4996);
nand U5393 (N_5393,N_4048,N_4467);
or U5394 (N_5394,N_4673,N_4696);
and U5395 (N_5395,N_4245,N_4195);
and U5396 (N_5396,N_4260,N_4741);
nand U5397 (N_5397,N_4625,N_4338);
nor U5398 (N_5398,N_4606,N_4658);
xor U5399 (N_5399,N_4457,N_4203);
nand U5400 (N_5400,N_4836,N_4579);
or U5401 (N_5401,N_4193,N_4703);
xnor U5402 (N_5402,N_4792,N_4797);
xor U5403 (N_5403,N_4475,N_4958);
or U5404 (N_5404,N_4170,N_4469);
nand U5405 (N_5405,N_4908,N_4821);
xnor U5406 (N_5406,N_4630,N_4143);
and U5407 (N_5407,N_4109,N_4098);
nand U5408 (N_5408,N_4535,N_4211);
and U5409 (N_5409,N_4018,N_4261);
and U5410 (N_5410,N_4453,N_4263);
nor U5411 (N_5411,N_4618,N_4158);
xnor U5412 (N_5412,N_4292,N_4937);
xnor U5413 (N_5413,N_4348,N_4545);
nor U5414 (N_5414,N_4378,N_4785);
nand U5415 (N_5415,N_4501,N_4621);
xor U5416 (N_5416,N_4711,N_4854);
and U5417 (N_5417,N_4984,N_4186);
or U5418 (N_5418,N_4820,N_4346);
xor U5419 (N_5419,N_4553,N_4494);
xnor U5420 (N_5420,N_4604,N_4282);
nand U5421 (N_5421,N_4178,N_4250);
or U5422 (N_5422,N_4390,N_4947);
nor U5423 (N_5423,N_4000,N_4229);
and U5424 (N_5424,N_4839,N_4623);
or U5425 (N_5425,N_4082,N_4189);
nand U5426 (N_5426,N_4989,N_4362);
xnor U5427 (N_5427,N_4622,N_4481);
xor U5428 (N_5428,N_4240,N_4351);
xor U5429 (N_5429,N_4843,N_4576);
nand U5430 (N_5430,N_4577,N_4962);
nor U5431 (N_5431,N_4071,N_4422);
nand U5432 (N_5432,N_4269,N_4751);
nor U5433 (N_5433,N_4561,N_4705);
nand U5434 (N_5434,N_4299,N_4670);
and U5435 (N_5435,N_4099,N_4486);
nand U5436 (N_5436,N_4825,N_4619);
and U5437 (N_5437,N_4578,N_4715);
nor U5438 (N_5438,N_4710,N_4026);
or U5439 (N_5439,N_4668,N_4073);
nor U5440 (N_5440,N_4092,N_4107);
nand U5441 (N_5441,N_4276,N_4712);
xor U5442 (N_5442,N_4802,N_4076);
and U5443 (N_5443,N_4774,N_4447);
nand U5444 (N_5444,N_4845,N_4842);
nand U5445 (N_5445,N_4271,N_4550);
nand U5446 (N_5446,N_4373,N_4776);
xor U5447 (N_5447,N_4944,N_4599);
xor U5448 (N_5448,N_4290,N_4851);
nand U5449 (N_5449,N_4177,N_4285);
nor U5450 (N_5450,N_4222,N_4114);
xnor U5451 (N_5451,N_4093,N_4175);
and U5452 (N_5452,N_4288,N_4352);
nand U5453 (N_5453,N_4032,N_4723);
or U5454 (N_5454,N_4675,N_4049);
nand U5455 (N_5455,N_4262,N_4873);
and U5456 (N_5456,N_4040,N_4889);
nand U5457 (N_5457,N_4722,N_4688);
nor U5458 (N_5458,N_4339,N_4956);
nand U5459 (N_5459,N_4498,N_4714);
nand U5460 (N_5460,N_4994,N_4759);
or U5461 (N_5461,N_4856,N_4227);
xnor U5462 (N_5462,N_4813,N_4575);
nor U5463 (N_5463,N_4928,N_4020);
nand U5464 (N_5464,N_4482,N_4401);
nand U5465 (N_5465,N_4320,N_4096);
nand U5466 (N_5466,N_4518,N_4769);
xnor U5467 (N_5467,N_4379,N_4916);
or U5468 (N_5468,N_4638,N_4456);
and U5469 (N_5469,N_4603,N_4079);
nand U5470 (N_5470,N_4397,N_4461);
nor U5471 (N_5471,N_4375,N_4118);
nor U5472 (N_5472,N_4041,N_4682);
and U5473 (N_5473,N_4172,N_4353);
xnor U5474 (N_5474,N_4230,N_4902);
or U5475 (N_5475,N_4357,N_4609);
nand U5476 (N_5476,N_4848,N_4332);
and U5477 (N_5477,N_4418,N_4086);
nor U5478 (N_5478,N_4965,N_4895);
nor U5479 (N_5479,N_4424,N_4416);
nor U5480 (N_5480,N_4121,N_4811);
and U5481 (N_5481,N_4733,N_4794);
nand U5482 (N_5482,N_4234,N_4992);
xnor U5483 (N_5483,N_4793,N_4090);
and U5484 (N_5484,N_4503,N_4226);
or U5485 (N_5485,N_4123,N_4133);
or U5486 (N_5486,N_4554,N_4363);
and U5487 (N_5487,N_4566,N_4374);
and U5488 (N_5488,N_4139,N_4054);
and U5489 (N_5489,N_4678,N_4015);
nor U5490 (N_5490,N_4182,N_4837);
xor U5491 (N_5491,N_4931,N_4954);
or U5492 (N_5492,N_4192,N_4145);
xnor U5493 (N_5493,N_4437,N_4730);
nand U5494 (N_5494,N_4036,N_4770);
or U5495 (N_5495,N_4404,N_4652);
or U5496 (N_5496,N_4055,N_4004);
nand U5497 (N_5497,N_4538,N_4626);
and U5498 (N_5498,N_4985,N_4249);
and U5499 (N_5499,N_4141,N_4735);
or U5500 (N_5500,N_4079,N_4702);
and U5501 (N_5501,N_4832,N_4152);
xnor U5502 (N_5502,N_4474,N_4287);
nor U5503 (N_5503,N_4699,N_4717);
or U5504 (N_5504,N_4348,N_4418);
or U5505 (N_5505,N_4525,N_4453);
nand U5506 (N_5506,N_4880,N_4471);
and U5507 (N_5507,N_4253,N_4587);
nand U5508 (N_5508,N_4610,N_4749);
xnor U5509 (N_5509,N_4593,N_4204);
or U5510 (N_5510,N_4412,N_4375);
or U5511 (N_5511,N_4339,N_4967);
nand U5512 (N_5512,N_4933,N_4466);
and U5513 (N_5513,N_4601,N_4780);
xnor U5514 (N_5514,N_4074,N_4241);
nand U5515 (N_5515,N_4732,N_4578);
xnor U5516 (N_5516,N_4570,N_4730);
nand U5517 (N_5517,N_4634,N_4538);
and U5518 (N_5518,N_4950,N_4160);
nand U5519 (N_5519,N_4860,N_4538);
xor U5520 (N_5520,N_4400,N_4728);
nand U5521 (N_5521,N_4477,N_4026);
or U5522 (N_5522,N_4473,N_4585);
and U5523 (N_5523,N_4520,N_4358);
and U5524 (N_5524,N_4061,N_4281);
nor U5525 (N_5525,N_4176,N_4287);
xnor U5526 (N_5526,N_4656,N_4970);
or U5527 (N_5527,N_4210,N_4793);
xnor U5528 (N_5528,N_4755,N_4213);
nor U5529 (N_5529,N_4272,N_4992);
nor U5530 (N_5530,N_4670,N_4744);
nand U5531 (N_5531,N_4721,N_4081);
and U5532 (N_5532,N_4045,N_4320);
xnor U5533 (N_5533,N_4468,N_4867);
or U5534 (N_5534,N_4980,N_4344);
nand U5535 (N_5535,N_4031,N_4317);
xnor U5536 (N_5536,N_4939,N_4538);
or U5537 (N_5537,N_4608,N_4290);
xnor U5538 (N_5538,N_4117,N_4358);
nor U5539 (N_5539,N_4528,N_4724);
nand U5540 (N_5540,N_4798,N_4402);
xor U5541 (N_5541,N_4600,N_4623);
nor U5542 (N_5542,N_4143,N_4521);
xor U5543 (N_5543,N_4018,N_4768);
nor U5544 (N_5544,N_4040,N_4980);
nor U5545 (N_5545,N_4594,N_4435);
nor U5546 (N_5546,N_4991,N_4506);
or U5547 (N_5547,N_4694,N_4855);
xor U5548 (N_5548,N_4772,N_4402);
nand U5549 (N_5549,N_4227,N_4167);
or U5550 (N_5550,N_4953,N_4076);
or U5551 (N_5551,N_4346,N_4497);
and U5552 (N_5552,N_4784,N_4363);
or U5553 (N_5553,N_4040,N_4495);
or U5554 (N_5554,N_4272,N_4276);
nor U5555 (N_5555,N_4831,N_4501);
xor U5556 (N_5556,N_4272,N_4453);
xor U5557 (N_5557,N_4663,N_4164);
nand U5558 (N_5558,N_4017,N_4283);
or U5559 (N_5559,N_4446,N_4027);
or U5560 (N_5560,N_4236,N_4778);
nor U5561 (N_5561,N_4116,N_4722);
xor U5562 (N_5562,N_4800,N_4825);
nor U5563 (N_5563,N_4700,N_4358);
or U5564 (N_5564,N_4826,N_4890);
and U5565 (N_5565,N_4118,N_4014);
and U5566 (N_5566,N_4655,N_4089);
nor U5567 (N_5567,N_4429,N_4264);
nor U5568 (N_5568,N_4574,N_4088);
nand U5569 (N_5569,N_4390,N_4095);
and U5570 (N_5570,N_4898,N_4022);
xnor U5571 (N_5571,N_4070,N_4587);
and U5572 (N_5572,N_4209,N_4416);
nor U5573 (N_5573,N_4413,N_4138);
and U5574 (N_5574,N_4219,N_4670);
or U5575 (N_5575,N_4747,N_4441);
or U5576 (N_5576,N_4553,N_4303);
or U5577 (N_5577,N_4392,N_4275);
and U5578 (N_5578,N_4243,N_4642);
and U5579 (N_5579,N_4921,N_4391);
and U5580 (N_5580,N_4355,N_4688);
xnor U5581 (N_5581,N_4318,N_4278);
nand U5582 (N_5582,N_4510,N_4528);
or U5583 (N_5583,N_4156,N_4147);
or U5584 (N_5584,N_4703,N_4211);
nand U5585 (N_5585,N_4562,N_4768);
or U5586 (N_5586,N_4733,N_4721);
and U5587 (N_5587,N_4532,N_4042);
nand U5588 (N_5588,N_4039,N_4818);
nand U5589 (N_5589,N_4975,N_4400);
nand U5590 (N_5590,N_4904,N_4261);
or U5591 (N_5591,N_4992,N_4123);
xor U5592 (N_5592,N_4274,N_4657);
nor U5593 (N_5593,N_4283,N_4697);
xnor U5594 (N_5594,N_4487,N_4385);
nor U5595 (N_5595,N_4916,N_4626);
nand U5596 (N_5596,N_4596,N_4916);
nor U5597 (N_5597,N_4441,N_4654);
and U5598 (N_5598,N_4271,N_4835);
nand U5599 (N_5599,N_4749,N_4765);
and U5600 (N_5600,N_4420,N_4704);
nor U5601 (N_5601,N_4233,N_4333);
nand U5602 (N_5602,N_4652,N_4959);
or U5603 (N_5603,N_4142,N_4556);
nor U5604 (N_5604,N_4865,N_4926);
or U5605 (N_5605,N_4744,N_4108);
xor U5606 (N_5606,N_4116,N_4675);
and U5607 (N_5607,N_4834,N_4195);
or U5608 (N_5608,N_4371,N_4079);
or U5609 (N_5609,N_4664,N_4650);
nand U5610 (N_5610,N_4314,N_4723);
or U5611 (N_5611,N_4557,N_4815);
or U5612 (N_5612,N_4555,N_4654);
nand U5613 (N_5613,N_4049,N_4320);
or U5614 (N_5614,N_4449,N_4076);
and U5615 (N_5615,N_4008,N_4458);
xnor U5616 (N_5616,N_4557,N_4118);
nand U5617 (N_5617,N_4262,N_4009);
nor U5618 (N_5618,N_4243,N_4177);
and U5619 (N_5619,N_4170,N_4377);
and U5620 (N_5620,N_4861,N_4289);
nand U5621 (N_5621,N_4486,N_4575);
or U5622 (N_5622,N_4283,N_4890);
nor U5623 (N_5623,N_4872,N_4995);
nand U5624 (N_5624,N_4750,N_4535);
nand U5625 (N_5625,N_4863,N_4399);
nor U5626 (N_5626,N_4439,N_4531);
xor U5627 (N_5627,N_4362,N_4463);
or U5628 (N_5628,N_4989,N_4726);
and U5629 (N_5629,N_4731,N_4219);
and U5630 (N_5630,N_4776,N_4447);
or U5631 (N_5631,N_4090,N_4371);
nand U5632 (N_5632,N_4197,N_4401);
or U5633 (N_5633,N_4941,N_4964);
or U5634 (N_5634,N_4357,N_4022);
nand U5635 (N_5635,N_4165,N_4615);
nand U5636 (N_5636,N_4817,N_4003);
xnor U5637 (N_5637,N_4169,N_4591);
nand U5638 (N_5638,N_4001,N_4431);
and U5639 (N_5639,N_4019,N_4745);
xor U5640 (N_5640,N_4689,N_4778);
nor U5641 (N_5641,N_4167,N_4749);
and U5642 (N_5642,N_4440,N_4666);
nand U5643 (N_5643,N_4529,N_4693);
nor U5644 (N_5644,N_4686,N_4605);
xnor U5645 (N_5645,N_4617,N_4120);
or U5646 (N_5646,N_4654,N_4117);
and U5647 (N_5647,N_4744,N_4572);
or U5648 (N_5648,N_4608,N_4350);
xnor U5649 (N_5649,N_4873,N_4746);
nand U5650 (N_5650,N_4457,N_4440);
nor U5651 (N_5651,N_4608,N_4614);
or U5652 (N_5652,N_4181,N_4375);
or U5653 (N_5653,N_4244,N_4115);
nand U5654 (N_5654,N_4118,N_4882);
or U5655 (N_5655,N_4042,N_4279);
nand U5656 (N_5656,N_4634,N_4313);
nor U5657 (N_5657,N_4726,N_4723);
or U5658 (N_5658,N_4857,N_4375);
and U5659 (N_5659,N_4491,N_4963);
or U5660 (N_5660,N_4361,N_4147);
or U5661 (N_5661,N_4905,N_4524);
nand U5662 (N_5662,N_4538,N_4829);
or U5663 (N_5663,N_4340,N_4915);
nor U5664 (N_5664,N_4113,N_4680);
nor U5665 (N_5665,N_4397,N_4449);
and U5666 (N_5666,N_4817,N_4790);
xor U5667 (N_5667,N_4902,N_4718);
or U5668 (N_5668,N_4670,N_4819);
xnor U5669 (N_5669,N_4731,N_4734);
nor U5670 (N_5670,N_4270,N_4303);
xor U5671 (N_5671,N_4068,N_4471);
or U5672 (N_5672,N_4118,N_4466);
nor U5673 (N_5673,N_4734,N_4160);
nand U5674 (N_5674,N_4333,N_4146);
nor U5675 (N_5675,N_4371,N_4711);
nor U5676 (N_5676,N_4115,N_4475);
nor U5677 (N_5677,N_4484,N_4538);
or U5678 (N_5678,N_4450,N_4560);
or U5679 (N_5679,N_4164,N_4981);
nor U5680 (N_5680,N_4200,N_4329);
nand U5681 (N_5681,N_4575,N_4012);
nand U5682 (N_5682,N_4219,N_4833);
and U5683 (N_5683,N_4140,N_4919);
nand U5684 (N_5684,N_4977,N_4732);
and U5685 (N_5685,N_4378,N_4533);
nand U5686 (N_5686,N_4838,N_4532);
xor U5687 (N_5687,N_4998,N_4378);
and U5688 (N_5688,N_4527,N_4422);
or U5689 (N_5689,N_4060,N_4631);
nand U5690 (N_5690,N_4073,N_4636);
xnor U5691 (N_5691,N_4298,N_4326);
xor U5692 (N_5692,N_4918,N_4046);
nor U5693 (N_5693,N_4746,N_4789);
nand U5694 (N_5694,N_4699,N_4253);
nand U5695 (N_5695,N_4557,N_4912);
or U5696 (N_5696,N_4657,N_4046);
nor U5697 (N_5697,N_4760,N_4263);
or U5698 (N_5698,N_4532,N_4132);
nor U5699 (N_5699,N_4073,N_4359);
nor U5700 (N_5700,N_4192,N_4938);
nand U5701 (N_5701,N_4278,N_4375);
nor U5702 (N_5702,N_4494,N_4631);
nor U5703 (N_5703,N_4448,N_4484);
xor U5704 (N_5704,N_4301,N_4891);
or U5705 (N_5705,N_4907,N_4732);
nand U5706 (N_5706,N_4548,N_4816);
and U5707 (N_5707,N_4363,N_4225);
or U5708 (N_5708,N_4625,N_4300);
nor U5709 (N_5709,N_4722,N_4785);
and U5710 (N_5710,N_4851,N_4752);
nor U5711 (N_5711,N_4316,N_4451);
nor U5712 (N_5712,N_4973,N_4578);
nor U5713 (N_5713,N_4768,N_4755);
nor U5714 (N_5714,N_4173,N_4894);
xor U5715 (N_5715,N_4169,N_4752);
nand U5716 (N_5716,N_4886,N_4953);
nor U5717 (N_5717,N_4972,N_4416);
nand U5718 (N_5718,N_4521,N_4209);
or U5719 (N_5719,N_4785,N_4304);
and U5720 (N_5720,N_4604,N_4019);
and U5721 (N_5721,N_4010,N_4554);
nor U5722 (N_5722,N_4897,N_4088);
or U5723 (N_5723,N_4422,N_4100);
nor U5724 (N_5724,N_4080,N_4256);
nand U5725 (N_5725,N_4638,N_4488);
or U5726 (N_5726,N_4833,N_4652);
nor U5727 (N_5727,N_4718,N_4977);
nor U5728 (N_5728,N_4624,N_4401);
nor U5729 (N_5729,N_4056,N_4529);
and U5730 (N_5730,N_4030,N_4792);
and U5731 (N_5731,N_4864,N_4084);
nor U5732 (N_5732,N_4953,N_4581);
nand U5733 (N_5733,N_4361,N_4396);
nor U5734 (N_5734,N_4038,N_4904);
nor U5735 (N_5735,N_4050,N_4287);
xnor U5736 (N_5736,N_4242,N_4155);
xor U5737 (N_5737,N_4041,N_4936);
nand U5738 (N_5738,N_4947,N_4574);
and U5739 (N_5739,N_4194,N_4577);
or U5740 (N_5740,N_4108,N_4259);
or U5741 (N_5741,N_4377,N_4076);
xor U5742 (N_5742,N_4649,N_4586);
nand U5743 (N_5743,N_4153,N_4378);
or U5744 (N_5744,N_4201,N_4218);
nand U5745 (N_5745,N_4686,N_4462);
or U5746 (N_5746,N_4008,N_4747);
nand U5747 (N_5747,N_4156,N_4954);
and U5748 (N_5748,N_4211,N_4280);
nor U5749 (N_5749,N_4140,N_4956);
or U5750 (N_5750,N_4177,N_4765);
nor U5751 (N_5751,N_4441,N_4819);
nor U5752 (N_5752,N_4294,N_4342);
nor U5753 (N_5753,N_4070,N_4090);
or U5754 (N_5754,N_4715,N_4138);
nand U5755 (N_5755,N_4489,N_4309);
or U5756 (N_5756,N_4096,N_4933);
and U5757 (N_5757,N_4326,N_4628);
nor U5758 (N_5758,N_4599,N_4234);
or U5759 (N_5759,N_4692,N_4315);
or U5760 (N_5760,N_4832,N_4851);
or U5761 (N_5761,N_4375,N_4133);
xnor U5762 (N_5762,N_4103,N_4849);
nor U5763 (N_5763,N_4556,N_4932);
nand U5764 (N_5764,N_4541,N_4321);
xor U5765 (N_5765,N_4481,N_4448);
nand U5766 (N_5766,N_4824,N_4939);
xor U5767 (N_5767,N_4259,N_4387);
xor U5768 (N_5768,N_4592,N_4775);
xnor U5769 (N_5769,N_4828,N_4502);
nand U5770 (N_5770,N_4364,N_4735);
nor U5771 (N_5771,N_4115,N_4337);
nor U5772 (N_5772,N_4577,N_4706);
nor U5773 (N_5773,N_4598,N_4664);
nor U5774 (N_5774,N_4571,N_4477);
xor U5775 (N_5775,N_4938,N_4331);
nor U5776 (N_5776,N_4073,N_4731);
nand U5777 (N_5777,N_4584,N_4610);
xnor U5778 (N_5778,N_4714,N_4323);
nand U5779 (N_5779,N_4231,N_4310);
nand U5780 (N_5780,N_4824,N_4581);
nor U5781 (N_5781,N_4060,N_4256);
xor U5782 (N_5782,N_4555,N_4152);
xnor U5783 (N_5783,N_4457,N_4955);
xnor U5784 (N_5784,N_4760,N_4271);
nor U5785 (N_5785,N_4963,N_4672);
or U5786 (N_5786,N_4945,N_4143);
xor U5787 (N_5787,N_4566,N_4527);
and U5788 (N_5788,N_4737,N_4197);
nor U5789 (N_5789,N_4098,N_4559);
xnor U5790 (N_5790,N_4445,N_4336);
or U5791 (N_5791,N_4970,N_4911);
or U5792 (N_5792,N_4775,N_4067);
or U5793 (N_5793,N_4497,N_4357);
xnor U5794 (N_5794,N_4211,N_4409);
xor U5795 (N_5795,N_4923,N_4333);
xor U5796 (N_5796,N_4211,N_4264);
or U5797 (N_5797,N_4233,N_4185);
xnor U5798 (N_5798,N_4434,N_4443);
and U5799 (N_5799,N_4199,N_4444);
nor U5800 (N_5800,N_4384,N_4199);
xnor U5801 (N_5801,N_4926,N_4737);
nand U5802 (N_5802,N_4495,N_4764);
and U5803 (N_5803,N_4871,N_4507);
or U5804 (N_5804,N_4951,N_4015);
and U5805 (N_5805,N_4448,N_4825);
nor U5806 (N_5806,N_4682,N_4736);
nor U5807 (N_5807,N_4241,N_4391);
or U5808 (N_5808,N_4925,N_4009);
xnor U5809 (N_5809,N_4141,N_4606);
nand U5810 (N_5810,N_4046,N_4423);
or U5811 (N_5811,N_4595,N_4788);
or U5812 (N_5812,N_4849,N_4859);
or U5813 (N_5813,N_4480,N_4676);
nor U5814 (N_5814,N_4928,N_4495);
and U5815 (N_5815,N_4422,N_4535);
nand U5816 (N_5816,N_4289,N_4655);
or U5817 (N_5817,N_4133,N_4458);
xnor U5818 (N_5818,N_4018,N_4666);
xnor U5819 (N_5819,N_4784,N_4222);
or U5820 (N_5820,N_4657,N_4993);
xnor U5821 (N_5821,N_4733,N_4432);
nor U5822 (N_5822,N_4177,N_4054);
or U5823 (N_5823,N_4059,N_4130);
and U5824 (N_5824,N_4498,N_4898);
xnor U5825 (N_5825,N_4739,N_4683);
or U5826 (N_5826,N_4804,N_4253);
nand U5827 (N_5827,N_4780,N_4001);
nand U5828 (N_5828,N_4407,N_4989);
nor U5829 (N_5829,N_4960,N_4542);
nor U5830 (N_5830,N_4609,N_4768);
or U5831 (N_5831,N_4194,N_4855);
nor U5832 (N_5832,N_4357,N_4695);
nand U5833 (N_5833,N_4820,N_4476);
or U5834 (N_5834,N_4259,N_4799);
and U5835 (N_5835,N_4031,N_4620);
nor U5836 (N_5836,N_4624,N_4498);
xnor U5837 (N_5837,N_4194,N_4985);
nand U5838 (N_5838,N_4530,N_4657);
and U5839 (N_5839,N_4951,N_4219);
nand U5840 (N_5840,N_4287,N_4227);
nand U5841 (N_5841,N_4184,N_4550);
xnor U5842 (N_5842,N_4014,N_4317);
or U5843 (N_5843,N_4494,N_4469);
nand U5844 (N_5844,N_4750,N_4890);
or U5845 (N_5845,N_4218,N_4235);
nand U5846 (N_5846,N_4406,N_4342);
or U5847 (N_5847,N_4141,N_4817);
nor U5848 (N_5848,N_4700,N_4395);
nand U5849 (N_5849,N_4412,N_4644);
nor U5850 (N_5850,N_4068,N_4972);
or U5851 (N_5851,N_4047,N_4818);
nand U5852 (N_5852,N_4761,N_4705);
xor U5853 (N_5853,N_4370,N_4253);
nand U5854 (N_5854,N_4737,N_4484);
and U5855 (N_5855,N_4455,N_4013);
nand U5856 (N_5856,N_4426,N_4499);
nor U5857 (N_5857,N_4976,N_4248);
nor U5858 (N_5858,N_4931,N_4543);
nor U5859 (N_5859,N_4828,N_4392);
and U5860 (N_5860,N_4075,N_4318);
nor U5861 (N_5861,N_4882,N_4039);
and U5862 (N_5862,N_4809,N_4959);
nor U5863 (N_5863,N_4827,N_4081);
and U5864 (N_5864,N_4710,N_4423);
and U5865 (N_5865,N_4654,N_4113);
nor U5866 (N_5866,N_4451,N_4681);
or U5867 (N_5867,N_4513,N_4822);
nor U5868 (N_5868,N_4443,N_4755);
xnor U5869 (N_5869,N_4086,N_4913);
nand U5870 (N_5870,N_4450,N_4770);
or U5871 (N_5871,N_4121,N_4795);
nand U5872 (N_5872,N_4605,N_4151);
xnor U5873 (N_5873,N_4258,N_4710);
and U5874 (N_5874,N_4091,N_4403);
nand U5875 (N_5875,N_4004,N_4936);
and U5876 (N_5876,N_4134,N_4144);
nor U5877 (N_5877,N_4679,N_4251);
nand U5878 (N_5878,N_4483,N_4234);
xnor U5879 (N_5879,N_4900,N_4906);
nand U5880 (N_5880,N_4666,N_4674);
xor U5881 (N_5881,N_4280,N_4875);
or U5882 (N_5882,N_4774,N_4828);
nand U5883 (N_5883,N_4124,N_4590);
or U5884 (N_5884,N_4698,N_4570);
nor U5885 (N_5885,N_4523,N_4328);
xor U5886 (N_5886,N_4824,N_4144);
or U5887 (N_5887,N_4562,N_4632);
xnor U5888 (N_5888,N_4320,N_4766);
nor U5889 (N_5889,N_4681,N_4150);
and U5890 (N_5890,N_4121,N_4214);
nor U5891 (N_5891,N_4981,N_4696);
nand U5892 (N_5892,N_4769,N_4905);
or U5893 (N_5893,N_4101,N_4408);
nand U5894 (N_5894,N_4356,N_4512);
nor U5895 (N_5895,N_4044,N_4186);
and U5896 (N_5896,N_4333,N_4380);
and U5897 (N_5897,N_4862,N_4632);
and U5898 (N_5898,N_4472,N_4936);
and U5899 (N_5899,N_4553,N_4039);
nor U5900 (N_5900,N_4426,N_4801);
xnor U5901 (N_5901,N_4870,N_4940);
nand U5902 (N_5902,N_4511,N_4891);
nand U5903 (N_5903,N_4317,N_4910);
xnor U5904 (N_5904,N_4908,N_4939);
nand U5905 (N_5905,N_4662,N_4960);
xnor U5906 (N_5906,N_4897,N_4723);
nor U5907 (N_5907,N_4123,N_4731);
xor U5908 (N_5908,N_4316,N_4559);
xor U5909 (N_5909,N_4131,N_4927);
or U5910 (N_5910,N_4883,N_4187);
nand U5911 (N_5911,N_4826,N_4611);
xnor U5912 (N_5912,N_4009,N_4266);
nand U5913 (N_5913,N_4770,N_4575);
nor U5914 (N_5914,N_4376,N_4019);
nand U5915 (N_5915,N_4495,N_4193);
xnor U5916 (N_5916,N_4523,N_4540);
nand U5917 (N_5917,N_4419,N_4496);
and U5918 (N_5918,N_4011,N_4988);
nand U5919 (N_5919,N_4949,N_4157);
nand U5920 (N_5920,N_4233,N_4040);
and U5921 (N_5921,N_4235,N_4882);
nor U5922 (N_5922,N_4366,N_4846);
and U5923 (N_5923,N_4734,N_4540);
and U5924 (N_5924,N_4965,N_4298);
and U5925 (N_5925,N_4689,N_4282);
and U5926 (N_5926,N_4049,N_4190);
xnor U5927 (N_5927,N_4595,N_4719);
nor U5928 (N_5928,N_4774,N_4910);
and U5929 (N_5929,N_4440,N_4418);
or U5930 (N_5930,N_4839,N_4969);
or U5931 (N_5931,N_4469,N_4192);
or U5932 (N_5932,N_4365,N_4454);
nand U5933 (N_5933,N_4128,N_4728);
nor U5934 (N_5934,N_4389,N_4446);
and U5935 (N_5935,N_4096,N_4894);
nand U5936 (N_5936,N_4778,N_4858);
xnor U5937 (N_5937,N_4037,N_4325);
xnor U5938 (N_5938,N_4573,N_4868);
nand U5939 (N_5939,N_4300,N_4761);
and U5940 (N_5940,N_4057,N_4757);
nand U5941 (N_5941,N_4225,N_4951);
nand U5942 (N_5942,N_4087,N_4747);
or U5943 (N_5943,N_4919,N_4621);
xnor U5944 (N_5944,N_4573,N_4365);
or U5945 (N_5945,N_4182,N_4300);
nor U5946 (N_5946,N_4225,N_4030);
nand U5947 (N_5947,N_4167,N_4107);
xor U5948 (N_5948,N_4963,N_4334);
xnor U5949 (N_5949,N_4763,N_4830);
nor U5950 (N_5950,N_4218,N_4800);
xnor U5951 (N_5951,N_4836,N_4154);
nor U5952 (N_5952,N_4643,N_4611);
xor U5953 (N_5953,N_4854,N_4363);
and U5954 (N_5954,N_4403,N_4201);
nor U5955 (N_5955,N_4744,N_4454);
nor U5956 (N_5956,N_4838,N_4450);
nand U5957 (N_5957,N_4070,N_4567);
xor U5958 (N_5958,N_4788,N_4144);
xor U5959 (N_5959,N_4297,N_4036);
and U5960 (N_5960,N_4507,N_4003);
nand U5961 (N_5961,N_4901,N_4246);
and U5962 (N_5962,N_4765,N_4932);
xor U5963 (N_5963,N_4060,N_4314);
xnor U5964 (N_5964,N_4491,N_4449);
nand U5965 (N_5965,N_4646,N_4249);
nand U5966 (N_5966,N_4924,N_4635);
nor U5967 (N_5967,N_4683,N_4427);
nand U5968 (N_5968,N_4193,N_4093);
or U5969 (N_5969,N_4868,N_4933);
xnor U5970 (N_5970,N_4420,N_4456);
xor U5971 (N_5971,N_4862,N_4786);
nand U5972 (N_5972,N_4500,N_4516);
or U5973 (N_5973,N_4179,N_4106);
and U5974 (N_5974,N_4392,N_4415);
nor U5975 (N_5975,N_4375,N_4261);
and U5976 (N_5976,N_4640,N_4357);
xnor U5977 (N_5977,N_4001,N_4215);
xor U5978 (N_5978,N_4643,N_4341);
and U5979 (N_5979,N_4676,N_4091);
and U5980 (N_5980,N_4734,N_4703);
xnor U5981 (N_5981,N_4543,N_4129);
nand U5982 (N_5982,N_4285,N_4476);
and U5983 (N_5983,N_4353,N_4207);
and U5984 (N_5984,N_4878,N_4236);
or U5985 (N_5985,N_4650,N_4875);
nor U5986 (N_5986,N_4627,N_4530);
xor U5987 (N_5987,N_4352,N_4858);
nand U5988 (N_5988,N_4686,N_4925);
nor U5989 (N_5989,N_4185,N_4525);
or U5990 (N_5990,N_4869,N_4381);
xor U5991 (N_5991,N_4852,N_4341);
nor U5992 (N_5992,N_4352,N_4093);
nor U5993 (N_5993,N_4166,N_4199);
nand U5994 (N_5994,N_4803,N_4263);
nand U5995 (N_5995,N_4238,N_4640);
or U5996 (N_5996,N_4684,N_4130);
nand U5997 (N_5997,N_4805,N_4365);
or U5998 (N_5998,N_4516,N_4385);
nor U5999 (N_5999,N_4990,N_4052);
and U6000 (N_6000,N_5018,N_5832);
xnor U6001 (N_6001,N_5881,N_5588);
and U6002 (N_6002,N_5309,N_5241);
nand U6003 (N_6003,N_5087,N_5504);
nor U6004 (N_6004,N_5636,N_5254);
nand U6005 (N_6005,N_5161,N_5474);
xnor U6006 (N_6006,N_5243,N_5691);
nand U6007 (N_6007,N_5886,N_5908);
or U6008 (N_6008,N_5767,N_5188);
xor U6009 (N_6009,N_5748,N_5863);
xnor U6010 (N_6010,N_5493,N_5484);
nor U6011 (N_6011,N_5920,N_5805);
xnor U6012 (N_6012,N_5895,N_5455);
nand U6013 (N_6013,N_5155,N_5487);
or U6014 (N_6014,N_5048,N_5926);
and U6015 (N_6015,N_5007,N_5220);
nor U6016 (N_6016,N_5657,N_5806);
nor U6017 (N_6017,N_5456,N_5903);
or U6018 (N_6018,N_5150,N_5503);
nand U6019 (N_6019,N_5202,N_5560);
nor U6020 (N_6020,N_5968,N_5777);
xor U6021 (N_6021,N_5131,N_5184);
nor U6022 (N_6022,N_5169,N_5800);
nand U6023 (N_6023,N_5702,N_5818);
nor U6024 (N_6024,N_5125,N_5675);
or U6025 (N_6025,N_5017,N_5962);
xor U6026 (N_6026,N_5052,N_5313);
xnor U6027 (N_6027,N_5529,N_5699);
or U6028 (N_6028,N_5878,N_5937);
and U6029 (N_6029,N_5979,N_5860);
and U6030 (N_6030,N_5797,N_5472);
and U6031 (N_6031,N_5583,N_5020);
xor U6032 (N_6032,N_5597,N_5251);
nor U6033 (N_6033,N_5779,N_5177);
nor U6034 (N_6034,N_5708,N_5183);
nor U6035 (N_6035,N_5667,N_5760);
nand U6036 (N_6036,N_5872,N_5585);
nand U6037 (N_6037,N_5110,N_5301);
xor U6038 (N_6038,N_5397,N_5332);
and U6039 (N_6039,N_5793,N_5807);
nand U6040 (N_6040,N_5275,N_5513);
xnor U6041 (N_6041,N_5726,N_5743);
or U6042 (N_6042,N_5115,N_5506);
or U6043 (N_6043,N_5442,N_5199);
xnor U6044 (N_6044,N_5796,N_5178);
nand U6045 (N_6045,N_5817,N_5428);
xor U6046 (N_6046,N_5620,N_5540);
nor U6047 (N_6047,N_5780,N_5972);
nor U6048 (N_6048,N_5095,N_5684);
or U6049 (N_6049,N_5292,N_5252);
xor U6050 (N_6050,N_5151,N_5546);
xnor U6051 (N_6051,N_5399,N_5043);
nor U6052 (N_6052,N_5923,N_5651);
xnor U6053 (N_6053,N_5812,N_5149);
and U6054 (N_6054,N_5305,N_5745);
nand U6055 (N_6055,N_5333,N_5512);
nand U6056 (N_6056,N_5711,N_5804);
and U6057 (N_6057,N_5545,N_5887);
or U6058 (N_6058,N_5065,N_5727);
nand U6059 (N_6059,N_5490,N_5893);
or U6060 (N_6060,N_5785,N_5899);
xor U6061 (N_6061,N_5417,N_5717);
nor U6062 (N_6062,N_5622,N_5280);
nor U6063 (N_6063,N_5447,N_5337);
xnor U6064 (N_6064,N_5344,N_5694);
xnor U6065 (N_6065,N_5104,N_5200);
or U6066 (N_6066,N_5931,N_5764);
nand U6067 (N_6067,N_5852,N_5094);
and U6068 (N_6068,N_5024,N_5845);
xor U6069 (N_6069,N_5720,N_5320);
nor U6070 (N_6070,N_5196,N_5627);
nor U6071 (N_6071,N_5993,N_5297);
and U6072 (N_6072,N_5075,N_5864);
xor U6073 (N_6073,N_5380,N_5262);
and U6074 (N_6074,N_5752,N_5963);
and U6075 (N_6075,N_5730,N_5370);
or U6076 (N_6076,N_5366,N_5426);
xnor U6077 (N_6077,N_5824,N_5444);
and U6078 (N_6078,N_5359,N_5693);
or U6079 (N_6079,N_5973,N_5132);
and U6080 (N_6080,N_5851,N_5965);
or U6081 (N_6081,N_5143,N_5971);
xnor U6082 (N_6082,N_5408,N_5910);
nor U6083 (N_6083,N_5820,N_5680);
nand U6084 (N_6084,N_5642,N_5737);
or U6085 (N_6085,N_5057,N_5165);
and U6086 (N_6086,N_5871,N_5100);
nor U6087 (N_6087,N_5282,N_5565);
xnor U6088 (N_6088,N_5286,N_5076);
or U6089 (N_6089,N_5544,N_5211);
and U6090 (N_6090,N_5757,N_5722);
nand U6091 (N_6091,N_5739,N_5314);
xor U6092 (N_6092,N_5413,N_5716);
or U6093 (N_6093,N_5228,N_5395);
nor U6094 (N_6094,N_5549,N_5698);
and U6095 (N_6095,N_5023,N_5083);
xor U6096 (N_6096,N_5495,N_5326);
and U6097 (N_6097,N_5610,N_5367);
nand U6098 (N_6098,N_5523,N_5579);
and U6099 (N_6099,N_5436,N_5203);
or U6100 (N_6100,N_5081,N_5144);
nor U6101 (N_6101,N_5728,N_5011);
nand U6102 (N_6102,N_5526,N_5233);
nand U6103 (N_6103,N_5040,N_5858);
nor U6104 (N_6104,N_5891,N_5128);
or U6105 (N_6105,N_5576,N_5129);
xor U6106 (N_6106,N_5875,N_5515);
nand U6107 (N_6107,N_5185,N_5488);
or U6108 (N_6108,N_5283,N_5437);
or U6109 (N_6109,N_5054,N_5400);
nor U6110 (N_6110,N_5058,N_5645);
nor U6111 (N_6111,N_5232,N_5460);
and U6112 (N_6112,N_5363,N_5371);
nor U6113 (N_6113,N_5612,N_5528);
xor U6114 (N_6114,N_5402,N_5833);
nor U6115 (N_6115,N_5267,N_5205);
and U6116 (N_6116,N_5913,N_5531);
nor U6117 (N_6117,N_5510,N_5568);
nand U6118 (N_6118,N_5704,N_5475);
nand U6119 (N_6119,N_5936,N_5263);
nand U6120 (N_6120,N_5646,N_5195);
xor U6121 (N_6121,N_5681,N_5525);
nor U6122 (N_6122,N_5856,N_5022);
or U6123 (N_6123,N_5640,N_5935);
xor U6124 (N_6124,N_5892,N_5587);
or U6125 (N_6125,N_5897,N_5520);
and U6126 (N_6126,N_5758,N_5900);
or U6127 (N_6127,N_5669,N_5257);
xnor U6128 (N_6128,N_5330,N_5270);
and U6129 (N_6129,N_5616,N_5407);
xor U6130 (N_6130,N_5733,N_5404);
nor U6131 (N_6131,N_5609,N_5079);
xnor U6132 (N_6132,N_5957,N_5319);
nor U6133 (N_6133,N_5683,N_5181);
xnor U6134 (N_6134,N_5514,N_5273);
nand U6135 (N_6135,N_5999,N_5922);
or U6136 (N_6136,N_5418,N_5072);
nand U6137 (N_6137,N_5209,N_5665);
nand U6138 (N_6138,N_5331,N_5192);
xnor U6139 (N_6139,N_5450,N_5360);
and U6140 (N_6140,N_5541,N_5561);
nor U6141 (N_6141,N_5406,N_5118);
xnor U6142 (N_6142,N_5461,N_5245);
or U6143 (N_6143,N_5677,N_5844);
nor U6144 (N_6144,N_5168,N_5857);
xnor U6145 (N_6145,N_5825,N_5039);
nand U6146 (N_6146,N_5225,N_5633);
xor U6147 (N_6147,N_5160,N_5814);
nand U6148 (N_6148,N_5906,N_5924);
xor U6149 (N_6149,N_5298,N_5953);
and U6150 (N_6150,N_5207,N_5927);
nor U6151 (N_6151,N_5994,N_5074);
and U6152 (N_6152,N_5284,N_5005);
and U6153 (N_6153,N_5898,N_5032);
nand U6154 (N_6154,N_5316,N_5194);
or U6155 (N_6155,N_5421,N_5302);
and U6156 (N_6156,N_5984,N_5639);
nor U6157 (N_6157,N_5130,N_5457);
or U6158 (N_6158,N_5463,N_5916);
xnor U6159 (N_6159,N_5580,N_5046);
xor U6160 (N_6160,N_5859,N_5438);
or U6161 (N_6161,N_5385,N_5027);
nand U6162 (N_6162,N_5664,N_5443);
nand U6163 (N_6163,N_5932,N_5422);
or U6164 (N_6164,N_5409,N_5381);
nor U6165 (N_6165,N_5247,N_5819);
nand U6166 (N_6166,N_5062,N_5044);
nand U6167 (N_6167,N_5288,N_5603);
or U6168 (N_6168,N_5338,N_5123);
nor U6169 (N_6169,N_5101,N_5358);
xnor U6170 (N_6170,N_5483,N_5649);
xnor U6171 (N_6171,N_5986,N_5445);
xnor U6172 (N_6172,N_5988,N_5507);
xnor U6173 (N_6173,N_5364,N_5635);
nor U6174 (N_6174,N_5272,N_5003);
nor U6175 (N_6175,N_5547,N_5117);
and U6176 (N_6176,N_5686,N_5035);
nor U6177 (N_6177,N_5294,N_5532);
nand U6178 (N_6178,N_5264,N_5398);
xor U6179 (N_6179,N_5287,N_5031);
xor U6180 (N_6180,N_5846,N_5481);
xor U6181 (N_6181,N_5989,N_5479);
and U6182 (N_6182,N_5174,N_5171);
or U6183 (N_6183,N_5111,N_5379);
or U6184 (N_6184,N_5659,N_5765);
and U6185 (N_6185,N_5368,N_5223);
nand U6186 (N_6186,N_5138,N_5768);
nor U6187 (N_6187,N_5106,N_5253);
nor U6188 (N_6188,N_5411,N_5028);
nand U6189 (N_6189,N_5029,N_5362);
and U6190 (N_6190,N_5942,N_5557);
nand U6191 (N_6191,N_5705,N_5630);
or U6192 (N_6192,N_5574,N_5831);
or U6193 (N_6193,N_5480,N_5153);
and U6194 (N_6194,N_5734,N_5112);
nand U6195 (N_6195,N_5628,N_5629);
xor U6196 (N_6196,N_5911,N_5901);
xnor U6197 (N_6197,N_5811,N_5465);
nand U6198 (N_6198,N_5862,N_5033);
nor U6199 (N_6199,N_5749,N_5041);
and U6200 (N_6200,N_5985,N_5602);
nand U6201 (N_6201,N_5499,N_5497);
xor U6202 (N_6202,N_5950,N_5189);
xor U6203 (N_6203,N_5548,N_5321);
or U6204 (N_6204,N_5242,N_5036);
or U6205 (N_6205,N_5582,N_5822);
or U6206 (N_6206,N_5378,N_5116);
and U6207 (N_6207,N_5449,N_5981);
nor U6208 (N_6208,N_5345,N_5788);
nor U6209 (N_6209,N_5204,N_5158);
nand U6210 (N_6210,N_5896,N_5212);
and U6211 (N_6211,N_5414,N_5290);
nand U6212 (N_6212,N_5751,N_5256);
nand U6213 (N_6213,N_5429,N_5682);
nor U6214 (N_6214,N_5030,N_5873);
nand U6215 (N_6215,N_5536,N_5277);
and U6216 (N_6216,N_5631,N_5388);
nor U6217 (N_6217,N_5415,N_5867);
xor U6218 (N_6218,N_5542,N_5060);
and U6219 (N_6219,N_5139,N_5231);
nor U6220 (N_6220,N_5391,N_5615);
or U6221 (N_6221,N_5315,N_5865);
and U6222 (N_6222,N_5424,N_5842);
or U6223 (N_6223,N_5237,N_5260);
and U6224 (N_6224,N_5919,N_5619);
xor U6225 (N_6225,N_5918,N_5712);
or U6226 (N_6226,N_5921,N_5431);
xnor U6227 (N_6227,N_5672,N_5834);
xor U6228 (N_6228,N_5763,N_5586);
nand U6229 (N_6229,N_5700,N_5671);
nand U6230 (N_6230,N_5435,N_5375);
and U6231 (N_6231,N_5666,N_5869);
nand U6232 (N_6232,N_5991,N_5471);
xor U6233 (N_6233,N_5823,N_5605);
nor U6234 (N_6234,N_5689,N_5240);
xnor U6235 (N_6235,N_5750,N_5961);
or U6236 (N_6236,N_5038,N_5626);
or U6237 (N_6237,N_5732,N_5740);
nor U6238 (N_6238,N_5410,N_5102);
xnor U6239 (N_6239,N_5070,N_5230);
or U6240 (N_6240,N_5098,N_5372);
xor U6241 (N_6241,N_5441,N_5761);
nor U6242 (N_6242,N_5782,N_5077);
and U6243 (N_6243,N_5509,N_5051);
and U6244 (N_6244,N_5608,N_5222);
xor U6245 (N_6245,N_5006,N_5591);
or U6246 (N_6246,N_5519,N_5721);
and U6247 (N_6247,N_5904,N_5325);
nor U6248 (N_6248,N_5328,N_5170);
xnor U6249 (N_6249,N_5047,N_5323);
and U6250 (N_6250,N_5839,N_5949);
and U6251 (N_6251,N_5976,N_5945);
xnor U6252 (N_6252,N_5952,N_5599);
nor U6253 (N_6253,N_5652,N_5634);
xor U6254 (N_6254,N_5607,N_5502);
xor U6255 (N_6255,N_5855,N_5791);
or U6256 (N_6256,N_5182,N_5322);
nand U6257 (N_6257,N_5725,N_5928);
or U6258 (N_6258,N_5056,N_5880);
or U6259 (N_6259,N_5987,N_5941);
and U6260 (N_6260,N_5145,N_5756);
nand U6261 (N_6261,N_5648,N_5688);
xor U6262 (N_6262,N_5632,N_5654);
xor U6263 (N_6263,N_5001,N_5295);
nand U6264 (N_6264,N_5890,N_5550);
nor U6265 (N_6265,N_5351,N_5946);
and U6266 (N_6266,N_5709,N_5224);
nand U6267 (N_6267,N_5710,N_5762);
nand U6268 (N_6268,N_5135,N_5369);
nand U6269 (N_6269,N_5010,N_5889);
or U6270 (N_6270,N_5008,N_5173);
nand U6271 (N_6271,N_5097,N_5840);
nor U6272 (N_6272,N_5226,N_5933);
nand U6273 (N_6273,N_5556,N_5522);
nor U6274 (N_6274,N_5090,N_5217);
nor U6275 (N_6275,N_5318,N_5141);
and U6276 (N_6276,N_5156,N_5494);
and U6277 (N_6277,N_5731,N_5795);
or U6278 (N_6278,N_5473,N_5405);
xor U6279 (N_6279,N_5154,N_5190);
and U6280 (N_6280,N_5193,N_5943);
or U6281 (N_6281,N_5312,N_5821);
nand U6282 (N_6282,N_5462,N_5572);
or U6283 (N_6283,N_5279,N_5816);
xnor U6284 (N_6284,N_5496,N_5179);
nor U6285 (N_6285,N_5974,N_5324);
and U6286 (N_6286,N_5433,N_5361);
nand U6287 (N_6287,N_5637,N_5970);
xor U6288 (N_6288,N_5978,N_5085);
nor U6289 (N_6289,N_5109,N_5430);
or U6290 (N_6290,N_5012,N_5434);
and U6291 (N_6291,N_5221,N_5969);
nor U6292 (N_6292,N_5747,N_5653);
nand U6293 (N_6293,N_5208,N_5355);
nand U6294 (N_6294,N_5053,N_5951);
xnor U6295 (N_6295,N_5589,N_5492);
xnor U6296 (N_6296,N_5299,N_5459);
nand U6297 (N_6297,N_5660,N_5336);
and U6298 (N_6298,N_5960,N_5148);
nor U6299 (N_6299,N_5934,N_5902);
xor U6300 (N_6300,N_5621,N_5849);
or U6301 (N_6301,N_5142,N_5269);
nand U6302 (N_6302,N_5837,N_5274);
and U6303 (N_6303,N_5882,N_5786);
nor U6304 (N_6304,N_5829,N_5458);
or U6305 (N_6305,N_5658,N_5261);
nor U6306 (N_6306,N_5317,N_5088);
and U6307 (N_6307,N_5581,N_5291);
xnor U6308 (N_6308,N_5781,N_5894);
or U6309 (N_6309,N_5392,N_5964);
or U6310 (N_6310,N_5180,N_5162);
nor U6311 (N_6311,N_5715,N_5050);
nor U6312 (N_6312,N_5573,N_5827);
nor U6313 (N_6313,N_5690,N_5468);
xor U6314 (N_6314,N_5229,N_5082);
and U6315 (N_6315,N_5218,N_5644);
and U6316 (N_6316,N_5707,N_5592);
or U6317 (N_6317,N_5771,N_5349);
and U6318 (N_6318,N_5466,N_5673);
xor U6319 (N_6319,N_5197,N_5239);
and U6320 (N_6320,N_5157,N_5662);
nor U6321 (N_6321,N_5244,N_5879);
nor U6322 (N_6322,N_5527,N_5356);
nand U6323 (N_6323,N_5877,N_5485);
or U6324 (N_6324,N_5977,N_5836);
or U6325 (N_6325,N_5306,N_5915);
nand U6326 (N_6326,N_5870,N_5425);
or U6327 (N_6327,N_5365,N_5719);
xnor U6328 (N_6328,N_5215,N_5692);
xnor U6329 (N_6329,N_5009,N_5099);
and U6330 (N_6330,N_5334,N_5186);
and U6331 (N_6331,N_5427,N_5346);
or U6332 (N_6332,N_5813,N_5501);
or U6333 (N_6333,N_5108,N_5802);
xor U6334 (N_6334,N_5478,N_5925);
and U6335 (N_6335,N_5755,N_5888);
or U6336 (N_6336,N_5784,N_5685);
nand U6337 (N_6337,N_5084,N_5464);
nor U6338 (N_6338,N_5152,N_5086);
xor U6339 (N_6339,N_5695,N_5068);
nand U6340 (N_6340,N_5140,N_5015);
or U6341 (N_6341,N_5394,N_5907);
xnor U6342 (N_6342,N_5975,N_5838);
or U6343 (N_6343,N_5533,N_5067);
or U6344 (N_6344,N_5656,N_5470);
nand U6345 (N_6345,N_5929,N_5939);
or U6346 (N_6346,N_5697,N_5403);
or U6347 (N_6347,N_5219,N_5055);
nand U6348 (N_6348,N_5310,N_5335);
nor U6349 (N_6349,N_5980,N_5311);
xor U6350 (N_6350,N_5059,N_5611);
nor U6351 (N_6351,N_5249,N_5227);
nor U6352 (N_6352,N_5567,N_5376);
xor U6353 (N_6353,N_5163,N_5191);
xor U6354 (N_6354,N_5069,N_5448);
nor U6355 (N_6355,N_5396,N_5278);
or U6356 (N_6356,N_5146,N_5787);
nor U6357 (N_6357,N_5909,N_5614);
and U6358 (N_6358,N_5558,N_5638);
or U6359 (N_6359,N_5440,N_5049);
nor U6360 (N_6360,N_5308,N_5955);
nand U6361 (N_6361,N_5940,N_5948);
xor U6362 (N_6362,N_5167,N_5511);
and U6363 (N_6363,N_5250,N_5026);
or U6364 (N_6364,N_5105,N_5944);
or U6365 (N_6365,N_5451,N_5905);
or U6366 (N_6366,N_5759,N_5650);
nand U6367 (N_6367,N_5354,N_5661);
nand U6368 (N_6368,N_5300,N_5535);
or U6369 (N_6369,N_5701,N_5538);
nand U6370 (N_6370,N_5930,N_5995);
or U6371 (N_6371,N_5735,N_5738);
nand U6372 (N_6372,N_5555,N_5678);
and U6373 (N_6373,N_5647,N_5350);
and U6374 (N_6374,N_5293,N_5500);
nor U6375 (N_6375,N_5382,N_5353);
and U6376 (N_6376,N_5491,N_5384);
nor U6377 (N_6377,N_5071,N_5198);
nand U6378 (N_6378,N_5446,N_5884);
nor U6379 (N_6379,N_5296,N_5798);
xor U6380 (N_6380,N_5347,N_5486);
nor U6381 (N_6381,N_5617,N_5854);
nand U6382 (N_6382,N_5593,N_5096);
nand U6383 (N_6383,N_5259,N_5718);
xor U6384 (N_6384,N_5841,N_5983);
nand U6385 (N_6385,N_5093,N_5956);
or U6386 (N_6386,N_5792,N_5377);
nor U6387 (N_6387,N_5679,N_5214);
xor U6388 (N_6388,N_5452,N_5386);
nand U6389 (N_6389,N_5477,N_5073);
and U6390 (N_6390,N_5271,N_5537);
or U6391 (N_6391,N_5596,N_5172);
or U6392 (N_6392,N_5453,N_5216);
and U6393 (N_6393,N_5126,N_5454);
nor U6394 (N_6394,N_5606,N_5947);
and U6395 (N_6395,N_5164,N_5843);
nand U6396 (N_6396,N_5553,N_5516);
xnor U6397 (N_6397,N_5655,N_5103);
or U6398 (N_6398,N_5966,N_5618);
xor U6399 (N_6399,N_5569,N_5518);
nand U6400 (N_6400,N_5187,N_5476);
xor U6401 (N_6401,N_5663,N_5340);
and U6402 (N_6402,N_5789,N_5285);
or U6403 (N_6403,N_5571,N_5874);
or U6404 (N_6404,N_5566,N_5248);
or U6405 (N_6405,N_5815,N_5121);
xor U6406 (N_6406,N_5136,N_5080);
and U6407 (N_6407,N_5590,N_5482);
and U6408 (N_6408,N_5625,N_5773);
and U6409 (N_6409,N_5601,N_5373);
or U6410 (N_6410,N_5061,N_5517);
xnor U6411 (N_6411,N_5914,N_5954);
xor U6412 (N_6412,N_5120,N_5670);
and U6413 (N_6413,N_5958,N_5004);
and U6414 (N_6414,N_5255,N_5769);
nand U6415 (N_6415,N_5623,N_5210);
xor U6416 (N_6416,N_5265,N_5774);
and U6417 (N_6417,N_5534,N_5744);
nand U6418 (N_6418,N_5866,N_5159);
nor U6419 (N_6419,N_5643,N_5530);
or U6420 (N_6420,N_5352,N_5577);
nand U6421 (N_6421,N_5676,N_5013);
nand U6422 (N_6422,N_5133,N_5176);
nor U6423 (N_6423,N_5034,N_5713);
nor U6424 (N_6424,N_5303,N_5124);
nand U6425 (N_6425,N_5122,N_5401);
nand U6426 (N_6426,N_5706,N_5064);
nand U6427 (N_6427,N_5674,N_5432);
nor U6428 (N_6428,N_5268,N_5357);
nor U6429 (N_6429,N_5343,N_5876);
xnor U6430 (N_6430,N_5754,N_5037);
nor U6431 (N_6431,N_5246,N_5772);
or U6432 (N_6432,N_5742,N_5967);
nand U6433 (N_6433,N_5341,N_5604);
nand U6434 (N_6434,N_5770,N_5420);
or U6435 (N_6435,N_5387,N_5508);
or U6436 (N_6436,N_5134,N_5575);
nand U6437 (N_6437,N_5724,N_5276);
or U6438 (N_6438,N_5808,N_5439);
nor U6439 (N_6439,N_5554,N_5753);
nand U6440 (N_6440,N_5137,N_5281);
nor U6441 (N_6441,N_5778,N_5883);
nor U6442 (N_6442,N_5019,N_5826);
and U6443 (N_6443,N_5998,N_5848);
or U6444 (N_6444,N_5114,N_5235);
xor U6445 (N_6445,N_5803,N_5783);
nand U6446 (N_6446,N_5938,N_5304);
and U6447 (N_6447,N_5119,N_5063);
and U6448 (N_6448,N_5078,N_5850);
nand U6449 (N_6449,N_5390,N_5595);
and U6450 (N_6450,N_5236,N_5594);
xor U6451 (N_6451,N_5696,N_5868);
nand U6452 (N_6452,N_5990,N_5000);
or U6453 (N_6453,N_5107,N_5810);
xor U6454 (N_6454,N_5912,N_5166);
nor U6455 (N_6455,N_5521,N_5042);
or U6456 (N_6456,N_5539,N_5348);
nand U6457 (N_6457,N_5289,N_5736);
xnor U6458 (N_6458,N_5578,N_5959);
and U6459 (N_6459,N_5543,N_5600);
xor U6460 (N_6460,N_5828,N_5147);
and U6461 (N_6461,N_5127,N_5835);
xor U6462 (N_6462,N_5861,N_5416);
nor U6463 (N_6463,N_5741,N_5258);
nor U6464 (N_6464,N_5498,N_5997);
nand U6465 (N_6465,N_5687,N_5584);
nor U6466 (N_6466,N_5801,N_5505);
xnor U6467 (N_6467,N_5563,N_5423);
nand U6468 (N_6468,N_5234,N_5982);
or U6469 (N_6469,N_5327,N_5393);
xor U6470 (N_6470,N_5342,N_5002);
nand U6471 (N_6471,N_5045,N_5552);
or U6472 (N_6472,N_5853,N_5489);
and U6473 (N_6473,N_5703,N_5089);
nor U6474 (N_6474,N_5014,N_5524);
or U6475 (N_6475,N_5266,N_5469);
and U6476 (N_6476,N_5917,N_5714);
and U6477 (N_6477,N_5794,N_5551);
and U6478 (N_6478,N_5809,N_5729);
nor U6479 (N_6479,N_5213,N_5790);
and U6480 (N_6480,N_5383,N_5723);
and U6481 (N_6481,N_5307,N_5412);
or U6482 (N_6482,N_5624,N_5374);
nor U6483 (N_6483,N_5996,N_5668);
and U6484 (N_6484,N_5847,N_5830);
xor U6485 (N_6485,N_5206,N_5992);
nor U6486 (N_6486,N_5613,N_5201);
and U6487 (N_6487,N_5113,N_5467);
nand U6488 (N_6488,N_5562,N_5025);
and U6489 (N_6489,N_5389,N_5175);
nor U6490 (N_6490,N_5021,N_5570);
nand U6491 (N_6491,N_5419,N_5598);
nor U6492 (N_6492,N_5776,N_5091);
nand U6493 (N_6493,N_5775,N_5092);
nor U6494 (N_6494,N_5559,N_5066);
or U6495 (N_6495,N_5746,N_5238);
or U6496 (N_6496,N_5885,N_5564);
or U6497 (N_6497,N_5339,N_5016);
xnor U6498 (N_6498,N_5641,N_5799);
nand U6499 (N_6499,N_5766,N_5329);
nor U6500 (N_6500,N_5097,N_5339);
xor U6501 (N_6501,N_5537,N_5247);
nand U6502 (N_6502,N_5941,N_5116);
or U6503 (N_6503,N_5583,N_5657);
xor U6504 (N_6504,N_5466,N_5461);
nor U6505 (N_6505,N_5144,N_5903);
xnor U6506 (N_6506,N_5068,N_5743);
nor U6507 (N_6507,N_5008,N_5038);
xnor U6508 (N_6508,N_5366,N_5045);
nand U6509 (N_6509,N_5921,N_5782);
and U6510 (N_6510,N_5527,N_5638);
or U6511 (N_6511,N_5203,N_5347);
or U6512 (N_6512,N_5969,N_5859);
nor U6513 (N_6513,N_5100,N_5046);
xor U6514 (N_6514,N_5005,N_5647);
or U6515 (N_6515,N_5359,N_5717);
or U6516 (N_6516,N_5461,N_5590);
or U6517 (N_6517,N_5862,N_5264);
and U6518 (N_6518,N_5108,N_5464);
or U6519 (N_6519,N_5289,N_5674);
xor U6520 (N_6520,N_5548,N_5999);
or U6521 (N_6521,N_5907,N_5779);
nand U6522 (N_6522,N_5054,N_5972);
nand U6523 (N_6523,N_5299,N_5412);
nand U6524 (N_6524,N_5993,N_5669);
nand U6525 (N_6525,N_5433,N_5605);
nor U6526 (N_6526,N_5051,N_5140);
nand U6527 (N_6527,N_5518,N_5510);
and U6528 (N_6528,N_5882,N_5694);
xor U6529 (N_6529,N_5736,N_5848);
xor U6530 (N_6530,N_5753,N_5243);
or U6531 (N_6531,N_5069,N_5472);
nor U6532 (N_6532,N_5662,N_5651);
nor U6533 (N_6533,N_5262,N_5080);
or U6534 (N_6534,N_5467,N_5090);
nor U6535 (N_6535,N_5806,N_5927);
and U6536 (N_6536,N_5241,N_5090);
xnor U6537 (N_6537,N_5761,N_5735);
nor U6538 (N_6538,N_5392,N_5849);
nand U6539 (N_6539,N_5642,N_5728);
or U6540 (N_6540,N_5970,N_5133);
and U6541 (N_6541,N_5472,N_5761);
xor U6542 (N_6542,N_5626,N_5472);
nor U6543 (N_6543,N_5542,N_5261);
nor U6544 (N_6544,N_5031,N_5401);
and U6545 (N_6545,N_5592,N_5309);
xor U6546 (N_6546,N_5859,N_5901);
xnor U6547 (N_6547,N_5503,N_5490);
or U6548 (N_6548,N_5418,N_5736);
nand U6549 (N_6549,N_5419,N_5205);
or U6550 (N_6550,N_5967,N_5316);
xnor U6551 (N_6551,N_5413,N_5431);
or U6552 (N_6552,N_5477,N_5838);
xor U6553 (N_6553,N_5100,N_5936);
nand U6554 (N_6554,N_5758,N_5844);
nor U6555 (N_6555,N_5165,N_5130);
nor U6556 (N_6556,N_5160,N_5247);
and U6557 (N_6557,N_5053,N_5579);
or U6558 (N_6558,N_5665,N_5838);
nand U6559 (N_6559,N_5337,N_5492);
nand U6560 (N_6560,N_5484,N_5943);
or U6561 (N_6561,N_5818,N_5365);
nand U6562 (N_6562,N_5928,N_5321);
and U6563 (N_6563,N_5238,N_5406);
or U6564 (N_6564,N_5194,N_5177);
nand U6565 (N_6565,N_5599,N_5311);
nand U6566 (N_6566,N_5832,N_5055);
or U6567 (N_6567,N_5943,N_5862);
xnor U6568 (N_6568,N_5971,N_5104);
nor U6569 (N_6569,N_5887,N_5287);
and U6570 (N_6570,N_5104,N_5276);
nand U6571 (N_6571,N_5760,N_5776);
and U6572 (N_6572,N_5676,N_5767);
or U6573 (N_6573,N_5122,N_5795);
nor U6574 (N_6574,N_5972,N_5150);
and U6575 (N_6575,N_5791,N_5298);
and U6576 (N_6576,N_5326,N_5702);
and U6577 (N_6577,N_5189,N_5045);
nor U6578 (N_6578,N_5851,N_5215);
and U6579 (N_6579,N_5975,N_5943);
nand U6580 (N_6580,N_5503,N_5292);
nand U6581 (N_6581,N_5579,N_5788);
nand U6582 (N_6582,N_5295,N_5719);
and U6583 (N_6583,N_5857,N_5496);
nor U6584 (N_6584,N_5765,N_5558);
xor U6585 (N_6585,N_5464,N_5394);
and U6586 (N_6586,N_5293,N_5699);
nor U6587 (N_6587,N_5753,N_5301);
and U6588 (N_6588,N_5085,N_5248);
xnor U6589 (N_6589,N_5554,N_5160);
or U6590 (N_6590,N_5513,N_5470);
nor U6591 (N_6591,N_5591,N_5025);
or U6592 (N_6592,N_5019,N_5040);
and U6593 (N_6593,N_5715,N_5635);
nand U6594 (N_6594,N_5016,N_5577);
nand U6595 (N_6595,N_5804,N_5663);
or U6596 (N_6596,N_5750,N_5766);
nor U6597 (N_6597,N_5771,N_5365);
nor U6598 (N_6598,N_5011,N_5589);
or U6599 (N_6599,N_5403,N_5580);
and U6600 (N_6600,N_5556,N_5789);
nor U6601 (N_6601,N_5137,N_5002);
and U6602 (N_6602,N_5884,N_5980);
or U6603 (N_6603,N_5693,N_5197);
or U6604 (N_6604,N_5538,N_5178);
nor U6605 (N_6605,N_5430,N_5196);
nand U6606 (N_6606,N_5817,N_5278);
nand U6607 (N_6607,N_5629,N_5960);
xor U6608 (N_6608,N_5581,N_5289);
or U6609 (N_6609,N_5987,N_5662);
or U6610 (N_6610,N_5430,N_5966);
xnor U6611 (N_6611,N_5043,N_5668);
xnor U6612 (N_6612,N_5265,N_5323);
and U6613 (N_6613,N_5363,N_5895);
and U6614 (N_6614,N_5566,N_5709);
and U6615 (N_6615,N_5778,N_5191);
or U6616 (N_6616,N_5628,N_5937);
xor U6617 (N_6617,N_5416,N_5169);
nand U6618 (N_6618,N_5665,N_5413);
and U6619 (N_6619,N_5435,N_5909);
xnor U6620 (N_6620,N_5060,N_5637);
nand U6621 (N_6621,N_5571,N_5750);
or U6622 (N_6622,N_5069,N_5981);
and U6623 (N_6623,N_5628,N_5183);
xor U6624 (N_6624,N_5112,N_5262);
xnor U6625 (N_6625,N_5894,N_5613);
or U6626 (N_6626,N_5861,N_5486);
nor U6627 (N_6627,N_5615,N_5564);
nor U6628 (N_6628,N_5141,N_5054);
nor U6629 (N_6629,N_5976,N_5234);
nand U6630 (N_6630,N_5178,N_5254);
nand U6631 (N_6631,N_5017,N_5597);
or U6632 (N_6632,N_5016,N_5277);
and U6633 (N_6633,N_5077,N_5242);
nand U6634 (N_6634,N_5613,N_5902);
or U6635 (N_6635,N_5950,N_5943);
xnor U6636 (N_6636,N_5073,N_5098);
nand U6637 (N_6637,N_5147,N_5622);
and U6638 (N_6638,N_5364,N_5124);
nand U6639 (N_6639,N_5939,N_5028);
or U6640 (N_6640,N_5340,N_5771);
xnor U6641 (N_6641,N_5827,N_5577);
nand U6642 (N_6642,N_5806,N_5612);
or U6643 (N_6643,N_5179,N_5057);
and U6644 (N_6644,N_5725,N_5025);
or U6645 (N_6645,N_5897,N_5472);
or U6646 (N_6646,N_5413,N_5008);
and U6647 (N_6647,N_5656,N_5069);
xor U6648 (N_6648,N_5557,N_5718);
or U6649 (N_6649,N_5061,N_5742);
xor U6650 (N_6650,N_5211,N_5997);
nand U6651 (N_6651,N_5387,N_5126);
nand U6652 (N_6652,N_5590,N_5831);
nand U6653 (N_6653,N_5859,N_5644);
and U6654 (N_6654,N_5194,N_5363);
nand U6655 (N_6655,N_5698,N_5154);
xnor U6656 (N_6656,N_5862,N_5212);
or U6657 (N_6657,N_5760,N_5240);
xnor U6658 (N_6658,N_5735,N_5034);
or U6659 (N_6659,N_5813,N_5154);
nand U6660 (N_6660,N_5885,N_5923);
nand U6661 (N_6661,N_5321,N_5282);
and U6662 (N_6662,N_5562,N_5260);
nor U6663 (N_6663,N_5686,N_5690);
nand U6664 (N_6664,N_5737,N_5932);
xor U6665 (N_6665,N_5344,N_5273);
and U6666 (N_6666,N_5288,N_5256);
or U6667 (N_6667,N_5012,N_5879);
nor U6668 (N_6668,N_5635,N_5020);
or U6669 (N_6669,N_5290,N_5064);
nand U6670 (N_6670,N_5472,N_5179);
xor U6671 (N_6671,N_5588,N_5627);
nand U6672 (N_6672,N_5827,N_5759);
nor U6673 (N_6673,N_5387,N_5599);
nor U6674 (N_6674,N_5761,N_5557);
or U6675 (N_6675,N_5716,N_5144);
xor U6676 (N_6676,N_5148,N_5752);
nand U6677 (N_6677,N_5649,N_5244);
nor U6678 (N_6678,N_5274,N_5553);
and U6679 (N_6679,N_5193,N_5881);
or U6680 (N_6680,N_5185,N_5112);
or U6681 (N_6681,N_5134,N_5821);
or U6682 (N_6682,N_5336,N_5734);
and U6683 (N_6683,N_5675,N_5177);
nor U6684 (N_6684,N_5105,N_5171);
or U6685 (N_6685,N_5532,N_5699);
and U6686 (N_6686,N_5321,N_5101);
or U6687 (N_6687,N_5403,N_5601);
nor U6688 (N_6688,N_5343,N_5621);
and U6689 (N_6689,N_5448,N_5954);
or U6690 (N_6690,N_5854,N_5712);
xor U6691 (N_6691,N_5525,N_5234);
and U6692 (N_6692,N_5147,N_5517);
nor U6693 (N_6693,N_5566,N_5930);
nor U6694 (N_6694,N_5830,N_5842);
nor U6695 (N_6695,N_5307,N_5732);
nor U6696 (N_6696,N_5879,N_5025);
nor U6697 (N_6697,N_5515,N_5795);
xnor U6698 (N_6698,N_5482,N_5415);
nand U6699 (N_6699,N_5346,N_5024);
or U6700 (N_6700,N_5776,N_5539);
nand U6701 (N_6701,N_5153,N_5666);
nor U6702 (N_6702,N_5221,N_5439);
xor U6703 (N_6703,N_5740,N_5469);
nor U6704 (N_6704,N_5606,N_5456);
nand U6705 (N_6705,N_5845,N_5884);
xor U6706 (N_6706,N_5751,N_5011);
nor U6707 (N_6707,N_5546,N_5672);
or U6708 (N_6708,N_5004,N_5337);
nor U6709 (N_6709,N_5826,N_5956);
nor U6710 (N_6710,N_5473,N_5608);
nor U6711 (N_6711,N_5536,N_5384);
or U6712 (N_6712,N_5344,N_5551);
or U6713 (N_6713,N_5944,N_5822);
or U6714 (N_6714,N_5906,N_5821);
nor U6715 (N_6715,N_5692,N_5539);
nor U6716 (N_6716,N_5233,N_5009);
nor U6717 (N_6717,N_5291,N_5316);
nor U6718 (N_6718,N_5194,N_5245);
nor U6719 (N_6719,N_5448,N_5607);
xnor U6720 (N_6720,N_5680,N_5386);
and U6721 (N_6721,N_5980,N_5299);
xnor U6722 (N_6722,N_5780,N_5108);
nand U6723 (N_6723,N_5507,N_5966);
nand U6724 (N_6724,N_5304,N_5642);
nand U6725 (N_6725,N_5385,N_5063);
and U6726 (N_6726,N_5745,N_5313);
or U6727 (N_6727,N_5657,N_5154);
nor U6728 (N_6728,N_5300,N_5876);
nand U6729 (N_6729,N_5925,N_5384);
xnor U6730 (N_6730,N_5221,N_5929);
and U6731 (N_6731,N_5122,N_5787);
nand U6732 (N_6732,N_5617,N_5579);
nand U6733 (N_6733,N_5986,N_5887);
or U6734 (N_6734,N_5104,N_5660);
nor U6735 (N_6735,N_5847,N_5320);
nor U6736 (N_6736,N_5746,N_5093);
nor U6737 (N_6737,N_5654,N_5928);
xor U6738 (N_6738,N_5518,N_5547);
nor U6739 (N_6739,N_5559,N_5903);
nor U6740 (N_6740,N_5181,N_5858);
nor U6741 (N_6741,N_5112,N_5699);
or U6742 (N_6742,N_5238,N_5205);
xor U6743 (N_6743,N_5988,N_5981);
and U6744 (N_6744,N_5667,N_5238);
nor U6745 (N_6745,N_5951,N_5879);
nand U6746 (N_6746,N_5161,N_5229);
nand U6747 (N_6747,N_5891,N_5532);
or U6748 (N_6748,N_5676,N_5459);
or U6749 (N_6749,N_5823,N_5496);
and U6750 (N_6750,N_5486,N_5028);
and U6751 (N_6751,N_5159,N_5954);
xor U6752 (N_6752,N_5958,N_5498);
nand U6753 (N_6753,N_5671,N_5956);
xnor U6754 (N_6754,N_5037,N_5851);
and U6755 (N_6755,N_5054,N_5613);
xor U6756 (N_6756,N_5298,N_5944);
or U6757 (N_6757,N_5314,N_5934);
and U6758 (N_6758,N_5617,N_5634);
and U6759 (N_6759,N_5379,N_5356);
nand U6760 (N_6760,N_5950,N_5455);
nand U6761 (N_6761,N_5022,N_5547);
xor U6762 (N_6762,N_5900,N_5586);
or U6763 (N_6763,N_5206,N_5813);
xnor U6764 (N_6764,N_5439,N_5396);
or U6765 (N_6765,N_5603,N_5008);
xnor U6766 (N_6766,N_5522,N_5160);
nor U6767 (N_6767,N_5721,N_5357);
nand U6768 (N_6768,N_5320,N_5525);
nor U6769 (N_6769,N_5480,N_5398);
nand U6770 (N_6770,N_5964,N_5199);
and U6771 (N_6771,N_5490,N_5577);
nand U6772 (N_6772,N_5027,N_5153);
nand U6773 (N_6773,N_5351,N_5825);
nor U6774 (N_6774,N_5044,N_5556);
and U6775 (N_6775,N_5896,N_5457);
and U6776 (N_6776,N_5607,N_5636);
or U6777 (N_6777,N_5202,N_5935);
and U6778 (N_6778,N_5130,N_5219);
or U6779 (N_6779,N_5416,N_5738);
and U6780 (N_6780,N_5300,N_5844);
xnor U6781 (N_6781,N_5928,N_5109);
or U6782 (N_6782,N_5157,N_5333);
and U6783 (N_6783,N_5787,N_5380);
or U6784 (N_6784,N_5215,N_5850);
nand U6785 (N_6785,N_5138,N_5869);
nand U6786 (N_6786,N_5368,N_5091);
and U6787 (N_6787,N_5956,N_5891);
and U6788 (N_6788,N_5727,N_5790);
or U6789 (N_6789,N_5571,N_5546);
nand U6790 (N_6790,N_5167,N_5036);
xor U6791 (N_6791,N_5296,N_5806);
nand U6792 (N_6792,N_5735,N_5326);
nand U6793 (N_6793,N_5816,N_5037);
nor U6794 (N_6794,N_5086,N_5480);
nand U6795 (N_6795,N_5523,N_5615);
nand U6796 (N_6796,N_5751,N_5734);
and U6797 (N_6797,N_5303,N_5384);
xor U6798 (N_6798,N_5192,N_5408);
and U6799 (N_6799,N_5687,N_5464);
nand U6800 (N_6800,N_5129,N_5398);
or U6801 (N_6801,N_5639,N_5902);
nor U6802 (N_6802,N_5444,N_5093);
or U6803 (N_6803,N_5846,N_5241);
nor U6804 (N_6804,N_5371,N_5074);
nand U6805 (N_6805,N_5981,N_5188);
nor U6806 (N_6806,N_5928,N_5476);
and U6807 (N_6807,N_5492,N_5976);
xor U6808 (N_6808,N_5238,N_5351);
xnor U6809 (N_6809,N_5836,N_5512);
and U6810 (N_6810,N_5726,N_5143);
nand U6811 (N_6811,N_5209,N_5945);
nand U6812 (N_6812,N_5318,N_5431);
xor U6813 (N_6813,N_5240,N_5403);
nand U6814 (N_6814,N_5872,N_5270);
or U6815 (N_6815,N_5497,N_5861);
xnor U6816 (N_6816,N_5263,N_5366);
or U6817 (N_6817,N_5730,N_5656);
and U6818 (N_6818,N_5480,N_5603);
nor U6819 (N_6819,N_5753,N_5273);
or U6820 (N_6820,N_5158,N_5260);
nor U6821 (N_6821,N_5474,N_5223);
and U6822 (N_6822,N_5966,N_5798);
nand U6823 (N_6823,N_5633,N_5921);
nor U6824 (N_6824,N_5894,N_5005);
nand U6825 (N_6825,N_5354,N_5537);
nand U6826 (N_6826,N_5470,N_5413);
nor U6827 (N_6827,N_5124,N_5756);
and U6828 (N_6828,N_5065,N_5825);
and U6829 (N_6829,N_5688,N_5633);
or U6830 (N_6830,N_5386,N_5798);
and U6831 (N_6831,N_5897,N_5533);
xor U6832 (N_6832,N_5487,N_5779);
or U6833 (N_6833,N_5130,N_5032);
or U6834 (N_6834,N_5241,N_5978);
nand U6835 (N_6835,N_5006,N_5483);
and U6836 (N_6836,N_5906,N_5175);
and U6837 (N_6837,N_5519,N_5457);
or U6838 (N_6838,N_5483,N_5922);
nand U6839 (N_6839,N_5177,N_5646);
or U6840 (N_6840,N_5707,N_5029);
or U6841 (N_6841,N_5616,N_5786);
and U6842 (N_6842,N_5476,N_5916);
nor U6843 (N_6843,N_5965,N_5288);
or U6844 (N_6844,N_5712,N_5025);
nand U6845 (N_6845,N_5208,N_5781);
nand U6846 (N_6846,N_5240,N_5914);
nor U6847 (N_6847,N_5393,N_5647);
and U6848 (N_6848,N_5467,N_5935);
nor U6849 (N_6849,N_5087,N_5391);
or U6850 (N_6850,N_5398,N_5158);
nand U6851 (N_6851,N_5094,N_5844);
nand U6852 (N_6852,N_5119,N_5804);
and U6853 (N_6853,N_5758,N_5666);
and U6854 (N_6854,N_5289,N_5132);
xnor U6855 (N_6855,N_5470,N_5244);
nand U6856 (N_6856,N_5517,N_5463);
or U6857 (N_6857,N_5183,N_5755);
xor U6858 (N_6858,N_5337,N_5780);
or U6859 (N_6859,N_5605,N_5546);
nor U6860 (N_6860,N_5325,N_5614);
xnor U6861 (N_6861,N_5227,N_5375);
or U6862 (N_6862,N_5962,N_5006);
and U6863 (N_6863,N_5199,N_5033);
xor U6864 (N_6864,N_5682,N_5586);
xor U6865 (N_6865,N_5118,N_5497);
nand U6866 (N_6866,N_5952,N_5204);
or U6867 (N_6867,N_5812,N_5900);
and U6868 (N_6868,N_5570,N_5916);
xnor U6869 (N_6869,N_5019,N_5152);
xnor U6870 (N_6870,N_5335,N_5624);
xnor U6871 (N_6871,N_5520,N_5997);
or U6872 (N_6872,N_5501,N_5420);
nor U6873 (N_6873,N_5103,N_5534);
or U6874 (N_6874,N_5573,N_5474);
nand U6875 (N_6875,N_5339,N_5476);
or U6876 (N_6876,N_5416,N_5558);
or U6877 (N_6877,N_5258,N_5541);
nand U6878 (N_6878,N_5842,N_5591);
and U6879 (N_6879,N_5647,N_5781);
and U6880 (N_6880,N_5559,N_5546);
nor U6881 (N_6881,N_5494,N_5885);
and U6882 (N_6882,N_5181,N_5536);
or U6883 (N_6883,N_5612,N_5448);
xor U6884 (N_6884,N_5174,N_5299);
nor U6885 (N_6885,N_5556,N_5294);
nand U6886 (N_6886,N_5201,N_5680);
nor U6887 (N_6887,N_5445,N_5007);
and U6888 (N_6888,N_5731,N_5420);
and U6889 (N_6889,N_5602,N_5709);
or U6890 (N_6890,N_5268,N_5013);
or U6891 (N_6891,N_5050,N_5813);
and U6892 (N_6892,N_5745,N_5288);
xor U6893 (N_6893,N_5952,N_5354);
nand U6894 (N_6894,N_5232,N_5995);
xnor U6895 (N_6895,N_5684,N_5778);
nand U6896 (N_6896,N_5370,N_5430);
xnor U6897 (N_6897,N_5027,N_5360);
nor U6898 (N_6898,N_5494,N_5209);
nand U6899 (N_6899,N_5904,N_5515);
and U6900 (N_6900,N_5282,N_5570);
nand U6901 (N_6901,N_5576,N_5156);
or U6902 (N_6902,N_5658,N_5511);
and U6903 (N_6903,N_5797,N_5713);
and U6904 (N_6904,N_5672,N_5095);
xor U6905 (N_6905,N_5413,N_5874);
and U6906 (N_6906,N_5367,N_5266);
nor U6907 (N_6907,N_5863,N_5064);
or U6908 (N_6908,N_5184,N_5588);
nor U6909 (N_6909,N_5743,N_5329);
xnor U6910 (N_6910,N_5021,N_5587);
nand U6911 (N_6911,N_5704,N_5742);
nor U6912 (N_6912,N_5142,N_5712);
nand U6913 (N_6913,N_5303,N_5192);
nand U6914 (N_6914,N_5609,N_5521);
or U6915 (N_6915,N_5136,N_5124);
nand U6916 (N_6916,N_5452,N_5325);
nand U6917 (N_6917,N_5744,N_5436);
nand U6918 (N_6918,N_5526,N_5364);
or U6919 (N_6919,N_5014,N_5425);
or U6920 (N_6920,N_5127,N_5008);
xor U6921 (N_6921,N_5779,N_5515);
or U6922 (N_6922,N_5018,N_5283);
nand U6923 (N_6923,N_5056,N_5238);
xor U6924 (N_6924,N_5747,N_5163);
nand U6925 (N_6925,N_5485,N_5923);
xnor U6926 (N_6926,N_5921,N_5239);
and U6927 (N_6927,N_5328,N_5906);
nand U6928 (N_6928,N_5295,N_5051);
and U6929 (N_6929,N_5779,N_5427);
xor U6930 (N_6930,N_5942,N_5881);
nor U6931 (N_6931,N_5594,N_5006);
or U6932 (N_6932,N_5839,N_5847);
nor U6933 (N_6933,N_5554,N_5051);
nor U6934 (N_6934,N_5875,N_5931);
and U6935 (N_6935,N_5099,N_5277);
or U6936 (N_6936,N_5457,N_5066);
nor U6937 (N_6937,N_5886,N_5007);
and U6938 (N_6938,N_5034,N_5229);
or U6939 (N_6939,N_5940,N_5587);
xor U6940 (N_6940,N_5465,N_5713);
and U6941 (N_6941,N_5865,N_5545);
nor U6942 (N_6942,N_5251,N_5352);
and U6943 (N_6943,N_5424,N_5533);
xor U6944 (N_6944,N_5592,N_5071);
nor U6945 (N_6945,N_5971,N_5985);
and U6946 (N_6946,N_5569,N_5798);
nand U6947 (N_6947,N_5370,N_5928);
nor U6948 (N_6948,N_5272,N_5517);
nor U6949 (N_6949,N_5514,N_5785);
nand U6950 (N_6950,N_5973,N_5151);
or U6951 (N_6951,N_5550,N_5889);
xnor U6952 (N_6952,N_5448,N_5819);
nor U6953 (N_6953,N_5607,N_5297);
xor U6954 (N_6954,N_5199,N_5952);
or U6955 (N_6955,N_5068,N_5996);
or U6956 (N_6956,N_5840,N_5121);
xor U6957 (N_6957,N_5716,N_5890);
or U6958 (N_6958,N_5723,N_5307);
nor U6959 (N_6959,N_5912,N_5051);
or U6960 (N_6960,N_5888,N_5876);
xor U6961 (N_6961,N_5600,N_5673);
or U6962 (N_6962,N_5338,N_5522);
nor U6963 (N_6963,N_5535,N_5596);
and U6964 (N_6964,N_5834,N_5446);
nand U6965 (N_6965,N_5629,N_5859);
xnor U6966 (N_6966,N_5680,N_5669);
or U6967 (N_6967,N_5740,N_5779);
or U6968 (N_6968,N_5760,N_5319);
nor U6969 (N_6969,N_5224,N_5050);
and U6970 (N_6970,N_5649,N_5133);
or U6971 (N_6971,N_5979,N_5877);
xnor U6972 (N_6972,N_5761,N_5482);
or U6973 (N_6973,N_5610,N_5659);
or U6974 (N_6974,N_5597,N_5952);
nand U6975 (N_6975,N_5725,N_5721);
nand U6976 (N_6976,N_5953,N_5968);
nand U6977 (N_6977,N_5642,N_5657);
nor U6978 (N_6978,N_5981,N_5053);
nand U6979 (N_6979,N_5424,N_5826);
and U6980 (N_6980,N_5271,N_5189);
xnor U6981 (N_6981,N_5238,N_5195);
or U6982 (N_6982,N_5052,N_5280);
xnor U6983 (N_6983,N_5427,N_5706);
or U6984 (N_6984,N_5833,N_5020);
nor U6985 (N_6985,N_5420,N_5393);
nor U6986 (N_6986,N_5267,N_5491);
and U6987 (N_6987,N_5278,N_5179);
or U6988 (N_6988,N_5980,N_5754);
xor U6989 (N_6989,N_5366,N_5688);
or U6990 (N_6990,N_5217,N_5192);
nor U6991 (N_6991,N_5061,N_5442);
and U6992 (N_6992,N_5367,N_5442);
and U6993 (N_6993,N_5267,N_5426);
nor U6994 (N_6994,N_5039,N_5674);
nand U6995 (N_6995,N_5267,N_5740);
nor U6996 (N_6996,N_5488,N_5242);
nor U6997 (N_6997,N_5572,N_5002);
nand U6998 (N_6998,N_5819,N_5619);
or U6999 (N_6999,N_5868,N_5979);
xor U7000 (N_7000,N_6796,N_6420);
nor U7001 (N_7001,N_6805,N_6424);
xnor U7002 (N_7002,N_6359,N_6211);
or U7003 (N_7003,N_6873,N_6586);
nor U7004 (N_7004,N_6109,N_6120);
or U7005 (N_7005,N_6015,N_6702);
or U7006 (N_7006,N_6752,N_6806);
or U7007 (N_7007,N_6325,N_6813);
and U7008 (N_7008,N_6934,N_6358);
or U7009 (N_7009,N_6923,N_6062);
nor U7010 (N_7010,N_6711,N_6701);
and U7011 (N_7011,N_6599,N_6123);
and U7012 (N_7012,N_6027,N_6587);
nor U7013 (N_7013,N_6496,N_6474);
and U7014 (N_7014,N_6432,N_6003);
and U7015 (N_7015,N_6994,N_6764);
and U7016 (N_7016,N_6465,N_6491);
or U7017 (N_7017,N_6938,N_6261);
or U7018 (N_7018,N_6052,N_6737);
nand U7019 (N_7019,N_6666,N_6126);
or U7020 (N_7020,N_6784,N_6925);
or U7021 (N_7021,N_6105,N_6088);
or U7022 (N_7022,N_6561,N_6556);
xnor U7023 (N_7023,N_6847,N_6384);
nor U7024 (N_7024,N_6210,N_6213);
xor U7025 (N_7025,N_6302,N_6115);
nand U7026 (N_7026,N_6636,N_6582);
xnor U7027 (N_7027,N_6960,N_6229);
xor U7028 (N_7028,N_6036,N_6795);
nand U7029 (N_7029,N_6481,N_6108);
nor U7030 (N_7030,N_6877,N_6060);
nand U7031 (N_7031,N_6324,N_6492);
nand U7032 (N_7032,N_6272,N_6695);
xor U7033 (N_7033,N_6131,N_6622);
and U7034 (N_7034,N_6292,N_6347);
xnor U7035 (N_7035,N_6043,N_6732);
and U7036 (N_7036,N_6346,N_6039);
nand U7037 (N_7037,N_6935,N_6146);
xor U7038 (N_7038,N_6137,N_6288);
nor U7039 (N_7039,N_6021,N_6722);
xnor U7040 (N_7040,N_6761,N_6687);
xor U7041 (N_7041,N_6768,N_6634);
nor U7042 (N_7042,N_6270,N_6117);
xnor U7043 (N_7043,N_6767,N_6281);
nand U7044 (N_7044,N_6755,N_6639);
nor U7045 (N_7045,N_6963,N_6215);
and U7046 (N_7046,N_6243,N_6940);
xor U7047 (N_7047,N_6607,N_6336);
or U7048 (N_7048,N_6199,N_6782);
and U7049 (N_7049,N_6204,N_6720);
xnor U7050 (N_7050,N_6476,N_6533);
nor U7051 (N_7051,N_6580,N_6590);
nor U7052 (N_7052,N_6071,N_6132);
nand U7053 (N_7053,N_6750,N_6462);
and U7054 (N_7054,N_6014,N_6408);
or U7055 (N_7055,N_6531,N_6896);
or U7056 (N_7056,N_6074,N_6611);
xor U7057 (N_7057,N_6901,N_6878);
or U7058 (N_7058,N_6852,N_6040);
or U7059 (N_7059,N_6827,N_6779);
and U7060 (N_7060,N_6808,N_6285);
xor U7061 (N_7061,N_6075,N_6621);
or U7062 (N_7062,N_6663,N_6678);
nand U7063 (N_7063,N_6328,N_6369);
xnor U7064 (N_7064,N_6943,N_6706);
nand U7065 (N_7065,N_6592,N_6684);
nor U7066 (N_7066,N_6958,N_6615);
xnor U7067 (N_7067,N_6274,N_6945);
nand U7068 (N_7068,N_6739,N_6380);
xor U7069 (N_7069,N_6151,N_6845);
and U7070 (N_7070,N_6828,N_6881);
nand U7071 (N_7071,N_6987,N_6600);
or U7072 (N_7072,N_6859,N_6220);
and U7073 (N_7073,N_6139,N_6961);
and U7074 (N_7074,N_6005,N_6522);
and U7075 (N_7075,N_6181,N_6682);
nor U7076 (N_7076,N_6889,N_6479);
xnor U7077 (N_7077,N_6754,N_6182);
nand U7078 (N_7078,N_6537,N_6501);
or U7079 (N_7079,N_6778,N_6447);
xnor U7080 (N_7080,N_6254,N_6050);
and U7081 (N_7081,N_6912,N_6564);
nand U7082 (N_7082,N_6147,N_6673);
or U7083 (N_7083,N_6967,N_6545);
and U7084 (N_7084,N_6977,N_6193);
nor U7085 (N_7085,N_6811,N_6023);
or U7086 (N_7086,N_6955,N_6936);
and U7087 (N_7087,N_6252,N_6797);
xnor U7088 (N_7088,N_6177,N_6295);
xnor U7089 (N_7089,N_6119,N_6649);
and U7090 (N_7090,N_6746,N_6077);
nand U7091 (N_7091,N_6762,N_6032);
and U7092 (N_7092,N_6233,N_6434);
or U7093 (N_7093,N_6583,N_6657);
nor U7094 (N_7094,N_6879,N_6905);
xnor U7095 (N_7095,N_6449,N_6268);
nand U7096 (N_7096,N_6148,N_6488);
and U7097 (N_7097,N_6831,N_6846);
nor U7098 (N_7098,N_6990,N_6662);
xnor U7099 (N_7099,N_6414,N_6610);
or U7100 (N_7100,N_6149,N_6171);
or U7101 (N_7101,N_6700,N_6323);
nand U7102 (N_7102,N_6184,N_6353);
nand U7103 (N_7103,N_6427,N_6020);
nand U7104 (N_7104,N_6874,N_6385);
or U7105 (N_7105,N_6947,N_6498);
nor U7106 (N_7106,N_6585,N_6511);
nor U7107 (N_7107,N_6224,N_6675);
xor U7108 (N_7108,N_6400,N_6532);
nand U7109 (N_7109,N_6225,N_6183);
nor U7110 (N_7110,N_6627,N_6195);
nor U7111 (N_7111,N_6697,N_6508);
or U7112 (N_7112,N_6815,N_6464);
nor U7113 (N_7113,N_6208,N_6708);
or U7114 (N_7114,N_6850,N_6266);
or U7115 (N_7115,N_6245,N_6275);
xor U7116 (N_7116,N_6058,N_6861);
and U7117 (N_7117,N_6306,N_6562);
or U7118 (N_7118,N_6355,N_6386);
nor U7119 (N_7119,N_6717,N_6076);
and U7120 (N_7120,N_6547,N_6396);
nor U7121 (N_7121,N_6168,N_6045);
xor U7122 (N_7122,N_6628,N_6357);
nor U7123 (N_7123,N_6853,N_6162);
xor U7124 (N_7124,N_6232,N_6127);
nor U7125 (N_7125,N_6202,N_6996);
nand U7126 (N_7126,N_6763,N_6188);
nand U7127 (N_7127,N_6803,N_6469);
nand U7128 (N_7128,N_6406,N_6944);
and U7129 (N_7129,N_6558,N_6055);
nor U7130 (N_7130,N_6291,N_6866);
nand U7131 (N_7131,N_6389,N_6696);
nand U7132 (N_7132,N_6267,N_6128);
or U7133 (N_7133,N_6626,N_6571);
or U7134 (N_7134,N_6167,N_6218);
nor U7135 (N_7135,N_6426,N_6235);
nand U7136 (N_7136,N_6569,N_6433);
nor U7137 (N_7137,N_6007,N_6000);
nor U7138 (N_7138,N_6789,N_6618);
nor U7139 (N_7139,N_6930,N_6614);
or U7140 (N_7140,N_6665,N_6284);
or U7141 (N_7141,N_6502,N_6373);
and U7142 (N_7142,N_6282,N_6051);
nand U7143 (N_7143,N_6388,N_6911);
or U7144 (N_7144,N_6589,N_6517);
or U7145 (N_7145,N_6379,N_6812);
nand U7146 (N_7146,N_6159,N_6951);
nand U7147 (N_7147,N_6334,N_6733);
nor U7148 (N_7148,N_6157,N_6054);
nor U7149 (N_7149,N_6907,N_6140);
nand U7150 (N_7150,N_6887,N_6487);
nor U7151 (N_7151,N_6500,N_6937);
nor U7152 (N_7152,N_6559,N_6613);
or U7153 (N_7153,N_6728,N_6271);
nand U7154 (N_7154,N_6772,N_6917);
or U7155 (N_7155,N_6402,N_6952);
nor U7156 (N_7156,N_6205,N_6982);
and U7157 (N_7157,N_6138,N_6608);
xor U7158 (N_7158,N_6953,N_6801);
nand U7159 (N_7159,N_6293,N_6770);
nand U7160 (N_7160,N_6651,N_6993);
nand U7161 (N_7161,N_6680,N_6578);
or U7162 (N_7162,N_6601,N_6099);
xnor U7163 (N_7163,N_6661,N_6056);
and U7164 (N_7164,N_6959,N_6361);
or U7165 (N_7165,N_6314,N_6290);
xnor U7166 (N_7166,N_6404,N_6693);
and U7167 (N_7167,N_6962,N_6834);
or U7168 (N_7168,N_6318,N_6134);
xnor U7169 (N_7169,N_6931,N_6011);
nor U7170 (N_7170,N_6572,N_6303);
and U7171 (N_7171,N_6593,N_6175);
xor U7172 (N_7172,N_6279,N_6774);
nand U7173 (N_7173,N_6124,N_6370);
and U7174 (N_7174,N_6121,N_6798);
nand U7175 (N_7175,N_6872,N_6928);
or U7176 (N_7176,N_6730,N_6226);
xor U7177 (N_7177,N_6342,N_6471);
nor U7178 (N_7178,N_6332,N_6046);
and U7179 (N_7179,N_6529,N_6247);
nor U7180 (N_7180,N_6942,N_6441);
nor U7181 (N_7181,N_6490,N_6360);
xnor U7182 (N_7182,N_6435,N_6929);
and U7183 (N_7183,N_6836,N_6786);
xnor U7184 (N_7184,N_6619,N_6024);
xor U7185 (N_7185,N_6956,N_6620);
and U7186 (N_7186,N_6681,N_6368);
nand U7187 (N_7187,N_6591,N_6891);
xor U7188 (N_7188,N_6659,N_6609);
xnor U7189 (N_7189,N_6350,N_6277);
xor U7190 (N_7190,N_6818,N_6102);
xnor U7191 (N_7191,N_6642,N_6792);
xor U7192 (N_7192,N_6849,N_6718);
nor U7193 (N_7193,N_6004,N_6486);
xor U7194 (N_7194,N_6315,N_6198);
nand U7195 (N_7195,N_6848,N_6504);
and U7196 (N_7196,N_6676,N_6297);
nor U7197 (N_7197,N_6894,N_6825);
nor U7198 (N_7198,N_6679,N_6044);
nand U7199 (N_7199,N_6807,N_6239);
nor U7200 (N_7200,N_6038,N_6069);
and U7201 (N_7201,N_6033,N_6524);
and U7202 (N_7202,N_6503,N_6214);
or U7203 (N_7203,N_6791,N_6799);
and U7204 (N_7204,N_6704,N_6908);
or U7205 (N_7205,N_6228,N_6317);
and U7206 (N_7206,N_6249,N_6641);
nor U7207 (N_7207,N_6841,N_6013);
or U7208 (N_7208,N_6209,N_6705);
or U7209 (N_7209,N_6244,N_6823);
or U7210 (N_7210,N_6440,N_6790);
xnor U7211 (N_7211,N_6523,N_6142);
or U7212 (N_7212,N_6345,N_6660);
and U7213 (N_7213,N_6640,N_6187);
and U7214 (N_7214,N_6480,N_6240);
nand U7215 (N_7215,N_6715,N_6566);
xnor U7216 (N_7216,N_6946,N_6727);
or U7217 (N_7217,N_6975,N_6869);
and U7218 (N_7218,N_6902,N_6731);
nand U7219 (N_7219,N_6810,N_6863);
or U7220 (N_7220,N_6231,N_6594);
nand U7221 (N_7221,N_6867,N_6478);
xnor U7222 (N_7222,N_6513,N_6716);
xnor U7223 (N_7223,N_6103,N_6802);
xor U7224 (N_7224,N_6100,N_6463);
or U7225 (N_7225,N_6816,N_6337);
nand U7226 (N_7226,N_6544,N_6253);
nor U7227 (N_7227,N_6352,N_6413);
xor U7228 (N_7228,N_6378,N_6980);
nor U7229 (N_7229,N_6506,N_6747);
nand U7230 (N_7230,N_6507,N_6703);
nand U7231 (N_7231,N_6179,N_6528);
nor U7232 (N_7232,N_6048,N_6821);
or U7233 (N_7233,N_6372,N_6410);
nand U7234 (N_7234,N_6312,N_6882);
or U7235 (N_7235,N_6387,N_6242);
or U7236 (N_7236,N_6976,N_6950);
nor U7237 (N_7237,N_6753,N_6114);
nor U7238 (N_7238,N_6992,N_6870);
and U7239 (N_7239,N_6824,N_6820);
xor U7240 (N_7240,N_6819,N_6629);
xnor U7241 (N_7241,N_6759,N_6073);
or U7242 (N_7242,N_6381,N_6065);
or U7243 (N_7243,N_6577,N_6444);
and U7244 (N_7244,N_6002,N_6264);
or U7245 (N_7245,N_6237,N_6677);
nand U7246 (N_7246,N_6542,N_6653);
nor U7247 (N_7247,N_6886,N_6319);
and U7248 (N_7248,N_6156,N_6596);
nor U7249 (N_7249,N_6671,N_6309);
nor U7250 (N_7250,N_6844,N_6223);
nor U7251 (N_7251,N_6757,N_6057);
and U7252 (N_7252,N_6258,N_6536);
xnor U7253 (N_7253,N_6383,N_6094);
nand U7254 (N_7254,N_6405,N_6415);
nand U7255 (N_7255,N_6246,N_6574);
nor U7256 (N_7256,N_6766,N_6751);
nand U7257 (N_7257,N_6407,N_6656);
nor U7258 (N_7258,N_6579,N_6448);
and U7259 (N_7259,N_6042,N_6316);
or U7260 (N_7260,N_6165,N_6203);
xor U7261 (N_7261,N_6145,N_6307);
nand U7262 (N_7262,N_6467,N_6118);
and U7263 (N_7263,N_6144,N_6829);
xnor U7264 (N_7264,N_6893,N_6106);
or U7265 (N_7265,N_6344,N_6161);
and U7266 (N_7266,N_6439,N_6280);
and U7267 (N_7267,N_6461,N_6493);
nand U7268 (N_7268,N_6672,N_6130);
or U7269 (N_7269,N_6445,N_6484);
nor U7270 (N_7270,N_6966,N_6351);
nor U7271 (N_7271,N_6550,N_6981);
or U7272 (N_7272,N_6918,N_6376);
nand U7273 (N_7273,N_6991,N_6670);
xor U7274 (N_7274,N_6890,N_6856);
nor U7275 (N_7275,N_6974,N_6921);
nor U7276 (N_7276,N_6397,N_6735);
or U7277 (N_7277,N_6540,N_6339);
or U7278 (N_7278,N_6089,N_6459);
nor U7279 (N_7279,N_6738,N_6301);
xnor U7280 (N_7280,N_6230,N_6749);
nor U7281 (N_7281,N_6296,N_6212);
xor U7282 (N_7282,N_6068,N_6926);
and U7283 (N_7283,N_6409,N_6690);
nand U7284 (N_7284,N_6260,N_6954);
nand U7285 (N_7285,N_6107,N_6541);
nand U7286 (N_7286,N_6969,N_6422);
or U7287 (N_7287,N_6826,N_6526);
xor U7288 (N_7288,N_6234,N_6416);
and U7289 (N_7289,N_6122,N_6565);
nand U7290 (N_7290,N_6257,N_6001);
or U7291 (N_7291,N_6173,N_6775);
nor U7292 (N_7292,N_6080,N_6914);
and U7293 (N_7293,N_6597,N_6605);
nor U7294 (N_7294,N_6860,N_6090);
nor U7295 (N_7295,N_6116,N_6986);
nand U7296 (N_7296,N_6871,N_6998);
and U7297 (N_7297,N_6273,N_6428);
xor U7298 (N_7298,N_6178,N_6645);
or U7299 (N_7299,N_6744,N_6830);
nor U7300 (N_7300,N_6129,N_6256);
or U7301 (N_7301,N_6606,N_6785);
or U7302 (N_7302,N_6341,N_6933);
nor U7303 (N_7303,N_6552,N_6190);
nor U7304 (N_7304,N_6340,N_6031);
or U7305 (N_7305,N_6322,N_6450);
nor U7306 (N_7306,N_6520,N_6059);
and U7307 (N_7307,N_6691,N_6644);
nand U7308 (N_7308,N_6236,N_6973);
or U7309 (N_7309,N_6294,N_6927);
nand U7310 (N_7310,N_6794,N_6398);
or U7311 (N_7311,N_6685,N_6028);
nor U7312 (N_7312,N_6989,N_6446);
and U7313 (N_7313,N_6141,N_6475);
or U7314 (N_7314,N_6984,N_6875);
nand U7315 (N_7315,N_6382,N_6516);
nor U7316 (N_7316,N_6452,N_6876);
nor U7317 (N_7317,N_6916,N_6771);
and U7318 (N_7318,N_6623,N_6192);
nand U7319 (N_7319,N_6391,N_6425);
and U7320 (N_7320,N_6091,N_6840);
nand U7321 (N_7321,N_6221,N_6421);
xor U7322 (N_7322,N_6988,N_6371);
xnor U7323 (N_7323,N_6308,N_6694);
nor U7324 (N_7324,N_6971,N_6842);
xor U7325 (N_7325,N_6723,N_6787);
or U7326 (N_7326,N_6631,N_6473);
or U7327 (N_7327,N_6919,N_6392);
and U7328 (N_7328,N_6979,N_6217);
and U7329 (N_7329,N_6985,N_6995);
xor U7330 (N_7330,N_6133,N_6009);
xor U7331 (N_7331,N_6393,N_6010);
nor U7332 (N_7332,N_6092,N_6897);
and U7333 (N_7333,N_6838,N_6299);
xnor U7334 (N_7334,N_6375,N_6111);
nor U7335 (N_7335,N_6788,N_6740);
nor U7336 (N_7336,N_6864,N_6843);
nand U7337 (N_7337,N_6457,N_6637);
or U7338 (N_7338,N_6166,N_6155);
nor U7339 (N_7339,N_6833,N_6983);
and U7340 (N_7340,N_6263,N_6535);
and U7341 (N_7341,N_6888,N_6412);
or U7342 (N_7342,N_6018,N_6783);
xnor U7343 (N_7343,N_6436,N_6904);
and U7344 (N_7344,N_6008,N_6241);
xor U7345 (N_7345,N_6250,N_6549);
xnor U7346 (N_7346,N_6468,N_6692);
and U7347 (N_7347,N_6868,N_6519);
or U7348 (N_7348,N_6910,N_6667);
or U7349 (N_7349,N_6510,N_6885);
or U7350 (N_7350,N_6632,N_6072);
or U7351 (N_7351,N_6278,N_6616);
and U7352 (N_7352,N_6742,N_6892);
or U7353 (N_7353,N_6276,N_6429);
or U7354 (N_7354,N_6049,N_6643);
xnor U7355 (N_7355,N_6403,N_6957);
nor U7356 (N_7356,N_6216,N_6712);
nor U7357 (N_7357,N_6721,N_6087);
and U7358 (N_7358,N_6924,N_6006);
nor U7359 (N_7359,N_6725,N_6136);
and U7360 (N_7360,N_6067,N_6814);
nand U7361 (N_7361,N_6758,N_6563);
xor U7362 (N_7362,N_6699,N_6084);
and U7363 (N_7363,N_6298,N_6689);
nand U7364 (N_7364,N_6800,N_6219);
and U7365 (N_7365,N_6365,N_6470);
nor U7366 (N_7366,N_6097,N_6698);
xor U7367 (N_7367,N_6553,N_6832);
or U7368 (N_7368,N_6970,N_6197);
xor U7369 (N_7369,N_6390,N_6070);
nor U7370 (N_7370,N_6654,N_6019);
nand U7371 (N_7371,N_6906,N_6576);
nor U7372 (N_7372,N_6238,N_6104);
or U7373 (N_7373,N_6624,N_6515);
and U7374 (N_7374,N_6017,N_6455);
and U7375 (N_7375,N_6079,N_6431);
xor U7376 (N_7376,N_6377,N_6186);
or U7377 (N_7377,N_6086,N_6153);
xor U7378 (N_7378,N_6858,N_6152);
nand U7379 (N_7379,N_6401,N_6207);
nand U7380 (N_7380,N_6809,N_6098);
or U7381 (N_7381,N_6169,N_6326);
or U7382 (N_7382,N_6939,N_6570);
nand U7383 (N_7383,N_6363,N_6330);
nor U7384 (N_7384,N_6898,N_6857);
and U7385 (N_7385,N_6456,N_6356);
or U7386 (N_7386,N_6736,N_6185);
and U7387 (N_7387,N_6546,N_6617);
or U7388 (N_7388,N_6367,N_6477);
or U7389 (N_7389,N_6743,N_6485);
nor U7390 (N_7390,N_6095,N_6313);
xnor U7391 (N_7391,N_6170,N_6082);
nand U7392 (N_7392,N_6534,N_6648);
nand U7393 (N_7393,N_6922,N_6612);
or U7394 (N_7394,N_6248,N_6012);
or U7395 (N_7395,N_6710,N_6063);
and U7396 (N_7396,N_6164,N_6729);
and U7397 (N_7397,N_6262,N_6555);
or U7398 (N_7398,N_6037,N_6997);
or U7399 (N_7399,N_6251,N_6652);
nand U7400 (N_7400,N_6430,N_6932);
or U7401 (N_7401,N_6920,N_6509);
nand U7402 (N_7402,N_6495,N_6411);
xor U7403 (N_7403,N_6756,N_6399);
nand U7404 (N_7404,N_6999,N_6568);
and U7405 (N_7405,N_6903,N_6349);
and U7406 (N_7406,N_6083,N_6965);
and U7407 (N_7407,N_6543,N_6304);
nand U7408 (N_7408,N_6438,N_6554);
nor U7409 (N_7409,N_6512,N_6530);
and U7410 (N_7410,N_6458,N_6518);
nand U7411 (N_7411,N_6968,N_6909);
or U7412 (N_7412,N_6683,N_6348);
nor U7413 (N_7413,N_6647,N_6707);
nand U7414 (N_7414,N_6595,N_6514);
nor U7415 (N_7415,N_6035,N_6061);
and U7416 (N_7416,N_6900,N_6964);
and U7417 (N_7417,N_6719,N_6598);
nand U7418 (N_7418,N_6442,N_6588);
xnor U7419 (N_7419,N_6135,N_6668);
nand U7420 (N_7420,N_6066,N_6200);
nor U7421 (N_7421,N_6113,N_6154);
xnor U7422 (N_7422,N_6047,N_6026);
nor U7423 (N_7423,N_6150,N_6854);
nand U7424 (N_7424,N_6776,N_6366);
xor U7425 (N_7425,N_6283,N_6305);
or U7426 (N_7426,N_6453,N_6822);
nand U7427 (N_7427,N_6745,N_6604);
nand U7428 (N_7428,N_6709,N_6201);
xnor U7429 (N_7429,N_6575,N_6483);
or U7430 (N_7430,N_6143,N_6472);
or U7431 (N_7431,N_6734,N_6669);
xor U7432 (N_7432,N_6034,N_6374);
and U7433 (N_7433,N_6194,N_6505);
or U7434 (N_7434,N_6286,N_6321);
and U7435 (N_7435,N_6658,N_6494);
xor U7436 (N_7436,N_6781,N_6913);
nand U7437 (N_7437,N_6206,N_6635);
xnor U7438 (N_7438,N_6338,N_6525);
or U7439 (N_7439,N_6101,N_6454);
xnor U7440 (N_7440,N_6176,N_6081);
and U7441 (N_7441,N_6567,N_6584);
nand U7442 (N_7442,N_6259,N_6551);
or U7443 (N_7443,N_6655,N_6110);
and U7444 (N_7444,N_6030,N_6633);
nand U7445 (N_7445,N_6630,N_6688);
nand U7446 (N_7446,N_6978,N_6343);
xor U7447 (N_7447,N_6418,N_6499);
nor U7448 (N_7448,N_6839,N_6741);
and U7449 (N_7449,N_6354,N_6310);
nor U7450 (N_7450,N_6451,N_6437);
nor U7451 (N_7451,N_6895,N_6760);
or U7452 (N_7452,N_6489,N_6646);
nor U7453 (N_7453,N_6602,N_6174);
or U7454 (N_7454,N_6603,N_6765);
and U7455 (N_7455,N_6329,N_6287);
nor U7456 (N_7456,N_6394,N_6016);
nand U7457 (N_7457,N_6674,N_6581);
nor U7458 (N_7458,N_6022,N_6748);
or U7459 (N_7459,N_6327,N_6265);
nand U7460 (N_7460,N_6053,N_6941);
or U7461 (N_7461,N_6064,N_6724);
or U7462 (N_7462,N_6899,N_6227);
xnor U7463 (N_7463,N_6527,N_6497);
xnor U7464 (N_7464,N_6096,N_6883);
xnor U7465 (N_7465,N_6180,N_6880);
and U7466 (N_7466,N_6112,N_6189);
nor U7467 (N_7467,N_6538,N_6865);
nand U7468 (N_7468,N_6364,N_6331);
and U7469 (N_7469,N_6638,N_6884);
xnor U7470 (N_7470,N_6196,N_6443);
nand U7471 (N_7471,N_6085,N_6466);
nor U7472 (N_7472,N_6125,N_6726);
or U7473 (N_7473,N_6686,N_6769);
or U7474 (N_7474,N_6158,N_6335);
or U7475 (N_7475,N_6333,N_6300);
nand U7476 (N_7476,N_6289,N_6191);
nor U7477 (N_7477,N_6862,N_6163);
nand U7478 (N_7478,N_6714,N_6650);
or U7479 (N_7479,N_6093,N_6172);
or U7480 (N_7480,N_6851,N_6419);
nor U7481 (N_7481,N_6460,N_6548);
xnor U7482 (N_7482,N_6949,N_6423);
nor U7483 (N_7483,N_6025,N_6539);
nor U7484 (N_7484,N_6713,N_6837);
nor U7485 (N_7485,N_6521,N_6972);
xnor U7486 (N_7486,N_6041,N_6417);
nor U7487 (N_7487,N_6777,N_6557);
or U7488 (N_7488,N_6804,N_6573);
or U7489 (N_7489,N_6780,N_6255);
nor U7490 (N_7490,N_6948,N_6773);
nand U7491 (N_7491,N_6362,N_6855);
or U7492 (N_7492,N_6311,N_6664);
and U7493 (N_7493,N_6160,N_6482);
nor U7494 (N_7494,N_6835,N_6029);
nand U7495 (N_7495,N_6395,N_6560);
xor U7496 (N_7496,N_6915,N_6320);
xor U7497 (N_7497,N_6625,N_6078);
xnor U7498 (N_7498,N_6793,N_6222);
and U7499 (N_7499,N_6269,N_6817);
or U7500 (N_7500,N_6458,N_6472);
and U7501 (N_7501,N_6691,N_6203);
nor U7502 (N_7502,N_6473,N_6742);
nand U7503 (N_7503,N_6814,N_6558);
nand U7504 (N_7504,N_6737,N_6764);
nor U7505 (N_7505,N_6497,N_6946);
and U7506 (N_7506,N_6589,N_6062);
nor U7507 (N_7507,N_6206,N_6017);
nand U7508 (N_7508,N_6797,N_6798);
and U7509 (N_7509,N_6316,N_6650);
xnor U7510 (N_7510,N_6550,N_6965);
nand U7511 (N_7511,N_6143,N_6905);
or U7512 (N_7512,N_6819,N_6990);
nor U7513 (N_7513,N_6698,N_6399);
nor U7514 (N_7514,N_6475,N_6747);
nor U7515 (N_7515,N_6158,N_6217);
or U7516 (N_7516,N_6620,N_6393);
nand U7517 (N_7517,N_6567,N_6926);
xor U7518 (N_7518,N_6764,N_6406);
nor U7519 (N_7519,N_6510,N_6137);
nand U7520 (N_7520,N_6281,N_6781);
or U7521 (N_7521,N_6294,N_6540);
and U7522 (N_7522,N_6772,N_6463);
nand U7523 (N_7523,N_6326,N_6537);
nand U7524 (N_7524,N_6100,N_6120);
xnor U7525 (N_7525,N_6748,N_6087);
xnor U7526 (N_7526,N_6965,N_6709);
and U7527 (N_7527,N_6925,N_6143);
nand U7528 (N_7528,N_6253,N_6813);
nor U7529 (N_7529,N_6047,N_6242);
nand U7530 (N_7530,N_6325,N_6217);
nand U7531 (N_7531,N_6664,N_6937);
nor U7532 (N_7532,N_6608,N_6408);
and U7533 (N_7533,N_6532,N_6071);
xnor U7534 (N_7534,N_6236,N_6827);
nand U7535 (N_7535,N_6330,N_6144);
nand U7536 (N_7536,N_6260,N_6478);
xnor U7537 (N_7537,N_6963,N_6591);
or U7538 (N_7538,N_6823,N_6998);
nor U7539 (N_7539,N_6142,N_6076);
nand U7540 (N_7540,N_6724,N_6333);
and U7541 (N_7541,N_6134,N_6594);
nor U7542 (N_7542,N_6099,N_6553);
xor U7543 (N_7543,N_6427,N_6443);
nand U7544 (N_7544,N_6406,N_6418);
and U7545 (N_7545,N_6705,N_6196);
nor U7546 (N_7546,N_6796,N_6506);
or U7547 (N_7547,N_6672,N_6836);
and U7548 (N_7548,N_6655,N_6237);
xnor U7549 (N_7549,N_6068,N_6996);
nor U7550 (N_7550,N_6746,N_6361);
and U7551 (N_7551,N_6546,N_6592);
and U7552 (N_7552,N_6739,N_6987);
nand U7553 (N_7553,N_6315,N_6314);
nand U7554 (N_7554,N_6368,N_6011);
nor U7555 (N_7555,N_6935,N_6003);
nor U7556 (N_7556,N_6516,N_6996);
nand U7557 (N_7557,N_6356,N_6148);
and U7558 (N_7558,N_6464,N_6805);
nor U7559 (N_7559,N_6784,N_6875);
nand U7560 (N_7560,N_6488,N_6410);
or U7561 (N_7561,N_6201,N_6952);
and U7562 (N_7562,N_6354,N_6905);
and U7563 (N_7563,N_6152,N_6513);
xnor U7564 (N_7564,N_6506,N_6391);
nor U7565 (N_7565,N_6310,N_6677);
and U7566 (N_7566,N_6747,N_6037);
or U7567 (N_7567,N_6142,N_6974);
xor U7568 (N_7568,N_6292,N_6283);
or U7569 (N_7569,N_6152,N_6966);
or U7570 (N_7570,N_6513,N_6818);
xnor U7571 (N_7571,N_6817,N_6522);
nor U7572 (N_7572,N_6922,N_6213);
nand U7573 (N_7573,N_6151,N_6542);
and U7574 (N_7574,N_6704,N_6601);
xnor U7575 (N_7575,N_6757,N_6078);
and U7576 (N_7576,N_6580,N_6106);
nand U7577 (N_7577,N_6368,N_6638);
xnor U7578 (N_7578,N_6078,N_6838);
nand U7579 (N_7579,N_6553,N_6158);
xnor U7580 (N_7580,N_6424,N_6085);
or U7581 (N_7581,N_6766,N_6021);
nand U7582 (N_7582,N_6985,N_6732);
nor U7583 (N_7583,N_6530,N_6466);
nand U7584 (N_7584,N_6210,N_6817);
or U7585 (N_7585,N_6680,N_6084);
nand U7586 (N_7586,N_6140,N_6416);
nand U7587 (N_7587,N_6465,N_6849);
xor U7588 (N_7588,N_6197,N_6326);
nand U7589 (N_7589,N_6707,N_6583);
xnor U7590 (N_7590,N_6899,N_6526);
and U7591 (N_7591,N_6509,N_6502);
nand U7592 (N_7592,N_6464,N_6867);
xor U7593 (N_7593,N_6550,N_6390);
and U7594 (N_7594,N_6554,N_6851);
or U7595 (N_7595,N_6870,N_6821);
xor U7596 (N_7596,N_6430,N_6941);
and U7597 (N_7597,N_6691,N_6823);
nand U7598 (N_7598,N_6959,N_6897);
xnor U7599 (N_7599,N_6700,N_6045);
nand U7600 (N_7600,N_6375,N_6564);
and U7601 (N_7601,N_6558,N_6982);
nand U7602 (N_7602,N_6902,N_6532);
nor U7603 (N_7603,N_6353,N_6234);
nor U7604 (N_7604,N_6781,N_6582);
xnor U7605 (N_7605,N_6734,N_6528);
nand U7606 (N_7606,N_6754,N_6574);
xor U7607 (N_7607,N_6729,N_6066);
and U7608 (N_7608,N_6901,N_6033);
or U7609 (N_7609,N_6655,N_6963);
and U7610 (N_7610,N_6727,N_6947);
nand U7611 (N_7611,N_6256,N_6662);
xor U7612 (N_7612,N_6643,N_6407);
or U7613 (N_7613,N_6975,N_6996);
nand U7614 (N_7614,N_6288,N_6800);
nand U7615 (N_7615,N_6335,N_6747);
xnor U7616 (N_7616,N_6701,N_6887);
xor U7617 (N_7617,N_6492,N_6762);
nand U7618 (N_7618,N_6703,N_6975);
nand U7619 (N_7619,N_6051,N_6089);
and U7620 (N_7620,N_6846,N_6888);
nor U7621 (N_7621,N_6786,N_6398);
or U7622 (N_7622,N_6161,N_6304);
nand U7623 (N_7623,N_6158,N_6077);
and U7624 (N_7624,N_6249,N_6841);
and U7625 (N_7625,N_6078,N_6953);
nor U7626 (N_7626,N_6239,N_6652);
and U7627 (N_7627,N_6300,N_6919);
or U7628 (N_7628,N_6131,N_6203);
and U7629 (N_7629,N_6241,N_6030);
nand U7630 (N_7630,N_6626,N_6235);
or U7631 (N_7631,N_6328,N_6900);
nor U7632 (N_7632,N_6073,N_6765);
xor U7633 (N_7633,N_6512,N_6207);
xnor U7634 (N_7634,N_6888,N_6072);
nor U7635 (N_7635,N_6007,N_6214);
nor U7636 (N_7636,N_6906,N_6622);
nor U7637 (N_7637,N_6025,N_6376);
nor U7638 (N_7638,N_6738,N_6851);
nand U7639 (N_7639,N_6734,N_6102);
and U7640 (N_7640,N_6580,N_6505);
xor U7641 (N_7641,N_6631,N_6477);
xnor U7642 (N_7642,N_6053,N_6664);
and U7643 (N_7643,N_6743,N_6028);
or U7644 (N_7644,N_6010,N_6043);
nor U7645 (N_7645,N_6794,N_6734);
nor U7646 (N_7646,N_6321,N_6590);
or U7647 (N_7647,N_6038,N_6121);
xnor U7648 (N_7648,N_6133,N_6199);
nor U7649 (N_7649,N_6774,N_6541);
and U7650 (N_7650,N_6141,N_6016);
xnor U7651 (N_7651,N_6427,N_6662);
or U7652 (N_7652,N_6656,N_6919);
nand U7653 (N_7653,N_6882,N_6979);
xor U7654 (N_7654,N_6587,N_6351);
nor U7655 (N_7655,N_6971,N_6295);
or U7656 (N_7656,N_6641,N_6305);
and U7657 (N_7657,N_6438,N_6824);
and U7658 (N_7658,N_6427,N_6111);
nand U7659 (N_7659,N_6769,N_6875);
nor U7660 (N_7660,N_6769,N_6855);
xnor U7661 (N_7661,N_6010,N_6979);
nor U7662 (N_7662,N_6036,N_6815);
or U7663 (N_7663,N_6142,N_6555);
nand U7664 (N_7664,N_6614,N_6243);
xor U7665 (N_7665,N_6276,N_6950);
and U7666 (N_7666,N_6054,N_6397);
and U7667 (N_7667,N_6588,N_6490);
and U7668 (N_7668,N_6076,N_6494);
or U7669 (N_7669,N_6074,N_6462);
nand U7670 (N_7670,N_6796,N_6094);
nand U7671 (N_7671,N_6779,N_6331);
xnor U7672 (N_7672,N_6908,N_6402);
and U7673 (N_7673,N_6081,N_6673);
and U7674 (N_7674,N_6391,N_6107);
or U7675 (N_7675,N_6744,N_6711);
xnor U7676 (N_7676,N_6812,N_6990);
nor U7677 (N_7677,N_6512,N_6770);
and U7678 (N_7678,N_6922,N_6128);
and U7679 (N_7679,N_6433,N_6508);
xor U7680 (N_7680,N_6635,N_6356);
xor U7681 (N_7681,N_6300,N_6882);
xnor U7682 (N_7682,N_6534,N_6817);
or U7683 (N_7683,N_6683,N_6182);
or U7684 (N_7684,N_6091,N_6636);
or U7685 (N_7685,N_6191,N_6595);
nand U7686 (N_7686,N_6598,N_6820);
and U7687 (N_7687,N_6507,N_6017);
nor U7688 (N_7688,N_6893,N_6637);
xor U7689 (N_7689,N_6173,N_6966);
or U7690 (N_7690,N_6279,N_6054);
nand U7691 (N_7691,N_6352,N_6619);
xnor U7692 (N_7692,N_6402,N_6440);
xor U7693 (N_7693,N_6180,N_6709);
and U7694 (N_7694,N_6957,N_6176);
xor U7695 (N_7695,N_6969,N_6544);
and U7696 (N_7696,N_6268,N_6959);
xnor U7697 (N_7697,N_6826,N_6832);
or U7698 (N_7698,N_6184,N_6439);
and U7699 (N_7699,N_6750,N_6891);
and U7700 (N_7700,N_6021,N_6038);
and U7701 (N_7701,N_6054,N_6879);
or U7702 (N_7702,N_6266,N_6775);
or U7703 (N_7703,N_6073,N_6672);
xnor U7704 (N_7704,N_6478,N_6669);
nand U7705 (N_7705,N_6771,N_6133);
or U7706 (N_7706,N_6369,N_6359);
or U7707 (N_7707,N_6708,N_6992);
xnor U7708 (N_7708,N_6556,N_6537);
or U7709 (N_7709,N_6927,N_6081);
nand U7710 (N_7710,N_6767,N_6302);
xnor U7711 (N_7711,N_6772,N_6957);
nor U7712 (N_7712,N_6192,N_6852);
xor U7713 (N_7713,N_6991,N_6136);
or U7714 (N_7714,N_6201,N_6022);
xnor U7715 (N_7715,N_6843,N_6283);
xor U7716 (N_7716,N_6959,N_6618);
nand U7717 (N_7717,N_6776,N_6352);
nand U7718 (N_7718,N_6696,N_6212);
nand U7719 (N_7719,N_6350,N_6204);
nor U7720 (N_7720,N_6126,N_6426);
xor U7721 (N_7721,N_6336,N_6149);
xor U7722 (N_7722,N_6441,N_6478);
nor U7723 (N_7723,N_6324,N_6744);
and U7724 (N_7724,N_6501,N_6214);
xor U7725 (N_7725,N_6014,N_6409);
and U7726 (N_7726,N_6649,N_6401);
nand U7727 (N_7727,N_6392,N_6442);
and U7728 (N_7728,N_6322,N_6457);
or U7729 (N_7729,N_6051,N_6236);
nor U7730 (N_7730,N_6786,N_6492);
xor U7731 (N_7731,N_6527,N_6980);
nor U7732 (N_7732,N_6532,N_6216);
and U7733 (N_7733,N_6593,N_6499);
nand U7734 (N_7734,N_6306,N_6529);
and U7735 (N_7735,N_6004,N_6964);
nand U7736 (N_7736,N_6735,N_6988);
and U7737 (N_7737,N_6498,N_6982);
xor U7738 (N_7738,N_6174,N_6534);
nand U7739 (N_7739,N_6019,N_6706);
or U7740 (N_7740,N_6955,N_6425);
nor U7741 (N_7741,N_6896,N_6619);
and U7742 (N_7742,N_6093,N_6561);
or U7743 (N_7743,N_6550,N_6702);
nor U7744 (N_7744,N_6526,N_6776);
and U7745 (N_7745,N_6735,N_6244);
or U7746 (N_7746,N_6610,N_6591);
and U7747 (N_7747,N_6403,N_6575);
or U7748 (N_7748,N_6739,N_6285);
or U7749 (N_7749,N_6500,N_6811);
xnor U7750 (N_7750,N_6239,N_6739);
xor U7751 (N_7751,N_6888,N_6400);
or U7752 (N_7752,N_6964,N_6200);
nand U7753 (N_7753,N_6962,N_6058);
and U7754 (N_7754,N_6974,N_6396);
nor U7755 (N_7755,N_6540,N_6764);
nor U7756 (N_7756,N_6536,N_6329);
nor U7757 (N_7757,N_6908,N_6293);
or U7758 (N_7758,N_6535,N_6670);
nor U7759 (N_7759,N_6432,N_6482);
nor U7760 (N_7760,N_6607,N_6182);
xor U7761 (N_7761,N_6984,N_6689);
or U7762 (N_7762,N_6655,N_6853);
and U7763 (N_7763,N_6227,N_6774);
xor U7764 (N_7764,N_6552,N_6085);
and U7765 (N_7765,N_6776,N_6406);
nand U7766 (N_7766,N_6786,N_6069);
or U7767 (N_7767,N_6323,N_6028);
or U7768 (N_7768,N_6209,N_6104);
nor U7769 (N_7769,N_6075,N_6779);
nand U7770 (N_7770,N_6361,N_6503);
nand U7771 (N_7771,N_6278,N_6797);
and U7772 (N_7772,N_6748,N_6576);
xnor U7773 (N_7773,N_6555,N_6560);
nor U7774 (N_7774,N_6643,N_6546);
and U7775 (N_7775,N_6073,N_6502);
or U7776 (N_7776,N_6677,N_6584);
nor U7777 (N_7777,N_6830,N_6416);
nand U7778 (N_7778,N_6343,N_6769);
xor U7779 (N_7779,N_6527,N_6113);
nand U7780 (N_7780,N_6417,N_6875);
nor U7781 (N_7781,N_6542,N_6232);
and U7782 (N_7782,N_6587,N_6071);
or U7783 (N_7783,N_6560,N_6435);
and U7784 (N_7784,N_6329,N_6827);
nor U7785 (N_7785,N_6839,N_6697);
and U7786 (N_7786,N_6137,N_6901);
nor U7787 (N_7787,N_6841,N_6494);
or U7788 (N_7788,N_6632,N_6832);
nor U7789 (N_7789,N_6677,N_6129);
nor U7790 (N_7790,N_6016,N_6718);
xnor U7791 (N_7791,N_6611,N_6597);
xor U7792 (N_7792,N_6438,N_6136);
and U7793 (N_7793,N_6776,N_6599);
xnor U7794 (N_7794,N_6753,N_6120);
nor U7795 (N_7795,N_6314,N_6276);
xnor U7796 (N_7796,N_6692,N_6361);
xor U7797 (N_7797,N_6972,N_6690);
nor U7798 (N_7798,N_6746,N_6899);
nor U7799 (N_7799,N_6155,N_6466);
xor U7800 (N_7800,N_6750,N_6819);
nand U7801 (N_7801,N_6662,N_6890);
nor U7802 (N_7802,N_6750,N_6990);
xnor U7803 (N_7803,N_6834,N_6938);
nand U7804 (N_7804,N_6175,N_6949);
and U7805 (N_7805,N_6991,N_6241);
or U7806 (N_7806,N_6877,N_6537);
xnor U7807 (N_7807,N_6024,N_6349);
nor U7808 (N_7808,N_6625,N_6970);
xnor U7809 (N_7809,N_6643,N_6024);
nand U7810 (N_7810,N_6286,N_6378);
nor U7811 (N_7811,N_6596,N_6334);
xor U7812 (N_7812,N_6461,N_6772);
nand U7813 (N_7813,N_6611,N_6931);
or U7814 (N_7814,N_6946,N_6577);
and U7815 (N_7815,N_6394,N_6330);
or U7816 (N_7816,N_6767,N_6936);
nor U7817 (N_7817,N_6357,N_6322);
xor U7818 (N_7818,N_6553,N_6435);
nand U7819 (N_7819,N_6475,N_6627);
nor U7820 (N_7820,N_6673,N_6597);
xor U7821 (N_7821,N_6356,N_6891);
or U7822 (N_7822,N_6672,N_6057);
and U7823 (N_7823,N_6304,N_6299);
and U7824 (N_7824,N_6254,N_6385);
nor U7825 (N_7825,N_6373,N_6332);
nor U7826 (N_7826,N_6636,N_6275);
or U7827 (N_7827,N_6346,N_6669);
nor U7828 (N_7828,N_6644,N_6498);
xnor U7829 (N_7829,N_6507,N_6251);
xor U7830 (N_7830,N_6528,N_6699);
xnor U7831 (N_7831,N_6143,N_6784);
and U7832 (N_7832,N_6722,N_6142);
xor U7833 (N_7833,N_6052,N_6048);
nor U7834 (N_7834,N_6939,N_6247);
or U7835 (N_7835,N_6882,N_6646);
nand U7836 (N_7836,N_6339,N_6156);
and U7837 (N_7837,N_6916,N_6946);
xor U7838 (N_7838,N_6778,N_6252);
or U7839 (N_7839,N_6602,N_6464);
or U7840 (N_7840,N_6845,N_6429);
xnor U7841 (N_7841,N_6218,N_6389);
or U7842 (N_7842,N_6448,N_6081);
nor U7843 (N_7843,N_6586,N_6441);
xnor U7844 (N_7844,N_6258,N_6347);
and U7845 (N_7845,N_6422,N_6674);
nand U7846 (N_7846,N_6493,N_6684);
xnor U7847 (N_7847,N_6159,N_6858);
and U7848 (N_7848,N_6003,N_6125);
nor U7849 (N_7849,N_6677,N_6906);
or U7850 (N_7850,N_6294,N_6620);
nor U7851 (N_7851,N_6279,N_6457);
and U7852 (N_7852,N_6858,N_6711);
or U7853 (N_7853,N_6091,N_6548);
xnor U7854 (N_7854,N_6901,N_6473);
nand U7855 (N_7855,N_6515,N_6763);
or U7856 (N_7856,N_6836,N_6756);
and U7857 (N_7857,N_6971,N_6764);
and U7858 (N_7858,N_6541,N_6816);
nor U7859 (N_7859,N_6076,N_6001);
and U7860 (N_7860,N_6390,N_6895);
and U7861 (N_7861,N_6437,N_6383);
nor U7862 (N_7862,N_6753,N_6629);
nand U7863 (N_7863,N_6029,N_6673);
nand U7864 (N_7864,N_6424,N_6806);
nor U7865 (N_7865,N_6711,N_6105);
and U7866 (N_7866,N_6034,N_6755);
and U7867 (N_7867,N_6002,N_6918);
and U7868 (N_7868,N_6209,N_6941);
and U7869 (N_7869,N_6174,N_6496);
xor U7870 (N_7870,N_6018,N_6753);
xor U7871 (N_7871,N_6942,N_6118);
or U7872 (N_7872,N_6818,N_6329);
nand U7873 (N_7873,N_6809,N_6774);
or U7874 (N_7874,N_6177,N_6886);
xor U7875 (N_7875,N_6556,N_6700);
or U7876 (N_7876,N_6116,N_6946);
xor U7877 (N_7877,N_6904,N_6047);
nand U7878 (N_7878,N_6201,N_6814);
or U7879 (N_7879,N_6583,N_6561);
nand U7880 (N_7880,N_6756,N_6468);
nor U7881 (N_7881,N_6965,N_6173);
or U7882 (N_7882,N_6058,N_6225);
and U7883 (N_7883,N_6061,N_6345);
xnor U7884 (N_7884,N_6154,N_6005);
or U7885 (N_7885,N_6847,N_6855);
nand U7886 (N_7886,N_6768,N_6970);
nor U7887 (N_7887,N_6261,N_6922);
or U7888 (N_7888,N_6424,N_6691);
nand U7889 (N_7889,N_6445,N_6130);
and U7890 (N_7890,N_6102,N_6090);
xor U7891 (N_7891,N_6284,N_6528);
or U7892 (N_7892,N_6473,N_6264);
xnor U7893 (N_7893,N_6512,N_6631);
xnor U7894 (N_7894,N_6709,N_6611);
or U7895 (N_7895,N_6575,N_6857);
nand U7896 (N_7896,N_6667,N_6331);
or U7897 (N_7897,N_6884,N_6817);
and U7898 (N_7898,N_6546,N_6106);
nor U7899 (N_7899,N_6295,N_6170);
xor U7900 (N_7900,N_6056,N_6919);
nor U7901 (N_7901,N_6129,N_6865);
nand U7902 (N_7902,N_6444,N_6699);
or U7903 (N_7903,N_6726,N_6955);
nand U7904 (N_7904,N_6546,N_6688);
nor U7905 (N_7905,N_6105,N_6668);
nand U7906 (N_7906,N_6763,N_6185);
and U7907 (N_7907,N_6554,N_6643);
and U7908 (N_7908,N_6545,N_6785);
and U7909 (N_7909,N_6930,N_6943);
or U7910 (N_7910,N_6406,N_6381);
nand U7911 (N_7911,N_6129,N_6959);
or U7912 (N_7912,N_6056,N_6885);
xor U7913 (N_7913,N_6108,N_6903);
nor U7914 (N_7914,N_6773,N_6909);
nor U7915 (N_7915,N_6812,N_6763);
nand U7916 (N_7916,N_6189,N_6595);
or U7917 (N_7917,N_6408,N_6332);
nand U7918 (N_7918,N_6074,N_6279);
and U7919 (N_7919,N_6488,N_6905);
nand U7920 (N_7920,N_6978,N_6874);
nor U7921 (N_7921,N_6910,N_6082);
nor U7922 (N_7922,N_6958,N_6468);
nor U7923 (N_7923,N_6469,N_6365);
and U7924 (N_7924,N_6495,N_6488);
and U7925 (N_7925,N_6694,N_6131);
xor U7926 (N_7926,N_6148,N_6708);
nor U7927 (N_7927,N_6528,N_6245);
nand U7928 (N_7928,N_6573,N_6119);
xor U7929 (N_7929,N_6288,N_6652);
xnor U7930 (N_7930,N_6014,N_6494);
xnor U7931 (N_7931,N_6853,N_6083);
nand U7932 (N_7932,N_6956,N_6189);
and U7933 (N_7933,N_6847,N_6730);
or U7934 (N_7934,N_6572,N_6660);
and U7935 (N_7935,N_6706,N_6379);
nor U7936 (N_7936,N_6512,N_6541);
or U7937 (N_7937,N_6660,N_6299);
nor U7938 (N_7938,N_6474,N_6354);
xnor U7939 (N_7939,N_6756,N_6630);
or U7940 (N_7940,N_6461,N_6306);
xnor U7941 (N_7941,N_6278,N_6376);
or U7942 (N_7942,N_6017,N_6332);
nor U7943 (N_7943,N_6887,N_6177);
and U7944 (N_7944,N_6741,N_6695);
nand U7945 (N_7945,N_6813,N_6930);
xor U7946 (N_7946,N_6451,N_6515);
or U7947 (N_7947,N_6192,N_6989);
nor U7948 (N_7948,N_6344,N_6705);
nand U7949 (N_7949,N_6855,N_6235);
xor U7950 (N_7950,N_6109,N_6292);
nor U7951 (N_7951,N_6612,N_6126);
xor U7952 (N_7952,N_6885,N_6185);
or U7953 (N_7953,N_6005,N_6432);
xor U7954 (N_7954,N_6130,N_6667);
and U7955 (N_7955,N_6752,N_6821);
nand U7956 (N_7956,N_6132,N_6610);
nand U7957 (N_7957,N_6096,N_6692);
nand U7958 (N_7958,N_6256,N_6808);
nor U7959 (N_7959,N_6202,N_6882);
or U7960 (N_7960,N_6841,N_6261);
nor U7961 (N_7961,N_6058,N_6103);
nand U7962 (N_7962,N_6376,N_6899);
xnor U7963 (N_7963,N_6620,N_6717);
xnor U7964 (N_7964,N_6538,N_6547);
and U7965 (N_7965,N_6911,N_6254);
nand U7966 (N_7966,N_6884,N_6361);
or U7967 (N_7967,N_6266,N_6917);
or U7968 (N_7968,N_6086,N_6634);
xnor U7969 (N_7969,N_6549,N_6777);
and U7970 (N_7970,N_6496,N_6988);
and U7971 (N_7971,N_6686,N_6394);
nor U7972 (N_7972,N_6249,N_6029);
nand U7973 (N_7973,N_6644,N_6953);
xnor U7974 (N_7974,N_6094,N_6700);
xnor U7975 (N_7975,N_6184,N_6523);
nand U7976 (N_7976,N_6225,N_6433);
nand U7977 (N_7977,N_6086,N_6478);
nor U7978 (N_7978,N_6618,N_6380);
nand U7979 (N_7979,N_6633,N_6048);
nor U7980 (N_7980,N_6093,N_6868);
xnor U7981 (N_7981,N_6968,N_6025);
nand U7982 (N_7982,N_6467,N_6505);
nor U7983 (N_7983,N_6277,N_6113);
nor U7984 (N_7984,N_6575,N_6830);
xor U7985 (N_7985,N_6448,N_6971);
and U7986 (N_7986,N_6488,N_6629);
nand U7987 (N_7987,N_6622,N_6118);
xnor U7988 (N_7988,N_6162,N_6030);
xnor U7989 (N_7989,N_6408,N_6107);
nand U7990 (N_7990,N_6908,N_6426);
nor U7991 (N_7991,N_6259,N_6199);
nor U7992 (N_7992,N_6653,N_6828);
nand U7993 (N_7993,N_6245,N_6494);
nand U7994 (N_7994,N_6863,N_6090);
and U7995 (N_7995,N_6576,N_6059);
and U7996 (N_7996,N_6689,N_6353);
and U7997 (N_7997,N_6162,N_6195);
xnor U7998 (N_7998,N_6737,N_6406);
and U7999 (N_7999,N_6273,N_6398);
and U8000 (N_8000,N_7764,N_7392);
and U8001 (N_8001,N_7444,N_7934);
nand U8002 (N_8002,N_7199,N_7698);
nand U8003 (N_8003,N_7667,N_7747);
and U8004 (N_8004,N_7555,N_7318);
and U8005 (N_8005,N_7672,N_7928);
or U8006 (N_8006,N_7918,N_7598);
or U8007 (N_8007,N_7761,N_7235);
nand U8008 (N_8008,N_7927,N_7691);
or U8009 (N_8009,N_7684,N_7080);
or U8010 (N_8010,N_7020,N_7053);
or U8011 (N_8011,N_7673,N_7134);
xnor U8012 (N_8012,N_7690,N_7793);
xor U8013 (N_8013,N_7363,N_7527);
or U8014 (N_8014,N_7828,N_7206);
nor U8015 (N_8015,N_7827,N_7586);
or U8016 (N_8016,N_7525,N_7337);
nor U8017 (N_8017,N_7822,N_7292);
or U8018 (N_8018,N_7696,N_7172);
xnor U8019 (N_8019,N_7613,N_7681);
nor U8020 (N_8020,N_7883,N_7563);
and U8021 (N_8021,N_7678,N_7721);
or U8022 (N_8022,N_7992,N_7432);
nand U8023 (N_8023,N_7834,N_7602);
xor U8024 (N_8024,N_7773,N_7825);
nor U8025 (N_8025,N_7163,N_7802);
xor U8026 (N_8026,N_7414,N_7329);
nand U8027 (N_8027,N_7325,N_7739);
and U8028 (N_8028,N_7469,N_7521);
nand U8029 (N_8029,N_7550,N_7608);
and U8030 (N_8030,N_7127,N_7588);
nor U8031 (N_8031,N_7366,N_7383);
and U8032 (N_8032,N_7263,N_7112);
nor U8033 (N_8033,N_7736,N_7400);
and U8034 (N_8034,N_7055,N_7359);
nor U8035 (N_8035,N_7137,N_7907);
xor U8036 (N_8036,N_7259,N_7767);
nand U8037 (N_8037,N_7955,N_7141);
nor U8038 (N_8038,N_7836,N_7451);
or U8039 (N_8039,N_7166,N_7906);
or U8040 (N_8040,N_7566,N_7036);
xnor U8041 (N_8041,N_7858,N_7242);
xor U8042 (N_8042,N_7880,N_7872);
nor U8043 (N_8043,N_7958,N_7731);
nand U8044 (N_8044,N_7984,N_7887);
nand U8045 (N_8045,N_7157,N_7323);
or U8046 (N_8046,N_7751,N_7252);
and U8047 (N_8047,N_7682,N_7531);
or U8048 (N_8048,N_7974,N_7683);
and U8049 (N_8049,N_7445,N_7636);
and U8050 (N_8050,N_7776,N_7993);
xnor U8051 (N_8051,N_7096,N_7968);
or U8052 (N_8052,N_7786,N_7988);
or U8053 (N_8053,N_7101,N_7475);
or U8054 (N_8054,N_7393,N_7851);
or U8055 (N_8055,N_7479,N_7915);
and U8056 (N_8056,N_7911,N_7717);
xor U8057 (N_8057,N_7500,N_7312);
nand U8058 (N_8058,N_7897,N_7399);
nor U8059 (N_8059,N_7877,N_7526);
and U8060 (N_8060,N_7917,N_7591);
nand U8061 (N_8061,N_7117,N_7255);
or U8062 (N_8062,N_7882,N_7311);
xnor U8063 (N_8063,N_7440,N_7631);
or U8064 (N_8064,N_7256,N_7351);
nor U8065 (N_8065,N_7951,N_7846);
and U8066 (N_8066,N_7943,N_7221);
and U8067 (N_8067,N_7493,N_7219);
or U8068 (N_8068,N_7027,N_7619);
xnor U8069 (N_8069,N_7743,N_7549);
xor U8070 (N_8070,N_7187,N_7540);
or U8071 (N_8071,N_7963,N_7015);
nand U8072 (N_8072,N_7775,N_7412);
nor U8073 (N_8073,N_7413,N_7178);
and U8074 (N_8074,N_7946,N_7277);
nor U8075 (N_8075,N_7810,N_7954);
nand U8076 (N_8076,N_7538,N_7085);
nand U8077 (N_8077,N_7823,N_7406);
nand U8078 (N_8078,N_7726,N_7885);
xor U8079 (N_8079,N_7929,N_7148);
or U8080 (N_8080,N_7948,N_7049);
and U8081 (N_8081,N_7111,N_7090);
nand U8082 (N_8082,N_7931,N_7102);
and U8083 (N_8083,N_7364,N_7048);
or U8084 (N_8084,N_7668,N_7059);
xnor U8085 (N_8085,N_7654,N_7628);
nand U8086 (N_8086,N_7795,N_7489);
and U8087 (N_8087,N_7468,N_7223);
or U8088 (N_8088,N_7863,N_7923);
or U8089 (N_8089,N_7217,N_7518);
xnor U8090 (N_8090,N_7706,N_7944);
and U8091 (N_8091,N_7068,N_7817);
xor U8092 (N_8092,N_7287,N_7142);
nand U8093 (N_8093,N_7675,N_7788);
and U8094 (N_8094,N_7818,N_7353);
or U8095 (N_8095,N_7711,N_7530);
nand U8096 (N_8096,N_7548,N_7921);
or U8097 (N_8097,N_7657,N_7703);
nand U8098 (N_8098,N_7727,N_7511);
or U8099 (N_8099,N_7322,N_7630);
and U8100 (N_8100,N_7030,N_7964);
nand U8101 (N_8101,N_7966,N_7644);
nand U8102 (N_8102,N_7539,N_7006);
or U8103 (N_8103,N_7575,N_7088);
xor U8104 (N_8104,N_7275,N_7170);
xor U8105 (N_8105,N_7331,N_7996);
nor U8106 (N_8106,N_7926,N_7434);
xor U8107 (N_8107,N_7179,N_7517);
nor U8108 (N_8108,N_7756,N_7597);
nand U8109 (N_8109,N_7758,N_7460);
and U8110 (N_8110,N_7182,N_7590);
nand U8111 (N_8111,N_7332,N_7176);
xnor U8112 (N_8112,N_7640,N_7976);
nor U8113 (N_8113,N_7431,N_7159);
nand U8114 (N_8114,N_7635,N_7940);
and U8115 (N_8115,N_7949,N_7158);
or U8116 (N_8116,N_7384,N_7483);
nand U8117 (N_8117,N_7796,N_7089);
or U8118 (N_8118,N_7319,N_7086);
nand U8119 (N_8119,N_7896,N_7745);
nand U8120 (N_8120,N_7553,N_7599);
nand U8121 (N_8121,N_7288,N_7133);
nor U8122 (N_8122,N_7038,N_7082);
nor U8123 (N_8123,N_7411,N_7961);
nand U8124 (N_8124,N_7019,N_7272);
nor U8125 (N_8125,N_7809,N_7371);
and U8126 (N_8126,N_7340,N_7334);
nand U8127 (N_8127,N_7234,N_7123);
nand U8128 (N_8128,N_7407,N_7894);
or U8129 (N_8129,N_7355,N_7589);
nor U8130 (N_8130,N_7680,N_7699);
xnor U8131 (N_8131,N_7103,N_7890);
nand U8132 (N_8132,N_7120,N_7935);
xnor U8133 (N_8133,N_7001,N_7495);
or U8134 (N_8134,N_7404,N_7965);
nand U8135 (N_8135,N_7016,N_7249);
xor U8136 (N_8136,N_7789,N_7670);
nand U8137 (N_8137,N_7336,N_7342);
xnor U8138 (N_8138,N_7033,N_7728);
and U8139 (N_8139,N_7343,N_7939);
and U8140 (N_8140,N_7648,N_7983);
xor U8141 (N_8141,N_7128,N_7637);
or U8142 (N_8142,N_7290,N_7744);
or U8143 (N_8143,N_7838,N_7945);
nand U8144 (N_8144,N_7310,N_7580);
xnor U8145 (N_8145,N_7456,N_7614);
and U8146 (N_8146,N_7567,N_7389);
or U8147 (N_8147,N_7953,N_7752);
nor U8148 (N_8148,N_7546,N_7909);
and U8149 (N_8149,N_7194,N_7625);
xnor U8150 (N_8150,N_7876,N_7046);
or U8151 (N_8151,N_7615,N_7778);
nand U8152 (N_8152,N_7829,N_7688);
and U8153 (N_8153,N_7121,N_7729);
or U8154 (N_8154,N_7346,N_7480);
and U8155 (N_8155,N_7065,N_7695);
and U8156 (N_8156,N_7233,N_7045);
nor U8157 (N_8157,N_7448,N_7064);
xnor U8158 (N_8158,N_7800,N_7427);
or U8159 (N_8159,N_7607,N_7126);
nand U8160 (N_8160,N_7874,N_7405);
nor U8161 (N_8161,N_7076,N_7560);
or U8162 (N_8162,N_7306,N_7627);
or U8163 (N_8163,N_7236,N_7373);
xor U8164 (N_8164,N_7150,N_7308);
nor U8165 (N_8165,N_7522,N_7058);
and U8166 (N_8166,N_7886,N_7060);
xnor U8167 (N_8167,N_7095,N_7136);
xnor U8168 (N_8168,N_7110,N_7017);
and U8169 (N_8169,N_7160,N_7061);
or U8170 (N_8170,N_7294,N_7193);
and U8171 (N_8171,N_7975,N_7532);
and U8172 (N_8172,N_7956,N_7330);
and U8173 (N_8173,N_7050,N_7647);
or U8174 (N_8174,N_7618,N_7768);
or U8175 (N_8175,N_7018,N_7642);
xor U8176 (N_8176,N_7506,N_7140);
nand U8177 (N_8177,N_7477,N_7665);
nor U8178 (N_8178,N_7645,N_7171);
and U8179 (N_8179,N_7488,N_7299);
nor U8180 (N_8180,N_7115,N_7771);
and U8181 (N_8181,N_7261,N_7307);
and U8182 (N_8182,N_7716,N_7908);
xnor U8183 (N_8183,N_7669,N_7621);
xor U8184 (N_8184,N_7382,N_7568);
or U8185 (N_8185,N_7715,N_7960);
and U8186 (N_8186,N_7655,N_7420);
and U8187 (N_8187,N_7660,N_7938);
and U8188 (N_8188,N_7562,N_7295);
nand U8189 (N_8189,N_7347,N_7433);
xnor U8190 (N_8190,N_7849,N_7189);
and U8191 (N_8191,N_7520,N_7959);
nand U8192 (N_8192,N_7408,N_7650);
nand U8193 (N_8193,N_7844,N_7692);
nor U8194 (N_8194,N_7097,N_7930);
nand U8195 (N_8195,N_7357,N_7978);
or U8196 (N_8196,N_7035,N_7398);
xnor U8197 (N_8197,N_7561,N_7358);
nand U8198 (N_8198,N_7165,N_7063);
or U8199 (N_8199,N_7501,N_7071);
or U8200 (N_8200,N_7824,N_7008);
or U8201 (N_8201,N_7418,N_7842);
nor U8202 (N_8202,N_7785,N_7354);
nor U8203 (N_8203,N_7376,N_7565);
xor U8204 (N_8204,N_7671,N_7865);
nor U8205 (N_8205,N_7899,N_7226);
xnor U8206 (N_8206,N_7903,N_7177);
or U8207 (N_8207,N_7545,N_7798);
and U8208 (N_8208,N_7596,N_7733);
nor U8209 (N_8209,N_7296,N_7845);
or U8210 (N_8210,N_7062,N_7072);
nor U8211 (N_8211,N_7230,N_7113);
nand U8212 (N_8212,N_7465,N_7719);
or U8213 (N_8213,N_7679,N_7026);
or U8214 (N_8214,N_7856,N_7155);
nand U8215 (N_8215,N_7864,N_7144);
nor U8216 (N_8216,N_7470,N_7689);
or U8217 (N_8217,N_7327,N_7649);
xnor U8218 (N_8218,N_7813,N_7740);
nand U8219 (N_8219,N_7381,N_7286);
nor U8220 (N_8220,N_7714,N_7854);
or U8221 (N_8221,N_7457,N_7153);
or U8222 (N_8222,N_7855,N_7471);
xnor U8223 (N_8223,N_7205,N_7264);
nand U8224 (N_8224,N_7125,N_7762);
and U8225 (N_8225,N_7443,N_7742);
or U8226 (N_8226,N_7447,N_7730);
nand U8227 (N_8227,N_7629,N_7620);
xor U8228 (N_8228,N_7138,N_7032);
xor U8229 (N_8229,N_7852,N_7499);
nor U8230 (N_8230,N_7034,N_7007);
or U8231 (N_8231,N_7051,N_7662);
or U8232 (N_8232,N_7587,N_7116);
xor U8233 (N_8233,N_7884,N_7476);
or U8234 (N_8234,N_7485,N_7833);
nor U8235 (N_8235,N_7512,N_7749);
or U8236 (N_8236,N_7375,N_7542);
xnor U8237 (N_8237,N_7603,N_7461);
nand U8238 (N_8238,N_7084,N_7238);
or U8239 (N_8239,N_7666,N_7794);
and U8240 (N_8240,N_7013,N_7969);
and U8241 (N_8241,N_7857,N_7821);
xor U8242 (N_8242,N_7578,N_7674);
xor U8243 (N_8243,N_7986,N_7350);
nor U8244 (N_8244,N_7388,N_7701);
xor U8245 (N_8245,N_7718,N_7487);
and U8246 (N_8246,N_7022,N_7188);
or U8247 (N_8247,N_7245,N_7801);
nor U8248 (N_8248,N_7409,N_7947);
nor U8249 (N_8249,N_7191,N_7284);
and U8250 (N_8250,N_7772,N_7643);
nor U8251 (N_8251,N_7991,N_7878);
and U8252 (N_8252,N_7901,N_7780);
xnor U8253 (N_8253,N_7228,N_7247);
xnor U8254 (N_8254,N_7551,N_7231);
nand U8255 (N_8255,N_7811,N_7871);
and U8256 (N_8256,N_7012,N_7380);
and U8257 (N_8257,N_7514,N_7920);
nand U8258 (N_8258,N_7401,N_7812);
nor U8259 (N_8259,N_7156,N_7362);
or U8260 (N_8260,N_7174,N_7616);
nand U8261 (N_8261,N_7604,N_7895);
xor U8262 (N_8262,N_7724,N_7516);
xor U8263 (N_8263,N_7529,N_7029);
nand U8264 (N_8264,N_7419,N_7543);
or U8265 (N_8265,N_7341,N_7459);
nor U8266 (N_8266,N_7151,N_7087);
or U8267 (N_8267,N_7003,N_7748);
and U8268 (N_8268,N_7685,N_7732);
and U8269 (N_8269,N_7079,N_7303);
or U8270 (N_8270,N_7094,N_7130);
nand U8271 (N_8271,N_7365,N_7011);
nand U8272 (N_8272,N_7709,N_7273);
xnor U8273 (N_8273,N_7344,N_7198);
nor U8274 (N_8274,N_7486,N_7766);
xor U8275 (N_8275,N_7820,N_7004);
and U8276 (N_8276,N_7651,N_7293);
nand U8277 (N_8277,N_7462,N_7270);
and U8278 (N_8278,N_7300,N_7202);
xnor U8279 (N_8279,N_7056,N_7175);
nand U8280 (N_8280,N_7279,N_7262);
nand U8281 (N_8281,N_7970,N_7547);
and U8282 (N_8282,N_7237,N_7143);
and U8283 (N_8283,N_7367,N_7124);
nor U8284 (N_8284,N_7266,N_7893);
and U8285 (N_8285,N_7652,N_7843);
nor U8286 (N_8286,N_7466,N_7131);
and U8287 (N_8287,N_7850,N_7735);
nor U8288 (N_8288,N_7712,N_7980);
xor U8289 (N_8289,N_7898,N_7149);
and U8290 (N_8290,N_7995,N_7866);
nand U8291 (N_8291,N_7807,N_7421);
xor U8292 (N_8292,N_7360,N_7098);
or U8293 (N_8293,N_7066,N_7967);
or U8294 (N_8294,N_7656,N_7464);
nand U8295 (N_8295,N_7556,N_7145);
and U8296 (N_8296,N_7478,N_7889);
xnor U8297 (N_8297,N_7267,N_7356);
xor U8298 (N_8298,N_7119,N_7248);
and U8299 (N_8299,N_7397,N_7722);
or U8300 (N_8300,N_7214,N_7246);
nand U8301 (N_8301,N_7338,N_7663);
nand U8302 (N_8302,N_7624,N_7559);
or U8303 (N_8303,N_7738,N_7741);
nand U8304 (N_8304,N_7515,N_7472);
nor U8305 (N_8305,N_7301,N_7862);
or U8306 (N_8306,N_7403,N_7760);
and U8307 (N_8307,N_7067,N_7564);
or U8308 (N_8308,N_7859,N_7075);
nor U8309 (N_8309,N_7435,N_7200);
or U8310 (N_8310,N_7369,N_7777);
nand U8311 (N_8311,N_7541,N_7250);
nand U8312 (N_8312,N_7240,N_7936);
xnor U8313 (N_8313,N_7534,N_7888);
xnor U8314 (N_8314,N_7998,N_7315);
xor U8315 (N_8315,N_7808,N_7806);
and U8316 (N_8316,N_7378,N_7557);
and U8317 (N_8317,N_7320,N_7490);
nor U8318 (N_8318,N_7819,N_7875);
or U8319 (N_8319,N_7291,N_7450);
and U8320 (N_8320,N_7326,N_7167);
nor U8321 (N_8321,N_7289,N_7870);
nor U8322 (N_8322,N_7083,N_7028);
or U8323 (N_8323,N_7841,N_7932);
nor U8324 (N_8324,N_7154,N_7641);
and U8325 (N_8325,N_7664,N_7129);
and U8326 (N_8326,N_7169,N_7423);
nor U8327 (N_8327,N_7227,N_7181);
nand U8328 (N_8328,N_7316,N_7609);
nand U8329 (N_8329,N_7574,N_7429);
nor U8330 (N_8330,N_7276,N_7892);
nand U8331 (N_8331,N_7577,N_7804);
nand U8332 (N_8332,N_7700,N_7044);
and U8333 (N_8333,N_7611,N_7508);
and U8334 (N_8334,N_7633,N_7328);
xnor U8335 (N_8335,N_7147,N_7239);
nand U8336 (N_8336,N_7391,N_7282);
xnor U8337 (N_8337,N_7746,N_7774);
or U8338 (N_8338,N_7987,N_7910);
nor U8339 (N_8339,N_7251,N_7192);
nand U8340 (N_8340,N_7676,N_7737);
nand U8341 (N_8341,N_7552,N_7449);
xor U8342 (N_8342,N_7606,N_7639);
or U8343 (N_8343,N_7070,N_7211);
or U8344 (N_8344,N_7659,N_7254);
nor U8345 (N_8345,N_7533,N_7913);
nor U8346 (N_8346,N_7152,N_7268);
and U8347 (N_8347,N_7074,N_7704);
or U8348 (N_8348,N_7207,N_7904);
or U8349 (N_8349,N_7430,N_7973);
nor U8350 (N_8350,N_7581,N_7569);
or U8351 (N_8351,N_7395,N_7041);
nand U8352 (N_8352,N_7994,N_7723);
nand U8353 (N_8353,N_7610,N_7304);
or U8354 (N_8354,N_7280,N_7091);
nor U8355 (N_8355,N_7314,N_7941);
and U8356 (N_8356,N_7962,N_7720);
and U8357 (N_8357,N_7694,N_7232);
and U8358 (N_8358,N_7769,N_7057);
nand U8359 (N_8359,N_7024,N_7209);
xor U8360 (N_8360,N_7990,N_7180);
or U8361 (N_8361,N_7831,N_7585);
or U8362 (N_8362,N_7805,N_7396);
xor U8363 (N_8363,N_7753,N_7507);
nor U8364 (N_8364,N_7919,N_7426);
and U8365 (N_8365,N_7523,N_7916);
or U8366 (N_8366,N_7368,N_7139);
and U8367 (N_8367,N_7162,N_7370);
xor U8368 (N_8368,N_7297,N_7950);
or U8369 (N_8369,N_7830,N_7069);
and U8370 (N_8370,N_7705,N_7377);
nand U8371 (N_8371,N_7224,N_7099);
or U8372 (N_8372,N_7754,N_7781);
nand U8373 (N_8373,N_7687,N_7661);
nor U8374 (N_8374,N_7891,N_7416);
and U8375 (N_8375,N_7867,N_7815);
nor U8376 (N_8376,N_7385,N_7442);
nand U8377 (N_8377,N_7361,N_7484);
and U8378 (N_8378,N_7535,N_7047);
or U8379 (N_8379,N_7977,N_7260);
or U8380 (N_8380,N_7554,N_7708);
nand U8381 (N_8381,N_7054,N_7455);
xnor U8382 (N_8382,N_7037,N_7173);
xnor U8383 (N_8383,N_7313,N_7881);
or U8384 (N_8384,N_7100,N_7321);
nor U8385 (N_8385,N_7039,N_7702);
or U8386 (N_8386,N_7164,N_7437);
nand U8387 (N_8387,N_7971,N_7879);
xnor U8388 (N_8388,N_7503,N_7757);
nand U8389 (N_8389,N_7600,N_7190);
and U8390 (N_8390,N_7784,N_7135);
nand U8391 (N_8391,N_7213,N_7040);
xor U8392 (N_8392,N_7186,N_7677);
nand U8393 (N_8393,N_7439,N_7942);
nor U8394 (N_8394,N_7622,N_7799);
nand U8395 (N_8395,N_7595,N_7241);
xor U8396 (N_8396,N_7106,N_7372);
nand U8397 (N_8397,N_7184,N_7697);
nand U8398 (N_8398,N_7118,N_7623);
nor U8399 (N_8399,N_7504,N_7146);
or U8400 (N_8400,N_7519,N_7424);
nor U8401 (N_8401,N_7782,N_7474);
nand U8402 (N_8402,N_7105,N_7210);
and U8403 (N_8403,N_7271,N_7298);
xnor U8404 (N_8404,N_7952,N_7002);
nand U8405 (N_8405,N_7605,N_7925);
and U8406 (N_8406,N_7285,N_7573);
nand U8407 (N_8407,N_7463,N_7212);
or U8408 (N_8408,N_7482,N_7803);
nor U8409 (N_8409,N_7216,N_7905);
xnor U8410 (N_8410,N_7014,N_7114);
and U8411 (N_8411,N_7626,N_7203);
or U8412 (N_8412,N_7632,N_7853);
and U8413 (N_8413,N_7265,N_7195);
and U8414 (N_8414,N_7571,N_7997);
nor U8415 (N_8415,N_7122,N_7755);
nand U8416 (N_8416,N_7208,N_7052);
or U8417 (N_8417,N_7073,N_7093);
and U8418 (N_8418,N_7107,N_7257);
nor U8419 (N_8419,N_7646,N_7594);
nand U8420 (N_8420,N_7196,N_7021);
or U8421 (N_8421,N_7713,N_7601);
and U8422 (N_8422,N_7814,N_7860);
nor U8423 (N_8423,N_7902,N_7912);
and U8424 (N_8424,N_7394,N_7985);
nor U8425 (N_8425,N_7494,N_7078);
or U8426 (N_8426,N_7937,N_7510);
xnor U8427 (N_8427,N_7787,N_7658);
nor U8428 (N_8428,N_7779,N_7417);
or U8429 (N_8429,N_7583,N_7274);
nand U8430 (N_8430,N_7108,N_7707);
or U8431 (N_8431,N_7592,N_7422);
nor U8432 (N_8432,N_7317,N_7759);
nand U8433 (N_8433,N_7900,N_7345);
and U8434 (N_8434,N_7348,N_7023);
xnor U8435 (N_8435,N_7979,N_7243);
or U8436 (N_8436,N_7000,N_7335);
xnor U8437 (N_8437,N_7302,N_7957);
xor U8438 (N_8438,N_7305,N_7570);
nand U8439 (N_8439,N_7081,N_7349);
nor U8440 (N_8440,N_7458,N_7379);
nor U8441 (N_8441,N_7505,N_7109);
xor U8442 (N_8442,N_7835,N_7765);
and U8443 (N_8443,N_7869,N_7868);
xor U8444 (N_8444,N_7933,N_7092);
or U8445 (N_8445,N_7582,N_7497);
nor U8446 (N_8446,N_7792,N_7763);
nand U8447 (N_8447,N_7425,N_7922);
or U8448 (N_8448,N_7847,N_7491);
and U8449 (N_8449,N_7324,N_7509);
nand U8450 (N_8450,N_7839,N_7593);
xor U8451 (N_8451,N_7686,N_7537);
xor U8452 (N_8452,N_7132,N_7387);
nand U8453 (N_8453,N_7498,N_7873);
nor U8454 (N_8454,N_7197,N_7402);
nand U8455 (N_8455,N_7244,N_7168);
and U8456 (N_8456,N_7576,N_7797);
and U8457 (N_8457,N_7215,N_7333);
or U8458 (N_8458,N_7225,N_7258);
nand U8459 (N_8459,N_7734,N_7579);
or U8460 (N_8460,N_7832,N_7278);
and U8461 (N_8461,N_7077,N_7031);
and U8462 (N_8462,N_7185,N_7220);
and U8463 (N_8463,N_7861,N_7837);
xnor U8464 (N_8464,N_7269,N_7229);
or U8465 (N_8465,N_7467,N_7410);
or U8466 (N_8466,N_7513,N_7783);
xor U8467 (N_8467,N_7452,N_7386);
nand U8468 (N_8468,N_7638,N_7204);
nand U8469 (N_8469,N_7816,N_7283);
or U8470 (N_8470,N_7253,N_7473);
and U8471 (N_8471,N_7428,N_7981);
xor U8472 (N_8472,N_7972,N_7339);
and U8473 (N_8473,N_7710,N_7536);
or U8474 (N_8474,N_7791,N_7982);
xor U8475 (N_8475,N_7989,N_7572);
xor U8476 (N_8476,N_7161,N_7558);
nand U8477 (N_8477,N_7914,N_7104);
and U8478 (N_8478,N_7009,N_7826);
or U8479 (N_8479,N_7725,N_7446);
xor U8480 (N_8480,N_7848,N_7281);
nand U8481 (N_8481,N_7453,N_7352);
xnor U8482 (N_8482,N_7043,N_7502);
xnor U8483 (N_8483,N_7201,N_7617);
nand U8484 (N_8484,N_7770,N_7924);
nand U8485 (N_8485,N_7309,N_7222);
nand U8486 (N_8486,N_7840,N_7492);
or U8487 (N_8487,N_7436,N_7693);
or U8488 (N_8488,N_7528,N_7025);
nor U8489 (N_8489,N_7374,N_7544);
nor U8490 (N_8490,N_7481,N_7612);
or U8491 (N_8491,N_7441,N_7999);
xor U8492 (N_8492,N_7390,N_7042);
nand U8493 (N_8493,N_7438,N_7524);
xnor U8494 (N_8494,N_7634,N_7218);
nor U8495 (N_8495,N_7653,N_7584);
or U8496 (N_8496,N_7496,N_7454);
or U8497 (N_8497,N_7183,N_7005);
and U8498 (N_8498,N_7415,N_7790);
xnor U8499 (N_8499,N_7010,N_7750);
or U8500 (N_8500,N_7293,N_7592);
xnor U8501 (N_8501,N_7281,N_7808);
xnor U8502 (N_8502,N_7776,N_7812);
nand U8503 (N_8503,N_7085,N_7677);
xor U8504 (N_8504,N_7731,N_7566);
or U8505 (N_8505,N_7189,N_7021);
nand U8506 (N_8506,N_7094,N_7150);
xnor U8507 (N_8507,N_7914,N_7557);
nand U8508 (N_8508,N_7964,N_7273);
nand U8509 (N_8509,N_7787,N_7909);
nand U8510 (N_8510,N_7799,N_7426);
xor U8511 (N_8511,N_7115,N_7076);
nor U8512 (N_8512,N_7161,N_7922);
nand U8513 (N_8513,N_7361,N_7301);
and U8514 (N_8514,N_7709,N_7081);
or U8515 (N_8515,N_7059,N_7831);
and U8516 (N_8516,N_7572,N_7715);
and U8517 (N_8517,N_7888,N_7599);
nand U8518 (N_8518,N_7831,N_7247);
and U8519 (N_8519,N_7814,N_7379);
xor U8520 (N_8520,N_7109,N_7154);
xnor U8521 (N_8521,N_7484,N_7134);
xnor U8522 (N_8522,N_7183,N_7981);
and U8523 (N_8523,N_7818,N_7601);
and U8524 (N_8524,N_7098,N_7722);
nand U8525 (N_8525,N_7108,N_7741);
nor U8526 (N_8526,N_7992,N_7986);
or U8527 (N_8527,N_7106,N_7236);
and U8528 (N_8528,N_7229,N_7257);
nor U8529 (N_8529,N_7833,N_7968);
and U8530 (N_8530,N_7226,N_7229);
and U8531 (N_8531,N_7191,N_7114);
nor U8532 (N_8532,N_7596,N_7598);
xor U8533 (N_8533,N_7624,N_7727);
or U8534 (N_8534,N_7597,N_7901);
nor U8535 (N_8535,N_7810,N_7632);
or U8536 (N_8536,N_7016,N_7107);
nor U8537 (N_8537,N_7412,N_7780);
nor U8538 (N_8538,N_7654,N_7184);
or U8539 (N_8539,N_7000,N_7946);
nand U8540 (N_8540,N_7346,N_7460);
nor U8541 (N_8541,N_7813,N_7880);
nand U8542 (N_8542,N_7210,N_7332);
or U8543 (N_8543,N_7967,N_7830);
and U8544 (N_8544,N_7634,N_7853);
or U8545 (N_8545,N_7694,N_7384);
nor U8546 (N_8546,N_7054,N_7338);
nor U8547 (N_8547,N_7803,N_7855);
xnor U8548 (N_8548,N_7671,N_7539);
nor U8549 (N_8549,N_7802,N_7430);
nor U8550 (N_8550,N_7273,N_7859);
or U8551 (N_8551,N_7490,N_7884);
xor U8552 (N_8552,N_7023,N_7435);
and U8553 (N_8553,N_7658,N_7833);
or U8554 (N_8554,N_7399,N_7719);
xnor U8555 (N_8555,N_7260,N_7619);
nand U8556 (N_8556,N_7994,N_7812);
nand U8557 (N_8557,N_7420,N_7208);
nor U8558 (N_8558,N_7457,N_7354);
xor U8559 (N_8559,N_7054,N_7918);
and U8560 (N_8560,N_7927,N_7363);
nor U8561 (N_8561,N_7905,N_7558);
nand U8562 (N_8562,N_7188,N_7254);
xor U8563 (N_8563,N_7888,N_7086);
or U8564 (N_8564,N_7196,N_7912);
nand U8565 (N_8565,N_7949,N_7656);
xor U8566 (N_8566,N_7004,N_7554);
or U8567 (N_8567,N_7400,N_7854);
nand U8568 (N_8568,N_7050,N_7428);
or U8569 (N_8569,N_7049,N_7988);
xor U8570 (N_8570,N_7597,N_7070);
and U8571 (N_8571,N_7631,N_7697);
nand U8572 (N_8572,N_7656,N_7045);
xor U8573 (N_8573,N_7344,N_7881);
xor U8574 (N_8574,N_7261,N_7524);
nor U8575 (N_8575,N_7577,N_7700);
xnor U8576 (N_8576,N_7063,N_7089);
and U8577 (N_8577,N_7191,N_7480);
xnor U8578 (N_8578,N_7631,N_7722);
or U8579 (N_8579,N_7914,N_7001);
or U8580 (N_8580,N_7619,N_7153);
or U8581 (N_8581,N_7108,N_7891);
or U8582 (N_8582,N_7751,N_7965);
and U8583 (N_8583,N_7337,N_7507);
xnor U8584 (N_8584,N_7291,N_7834);
and U8585 (N_8585,N_7401,N_7356);
nor U8586 (N_8586,N_7600,N_7841);
nor U8587 (N_8587,N_7939,N_7602);
nor U8588 (N_8588,N_7868,N_7821);
xor U8589 (N_8589,N_7342,N_7206);
or U8590 (N_8590,N_7605,N_7568);
xnor U8591 (N_8591,N_7116,N_7991);
or U8592 (N_8592,N_7406,N_7968);
nor U8593 (N_8593,N_7667,N_7555);
nand U8594 (N_8594,N_7709,N_7008);
or U8595 (N_8595,N_7585,N_7770);
nor U8596 (N_8596,N_7984,N_7379);
or U8597 (N_8597,N_7666,N_7700);
and U8598 (N_8598,N_7732,N_7739);
nor U8599 (N_8599,N_7513,N_7390);
or U8600 (N_8600,N_7510,N_7333);
nor U8601 (N_8601,N_7132,N_7233);
nor U8602 (N_8602,N_7272,N_7132);
xnor U8603 (N_8603,N_7886,N_7926);
and U8604 (N_8604,N_7799,N_7924);
xor U8605 (N_8605,N_7312,N_7655);
nor U8606 (N_8606,N_7428,N_7729);
xor U8607 (N_8607,N_7718,N_7924);
and U8608 (N_8608,N_7517,N_7266);
nor U8609 (N_8609,N_7037,N_7096);
or U8610 (N_8610,N_7436,N_7612);
xor U8611 (N_8611,N_7857,N_7188);
nand U8612 (N_8612,N_7009,N_7300);
and U8613 (N_8613,N_7197,N_7430);
or U8614 (N_8614,N_7518,N_7886);
or U8615 (N_8615,N_7403,N_7972);
xnor U8616 (N_8616,N_7687,N_7916);
nand U8617 (N_8617,N_7037,N_7565);
nor U8618 (N_8618,N_7289,N_7118);
or U8619 (N_8619,N_7642,N_7007);
xnor U8620 (N_8620,N_7890,N_7910);
nand U8621 (N_8621,N_7382,N_7071);
and U8622 (N_8622,N_7542,N_7337);
nor U8623 (N_8623,N_7515,N_7345);
and U8624 (N_8624,N_7623,N_7387);
xor U8625 (N_8625,N_7651,N_7171);
or U8626 (N_8626,N_7579,N_7218);
nand U8627 (N_8627,N_7856,N_7628);
or U8628 (N_8628,N_7052,N_7330);
nand U8629 (N_8629,N_7209,N_7661);
or U8630 (N_8630,N_7385,N_7523);
and U8631 (N_8631,N_7519,N_7347);
nand U8632 (N_8632,N_7271,N_7207);
and U8633 (N_8633,N_7783,N_7084);
nor U8634 (N_8634,N_7052,N_7594);
or U8635 (N_8635,N_7306,N_7677);
nor U8636 (N_8636,N_7718,N_7810);
xnor U8637 (N_8637,N_7760,N_7015);
and U8638 (N_8638,N_7264,N_7521);
xor U8639 (N_8639,N_7145,N_7577);
and U8640 (N_8640,N_7551,N_7953);
and U8641 (N_8641,N_7782,N_7459);
nand U8642 (N_8642,N_7640,N_7255);
nor U8643 (N_8643,N_7141,N_7540);
xnor U8644 (N_8644,N_7381,N_7586);
nand U8645 (N_8645,N_7827,N_7690);
nand U8646 (N_8646,N_7760,N_7632);
nor U8647 (N_8647,N_7822,N_7415);
nand U8648 (N_8648,N_7842,N_7911);
nor U8649 (N_8649,N_7967,N_7615);
and U8650 (N_8650,N_7571,N_7204);
nor U8651 (N_8651,N_7614,N_7450);
nor U8652 (N_8652,N_7504,N_7479);
nand U8653 (N_8653,N_7532,N_7887);
xnor U8654 (N_8654,N_7349,N_7003);
or U8655 (N_8655,N_7634,N_7855);
nor U8656 (N_8656,N_7115,N_7250);
and U8657 (N_8657,N_7354,N_7430);
and U8658 (N_8658,N_7048,N_7677);
and U8659 (N_8659,N_7582,N_7984);
xnor U8660 (N_8660,N_7640,N_7211);
nand U8661 (N_8661,N_7524,N_7626);
nand U8662 (N_8662,N_7287,N_7626);
and U8663 (N_8663,N_7991,N_7671);
nor U8664 (N_8664,N_7809,N_7364);
nor U8665 (N_8665,N_7875,N_7110);
and U8666 (N_8666,N_7833,N_7634);
nor U8667 (N_8667,N_7386,N_7936);
nand U8668 (N_8668,N_7793,N_7321);
nor U8669 (N_8669,N_7493,N_7698);
xor U8670 (N_8670,N_7335,N_7430);
or U8671 (N_8671,N_7550,N_7835);
and U8672 (N_8672,N_7458,N_7555);
or U8673 (N_8673,N_7620,N_7638);
and U8674 (N_8674,N_7280,N_7262);
or U8675 (N_8675,N_7316,N_7635);
nand U8676 (N_8676,N_7069,N_7567);
nor U8677 (N_8677,N_7746,N_7976);
xnor U8678 (N_8678,N_7241,N_7037);
nand U8679 (N_8679,N_7832,N_7055);
and U8680 (N_8680,N_7475,N_7360);
xor U8681 (N_8681,N_7168,N_7508);
or U8682 (N_8682,N_7011,N_7672);
xor U8683 (N_8683,N_7640,N_7905);
and U8684 (N_8684,N_7986,N_7416);
nand U8685 (N_8685,N_7468,N_7277);
xor U8686 (N_8686,N_7079,N_7213);
xor U8687 (N_8687,N_7929,N_7123);
xnor U8688 (N_8688,N_7890,N_7323);
and U8689 (N_8689,N_7121,N_7537);
nand U8690 (N_8690,N_7027,N_7217);
xor U8691 (N_8691,N_7820,N_7407);
and U8692 (N_8692,N_7083,N_7322);
or U8693 (N_8693,N_7126,N_7560);
nand U8694 (N_8694,N_7887,N_7518);
or U8695 (N_8695,N_7718,N_7537);
xnor U8696 (N_8696,N_7483,N_7980);
nor U8697 (N_8697,N_7782,N_7413);
or U8698 (N_8698,N_7397,N_7449);
xnor U8699 (N_8699,N_7241,N_7390);
or U8700 (N_8700,N_7828,N_7591);
nor U8701 (N_8701,N_7194,N_7638);
nor U8702 (N_8702,N_7742,N_7946);
xor U8703 (N_8703,N_7786,N_7284);
or U8704 (N_8704,N_7069,N_7598);
xor U8705 (N_8705,N_7873,N_7172);
and U8706 (N_8706,N_7925,N_7274);
nor U8707 (N_8707,N_7251,N_7214);
xnor U8708 (N_8708,N_7937,N_7217);
and U8709 (N_8709,N_7915,N_7121);
or U8710 (N_8710,N_7555,N_7545);
or U8711 (N_8711,N_7904,N_7537);
nor U8712 (N_8712,N_7270,N_7563);
xor U8713 (N_8713,N_7313,N_7269);
nor U8714 (N_8714,N_7845,N_7813);
nor U8715 (N_8715,N_7226,N_7241);
xnor U8716 (N_8716,N_7643,N_7238);
or U8717 (N_8717,N_7292,N_7195);
and U8718 (N_8718,N_7554,N_7661);
nand U8719 (N_8719,N_7445,N_7064);
or U8720 (N_8720,N_7845,N_7164);
or U8721 (N_8721,N_7086,N_7991);
xnor U8722 (N_8722,N_7003,N_7184);
or U8723 (N_8723,N_7895,N_7869);
nand U8724 (N_8724,N_7792,N_7814);
xnor U8725 (N_8725,N_7699,N_7315);
and U8726 (N_8726,N_7707,N_7781);
and U8727 (N_8727,N_7657,N_7254);
or U8728 (N_8728,N_7663,N_7941);
and U8729 (N_8729,N_7788,N_7200);
nor U8730 (N_8730,N_7165,N_7609);
nor U8731 (N_8731,N_7038,N_7411);
xor U8732 (N_8732,N_7189,N_7903);
nor U8733 (N_8733,N_7899,N_7034);
and U8734 (N_8734,N_7089,N_7078);
nand U8735 (N_8735,N_7952,N_7275);
xnor U8736 (N_8736,N_7068,N_7531);
nand U8737 (N_8737,N_7778,N_7369);
xnor U8738 (N_8738,N_7343,N_7576);
nand U8739 (N_8739,N_7542,N_7857);
xnor U8740 (N_8740,N_7477,N_7690);
nand U8741 (N_8741,N_7459,N_7599);
nand U8742 (N_8742,N_7538,N_7874);
nand U8743 (N_8743,N_7101,N_7633);
xnor U8744 (N_8744,N_7908,N_7079);
xor U8745 (N_8745,N_7882,N_7797);
xor U8746 (N_8746,N_7585,N_7812);
nand U8747 (N_8747,N_7148,N_7289);
xor U8748 (N_8748,N_7675,N_7076);
xor U8749 (N_8749,N_7692,N_7277);
and U8750 (N_8750,N_7758,N_7395);
and U8751 (N_8751,N_7342,N_7710);
and U8752 (N_8752,N_7956,N_7856);
xnor U8753 (N_8753,N_7997,N_7533);
xor U8754 (N_8754,N_7321,N_7400);
and U8755 (N_8755,N_7521,N_7283);
xnor U8756 (N_8756,N_7069,N_7187);
nor U8757 (N_8757,N_7955,N_7291);
nor U8758 (N_8758,N_7540,N_7107);
and U8759 (N_8759,N_7966,N_7559);
xnor U8760 (N_8760,N_7527,N_7884);
nand U8761 (N_8761,N_7945,N_7804);
nor U8762 (N_8762,N_7705,N_7876);
nor U8763 (N_8763,N_7671,N_7276);
nand U8764 (N_8764,N_7606,N_7291);
or U8765 (N_8765,N_7235,N_7634);
nand U8766 (N_8766,N_7882,N_7423);
and U8767 (N_8767,N_7541,N_7757);
nand U8768 (N_8768,N_7609,N_7058);
or U8769 (N_8769,N_7803,N_7786);
xor U8770 (N_8770,N_7704,N_7783);
or U8771 (N_8771,N_7490,N_7252);
and U8772 (N_8772,N_7276,N_7468);
or U8773 (N_8773,N_7859,N_7416);
nand U8774 (N_8774,N_7421,N_7787);
xor U8775 (N_8775,N_7398,N_7763);
and U8776 (N_8776,N_7729,N_7483);
or U8777 (N_8777,N_7425,N_7047);
or U8778 (N_8778,N_7749,N_7584);
or U8779 (N_8779,N_7056,N_7067);
nor U8780 (N_8780,N_7460,N_7340);
nor U8781 (N_8781,N_7700,N_7562);
xor U8782 (N_8782,N_7924,N_7832);
xor U8783 (N_8783,N_7381,N_7896);
xnor U8784 (N_8784,N_7045,N_7419);
or U8785 (N_8785,N_7665,N_7992);
and U8786 (N_8786,N_7320,N_7143);
nor U8787 (N_8787,N_7280,N_7704);
nand U8788 (N_8788,N_7838,N_7909);
or U8789 (N_8789,N_7332,N_7620);
nand U8790 (N_8790,N_7568,N_7160);
nor U8791 (N_8791,N_7412,N_7347);
and U8792 (N_8792,N_7955,N_7002);
nor U8793 (N_8793,N_7917,N_7497);
xnor U8794 (N_8794,N_7762,N_7601);
nor U8795 (N_8795,N_7054,N_7565);
or U8796 (N_8796,N_7586,N_7077);
xnor U8797 (N_8797,N_7137,N_7890);
nand U8798 (N_8798,N_7885,N_7609);
xor U8799 (N_8799,N_7658,N_7211);
or U8800 (N_8800,N_7830,N_7842);
nand U8801 (N_8801,N_7860,N_7683);
and U8802 (N_8802,N_7613,N_7899);
nor U8803 (N_8803,N_7811,N_7110);
or U8804 (N_8804,N_7132,N_7985);
and U8805 (N_8805,N_7547,N_7961);
xor U8806 (N_8806,N_7376,N_7734);
nor U8807 (N_8807,N_7662,N_7262);
xor U8808 (N_8808,N_7019,N_7972);
nor U8809 (N_8809,N_7958,N_7772);
and U8810 (N_8810,N_7785,N_7546);
nor U8811 (N_8811,N_7910,N_7208);
xnor U8812 (N_8812,N_7506,N_7745);
and U8813 (N_8813,N_7824,N_7949);
and U8814 (N_8814,N_7903,N_7411);
nor U8815 (N_8815,N_7747,N_7878);
xor U8816 (N_8816,N_7401,N_7896);
and U8817 (N_8817,N_7468,N_7258);
or U8818 (N_8818,N_7884,N_7350);
or U8819 (N_8819,N_7254,N_7383);
or U8820 (N_8820,N_7627,N_7728);
and U8821 (N_8821,N_7858,N_7172);
nor U8822 (N_8822,N_7308,N_7909);
or U8823 (N_8823,N_7606,N_7738);
nand U8824 (N_8824,N_7994,N_7997);
xor U8825 (N_8825,N_7377,N_7755);
and U8826 (N_8826,N_7296,N_7878);
nand U8827 (N_8827,N_7440,N_7128);
and U8828 (N_8828,N_7399,N_7570);
xnor U8829 (N_8829,N_7204,N_7304);
nand U8830 (N_8830,N_7389,N_7215);
and U8831 (N_8831,N_7259,N_7969);
nor U8832 (N_8832,N_7894,N_7801);
and U8833 (N_8833,N_7409,N_7413);
xor U8834 (N_8834,N_7778,N_7013);
xor U8835 (N_8835,N_7448,N_7368);
nand U8836 (N_8836,N_7536,N_7623);
nor U8837 (N_8837,N_7716,N_7580);
and U8838 (N_8838,N_7919,N_7543);
xor U8839 (N_8839,N_7415,N_7568);
nand U8840 (N_8840,N_7497,N_7963);
and U8841 (N_8841,N_7138,N_7395);
nor U8842 (N_8842,N_7743,N_7514);
xnor U8843 (N_8843,N_7563,N_7135);
and U8844 (N_8844,N_7620,N_7731);
or U8845 (N_8845,N_7173,N_7143);
nor U8846 (N_8846,N_7678,N_7074);
and U8847 (N_8847,N_7740,N_7043);
or U8848 (N_8848,N_7201,N_7110);
and U8849 (N_8849,N_7140,N_7691);
and U8850 (N_8850,N_7902,N_7773);
and U8851 (N_8851,N_7145,N_7711);
nand U8852 (N_8852,N_7654,N_7093);
xor U8853 (N_8853,N_7523,N_7718);
nand U8854 (N_8854,N_7640,N_7636);
and U8855 (N_8855,N_7092,N_7562);
xor U8856 (N_8856,N_7505,N_7070);
nand U8857 (N_8857,N_7623,N_7775);
and U8858 (N_8858,N_7805,N_7116);
xor U8859 (N_8859,N_7955,N_7275);
nor U8860 (N_8860,N_7749,N_7138);
or U8861 (N_8861,N_7287,N_7674);
nand U8862 (N_8862,N_7383,N_7757);
and U8863 (N_8863,N_7891,N_7155);
xor U8864 (N_8864,N_7438,N_7226);
nand U8865 (N_8865,N_7053,N_7762);
xor U8866 (N_8866,N_7455,N_7236);
xor U8867 (N_8867,N_7060,N_7743);
xnor U8868 (N_8868,N_7571,N_7401);
nand U8869 (N_8869,N_7582,N_7564);
or U8870 (N_8870,N_7666,N_7866);
and U8871 (N_8871,N_7393,N_7960);
and U8872 (N_8872,N_7761,N_7075);
or U8873 (N_8873,N_7353,N_7705);
xnor U8874 (N_8874,N_7985,N_7832);
or U8875 (N_8875,N_7513,N_7866);
nand U8876 (N_8876,N_7254,N_7466);
nor U8877 (N_8877,N_7614,N_7648);
nor U8878 (N_8878,N_7594,N_7306);
xor U8879 (N_8879,N_7052,N_7131);
nor U8880 (N_8880,N_7338,N_7782);
nor U8881 (N_8881,N_7190,N_7375);
nand U8882 (N_8882,N_7004,N_7563);
nand U8883 (N_8883,N_7643,N_7399);
nor U8884 (N_8884,N_7416,N_7187);
nand U8885 (N_8885,N_7857,N_7239);
nand U8886 (N_8886,N_7877,N_7691);
and U8887 (N_8887,N_7355,N_7559);
nor U8888 (N_8888,N_7542,N_7914);
and U8889 (N_8889,N_7701,N_7608);
nand U8890 (N_8890,N_7545,N_7788);
or U8891 (N_8891,N_7711,N_7956);
and U8892 (N_8892,N_7618,N_7185);
xor U8893 (N_8893,N_7674,N_7395);
or U8894 (N_8894,N_7836,N_7702);
or U8895 (N_8895,N_7816,N_7018);
nor U8896 (N_8896,N_7989,N_7943);
or U8897 (N_8897,N_7443,N_7369);
or U8898 (N_8898,N_7993,N_7399);
and U8899 (N_8899,N_7723,N_7785);
or U8900 (N_8900,N_7388,N_7566);
nor U8901 (N_8901,N_7508,N_7813);
nor U8902 (N_8902,N_7969,N_7878);
nand U8903 (N_8903,N_7602,N_7892);
nor U8904 (N_8904,N_7756,N_7170);
and U8905 (N_8905,N_7224,N_7076);
xor U8906 (N_8906,N_7992,N_7538);
nor U8907 (N_8907,N_7104,N_7325);
and U8908 (N_8908,N_7589,N_7705);
xor U8909 (N_8909,N_7514,N_7324);
nand U8910 (N_8910,N_7633,N_7212);
and U8911 (N_8911,N_7908,N_7929);
nor U8912 (N_8912,N_7410,N_7005);
nor U8913 (N_8913,N_7386,N_7587);
or U8914 (N_8914,N_7448,N_7197);
nand U8915 (N_8915,N_7645,N_7084);
nor U8916 (N_8916,N_7716,N_7429);
nand U8917 (N_8917,N_7280,N_7290);
nand U8918 (N_8918,N_7821,N_7168);
nand U8919 (N_8919,N_7704,N_7161);
and U8920 (N_8920,N_7042,N_7241);
nor U8921 (N_8921,N_7612,N_7813);
or U8922 (N_8922,N_7435,N_7372);
and U8923 (N_8923,N_7619,N_7374);
and U8924 (N_8924,N_7868,N_7783);
and U8925 (N_8925,N_7731,N_7685);
nand U8926 (N_8926,N_7436,N_7913);
and U8927 (N_8927,N_7821,N_7898);
nand U8928 (N_8928,N_7769,N_7556);
xor U8929 (N_8929,N_7769,N_7590);
xnor U8930 (N_8930,N_7181,N_7379);
and U8931 (N_8931,N_7699,N_7134);
nand U8932 (N_8932,N_7953,N_7805);
nand U8933 (N_8933,N_7831,N_7829);
nor U8934 (N_8934,N_7654,N_7794);
and U8935 (N_8935,N_7514,N_7096);
and U8936 (N_8936,N_7406,N_7964);
or U8937 (N_8937,N_7837,N_7534);
or U8938 (N_8938,N_7428,N_7994);
nor U8939 (N_8939,N_7920,N_7862);
xor U8940 (N_8940,N_7379,N_7772);
or U8941 (N_8941,N_7675,N_7593);
nand U8942 (N_8942,N_7806,N_7972);
or U8943 (N_8943,N_7329,N_7277);
and U8944 (N_8944,N_7356,N_7623);
xnor U8945 (N_8945,N_7808,N_7756);
xor U8946 (N_8946,N_7126,N_7858);
or U8947 (N_8947,N_7860,N_7775);
xor U8948 (N_8948,N_7518,N_7235);
nand U8949 (N_8949,N_7480,N_7183);
nor U8950 (N_8950,N_7459,N_7148);
and U8951 (N_8951,N_7151,N_7423);
nor U8952 (N_8952,N_7994,N_7649);
or U8953 (N_8953,N_7174,N_7946);
and U8954 (N_8954,N_7441,N_7387);
or U8955 (N_8955,N_7728,N_7432);
nor U8956 (N_8956,N_7182,N_7880);
and U8957 (N_8957,N_7592,N_7579);
xnor U8958 (N_8958,N_7031,N_7750);
or U8959 (N_8959,N_7704,N_7088);
or U8960 (N_8960,N_7640,N_7024);
or U8961 (N_8961,N_7658,N_7175);
nor U8962 (N_8962,N_7380,N_7118);
nand U8963 (N_8963,N_7947,N_7880);
and U8964 (N_8964,N_7513,N_7894);
or U8965 (N_8965,N_7223,N_7452);
and U8966 (N_8966,N_7274,N_7700);
xor U8967 (N_8967,N_7513,N_7042);
or U8968 (N_8968,N_7582,N_7239);
nor U8969 (N_8969,N_7088,N_7411);
nor U8970 (N_8970,N_7114,N_7741);
nor U8971 (N_8971,N_7852,N_7784);
xnor U8972 (N_8972,N_7937,N_7835);
or U8973 (N_8973,N_7720,N_7999);
nor U8974 (N_8974,N_7554,N_7091);
or U8975 (N_8975,N_7691,N_7821);
and U8976 (N_8976,N_7602,N_7441);
and U8977 (N_8977,N_7623,N_7218);
and U8978 (N_8978,N_7478,N_7086);
and U8979 (N_8979,N_7978,N_7390);
nand U8980 (N_8980,N_7153,N_7017);
and U8981 (N_8981,N_7529,N_7128);
and U8982 (N_8982,N_7119,N_7927);
nor U8983 (N_8983,N_7212,N_7931);
nor U8984 (N_8984,N_7218,N_7171);
nand U8985 (N_8985,N_7933,N_7101);
nand U8986 (N_8986,N_7900,N_7720);
or U8987 (N_8987,N_7041,N_7465);
xnor U8988 (N_8988,N_7615,N_7218);
or U8989 (N_8989,N_7936,N_7023);
or U8990 (N_8990,N_7997,N_7174);
and U8991 (N_8991,N_7726,N_7910);
and U8992 (N_8992,N_7384,N_7764);
and U8993 (N_8993,N_7951,N_7620);
nand U8994 (N_8994,N_7914,N_7726);
nand U8995 (N_8995,N_7214,N_7980);
nand U8996 (N_8996,N_7002,N_7162);
and U8997 (N_8997,N_7978,N_7612);
or U8998 (N_8998,N_7893,N_7722);
and U8999 (N_8999,N_7544,N_7917);
xnor U9000 (N_9000,N_8031,N_8549);
nand U9001 (N_9001,N_8240,N_8003);
and U9002 (N_9002,N_8650,N_8762);
or U9003 (N_9003,N_8290,N_8786);
nor U9004 (N_9004,N_8953,N_8531);
and U9005 (N_9005,N_8026,N_8716);
xnor U9006 (N_9006,N_8485,N_8873);
and U9007 (N_9007,N_8360,N_8681);
nor U9008 (N_9008,N_8028,N_8570);
xnor U9009 (N_9009,N_8179,N_8283);
nand U9010 (N_9010,N_8673,N_8637);
nor U9011 (N_9011,N_8501,N_8864);
xnor U9012 (N_9012,N_8265,N_8508);
and U9013 (N_9013,N_8550,N_8809);
xor U9014 (N_9014,N_8312,N_8876);
or U9015 (N_9015,N_8958,N_8436);
xnor U9016 (N_9016,N_8229,N_8241);
or U9017 (N_9017,N_8074,N_8203);
nor U9018 (N_9018,N_8815,N_8005);
or U9019 (N_9019,N_8522,N_8424);
and U9020 (N_9020,N_8530,N_8445);
xor U9021 (N_9021,N_8612,N_8085);
or U9022 (N_9022,N_8606,N_8390);
xnor U9023 (N_9023,N_8210,N_8342);
nor U9024 (N_9024,N_8202,N_8347);
nand U9025 (N_9025,N_8954,N_8106);
and U9026 (N_9026,N_8687,N_8351);
and U9027 (N_9027,N_8785,N_8423);
nand U9028 (N_9028,N_8669,N_8759);
or U9029 (N_9029,N_8946,N_8220);
or U9030 (N_9030,N_8327,N_8111);
xor U9031 (N_9031,N_8126,N_8438);
and U9032 (N_9032,N_8469,N_8150);
and U9033 (N_9033,N_8533,N_8018);
nor U9034 (N_9034,N_8472,N_8398);
nor U9035 (N_9035,N_8734,N_8224);
xor U9036 (N_9036,N_8409,N_8050);
nand U9037 (N_9037,N_8643,N_8113);
or U9038 (N_9038,N_8845,N_8162);
xnor U9039 (N_9039,N_8857,N_8729);
nor U9040 (N_9040,N_8990,N_8339);
nand U9041 (N_9041,N_8260,N_8965);
xor U9042 (N_9042,N_8594,N_8223);
and U9043 (N_9043,N_8581,N_8082);
nand U9044 (N_9044,N_8844,N_8127);
nand U9045 (N_9045,N_8000,N_8035);
and U9046 (N_9046,N_8623,N_8338);
nand U9047 (N_9047,N_8110,N_8410);
or U9048 (N_9048,N_8186,N_8727);
nand U9049 (N_9049,N_8546,N_8077);
nand U9050 (N_9050,N_8197,N_8417);
or U9051 (N_9051,N_8731,N_8314);
or U9052 (N_9052,N_8289,N_8416);
nand U9053 (N_9053,N_8025,N_8929);
xnor U9054 (N_9054,N_8306,N_8776);
nand U9055 (N_9055,N_8945,N_8340);
nand U9056 (N_9056,N_8405,N_8739);
nand U9057 (N_9057,N_8829,N_8732);
and U9058 (N_9058,N_8333,N_8832);
nand U9059 (N_9059,N_8964,N_8935);
and U9060 (N_9060,N_8822,N_8872);
xnor U9061 (N_9061,N_8835,N_8985);
nand U9062 (N_9062,N_8824,N_8242);
nor U9063 (N_9063,N_8638,N_8881);
nand U9064 (N_9064,N_8529,N_8853);
nor U9065 (N_9065,N_8118,N_8366);
and U9066 (N_9066,N_8038,N_8123);
nand U9067 (N_9067,N_8651,N_8419);
and U9068 (N_9068,N_8209,N_8067);
or U9069 (N_9069,N_8457,N_8898);
or U9070 (N_9070,N_8742,N_8816);
nor U9071 (N_9071,N_8023,N_8052);
nand U9072 (N_9072,N_8747,N_8310);
nor U9073 (N_9073,N_8622,N_8129);
and U9074 (N_9074,N_8486,N_8072);
nor U9075 (N_9075,N_8323,N_8171);
and U9076 (N_9076,N_8010,N_8942);
xnor U9077 (N_9077,N_8849,N_8497);
or U9078 (N_9078,N_8591,N_8773);
nor U9079 (N_9079,N_8795,N_8659);
xnor U9080 (N_9080,N_8578,N_8244);
or U9081 (N_9081,N_8138,N_8620);
xor U9082 (N_9082,N_8356,N_8281);
and U9083 (N_9083,N_8452,N_8218);
or U9084 (N_9084,N_8839,N_8427);
nor U9085 (N_9085,N_8752,N_8167);
or U9086 (N_9086,N_8108,N_8482);
and U9087 (N_9087,N_8598,N_8924);
and U9088 (N_9088,N_8198,N_8459);
xnor U9089 (N_9089,N_8880,N_8913);
nand U9090 (N_9090,N_8928,N_8668);
nand U9091 (N_9091,N_8719,N_8093);
xnor U9092 (N_9092,N_8922,N_8261);
and U9093 (N_9093,N_8502,N_8274);
and U9094 (N_9094,N_8429,N_8784);
and U9095 (N_9095,N_8304,N_8733);
or U9096 (N_9096,N_8861,N_8201);
nand U9097 (N_9097,N_8048,N_8233);
xor U9098 (N_9098,N_8678,N_8315);
nand U9099 (N_9099,N_8647,N_8331);
and U9100 (N_9100,N_8053,N_8661);
xor U9101 (N_9101,N_8599,N_8217);
nor U9102 (N_9102,N_8547,N_8316);
nor U9103 (N_9103,N_8807,N_8634);
nor U9104 (N_9104,N_8148,N_8700);
or U9105 (N_9105,N_8563,N_8385);
and U9106 (N_9106,N_8640,N_8483);
xor U9107 (N_9107,N_8041,N_8827);
nor U9108 (N_9108,N_8032,N_8136);
nor U9109 (N_9109,N_8828,N_8925);
nand U9110 (N_9110,N_8934,N_8181);
xor U9111 (N_9111,N_8278,N_8516);
nand U9112 (N_9112,N_8037,N_8627);
nor U9113 (N_9113,N_8979,N_8866);
xor U9114 (N_9114,N_8101,N_8595);
and U9115 (N_9115,N_8628,N_8500);
xor U9116 (N_9116,N_8395,N_8291);
nand U9117 (N_9117,N_8400,N_8768);
or U9118 (N_9118,N_8158,N_8247);
nand U9119 (N_9119,N_8653,N_8104);
and U9120 (N_9120,N_8286,N_8205);
nor U9121 (N_9121,N_8751,N_8115);
xnor U9122 (N_9122,N_8860,N_8213);
nor U9123 (N_9123,N_8112,N_8960);
xnor U9124 (N_9124,N_8195,N_8470);
xnor U9125 (N_9125,N_8166,N_8036);
nand U9126 (N_9126,N_8130,N_8941);
nand U9127 (N_9127,N_8649,N_8276);
xnor U9128 (N_9128,N_8488,N_8963);
nand U9129 (N_9129,N_8103,N_8272);
and U9130 (N_9130,N_8362,N_8883);
and U9131 (N_9131,N_8034,N_8114);
and U9132 (N_9132,N_8094,N_8422);
nand U9133 (N_9133,N_8042,N_8294);
nand U9134 (N_9134,N_8474,N_8688);
nor U9135 (N_9135,N_8617,N_8808);
nor U9136 (N_9136,N_8091,N_8630);
xor U9137 (N_9137,N_8803,N_8430);
nor U9138 (N_9138,N_8080,N_8001);
and U9139 (N_9139,N_8345,N_8813);
xnor U9140 (N_9140,N_8792,N_8788);
or U9141 (N_9141,N_8851,N_8690);
xor U9142 (N_9142,N_8939,N_8479);
xnor U9143 (N_9143,N_8874,N_8288);
or U9144 (N_9144,N_8192,N_8543);
xor U9145 (N_9145,N_8377,N_8368);
nand U9146 (N_9146,N_8277,N_8884);
nand U9147 (N_9147,N_8043,N_8841);
xnor U9148 (N_9148,N_8680,N_8583);
nand U9149 (N_9149,N_8267,N_8567);
xor U9150 (N_9150,N_8301,N_8391);
or U9151 (N_9151,N_8441,N_8341);
xor U9152 (N_9152,N_8433,N_8088);
nand U9153 (N_9153,N_8949,N_8648);
xnor U9154 (N_9154,N_8825,N_8380);
nand U9155 (N_9155,N_8014,N_8475);
or U9156 (N_9156,N_8151,N_8105);
or U9157 (N_9157,N_8473,N_8319);
and U9158 (N_9158,N_8476,N_8125);
xnor U9159 (N_9159,N_8145,N_8877);
xor U9160 (N_9160,N_8756,N_8976);
and U9161 (N_9161,N_8216,N_8777);
nand U9162 (N_9162,N_8057,N_8592);
and U9163 (N_9163,N_8477,N_8968);
nand U9164 (N_9164,N_8449,N_8701);
nand U9165 (N_9165,N_8789,N_8525);
xnor U9166 (N_9166,N_8830,N_8079);
nor U9167 (N_9167,N_8749,N_8697);
xor U9168 (N_9168,N_8305,N_8453);
xor U9169 (N_9169,N_8714,N_8448);
nor U9170 (N_9170,N_8682,N_8631);
or U9171 (N_9171,N_8590,N_8487);
and U9172 (N_9172,N_8748,N_8607);
or U9173 (N_9173,N_8962,N_8320);
xor U9174 (N_9174,N_8442,N_8551);
nand U9175 (N_9175,N_8520,N_8615);
or U9176 (N_9176,N_8293,N_8540);
nor U9177 (N_9177,N_8843,N_8373);
or U9178 (N_9178,N_8047,N_8977);
nand U9179 (N_9179,N_8646,N_8624);
or U9180 (N_9180,N_8246,N_8299);
nor U9181 (N_9181,N_8667,N_8464);
nand U9182 (N_9182,N_8806,N_8699);
nor U9183 (N_9183,N_8772,N_8725);
xor U9184 (N_9184,N_8582,N_8914);
or U9185 (N_9185,N_8255,N_8413);
nand U9186 (N_9186,N_8619,N_8322);
nor U9187 (N_9187,N_8693,N_8975);
or U9188 (N_9188,N_8794,N_8002);
nand U9189 (N_9189,N_8579,N_8292);
or U9190 (N_9190,N_8737,N_8495);
or U9191 (N_9191,N_8109,N_8616);
and U9192 (N_9192,N_8444,N_8758);
and U9193 (N_9193,N_8344,N_8403);
or U9194 (N_9194,N_8394,N_8933);
xnor U9195 (N_9195,N_8326,N_8662);
xnor U9196 (N_9196,N_8039,N_8134);
nand U9197 (N_9197,N_8801,N_8484);
or U9198 (N_9198,N_8371,N_8774);
nand U9199 (N_9199,N_8099,N_8092);
nand U9200 (N_9200,N_8059,N_8013);
and U9201 (N_9201,N_8262,N_8852);
or U9202 (N_9202,N_8219,N_8698);
nor U9203 (N_9203,N_8415,N_8709);
xnor U9204 (N_9204,N_8566,N_8076);
or U9205 (N_9205,N_8764,N_8863);
nor U9206 (N_9206,N_8585,N_8251);
nor U9207 (N_9207,N_8258,N_8902);
nand U9208 (N_9208,N_8871,N_8257);
nor U9209 (N_9209,N_8143,N_8055);
xnor U9210 (N_9210,N_8402,N_8885);
or U9211 (N_9211,N_8797,N_8544);
nand U9212 (N_9212,N_8334,N_8995);
and U9213 (N_9213,N_8660,N_8707);
nor U9214 (N_9214,N_8069,N_8770);
and U9215 (N_9215,N_8819,N_8608);
nand U9216 (N_9216,N_8689,N_8703);
or U9217 (N_9217,N_8943,N_8308);
nand U9218 (N_9218,N_8626,N_8528);
or U9219 (N_9219,N_8019,N_8955);
nand U9220 (N_9220,N_8587,N_8896);
or U9221 (N_9221,N_8364,N_8180);
or U9222 (N_9222,N_8918,N_8895);
and U9223 (N_9223,N_8576,N_8404);
nand U9224 (N_9224,N_8900,N_8554);
nor U9225 (N_9225,N_8972,N_8679);
nor U9226 (N_9226,N_8033,N_8812);
or U9227 (N_9227,N_8992,N_8800);
and U9228 (N_9228,N_8172,N_8024);
nor U9229 (N_9229,N_8798,N_8083);
or U9230 (N_9230,N_8128,N_8793);
nand U9231 (N_9231,N_8639,N_8119);
and U9232 (N_9232,N_8512,N_8636);
nor U9233 (N_9233,N_8058,N_8771);
or U9234 (N_9234,N_8905,N_8597);
nand U9235 (N_9235,N_8046,N_8996);
or U9236 (N_9236,N_8169,N_8685);
or U9237 (N_9237,N_8984,N_8834);
nor U9238 (N_9238,N_8361,N_8894);
xnor U9239 (N_9239,N_8600,N_8517);
and U9240 (N_9240,N_8147,N_8817);
xnor U9241 (N_9241,N_8221,N_8666);
xnor U9242 (N_9242,N_8102,N_8153);
or U9243 (N_9243,N_8514,N_8753);
xnor U9244 (N_9244,N_8354,N_8761);
nand U9245 (N_9245,N_8414,N_8357);
xnor U9246 (N_9246,N_8492,N_8769);
or U9247 (N_9247,N_8621,N_8947);
and U9248 (N_9248,N_8062,N_8865);
nand U9249 (N_9249,N_8467,N_8051);
nand U9250 (N_9250,N_8190,N_8132);
or U9251 (N_9251,N_8967,N_8207);
and U9252 (N_9252,N_8892,N_8012);
and U9253 (N_9253,N_8389,N_8736);
or U9254 (N_9254,N_8948,N_8904);
or U9255 (N_9255,N_8826,N_8493);
xnor U9256 (N_9256,N_8847,N_8565);
and U9257 (N_9257,N_8559,N_8738);
xor U9258 (N_9258,N_8527,N_8743);
nor U9259 (N_9259,N_8225,N_8642);
xor U9260 (N_9260,N_8746,N_8674);
nor U9261 (N_9261,N_8157,N_8907);
nor U9262 (N_9262,N_8382,N_8252);
or U9263 (N_9263,N_8135,N_8496);
nor U9264 (N_9264,N_8713,N_8574);
or U9265 (N_9265,N_8396,N_8886);
nand U9266 (N_9266,N_8609,N_8586);
nand U9267 (N_9267,N_8564,N_8555);
nand U9268 (N_9268,N_8952,N_8061);
or U9269 (N_9269,N_8426,N_8683);
nor U9270 (N_9270,N_8121,N_8471);
or U9271 (N_9271,N_8878,N_8236);
and U9272 (N_9272,N_8481,N_8071);
or U9273 (N_9273,N_8889,N_8245);
nand U9274 (N_9274,N_8399,N_8718);
or U9275 (N_9275,N_8654,N_8658);
or U9276 (N_9276,N_8912,N_8098);
and U9277 (N_9277,N_8726,N_8780);
nor U9278 (N_9278,N_8401,N_8836);
xor U9279 (N_9279,N_8275,N_8020);
xor U9280 (N_9280,N_8927,N_8359);
nand U9281 (N_9281,N_8144,N_8117);
nand U9282 (N_9282,N_8614,N_8087);
or U9283 (N_9283,N_8397,N_8178);
xnor U9284 (N_9284,N_8328,N_8060);
nor U9285 (N_9285,N_8657,N_8859);
and U9286 (N_9286,N_8970,N_8412);
and U9287 (N_9287,N_8264,N_8532);
xnor U9288 (N_9288,N_8572,N_8930);
xor U9289 (N_9289,N_8577,N_8722);
or U9290 (N_9290,N_8352,N_8466);
xnor U9291 (N_9291,N_8384,N_8802);
and U9292 (N_9292,N_8421,N_8510);
nand U9293 (N_9293,N_8163,N_8096);
xnor U9294 (N_9294,N_8519,N_8507);
or U9295 (N_9295,N_8675,N_8804);
xnor U9296 (N_9296,N_8450,N_8686);
or U9297 (N_9297,N_8008,N_8165);
and U9298 (N_9298,N_8056,N_8363);
nand U9299 (N_9299,N_8021,N_8189);
or U9300 (N_9300,N_8980,N_8222);
nor U9301 (N_9301,N_8956,N_8386);
and U9302 (N_9302,N_8916,N_8664);
xnor U9303 (N_9303,N_8440,N_8022);
xnor U9304 (N_9304,N_8387,N_8271);
or U9305 (N_9305,N_8537,N_8692);
or U9306 (N_9306,N_8044,N_8081);
and U9307 (N_9307,N_8282,N_8856);
or U9308 (N_9308,N_8461,N_8875);
and U9309 (N_9309,N_8437,N_8232);
or U9310 (N_9310,N_8456,N_8903);
or U9311 (N_9311,N_8355,N_8137);
xnor U9312 (N_9312,N_8455,N_8750);
and U9313 (N_9313,N_8318,N_8879);
xor U9314 (N_9314,N_8296,N_8671);
nor U9315 (N_9315,N_8848,N_8173);
xnor U9316 (N_9316,N_8635,N_8765);
nor U9317 (N_9317,N_8238,N_8840);
and U9318 (N_9318,N_8231,N_8330);
xnor U9319 (N_9319,N_8006,N_8040);
xnor U9320 (N_9320,N_8677,N_8237);
nand U9321 (N_9321,N_8505,N_8655);
or U9322 (N_9322,N_8349,N_8432);
or U9323 (N_9323,N_8155,N_8175);
or U9324 (N_9324,N_8994,N_8618);
nand U9325 (N_9325,N_8915,N_8858);
and U9326 (N_9326,N_8862,N_8775);
nand U9327 (N_9327,N_8131,N_8270);
xnor U9328 (N_9328,N_8183,N_8346);
or U9329 (N_9329,N_8263,N_8004);
or U9330 (N_9330,N_8989,N_8506);
or U9331 (N_9331,N_8446,N_8029);
nand U9332 (N_9332,N_8372,N_8250);
and U9333 (N_9333,N_8589,N_8632);
nor U9334 (N_9334,N_8468,N_8523);
or U9335 (N_9335,N_8498,N_8604);
nor U9336 (N_9336,N_8909,N_8521);
nor U9337 (N_9337,N_8285,N_8249);
or U9338 (N_9338,N_8336,N_8447);
nor U9339 (N_9339,N_8141,N_8268);
xnor U9340 (N_9340,N_8230,N_8920);
or U9341 (N_9341,N_8782,N_8712);
xnor U9342 (N_9342,N_8937,N_8324);
or U9343 (N_9343,N_8309,N_8458);
nor U9344 (N_9344,N_8494,N_8159);
and U9345 (N_9345,N_8227,N_8708);
nor U9346 (N_9346,N_8116,N_8961);
and U9347 (N_9347,N_8694,N_8870);
xor U9348 (N_9348,N_8297,N_8078);
and U9349 (N_9349,N_8100,N_8228);
and U9350 (N_9350,N_8027,N_8571);
and U9351 (N_9351,N_8676,N_8931);
and U9352 (N_9352,N_8706,N_8374);
nand U9353 (N_9353,N_8451,N_8735);
or U9354 (N_9354,N_8139,N_8140);
xor U9355 (N_9355,N_8066,N_8997);
or U9356 (N_9356,N_8787,N_8569);
xnor U9357 (N_9357,N_8462,N_8406);
and U9358 (N_9358,N_8411,N_8204);
or U9359 (N_9359,N_8901,N_8791);
and U9360 (N_9360,N_8392,N_8534);
and U9361 (N_9361,N_8810,N_8820);
nand U9362 (N_9362,N_8882,N_8212);
nor U9363 (N_9363,N_8465,N_8613);
nand U9364 (N_9364,N_8435,N_8524);
xnor U9365 (N_9365,N_8538,N_8652);
and U9366 (N_9366,N_8542,N_8783);
nor U9367 (N_9367,N_8710,N_8358);
or U9368 (N_9368,N_8420,N_8974);
nand U9369 (N_9369,N_8545,N_8084);
xnor U9370 (N_9370,N_8723,N_8663);
or U9371 (N_9371,N_8645,N_8717);
or U9372 (N_9372,N_8971,N_8408);
xor U9373 (N_9373,N_8015,N_8379);
nand U9374 (N_9374,N_8656,N_8187);
nand U9375 (N_9375,N_8161,N_8378);
nand U9376 (N_9376,N_8325,N_8846);
and U9377 (N_9377,N_8910,N_8388);
nand U9378 (N_9378,N_8065,N_8821);
nor U9379 (N_9379,N_8174,N_8369);
xnor U9380 (N_9380,N_8383,N_8206);
xor U9381 (N_9381,N_8625,N_8199);
nand U9382 (N_9382,N_8503,N_8248);
and U9383 (N_9383,N_8226,N_8923);
and U9384 (N_9384,N_8665,N_8568);
or U9385 (N_9385,N_8811,N_8313);
and U9386 (N_9386,N_8329,N_8350);
and U9387 (N_9387,N_8603,N_8715);
or U9388 (N_9388,N_8269,N_8767);
xor U9389 (N_9389,N_8182,N_8781);
nor U9390 (N_9390,N_8644,N_8234);
or U9391 (N_9391,N_8991,N_8478);
and U9392 (N_9392,N_8156,N_8208);
or U9393 (N_9393,N_8796,N_8443);
and U9394 (N_9394,N_8348,N_8584);
xor U9395 (N_9395,N_8575,N_8300);
xor U9396 (N_9396,N_8375,N_8343);
or U9397 (N_9397,N_8670,N_8254);
and U9398 (N_9398,N_8431,N_8705);
nor U9399 (N_9399,N_8951,N_8818);
and U9400 (N_9400,N_8321,N_8897);
nor U9401 (N_9401,N_8766,N_8823);
or U9402 (N_9402,N_8454,N_8588);
or U9403 (N_9403,N_8917,N_8239);
nor U9404 (N_9404,N_8491,N_8298);
or U9405 (N_9405,N_8214,N_8302);
and U9406 (N_9406,N_8691,N_8370);
xnor U9407 (N_9407,N_8287,N_8741);
and U9408 (N_9408,N_8799,N_8704);
nand U9409 (N_9409,N_8504,N_8256);
nand U9410 (N_9410,N_8535,N_8908);
nand U9411 (N_9411,N_8463,N_8016);
xnor U9412 (N_9412,N_8740,N_8966);
or U9413 (N_9413,N_8728,N_8911);
nor U9414 (N_9414,N_8999,N_8556);
and U9415 (N_9415,N_8191,N_8253);
and U9416 (N_9416,N_8778,N_8526);
xor U9417 (N_9417,N_8200,N_8950);
nor U9418 (N_9418,N_8007,N_8779);
or U9419 (N_9419,N_8596,N_8899);
or U9420 (N_9420,N_8188,N_8986);
xor U9421 (N_9421,N_8009,N_8120);
or U9422 (N_9422,N_8295,N_8185);
or U9423 (N_9423,N_8696,N_8702);
xor U9424 (N_9424,N_8610,N_8850);
xnor U9425 (N_9425,N_8365,N_8407);
nand U9426 (N_9426,N_8196,N_8434);
and U9427 (N_9427,N_8097,N_8168);
nor U9428 (N_9428,N_8938,N_8154);
nand U9429 (N_9429,N_8919,N_8284);
or U9430 (N_9430,N_8307,N_8605);
or U9431 (N_9431,N_8558,N_8303);
and U9432 (N_9432,N_8317,N_8353);
or U9433 (N_9433,N_8944,N_8982);
or U9434 (N_9434,N_8593,N_8460);
nand U9435 (N_9435,N_8633,N_8867);
nor U9436 (N_9436,N_8418,N_8489);
nand U9437 (N_9437,N_8641,N_8215);
nand U9438 (N_9438,N_8393,N_8981);
xnor U9439 (N_9439,N_8754,N_8073);
nand U9440 (N_9440,N_8509,N_8932);
or U9441 (N_9441,N_8539,N_8011);
nand U9442 (N_9442,N_8601,N_8367);
nor U9443 (N_9443,N_8017,N_8720);
or U9444 (N_9444,N_8695,N_8573);
nor U9445 (N_9445,N_8054,N_8064);
xor U9446 (N_9446,N_8959,N_8757);
nor U9447 (N_9447,N_8518,N_8998);
or U9448 (N_9448,N_8763,N_8439);
nor U9449 (N_9449,N_8611,N_8152);
and U9450 (N_9450,N_8160,N_8854);
nand U9451 (N_9451,N_8211,N_8095);
xor U9452 (N_9452,N_8721,N_8869);
nor U9453 (N_9453,N_8887,N_8833);
nand U9454 (N_9454,N_8122,N_8133);
nor U9455 (N_9455,N_8973,N_8089);
and U9456 (N_9456,N_8030,N_8906);
and U9457 (N_9457,N_8730,N_8480);
nand U9458 (N_9458,N_8711,N_8243);
and U9459 (N_9459,N_8890,N_8259);
xnor U9460 (N_9460,N_8045,N_8553);
nor U9461 (N_9461,N_8602,N_8988);
xor U9462 (N_9462,N_8490,N_8337);
and U9463 (N_9463,N_8983,N_8993);
nand U9464 (N_9464,N_8760,N_8838);
nor U9465 (N_9465,N_8149,N_8273);
or U9466 (N_9466,N_8888,N_8266);
nand U9467 (N_9467,N_8170,N_8376);
xor U9468 (N_9468,N_8744,N_8684);
nor U9469 (N_9469,N_8957,N_8969);
nand U9470 (N_9470,N_8536,N_8831);
and U9471 (N_9471,N_8755,N_8049);
and U9472 (N_9472,N_8311,N_8560);
or U9473 (N_9473,N_8107,N_8515);
or U9474 (N_9474,N_8842,N_8561);
nand U9475 (N_9475,N_8177,N_8562);
nand U9476 (N_9476,N_8552,N_8629);
or U9477 (N_9477,N_8541,N_8837);
nor U9478 (N_9478,N_8511,N_8235);
nor U9479 (N_9479,N_8280,N_8332);
nand U9480 (N_9480,N_8987,N_8855);
nor U9481 (N_9481,N_8893,N_8194);
nor U9482 (N_9482,N_8921,N_8279);
nor U9483 (N_9483,N_8580,N_8724);
xnor U9484 (N_9484,N_8513,N_8335);
xor U9485 (N_9485,N_8090,N_8164);
nand U9486 (N_9486,N_8063,N_8557);
nor U9487 (N_9487,N_8075,N_8978);
nor U9488 (N_9488,N_8176,N_8745);
xor U9489 (N_9489,N_8184,N_8381);
or U9490 (N_9490,N_8814,N_8868);
xor U9491 (N_9491,N_8891,N_8805);
or U9492 (N_9492,N_8142,N_8672);
or U9493 (N_9493,N_8790,N_8936);
and U9494 (N_9494,N_8070,N_8068);
xnor U9495 (N_9495,N_8124,N_8926);
and U9496 (N_9496,N_8499,N_8940);
and U9497 (N_9497,N_8086,N_8425);
xnor U9498 (N_9498,N_8428,N_8146);
or U9499 (N_9499,N_8548,N_8193);
or U9500 (N_9500,N_8061,N_8074);
or U9501 (N_9501,N_8245,N_8810);
and U9502 (N_9502,N_8301,N_8895);
nor U9503 (N_9503,N_8418,N_8122);
nor U9504 (N_9504,N_8265,N_8852);
nand U9505 (N_9505,N_8145,N_8393);
nor U9506 (N_9506,N_8861,N_8483);
or U9507 (N_9507,N_8735,N_8247);
or U9508 (N_9508,N_8611,N_8564);
xnor U9509 (N_9509,N_8837,N_8959);
or U9510 (N_9510,N_8865,N_8080);
and U9511 (N_9511,N_8075,N_8135);
nand U9512 (N_9512,N_8132,N_8594);
and U9513 (N_9513,N_8861,N_8430);
nand U9514 (N_9514,N_8358,N_8351);
nor U9515 (N_9515,N_8061,N_8700);
nor U9516 (N_9516,N_8348,N_8726);
xnor U9517 (N_9517,N_8412,N_8026);
or U9518 (N_9518,N_8372,N_8578);
xnor U9519 (N_9519,N_8590,N_8257);
or U9520 (N_9520,N_8283,N_8941);
nand U9521 (N_9521,N_8016,N_8336);
nand U9522 (N_9522,N_8965,N_8152);
nand U9523 (N_9523,N_8656,N_8482);
xnor U9524 (N_9524,N_8237,N_8540);
xor U9525 (N_9525,N_8914,N_8462);
nor U9526 (N_9526,N_8546,N_8161);
or U9527 (N_9527,N_8592,N_8207);
or U9528 (N_9528,N_8166,N_8377);
nand U9529 (N_9529,N_8540,N_8001);
and U9530 (N_9530,N_8004,N_8421);
and U9531 (N_9531,N_8200,N_8408);
xor U9532 (N_9532,N_8768,N_8010);
nor U9533 (N_9533,N_8102,N_8187);
nand U9534 (N_9534,N_8677,N_8059);
xnor U9535 (N_9535,N_8819,N_8568);
xnor U9536 (N_9536,N_8834,N_8364);
xor U9537 (N_9537,N_8989,N_8420);
nand U9538 (N_9538,N_8901,N_8517);
nand U9539 (N_9539,N_8394,N_8058);
nand U9540 (N_9540,N_8662,N_8363);
and U9541 (N_9541,N_8396,N_8813);
and U9542 (N_9542,N_8594,N_8030);
or U9543 (N_9543,N_8979,N_8017);
and U9544 (N_9544,N_8289,N_8551);
nand U9545 (N_9545,N_8453,N_8210);
xnor U9546 (N_9546,N_8428,N_8904);
and U9547 (N_9547,N_8727,N_8817);
and U9548 (N_9548,N_8156,N_8511);
and U9549 (N_9549,N_8181,N_8147);
xnor U9550 (N_9550,N_8771,N_8067);
and U9551 (N_9551,N_8523,N_8111);
nor U9552 (N_9552,N_8329,N_8724);
xor U9553 (N_9553,N_8279,N_8739);
or U9554 (N_9554,N_8449,N_8196);
xnor U9555 (N_9555,N_8869,N_8989);
nor U9556 (N_9556,N_8202,N_8483);
nand U9557 (N_9557,N_8170,N_8742);
xnor U9558 (N_9558,N_8545,N_8298);
or U9559 (N_9559,N_8412,N_8758);
nor U9560 (N_9560,N_8395,N_8142);
xor U9561 (N_9561,N_8688,N_8877);
nor U9562 (N_9562,N_8004,N_8923);
nor U9563 (N_9563,N_8993,N_8669);
or U9564 (N_9564,N_8681,N_8773);
xor U9565 (N_9565,N_8123,N_8076);
nand U9566 (N_9566,N_8376,N_8080);
xor U9567 (N_9567,N_8668,N_8933);
or U9568 (N_9568,N_8065,N_8738);
nor U9569 (N_9569,N_8534,N_8174);
xor U9570 (N_9570,N_8622,N_8968);
nor U9571 (N_9571,N_8252,N_8933);
and U9572 (N_9572,N_8782,N_8292);
nand U9573 (N_9573,N_8545,N_8823);
nor U9574 (N_9574,N_8937,N_8163);
and U9575 (N_9575,N_8440,N_8961);
nand U9576 (N_9576,N_8904,N_8325);
and U9577 (N_9577,N_8147,N_8691);
and U9578 (N_9578,N_8956,N_8862);
nor U9579 (N_9579,N_8739,N_8696);
and U9580 (N_9580,N_8086,N_8779);
or U9581 (N_9581,N_8545,N_8111);
and U9582 (N_9582,N_8516,N_8007);
or U9583 (N_9583,N_8599,N_8343);
nor U9584 (N_9584,N_8757,N_8590);
nor U9585 (N_9585,N_8905,N_8075);
or U9586 (N_9586,N_8715,N_8023);
or U9587 (N_9587,N_8163,N_8578);
or U9588 (N_9588,N_8399,N_8935);
and U9589 (N_9589,N_8928,N_8743);
nand U9590 (N_9590,N_8435,N_8706);
nand U9591 (N_9591,N_8066,N_8400);
and U9592 (N_9592,N_8198,N_8957);
and U9593 (N_9593,N_8627,N_8803);
and U9594 (N_9594,N_8983,N_8710);
or U9595 (N_9595,N_8729,N_8270);
xnor U9596 (N_9596,N_8990,N_8161);
nor U9597 (N_9597,N_8020,N_8332);
nand U9598 (N_9598,N_8418,N_8200);
nand U9599 (N_9599,N_8981,N_8874);
xor U9600 (N_9600,N_8978,N_8773);
nor U9601 (N_9601,N_8181,N_8058);
nand U9602 (N_9602,N_8086,N_8126);
nand U9603 (N_9603,N_8164,N_8524);
xnor U9604 (N_9604,N_8144,N_8215);
nor U9605 (N_9605,N_8182,N_8191);
nand U9606 (N_9606,N_8438,N_8741);
or U9607 (N_9607,N_8331,N_8708);
and U9608 (N_9608,N_8420,N_8723);
or U9609 (N_9609,N_8807,N_8090);
xnor U9610 (N_9610,N_8091,N_8380);
or U9611 (N_9611,N_8821,N_8153);
xnor U9612 (N_9612,N_8099,N_8352);
or U9613 (N_9613,N_8451,N_8539);
or U9614 (N_9614,N_8339,N_8514);
xor U9615 (N_9615,N_8440,N_8350);
or U9616 (N_9616,N_8247,N_8174);
nand U9617 (N_9617,N_8543,N_8024);
nor U9618 (N_9618,N_8863,N_8545);
nor U9619 (N_9619,N_8697,N_8087);
nor U9620 (N_9620,N_8617,N_8429);
nor U9621 (N_9621,N_8443,N_8259);
and U9622 (N_9622,N_8429,N_8223);
or U9623 (N_9623,N_8233,N_8409);
or U9624 (N_9624,N_8521,N_8991);
nor U9625 (N_9625,N_8868,N_8562);
xor U9626 (N_9626,N_8357,N_8472);
or U9627 (N_9627,N_8535,N_8057);
xnor U9628 (N_9628,N_8669,N_8170);
and U9629 (N_9629,N_8464,N_8316);
nor U9630 (N_9630,N_8341,N_8469);
nor U9631 (N_9631,N_8687,N_8921);
nand U9632 (N_9632,N_8260,N_8485);
and U9633 (N_9633,N_8308,N_8497);
xor U9634 (N_9634,N_8364,N_8264);
nor U9635 (N_9635,N_8289,N_8575);
and U9636 (N_9636,N_8260,N_8820);
and U9637 (N_9637,N_8401,N_8260);
or U9638 (N_9638,N_8946,N_8348);
nand U9639 (N_9639,N_8986,N_8598);
nor U9640 (N_9640,N_8723,N_8653);
nor U9641 (N_9641,N_8780,N_8578);
nor U9642 (N_9642,N_8846,N_8798);
or U9643 (N_9643,N_8317,N_8464);
or U9644 (N_9644,N_8910,N_8689);
nor U9645 (N_9645,N_8872,N_8830);
xnor U9646 (N_9646,N_8605,N_8192);
xor U9647 (N_9647,N_8178,N_8980);
or U9648 (N_9648,N_8758,N_8247);
nor U9649 (N_9649,N_8953,N_8599);
or U9650 (N_9650,N_8067,N_8617);
and U9651 (N_9651,N_8340,N_8975);
xnor U9652 (N_9652,N_8974,N_8352);
nor U9653 (N_9653,N_8494,N_8239);
nor U9654 (N_9654,N_8976,N_8220);
xnor U9655 (N_9655,N_8832,N_8481);
nand U9656 (N_9656,N_8375,N_8165);
nand U9657 (N_9657,N_8115,N_8408);
nor U9658 (N_9658,N_8012,N_8388);
nor U9659 (N_9659,N_8561,N_8513);
nand U9660 (N_9660,N_8254,N_8649);
nand U9661 (N_9661,N_8901,N_8764);
nand U9662 (N_9662,N_8008,N_8980);
nor U9663 (N_9663,N_8711,N_8366);
nand U9664 (N_9664,N_8931,N_8872);
nor U9665 (N_9665,N_8525,N_8007);
xnor U9666 (N_9666,N_8517,N_8812);
nor U9667 (N_9667,N_8666,N_8436);
and U9668 (N_9668,N_8696,N_8142);
or U9669 (N_9669,N_8695,N_8338);
and U9670 (N_9670,N_8549,N_8727);
and U9671 (N_9671,N_8830,N_8661);
nor U9672 (N_9672,N_8133,N_8095);
nor U9673 (N_9673,N_8623,N_8663);
nand U9674 (N_9674,N_8350,N_8632);
and U9675 (N_9675,N_8589,N_8260);
and U9676 (N_9676,N_8312,N_8744);
or U9677 (N_9677,N_8967,N_8799);
xor U9678 (N_9678,N_8729,N_8179);
xor U9679 (N_9679,N_8922,N_8192);
xnor U9680 (N_9680,N_8029,N_8975);
nand U9681 (N_9681,N_8068,N_8495);
or U9682 (N_9682,N_8333,N_8923);
or U9683 (N_9683,N_8660,N_8455);
nand U9684 (N_9684,N_8125,N_8417);
and U9685 (N_9685,N_8757,N_8688);
and U9686 (N_9686,N_8840,N_8344);
xnor U9687 (N_9687,N_8548,N_8333);
and U9688 (N_9688,N_8083,N_8737);
nand U9689 (N_9689,N_8817,N_8919);
nor U9690 (N_9690,N_8768,N_8537);
and U9691 (N_9691,N_8529,N_8488);
xor U9692 (N_9692,N_8536,N_8720);
or U9693 (N_9693,N_8399,N_8388);
xor U9694 (N_9694,N_8755,N_8333);
or U9695 (N_9695,N_8989,N_8131);
nand U9696 (N_9696,N_8329,N_8692);
and U9697 (N_9697,N_8973,N_8833);
nor U9698 (N_9698,N_8266,N_8804);
nand U9699 (N_9699,N_8519,N_8023);
nand U9700 (N_9700,N_8105,N_8483);
and U9701 (N_9701,N_8703,N_8182);
nor U9702 (N_9702,N_8257,N_8439);
nand U9703 (N_9703,N_8485,N_8812);
and U9704 (N_9704,N_8900,N_8187);
xor U9705 (N_9705,N_8253,N_8807);
nand U9706 (N_9706,N_8212,N_8684);
xnor U9707 (N_9707,N_8677,N_8848);
nand U9708 (N_9708,N_8800,N_8859);
or U9709 (N_9709,N_8230,N_8108);
and U9710 (N_9710,N_8955,N_8575);
nand U9711 (N_9711,N_8477,N_8849);
and U9712 (N_9712,N_8370,N_8045);
nor U9713 (N_9713,N_8217,N_8278);
xnor U9714 (N_9714,N_8428,N_8510);
nand U9715 (N_9715,N_8868,N_8811);
nor U9716 (N_9716,N_8766,N_8350);
nor U9717 (N_9717,N_8447,N_8140);
nand U9718 (N_9718,N_8624,N_8736);
xnor U9719 (N_9719,N_8870,N_8856);
xnor U9720 (N_9720,N_8290,N_8940);
or U9721 (N_9721,N_8456,N_8442);
or U9722 (N_9722,N_8847,N_8468);
or U9723 (N_9723,N_8385,N_8191);
or U9724 (N_9724,N_8362,N_8484);
nand U9725 (N_9725,N_8611,N_8715);
or U9726 (N_9726,N_8663,N_8712);
and U9727 (N_9727,N_8330,N_8728);
or U9728 (N_9728,N_8745,N_8140);
nand U9729 (N_9729,N_8193,N_8439);
xor U9730 (N_9730,N_8393,N_8743);
xnor U9731 (N_9731,N_8651,N_8098);
or U9732 (N_9732,N_8780,N_8001);
or U9733 (N_9733,N_8085,N_8313);
and U9734 (N_9734,N_8718,N_8786);
nand U9735 (N_9735,N_8748,N_8624);
and U9736 (N_9736,N_8060,N_8325);
nor U9737 (N_9737,N_8844,N_8248);
xor U9738 (N_9738,N_8813,N_8382);
or U9739 (N_9739,N_8128,N_8067);
nor U9740 (N_9740,N_8992,N_8519);
nand U9741 (N_9741,N_8017,N_8495);
xor U9742 (N_9742,N_8230,N_8354);
and U9743 (N_9743,N_8378,N_8775);
and U9744 (N_9744,N_8565,N_8678);
and U9745 (N_9745,N_8051,N_8470);
xnor U9746 (N_9746,N_8000,N_8372);
nand U9747 (N_9747,N_8335,N_8228);
or U9748 (N_9748,N_8591,N_8909);
and U9749 (N_9749,N_8531,N_8437);
nor U9750 (N_9750,N_8940,N_8682);
xnor U9751 (N_9751,N_8614,N_8340);
nor U9752 (N_9752,N_8240,N_8254);
nand U9753 (N_9753,N_8418,N_8710);
xnor U9754 (N_9754,N_8440,N_8880);
nand U9755 (N_9755,N_8984,N_8964);
nor U9756 (N_9756,N_8401,N_8200);
xor U9757 (N_9757,N_8167,N_8081);
or U9758 (N_9758,N_8523,N_8285);
nor U9759 (N_9759,N_8110,N_8826);
and U9760 (N_9760,N_8688,N_8675);
nand U9761 (N_9761,N_8539,N_8368);
and U9762 (N_9762,N_8293,N_8003);
xor U9763 (N_9763,N_8370,N_8435);
nor U9764 (N_9764,N_8772,N_8785);
xnor U9765 (N_9765,N_8399,N_8517);
nor U9766 (N_9766,N_8398,N_8985);
and U9767 (N_9767,N_8494,N_8390);
and U9768 (N_9768,N_8829,N_8259);
or U9769 (N_9769,N_8258,N_8457);
nand U9770 (N_9770,N_8407,N_8674);
or U9771 (N_9771,N_8906,N_8709);
nand U9772 (N_9772,N_8533,N_8287);
and U9773 (N_9773,N_8336,N_8892);
nor U9774 (N_9774,N_8178,N_8253);
or U9775 (N_9775,N_8870,N_8007);
or U9776 (N_9776,N_8780,N_8596);
nand U9777 (N_9777,N_8896,N_8379);
or U9778 (N_9778,N_8424,N_8178);
or U9779 (N_9779,N_8171,N_8850);
or U9780 (N_9780,N_8611,N_8149);
and U9781 (N_9781,N_8045,N_8603);
xor U9782 (N_9782,N_8742,N_8654);
and U9783 (N_9783,N_8038,N_8503);
and U9784 (N_9784,N_8960,N_8528);
nor U9785 (N_9785,N_8240,N_8436);
nand U9786 (N_9786,N_8514,N_8358);
xor U9787 (N_9787,N_8962,N_8426);
or U9788 (N_9788,N_8652,N_8346);
nand U9789 (N_9789,N_8160,N_8313);
and U9790 (N_9790,N_8276,N_8507);
nand U9791 (N_9791,N_8095,N_8983);
xor U9792 (N_9792,N_8768,N_8193);
nand U9793 (N_9793,N_8326,N_8139);
and U9794 (N_9794,N_8067,N_8311);
nand U9795 (N_9795,N_8060,N_8824);
nand U9796 (N_9796,N_8054,N_8765);
and U9797 (N_9797,N_8792,N_8001);
xor U9798 (N_9798,N_8859,N_8592);
xnor U9799 (N_9799,N_8797,N_8181);
nor U9800 (N_9800,N_8218,N_8599);
nor U9801 (N_9801,N_8733,N_8163);
and U9802 (N_9802,N_8399,N_8942);
xnor U9803 (N_9803,N_8540,N_8629);
xor U9804 (N_9804,N_8613,N_8956);
nor U9805 (N_9805,N_8267,N_8183);
nand U9806 (N_9806,N_8994,N_8064);
nand U9807 (N_9807,N_8011,N_8787);
or U9808 (N_9808,N_8298,N_8543);
nor U9809 (N_9809,N_8840,N_8269);
nor U9810 (N_9810,N_8302,N_8322);
and U9811 (N_9811,N_8107,N_8677);
or U9812 (N_9812,N_8884,N_8657);
nor U9813 (N_9813,N_8336,N_8141);
or U9814 (N_9814,N_8714,N_8728);
and U9815 (N_9815,N_8461,N_8666);
and U9816 (N_9816,N_8765,N_8572);
or U9817 (N_9817,N_8097,N_8969);
and U9818 (N_9818,N_8821,N_8787);
nor U9819 (N_9819,N_8936,N_8546);
nor U9820 (N_9820,N_8279,N_8037);
xor U9821 (N_9821,N_8086,N_8011);
nor U9822 (N_9822,N_8786,N_8507);
xnor U9823 (N_9823,N_8777,N_8282);
and U9824 (N_9824,N_8512,N_8610);
nand U9825 (N_9825,N_8776,N_8068);
or U9826 (N_9826,N_8493,N_8182);
and U9827 (N_9827,N_8772,N_8122);
xnor U9828 (N_9828,N_8610,N_8191);
or U9829 (N_9829,N_8353,N_8587);
nand U9830 (N_9830,N_8790,N_8354);
xor U9831 (N_9831,N_8337,N_8734);
nand U9832 (N_9832,N_8609,N_8643);
or U9833 (N_9833,N_8030,N_8513);
nor U9834 (N_9834,N_8695,N_8588);
nand U9835 (N_9835,N_8893,N_8503);
and U9836 (N_9836,N_8764,N_8209);
or U9837 (N_9837,N_8842,N_8475);
nor U9838 (N_9838,N_8035,N_8536);
or U9839 (N_9839,N_8930,N_8184);
nand U9840 (N_9840,N_8369,N_8165);
or U9841 (N_9841,N_8815,N_8329);
nand U9842 (N_9842,N_8653,N_8572);
nand U9843 (N_9843,N_8758,N_8604);
nand U9844 (N_9844,N_8052,N_8698);
and U9845 (N_9845,N_8713,N_8157);
nor U9846 (N_9846,N_8406,N_8555);
or U9847 (N_9847,N_8775,N_8629);
xor U9848 (N_9848,N_8940,N_8838);
or U9849 (N_9849,N_8899,N_8728);
nand U9850 (N_9850,N_8464,N_8084);
nor U9851 (N_9851,N_8389,N_8666);
or U9852 (N_9852,N_8688,N_8822);
nor U9853 (N_9853,N_8977,N_8825);
xor U9854 (N_9854,N_8221,N_8375);
nor U9855 (N_9855,N_8591,N_8413);
nand U9856 (N_9856,N_8743,N_8029);
or U9857 (N_9857,N_8045,N_8945);
nor U9858 (N_9858,N_8164,N_8637);
or U9859 (N_9859,N_8026,N_8591);
nor U9860 (N_9860,N_8065,N_8552);
or U9861 (N_9861,N_8127,N_8060);
nor U9862 (N_9862,N_8817,N_8836);
xnor U9863 (N_9863,N_8338,N_8154);
nand U9864 (N_9864,N_8456,N_8065);
nand U9865 (N_9865,N_8011,N_8718);
or U9866 (N_9866,N_8570,N_8037);
and U9867 (N_9867,N_8155,N_8566);
nor U9868 (N_9868,N_8621,N_8006);
nand U9869 (N_9869,N_8780,N_8272);
and U9870 (N_9870,N_8576,N_8310);
and U9871 (N_9871,N_8019,N_8477);
xor U9872 (N_9872,N_8928,N_8669);
nor U9873 (N_9873,N_8055,N_8754);
nor U9874 (N_9874,N_8459,N_8791);
or U9875 (N_9875,N_8067,N_8081);
nor U9876 (N_9876,N_8118,N_8768);
nor U9877 (N_9877,N_8347,N_8396);
and U9878 (N_9878,N_8968,N_8412);
nor U9879 (N_9879,N_8923,N_8970);
nor U9880 (N_9880,N_8754,N_8953);
and U9881 (N_9881,N_8672,N_8485);
and U9882 (N_9882,N_8070,N_8654);
and U9883 (N_9883,N_8146,N_8035);
and U9884 (N_9884,N_8396,N_8981);
nor U9885 (N_9885,N_8325,N_8340);
nand U9886 (N_9886,N_8499,N_8925);
nor U9887 (N_9887,N_8339,N_8118);
nor U9888 (N_9888,N_8207,N_8520);
nor U9889 (N_9889,N_8625,N_8549);
and U9890 (N_9890,N_8529,N_8365);
xnor U9891 (N_9891,N_8772,N_8540);
nor U9892 (N_9892,N_8704,N_8323);
xnor U9893 (N_9893,N_8740,N_8202);
or U9894 (N_9894,N_8848,N_8051);
xor U9895 (N_9895,N_8960,N_8014);
xor U9896 (N_9896,N_8183,N_8418);
or U9897 (N_9897,N_8153,N_8869);
and U9898 (N_9898,N_8640,N_8208);
xnor U9899 (N_9899,N_8946,N_8029);
nand U9900 (N_9900,N_8479,N_8049);
xnor U9901 (N_9901,N_8747,N_8322);
or U9902 (N_9902,N_8874,N_8880);
nor U9903 (N_9903,N_8936,N_8946);
nand U9904 (N_9904,N_8562,N_8287);
nand U9905 (N_9905,N_8693,N_8567);
nor U9906 (N_9906,N_8502,N_8624);
and U9907 (N_9907,N_8777,N_8232);
xor U9908 (N_9908,N_8656,N_8659);
and U9909 (N_9909,N_8457,N_8060);
and U9910 (N_9910,N_8782,N_8748);
nand U9911 (N_9911,N_8942,N_8304);
or U9912 (N_9912,N_8329,N_8448);
nand U9913 (N_9913,N_8432,N_8998);
xor U9914 (N_9914,N_8070,N_8583);
nand U9915 (N_9915,N_8769,N_8132);
nor U9916 (N_9916,N_8561,N_8772);
xor U9917 (N_9917,N_8577,N_8135);
nor U9918 (N_9918,N_8443,N_8417);
nand U9919 (N_9919,N_8498,N_8149);
or U9920 (N_9920,N_8373,N_8311);
xnor U9921 (N_9921,N_8763,N_8037);
xnor U9922 (N_9922,N_8382,N_8795);
xnor U9923 (N_9923,N_8408,N_8466);
nand U9924 (N_9924,N_8843,N_8699);
nor U9925 (N_9925,N_8381,N_8021);
xnor U9926 (N_9926,N_8338,N_8314);
xor U9927 (N_9927,N_8774,N_8824);
or U9928 (N_9928,N_8414,N_8034);
nand U9929 (N_9929,N_8888,N_8643);
nor U9930 (N_9930,N_8019,N_8035);
nor U9931 (N_9931,N_8984,N_8624);
xnor U9932 (N_9932,N_8565,N_8773);
xnor U9933 (N_9933,N_8763,N_8284);
or U9934 (N_9934,N_8646,N_8443);
or U9935 (N_9935,N_8403,N_8949);
or U9936 (N_9936,N_8321,N_8765);
xor U9937 (N_9937,N_8473,N_8898);
nand U9938 (N_9938,N_8325,N_8291);
and U9939 (N_9939,N_8268,N_8997);
nand U9940 (N_9940,N_8297,N_8507);
or U9941 (N_9941,N_8535,N_8838);
nor U9942 (N_9942,N_8097,N_8999);
or U9943 (N_9943,N_8032,N_8995);
nor U9944 (N_9944,N_8346,N_8483);
and U9945 (N_9945,N_8194,N_8616);
or U9946 (N_9946,N_8334,N_8353);
xnor U9947 (N_9947,N_8368,N_8094);
or U9948 (N_9948,N_8121,N_8181);
or U9949 (N_9949,N_8726,N_8060);
and U9950 (N_9950,N_8110,N_8418);
and U9951 (N_9951,N_8597,N_8931);
nor U9952 (N_9952,N_8202,N_8749);
and U9953 (N_9953,N_8494,N_8560);
and U9954 (N_9954,N_8458,N_8894);
nand U9955 (N_9955,N_8239,N_8705);
nor U9956 (N_9956,N_8739,N_8197);
nor U9957 (N_9957,N_8782,N_8319);
xnor U9958 (N_9958,N_8585,N_8013);
xnor U9959 (N_9959,N_8507,N_8028);
nand U9960 (N_9960,N_8676,N_8781);
xnor U9961 (N_9961,N_8244,N_8274);
and U9962 (N_9962,N_8136,N_8864);
nand U9963 (N_9963,N_8699,N_8891);
nand U9964 (N_9964,N_8557,N_8133);
or U9965 (N_9965,N_8419,N_8735);
or U9966 (N_9966,N_8385,N_8050);
nor U9967 (N_9967,N_8341,N_8856);
xnor U9968 (N_9968,N_8171,N_8845);
or U9969 (N_9969,N_8977,N_8293);
xnor U9970 (N_9970,N_8173,N_8510);
nand U9971 (N_9971,N_8495,N_8833);
or U9972 (N_9972,N_8905,N_8740);
or U9973 (N_9973,N_8973,N_8904);
nor U9974 (N_9974,N_8287,N_8945);
xor U9975 (N_9975,N_8619,N_8392);
and U9976 (N_9976,N_8925,N_8895);
xnor U9977 (N_9977,N_8464,N_8761);
nor U9978 (N_9978,N_8457,N_8023);
nand U9979 (N_9979,N_8385,N_8293);
or U9980 (N_9980,N_8308,N_8026);
or U9981 (N_9981,N_8639,N_8276);
and U9982 (N_9982,N_8960,N_8555);
nand U9983 (N_9983,N_8649,N_8631);
nor U9984 (N_9984,N_8512,N_8698);
xnor U9985 (N_9985,N_8608,N_8254);
xor U9986 (N_9986,N_8952,N_8729);
nand U9987 (N_9987,N_8119,N_8428);
nand U9988 (N_9988,N_8177,N_8449);
and U9989 (N_9989,N_8519,N_8455);
or U9990 (N_9990,N_8053,N_8232);
and U9991 (N_9991,N_8394,N_8314);
xnor U9992 (N_9992,N_8938,N_8846);
nor U9993 (N_9993,N_8344,N_8547);
or U9994 (N_9994,N_8600,N_8516);
xnor U9995 (N_9995,N_8914,N_8847);
or U9996 (N_9996,N_8579,N_8563);
and U9997 (N_9997,N_8092,N_8683);
or U9998 (N_9998,N_8769,N_8398);
nand U9999 (N_9999,N_8932,N_8085);
xor U10000 (N_10000,N_9563,N_9216);
nand U10001 (N_10001,N_9496,N_9814);
nand U10002 (N_10002,N_9544,N_9253);
or U10003 (N_10003,N_9238,N_9324);
or U10004 (N_10004,N_9803,N_9381);
nand U10005 (N_10005,N_9375,N_9647);
nor U10006 (N_10006,N_9414,N_9602);
nand U10007 (N_10007,N_9157,N_9150);
xnor U10008 (N_10008,N_9540,N_9278);
nor U10009 (N_10009,N_9223,N_9861);
or U10010 (N_10010,N_9639,N_9985);
and U10011 (N_10011,N_9107,N_9329);
and U10012 (N_10012,N_9296,N_9227);
nor U10013 (N_10013,N_9973,N_9418);
and U10014 (N_10014,N_9705,N_9608);
nand U10015 (N_10015,N_9146,N_9117);
or U10016 (N_10016,N_9516,N_9443);
nor U10017 (N_10017,N_9979,N_9844);
nor U10018 (N_10018,N_9090,N_9987);
nand U10019 (N_10019,N_9636,N_9458);
xor U10020 (N_10020,N_9135,N_9561);
xor U10021 (N_10021,N_9908,N_9272);
nand U10022 (N_10022,N_9930,N_9522);
xor U10023 (N_10023,N_9752,N_9520);
nand U10024 (N_10024,N_9849,N_9420);
nor U10025 (N_10025,N_9954,N_9098);
and U10026 (N_10026,N_9269,N_9836);
nand U10027 (N_10027,N_9758,N_9975);
xnor U10028 (N_10028,N_9993,N_9548);
and U10029 (N_10029,N_9552,N_9620);
nor U10030 (N_10030,N_9457,N_9753);
or U10031 (N_10031,N_9615,N_9093);
nand U10032 (N_10032,N_9816,N_9601);
xnor U10033 (N_10033,N_9156,N_9184);
xor U10034 (N_10034,N_9404,N_9222);
and U10035 (N_10035,N_9197,N_9472);
nand U10036 (N_10036,N_9110,N_9890);
nand U10037 (N_10037,N_9568,N_9576);
nor U10038 (N_10038,N_9688,N_9124);
and U10039 (N_10039,N_9657,N_9668);
or U10040 (N_10040,N_9796,N_9815);
nor U10041 (N_10041,N_9410,N_9252);
and U10042 (N_10042,N_9046,N_9255);
nor U10043 (N_10043,N_9559,N_9043);
xor U10044 (N_10044,N_9052,N_9318);
or U10045 (N_10045,N_9773,N_9310);
nor U10046 (N_10046,N_9500,N_9995);
or U10047 (N_10047,N_9256,N_9512);
xor U10048 (N_10048,N_9190,N_9183);
nand U10049 (N_10049,N_9123,N_9536);
and U10050 (N_10050,N_9042,N_9679);
nor U10051 (N_10051,N_9630,N_9359);
or U10052 (N_10052,N_9943,N_9575);
and U10053 (N_10053,N_9888,N_9514);
xor U10054 (N_10054,N_9231,N_9365);
xor U10055 (N_10055,N_9170,N_9694);
nand U10056 (N_10056,N_9030,N_9645);
or U10057 (N_10057,N_9698,N_9840);
xor U10058 (N_10058,N_9392,N_9407);
xor U10059 (N_10059,N_9137,N_9994);
xnor U10060 (N_10060,N_9813,N_9573);
xnor U10061 (N_10061,N_9416,N_9703);
nor U10062 (N_10062,N_9887,N_9261);
nor U10063 (N_10063,N_9564,N_9185);
xnor U10064 (N_10064,N_9009,N_9940);
nand U10065 (N_10065,N_9293,N_9062);
nor U10066 (N_10066,N_9149,N_9907);
or U10067 (N_10067,N_9026,N_9785);
nor U10068 (N_10068,N_9933,N_9167);
nor U10069 (N_10069,N_9492,N_9367);
or U10070 (N_10070,N_9397,N_9160);
nor U10071 (N_10071,N_9951,N_9208);
xnor U10072 (N_10072,N_9068,N_9533);
and U10073 (N_10073,N_9812,N_9881);
nor U10074 (N_10074,N_9074,N_9133);
and U10075 (N_10075,N_9587,N_9205);
xor U10076 (N_10076,N_9154,N_9718);
xor U10077 (N_10077,N_9019,N_9724);
nand U10078 (N_10078,N_9398,N_9386);
nand U10079 (N_10079,N_9875,N_9424);
nor U10080 (N_10080,N_9323,N_9931);
or U10081 (N_10081,N_9733,N_9274);
xor U10082 (N_10082,N_9543,N_9012);
nand U10083 (N_10083,N_9715,N_9676);
xor U10084 (N_10084,N_9966,N_9389);
nand U10085 (N_10085,N_9851,N_9554);
xnor U10086 (N_10086,N_9437,N_9779);
nor U10087 (N_10087,N_9946,N_9749);
nand U10088 (N_10088,N_9339,N_9145);
or U10089 (N_10089,N_9142,N_9258);
nand U10090 (N_10090,N_9671,N_9164);
or U10091 (N_10091,N_9710,N_9672);
or U10092 (N_10092,N_9955,N_9203);
nand U10093 (N_10093,N_9104,N_9904);
or U10094 (N_10094,N_9945,N_9806);
nor U10095 (N_10095,N_9607,N_9736);
nand U10096 (N_10096,N_9936,N_9187);
xnor U10097 (N_10097,N_9596,N_9867);
and U10098 (N_10098,N_9342,N_9571);
xor U10099 (N_10099,N_9405,N_9096);
nand U10100 (N_10100,N_9592,N_9442);
xor U10101 (N_10101,N_9726,N_9474);
nand U10102 (N_10102,N_9388,N_9115);
nor U10103 (N_10103,N_9864,N_9447);
or U10104 (N_10104,N_9366,N_9619);
or U10105 (N_10105,N_9082,N_9807);
xor U10106 (N_10106,N_9532,N_9010);
nand U10107 (N_10107,N_9317,N_9834);
and U10108 (N_10108,N_9495,N_9210);
nor U10109 (N_10109,N_9067,N_9163);
nor U10110 (N_10110,N_9562,N_9605);
nand U10111 (N_10111,N_9949,N_9200);
nand U10112 (N_10112,N_9081,N_9111);
and U10113 (N_10113,N_9859,N_9958);
xnor U10114 (N_10114,N_9744,N_9413);
nor U10115 (N_10115,N_9644,N_9618);
and U10116 (N_10116,N_9105,N_9064);
xor U10117 (N_10117,N_9862,N_9920);
nand U10118 (N_10118,N_9285,N_9409);
nand U10119 (N_10119,N_9924,N_9557);
nor U10120 (N_10120,N_9700,N_9621);
or U10121 (N_10121,N_9266,N_9438);
nand U10122 (N_10122,N_9505,N_9417);
or U10123 (N_10123,N_9066,N_9423);
nand U10124 (N_10124,N_9327,N_9761);
nand U10125 (N_10125,N_9427,N_9631);
xnor U10126 (N_10126,N_9750,N_9182);
nor U10127 (N_10127,N_9034,N_9531);
xor U10128 (N_10128,N_9546,N_9013);
and U10129 (N_10129,N_9800,N_9101);
and U10130 (N_10130,N_9054,N_9383);
and U10131 (N_10131,N_9415,N_9534);
nand U10132 (N_10132,N_9787,N_9048);
or U10133 (N_10133,N_9884,N_9517);
and U10134 (N_10134,N_9590,N_9049);
nand U10135 (N_10135,N_9132,N_9060);
or U10136 (N_10136,N_9071,N_9569);
or U10137 (N_10137,N_9691,N_9574);
or U10138 (N_10138,N_9802,N_9250);
nor U10139 (N_10139,N_9330,N_9378);
nor U10140 (N_10140,N_9035,N_9848);
xor U10141 (N_10141,N_9612,N_9314);
and U10142 (N_10142,N_9411,N_9869);
nand U10143 (N_10143,N_9777,N_9856);
or U10144 (N_10144,N_9491,N_9391);
nor U10145 (N_10145,N_9380,N_9294);
or U10146 (N_10146,N_9600,N_9055);
and U10147 (N_10147,N_9088,N_9309);
or U10148 (N_10148,N_9739,N_9942);
xnor U10149 (N_10149,N_9482,N_9570);
nand U10150 (N_10150,N_9358,N_9229);
or U10151 (N_10151,N_9125,N_9089);
nor U10152 (N_10152,N_9905,N_9304);
or U10153 (N_10153,N_9284,N_9077);
xor U10154 (N_10154,N_9198,N_9501);
xor U10155 (N_10155,N_9696,N_9095);
nand U10156 (N_10156,N_9481,N_9738);
or U10157 (N_10157,N_9345,N_9390);
and U10158 (N_10158,N_9239,N_9820);
nand U10159 (N_10159,N_9640,N_9152);
nand U10160 (N_10160,N_9911,N_9159);
nand U10161 (N_10161,N_9504,N_9595);
nor U10162 (N_10162,N_9385,N_9537);
nor U10163 (N_10163,N_9650,N_9100);
and U10164 (N_10164,N_9850,N_9801);
xor U10165 (N_10165,N_9017,N_9045);
nand U10166 (N_10166,N_9527,N_9956);
and U10167 (N_10167,N_9332,N_9195);
nor U10168 (N_10168,N_9720,N_9259);
or U10169 (N_10169,N_9387,N_9161);
nand U10170 (N_10170,N_9106,N_9007);
or U10171 (N_10171,N_9031,N_9871);
nand U10172 (N_10172,N_9086,N_9439);
nand U10173 (N_10173,N_9033,N_9843);
nand U10174 (N_10174,N_9965,N_9232);
and U10175 (N_10175,N_9877,N_9153);
nor U10176 (N_10176,N_9245,N_9044);
nand U10177 (N_10177,N_9879,N_9246);
nand U10178 (N_10178,N_9690,N_9097);
or U10179 (N_10179,N_9996,N_9972);
nor U10180 (N_10180,N_9488,N_9586);
xnor U10181 (N_10181,N_9717,N_9662);
nor U10182 (N_10182,N_9889,N_9301);
and U10183 (N_10183,N_9058,N_9464);
or U10184 (N_10184,N_9742,N_9782);
nand U10185 (N_10185,N_9830,N_9057);
and U10186 (N_10186,N_9158,N_9363);
nor U10187 (N_10187,N_9654,N_9827);
nor U10188 (N_10188,N_9934,N_9992);
nor U10189 (N_10189,N_9661,N_9288);
or U10190 (N_10190,N_9968,N_9556);
xnor U10191 (N_10191,N_9845,N_9087);
nand U10192 (N_10192,N_9461,N_9050);
xor U10193 (N_10193,N_9355,N_9273);
xor U10194 (N_10194,N_9118,N_9311);
nor U10195 (N_10195,N_9865,N_9193);
nand U10196 (N_10196,N_9759,N_9876);
or U10197 (N_10197,N_9094,N_9240);
xor U10198 (N_10198,N_9673,N_9810);
xor U10199 (N_10199,N_9373,N_9823);
xnor U10200 (N_10200,N_9541,N_9664);
nand U10201 (N_10201,N_9073,N_9497);
and U10202 (N_10202,N_9213,N_9633);
and U10203 (N_10203,N_9912,N_9891);
nor U10204 (N_10204,N_9970,N_9914);
nand U10205 (N_10205,N_9950,N_9680);
or U10206 (N_10206,N_9333,N_9896);
or U10207 (N_10207,N_9990,N_9412);
nand U10208 (N_10208,N_9948,N_9999);
nand U10209 (N_10209,N_9938,N_9772);
and U10210 (N_10210,N_9670,N_9286);
nor U10211 (N_10211,N_9344,N_9446);
nand U10212 (N_10212,N_9766,N_9883);
xnor U10213 (N_10213,N_9341,N_9583);
or U10214 (N_10214,N_9741,N_9312);
or U10215 (N_10215,N_9658,N_9775);
and U10216 (N_10216,N_9632,N_9138);
xor U10217 (N_10217,N_9725,N_9530);
and U10218 (N_10218,N_9704,N_9141);
or U10219 (N_10219,N_9788,N_9895);
and U10220 (N_10220,N_9598,N_9277);
nand U10221 (N_10221,N_9635,N_9173);
nor U10222 (N_10222,N_9006,N_9393);
nor U10223 (N_10223,N_9892,N_9235);
nand U10224 (N_10224,N_9102,N_9751);
nor U10225 (N_10225,N_9027,N_9428);
nand U10226 (N_10226,N_9291,N_9131);
nor U10227 (N_10227,N_9490,N_9168);
xor U10228 (N_10228,N_9120,N_9747);
nor U10229 (N_10229,N_9578,N_9028);
and U10230 (N_10230,N_9832,N_9070);
and U10231 (N_10231,N_9178,N_9003);
nand U10232 (N_10232,N_9267,N_9307);
or U10233 (N_10233,N_9292,N_9456);
nor U10234 (N_10234,N_9244,N_9436);
and U10235 (N_10235,N_9722,N_9964);
nor U10236 (N_10236,N_9666,N_9901);
and U10237 (N_10237,N_9004,N_9254);
nor U10238 (N_10238,N_9024,N_9233);
nand U10239 (N_10239,N_9065,N_9727);
nor U10240 (N_10240,N_9511,N_9155);
or U10241 (N_10241,N_9900,N_9040);
xnor U10242 (N_10242,N_9171,N_9821);
nand U10243 (N_10243,N_9743,N_9368);
nor U10244 (N_10244,N_9280,N_9321);
or U10245 (N_10245,N_9984,N_9915);
and U10246 (N_10246,N_9475,N_9452);
and U10247 (N_10247,N_9289,N_9684);
nor U10248 (N_10248,N_9349,N_9053);
nor U10249 (N_10249,N_9455,N_9376);
and U10250 (N_10250,N_9708,N_9473);
nor U10251 (N_10251,N_9176,N_9029);
or U10252 (N_10252,N_9140,N_9435);
and U10253 (N_10253,N_9147,N_9963);
xor U10254 (N_10254,N_9909,N_9305);
and U10255 (N_10255,N_9212,N_9880);
or U10256 (N_10256,N_9480,N_9593);
or U10257 (N_10257,N_9509,N_9038);
or U10258 (N_10258,N_9112,N_9037);
nand U10259 (N_10259,N_9919,N_9025);
and U10260 (N_10260,N_9510,N_9370);
nor U10261 (N_10261,N_9144,N_9300);
xor U10262 (N_10262,N_9603,N_9271);
and U10263 (N_10263,N_9350,N_9989);
and U10264 (N_10264,N_9484,N_9737);
and U10265 (N_10265,N_9351,N_9174);
or U10266 (N_10266,N_9306,N_9776);
or U10267 (N_10267,N_9641,N_9263);
xnor U10268 (N_10268,N_9507,N_9822);
xnor U10269 (N_10269,N_9188,N_9594);
xnor U10270 (N_10270,N_9357,N_9316);
and U10271 (N_10271,N_9701,N_9652);
or U10272 (N_10272,N_9348,N_9937);
nor U10273 (N_10273,N_9426,N_9196);
nor U10274 (N_10274,N_9780,N_9218);
and U10275 (N_10275,N_9719,N_9281);
or U10276 (N_10276,N_9237,N_9275);
and U10277 (N_10277,N_9853,N_9921);
xnor U10278 (N_10278,N_9611,N_9697);
xnor U10279 (N_10279,N_9018,N_9331);
or U10280 (N_10280,N_9898,N_9078);
and U10281 (N_10281,N_9616,N_9448);
and U10282 (N_10282,N_9613,N_9005);
xnor U10283 (N_10283,N_9986,N_9328);
xnor U10284 (N_10284,N_9211,N_9186);
xnor U10285 (N_10285,N_9625,N_9394);
and U10286 (N_10286,N_9194,N_9846);
nand U10287 (N_10287,N_9799,N_9545);
nand U10288 (N_10288,N_9833,N_9916);
and U10289 (N_10289,N_9011,N_9525);
or U10290 (N_10290,N_9128,N_9885);
nand U10291 (N_10291,N_9765,N_9874);
or U10292 (N_10292,N_9922,N_9444);
and U10293 (N_10293,N_9714,N_9678);
or U10294 (N_10294,N_9695,N_9468);
nor U10295 (N_10295,N_9039,N_9347);
nor U10296 (N_10296,N_9648,N_9841);
and U10297 (N_10297,N_9872,N_9471);
nand U10298 (N_10298,N_9660,N_9935);
or U10299 (N_10299,N_9395,N_9466);
nor U10300 (N_10300,N_9108,N_9610);
or U10301 (N_10301,N_9109,N_9283);
and U10302 (N_10302,N_9224,N_9091);
or U10303 (N_10303,N_9083,N_9926);
nand U10304 (N_10304,N_9303,N_9508);
or U10305 (N_10305,N_9202,N_9981);
nor U10306 (N_10306,N_9798,N_9364);
nor U10307 (N_10307,N_9689,N_9629);
and U10308 (N_10308,N_9837,N_9623);
or U10309 (N_10309,N_9535,N_9489);
nand U10310 (N_10310,N_9234,N_9925);
and U10311 (N_10311,N_9831,N_9804);
nand U10312 (N_10312,N_9346,N_9265);
and U10313 (N_10313,N_9297,N_9002);
or U10314 (N_10314,N_9079,N_9817);
nor U10315 (N_10315,N_9783,N_9767);
nand U10316 (N_10316,N_9463,N_9971);
nand U10317 (N_10317,N_9923,N_9811);
xnor U10318 (N_10318,N_9264,N_9126);
xnor U10319 (N_10319,N_9624,N_9519);
xor U10320 (N_10320,N_9217,N_9433);
and U10321 (N_10321,N_9260,N_9702);
nor U10322 (N_10322,N_9276,N_9808);
nand U10323 (N_10323,N_9014,N_9236);
nor U10324 (N_10324,N_9771,N_9609);
nor U10325 (N_10325,N_9116,N_9939);
or U10326 (N_10326,N_9790,N_9962);
and U10327 (N_10327,N_9838,N_9215);
xnor U10328 (N_10328,N_9020,N_9361);
and U10329 (N_10329,N_9656,N_9477);
nand U10330 (N_10330,N_9228,N_9959);
and U10331 (N_10331,N_9099,N_9372);
xnor U10332 (N_10332,N_9494,N_9565);
or U10333 (N_10333,N_9084,N_9567);
and U10334 (N_10334,N_9542,N_9063);
or U10335 (N_10335,N_9952,N_9634);
nand U10336 (N_10336,N_9716,N_9795);
and U10337 (N_10337,N_9059,N_9980);
xnor U10338 (N_10338,N_9614,N_9745);
nor U10339 (N_10339,N_9659,N_9369);
and U10340 (N_10340,N_9655,N_9175);
xor U10341 (N_10341,N_9180,N_9918);
xnor U10342 (N_10342,N_9319,N_9022);
nor U10343 (N_10343,N_9762,N_9893);
or U10344 (N_10344,N_9498,N_9247);
xnor U10345 (N_10345,N_9001,N_9735);
and U10346 (N_10346,N_9356,N_9675);
xor U10347 (N_10347,N_9860,N_9431);
and U10348 (N_10348,N_9529,N_9421);
nor U10349 (N_10349,N_9041,N_9047);
or U10350 (N_10350,N_9910,N_9746);
and U10351 (N_10351,N_9169,N_9663);
nand U10352 (N_10352,N_9707,N_9023);
nand U10353 (N_10353,N_9682,N_9320);
nand U10354 (N_10354,N_9230,N_9826);
or U10355 (N_10355,N_9687,N_9335);
nand U10356 (N_10356,N_9969,N_9755);
xnor U10357 (N_10357,N_9401,N_9295);
nor U10358 (N_10358,N_9219,N_9402);
nor U10359 (N_10359,N_9786,N_9711);
nand U10360 (N_10360,N_9524,N_9549);
xnor U10361 (N_10361,N_9441,N_9399);
and U10362 (N_10362,N_9179,N_9374);
xnor U10363 (N_10363,N_9340,N_9419);
and U10364 (N_10364,N_9729,N_9878);
and U10365 (N_10365,N_9430,N_9051);
and U10366 (N_10366,N_9015,N_9226);
nor U10367 (N_10367,N_9677,N_9282);
and U10368 (N_10368,N_9906,N_9582);
and U10369 (N_10369,N_9917,N_9947);
or U10370 (N_10370,N_9539,N_9792);
and U10371 (N_10371,N_9432,N_9445);
nor U10372 (N_10372,N_9774,N_9201);
nand U10373 (N_10373,N_9852,N_9997);
or U10374 (N_10374,N_9204,N_9731);
or U10375 (N_10375,N_9768,N_9130);
xor U10376 (N_10376,N_9422,N_9449);
nor U10377 (N_10377,N_9287,N_9847);
nand U10378 (N_10378,N_9791,N_9839);
xnor U10379 (N_10379,N_9982,N_9903);
xor U10380 (N_10380,N_9462,N_9643);
and U10381 (N_10381,N_9858,N_9248);
or U10382 (N_10382,N_9406,N_9683);
nor U10383 (N_10383,N_9075,N_9740);
nand U10384 (N_10384,N_9486,N_9597);
and U10385 (N_10385,N_9523,N_9538);
xnor U10386 (N_10386,N_9470,N_9450);
and U10387 (N_10387,N_9998,N_9487);
or U10388 (N_10388,N_9882,N_9555);
nor U10389 (N_10389,N_9478,N_9249);
xor U10390 (N_10390,N_9870,N_9854);
and U10391 (N_10391,N_9585,N_9626);
or U10392 (N_10392,N_9604,N_9721);
and U10393 (N_10393,N_9957,N_9377);
nor U10394 (N_10394,N_9770,N_9809);
xor U10395 (N_10395,N_9521,N_9451);
xor U10396 (N_10396,N_9460,N_9166);
and U10397 (N_10397,N_9805,N_9638);
or U10398 (N_10398,N_9476,N_9894);
nand U10399 (N_10399,N_9941,N_9103);
xor U10400 (N_10400,N_9978,N_9262);
and U10401 (N_10401,N_9379,N_9192);
xor U10402 (N_10402,N_9789,N_9465);
or U10403 (N_10403,N_9976,N_9008);
or U10404 (N_10404,N_9313,N_9769);
nand U10405 (N_10405,N_9493,N_9325);
or U10406 (N_10406,N_9902,N_9960);
nor U10407 (N_10407,N_9579,N_9622);
or U10408 (N_10408,N_9967,N_9829);
xnor U10409 (N_10409,N_9828,N_9669);
nand U10410 (N_10410,N_9279,N_9617);
and U10411 (N_10411,N_9897,N_9114);
xnor U10412 (N_10412,N_9692,N_9572);
or U10413 (N_10413,N_9113,N_9085);
nand U10414 (N_10414,N_9693,N_9646);
nand U10415 (N_10415,N_9974,N_9151);
or U10416 (N_10416,N_9929,N_9360);
and U10417 (N_10417,N_9547,N_9453);
and U10418 (N_10418,N_9209,N_9651);
nor U10419 (N_10419,N_9396,N_9712);
xnor U10420 (N_10420,N_9553,N_9302);
and U10421 (N_10421,N_9032,N_9298);
xor U10422 (N_10422,N_9199,N_9136);
xnor U10423 (N_10423,N_9122,N_9299);
nand U10424 (N_10424,N_9076,N_9513);
xor U10425 (N_10425,N_9354,N_9400);
nor U10426 (N_10426,N_9092,N_9732);
xnor U10427 (N_10427,N_9763,N_9589);
nor U10428 (N_10428,N_9824,N_9754);
or U10429 (N_10429,N_9021,N_9384);
nand U10430 (N_10430,N_9842,N_9241);
and U10431 (N_10431,N_9251,N_9127);
xor U10432 (N_10432,N_9434,N_9866);
and U10433 (N_10433,N_9036,N_9818);
or U10434 (N_10434,N_9606,N_9080);
and U10435 (N_10435,N_9343,N_9953);
nand U10436 (N_10436,N_9000,N_9129);
xor U10437 (N_10437,N_9352,N_9526);
or U10438 (N_10438,N_9709,N_9528);
and U10439 (N_10439,N_9061,N_9584);
or U10440 (N_10440,N_9599,N_9873);
xor U10441 (N_10441,N_9778,N_9713);
nor U10442 (N_10442,N_9855,N_9121);
or U10443 (N_10443,N_9467,N_9886);
nand U10444 (N_10444,N_9913,N_9653);
or U10445 (N_10445,N_9148,N_9674);
and U10446 (N_10446,N_9483,N_9172);
nor U10447 (N_10447,N_9336,N_9685);
nor U10448 (N_10448,N_9991,N_9207);
nand U10449 (N_10449,N_9628,N_9242);
xor U10450 (N_10450,N_9334,N_9206);
and U10451 (N_10451,N_9485,N_9988);
and U10452 (N_10452,N_9337,N_9518);
xnor U10453 (N_10453,N_9764,N_9793);
or U10454 (N_10454,N_9560,N_9403);
xor U10455 (N_10455,N_9429,N_9756);
and U10456 (N_10456,N_9479,N_9191);
and U10457 (N_10457,N_9270,N_9723);
nand U10458 (N_10458,N_9225,N_9699);
nand U10459 (N_10459,N_9706,N_9667);
or U10460 (N_10460,N_9637,N_9863);
nor U10461 (N_10461,N_9425,N_9165);
nor U10462 (N_10462,N_9665,N_9797);
nand U10463 (N_10463,N_9835,N_9469);
nor U10464 (N_10464,N_9857,N_9515);
xor U10465 (N_10465,N_9499,N_9177);
and U10466 (N_10466,N_9730,N_9781);
xor U10467 (N_10467,N_9162,N_9440);
xor U10468 (N_10468,N_9214,N_9588);
nor U10469 (N_10469,N_9308,N_9757);
and U10470 (N_10470,N_9944,N_9566);
or U10471 (N_10471,N_9382,N_9642);
xor U10472 (N_10472,N_9134,N_9558);
nor U10473 (N_10473,N_9362,N_9649);
xnor U10474 (N_10474,N_9072,N_9220);
and U10475 (N_10475,N_9961,N_9069);
xnor U10476 (N_10476,N_9353,N_9825);
xor U10477 (N_10477,N_9794,N_9139);
xor U10478 (N_10478,N_9221,N_9243);
and U10479 (N_10479,N_9268,N_9728);
xnor U10480 (N_10480,N_9290,N_9459);
nand U10481 (N_10481,N_9580,N_9551);
xnor U10482 (N_10482,N_9326,N_9577);
or U10483 (N_10483,N_9371,N_9927);
nor U10484 (N_10484,N_9928,N_9143);
nor U10485 (N_10485,N_9581,N_9408);
nand U10486 (N_10486,N_9257,N_9016);
nor U10487 (N_10487,N_9932,N_9591);
or U10488 (N_10488,N_9734,N_9748);
nand U10489 (N_10489,N_9506,N_9454);
and U10490 (N_10490,N_9338,N_9627);
nor U10491 (N_10491,N_9056,N_9899);
xnor U10492 (N_10492,N_9315,N_9502);
or U10493 (N_10493,N_9681,N_9503);
or U10494 (N_10494,N_9686,N_9868);
nand U10495 (N_10495,N_9784,N_9977);
nor U10496 (N_10496,N_9760,N_9819);
or U10497 (N_10497,N_9119,N_9550);
xnor U10498 (N_10498,N_9189,N_9322);
nor U10499 (N_10499,N_9181,N_9983);
nor U10500 (N_10500,N_9361,N_9829);
and U10501 (N_10501,N_9865,N_9257);
xor U10502 (N_10502,N_9889,N_9270);
nand U10503 (N_10503,N_9707,N_9109);
and U10504 (N_10504,N_9483,N_9890);
xor U10505 (N_10505,N_9269,N_9689);
xnor U10506 (N_10506,N_9769,N_9187);
nor U10507 (N_10507,N_9860,N_9960);
and U10508 (N_10508,N_9012,N_9104);
and U10509 (N_10509,N_9666,N_9909);
or U10510 (N_10510,N_9567,N_9918);
nor U10511 (N_10511,N_9346,N_9577);
nor U10512 (N_10512,N_9582,N_9936);
and U10513 (N_10513,N_9740,N_9564);
xnor U10514 (N_10514,N_9921,N_9183);
nand U10515 (N_10515,N_9345,N_9185);
or U10516 (N_10516,N_9397,N_9522);
or U10517 (N_10517,N_9453,N_9195);
and U10518 (N_10518,N_9246,N_9848);
and U10519 (N_10519,N_9691,N_9682);
or U10520 (N_10520,N_9847,N_9874);
nand U10521 (N_10521,N_9620,N_9534);
xnor U10522 (N_10522,N_9096,N_9480);
nand U10523 (N_10523,N_9079,N_9690);
or U10524 (N_10524,N_9099,N_9777);
nor U10525 (N_10525,N_9273,N_9667);
nor U10526 (N_10526,N_9795,N_9744);
or U10527 (N_10527,N_9987,N_9736);
nand U10528 (N_10528,N_9304,N_9675);
or U10529 (N_10529,N_9656,N_9133);
xor U10530 (N_10530,N_9376,N_9812);
nand U10531 (N_10531,N_9368,N_9033);
and U10532 (N_10532,N_9738,N_9833);
or U10533 (N_10533,N_9767,N_9195);
and U10534 (N_10534,N_9285,N_9191);
nor U10535 (N_10535,N_9120,N_9663);
nand U10536 (N_10536,N_9525,N_9394);
or U10537 (N_10537,N_9713,N_9368);
or U10538 (N_10538,N_9685,N_9508);
nand U10539 (N_10539,N_9645,N_9418);
or U10540 (N_10540,N_9132,N_9834);
nor U10541 (N_10541,N_9333,N_9862);
or U10542 (N_10542,N_9644,N_9621);
xor U10543 (N_10543,N_9906,N_9096);
xor U10544 (N_10544,N_9412,N_9676);
nor U10545 (N_10545,N_9104,N_9841);
nand U10546 (N_10546,N_9309,N_9583);
nand U10547 (N_10547,N_9261,N_9577);
or U10548 (N_10548,N_9471,N_9708);
or U10549 (N_10549,N_9467,N_9737);
nand U10550 (N_10550,N_9057,N_9214);
and U10551 (N_10551,N_9036,N_9561);
xnor U10552 (N_10552,N_9970,N_9614);
nor U10553 (N_10553,N_9703,N_9896);
nand U10554 (N_10554,N_9304,N_9929);
nand U10555 (N_10555,N_9053,N_9785);
and U10556 (N_10556,N_9581,N_9450);
nand U10557 (N_10557,N_9363,N_9198);
and U10558 (N_10558,N_9190,N_9734);
or U10559 (N_10559,N_9434,N_9457);
xor U10560 (N_10560,N_9181,N_9312);
xnor U10561 (N_10561,N_9959,N_9353);
xnor U10562 (N_10562,N_9701,N_9019);
or U10563 (N_10563,N_9794,N_9541);
and U10564 (N_10564,N_9117,N_9296);
nand U10565 (N_10565,N_9000,N_9628);
or U10566 (N_10566,N_9558,N_9570);
and U10567 (N_10567,N_9282,N_9237);
nor U10568 (N_10568,N_9470,N_9405);
nor U10569 (N_10569,N_9411,N_9317);
nor U10570 (N_10570,N_9182,N_9062);
xor U10571 (N_10571,N_9366,N_9306);
xor U10572 (N_10572,N_9703,N_9254);
or U10573 (N_10573,N_9709,N_9193);
nor U10574 (N_10574,N_9498,N_9508);
or U10575 (N_10575,N_9633,N_9001);
and U10576 (N_10576,N_9939,N_9515);
nand U10577 (N_10577,N_9642,N_9134);
nor U10578 (N_10578,N_9383,N_9248);
or U10579 (N_10579,N_9673,N_9657);
xor U10580 (N_10580,N_9202,N_9283);
xnor U10581 (N_10581,N_9698,N_9873);
xor U10582 (N_10582,N_9686,N_9761);
or U10583 (N_10583,N_9037,N_9161);
nand U10584 (N_10584,N_9031,N_9646);
or U10585 (N_10585,N_9449,N_9660);
and U10586 (N_10586,N_9932,N_9808);
and U10587 (N_10587,N_9240,N_9578);
nand U10588 (N_10588,N_9784,N_9674);
and U10589 (N_10589,N_9962,N_9147);
nand U10590 (N_10590,N_9932,N_9229);
or U10591 (N_10591,N_9224,N_9545);
and U10592 (N_10592,N_9778,N_9226);
and U10593 (N_10593,N_9741,N_9255);
nor U10594 (N_10594,N_9037,N_9046);
or U10595 (N_10595,N_9322,N_9068);
nor U10596 (N_10596,N_9496,N_9934);
nand U10597 (N_10597,N_9529,N_9479);
xor U10598 (N_10598,N_9100,N_9131);
xnor U10599 (N_10599,N_9747,N_9323);
xor U10600 (N_10600,N_9482,N_9830);
and U10601 (N_10601,N_9213,N_9362);
and U10602 (N_10602,N_9068,N_9345);
xnor U10603 (N_10603,N_9071,N_9375);
or U10604 (N_10604,N_9242,N_9339);
or U10605 (N_10605,N_9661,N_9837);
nor U10606 (N_10606,N_9943,N_9053);
xnor U10607 (N_10607,N_9154,N_9700);
nand U10608 (N_10608,N_9900,N_9782);
and U10609 (N_10609,N_9032,N_9841);
nand U10610 (N_10610,N_9984,N_9657);
xnor U10611 (N_10611,N_9213,N_9684);
xor U10612 (N_10612,N_9711,N_9234);
nand U10613 (N_10613,N_9723,N_9359);
or U10614 (N_10614,N_9981,N_9982);
or U10615 (N_10615,N_9093,N_9672);
or U10616 (N_10616,N_9345,N_9516);
or U10617 (N_10617,N_9131,N_9463);
xnor U10618 (N_10618,N_9054,N_9640);
nor U10619 (N_10619,N_9692,N_9082);
nand U10620 (N_10620,N_9447,N_9386);
or U10621 (N_10621,N_9277,N_9629);
or U10622 (N_10622,N_9598,N_9312);
and U10623 (N_10623,N_9503,N_9261);
nor U10624 (N_10624,N_9253,N_9454);
xor U10625 (N_10625,N_9934,N_9117);
and U10626 (N_10626,N_9479,N_9579);
or U10627 (N_10627,N_9695,N_9771);
or U10628 (N_10628,N_9968,N_9496);
nand U10629 (N_10629,N_9915,N_9081);
and U10630 (N_10630,N_9633,N_9568);
and U10631 (N_10631,N_9671,N_9455);
or U10632 (N_10632,N_9579,N_9366);
nor U10633 (N_10633,N_9814,N_9248);
xor U10634 (N_10634,N_9498,N_9195);
nor U10635 (N_10635,N_9456,N_9525);
or U10636 (N_10636,N_9622,N_9070);
nor U10637 (N_10637,N_9725,N_9589);
xnor U10638 (N_10638,N_9358,N_9013);
or U10639 (N_10639,N_9072,N_9515);
and U10640 (N_10640,N_9058,N_9554);
and U10641 (N_10641,N_9145,N_9371);
and U10642 (N_10642,N_9672,N_9630);
or U10643 (N_10643,N_9875,N_9190);
nand U10644 (N_10644,N_9895,N_9768);
xor U10645 (N_10645,N_9995,N_9603);
and U10646 (N_10646,N_9904,N_9327);
nand U10647 (N_10647,N_9283,N_9323);
and U10648 (N_10648,N_9068,N_9264);
nor U10649 (N_10649,N_9127,N_9808);
xor U10650 (N_10650,N_9878,N_9774);
nand U10651 (N_10651,N_9303,N_9668);
xor U10652 (N_10652,N_9034,N_9508);
nor U10653 (N_10653,N_9375,N_9202);
xor U10654 (N_10654,N_9403,N_9217);
nor U10655 (N_10655,N_9641,N_9851);
and U10656 (N_10656,N_9617,N_9310);
and U10657 (N_10657,N_9600,N_9404);
xor U10658 (N_10658,N_9088,N_9649);
xnor U10659 (N_10659,N_9627,N_9846);
nand U10660 (N_10660,N_9937,N_9328);
xor U10661 (N_10661,N_9232,N_9823);
xnor U10662 (N_10662,N_9584,N_9063);
and U10663 (N_10663,N_9489,N_9669);
nor U10664 (N_10664,N_9916,N_9095);
and U10665 (N_10665,N_9155,N_9911);
xnor U10666 (N_10666,N_9467,N_9572);
and U10667 (N_10667,N_9893,N_9456);
nand U10668 (N_10668,N_9107,N_9379);
xor U10669 (N_10669,N_9844,N_9059);
nand U10670 (N_10670,N_9608,N_9875);
and U10671 (N_10671,N_9480,N_9713);
nand U10672 (N_10672,N_9293,N_9291);
nor U10673 (N_10673,N_9903,N_9272);
or U10674 (N_10674,N_9663,N_9714);
nand U10675 (N_10675,N_9642,N_9324);
xnor U10676 (N_10676,N_9583,N_9278);
or U10677 (N_10677,N_9545,N_9783);
or U10678 (N_10678,N_9072,N_9849);
or U10679 (N_10679,N_9773,N_9415);
nor U10680 (N_10680,N_9775,N_9705);
or U10681 (N_10681,N_9187,N_9734);
xnor U10682 (N_10682,N_9083,N_9811);
nor U10683 (N_10683,N_9073,N_9508);
nor U10684 (N_10684,N_9493,N_9781);
and U10685 (N_10685,N_9172,N_9624);
and U10686 (N_10686,N_9905,N_9005);
nand U10687 (N_10687,N_9073,N_9486);
or U10688 (N_10688,N_9540,N_9852);
or U10689 (N_10689,N_9613,N_9509);
nand U10690 (N_10690,N_9854,N_9431);
xnor U10691 (N_10691,N_9572,N_9596);
xor U10692 (N_10692,N_9833,N_9084);
xnor U10693 (N_10693,N_9316,N_9452);
nand U10694 (N_10694,N_9559,N_9922);
xnor U10695 (N_10695,N_9052,N_9642);
nor U10696 (N_10696,N_9912,N_9587);
nor U10697 (N_10697,N_9251,N_9125);
xnor U10698 (N_10698,N_9173,N_9777);
or U10699 (N_10699,N_9646,N_9665);
xor U10700 (N_10700,N_9118,N_9240);
nor U10701 (N_10701,N_9065,N_9774);
xor U10702 (N_10702,N_9279,N_9674);
nand U10703 (N_10703,N_9990,N_9938);
nand U10704 (N_10704,N_9985,N_9781);
or U10705 (N_10705,N_9790,N_9297);
nand U10706 (N_10706,N_9293,N_9972);
nand U10707 (N_10707,N_9803,N_9608);
xor U10708 (N_10708,N_9876,N_9713);
nor U10709 (N_10709,N_9249,N_9971);
nor U10710 (N_10710,N_9684,N_9329);
and U10711 (N_10711,N_9630,N_9758);
xnor U10712 (N_10712,N_9256,N_9868);
xnor U10713 (N_10713,N_9236,N_9700);
or U10714 (N_10714,N_9545,N_9803);
nand U10715 (N_10715,N_9529,N_9778);
nand U10716 (N_10716,N_9302,N_9242);
nand U10717 (N_10717,N_9018,N_9713);
and U10718 (N_10718,N_9933,N_9130);
xor U10719 (N_10719,N_9418,N_9996);
or U10720 (N_10720,N_9860,N_9848);
nor U10721 (N_10721,N_9342,N_9407);
or U10722 (N_10722,N_9147,N_9505);
nand U10723 (N_10723,N_9982,N_9775);
or U10724 (N_10724,N_9219,N_9192);
nand U10725 (N_10725,N_9231,N_9369);
xnor U10726 (N_10726,N_9313,N_9527);
nand U10727 (N_10727,N_9909,N_9280);
nor U10728 (N_10728,N_9807,N_9972);
xor U10729 (N_10729,N_9250,N_9654);
or U10730 (N_10730,N_9411,N_9600);
or U10731 (N_10731,N_9833,N_9279);
nor U10732 (N_10732,N_9433,N_9794);
nand U10733 (N_10733,N_9750,N_9463);
xnor U10734 (N_10734,N_9918,N_9887);
and U10735 (N_10735,N_9153,N_9680);
nand U10736 (N_10736,N_9611,N_9287);
nor U10737 (N_10737,N_9918,N_9230);
nor U10738 (N_10738,N_9689,N_9135);
nor U10739 (N_10739,N_9970,N_9552);
nor U10740 (N_10740,N_9748,N_9252);
nand U10741 (N_10741,N_9226,N_9784);
or U10742 (N_10742,N_9935,N_9828);
or U10743 (N_10743,N_9337,N_9014);
nand U10744 (N_10744,N_9691,N_9594);
nor U10745 (N_10745,N_9399,N_9818);
nand U10746 (N_10746,N_9317,N_9944);
and U10747 (N_10747,N_9556,N_9264);
nand U10748 (N_10748,N_9075,N_9475);
nand U10749 (N_10749,N_9884,N_9738);
and U10750 (N_10750,N_9721,N_9755);
xnor U10751 (N_10751,N_9607,N_9472);
nand U10752 (N_10752,N_9617,N_9794);
xor U10753 (N_10753,N_9098,N_9155);
nand U10754 (N_10754,N_9456,N_9887);
nor U10755 (N_10755,N_9663,N_9415);
and U10756 (N_10756,N_9877,N_9053);
or U10757 (N_10757,N_9514,N_9636);
or U10758 (N_10758,N_9784,N_9571);
xor U10759 (N_10759,N_9904,N_9840);
or U10760 (N_10760,N_9827,N_9527);
or U10761 (N_10761,N_9240,N_9386);
or U10762 (N_10762,N_9014,N_9587);
nor U10763 (N_10763,N_9121,N_9148);
xnor U10764 (N_10764,N_9617,N_9168);
nor U10765 (N_10765,N_9468,N_9220);
xor U10766 (N_10766,N_9458,N_9493);
nand U10767 (N_10767,N_9773,N_9214);
and U10768 (N_10768,N_9747,N_9339);
and U10769 (N_10769,N_9717,N_9675);
or U10770 (N_10770,N_9380,N_9560);
nand U10771 (N_10771,N_9155,N_9730);
xor U10772 (N_10772,N_9765,N_9141);
and U10773 (N_10773,N_9236,N_9113);
xor U10774 (N_10774,N_9961,N_9678);
nor U10775 (N_10775,N_9465,N_9023);
nor U10776 (N_10776,N_9359,N_9580);
and U10777 (N_10777,N_9110,N_9402);
and U10778 (N_10778,N_9359,N_9026);
nand U10779 (N_10779,N_9305,N_9452);
nand U10780 (N_10780,N_9730,N_9613);
and U10781 (N_10781,N_9327,N_9070);
xnor U10782 (N_10782,N_9701,N_9427);
nand U10783 (N_10783,N_9879,N_9179);
and U10784 (N_10784,N_9948,N_9846);
xnor U10785 (N_10785,N_9799,N_9066);
or U10786 (N_10786,N_9650,N_9065);
and U10787 (N_10787,N_9588,N_9745);
nand U10788 (N_10788,N_9036,N_9944);
or U10789 (N_10789,N_9771,N_9735);
nor U10790 (N_10790,N_9623,N_9278);
and U10791 (N_10791,N_9691,N_9229);
nor U10792 (N_10792,N_9377,N_9588);
xnor U10793 (N_10793,N_9016,N_9080);
and U10794 (N_10794,N_9527,N_9973);
or U10795 (N_10795,N_9194,N_9436);
or U10796 (N_10796,N_9155,N_9179);
and U10797 (N_10797,N_9878,N_9152);
and U10798 (N_10798,N_9406,N_9257);
or U10799 (N_10799,N_9577,N_9625);
or U10800 (N_10800,N_9908,N_9898);
xnor U10801 (N_10801,N_9174,N_9877);
xnor U10802 (N_10802,N_9223,N_9051);
nand U10803 (N_10803,N_9785,N_9364);
nor U10804 (N_10804,N_9425,N_9233);
nand U10805 (N_10805,N_9003,N_9597);
and U10806 (N_10806,N_9233,N_9331);
or U10807 (N_10807,N_9415,N_9935);
nand U10808 (N_10808,N_9260,N_9169);
or U10809 (N_10809,N_9960,N_9818);
or U10810 (N_10810,N_9032,N_9371);
or U10811 (N_10811,N_9367,N_9277);
xnor U10812 (N_10812,N_9319,N_9229);
xor U10813 (N_10813,N_9080,N_9181);
or U10814 (N_10814,N_9081,N_9182);
xnor U10815 (N_10815,N_9722,N_9580);
or U10816 (N_10816,N_9279,N_9085);
xnor U10817 (N_10817,N_9920,N_9706);
and U10818 (N_10818,N_9115,N_9295);
and U10819 (N_10819,N_9992,N_9307);
xor U10820 (N_10820,N_9199,N_9066);
and U10821 (N_10821,N_9821,N_9686);
and U10822 (N_10822,N_9152,N_9642);
nor U10823 (N_10823,N_9814,N_9927);
nor U10824 (N_10824,N_9990,N_9124);
nand U10825 (N_10825,N_9479,N_9716);
or U10826 (N_10826,N_9498,N_9136);
or U10827 (N_10827,N_9971,N_9224);
and U10828 (N_10828,N_9603,N_9397);
or U10829 (N_10829,N_9670,N_9651);
nand U10830 (N_10830,N_9394,N_9819);
and U10831 (N_10831,N_9047,N_9879);
and U10832 (N_10832,N_9949,N_9722);
or U10833 (N_10833,N_9164,N_9085);
and U10834 (N_10834,N_9633,N_9650);
xor U10835 (N_10835,N_9625,N_9671);
nand U10836 (N_10836,N_9370,N_9066);
and U10837 (N_10837,N_9976,N_9947);
xnor U10838 (N_10838,N_9364,N_9862);
nand U10839 (N_10839,N_9822,N_9062);
or U10840 (N_10840,N_9686,N_9006);
or U10841 (N_10841,N_9879,N_9146);
nor U10842 (N_10842,N_9644,N_9154);
xnor U10843 (N_10843,N_9309,N_9027);
nor U10844 (N_10844,N_9214,N_9131);
or U10845 (N_10845,N_9858,N_9759);
xor U10846 (N_10846,N_9872,N_9498);
and U10847 (N_10847,N_9206,N_9649);
nor U10848 (N_10848,N_9198,N_9188);
nand U10849 (N_10849,N_9449,N_9706);
nand U10850 (N_10850,N_9780,N_9478);
and U10851 (N_10851,N_9015,N_9496);
or U10852 (N_10852,N_9988,N_9459);
or U10853 (N_10853,N_9080,N_9136);
or U10854 (N_10854,N_9669,N_9990);
and U10855 (N_10855,N_9258,N_9299);
nor U10856 (N_10856,N_9884,N_9174);
and U10857 (N_10857,N_9704,N_9092);
and U10858 (N_10858,N_9125,N_9970);
nor U10859 (N_10859,N_9771,N_9051);
or U10860 (N_10860,N_9449,N_9527);
xor U10861 (N_10861,N_9959,N_9272);
or U10862 (N_10862,N_9667,N_9438);
or U10863 (N_10863,N_9826,N_9895);
or U10864 (N_10864,N_9367,N_9546);
or U10865 (N_10865,N_9634,N_9414);
xor U10866 (N_10866,N_9913,N_9662);
and U10867 (N_10867,N_9777,N_9049);
xor U10868 (N_10868,N_9701,N_9194);
and U10869 (N_10869,N_9415,N_9130);
nand U10870 (N_10870,N_9262,N_9695);
nor U10871 (N_10871,N_9442,N_9556);
xor U10872 (N_10872,N_9315,N_9354);
nand U10873 (N_10873,N_9909,N_9579);
and U10874 (N_10874,N_9783,N_9184);
xnor U10875 (N_10875,N_9156,N_9816);
nand U10876 (N_10876,N_9479,N_9655);
or U10877 (N_10877,N_9689,N_9396);
or U10878 (N_10878,N_9502,N_9513);
nand U10879 (N_10879,N_9614,N_9317);
nand U10880 (N_10880,N_9720,N_9308);
or U10881 (N_10881,N_9112,N_9931);
xor U10882 (N_10882,N_9865,N_9445);
nand U10883 (N_10883,N_9423,N_9614);
nor U10884 (N_10884,N_9455,N_9766);
nand U10885 (N_10885,N_9741,N_9033);
or U10886 (N_10886,N_9398,N_9618);
nor U10887 (N_10887,N_9037,N_9964);
nand U10888 (N_10888,N_9079,N_9062);
xor U10889 (N_10889,N_9315,N_9622);
and U10890 (N_10890,N_9809,N_9078);
nor U10891 (N_10891,N_9867,N_9572);
xor U10892 (N_10892,N_9947,N_9636);
and U10893 (N_10893,N_9769,N_9726);
nor U10894 (N_10894,N_9783,N_9428);
nand U10895 (N_10895,N_9969,N_9135);
xnor U10896 (N_10896,N_9488,N_9622);
nand U10897 (N_10897,N_9198,N_9884);
nand U10898 (N_10898,N_9190,N_9630);
nand U10899 (N_10899,N_9997,N_9008);
or U10900 (N_10900,N_9914,N_9896);
xor U10901 (N_10901,N_9036,N_9298);
or U10902 (N_10902,N_9309,N_9632);
and U10903 (N_10903,N_9387,N_9206);
nand U10904 (N_10904,N_9113,N_9300);
or U10905 (N_10905,N_9761,N_9499);
or U10906 (N_10906,N_9792,N_9490);
nor U10907 (N_10907,N_9612,N_9823);
and U10908 (N_10908,N_9402,N_9531);
xnor U10909 (N_10909,N_9086,N_9565);
nand U10910 (N_10910,N_9344,N_9923);
xnor U10911 (N_10911,N_9251,N_9457);
or U10912 (N_10912,N_9684,N_9956);
and U10913 (N_10913,N_9965,N_9564);
and U10914 (N_10914,N_9373,N_9304);
or U10915 (N_10915,N_9365,N_9753);
nor U10916 (N_10916,N_9022,N_9602);
and U10917 (N_10917,N_9375,N_9775);
and U10918 (N_10918,N_9677,N_9373);
or U10919 (N_10919,N_9829,N_9596);
xor U10920 (N_10920,N_9580,N_9092);
nor U10921 (N_10921,N_9670,N_9366);
and U10922 (N_10922,N_9096,N_9771);
xnor U10923 (N_10923,N_9996,N_9441);
xor U10924 (N_10924,N_9047,N_9368);
nor U10925 (N_10925,N_9158,N_9201);
and U10926 (N_10926,N_9649,N_9814);
nand U10927 (N_10927,N_9688,N_9919);
xor U10928 (N_10928,N_9672,N_9170);
or U10929 (N_10929,N_9574,N_9990);
nor U10930 (N_10930,N_9571,N_9455);
nand U10931 (N_10931,N_9750,N_9325);
nand U10932 (N_10932,N_9302,N_9230);
or U10933 (N_10933,N_9813,N_9315);
xor U10934 (N_10934,N_9576,N_9777);
and U10935 (N_10935,N_9271,N_9210);
or U10936 (N_10936,N_9311,N_9379);
nand U10937 (N_10937,N_9438,N_9101);
nor U10938 (N_10938,N_9202,N_9820);
and U10939 (N_10939,N_9152,N_9619);
nor U10940 (N_10940,N_9871,N_9940);
nor U10941 (N_10941,N_9303,N_9138);
xor U10942 (N_10942,N_9114,N_9862);
and U10943 (N_10943,N_9031,N_9954);
nor U10944 (N_10944,N_9084,N_9351);
or U10945 (N_10945,N_9044,N_9648);
or U10946 (N_10946,N_9226,N_9844);
or U10947 (N_10947,N_9858,N_9468);
and U10948 (N_10948,N_9872,N_9214);
nor U10949 (N_10949,N_9994,N_9975);
nor U10950 (N_10950,N_9466,N_9875);
nand U10951 (N_10951,N_9725,N_9417);
nand U10952 (N_10952,N_9664,N_9608);
or U10953 (N_10953,N_9133,N_9786);
nor U10954 (N_10954,N_9923,N_9468);
nand U10955 (N_10955,N_9580,N_9382);
and U10956 (N_10956,N_9228,N_9602);
or U10957 (N_10957,N_9047,N_9737);
or U10958 (N_10958,N_9771,N_9404);
xor U10959 (N_10959,N_9178,N_9181);
and U10960 (N_10960,N_9795,N_9568);
nand U10961 (N_10961,N_9877,N_9582);
xnor U10962 (N_10962,N_9749,N_9456);
nand U10963 (N_10963,N_9226,N_9008);
nor U10964 (N_10964,N_9366,N_9255);
or U10965 (N_10965,N_9770,N_9305);
or U10966 (N_10966,N_9179,N_9199);
nand U10967 (N_10967,N_9293,N_9342);
xnor U10968 (N_10968,N_9530,N_9939);
and U10969 (N_10969,N_9674,N_9499);
xor U10970 (N_10970,N_9418,N_9861);
xnor U10971 (N_10971,N_9502,N_9344);
nand U10972 (N_10972,N_9754,N_9745);
nor U10973 (N_10973,N_9853,N_9550);
xor U10974 (N_10974,N_9718,N_9171);
and U10975 (N_10975,N_9606,N_9288);
or U10976 (N_10976,N_9173,N_9773);
xor U10977 (N_10977,N_9576,N_9242);
nor U10978 (N_10978,N_9859,N_9122);
and U10979 (N_10979,N_9818,N_9770);
and U10980 (N_10980,N_9779,N_9962);
xnor U10981 (N_10981,N_9535,N_9842);
and U10982 (N_10982,N_9247,N_9659);
nand U10983 (N_10983,N_9650,N_9698);
or U10984 (N_10984,N_9597,N_9227);
and U10985 (N_10985,N_9061,N_9082);
or U10986 (N_10986,N_9889,N_9734);
xnor U10987 (N_10987,N_9775,N_9601);
nand U10988 (N_10988,N_9207,N_9512);
or U10989 (N_10989,N_9373,N_9147);
and U10990 (N_10990,N_9842,N_9110);
xnor U10991 (N_10991,N_9034,N_9671);
or U10992 (N_10992,N_9104,N_9128);
or U10993 (N_10993,N_9478,N_9048);
or U10994 (N_10994,N_9346,N_9631);
nand U10995 (N_10995,N_9899,N_9246);
or U10996 (N_10996,N_9345,N_9971);
and U10997 (N_10997,N_9085,N_9802);
or U10998 (N_10998,N_9344,N_9471);
or U10999 (N_10999,N_9442,N_9346);
nand U11000 (N_11000,N_10311,N_10189);
and U11001 (N_11001,N_10441,N_10392);
and U11002 (N_11002,N_10049,N_10201);
and U11003 (N_11003,N_10591,N_10741);
and U11004 (N_11004,N_10032,N_10157);
nand U11005 (N_11005,N_10621,N_10462);
nand U11006 (N_11006,N_10676,N_10380);
nor U11007 (N_11007,N_10274,N_10921);
or U11008 (N_11008,N_10858,N_10545);
and U11009 (N_11009,N_10335,N_10994);
nand U11010 (N_11010,N_10439,N_10064);
or U11011 (N_11011,N_10907,N_10326);
nand U11012 (N_11012,N_10233,N_10885);
and U11013 (N_11013,N_10565,N_10323);
and U11014 (N_11014,N_10758,N_10127);
nand U11015 (N_11015,N_10953,N_10530);
nand U11016 (N_11016,N_10753,N_10417);
nand U11017 (N_11017,N_10416,N_10261);
and U11018 (N_11018,N_10175,N_10241);
nor U11019 (N_11019,N_10273,N_10935);
nor U11020 (N_11020,N_10160,N_10276);
and U11021 (N_11021,N_10998,N_10493);
or U11022 (N_11022,N_10247,N_10902);
nor U11023 (N_11023,N_10908,N_10029);
nor U11024 (N_11024,N_10541,N_10559);
and U11025 (N_11025,N_10289,N_10697);
xor U11026 (N_11026,N_10632,N_10734);
nor U11027 (N_11027,N_10942,N_10711);
and U11028 (N_11028,N_10874,N_10020);
and U11029 (N_11029,N_10117,N_10245);
or U11030 (N_11030,N_10950,N_10044);
or U11031 (N_11031,N_10546,N_10456);
or U11032 (N_11032,N_10444,N_10321);
nor U11033 (N_11033,N_10582,N_10988);
and U11034 (N_11034,N_10387,N_10472);
and U11035 (N_11035,N_10230,N_10534);
or U11036 (N_11036,N_10768,N_10001);
xnor U11037 (N_11037,N_10759,N_10033);
nor U11038 (N_11038,N_10128,N_10926);
or U11039 (N_11039,N_10188,N_10978);
xor U11040 (N_11040,N_10549,N_10058);
xnor U11041 (N_11041,N_10592,N_10821);
nor U11042 (N_11042,N_10060,N_10014);
and U11043 (N_11043,N_10543,N_10126);
nor U11044 (N_11044,N_10367,N_10186);
and U11045 (N_11045,N_10460,N_10750);
and U11046 (N_11046,N_10699,N_10832);
nand U11047 (N_11047,N_10536,N_10771);
xnor U11048 (N_11048,N_10966,N_10067);
xor U11049 (N_11049,N_10529,N_10584);
nand U11050 (N_11050,N_10791,N_10349);
xor U11051 (N_11051,N_10022,N_10041);
nand U11052 (N_11052,N_10042,N_10708);
xor U11053 (N_11053,N_10286,N_10211);
and U11054 (N_11054,N_10776,N_10903);
nor U11055 (N_11055,N_10923,N_10225);
and U11056 (N_11056,N_10388,N_10912);
nand U11057 (N_11057,N_10946,N_10431);
and U11058 (N_11058,N_10655,N_10981);
nor U11059 (N_11059,N_10607,N_10598);
nor U11060 (N_11060,N_10159,N_10544);
or U11061 (N_11061,N_10085,N_10364);
nand U11062 (N_11062,N_10046,N_10149);
or U11063 (N_11063,N_10875,N_10958);
or U11064 (N_11064,N_10114,N_10499);
xnor U11065 (N_11065,N_10019,N_10644);
nor U11066 (N_11066,N_10865,N_10666);
nor U11067 (N_11067,N_10897,N_10556);
nand U11068 (N_11068,N_10538,N_10939);
and U11069 (N_11069,N_10673,N_10773);
xor U11070 (N_11070,N_10742,N_10688);
xnor U11071 (N_11071,N_10103,N_10518);
or U11072 (N_11072,N_10015,N_10879);
xnor U11073 (N_11073,N_10191,N_10051);
nor U11074 (N_11074,N_10516,N_10365);
nor U11075 (N_11075,N_10256,N_10514);
and U11076 (N_11076,N_10890,N_10037);
and U11077 (N_11077,N_10389,N_10914);
nand U11078 (N_11078,N_10137,N_10925);
nor U11079 (N_11079,N_10146,N_10251);
or U11080 (N_11080,N_10864,N_10457);
or U11081 (N_11081,N_10463,N_10745);
and U11082 (N_11082,N_10718,N_10652);
or U11083 (N_11083,N_10706,N_10415);
nand U11084 (N_11084,N_10096,N_10839);
and U11085 (N_11085,N_10719,N_10316);
xor U11086 (N_11086,N_10943,N_10291);
nor U11087 (N_11087,N_10927,N_10532);
nand U11088 (N_11088,N_10635,N_10449);
nand U11089 (N_11089,N_10731,N_10496);
nor U11090 (N_11090,N_10094,N_10048);
nor U11091 (N_11091,N_10590,N_10356);
or U11092 (N_11092,N_10110,N_10275);
or U11093 (N_11093,N_10278,N_10608);
or U11094 (N_11094,N_10782,N_10414);
or U11095 (N_11095,N_10521,N_10002);
nor U11096 (N_11096,N_10008,N_10694);
nor U11097 (N_11097,N_10976,N_10100);
nand U11098 (N_11098,N_10420,N_10007);
nor U11099 (N_11099,N_10374,N_10980);
and U11100 (N_11100,N_10234,N_10983);
or U11101 (N_11101,N_10979,N_10640);
or U11102 (N_11102,N_10789,N_10259);
xnor U11103 (N_11103,N_10267,N_10740);
nor U11104 (N_11104,N_10111,N_10937);
nor U11105 (N_11105,N_10491,N_10558);
or U11106 (N_11106,N_10329,N_10270);
nand U11107 (N_11107,N_10167,N_10062);
xor U11108 (N_11108,N_10605,N_10038);
nand U11109 (N_11109,N_10299,N_10547);
and U11110 (N_11110,N_10682,N_10393);
nor U11111 (N_11111,N_10124,N_10492);
nand U11112 (N_11112,N_10630,N_10345);
nand U11113 (N_11113,N_10887,N_10170);
xnor U11114 (N_11114,N_10105,N_10113);
xnor U11115 (N_11115,N_10669,N_10373);
or U11116 (N_11116,N_10469,N_10985);
xnor U11117 (N_11117,N_10339,N_10969);
and U11118 (N_11118,N_10869,N_10495);
nand U11119 (N_11119,N_10235,N_10964);
xnor U11120 (N_11120,N_10639,N_10991);
xor U11121 (N_11121,N_10550,N_10264);
xor U11122 (N_11122,N_10130,N_10451);
and U11123 (N_11123,N_10917,N_10760);
nand U11124 (N_11124,N_10799,N_10977);
or U11125 (N_11125,N_10646,N_10295);
or U11126 (N_11126,N_10053,N_10066);
nor U11127 (N_11127,N_10602,N_10184);
or U11128 (N_11128,N_10569,N_10604);
xnor U11129 (N_11129,N_10447,N_10774);
and U11130 (N_11130,N_10829,N_10243);
nand U11131 (N_11131,N_10351,N_10767);
nor U11132 (N_11132,N_10513,N_10886);
nand U11133 (N_11133,N_10575,N_10056);
xor U11134 (N_11134,N_10017,N_10647);
and U11135 (N_11135,N_10272,N_10045);
or U11136 (N_11136,N_10878,N_10656);
or U11137 (N_11137,N_10871,N_10346);
nand U11138 (N_11138,N_10072,N_10433);
or U11139 (N_11139,N_10471,N_10302);
nand U11140 (N_11140,N_10928,N_10982);
nand U11141 (N_11141,N_10715,N_10770);
nor U11142 (N_11142,N_10486,N_10593);
and U11143 (N_11143,N_10571,N_10348);
nand U11144 (N_11144,N_10848,N_10271);
or U11145 (N_11145,N_10827,N_10781);
xnor U11146 (N_11146,N_10717,N_10999);
nand U11147 (N_11147,N_10476,N_10281);
and U11148 (N_11148,N_10319,N_10122);
nor U11149 (N_11149,N_10421,N_10379);
xnor U11150 (N_11150,N_10728,N_10624);
nand U11151 (N_11151,N_10083,N_10301);
nand U11152 (N_11152,N_10689,N_10654);
and U11153 (N_11153,N_10063,N_10138);
nor U11154 (N_11154,N_10509,N_10617);
xor U11155 (N_11155,N_10405,N_10819);
or U11156 (N_11156,N_10406,N_10112);
or U11157 (N_11157,N_10010,N_10880);
and U11158 (N_11158,N_10814,N_10080);
nand U11159 (N_11159,N_10594,N_10280);
nand U11160 (N_11160,N_10342,N_10086);
or U11161 (N_11161,N_10574,N_10338);
or U11162 (N_11162,N_10250,N_10504);
nand U11163 (N_11163,N_10714,N_10034);
or U11164 (N_11164,N_10068,N_10418);
or U11165 (N_11165,N_10199,N_10766);
and U11166 (N_11166,N_10055,N_10363);
xnor U11167 (N_11167,N_10906,N_10336);
and U11168 (N_11168,N_10372,N_10817);
or U11169 (N_11169,N_10485,N_10487);
nor U11170 (N_11170,N_10482,N_10949);
and U11171 (N_11171,N_10992,N_10801);
and U11172 (N_11172,N_10361,N_10526);
or U11173 (N_11173,N_10101,N_10479);
or U11174 (N_11174,N_10400,N_10973);
and U11175 (N_11175,N_10798,N_10169);
nor U11176 (N_11176,N_10077,N_10653);
xor U11177 (N_11177,N_10628,N_10325);
xor U11178 (N_11178,N_10721,N_10833);
or U11179 (N_11179,N_10026,N_10187);
nor U11180 (N_11180,N_10207,N_10733);
nand U11181 (N_11181,N_10023,N_10828);
nand U11182 (N_11182,N_10109,N_10967);
nand U11183 (N_11183,N_10643,N_10129);
nor U11184 (N_11184,N_10665,N_10783);
and U11185 (N_11185,N_10986,N_10573);
nor U11186 (N_11186,N_10877,N_10772);
and U11187 (N_11187,N_10580,N_10788);
and U11188 (N_11188,N_10279,N_10432);
nor U11189 (N_11189,N_10488,N_10362);
and U11190 (N_11190,N_10039,N_10586);
and U11191 (N_11191,N_10309,N_10030);
and U11192 (N_11192,N_10830,N_10151);
nand U11193 (N_11193,N_10841,N_10754);
xnor U11194 (N_11194,N_10443,N_10929);
xnor U11195 (N_11195,N_10383,N_10528);
nand U11196 (N_11196,N_10036,N_10687);
or U11197 (N_11197,N_10857,N_10566);
xnor U11198 (N_11198,N_10107,N_10568);
nor U11199 (N_11199,N_10428,N_10990);
nor U11200 (N_11200,N_10664,N_10555);
nand U11201 (N_11201,N_10614,N_10438);
and U11202 (N_11202,N_10872,N_10458);
nand U11203 (N_11203,N_10401,N_10497);
nor U11204 (N_11204,N_10494,N_10436);
and U11205 (N_11205,N_10695,N_10779);
and U11206 (N_11206,N_10920,N_10623);
or U11207 (N_11207,N_10206,N_10856);
xnor U11208 (N_11208,N_10308,N_10963);
xor U11209 (N_11209,N_10563,N_10394);
nor U11210 (N_11210,N_10061,N_10752);
nor U11211 (N_11211,N_10993,N_10587);
or U11212 (N_11212,N_10320,N_10501);
or U11213 (N_11213,N_10370,N_10961);
or U11214 (N_11214,N_10738,N_10317);
xnor U11215 (N_11215,N_10355,N_10181);
nor U11216 (N_11216,N_10422,N_10629);
xor U11217 (N_11217,N_10411,N_10163);
nor U11218 (N_11218,N_10508,N_10088);
xnor U11219 (N_11219,N_10054,N_10746);
or U11220 (N_11220,N_10262,N_10284);
and U11221 (N_11221,N_10304,N_10765);
or U11222 (N_11222,N_10919,N_10884);
nand U11223 (N_11223,N_10288,N_10334);
nand U11224 (N_11224,N_10135,N_10076);
nand U11225 (N_11225,N_10900,N_10174);
nor U11226 (N_11226,N_10164,N_10627);
nand U11227 (N_11227,N_10681,N_10385);
nand U11228 (N_11228,N_10337,N_10940);
xnor U11229 (N_11229,N_10260,N_10596);
nand U11230 (N_11230,N_10358,N_10778);
xnor U11231 (N_11231,N_10984,N_10232);
and U11232 (N_11232,N_10330,N_10567);
xnor U11233 (N_11233,N_10747,N_10579);
nand U11234 (N_11234,N_10470,N_10947);
xnor U11235 (N_11235,N_10474,N_10924);
or U11236 (N_11236,N_10217,N_10661);
and U11237 (N_11237,N_10231,N_10934);
nand U11238 (N_11238,N_10769,N_10141);
or U11239 (N_11239,N_10298,N_10861);
nand U11240 (N_11240,N_10527,N_10836);
nand U11241 (N_11241,N_10484,N_10564);
nand U11242 (N_11242,N_10266,N_10743);
nand U11243 (N_11243,N_10720,N_10576);
nand U11244 (N_11244,N_10822,N_10737);
or U11245 (N_11245,N_10246,N_10294);
nand U11246 (N_11246,N_10540,N_10227);
nand U11247 (N_11247,N_10248,N_10390);
nand U11248 (N_11248,N_10180,N_10177);
nor U11249 (N_11249,N_10209,N_10148);
and U11250 (N_11250,N_10686,N_10183);
nand U11251 (N_11251,N_10889,N_10079);
nand U11252 (N_11252,N_10219,N_10483);
nor U11253 (N_11253,N_10490,N_10677);
or U11254 (N_11254,N_10888,N_10143);
and U11255 (N_11255,N_10818,N_10704);
and U11256 (N_11256,N_10905,N_10794);
nor U11257 (N_11257,N_10703,N_10396);
and U11258 (N_11258,N_10852,N_10601);
nor U11259 (N_11259,N_10867,N_10178);
nor U11260 (N_11260,N_10360,N_10730);
or U11261 (N_11261,N_10615,N_10222);
nand U11262 (N_11262,N_10645,N_10659);
nor U11263 (N_11263,N_10723,N_10854);
and U11264 (N_11264,N_10724,N_10748);
xor U11265 (N_11265,N_10005,N_10764);
nand U11266 (N_11266,N_10312,N_10739);
and U11267 (N_11267,N_10347,N_10324);
and U11268 (N_11268,N_10554,N_10932);
nor U11269 (N_11269,N_10793,N_10027);
nor U11270 (N_11270,N_10812,N_10354);
and U11271 (N_11271,N_10249,N_10402);
nor U11272 (N_11272,N_10826,N_10369);
and U11273 (N_11273,N_10156,N_10104);
nor U11274 (N_11274,N_10296,N_10603);
nor U11275 (N_11275,N_10589,N_10391);
nand U11276 (N_11276,N_10909,N_10059);
and U11277 (N_11277,N_10016,N_10705);
xnor U11278 (N_11278,N_10140,N_10203);
xnor U11279 (N_11279,N_10423,N_10384);
xnor U11280 (N_11280,N_10445,N_10680);
xnor U11281 (N_11281,N_10252,N_10712);
nor U11282 (N_11282,N_10331,N_10253);
nor U11283 (N_11283,N_10859,N_10892);
nand U11284 (N_11284,N_10366,N_10710);
xnor U11285 (N_11285,N_10408,N_10155);
and U11286 (N_11286,N_10805,N_10226);
or U11287 (N_11287,N_10552,N_10519);
nor U11288 (N_11288,N_10663,N_10620);
xor U11289 (N_11289,N_10820,N_10202);
xor U11290 (N_11290,N_10609,N_10860);
xnor U11291 (N_11291,N_10168,N_10018);
nor U11292 (N_11292,N_10883,N_10955);
nor U11293 (N_11293,N_10310,N_10065);
or U11294 (N_11294,N_10314,N_10473);
xor U11295 (N_11295,N_10700,N_10690);
or U11296 (N_11296,N_10638,N_10244);
nor U11297 (N_11297,N_10825,N_10404);
and U11298 (N_11298,N_10397,N_10965);
nand U11299 (N_11299,N_10084,N_10726);
or U11300 (N_11300,N_10702,N_10631);
xnor U11301 (N_11301,N_10553,N_10729);
nand U11302 (N_11302,N_10727,N_10378);
xnor U11303 (N_11303,N_10954,N_10678);
nor U11304 (N_11304,N_10693,N_10333);
or U11305 (N_11305,N_10399,N_10268);
nand U11306 (N_11306,N_10523,N_10971);
nor U11307 (N_11307,N_10386,N_10255);
nor U11308 (N_11308,N_10960,N_10489);
and U11309 (N_11309,N_10823,N_10834);
nor U11310 (N_11310,N_10208,N_10802);
or U11311 (N_11311,N_10240,N_10093);
and U11312 (N_11312,N_10307,N_10698);
nand U11313 (N_11313,N_10173,N_10938);
and U11314 (N_11314,N_10870,N_10855);
nor U11315 (N_11315,N_10835,N_10707);
or U11316 (N_11316,N_10735,N_10882);
nand U11317 (N_11317,N_10011,N_10548);
nor U11318 (N_11318,N_10918,N_10775);
and U11319 (N_11319,N_10134,N_10377);
and U11320 (N_11320,N_10916,N_10679);
or U11321 (N_11321,N_10749,N_10375);
nor U11322 (N_11322,N_10931,N_10896);
nand U11323 (N_11323,N_10132,N_10756);
and U11324 (N_11324,N_10468,N_10071);
or U11325 (N_11325,N_10413,N_10811);
nand U11326 (N_11326,N_10442,N_10962);
or U11327 (N_11327,N_10637,N_10006);
nand U11328 (N_11328,N_10292,N_10099);
xnor U11329 (N_11329,N_10282,N_10236);
xnor U11330 (N_11330,N_10322,N_10344);
nor U11331 (N_11331,N_10481,N_10263);
nand U11332 (N_11332,N_10784,N_10172);
nor U11333 (N_11333,N_10816,N_10102);
nor U11334 (N_11334,N_10618,N_10082);
and U11335 (N_11335,N_10987,N_10806);
nor U11336 (N_11336,N_10277,N_10095);
nand U11337 (N_11337,N_10303,N_10641);
xor U11338 (N_11338,N_10936,N_10585);
nor U11339 (N_11339,N_10464,N_10824);
or U11340 (N_11340,N_10459,N_10813);
or U11341 (N_11341,N_10893,N_10097);
and U11342 (N_11342,N_10193,N_10692);
nand U11343 (N_11343,N_10634,N_10520);
and U11344 (N_11344,N_10945,N_10315);
xnor U11345 (N_11345,N_10911,N_10013);
nand U11346 (N_11346,N_10531,N_10974);
nor U11347 (N_11347,N_10803,N_10616);
xnor U11348 (N_11348,N_10507,N_10198);
or U11349 (N_11349,N_10121,N_10777);
nor U11350 (N_11350,N_10670,N_10948);
nand U11351 (N_11351,N_10158,N_10257);
and U11352 (N_11352,N_10522,N_10133);
nand U11353 (N_11353,N_10283,N_10658);
nand U11354 (N_11354,N_10505,N_10838);
and U11355 (N_11355,N_10787,N_10040);
nand U11356 (N_11356,N_10997,N_10578);
and U11357 (N_11357,N_10762,N_10142);
or U11358 (N_11358,N_10732,N_10480);
and U11359 (N_11359,N_10668,N_10419);
and U11360 (N_11360,N_10000,N_10780);
nand U11361 (N_11361,N_10503,N_10959);
or U11362 (N_11362,N_10525,N_10403);
nand U11363 (N_11363,N_10152,N_10810);
nor U11364 (N_11364,N_10150,N_10581);
xnor U11365 (N_11365,N_10891,N_10506);
or U11366 (N_11366,N_10357,N_10238);
xnor U11367 (N_11367,N_10613,N_10537);
xor U11368 (N_11368,N_10290,N_10098);
nor U11369 (N_11369,N_10131,N_10570);
xor U11370 (N_11370,N_10951,N_10287);
nand U11371 (N_11371,N_10381,N_10179);
nor U11372 (N_11372,N_10145,N_10642);
and U11373 (N_11373,N_10269,N_10873);
nor U11374 (N_11374,N_10561,N_10736);
nand U11375 (N_11375,N_10437,N_10434);
xor U11376 (N_11376,N_10119,N_10265);
xor U11377 (N_11377,N_10081,N_10674);
or U11378 (N_11378,N_10043,N_10972);
nand U11379 (N_11379,N_10847,N_10341);
and U11380 (N_11380,N_10595,N_10807);
xor U11381 (N_11381,N_10205,N_10751);
or U11382 (N_11382,N_10619,N_10868);
or U11383 (N_11383,N_10722,N_10995);
nor U11384 (N_11384,N_10125,N_10024);
nand U11385 (N_11385,N_10667,N_10218);
nor U11386 (N_11386,N_10849,N_10427);
xor U11387 (N_11387,N_10808,N_10210);
xor U11388 (N_11388,N_10190,N_10539);
and U11389 (N_11389,N_10498,N_10144);
xnor U11390 (N_11390,N_10691,N_10057);
and U11391 (N_11391,N_10551,N_10475);
nand U11392 (N_11392,N_10410,N_10376);
and U11393 (N_11393,N_10657,N_10612);
and U11394 (N_11394,N_10597,N_10904);
and U11395 (N_11395,N_10610,N_10254);
nand U11396 (N_11396,N_10293,N_10957);
xnor U11397 (N_11397,N_10467,N_10662);
and U11398 (N_11398,N_10328,N_10047);
nand U11399 (N_11399,N_10910,N_10116);
nand U11400 (N_11400,N_10672,N_10761);
nand U11401 (N_11401,N_10685,N_10862);
or U11402 (N_11402,N_10606,N_10340);
nand U11403 (N_11403,N_10863,N_10542);
xnor U11404 (N_11404,N_10285,N_10196);
or U11405 (N_11405,N_10162,N_10424);
or U11406 (N_11406,N_10757,N_10166);
nor U11407 (N_11407,N_10200,N_10407);
or U11408 (N_11408,N_10785,N_10881);
xor U11409 (N_11409,N_10792,N_10840);
or U11410 (N_11410,N_10306,N_10352);
nand U11411 (N_11411,N_10989,N_10915);
or U11412 (N_11412,N_10028,N_10696);
xnor U11413 (N_11413,N_10996,N_10395);
nor U11414 (N_11414,N_10300,N_10465);
nand U11415 (N_11415,N_10089,N_10895);
nor U11416 (N_11416,N_10115,N_10412);
nand U11417 (N_11417,N_10052,N_10454);
nor U11418 (N_11418,N_10012,N_10583);
xor U11419 (N_11419,N_10165,N_10429);
and U11420 (N_11420,N_10683,N_10195);
nor U11421 (N_11421,N_10185,N_10804);
xnor U11422 (N_11422,N_10837,N_10633);
and U11423 (N_11423,N_10648,N_10239);
xor U11424 (N_11424,N_10409,N_10216);
nor U11425 (N_11425,N_10371,N_10327);
and U11426 (N_11426,N_10078,N_10073);
and U11427 (N_11427,N_10572,N_10069);
xor U11428 (N_11428,N_10229,N_10204);
xor U11429 (N_11429,N_10511,N_10297);
or U11430 (N_11430,N_10332,N_10074);
nand U11431 (N_11431,N_10557,N_10343);
nor U11432 (N_11432,N_10588,N_10035);
xnor U11433 (N_11433,N_10025,N_10197);
nor U11434 (N_11434,N_10398,N_10368);
nand U11435 (N_11435,N_10651,N_10933);
nand U11436 (N_11436,N_10123,N_10853);
and U11437 (N_11437,N_10182,N_10899);
nor U11438 (N_11438,N_10725,N_10220);
or U11439 (N_11439,N_10430,N_10258);
or U11440 (N_11440,N_10815,N_10795);
nand U11441 (N_11441,N_10831,N_10176);
and U11442 (N_11442,N_10154,N_10913);
nand U11443 (N_11443,N_10562,N_10215);
and U11444 (N_11444,N_10139,N_10500);
nand U11445 (N_11445,N_10626,N_10213);
or U11446 (N_11446,N_10599,N_10050);
nand U11447 (N_11447,N_10510,N_10461);
and U11448 (N_11448,N_10382,N_10224);
nand U11449 (N_11449,N_10452,N_10106);
and U11450 (N_11450,N_10212,N_10577);
and U11451 (N_11451,N_10090,N_10003);
or U11452 (N_11452,N_10517,N_10786);
or U11453 (N_11453,N_10763,N_10161);
or U11454 (N_11454,N_10649,N_10956);
xor U11455 (N_11455,N_10466,N_10313);
and U11456 (N_11456,N_10350,N_10560);
nor U11457 (N_11457,N_10171,N_10031);
nor U11458 (N_11458,N_10426,N_10087);
or U11459 (N_11459,N_10075,N_10660);
nand U11460 (N_11460,N_10533,N_10894);
or U11461 (N_11461,N_10446,N_10070);
or U11462 (N_11462,N_10502,N_10851);
and U11463 (N_11463,N_10194,N_10975);
nor U11464 (N_11464,N_10228,N_10713);
nor U11465 (N_11465,N_10636,N_10448);
nand U11466 (N_11466,N_10535,N_10515);
nor U11467 (N_11467,N_10092,N_10952);
or U11468 (N_11468,N_10930,N_10425);
nand U11469 (N_11469,N_10800,N_10625);
or U11470 (N_11470,N_10009,N_10091);
and U11471 (N_11471,N_10922,N_10845);
nand U11472 (N_11472,N_10136,N_10843);
nand U11473 (N_11473,N_10004,N_10866);
and U11474 (N_11474,N_10223,N_10842);
nor U11475 (N_11475,N_10844,N_10192);
xor U11476 (N_11476,N_10675,N_10237);
nor U11477 (N_11477,N_10901,N_10755);
and U11478 (N_11478,N_10944,N_10650);
and U11479 (N_11479,N_10242,N_10898);
nand U11480 (N_11480,N_10744,N_10611);
xor U11481 (N_11481,N_10477,N_10435);
or U11482 (N_11482,N_10478,N_10359);
nor U11483 (N_11483,N_10797,N_10147);
nor U11484 (N_11484,N_10790,N_10968);
or U11485 (N_11485,N_10524,N_10021);
nor U11486 (N_11486,N_10455,N_10701);
nor U11487 (N_11487,N_10118,N_10716);
xor U11488 (N_11488,N_10846,N_10153);
xor U11489 (N_11489,N_10876,N_10941);
xor U11490 (N_11490,N_10709,N_10450);
nand U11491 (N_11491,N_10809,N_10684);
nor U11492 (N_11492,N_10440,N_10453);
and U11493 (N_11493,N_10671,N_10850);
nand U11494 (N_11494,N_10221,N_10970);
nand U11495 (N_11495,N_10120,N_10214);
and U11496 (N_11496,N_10512,N_10622);
or U11497 (N_11497,N_10796,N_10600);
or U11498 (N_11498,N_10318,N_10108);
and U11499 (N_11499,N_10353,N_10305);
or U11500 (N_11500,N_10212,N_10640);
xnor U11501 (N_11501,N_10373,N_10286);
xor U11502 (N_11502,N_10273,N_10472);
nor U11503 (N_11503,N_10554,N_10824);
nor U11504 (N_11504,N_10264,N_10770);
and U11505 (N_11505,N_10088,N_10044);
nand U11506 (N_11506,N_10274,N_10781);
or U11507 (N_11507,N_10528,N_10051);
nand U11508 (N_11508,N_10127,N_10926);
xor U11509 (N_11509,N_10921,N_10504);
nor U11510 (N_11510,N_10625,N_10401);
or U11511 (N_11511,N_10545,N_10426);
nor U11512 (N_11512,N_10857,N_10879);
nor U11513 (N_11513,N_10528,N_10482);
or U11514 (N_11514,N_10688,N_10770);
nand U11515 (N_11515,N_10587,N_10622);
nor U11516 (N_11516,N_10312,N_10298);
xnor U11517 (N_11517,N_10422,N_10853);
nor U11518 (N_11518,N_10779,N_10102);
or U11519 (N_11519,N_10463,N_10196);
nor U11520 (N_11520,N_10130,N_10332);
or U11521 (N_11521,N_10351,N_10735);
and U11522 (N_11522,N_10426,N_10526);
or U11523 (N_11523,N_10054,N_10922);
or U11524 (N_11524,N_10534,N_10870);
xnor U11525 (N_11525,N_10580,N_10526);
and U11526 (N_11526,N_10027,N_10260);
nand U11527 (N_11527,N_10693,N_10387);
xnor U11528 (N_11528,N_10728,N_10339);
nand U11529 (N_11529,N_10974,N_10406);
or U11530 (N_11530,N_10915,N_10690);
nand U11531 (N_11531,N_10988,N_10746);
or U11532 (N_11532,N_10846,N_10309);
or U11533 (N_11533,N_10094,N_10288);
nor U11534 (N_11534,N_10392,N_10262);
nor U11535 (N_11535,N_10003,N_10556);
and U11536 (N_11536,N_10579,N_10294);
or U11537 (N_11537,N_10498,N_10935);
nor U11538 (N_11538,N_10078,N_10117);
nor U11539 (N_11539,N_10525,N_10607);
nand U11540 (N_11540,N_10149,N_10782);
xnor U11541 (N_11541,N_10550,N_10987);
and U11542 (N_11542,N_10688,N_10019);
nor U11543 (N_11543,N_10920,N_10707);
xnor U11544 (N_11544,N_10298,N_10745);
and U11545 (N_11545,N_10646,N_10206);
nand U11546 (N_11546,N_10094,N_10753);
nor U11547 (N_11547,N_10138,N_10002);
xor U11548 (N_11548,N_10245,N_10553);
or U11549 (N_11549,N_10819,N_10631);
nor U11550 (N_11550,N_10329,N_10526);
xor U11551 (N_11551,N_10759,N_10317);
or U11552 (N_11552,N_10617,N_10951);
xor U11553 (N_11553,N_10204,N_10351);
and U11554 (N_11554,N_10058,N_10433);
and U11555 (N_11555,N_10616,N_10723);
and U11556 (N_11556,N_10024,N_10373);
nor U11557 (N_11557,N_10311,N_10354);
nand U11558 (N_11558,N_10518,N_10892);
or U11559 (N_11559,N_10727,N_10177);
and U11560 (N_11560,N_10343,N_10672);
nand U11561 (N_11561,N_10177,N_10349);
or U11562 (N_11562,N_10914,N_10710);
nor U11563 (N_11563,N_10362,N_10616);
nor U11564 (N_11564,N_10083,N_10672);
or U11565 (N_11565,N_10032,N_10319);
or U11566 (N_11566,N_10783,N_10522);
or U11567 (N_11567,N_10387,N_10398);
nor U11568 (N_11568,N_10322,N_10501);
xnor U11569 (N_11569,N_10484,N_10551);
nand U11570 (N_11570,N_10558,N_10949);
nand U11571 (N_11571,N_10514,N_10100);
and U11572 (N_11572,N_10784,N_10527);
xnor U11573 (N_11573,N_10150,N_10139);
nand U11574 (N_11574,N_10898,N_10459);
nand U11575 (N_11575,N_10619,N_10101);
or U11576 (N_11576,N_10785,N_10058);
xnor U11577 (N_11577,N_10783,N_10876);
or U11578 (N_11578,N_10234,N_10871);
and U11579 (N_11579,N_10789,N_10952);
xor U11580 (N_11580,N_10660,N_10192);
xor U11581 (N_11581,N_10978,N_10118);
and U11582 (N_11582,N_10006,N_10808);
nand U11583 (N_11583,N_10936,N_10348);
nor U11584 (N_11584,N_10735,N_10430);
and U11585 (N_11585,N_10651,N_10047);
and U11586 (N_11586,N_10473,N_10317);
or U11587 (N_11587,N_10441,N_10806);
nand U11588 (N_11588,N_10765,N_10725);
nand U11589 (N_11589,N_10743,N_10960);
or U11590 (N_11590,N_10551,N_10197);
and U11591 (N_11591,N_10462,N_10389);
xor U11592 (N_11592,N_10052,N_10838);
nor U11593 (N_11593,N_10886,N_10287);
xor U11594 (N_11594,N_10536,N_10650);
xnor U11595 (N_11595,N_10306,N_10454);
and U11596 (N_11596,N_10076,N_10334);
xnor U11597 (N_11597,N_10566,N_10498);
and U11598 (N_11598,N_10892,N_10103);
nor U11599 (N_11599,N_10654,N_10814);
xnor U11600 (N_11600,N_10845,N_10302);
nand U11601 (N_11601,N_10648,N_10204);
nand U11602 (N_11602,N_10134,N_10707);
xnor U11603 (N_11603,N_10555,N_10798);
nor U11604 (N_11604,N_10985,N_10202);
nor U11605 (N_11605,N_10744,N_10524);
or U11606 (N_11606,N_10341,N_10012);
nand U11607 (N_11607,N_10555,N_10684);
or U11608 (N_11608,N_10476,N_10884);
nand U11609 (N_11609,N_10067,N_10667);
or U11610 (N_11610,N_10033,N_10501);
or U11611 (N_11611,N_10160,N_10665);
nor U11612 (N_11612,N_10518,N_10743);
nand U11613 (N_11613,N_10987,N_10696);
and U11614 (N_11614,N_10365,N_10972);
and U11615 (N_11615,N_10706,N_10608);
nor U11616 (N_11616,N_10337,N_10853);
xor U11617 (N_11617,N_10073,N_10860);
nand U11618 (N_11618,N_10326,N_10837);
nand U11619 (N_11619,N_10718,N_10663);
nor U11620 (N_11620,N_10931,N_10510);
or U11621 (N_11621,N_10694,N_10606);
nand U11622 (N_11622,N_10915,N_10391);
and U11623 (N_11623,N_10744,N_10319);
xor U11624 (N_11624,N_10809,N_10144);
nor U11625 (N_11625,N_10669,N_10000);
or U11626 (N_11626,N_10193,N_10020);
xnor U11627 (N_11627,N_10920,N_10270);
and U11628 (N_11628,N_10631,N_10244);
nor U11629 (N_11629,N_10394,N_10779);
and U11630 (N_11630,N_10785,N_10470);
xnor U11631 (N_11631,N_10817,N_10332);
nor U11632 (N_11632,N_10382,N_10377);
and U11633 (N_11633,N_10260,N_10788);
xor U11634 (N_11634,N_10384,N_10560);
nand U11635 (N_11635,N_10162,N_10734);
nor U11636 (N_11636,N_10957,N_10386);
nor U11637 (N_11637,N_10124,N_10608);
and U11638 (N_11638,N_10157,N_10432);
and U11639 (N_11639,N_10144,N_10293);
xor U11640 (N_11640,N_10395,N_10273);
and U11641 (N_11641,N_10532,N_10878);
nor U11642 (N_11642,N_10027,N_10288);
nor U11643 (N_11643,N_10021,N_10729);
nand U11644 (N_11644,N_10498,N_10923);
or U11645 (N_11645,N_10693,N_10278);
xor U11646 (N_11646,N_10488,N_10639);
nor U11647 (N_11647,N_10155,N_10311);
and U11648 (N_11648,N_10599,N_10627);
or U11649 (N_11649,N_10836,N_10602);
or U11650 (N_11650,N_10759,N_10639);
or U11651 (N_11651,N_10098,N_10610);
or U11652 (N_11652,N_10669,N_10661);
or U11653 (N_11653,N_10882,N_10364);
nand U11654 (N_11654,N_10688,N_10769);
nand U11655 (N_11655,N_10213,N_10008);
and U11656 (N_11656,N_10079,N_10438);
and U11657 (N_11657,N_10266,N_10899);
or U11658 (N_11658,N_10493,N_10910);
nand U11659 (N_11659,N_10380,N_10982);
nor U11660 (N_11660,N_10748,N_10813);
or U11661 (N_11661,N_10500,N_10585);
nand U11662 (N_11662,N_10578,N_10228);
nand U11663 (N_11663,N_10173,N_10006);
or U11664 (N_11664,N_10172,N_10290);
xor U11665 (N_11665,N_10397,N_10299);
xnor U11666 (N_11666,N_10758,N_10598);
nand U11667 (N_11667,N_10467,N_10698);
xor U11668 (N_11668,N_10826,N_10442);
xnor U11669 (N_11669,N_10862,N_10098);
and U11670 (N_11670,N_10461,N_10183);
and U11671 (N_11671,N_10207,N_10483);
or U11672 (N_11672,N_10453,N_10457);
nor U11673 (N_11673,N_10383,N_10829);
nor U11674 (N_11674,N_10337,N_10282);
nand U11675 (N_11675,N_10025,N_10341);
xnor U11676 (N_11676,N_10832,N_10337);
xnor U11677 (N_11677,N_10822,N_10550);
xor U11678 (N_11678,N_10546,N_10234);
xor U11679 (N_11679,N_10850,N_10463);
nand U11680 (N_11680,N_10498,N_10681);
and U11681 (N_11681,N_10546,N_10312);
and U11682 (N_11682,N_10394,N_10597);
and U11683 (N_11683,N_10996,N_10533);
xor U11684 (N_11684,N_10970,N_10973);
and U11685 (N_11685,N_10114,N_10846);
nor U11686 (N_11686,N_10762,N_10377);
nand U11687 (N_11687,N_10113,N_10467);
xor U11688 (N_11688,N_10195,N_10922);
nand U11689 (N_11689,N_10730,N_10461);
nor U11690 (N_11690,N_10950,N_10694);
or U11691 (N_11691,N_10551,N_10058);
and U11692 (N_11692,N_10471,N_10670);
nor U11693 (N_11693,N_10262,N_10237);
nor U11694 (N_11694,N_10029,N_10307);
or U11695 (N_11695,N_10956,N_10911);
and U11696 (N_11696,N_10393,N_10565);
and U11697 (N_11697,N_10165,N_10676);
or U11698 (N_11698,N_10022,N_10062);
or U11699 (N_11699,N_10927,N_10515);
xnor U11700 (N_11700,N_10012,N_10058);
xnor U11701 (N_11701,N_10650,N_10619);
and U11702 (N_11702,N_10368,N_10761);
nand U11703 (N_11703,N_10607,N_10300);
or U11704 (N_11704,N_10612,N_10595);
nand U11705 (N_11705,N_10872,N_10428);
nor U11706 (N_11706,N_10613,N_10085);
nand U11707 (N_11707,N_10816,N_10494);
and U11708 (N_11708,N_10783,N_10924);
xor U11709 (N_11709,N_10065,N_10275);
xnor U11710 (N_11710,N_10797,N_10365);
nor U11711 (N_11711,N_10509,N_10182);
and U11712 (N_11712,N_10971,N_10798);
nor U11713 (N_11713,N_10597,N_10341);
nand U11714 (N_11714,N_10192,N_10172);
or U11715 (N_11715,N_10521,N_10539);
xnor U11716 (N_11716,N_10117,N_10379);
xor U11717 (N_11717,N_10214,N_10552);
or U11718 (N_11718,N_10493,N_10539);
nor U11719 (N_11719,N_10639,N_10240);
and U11720 (N_11720,N_10577,N_10769);
nor U11721 (N_11721,N_10455,N_10423);
xnor U11722 (N_11722,N_10848,N_10257);
and U11723 (N_11723,N_10911,N_10601);
xor U11724 (N_11724,N_10222,N_10267);
and U11725 (N_11725,N_10303,N_10602);
nand U11726 (N_11726,N_10556,N_10751);
nand U11727 (N_11727,N_10340,N_10125);
nand U11728 (N_11728,N_10373,N_10589);
xnor U11729 (N_11729,N_10345,N_10434);
xnor U11730 (N_11730,N_10899,N_10701);
xor U11731 (N_11731,N_10042,N_10938);
xnor U11732 (N_11732,N_10480,N_10709);
or U11733 (N_11733,N_10525,N_10072);
or U11734 (N_11734,N_10067,N_10921);
xor U11735 (N_11735,N_10360,N_10682);
or U11736 (N_11736,N_10246,N_10206);
xor U11737 (N_11737,N_10104,N_10985);
nor U11738 (N_11738,N_10868,N_10547);
nand U11739 (N_11739,N_10241,N_10059);
nand U11740 (N_11740,N_10512,N_10854);
nor U11741 (N_11741,N_10258,N_10644);
nand U11742 (N_11742,N_10425,N_10214);
or U11743 (N_11743,N_10881,N_10435);
xor U11744 (N_11744,N_10612,N_10220);
and U11745 (N_11745,N_10456,N_10899);
nor U11746 (N_11746,N_10923,N_10340);
xnor U11747 (N_11747,N_10688,N_10347);
and U11748 (N_11748,N_10706,N_10861);
and U11749 (N_11749,N_10955,N_10528);
nor U11750 (N_11750,N_10210,N_10828);
nor U11751 (N_11751,N_10815,N_10350);
or U11752 (N_11752,N_10811,N_10996);
nor U11753 (N_11753,N_10325,N_10287);
or U11754 (N_11754,N_10634,N_10600);
or U11755 (N_11755,N_10505,N_10354);
nand U11756 (N_11756,N_10410,N_10880);
and U11757 (N_11757,N_10607,N_10447);
and U11758 (N_11758,N_10199,N_10941);
or U11759 (N_11759,N_10635,N_10000);
nor U11760 (N_11760,N_10576,N_10381);
nand U11761 (N_11761,N_10395,N_10609);
nor U11762 (N_11762,N_10141,N_10613);
nand U11763 (N_11763,N_10922,N_10130);
xnor U11764 (N_11764,N_10736,N_10385);
nor U11765 (N_11765,N_10252,N_10688);
xnor U11766 (N_11766,N_10744,N_10214);
xor U11767 (N_11767,N_10689,N_10521);
nor U11768 (N_11768,N_10332,N_10527);
xor U11769 (N_11769,N_10750,N_10529);
or U11770 (N_11770,N_10827,N_10119);
nand U11771 (N_11771,N_10610,N_10154);
or U11772 (N_11772,N_10391,N_10116);
xor U11773 (N_11773,N_10715,N_10702);
or U11774 (N_11774,N_10940,N_10895);
or U11775 (N_11775,N_10589,N_10257);
or U11776 (N_11776,N_10211,N_10145);
or U11777 (N_11777,N_10613,N_10912);
xnor U11778 (N_11778,N_10725,N_10752);
nand U11779 (N_11779,N_10101,N_10719);
xnor U11780 (N_11780,N_10989,N_10529);
xor U11781 (N_11781,N_10671,N_10020);
xor U11782 (N_11782,N_10495,N_10741);
xor U11783 (N_11783,N_10849,N_10096);
or U11784 (N_11784,N_10287,N_10410);
or U11785 (N_11785,N_10975,N_10338);
nand U11786 (N_11786,N_10739,N_10428);
and U11787 (N_11787,N_10756,N_10510);
or U11788 (N_11788,N_10735,N_10892);
and U11789 (N_11789,N_10062,N_10556);
or U11790 (N_11790,N_10107,N_10328);
xor U11791 (N_11791,N_10097,N_10464);
xor U11792 (N_11792,N_10104,N_10284);
nand U11793 (N_11793,N_10466,N_10343);
and U11794 (N_11794,N_10396,N_10303);
and U11795 (N_11795,N_10755,N_10471);
nand U11796 (N_11796,N_10844,N_10629);
and U11797 (N_11797,N_10464,N_10432);
xor U11798 (N_11798,N_10415,N_10731);
or U11799 (N_11799,N_10694,N_10360);
nor U11800 (N_11800,N_10430,N_10551);
nor U11801 (N_11801,N_10443,N_10291);
or U11802 (N_11802,N_10782,N_10361);
or U11803 (N_11803,N_10864,N_10992);
nor U11804 (N_11804,N_10987,N_10710);
or U11805 (N_11805,N_10172,N_10508);
xnor U11806 (N_11806,N_10079,N_10785);
and U11807 (N_11807,N_10825,N_10994);
nand U11808 (N_11808,N_10943,N_10167);
xor U11809 (N_11809,N_10349,N_10306);
nand U11810 (N_11810,N_10597,N_10999);
nor U11811 (N_11811,N_10951,N_10597);
xor U11812 (N_11812,N_10101,N_10408);
nor U11813 (N_11813,N_10889,N_10657);
nand U11814 (N_11814,N_10524,N_10743);
nor U11815 (N_11815,N_10680,N_10702);
nand U11816 (N_11816,N_10889,N_10040);
xnor U11817 (N_11817,N_10552,N_10154);
or U11818 (N_11818,N_10347,N_10617);
and U11819 (N_11819,N_10414,N_10364);
nand U11820 (N_11820,N_10211,N_10959);
and U11821 (N_11821,N_10444,N_10311);
or U11822 (N_11822,N_10164,N_10094);
xnor U11823 (N_11823,N_10326,N_10590);
nor U11824 (N_11824,N_10412,N_10851);
xnor U11825 (N_11825,N_10193,N_10640);
nand U11826 (N_11826,N_10386,N_10080);
or U11827 (N_11827,N_10936,N_10626);
nor U11828 (N_11828,N_10458,N_10606);
nor U11829 (N_11829,N_10178,N_10037);
or U11830 (N_11830,N_10626,N_10183);
xor U11831 (N_11831,N_10401,N_10195);
nand U11832 (N_11832,N_10577,N_10390);
or U11833 (N_11833,N_10469,N_10731);
nand U11834 (N_11834,N_10313,N_10248);
xnor U11835 (N_11835,N_10102,N_10040);
nand U11836 (N_11836,N_10667,N_10834);
and U11837 (N_11837,N_10296,N_10285);
nand U11838 (N_11838,N_10372,N_10126);
and U11839 (N_11839,N_10398,N_10083);
xor U11840 (N_11840,N_10581,N_10639);
nand U11841 (N_11841,N_10578,N_10490);
nor U11842 (N_11842,N_10970,N_10593);
and U11843 (N_11843,N_10895,N_10965);
nand U11844 (N_11844,N_10126,N_10997);
nor U11845 (N_11845,N_10438,N_10769);
nor U11846 (N_11846,N_10966,N_10573);
or U11847 (N_11847,N_10791,N_10007);
or U11848 (N_11848,N_10898,N_10271);
nor U11849 (N_11849,N_10646,N_10405);
and U11850 (N_11850,N_10321,N_10541);
nor U11851 (N_11851,N_10803,N_10756);
or U11852 (N_11852,N_10386,N_10821);
nand U11853 (N_11853,N_10241,N_10506);
nand U11854 (N_11854,N_10213,N_10384);
nor U11855 (N_11855,N_10873,N_10100);
nand U11856 (N_11856,N_10457,N_10994);
or U11857 (N_11857,N_10153,N_10193);
and U11858 (N_11858,N_10010,N_10046);
nand U11859 (N_11859,N_10286,N_10911);
or U11860 (N_11860,N_10624,N_10838);
or U11861 (N_11861,N_10085,N_10646);
nor U11862 (N_11862,N_10291,N_10099);
or U11863 (N_11863,N_10435,N_10729);
or U11864 (N_11864,N_10836,N_10687);
xor U11865 (N_11865,N_10766,N_10654);
xnor U11866 (N_11866,N_10214,N_10140);
nor U11867 (N_11867,N_10026,N_10198);
xor U11868 (N_11868,N_10906,N_10625);
and U11869 (N_11869,N_10863,N_10447);
nand U11870 (N_11870,N_10401,N_10559);
or U11871 (N_11871,N_10292,N_10815);
and U11872 (N_11872,N_10459,N_10925);
or U11873 (N_11873,N_10815,N_10799);
xnor U11874 (N_11874,N_10097,N_10285);
nand U11875 (N_11875,N_10300,N_10691);
nand U11876 (N_11876,N_10012,N_10380);
nor U11877 (N_11877,N_10518,N_10606);
nor U11878 (N_11878,N_10693,N_10356);
and U11879 (N_11879,N_10678,N_10020);
and U11880 (N_11880,N_10461,N_10431);
and U11881 (N_11881,N_10720,N_10647);
nor U11882 (N_11882,N_10381,N_10183);
nand U11883 (N_11883,N_10880,N_10138);
or U11884 (N_11884,N_10873,N_10216);
xnor U11885 (N_11885,N_10218,N_10882);
nand U11886 (N_11886,N_10213,N_10376);
nor U11887 (N_11887,N_10372,N_10024);
xnor U11888 (N_11888,N_10114,N_10686);
and U11889 (N_11889,N_10434,N_10130);
and U11890 (N_11890,N_10607,N_10524);
xor U11891 (N_11891,N_10969,N_10338);
nand U11892 (N_11892,N_10942,N_10782);
nand U11893 (N_11893,N_10506,N_10135);
nand U11894 (N_11894,N_10245,N_10752);
nor U11895 (N_11895,N_10758,N_10815);
nor U11896 (N_11896,N_10218,N_10388);
xor U11897 (N_11897,N_10691,N_10185);
nand U11898 (N_11898,N_10507,N_10956);
xnor U11899 (N_11899,N_10425,N_10134);
and U11900 (N_11900,N_10673,N_10891);
nor U11901 (N_11901,N_10556,N_10112);
xor U11902 (N_11902,N_10671,N_10446);
and U11903 (N_11903,N_10607,N_10866);
xor U11904 (N_11904,N_10305,N_10490);
xnor U11905 (N_11905,N_10055,N_10232);
nor U11906 (N_11906,N_10755,N_10717);
nand U11907 (N_11907,N_10638,N_10885);
or U11908 (N_11908,N_10149,N_10784);
xor U11909 (N_11909,N_10924,N_10714);
and U11910 (N_11910,N_10185,N_10258);
and U11911 (N_11911,N_10421,N_10611);
xnor U11912 (N_11912,N_10661,N_10547);
or U11913 (N_11913,N_10725,N_10559);
xnor U11914 (N_11914,N_10713,N_10176);
xor U11915 (N_11915,N_10299,N_10106);
nor U11916 (N_11916,N_10734,N_10671);
nor U11917 (N_11917,N_10437,N_10886);
nand U11918 (N_11918,N_10220,N_10735);
or U11919 (N_11919,N_10549,N_10477);
xnor U11920 (N_11920,N_10892,N_10524);
or U11921 (N_11921,N_10354,N_10437);
nor U11922 (N_11922,N_10134,N_10131);
nor U11923 (N_11923,N_10898,N_10924);
nand U11924 (N_11924,N_10608,N_10207);
nand U11925 (N_11925,N_10644,N_10815);
xor U11926 (N_11926,N_10652,N_10304);
or U11927 (N_11927,N_10621,N_10867);
and U11928 (N_11928,N_10216,N_10569);
nand U11929 (N_11929,N_10386,N_10564);
or U11930 (N_11930,N_10312,N_10898);
xnor U11931 (N_11931,N_10578,N_10747);
nand U11932 (N_11932,N_10585,N_10275);
or U11933 (N_11933,N_10736,N_10726);
or U11934 (N_11934,N_10095,N_10909);
nor U11935 (N_11935,N_10498,N_10651);
nand U11936 (N_11936,N_10476,N_10017);
xor U11937 (N_11937,N_10042,N_10696);
or U11938 (N_11938,N_10058,N_10324);
nor U11939 (N_11939,N_10397,N_10593);
nand U11940 (N_11940,N_10162,N_10346);
or U11941 (N_11941,N_10574,N_10463);
or U11942 (N_11942,N_10908,N_10154);
or U11943 (N_11943,N_10065,N_10628);
nand U11944 (N_11944,N_10853,N_10174);
nor U11945 (N_11945,N_10696,N_10939);
or U11946 (N_11946,N_10983,N_10728);
and U11947 (N_11947,N_10992,N_10132);
xor U11948 (N_11948,N_10170,N_10295);
nor U11949 (N_11949,N_10536,N_10169);
nor U11950 (N_11950,N_10926,N_10778);
nand U11951 (N_11951,N_10940,N_10226);
or U11952 (N_11952,N_10080,N_10620);
or U11953 (N_11953,N_10671,N_10490);
xor U11954 (N_11954,N_10685,N_10891);
and U11955 (N_11955,N_10958,N_10234);
or U11956 (N_11956,N_10758,N_10041);
or U11957 (N_11957,N_10561,N_10898);
xnor U11958 (N_11958,N_10930,N_10779);
and U11959 (N_11959,N_10594,N_10217);
nand U11960 (N_11960,N_10187,N_10994);
or U11961 (N_11961,N_10030,N_10701);
nand U11962 (N_11962,N_10956,N_10059);
nand U11963 (N_11963,N_10506,N_10895);
nor U11964 (N_11964,N_10183,N_10670);
nor U11965 (N_11965,N_10725,N_10393);
and U11966 (N_11966,N_10345,N_10979);
nor U11967 (N_11967,N_10631,N_10146);
nor U11968 (N_11968,N_10002,N_10298);
xnor U11969 (N_11969,N_10522,N_10247);
nor U11970 (N_11970,N_10475,N_10327);
nand U11971 (N_11971,N_10035,N_10875);
nand U11972 (N_11972,N_10537,N_10172);
and U11973 (N_11973,N_10443,N_10899);
nor U11974 (N_11974,N_10281,N_10072);
or U11975 (N_11975,N_10399,N_10970);
nand U11976 (N_11976,N_10954,N_10294);
nand U11977 (N_11977,N_10793,N_10379);
nor U11978 (N_11978,N_10641,N_10116);
and U11979 (N_11979,N_10692,N_10487);
nor U11980 (N_11980,N_10816,N_10046);
and U11981 (N_11981,N_10462,N_10862);
xnor U11982 (N_11982,N_10512,N_10574);
and U11983 (N_11983,N_10086,N_10147);
or U11984 (N_11984,N_10960,N_10512);
or U11985 (N_11985,N_10767,N_10850);
and U11986 (N_11986,N_10550,N_10720);
xor U11987 (N_11987,N_10384,N_10011);
and U11988 (N_11988,N_10949,N_10769);
and U11989 (N_11989,N_10750,N_10051);
xnor U11990 (N_11990,N_10167,N_10777);
or U11991 (N_11991,N_10765,N_10715);
xor U11992 (N_11992,N_10191,N_10299);
nor U11993 (N_11993,N_10521,N_10625);
and U11994 (N_11994,N_10644,N_10236);
and U11995 (N_11995,N_10719,N_10189);
or U11996 (N_11996,N_10115,N_10215);
nand U11997 (N_11997,N_10639,N_10299);
or U11998 (N_11998,N_10938,N_10114);
and U11999 (N_11999,N_10211,N_10419);
nand U12000 (N_12000,N_11155,N_11583);
nor U12001 (N_12001,N_11611,N_11331);
nand U12002 (N_12002,N_11567,N_11685);
xor U12003 (N_12003,N_11867,N_11191);
xnor U12004 (N_12004,N_11555,N_11767);
xnor U12005 (N_12005,N_11438,N_11037);
xnor U12006 (N_12006,N_11104,N_11640);
nor U12007 (N_12007,N_11241,N_11355);
or U12008 (N_12008,N_11282,N_11718);
nor U12009 (N_12009,N_11961,N_11372);
xnor U12010 (N_12010,N_11008,N_11986);
or U12011 (N_12011,N_11928,N_11023);
nand U12012 (N_12012,N_11464,N_11553);
xnor U12013 (N_12013,N_11073,N_11277);
or U12014 (N_12014,N_11914,N_11145);
nor U12015 (N_12015,N_11550,N_11947);
or U12016 (N_12016,N_11100,N_11044);
xor U12017 (N_12017,N_11667,N_11076);
nor U12018 (N_12018,N_11597,N_11060);
nor U12019 (N_12019,N_11637,N_11224);
nor U12020 (N_12020,N_11662,N_11527);
nor U12021 (N_12021,N_11210,N_11967);
or U12022 (N_12022,N_11619,N_11242);
and U12023 (N_12023,N_11883,N_11252);
and U12024 (N_12024,N_11546,N_11432);
and U12025 (N_12025,N_11433,N_11194);
xnor U12026 (N_12026,N_11134,N_11494);
xnor U12027 (N_12027,N_11805,N_11370);
xor U12028 (N_12028,N_11906,N_11946);
or U12029 (N_12029,N_11207,N_11084);
and U12030 (N_12030,N_11554,N_11700);
nand U12031 (N_12031,N_11781,N_11657);
and U12032 (N_12032,N_11113,N_11186);
nor U12033 (N_12033,N_11047,N_11660);
or U12034 (N_12034,N_11424,N_11580);
and U12035 (N_12035,N_11158,N_11212);
xor U12036 (N_12036,N_11358,N_11603);
and U12037 (N_12037,N_11740,N_11534);
or U12038 (N_12038,N_11369,N_11541);
nor U12039 (N_12039,N_11639,N_11498);
nand U12040 (N_12040,N_11617,N_11146);
or U12041 (N_12041,N_11049,N_11788);
nand U12042 (N_12042,N_11338,N_11397);
nand U12043 (N_12043,N_11074,N_11556);
xor U12044 (N_12044,N_11579,N_11670);
nor U12045 (N_12045,N_11663,N_11326);
xor U12046 (N_12046,N_11343,N_11653);
xor U12047 (N_12047,N_11709,N_11460);
or U12048 (N_12048,N_11209,N_11802);
or U12049 (N_12049,N_11320,N_11190);
xnor U12050 (N_12050,N_11441,N_11193);
or U12051 (N_12051,N_11835,N_11184);
xor U12052 (N_12052,N_11834,N_11121);
nand U12053 (N_12053,N_11226,N_11129);
xor U12054 (N_12054,N_11022,N_11264);
xnor U12055 (N_12055,N_11631,N_11988);
nor U12056 (N_12056,N_11148,N_11801);
xor U12057 (N_12057,N_11674,N_11466);
or U12058 (N_12058,N_11572,N_11062);
or U12059 (N_12059,N_11087,N_11502);
xor U12060 (N_12060,N_11717,N_11010);
and U12061 (N_12061,N_11292,N_11475);
xor U12062 (N_12062,N_11566,N_11719);
nor U12063 (N_12063,N_11707,N_11735);
or U12064 (N_12064,N_11691,N_11544);
nor U12065 (N_12065,N_11123,N_11283);
or U12066 (N_12066,N_11849,N_11228);
or U12067 (N_12067,N_11564,N_11658);
and U12068 (N_12068,N_11253,N_11759);
or U12069 (N_12069,N_11723,N_11540);
nor U12070 (N_12070,N_11783,N_11257);
nor U12071 (N_12071,N_11858,N_11793);
nand U12072 (N_12072,N_11319,N_11995);
or U12073 (N_12073,N_11911,N_11945);
nor U12074 (N_12074,N_11205,N_11161);
and U12075 (N_12075,N_11736,N_11482);
or U12076 (N_12076,N_11059,N_11144);
xnor U12077 (N_12077,N_11888,N_11633);
and U12078 (N_12078,N_11672,N_11978);
xor U12079 (N_12079,N_11636,N_11795);
nor U12080 (N_12080,N_11837,N_11462);
nor U12081 (N_12081,N_11714,N_11818);
nor U12082 (N_12082,N_11671,N_11913);
xnor U12083 (N_12083,N_11558,N_11728);
xor U12084 (N_12084,N_11430,N_11752);
xnor U12085 (N_12085,N_11233,N_11125);
and U12086 (N_12086,N_11627,N_11136);
or U12087 (N_12087,N_11428,N_11015);
and U12088 (N_12088,N_11598,N_11479);
xnor U12089 (N_12089,N_11698,N_11530);
and U12090 (N_12090,N_11846,N_11298);
or U12091 (N_12091,N_11042,N_11046);
or U12092 (N_12092,N_11970,N_11181);
and U12093 (N_12093,N_11313,N_11293);
nor U12094 (N_12094,N_11920,N_11061);
xnor U12095 (N_12095,N_11923,N_11153);
nand U12096 (N_12096,N_11632,N_11289);
xnor U12097 (N_12097,N_11827,N_11528);
nand U12098 (N_12098,N_11962,N_11826);
and U12099 (N_12099,N_11879,N_11526);
and U12100 (N_12100,N_11615,N_11870);
or U12101 (N_12101,N_11532,N_11993);
nand U12102 (N_12102,N_11085,N_11725);
or U12103 (N_12103,N_11236,N_11905);
nor U12104 (N_12104,N_11608,N_11654);
nor U12105 (N_12105,N_11418,N_11976);
nand U12106 (N_12106,N_11072,N_11692);
or U12107 (N_12107,N_11545,N_11756);
nand U12108 (N_12108,N_11940,N_11377);
nor U12109 (N_12109,N_11106,N_11206);
nand U12110 (N_12110,N_11089,N_11351);
or U12111 (N_12111,N_11130,N_11864);
or U12112 (N_12112,N_11394,N_11956);
or U12113 (N_12113,N_11465,N_11291);
or U12114 (N_12114,N_11529,N_11794);
nor U12115 (N_12115,N_11701,N_11081);
and U12116 (N_12116,N_11522,N_11889);
or U12117 (N_12117,N_11408,N_11804);
or U12118 (N_12118,N_11678,N_11609);
nand U12119 (N_12119,N_11406,N_11285);
nand U12120 (N_12120,N_11222,N_11025);
or U12121 (N_12121,N_11679,N_11485);
nor U12122 (N_12122,N_11099,N_11594);
or U12123 (N_12123,N_11885,N_11859);
xnor U12124 (N_12124,N_11776,N_11684);
and U12125 (N_12125,N_11996,N_11028);
nor U12126 (N_12126,N_11635,N_11014);
and U12127 (N_12127,N_11551,N_11387);
or U12128 (N_12128,N_11624,N_11862);
xnor U12129 (N_12129,N_11668,N_11899);
and U12130 (N_12130,N_11588,N_11830);
nand U12131 (N_12131,N_11401,N_11216);
nor U12132 (N_12132,N_11951,N_11132);
or U12133 (N_12133,N_11949,N_11872);
or U12134 (N_12134,N_11841,N_11822);
xor U12135 (N_12135,N_11751,N_11021);
nand U12136 (N_12136,N_11045,N_11012);
nor U12137 (N_12137,N_11708,N_11673);
and U12138 (N_12138,N_11223,N_11798);
nand U12139 (N_12139,N_11971,N_11703);
xor U12140 (N_12140,N_11601,N_11655);
nor U12141 (N_12141,N_11890,N_11080);
or U12142 (N_12142,N_11437,N_11417);
nand U12143 (N_12143,N_11459,N_11542);
or U12144 (N_12144,N_11771,N_11218);
nand U12145 (N_12145,N_11427,N_11070);
nand U12146 (N_12146,N_11071,N_11489);
nor U12147 (N_12147,N_11543,N_11288);
xor U12148 (N_12148,N_11449,N_11569);
nand U12149 (N_12149,N_11120,N_11515);
nor U12150 (N_12150,N_11024,N_11237);
or U12151 (N_12151,N_11434,N_11690);
nor U12152 (N_12152,N_11274,N_11742);
or U12153 (N_12153,N_11832,N_11367);
nand U12154 (N_12154,N_11450,N_11315);
and U12155 (N_12155,N_11296,N_11769);
nand U12156 (N_12156,N_11651,N_11182);
xnor U12157 (N_12157,N_11931,N_11112);
nand U12158 (N_12158,N_11816,N_11322);
or U12159 (N_12159,N_11164,N_11918);
and U12160 (N_12160,N_11360,N_11741);
xor U12161 (N_12161,N_11357,N_11792);
xor U12162 (N_12162,N_11552,N_11189);
xnor U12163 (N_12163,N_11470,N_11912);
nand U12164 (N_12164,N_11431,N_11626);
nor U12165 (N_12165,N_11170,N_11269);
nand U12166 (N_12166,N_11254,N_11681);
nand U12167 (N_12167,N_11704,N_11699);
or U12168 (N_12168,N_11166,N_11768);
or U12169 (N_12169,N_11629,N_11442);
xnor U12170 (N_12170,N_11991,N_11812);
nor U12171 (N_12171,N_11900,N_11981);
nor U12172 (N_12172,N_11052,N_11443);
nor U12173 (N_12173,N_11304,N_11004);
and U12174 (N_12174,N_11131,N_11686);
nand U12175 (N_12175,N_11126,N_11957);
or U12176 (N_12176,N_11151,N_11796);
and U12177 (N_12177,N_11732,N_11456);
nand U12178 (N_12178,N_11229,N_11235);
nor U12179 (N_12179,N_11371,N_11623);
or U12180 (N_12180,N_11875,N_11921);
or U12181 (N_12181,N_11138,N_11032);
and U12182 (N_12182,N_11458,N_11874);
or U12183 (N_12183,N_11392,N_11180);
nand U12184 (N_12184,N_11279,N_11263);
nor U12185 (N_12185,N_11001,N_11851);
nor U12186 (N_12186,N_11806,N_11917);
nor U12187 (N_12187,N_11219,N_11018);
xor U12188 (N_12188,N_11747,N_11095);
nor U12189 (N_12189,N_11630,N_11203);
nand U12190 (N_12190,N_11341,N_11535);
nor U12191 (N_12191,N_11390,N_11117);
nand U12192 (N_12192,N_11969,N_11848);
xnor U12193 (N_12193,N_11726,N_11102);
xnor U12194 (N_12194,N_11512,N_11782);
and U12195 (N_12195,N_11273,N_11097);
nand U12196 (N_12196,N_11472,N_11185);
and U12197 (N_12197,N_11380,N_11828);
xnor U12198 (N_12198,N_11077,N_11634);
nand U12199 (N_12199,N_11362,N_11628);
or U12200 (N_12200,N_11780,N_11810);
nor U12201 (N_12201,N_11706,N_11041);
nand U12202 (N_12202,N_11952,N_11038);
and U12203 (N_12203,N_11729,N_11960);
nand U12204 (N_12204,N_11347,N_11169);
and U12205 (N_12205,N_11399,N_11737);
nand U12206 (N_12206,N_11549,N_11262);
xnor U12207 (N_12207,N_11944,N_11666);
nor U12208 (N_12208,N_11075,N_11027);
nor U12209 (N_12209,N_11348,N_11410);
nor U12210 (N_12210,N_11589,N_11333);
or U12211 (N_12211,N_11255,N_11391);
nand U12212 (N_12212,N_11019,N_11559);
xnor U12213 (N_12213,N_11402,N_11215);
xor U12214 (N_12214,N_11510,N_11919);
nand U12215 (N_12215,N_11924,N_11114);
nand U12216 (N_12216,N_11335,N_11689);
or U12217 (N_12217,N_11163,N_11328);
or U12218 (N_12218,N_11090,N_11855);
xnor U12219 (N_12219,N_11484,N_11268);
nor U12220 (N_12220,N_11429,N_11213);
nand U12221 (N_12221,N_11620,N_11468);
nand U12222 (N_12222,N_11746,N_11982);
nor U12223 (N_12223,N_11734,N_11648);
nand U12224 (N_12224,N_11111,N_11448);
nor U12225 (N_12225,N_11499,N_11492);
or U12226 (N_12226,N_11514,N_11451);
nand U12227 (N_12227,N_11755,N_11260);
nand U12228 (N_12228,N_11122,N_11842);
xor U12229 (N_12229,N_11426,N_11115);
nor U12230 (N_12230,N_11356,N_11403);
xnor U12231 (N_12231,N_11378,N_11892);
or U12232 (N_12232,N_11000,N_11656);
xor U12233 (N_12233,N_11150,N_11318);
and U12234 (N_12234,N_11440,N_11258);
nand U12235 (N_12235,N_11251,N_11325);
nand U12236 (N_12236,N_11301,N_11705);
or U12237 (N_12237,N_11720,N_11474);
or U12238 (N_12238,N_11645,N_11927);
or U12239 (N_12239,N_11584,N_11244);
nand U12240 (N_12240,N_11531,N_11230);
or U12241 (N_12241,N_11606,N_11607);
and U12242 (N_12242,N_11329,N_11141);
xnor U12243 (N_12243,N_11006,N_11710);
xnor U12244 (N_12244,N_11571,N_11772);
or U12245 (N_12245,N_11058,N_11143);
nand U12246 (N_12246,N_11473,N_11382);
xor U12247 (N_12247,N_11963,N_11715);
nand U12248 (N_12248,N_11523,N_11702);
or U12249 (N_12249,N_11724,N_11647);
or U12250 (N_12250,N_11649,N_11513);
nand U12251 (N_12251,N_11777,N_11078);
nor U12252 (N_12252,N_11953,N_11094);
xor U12253 (N_12253,N_11677,N_11965);
nor U12254 (N_12254,N_11831,N_11248);
nand U12255 (N_12255,N_11891,N_11204);
xor U12256 (N_12256,N_11033,N_11487);
xor U12257 (N_12257,N_11561,N_11933);
nand U12258 (N_12258,N_11789,N_11172);
and U12259 (N_12259,N_11659,N_11261);
or U12260 (N_12260,N_11761,N_11035);
and U12261 (N_12261,N_11415,N_11560);
nor U12262 (N_12262,N_11147,N_11086);
and U12263 (N_12263,N_11939,N_11625);
nor U12264 (N_12264,N_11853,N_11435);
xor U12265 (N_12265,N_11275,N_11152);
nand U12266 (N_12266,N_11198,N_11687);
xor U12267 (N_12267,N_11570,N_11770);
and U12268 (N_12268,N_11524,N_11446);
nor U12269 (N_12269,N_11844,N_11766);
nor U12270 (N_12270,N_11056,N_11250);
and U12271 (N_12271,N_11866,N_11124);
nor U12272 (N_12272,N_11276,N_11243);
nand U12273 (N_12273,N_11290,N_11165);
xnor U12274 (N_12274,N_11160,N_11385);
nand U12275 (N_12275,N_11861,N_11488);
xor U12276 (N_12276,N_11299,N_11171);
nand U12277 (N_12277,N_11503,N_11868);
nor U12278 (N_12278,N_11508,N_11950);
xnor U12279 (N_12279,N_11716,N_11463);
nor U12280 (N_12280,N_11157,N_11800);
or U12281 (N_12281,N_11817,N_11994);
xnor U12282 (N_12282,N_11383,N_11066);
nand U12283 (N_12283,N_11587,N_11833);
nor U12284 (N_12284,N_11353,N_11799);
xnor U12285 (N_12285,N_11763,N_11652);
nor U12286 (N_12286,N_11865,N_11774);
or U12287 (N_12287,N_11187,N_11232);
and U12288 (N_12288,N_11154,N_11936);
xor U12289 (N_12289,N_11003,N_11398);
nand U12290 (N_12290,N_11031,N_11739);
nand U12291 (N_12291,N_11054,N_11665);
nor U12292 (N_12292,N_11361,N_11188);
and U12293 (N_12293,N_11365,N_11178);
or U12294 (N_12294,N_11309,N_11231);
xnor U12295 (N_12295,N_11536,N_11803);
nor U12296 (N_12296,N_11682,N_11156);
nand U12297 (N_12297,N_11096,N_11176);
nor U12298 (N_12298,N_11688,N_11174);
nor U12299 (N_12299,N_11083,N_11177);
xor U12300 (N_12300,N_11352,N_11979);
and U12301 (N_12301,N_11020,N_11893);
nand U12302 (N_12302,N_11926,N_11646);
xor U12303 (N_12303,N_11311,N_11305);
and U12304 (N_12304,N_11461,N_11310);
nand U12305 (N_12305,N_11297,N_11932);
nor U12306 (N_12306,N_11467,N_11887);
or U12307 (N_12307,N_11878,N_11985);
or U12308 (N_12308,N_11909,N_11200);
nor U12309 (N_12309,N_11839,N_11040);
and U12310 (N_12310,N_11373,N_11116);
nand U12311 (N_12311,N_11696,N_11501);
nor U12312 (N_12312,N_11139,N_11057);
or U12313 (N_12313,N_11234,N_11324);
or U12314 (N_12314,N_11405,N_11471);
nor U12315 (N_12315,N_11481,N_11693);
or U12316 (N_12316,N_11695,N_11504);
and U12317 (N_12317,N_11168,N_11330);
nand U12318 (N_12318,N_11088,N_11421);
nand U12319 (N_12319,N_11053,N_11517);
nand U12320 (N_12320,N_11642,N_11337);
nand U12321 (N_12321,N_11622,N_11539);
and U12322 (N_12322,N_11030,N_11857);
or U12323 (N_12323,N_11109,N_11439);
nor U12324 (N_12324,N_11955,N_11175);
or U12325 (N_12325,N_11069,N_11135);
nor U12326 (N_12326,N_11342,N_11880);
and U12327 (N_12327,N_11916,N_11368);
nand U12328 (N_12328,N_11786,N_11643);
and U12329 (N_12329,N_11675,N_11287);
nor U12330 (N_12330,N_11295,N_11445);
nand U12331 (N_12331,N_11613,N_11847);
nor U12332 (N_12332,N_11730,N_11454);
nor U12333 (N_12333,N_11101,N_11596);
or U12334 (N_12334,N_11127,N_11974);
xnor U12335 (N_12335,N_11413,N_11948);
or U12336 (N_12336,N_11904,N_11850);
nand U12337 (N_12337,N_11079,N_11349);
xnor U12338 (N_12338,N_11563,N_11807);
and U12339 (N_12339,N_11029,N_11201);
nor U12340 (N_12340,N_11221,N_11829);
xor U12341 (N_12341,N_11159,N_11068);
nor U12342 (N_12342,N_11860,N_11749);
nand U12343 (N_12343,N_11898,N_11323);
nor U12344 (N_12344,N_11825,N_11050);
or U12345 (N_12345,N_11843,N_11882);
and U12346 (N_12346,N_11496,N_11345);
xor U12347 (N_12347,N_11453,N_11067);
xor U12348 (N_12348,N_11266,N_11676);
or U12349 (N_12349,N_11196,N_11091);
nand U12350 (N_12350,N_11336,N_11217);
nor U12351 (N_12351,N_11854,N_11618);
nor U12352 (N_12352,N_11975,N_11903);
and U12353 (N_12353,N_11308,N_11452);
nand U12354 (N_12354,N_11821,N_11002);
or U12355 (N_12355,N_11977,N_11162);
xnor U12356 (N_12356,N_11350,N_11108);
nor U12357 (N_12357,N_11585,N_11744);
nand U12358 (N_12358,N_11983,N_11354);
nand U12359 (N_12359,N_11852,N_11519);
xor U12360 (N_12360,N_11602,N_11173);
or U12361 (N_12361,N_11884,N_11455);
nand U12362 (N_12362,N_11745,N_11007);
nor U12363 (N_12363,N_11300,N_11412);
or U12364 (N_12364,N_11576,N_11376);
nor U12365 (N_12365,N_11110,N_11396);
xnor U12366 (N_12366,N_11959,N_11954);
xor U12367 (N_12367,N_11925,N_11063);
nor U12368 (N_12368,N_11199,N_11593);
nand U12369 (N_12369,N_11938,N_11980);
nor U12370 (N_12370,N_11284,N_11722);
nand U12371 (N_12371,N_11896,N_11227);
nor U12372 (N_12372,N_11265,N_11819);
and U12373 (N_12373,N_11727,N_11506);
or U12374 (N_12374,N_11476,N_11312);
nor U12375 (N_12375,N_11547,N_11838);
nor U12376 (N_12376,N_11537,N_11098);
xnor U12377 (N_12377,N_11915,N_11516);
nand U12378 (N_12378,N_11208,N_11497);
or U12379 (N_12379,N_11582,N_11239);
or U12380 (N_12380,N_11565,N_11784);
xnor U12381 (N_12381,N_11605,N_11886);
nor U12382 (N_12382,N_11824,N_11743);
nand U12383 (N_12383,N_11409,N_11366);
or U12384 (N_12384,N_11638,N_11895);
nor U12385 (N_12385,N_11964,N_11422);
and U12386 (N_12386,N_11577,N_11968);
and U12387 (N_12387,N_11256,N_11493);
nand U12388 (N_12388,N_11048,N_11259);
xnor U12389 (N_12389,N_11307,N_11192);
nor U12390 (N_12390,N_11065,N_11036);
and U12391 (N_12391,N_11505,N_11992);
or U12392 (N_12392,N_11581,N_11270);
xnor U12393 (N_12393,N_11480,N_11486);
nand U12394 (N_12394,N_11034,N_11721);
xor U12395 (N_12395,N_11574,N_11005);
or U12396 (N_12396,N_11578,N_11404);
or U12397 (N_12397,N_11103,N_11621);
nor U12398 (N_12398,N_11267,N_11738);
and U12399 (N_12399,N_11026,N_11495);
nor U12400 (N_12400,N_11321,N_11332);
or U12401 (N_12401,N_11317,N_11990);
xnor U12402 (N_12402,N_11764,N_11384);
nand U12403 (N_12403,N_11507,N_11225);
nor U12404 (N_12404,N_11051,N_11140);
nor U12405 (N_12405,N_11416,N_11245);
xor U12406 (N_12406,N_11680,N_11573);
or U12407 (N_12407,N_11082,N_11302);
and U12408 (N_12408,N_11779,N_11910);
xor U12409 (N_12409,N_11568,N_11845);
and U12410 (N_12410,N_11444,N_11610);
and U12411 (N_12411,N_11599,N_11500);
nor U12412 (N_12412,N_11694,N_11395);
xor U12413 (N_12413,N_11214,N_11644);
nor U12414 (N_12414,N_11787,N_11294);
or U12415 (N_12415,N_11303,N_11871);
nor U12416 (N_12416,N_11013,N_11922);
xor U12417 (N_12417,N_11836,N_11873);
nor U12418 (N_12418,N_11591,N_11869);
or U12419 (N_12419,N_11901,N_11105);
xor U12420 (N_12420,N_11881,N_11375);
or U12421 (N_12421,N_11809,N_11785);
nor U12422 (N_12422,N_11436,N_11278);
and U12423 (N_12423,N_11183,N_11491);
nor U12424 (N_12424,N_11423,N_11929);
nand U12425 (N_12425,N_11363,N_11897);
nor U12426 (N_12426,N_11316,N_11935);
nand U12427 (N_12427,N_11790,N_11943);
or U12428 (N_12428,N_11364,N_11483);
and U12429 (N_12429,N_11997,N_11958);
xor U12430 (N_12430,N_11907,N_11934);
and U12431 (N_12431,N_11388,N_11757);
nor U12432 (N_12432,N_11521,N_11937);
nor U12433 (N_12433,N_11393,N_11195);
nor U12434 (N_12434,N_11762,N_11359);
or U12435 (N_12435,N_11733,N_11509);
nor U12436 (N_12436,N_11477,N_11211);
xor U12437 (N_12437,N_11490,N_11791);
nand U12438 (N_12438,N_11856,N_11064);
xor U12439 (N_12439,N_11016,N_11661);
and U12440 (N_12440,N_11586,N_11093);
xnor U12441 (N_12441,N_11683,N_11039);
and U12442 (N_12442,N_11840,N_11966);
or U12443 (N_12443,N_11246,N_11760);
and U12444 (N_12444,N_11815,N_11137);
nand U12445 (N_12445,N_11107,N_11055);
nand U12446 (N_12446,N_11820,N_11011);
and U12447 (N_12447,N_11457,N_11149);
nand U12448 (N_12448,N_11314,N_11179);
xnor U12449 (N_12449,N_11711,N_11592);
xor U12450 (N_12450,N_11469,N_11411);
or U12451 (N_12451,N_11754,N_11972);
or U12452 (N_12452,N_11425,N_11281);
or U12453 (N_12453,N_11043,N_11984);
and U12454 (N_12454,N_11942,N_11750);
nor U12455 (N_12455,N_11520,N_11327);
xor U12456 (N_12456,N_11518,N_11389);
nor U12457 (N_12457,N_11773,N_11557);
and U12458 (N_12458,N_11753,N_11202);
nand U12459 (N_12459,N_11344,N_11220);
nand U12460 (N_12460,N_11346,N_11197);
nor U12461 (N_12461,N_11511,N_11877);
nor U12462 (N_12462,N_11876,N_11538);
and U12463 (N_12463,N_11811,N_11562);
nand U12464 (N_12464,N_11009,N_11590);
xnor U12465 (N_12465,N_11650,N_11271);
nor U12466 (N_12466,N_11758,N_11616);
nand U12467 (N_12467,N_11533,N_11600);
xnor U12468 (N_12468,N_11930,N_11167);
xor U12469 (N_12469,N_11669,N_11697);
nor U12470 (N_12470,N_11419,N_11973);
nor U12471 (N_12471,N_11386,N_11092);
nand U12472 (N_12472,N_11713,N_11614);
or U12473 (N_12473,N_11340,N_11118);
nor U12474 (N_12474,N_11414,N_11612);
nor U12475 (N_12475,N_11119,N_11379);
nor U12476 (N_12476,N_11142,N_11778);
nor U12477 (N_12477,N_11775,N_11420);
and U12478 (N_12478,N_11823,N_11249);
or U12479 (N_12479,N_11731,N_11797);
and U12480 (N_12480,N_11447,N_11133);
xnor U12481 (N_12481,N_11999,N_11575);
xor U12482 (N_12482,N_11664,N_11908);
nor U12483 (N_12483,N_11813,N_11765);
xor U12484 (N_12484,N_11604,N_11478);
xor U12485 (N_12485,N_11548,N_11240);
nand U12486 (N_12486,N_11339,N_11238);
nor U12487 (N_12487,N_11808,N_11863);
nand U12488 (N_12488,N_11272,N_11941);
or U12489 (N_12489,N_11525,N_11998);
xnor U12490 (N_12490,N_11374,N_11128);
nand U12491 (N_12491,N_11381,N_11902);
and U12492 (N_12492,N_11407,N_11400);
xnor U12493 (N_12493,N_11894,N_11987);
or U12494 (N_12494,N_11712,N_11814);
nand U12495 (N_12495,N_11595,N_11280);
nand U12496 (N_12496,N_11306,N_11989);
xor U12497 (N_12497,N_11017,N_11641);
or U12498 (N_12498,N_11247,N_11286);
nor U12499 (N_12499,N_11748,N_11334);
nand U12500 (N_12500,N_11864,N_11561);
or U12501 (N_12501,N_11455,N_11619);
or U12502 (N_12502,N_11669,N_11821);
nor U12503 (N_12503,N_11722,N_11498);
or U12504 (N_12504,N_11874,N_11548);
nor U12505 (N_12505,N_11068,N_11644);
nor U12506 (N_12506,N_11906,N_11024);
or U12507 (N_12507,N_11257,N_11207);
or U12508 (N_12508,N_11287,N_11460);
xor U12509 (N_12509,N_11747,N_11124);
or U12510 (N_12510,N_11407,N_11833);
xnor U12511 (N_12511,N_11480,N_11643);
xor U12512 (N_12512,N_11994,N_11500);
xor U12513 (N_12513,N_11568,N_11883);
xnor U12514 (N_12514,N_11532,N_11794);
xnor U12515 (N_12515,N_11428,N_11693);
nor U12516 (N_12516,N_11052,N_11284);
nand U12517 (N_12517,N_11028,N_11781);
nor U12518 (N_12518,N_11628,N_11291);
xnor U12519 (N_12519,N_11405,N_11376);
nor U12520 (N_12520,N_11251,N_11361);
xnor U12521 (N_12521,N_11789,N_11323);
and U12522 (N_12522,N_11444,N_11254);
xor U12523 (N_12523,N_11129,N_11344);
and U12524 (N_12524,N_11590,N_11534);
nor U12525 (N_12525,N_11780,N_11717);
and U12526 (N_12526,N_11530,N_11152);
or U12527 (N_12527,N_11874,N_11780);
nand U12528 (N_12528,N_11794,N_11278);
nand U12529 (N_12529,N_11805,N_11248);
nand U12530 (N_12530,N_11597,N_11385);
or U12531 (N_12531,N_11212,N_11121);
nand U12532 (N_12532,N_11806,N_11317);
nand U12533 (N_12533,N_11967,N_11102);
and U12534 (N_12534,N_11327,N_11212);
nand U12535 (N_12535,N_11456,N_11385);
xnor U12536 (N_12536,N_11764,N_11787);
or U12537 (N_12537,N_11736,N_11305);
xor U12538 (N_12538,N_11315,N_11674);
nor U12539 (N_12539,N_11079,N_11898);
and U12540 (N_12540,N_11744,N_11919);
nand U12541 (N_12541,N_11322,N_11694);
nand U12542 (N_12542,N_11278,N_11833);
or U12543 (N_12543,N_11474,N_11775);
or U12544 (N_12544,N_11332,N_11625);
or U12545 (N_12545,N_11153,N_11366);
nand U12546 (N_12546,N_11121,N_11264);
xnor U12547 (N_12547,N_11766,N_11353);
xnor U12548 (N_12548,N_11102,N_11581);
and U12549 (N_12549,N_11896,N_11785);
nand U12550 (N_12550,N_11836,N_11474);
and U12551 (N_12551,N_11778,N_11506);
or U12552 (N_12552,N_11538,N_11665);
nor U12553 (N_12553,N_11148,N_11909);
nand U12554 (N_12554,N_11537,N_11368);
xor U12555 (N_12555,N_11063,N_11833);
or U12556 (N_12556,N_11454,N_11838);
and U12557 (N_12557,N_11292,N_11061);
and U12558 (N_12558,N_11661,N_11640);
and U12559 (N_12559,N_11711,N_11832);
nand U12560 (N_12560,N_11080,N_11565);
xor U12561 (N_12561,N_11568,N_11171);
nor U12562 (N_12562,N_11625,N_11976);
nand U12563 (N_12563,N_11176,N_11196);
nor U12564 (N_12564,N_11527,N_11032);
and U12565 (N_12565,N_11199,N_11533);
xnor U12566 (N_12566,N_11582,N_11082);
or U12567 (N_12567,N_11411,N_11977);
xor U12568 (N_12568,N_11974,N_11958);
or U12569 (N_12569,N_11440,N_11458);
and U12570 (N_12570,N_11760,N_11277);
or U12571 (N_12571,N_11090,N_11116);
nor U12572 (N_12572,N_11534,N_11396);
nor U12573 (N_12573,N_11035,N_11092);
and U12574 (N_12574,N_11534,N_11565);
nor U12575 (N_12575,N_11178,N_11212);
nor U12576 (N_12576,N_11817,N_11419);
or U12577 (N_12577,N_11474,N_11591);
xnor U12578 (N_12578,N_11504,N_11725);
nor U12579 (N_12579,N_11162,N_11231);
or U12580 (N_12580,N_11631,N_11496);
or U12581 (N_12581,N_11675,N_11434);
or U12582 (N_12582,N_11539,N_11399);
nor U12583 (N_12583,N_11625,N_11278);
nand U12584 (N_12584,N_11620,N_11491);
nor U12585 (N_12585,N_11931,N_11318);
nor U12586 (N_12586,N_11301,N_11557);
or U12587 (N_12587,N_11984,N_11979);
nor U12588 (N_12588,N_11953,N_11128);
nor U12589 (N_12589,N_11128,N_11439);
nand U12590 (N_12590,N_11584,N_11623);
or U12591 (N_12591,N_11186,N_11467);
nor U12592 (N_12592,N_11852,N_11792);
nand U12593 (N_12593,N_11383,N_11171);
nand U12594 (N_12594,N_11999,N_11791);
nand U12595 (N_12595,N_11286,N_11107);
or U12596 (N_12596,N_11918,N_11206);
or U12597 (N_12597,N_11068,N_11611);
nand U12598 (N_12598,N_11697,N_11019);
nand U12599 (N_12599,N_11521,N_11447);
nand U12600 (N_12600,N_11281,N_11176);
and U12601 (N_12601,N_11277,N_11382);
xor U12602 (N_12602,N_11974,N_11404);
nand U12603 (N_12603,N_11231,N_11312);
nand U12604 (N_12604,N_11667,N_11640);
xor U12605 (N_12605,N_11614,N_11883);
or U12606 (N_12606,N_11420,N_11519);
or U12607 (N_12607,N_11180,N_11954);
nand U12608 (N_12608,N_11285,N_11353);
nor U12609 (N_12609,N_11910,N_11728);
and U12610 (N_12610,N_11343,N_11028);
nor U12611 (N_12611,N_11402,N_11346);
nand U12612 (N_12612,N_11451,N_11526);
nor U12613 (N_12613,N_11070,N_11320);
xor U12614 (N_12614,N_11331,N_11231);
nand U12615 (N_12615,N_11167,N_11670);
nand U12616 (N_12616,N_11784,N_11332);
nand U12617 (N_12617,N_11459,N_11266);
nand U12618 (N_12618,N_11863,N_11533);
and U12619 (N_12619,N_11707,N_11788);
xnor U12620 (N_12620,N_11872,N_11868);
nand U12621 (N_12621,N_11579,N_11201);
nand U12622 (N_12622,N_11393,N_11776);
nand U12623 (N_12623,N_11219,N_11464);
or U12624 (N_12624,N_11404,N_11055);
nand U12625 (N_12625,N_11628,N_11959);
or U12626 (N_12626,N_11110,N_11440);
or U12627 (N_12627,N_11249,N_11074);
nand U12628 (N_12628,N_11833,N_11491);
xnor U12629 (N_12629,N_11036,N_11681);
xnor U12630 (N_12630,N_11439,N_11646);
nand U12631 (N_12631,N_11455,N_11715);
nor U12632 (N_12632,N_11410,N_11083);
xor U12633 (N_12633,N_11102,N_11768);
xnor U12634 (N_12634,N_11477,N_11501);
and U12635 (N_12635,N_11960,N_11721);
or U12636 (N_12636,N_11810,N_11311);
and U12637 (N_12637,N_11702,N_11142);
xnor U12638 (N_12638,N_11848,N_11557);
xnor U12639 (N_12639,N_11100,N_11795);
and U12640 (N_12640,N_11713,N_11703);
nor U12641 (N_12641,N_11087,N_11101);
nand U12642 (N_12642,N_11267,N_11390);
xnor U12643 (N_12643,N_11031,N_11893);
nand U12644 (N_12644,N_11587,N_11635);
or U12645 (N_12645,N_11881,N_11945);
nor U12646 (N_12646,N_11400,N_11804);
nand U12647 (N_12647,N_11016,N_11713);
nor U12648 (N_12648,N_11832,N_11106);
nand U12649 (N_12649,N_11606,N_11745);
or U12650 (N_12650,N_11059,N_11441);
or U12651 (N_12651,N_11897,N_11158);
xor U12652 (N_12652,N_11509,N_11625);
nand U12653 (N_12653,N_11018,N_11893);
xor U12654 (N_12654,N_11530,N_11037);
nor U12655 (N_12655,N_11352,N_11307);
nand U12656 (N_12656,N_11267,N_11600);
nor U12657 (N_12657,N_11253,N_11521);
xnor U12658 (N_12658,N_11783,N_11217);
or U12659 (N_12659,N_11585,N_11718);
or U12660 (N_12660,N_11737,N_11395);
and U12661 (N_12661,N_11834,N_11659);
or U12662 (N_12662,N_11196,N_11933);
xor U12663 (N_12663,N_11332,N_11188);
nor U12664 (N_12664,N_11653,N_11124);
nand U12665 (N_12665,N_11717,N_11236);
or U12666 (N_12666,N_11856,N_11257);
nand U12667 (N_12667,N_11342,N_11355);
nand U12668 (N_12668,N_11494,N_11952);
and U12669 (N_12669,N_11182,N_11575);
xor U12670 (N_12670,N_11658,N_11541);
and U12671 (N_12671,N_11875,N_11701);
and U12672 (N_12672,N_11992,N_11392);
nand U12673 (N_12673,N_11786,N_11524);
and U12674 (N_12674,N_11368,N_11541);
or U12675 (N_12675,N_11705,N_11716);
nor U12676 (N_12676,N_11862,N_11212);
nand U12677 (N_12677,N_11095,N_11416);
nand U12678 (N_12678,N_11982,N_11456);
nor U12679 (N_12679,N_11963,N_11354);
nor U12680 (N_12680,N_11068,N_11417);
and U12681 (N_12681,N_11666,N_11505);
nand U12682 (N_12682,N_11953,N_11114);
xnor U12683 (N_12683,N_11986,N_11469);
nor U12684 (N_12684,N_11638,N_11325);
or U12685 (N_12685,N_11310,N_11792);
or U12686 (N_12686,N_11179,N_11512);
nor U12687 (N_12687,N_11422,N_11999);
nor U12688 (N_12688,N_11809,N_11748);
and U12689 (N_12689,N_11896,N_11293);
nor U12690 (N_12690,N_11977,N_11985);
xnor U12691 (N_12691,N_11514,N_11578);
nand U12692 (N_12692,N_11985,N_11715);
xor U12693 (N_12693,N_11744,N_11929);
nand U12694 (N_12694,N_11842,N_11305);
xnor U12695 (N_12695,N_11754,N_11916);
xnor U12696 (N_12696,N_11637,N_11677);
nand U12697 (N_12697,N_11795,N_11822);
or U12698 (N_12698,N_11037,N_11787);
xor U12699 (N_12699,N_11308,N_11007);
and U12700 (N_12700,N_11409,N_11403);
nand U12701 (N_12701,N_11931,N_11441);
nor U12702 (N_12702,N_11121,N_11211);
xnor U12703 (N_12703,N_11854,N_11375);
and U12704 (N_12704,N_11868,N_11569);
nor U12705 (N_12705,N_11229,N_11980);
xor U12706 (N_12706,N_11276,N_11899);
and U12707 (N_12707,N_11269,N_11299);
nor U12708 (N_12708,N_11935,N_11777);
nand U12709 (N_12709,N_11694,N_11128);
nand U12710 (N_12710,N_11727,N_11223);
nand U12711 (N_12711,N_11924,N_11330);
nor U12712 (N_12712,N_11451,N_11544);
or U12713 (N_12713,N_11505,N_11336);
xnor U12714 (N_12714,N_11862,N_11041);
or U12715 (N_12715,N_11417,N_11823);
xnor U12716 (N_12716,N_11663,N_11386);
nand U12717 (N_12717,N_11917,N_11498);
nor U12718 (N_12718,N_11566,N_11322);
and U12719 (N_12719,N_11883,N_11801);
and U12720 (N_12720,N_11406,N_11612);
nor U12721 (N_12721,N_11648,N_11505);
nand U12722 (N_12722,N_11772,N_11901);
nor U12723 (N_12723,N_11860,N_11253);
nor U12724 (N_12724,N_11434,N_11061);
or U12725 (N_12725,N_11829,N_11975);
or U12726 (N_12726,N_11373,N_11872);
and U12727 (N_12727,N_11418,N_11398);
xor U12728 (N_12728,N_11326,N_11877);
xnor U12729 (N_12729,N_11634,N_11322);
nor U12730 (N_12730,N_11169,N_11613);
or U12731 (N_12731,N_11417,N_11554);
and U12732 (N_12732,N_11934,N_11051);
nand U12733 (N_12733,N_11007,N_11808);
and U12734 (N_12734,N_11484,N_11085);
nor U12735 (N_12735,N_11904,N_11362);
and U12736 (N_12736,N_11008,N_11644);
nand U12737 (N_12737,N_11279,N_11511);
and U12738 (N_12738,N_11539,N_11595);
and U12739 (N_12739,N_11130,N_11700);
and U12740 (N_12740,N_11634,N_11794);
nor U12741 (N_12741,N_11493,N_11134);
and U12742 (N_12742,N_11874,N_11109);
nand U12743 (N_12743,N_11756,N_11723);
nand U12744 (N_12744,N_11611,N_11200);
and U12745 (N_12745,N_11178,N_11856);
nand U12746 (N_12746,N_11259,N_11819);
or U12747 (N_12747,N_11438,N_11968);
or U12748 (N_12748,N_11286,N_11859);
or U12749 (N_12749,N_11827,N_11681);
xor U12750 (N_12750,N_11298,N_11695);
and U12751 (N_12751,N_11336,N_11041);
nand U12752 (N_12752,N_11046,N_11167);
xor U12753 (N_12753,N_11898,N_11447);
and U12754 (N_12754,N_11894,N_11683);
xor U12755 (N_12755,N_11713,N_11017);
nand U12756 (N_12756,N_11977,N_11595);
nor U12757 (N_12757,N_11703,N_11706);
nand U12758 (N_12758,N_11556,N_11927);
and U12759 (N_12759,N_11162,N_11120);
nand U12760 (N_12760,N_11877,N_11615);
and U12761 (N_12761,N_11760,N_11320);
or U12762 (N_12762,N_11974,N_11571);
nand U12763 (N_12763,N_11132,N_11408);
xnor U12764 (N_12764,N_11434,N_11813);
or U12765 (N_12765,N_11265,N_11851);
xor U12766 (N_12766,N_11513,N_11499);
nor U12767 (N_12767,N_11105,N_11713);
or U12768 (N_12768,N_11226,N_11281);
and U12769 (N_12769,N_11518,N_11293);
nor U12770 (N_12770,N_11941,N_11085);
xnor U12771 (N_12771,N_11044,N_11403);
nor U12772 (N_12772,N_11345,N_11845);
and U12773 (N_12773,N_11902,N_11665);
xnor U12774 (N_12774,N_11918,N_11128);
nand U12775 (N_12775,N_11128,N_11161);
nand U12776 (N_12776,N_11436,N_11327);
or U12777 (N_12777,N_11145,N_11503);
nor U12778 (N_12778,N_11890,N_11124);
nand U12779 (N_12779,N_11061,N_11733);
nor U12780 (N_12780,N_11226,N_11921);
or U12781 (N_12781,N_11717,N_11608);
nor U12782 (N_12782,N_11083,N_11145);
and U12783 (N_12783,N_11022,N_11647);
or U12784 (N_12784,N_11981,N_11982);
or U12785 (N_12785,N_11040,N_11736);
nand U12786 (N_12786,N_11153,N_11606);
nand U12787 (N_12787,N_11951,N_11025);
and U12788 (N_12788,N_11244,N_11104);
nand U12789 (N_12789,N_11685,N_11494);
nor U12790 (N_12790,N_11727,N_11841);
or U12791 (N_12791,N_11201,N_11768);
and U12792 (N_12792,N_11878,N_11254);
nor U12793 (N_12793,N_11958,N_11124);
nand U12794 (N_12794,N_11401,N_11147);
nand U12795 (N_12795,N_11997,N_11266);
or U12796 (N_12796,N_11103,N_11414);
nor U12797 (N_12797,N_11602,N_11646);
xor U12798 (N_12798,N_11224,N_11932);
or U12799 (N_12799,N_11011,N_11809);
nor U12800 (N_12800,N_11610,N_11596);
or U12801 (N_12801,N_11096,N_11405);
nand U12802 (N_12802,N_11173,N_11790);
or U12803 (N_12803,N_11920,N_11346);
or U12804 (N_12804,N_11162,N_11389);
nand U12805 (N_12805,N_11403,N_11197);
and U12806 (N_12806,N_11272,N_11883);
or U12807 (N_12807,N_11182,N_11312);
or U12808 (N_12808,N_11986,N_11496);
xnor U12809 (N_12809,N_11661,N_11009);
and U12810 (N_12810,N_11430,N_11194);
or U12811 (N_12811,N_11455,N_11532);
nor U12812 (N_12812,N_11002,N_11657);
nor U12813 (N_12813,N_11068,N_11928);
nand U12814 (N_12814,N_11659,N_11215);
nand U12815 (N_12815,N_11206,N_11664);
xor U12816 (N_12816,N_11241,N_11679);
or U12817 (N_12817,N_11957,N_11327);
xnor U12818 (N_12818,N_11084,N_11851);
nand U12819 (N_12819,N_11390,N_11691);
nor U12820 (N_12820,N_11872,N_11414);
nor U12821 (N_12821,N_11692,N_11825);
or U12822 (N_12822,N_11661,N_11755);
nor U12823 (N_12823,N_11871,N_11365);
or U12824 (N_12824,N_11646,N_11731);
xor U12825 (N_12825,N_11494,N_11013);
xnor U12826 (N_12826,N_11246,N_11581);
and U12827 (N_12827,N_11083,N_11740);
nor U12828 (N_12828,N_11819,N_11181);
nand U12829 (N_12829,N_11819,N_11139);
xnor U12830 (N_12830,N_11954,N_11479);
xnor U12831 (N_12831,N_11159,N_11342);
nand U12832 (N_12832,N_11537,N_11028);
nor U12833 (N_12833,N_11147,N_11309);
nand U12834 (N_12834,N_11358,N_11273);
and U12835 (N_12835,N_11373,N_11612);
and U12836 (N_12836,N_11546,N_11681);
and U12837 (N_12837,N_11275,N_11048);
xnor U12838 (N_12838,N_11310,N_11437);
or U12839 (N_12839,N_11533,N_11739);
nor U12840 (N_12840,N_11380,N_11507);
or U12841 (N_12841,N_11224,N_11711);
and U12842 (N_12842,N_11774,N_11789);
nand U12843 (N_12843,N_11151,N_11749);
or U12844 (N_12844,N_11738,N_11594);
and U12845 (N_12845,N_11148,N_11884);
xor U12846 (N_12846,N_11820,N_11695);
and U12847 (N_12847,N_11787,N_11949);
nor U12848 (N_12848,N_11623,N_11034);
nand U12849 (N_12849,N_11178,N_11685);
xor U12850 (N_12850,N_11595,N_11772);
and U12851 (N_12851,N_11481,N_11807);
or U12852 (N_12852,N_11856,N_11854);
nor U12853 (N_12853,N_11633,N_11382);
nor U12854 (N_12854,N_11738,N_11812);
and U12855 (N_12855,N_11978,N_11732);
or U12856 (N_12856,N_11300,N_11131);
xor U12857 (N_12857,N_11066,N_11396);
xnor U12858 (N_12858,N_11188,N_11733);
and U12859 (N_12859,N_11855,N_11092);
xnor U12860 (N_12860,N_11783,N_11142);
nor U12861 (N_12861,N_11157,N_11807);
nor U12862 (N_12862,N_11934,N_11687);
and U12863 (N_12863,N_11841,N_11496);
nor U12864 (N_12864,N_11962,N_11615);
xnor U12865 (N_12865,N_11098,N_11955);
xnor U12866 (N_12866,N_11581,N_11949);
nand U12867 (N_12867,N_11394,N_11892);
or U12868 (N_12868,N_11894,N_11496);
and U12869 (N_12869,N_11803,N_11817);
nor U12870 (N_12870,N_11690,N_11050);
nor U12871 (N_12871,N_11235,N_11324);
nor U12872 (N_12872,N_11561,N_11903);
and U12873 (N_12873,N_11337,N_11137);
and U12874 (N_12874,N_11437,N_11988);
nor U12875 (N_12875,N_11961,N_11715);
nand U12876 (N_12876,N_11311,N_11221);
nor U12877 (N_12877,N_11937,N_11362);
nand U12878 (N_12878,N_11717,N_11269);
or U12879 (N_12879,N_11010,N_11124);
nor U12880 (N_12880,N_11760,N_11366);
xnor U12881 (N_12881,N_11949,N_11637);
nor U12882 (N_12882,N_11192,N_11009);
and U12883 (N_12883,N_11361,N_11160);
xor U12884 (N_12884,N_11545,N_11326);
and U12885 (N_12885,N_11161,N_11407);
and U12886 (N_12886,N_11374,N_11124);
nor U12887 (N_12887,N_11128,N_11179);
and U12888 (N_12888,N_11258,N_11988);
nand U12889 (N_12889,N_11026,N_11146);
or U12890 (N_12890,N_11863,N_11748);
or U12891 (N_12891,N_11423,N_11959);
or U12892 (N_12892,N_11735,N_11796);
or U12893 (N_12893,N_11450,N_11057);
nor U12894 (N_12894,N_11309,N_11646);
nand U12895 (N_12895,N_11145,N_11058);
nor U12896 (N_12896,N_11220,N_11244);
and U12897 (N_12897,N_11341,N_11024);
nand U12898 (N_12898,N_11398,N_11845);
or U12899 (N_12899,N_11314,N_11492);
nor U12900 (N_12900,N_11962,N_11608);
xor U12901 (N_12901,N_11167,N_11053);
and U12902 (N_12902,N_11334,N_11668);
or U12903 (N_12903,N_11686,N_11077);
nor U12904 (N_12904,N_11329,N_11835);
and U12905 (N_12905,N_11901,N_11290);
and U12906 (N_12906,N_11090,N_11428);
and U12907 (N_12907,N_11734,N_11135);
or U12908 (N_12908,N_11641,N_11394);
xnor U12909 (N_12909,N_11420,N_11045);
nand U12910 (N_12910,N_11353,N_11196);
or U12911 (N_12911,N_11435,N_11852);
nor U12912 (N_12912,N_11722,N_11114);
or U12913 (N_12913,N_11615,N_11729);
or U12914 (N_12914,N_11136,N_11067);
nor U12915 (N_12915,N_11072,N_11538);
xor U12916 (N_12916,N_11741,N_11351);
xor U12917 (N_12917,N_11962,N_11368);
nor U12918 (N_12918,N_11655,N_11404);
or U12919 (N_12919,N_11869,N_11573);
or U12920 (N_12920,N_11282,N_11631);
or U12921 (N_12921,N_11110,N_11552);
and U12922 (N_12922,N_11304,N_11858);
nand U12923 (N_12923,N_11844,N_11619);
or U12924 (N_12924,N_11363,N_11240);
nor U12925 (N_12925,N_11885,N_11486);
nand U12926 (N_12926,N_11740,N_11624);
xnor U12927 (N_12927,N_11352,N_11427);
nor U12928 (N_12928,N_11996,N_11464);
nand U12929 (N_12929,N_11824,N_11448);
nand U12930 (N_12930,N_11579,N_11782);
nand U12931 (N_12931,N_11887,N_11096);
and U12932 (N_12932,N_11758,N_11668);
nand U12933 (N_12933,N_11255,N_11895);
or U12934 (N_12934,N_11927,N_11191);
and U12935 (N_12935,N_11536,N_11570);
or U12936 (N_12936,N_11165,N_11449);
xor U12937 (N_12937,N_11696,N_11419);
nor U12938 (N_12938,N_11300,N_11051);
or U12939 (N_12939,N_11903,N_11859);
nor U12940 (N_12940,N_11157,N_11439);
or U12941 (N_12941,N_11260,N_11604);
or U12942 (N_12942,N_11553,N_11692);
and U12943 (N_12943,N_11864,N_11289);
and U12944 (N_12944,N_11133,N_11496);
nor U12945 (N_12945,N_11418,N_11586);
or U12946 (N_12946,N_11772,N_11332);
or U12947 (N_12947,N_11423,N_11347);
nand U12948 (N_12948,N_11858,N_11680);
nor U12949 (N_12949,N_11253,N_11616);
nor U12950 (N_12950,N_11633,N_11294);
and U12951 (N_12951,N_11893,N_11739);
xnor U12952 (N_12952,N_11696,N_11822);
and U12953 (N_12953,N_11992,N_11149);
nand U12954 (N_12954,N_11795,N_11024);
xnor U12955 (N_12955,N_11591,N_11091);
xor U12956 (N_12956,N_11239,N_11786);
nor U12957 (N_12957,N_11671,N_11628);
or U12958 (N_12958,N_11214,N_11893);
and U12959 (N_12959,N_11244,N_11016);
nand U12960 (N_12960,N_11321,N_11500);
nand U12961 (N_12961,N_11365,N_11958);
and U12962 (N_12962,N_11293,N_11231);
and U12963 (N_12963,N_11411,N_11220);
and U12964 (N_12964,N_11698,N_11117);
xor U12965 (N_12965,N_11970,N_11023);
xor U12966 (N_12966,N_11472,N_11044);
xnor U12967 (N_12967,N_11364,N_11719);
or U12968 (N_12968,N_11091,N_11086);
and U12969 (N_12969,N_11717,N_11204);
and U12970 (N_12970,N_11213,N_11778);
and U12971 (N_12971,N_11821,N_11538);
nor U12972 (N_12972,N_11838,N_11064);
and U12973 (N_12973,N_11069,N_11343);
and U12974 (N_12974,N_11251,N_11117);
nand U12975 (N_12975,N_11333,N_11980);
or U12976 (N_12976,N_11304,N_11395);
nor U12977 (N_12977,N_11808,N_11870);
nand U12978 (N_12978,N_11039,N_11809);
nor U12979 (N_12979,N_11592,N_11112);
nor U12980 (N_12980,N_11628,N_11997);
nor U12981 (N_12981,N_11925,N_11857);
nand U12982 (N_12982,N_11735,N_11835);
nor U12983 (N_12983,N_11106,N_11845);
nand U12984 (N_12984,N_11613,N_11700);
nor U12985 (N_12985,N_11521,N_11869);
nand U12986 (N_12986,N_11574,N_11954);
and U12987 (N_12987,N_11018,N_11042);
nand U12988 (N_12988,N_11187,N_11090);
xor U12989 (N_12989,N_11093,N_11997);
nand U12990 (N_12990,N_11964,N_11623);
nand U12991 (N_12991,N_11628,N_11741);
xor U12992 (N_12992,N_11247,N_11410);
and U12993 (N_12993,N_11284,N_11706);
and U12994 (N_12994,N_11891,N_11120);
nor U12995 (N_12995,N_11905,N_11823);
or U12996 (N_12996,N_11853,N_11177);
or U12997 (N_12997,N_11937,N_11777);
xnor U12998 (N_12998,N_11604,N_11846);
nand U12999 (N_12999,N_11352,N_11384);
or U13000 (N_13000,N_12318,N_12814);
xor U13001 (N_13001,N_12249,N_12323);
xor U13002 (N_13002,N_12012,N_12632);
or U13003 (N_13003,N_12830,N_12892);
nand U13004 (N_13004,N_12224,N_12669);
xnor U13005 (N_13005,N_12275,N_12435);
xnor U13006 (N_13006,N_12715,N_12545);
nand U13007 (N_13007,N_12358,N_12534);
nand U13008 (N_13008,N_12480,N_12753);
xor U13009 (N_13009,N_12344,N_12822);
or U13010 (N_13010,N_12646,N_12720);
and U13011 (N_13011,N_12512,N_12146);
or U13012 (N_13012,N_12272,N_12165);
nor U13013 (N_13013,N_12305,N_12621);
or U13014 (N_13014,N_12879,N_12543);
or U13015 (N_13015,N_12843,N_12353);
or U13016 (N_13016,N_12234,N_12216);
and U13017 (N_13017,N_12135,N_12619);
and U13018 (N_13018,N_12981,N_12985);
and U13019 (N_13019,N_12977,N_12885);
nor U13020 (N_13020,N_12335,N_12020);
nor U13021 (N_13021,N_12935,N_12766);
nor U13022 (N_13022,N_12898,N_12517);
nand U13023 (N_13023,N_12150,N_12682);
xnor U13024 (N_13024,N_12640,N_12235);
and U13025 (N_13025,N_12666,N_12732);
or U13026 (N_13026,N_12927,N_12837);
nor U13027 (N_13027,N_12198,N_12900);
xor U13028 (N_13028,N_12210,N_12613);
and U13029 (N_13029,N_12908,N_12933);
or U13030 (N_13030,N_12005,N_12507);
nor U13031 (N_13031,N_12737,N_12127);
xor U13032 (N_13032,N_12698,N_12696);
or U13033 (N_13033,N_12735,N_12411);
and U13034 (N_13034,N_12452,N_12761);
and U13035 (N_13035,N_12571,N_12492);
or U13036 (N_13036,N_12468,N_12805);
or U13037 (N_13037,N_12428,N_12767);
xnor U13038 (N_13038,N_12776,N_12228);
or U13039 (N_13039,N_12410,N_12462);
xnor U13040 (N_13040,N_12376,N_12844);
nand U13041 (N_13041,N_12333,N_12845);
nand U13042 (N_13042,N_12838,N_12481);
xnor U13043 (N_13043,N_12651,N_12848);
xor U13044 (N_13044,N_12929,N_12582);
and U13045 (N_13045,N_12361,N_12158);
and U13046 (N_13046,N_12606,N_12662);
nand U13047 (N_13047,N_12971,N_12099);
or U13048 (N_13048,N_12655,N_12577);
and U13049 (N_13049,N_12060,N_12231);
nor U13050 (N_13050,N_12192,N_12194);
nand U13051 (N_13051,N_12564,N_12710);
or U13052 (N_13052,N_12591,N_12009);
nor U13053 (N_13053,N_12775,N_12033);
and U13054 (N_13054,N_12920,N_12628);
xor U13055 (N_13055,N_12834,N_12040);
and U13056 (N_13056,N_12878,N_12405);
nor U13057 (N_13057,N_12043,N_12185);
xor U13058 (N_13058,N_12260,N_12679);
and U13059 (N_13059,N_12697,N_12759);
or U13060 (N_13060,N_12490,N_12291);
nor U13061 (N_13061,N_12093,N_12211);
nor U13062 (N_13062,N_12736,N_12849);
or U13063 (N_13063,N_12113,N_12245);
nor U13064 (N_13064,N_12811,N_12239);
nor U13065 (N_13065,N_12531,N_12392);
and U13066 (N_13066,N_12065,N_12128);
or U13067 (N_13067,N_12107,N_12401);
nor U13068 (N_13068,N_12382,N_12523);
xnor U13069 (N_13069,N_12626,N_12755);
xnor U13070 (N_13070,N_12731,N_12054);
nor U13071 (N_13071,N_12220,N_12835);
and U13072 (N_13072,N_12765,N_12876);
nand U13073 (N_13073,N_12899,N_12684);
and U13074 (N_13074,N_12456,N_12177);
or U13075 (N_13075,N_12675,N_12728);
and U13076 (N_13076,N_12576,N_12783);
or U13077 (N_13077,N_12637,N_12357);
and U13078 (N_13078,N_12151,N_12926);
xor U13079 (N_13079,N_12088,N_12082);
or U13080 (N_13080,N_12597,N_12790);
nor U13081 (N_13081,N_12037,N_12259);
xor U13082 (N_13082,N_12617,N_12573);
nand U13083 (N_13083,N_12520,N_12529);
or U13084 (N_13084,N_12180,N_12760);
xor U13085 (N_13085,N_12308,N_12421);
or U13086 (N_13086,N_12429,N_12251);
nor U13087 (N_13087,N_12189,N_12586);
nor U13088 (N_13088,N_12992,N_12544);
nand U13089 (N_13089,N_12290,N_12071);
or U13090 (N_13090,N_12021,N_12079);
or U13091 (N_13091,N_12562,N_12580);
or U13092 (N_13092,N_12351,N_12853);
xnor U13093 (N_13093,N_12579,N_12942);
xor U13094 (N_13094,N_12989,N_12585);
nor U13095 (N_13095,N_12890,N_12130);
and U13096 (N_13096,N_12129,N_12048);
or U13097 (N_13097,N_12945,N_12859);
nand U13098 (N_13098,N_12252,N_12758);
nand U13099 (N_13099,N_12340,N_12799);
or U13100 (N_13100,N_12553,N_12074);
and U13101 (N_13101,N_12886,N_12858);
nor U13102 (N_13102,N_12714,N_12727);
xor U13103 (N_13103,N_12800,N_12236);
and U13104 (N_13104,N_12739,N_12700);
nand U13105 (N_13105,N_12306,N_12982);
and U13106 (N_13106,N_12638,N_12824);
nor U13107 (N_13107,N_12796,N_12540);
nand U13108 (N_13108,N_12869,N_12689);
nand U13109 (N_13109,N_12903,N_12087);
and U13110 (N_13110,N_12653,N_12706);
nand U13111 (N_13111,N_12393,N_12491);
and U13112 (N_13112,N_12257,N_12705);
nor U13113 (N_13113,N_12371,N_12485);
xnor U13114 (N_13114,N_12536,N_12804);
nand U13115 (N_13115,N_12311,N_12167);
nor U13116 (N_13116,N_12524,N_12851);
or U13117 (N_13117,N_12703,N_12574);
nor U13118 (N_13118,N_12073,N_12538);
nand U13119 (N_13119,N_12961,N_12394);
xor U13120 (N_13120,N_12144,N_12503);
or U13121 (N_13121,N_12823,N_12865);
xor U13122 (N_13122,N_12059,N_12443);
or U13123 (N_13123,N_12064,N_12668);
and U13124 (N_13124,N_12449,N_12408);
nor U13125 (N_13125,N_12506,N_12042);
or U13126 (N_13126,N_12242,N_12687);
xor U13127 (N_13127,N_12115,N_12537);
and U13128 (N_13128,N_12578,N_12232);
nand U13129 (N_13129,N_12279,N_12554);
xor U13130 (N_13130,N_12195,N_12183);
nand U13131 (N_13131,N_12560,N_12988);
nor U13132 (N_13132,N_12077,N_12356);
xor U13133 (N_13133,N_12599,N_12609);
or U13134 (N_13134,N_12207,N_12522);
nor U13135 (N_13135,N_12779,N_12916);
or U13136 (N_13136,N_12169,N_12661);
nor U13137 (N_13137,N_12980,N_12432);
and U13138 (N_13138,N_12930,N_12999);
nand U13139 (N_13139,N_12950,N_12136);
nor U13140 (N_13140,N_12350,N_12894);
or U13141 (N_13141,N_12583,N_12409);
and U13142 (N_13142,N_12874,N_12388);
nor U13143 (N_13143,N_12566,N_12665);
nand U13144 (N_13144,N_12383,N_12826);
and U13145 (N_13145,N_12996,N_12200);
nor U13146 (N_13146,N_12702,N_12521);
nand U13147 (N_13147,N_12801,N_12178);
nand U13148 (N_13148,N_12026,N_12633);
or U13149 (N_13149,N_12749,N_12764);
nor U13150 (N_13150,N_12442,N_12162);
nand U13151 (N_13151,N_12484,N_12611);
and U13152 (N_13152,N_12444,N_12300);
nand U13153 (N_13153,N_12784,N_12918);
and U13154 (N_13154,N_12482,N_12891);
nand U13155 (N_13155,N_12078,N_12307);
and U13156 (N_13156,N_12086,N_12607);
nor U13157 (N_13157,N_12352,N_12096);
nor U13158 (N_13158,N_12140,N_12551);
nor U13159 (N_13159,N_12670,N_12047);
or U13160 (N_13160,N_12778,N_12615);
nand U13161 (N_13161,N_12230,N_12959);
xnor U13162 (N_13162,N_12893,N_12412);
nor U13163 (N_13163,N_12555,N_12172);
xor U13164 (N_13164,N_12139,N_12282);
or U13165 (N_13165,N_12802,N_12299);
nor U13166 (N_13166,N_12125,N_12631);
nor U13167 (N_13167,N_12550,N_12499);
nor U13168 (N_13168,N_12332,N_12363);
xnor U13169 (N_13169,N_12329,N_12664);
nor U13170 (N_13170,N_12769,N_12464);
nand U13171 (N_13171,N_12258,N_12004);
or U13172 (N_13172,N_12053,N_12692);
xor U13173 (N_13173,N_12287,N_12884);
or U13174 (N_13174,N_12241,N_12816);
xnor U13175 (N_13175,N_12827,N_12046);
nor U13176 (N_13176,N_12743,N_12747);
and U13177 (N_13177,N_12349,N_12247);
nor U13178 (N_13178,N_12474,N_12273);
nand U13179 (N_13179,N_12190,N_12062);
and U13180 (N_13180,N_12209,N_12000);
xor U13181 (N_13181,N_12268,N_12148);
or U13182 (N_13182,N_12075,N_12124);
or U13183 (N_13183,N_12833,N_12322);
or U13184 (N_13184,N_12288,N_12969);
or U13185 (N_13185,N_12437,N_12066);
or U13186 (N_13186,N_12440,N_12475);
and U13187 (N_13187,N_12445,N_12535);
and U13188 (N_13188,N_12106,N_12181);
nor U13189 (N_13189,N_12108,N_12016);
nor U13190 (N_13190,N_12419,N_12708);
and U13191 (N_13191,N_12203,N_12069);
nor U13192 (N_13192,N_12295,N_12153);
nand U13193 (N_13193,N_12725,N_12310);
xnor U13194 (N_13194,N_12023,N_12772);
nor U13195 (N_13195,N_12184,N_12339);
xor U13196 (N_13196,N_12673,N_12173);
and U13197 (N_13197,N_12379,N_12721);
nand U13198 (N_13198,N_12647,N_12425);
or U13199 (N_13199,N_12457,N_12154);
or U13200 (N_13200,N_12164,N_12212);
and U13201 (N_13201,N_12406,N_12463);
nand U13202 (N_13202,N_12501,N_12430);
nand U13203 (N_13203,N_12997,N_12119);
nand U13204 (N_13204,N_12187,N_12270);
and U13205 (N_13205,N_12722,N_12374);
and U13206 (N_13206,N_12623,N_12375);
and U13207 (N_13207,N_12365,N_12313);
or U13208 (N_13208,N_12603,N_12966);
nor U13209 (N_13209,N_12965,N_12547);
and U13210 (N_13210,N_12057,N_12386);
xor U13211 (N_13211,N_12568,N_12716);
xor U13212 (N_13212,N_12269,N_12711);
or U13213 (N_13213,N_12325,N_12174);
nor U13214 (N_13214,N_12598,N_12396);
and U13215 (N_13215,N_12789,N_12041);
or U13216 (N_13216,N_12176,N_12909);
or U13217 (N_13217,N_12745,N_12246);
nand U13218 (N_13218,N_12314,N_12122);
and U13219 (N_13219,N_12202,N_12347);
and U13220 (N_13220,N_12587,N_12559);
and U13221 (N_13221,N_12847,N_12451);
xor U13222 (N_13222,N_12785,N_12624);
xnor U13223 (N_13223,N_12302,N_12321);
nor U13224 (N_13224,N_12360,N_12159);
xnor U13225 (N_13225,N_12751,N_12389);
nor U13226 (N_13226,N_12362,N_12157);
or U13227 (N_13227,N_12941,N_12105);
or U13228 (N_13228,N_12565,N_12256);
and U13229 (N_13229,N_12188,N_12101);
or U13230 (N_13230,N_12511,N_12024);
nor U13231 (N_13231,N_12584,N_12953);
or U13232 (N_13232,N_12447,N_12552);
xnor U13233 (N_13233,N_12709,N_12143);
and U13234 (N_13234,N_12342,N_12690);
nor U13235 (N_13235,N_12348,N_12284);
and U13236 (N_13236,N_12793,N_12515);
nor U13237 (N_13237,N_12514,N_12880);
nand U13238 (N_13238,N_12791,N_12642);
or U13239 (N_13239,N_12262,N_12380);
xnor U13240 (N_13240,N_12455,N_12654);
and U13241 (N_13241,N_12635,N_12556);
nand U13242 (N_13242,N_12962,N_12116);
nand U13243 (N_13243,N_12656,N_12391);
or U13244 (N_13244,N_12919,N_12712);
or U13245 (N_13245,N_12671,N_12370);
or U13246 (N_13246,N_12987,N_12910);
or U13247 (N_13247,N_12806,N_12610);
or U13248 (N_13248,N_12494,N_12229);
nor U13249 (N_13249,N_12842,N_12533);
or U13250 (N_13250,N_12592,N_12897);
nor U13251 (N_13251,N_12952,N_12068);
or U13252 (N_13252,N_12864,N_12424);
or U13253 (N_13253,N_12384,N_12889);
nor U13254 (N_13254,N_12660,N_12770);
nand U13255 (N_13255,N_12820,N_12590);
or U13256 (N_13256,N_12530,N_12215);
and U13257 (N_13257,N_12001,N_12601);
nand U13258 (N_13258,N_12372,N_12469);
and U13259 (N_13259,N_12922,N_12439);
and U13260 (N_13260,N_12558,N_12338);
nor U13261 (N_13261,N_12142,N_12182);
nand U13262 (N_13262,N_12676,N_12780);
and U13263 (N_13263,N_12648,N_12828);
and U13264 (N_13264,N_12373,N_12984);
nand U13265 (N_13265,N_12070,N_12420);
or U13266 (N_13266,N_12588,N_12309);
nand U13267 (N_13267,N_12050,N_12354);
or U13268 (N_13268,N_12083,N_12652);
or U13269 (N_13269,N_12044,N_12875);
nor U13270 (N_13270,N_12002,N_12281);
nand U13271 (N_13271,N_12137,N_12787);
nor U13272 (N_13272,N_12657,N_12978);
nor U13273 (N_13273,N_12114,N_12602);
or U13274 (N_13274,N_12774,N_12508);
nor U13275 (N_13275,N_12301,N_12103);
or U13276 (N_13276,N_12525,N_12015);
nand U13277 (N_13277,N_12539,N_12091);
nor U13278 (N_13278,N_12902,N_12303);
or U13279 (N_13279,N_12931,N_12081);
or U13280 (N_13280,N_12199,N_12326);
nor U13281 (N_13281,N_12019,N_12809);
and U13282 (N_13282,N_12733,N_12126);
xnor U13283 (N_13283,N_12417,N_12912);
nand U13284 (N_13284,N_12090,N_12913);
nand U13285 (N_13285,N_12271,N_12250);
xor U13286 (N_13286,N_12297,N_12616);
nand U13287 (N_13287,N_12549,N_12111);
nor U13288 (N_13288,N_12713,N_12807);
or U13289 (N_13289,N_12404,N_12688);
or U13290 (N_13290,N_12862,N_12413);
xor U13291 (N_13291,N_12955,N_12487);
nand U13292 (N_13292,N_12681,N_12788);
nand U13293 (N_13293,N_12757,N_12120);
nor U13294 (N_13294,N_12527,N_12039);
nor U13295 (N_13295,N_12724,N_12940);
nand U13296 (N_13296,N_12943,N_12921);
xor U13297 (N_13297,N_12883,N_12958);
and U13298 (N_13298,N_12873,N_12014);
nand U13299 (N_13299,N_12888,N_12707);
xnor U13300 (N_13300,N_12841,N_12691);
nor U13301 (N_13301,N_12868,N_12097);
and U13302 (N_13302,N_12620,N_12699);
and U13303 (N_13303,N_12175,N_12528);
and U13304 (N_13304,N_12680,N_12771);
nand U13305 (N_13305,N_12505,N_12548);
and U13306 (N_13306,N_12650,N_12644);
and U13307 (N_13307,N_12949,N_12385);
and U13308 (N_13308,N_12109,N_12589);
nor U13309 (N_13309,N_12840,N_12618);
xnor U13310 (N_13310,N_12415,N_12836);
or U13311 (N_13311,N_12472,N_12267);
nor U13312 (N_13312,N_12990,N_12854);
nand U13313 (N_13313,N_12067,N_12346);
nand U13314 (N_13314,N_12240,N_12782);
and U13315 (N_13315,N_12399,N_12493);
and U13316 (N_13316,N_12817,N_12768);
nand U13317 (N_13317,N_12608,N_12718);
xor U13318 (N_13318,N_12133,N_12438);
or U13319 (N_13319,N_12867,N_12032);
xor U13320 (N_13320,N_12450,N_12911);
or U13321 (N_13321,N_12477,N_12035);
or U13322 (N_13322,N_12719,N_12238);
or U13323 (N_13323,N_12488,N_12092);
nor U13324 (N_13324,N_12798,N_12022);
and U13325 (N_13325,N_12740,N_12289);
and U13326 (N_13326,N_12118,N_12274);
xor U13327 (N_13327,N_12701,N_12968);
nand U13328 (N_13328,N_12331,N_12629);
nor U13329 (N_13329,N_12526,N_12055);
or U13330 (N_13330,N_12596,N_12294);
xnor U13331 (N_13331,N_12213,N_12423);
nand U13332 (N_13332,N_12860,N_12197);
nand U13333 (N_13333,N_12206,N_12237);
xnor U13334 (N_13334,N_12052,N_12896);
and U13335 (N_13335,N_12317,N_12089);
and U13336 (N_13336,N_12763,N_12003);
or U13337 (N_13337,N_12471,N_12147);
nor U13338 (N_13338,N_12663,N_12748);
and U13339 (N_13339,N_12027,N_12730);
xor U13340 (N_13340,N_12034,N_12928);
nor U13341 (N_13341,N_12557,N_12084);
xor U13342 (N_13342,N_12497,N_12466);
xnor U13343 (N_13343,N_12625,N_12217);
and U13344 (N_13344,N_12907,N_12255);
or U13345 (N_13345,N_12643,N_12476);
nand U13346 (N_13346,N_12575,N_12264);
or U13347 (N_13347,N_12341,N_12458);
or U13348 (N_13348,N_12917,N_12168);
xor U13349 (N_13349,N_12532,N_12937);
or U13350 (N_13350,N_12025,N_12744);
nand U13351 (N_13351,N_12193,N_12156);
or U13352 (N_13352,N_12446,N_12433);
or U13353 (N_13353,N_12479,N_12674);
nor U13354 (N_13354,N_12993,N_12612);
nor U13355 (N_13355,N_12460,N_12924);
or U13356 (N_13356,N_12914,N_12546);
or U13357 (N_13357,N_12773,N_12995);
xor U13358 (N_13358,N_12762,N_12972);
xnor U13359 (N_13359,N_12286,N_12881);
nand U13360 (N_13360,N_12387,N_12312);
nand U13361 (N_13361,N_12483,N_12658);
and U13362 (N_13362,N_12145,N_12453);
or U13363 (N_13363,N_12500,N_12756);
nor U13364 (N_13364,N_12645,N_12400);
nor U13365 (N_13365,N_12604,N_12542);
or U13366 (N_13366,N_12797,N_12316);
nor U13367 (N_13367,N_12418,N_12819);
or U13368 (N_13368,N_12416,N_12226);
xnor U13369 (N_13369,N_12201,N_12832);
nand U13370 (N_13370,N_12998,N_12395);
nand U13371 (N_13371,N_12112,N_12364);
nor U13372 (N_13372,N_12277,N_12976);
and U13373 (N_13373,N_12243,N_12498);
nand U13374 (N_13374,N_12011,N_12882);
nand U13375 (N_13375,N_12677,N_12315);
xnor U13376 (N_13376,N_12149,N_12355);
or U13377 (N_13377,N_12777,N_12948);
and U13378 (N_13378,N_12161,N_12821);
nor U13379 (N_13379,N_12298,N_12963);
nor U13380 (N_13380,N_12334,N_12141);
nand U13381 (N_13381,N_12327,N_12857);
xnor U13382 (N_13382,N_12695,N_12138);
and U13383 (N_13383,N_12939,N_12979);
xnor U13384 (N_13384,N_12672,N_12856);
nand U13385 (N_13385,N_12152,N_12072);
and U13386 (N_13386,N_12085,N_12678);
xnor U13387 (N_13387,N_12098,N_12818);
or U13388 (N_13388,N_12872,N_12381);
nand U13389 (N_13389,N_12754,N_12947);
or U13390 (N_13390,N_12486,N_12956);
and U13391 (N_13391,N_12983,N_12752);
nor U13392 (N_13392,N_12904,N_12970);
nand U13393 (N_13393,N_12171,N_12434);
xor U13394 (N_13394,N_12467,N_12038);
nand U13395 (N_13395,N_12516,N_12634);
xnor U13396 (N_13396,N_12008,N_12593);
or U13397 (N_13397,N_12649,N_12366);
xor U13398 (N_13398,N_12328,N_12470);
and U13399 (N_13399,N_12863,N_12541);
xnor U13400 (N_13400,N_12831,N_12726);
nor U13401 (N_13401,N_12923,N_12495);
and U13402 (N_13402,N_12991,N_12954);
xor U13403 (N_13403,N_12368,N_12685);
and U13404 (N_13404,N_12510,N_12861);
or U13405 (N_13405,N_12223,N_12013);
nor U13406 (N_13406,N_12123,N_12441);
nor U13407 (N_13407,N_12627,N_12131);
xor U13408 (N_13408,N_12825,N_12402);
nand U13409 (N_13409,N_12102,N_12887);
xor U13410 (N_13410,N_12426,N_12723);
and U13411 (N_13411,N_12283,N_12398);
nand U13412 (N_13412,N_12397,N_12227);
nor U13413 (N_13413,N_12938,N_12320);
nor U13414 (N_13414,N_12519,N_12218);
nand U13415 (N_13415,N_12160,N_12855);
or U13416 (N_13416,N_12006,N_12454);
nand U13417 (N_13417,N_12812,N_12063);
nand U13418 (N_13418,N_12792,N_12292);
and U13419 (N_13419,N_12594,N_12436);
nor U13420 (N_13420,N_12569,N_12278);
or U13421 (N_13421,N_12786,N_12390);
nand U13422 (N_13422,N_12489,N_12076);
xor U13423 (N_13423,N_12986,N_12906);
or U13424 (N_13424,N_12427,N_12049);
xor U13425 (N_13425,N_12581,N_12028);
xor U13426 (N_13426,N_12870,N_12448);
nor U13427 (N_13427,N_12877,N_12803);
nand U13428 (N_13428,N_12422,N_12905);
and U13429 (N_13429,N_12254,N_12957);
nor U13430 (N_13430,N_12901,N_12850);
or U13431 (N_13431,N_12829,N_12694);
or U13432 (N_13432,N_12017,N_12058);
nand U13433 (N_13433,N_12946,N_12407);
nor U13434 (N_13434,N_12994,N_12866);
xor U13435 (N_13435,N_12007,N_12852);
or U13436 (N_13436,N_12936,N_12742);
or U13437 (N_13437,N_12324,N_12051);
xnor U13438 (N_13438,N_12595,N_12461);
and U13439 (N_13439,N_12191,N_12170);
nor U13440 (N_13440,N_12233,N_12561);
nor U13441 (N_13441,N_12693,N_12513);
nor U13442 (N_13442,N_12163,N_12974);
nor U13443 (N_13443,N_12605,N_12359);
and U13444 (N_13444,N_12659,N_12925);
or U13445 (N_13445,N_12166,N_12155);
nand U13446 (N_13446,N_12330,N_12600);
and U13447 (N_13447,N_12337,N_12345);
or U13448 (N_13448,N_12186,N_12686);
and U13449 (N_13449,N_12496,N_12895);
nand U13450 (N_13450,N_12117,N_12095);
nor U13451 (N_13451,N_12932,N_12871);
nand U13452 (N_13452,N_12196,N_12810);
nand U13453 (N_13453,N_12639,N_12934);
nor U13454 (N_13454,N_12738,N_12944);
xnor U13455 (N_13455,N_12222,N_12964);
xor U13456 (N_13456,N_12293,N_12622);
nor U13457 (N_13457,N_12304,N_12518);
nand U13458 (N_13458,N_12502,N_12795);
and U13459 (N_13459,N_12459,N_12263);
nor U13460 (N_13460,N_12431,N_12614);
and U13461 (N_13461,N_12967,N_12951);
xnor U13462 (N_13462,N_12570,N_12846);
nor U13463 (N_13463,N_12815,N_12975);
nand U13464 (N_13464,N_12336,N_12734);
nor U13465 (N_13465,N_12030,N_12478);
xnor U13466 (N_13466,N_12036,N_12369);
or U13467 (N_13467,N_12121,N_12473);
xor U13468 (N_13468,N_12319,N_12221);
and U13469 (N_13469,N_12741,N_12973);
xnor U13470 (N_13470,N_12225,N_12403);
and U13471 (N_13471,N_12031,N_12261);
nand U13472 (N_13472,N_12029,N_12641);
or U13473 (N_13473,N_12414,N_12377);
and U13474 (N_13474,N_12205,N_12367);
xor U13475 (N_13475,N_12214,N_12100);
nor U13476 (N_13476,N_12572,N_12960);
nor U13477 (N_13477,N_12094,N_12808);
nor U13478 (N_13478,N_12630,N_12567);
or U13479 (N_13479,N_12276,N_12509);
nor U13480 (N_13480,N_12794,N_12285);
and U13481 (N_13481,N_12704,N_12104);
xnor U13482 (N_13482,N_12378,N_12056);
nand U13483 (N_13483,N_12266,N_12729);
and U13484 (N_13484,N_12265,N_12683);
nand U13485 (N_13485,N_12504,N_12717);
or U13486 (N_13486,N_12253,N_12839);
and U13487 (N_13487,N_12110,N_12248);
nand U13488 (N_13488,N_12244,N_12563);
and U13489 (N_13489,N_12915,N_12204);
nor U13490 (N_13490,N_12781,N_12018);
xor U13491 (N_13491,N_12010,N_12208);
nor U13492 (N_13492,N_12132,N_12296);
nor U13493 (N_13493,N_12061,N_12219);
and U13494 (N_13494,N_12667,N_12080);
nand U13495 (N_13495,N_12746,N_12045);
xnor U13496 (N_13496,N_12134,N_12636);
xor U13497 (N_13497,N_12343,N_12813);
and U13498 (N_13498,N_12280,N_12465);
or U13499 (N_13499,N_12750,N_12179);
nand U13500 (N_13500,N_12205,N_12161);
nor U13501 (N_13501,N_12858,N_12752);
xor U13502 (N_13502,N_12675,N_12983);
nor U13503 (N_13503,N_12198,N_12843);
xnor U13504 (N_13504,N_12385,N_12581);
nand U13505 (N_13505,N_12796,N_12315);
nor U13506 (N_13506,N_12735,N_12342);
nand U13507 (N_13507,N_12813,N_12973);
xnor U13508 (N_13508,N_12969,N_12203);
nand U13509 (N_13509,N_12144,N_12690);
or U13510 (N_13510,N_12692,N_12543);
nand U13511 (N_13511,N_12350,N_12034);
nand U13512 (N_13512,N_12320,N_12436);
or U13513 (N_13513,N_12145,N_12929);
or U13514 (N_13514,N_12491,N_12888);
or U13515 (N_13515,N_12253,N_12403);
nor U13516 (N_13516,N_12518,N_12253);
nor U13517 (N_13517,N_12814,N_12137);
xnor U13518 (N_13518,N_12821,N_12741);
and U13519 (N_13519,N_12824,N_12988);
or U13520 (N_13520,N_12429,N_12602);
nand U13521 (N_13521,N_12283,N_12785);
nor U13522 (N_13522,N_12770,N_12878);
xnor U13523 (N_13523,N_12997,N_12804);
and U13524 (N_13524,N_12553,N_12676);
and U13525 (N_13525,N_12210,N_12498);
or U13526 (N_13526,N_12276,N_12988);
xor U13527 (N_13527,N_12957,N_12240);
or U13528 (N_13528,N_12202,N_12588);
and U13529 (N_13529,N_12914,N_12852);
or U13530 (N_13530,N_12101,N_12360);
or U13531 (N_13531,N_12179,N_12784);
nor U13532 (N_13532,N_12186,N_12890);
nor U13533 (N_13533,N_12995,N_12186);
xnor U13534 (N_13534,N_12356,N_12094);
and U13535 (N_13535,N_12593,N_12030);
and U13536 (N_13536,N_12933,N_12911);
or U13537 (N_13537,N_12168,N_12973);
or U13538 (N_13538,N_12412,N_12620);
nor U13539 (N_13539,N_12551,N_12682);
and U13540 (N_13540,N_12339,N_12507);
and U13541 (N_13541,N_12336,N_12826);
xnor U13542 (N_13542,N_12154,N_12970);
nor U13543 (N_13543,N_12864,N_12904);
and U13544 (N_13544,N_12623,N_12941);
and U13545 (N_13545,N_12455,N_12555);
xor U13546 (N_13546,N_12774,N_12016);
nand U13547 (N_13547,N_12210,N_12983);
nor U13548 (N_13548,N_12136,N_12174);
and U13549 (N_13549,N_12876,N_12286);
or U13550 (N_13550,N_12602,N_12853);
and U13551 (N_13551,N_12051,N_12349);
xor U13552 (N_13552,N_12873,N_12118);
and U13553 (N_13553,N_12706,N_12450);
xor U13554 (N_13554,N_12507,N_12412);
and U13555 (N_13555,N_12157,N_12550);
nand U13556 (N_13556,N_12857,N_12256);
xor U13557 (N_13557,N_12862,N_12264);
nor U13558 (N_13558,N_12343,N_12198);
nand U13559 (N_13559,N_12062,N_12993);
nor U13560 (N_13560,N_12192,N_12068);
and U13561 (N_13561,N_12983,N_12915);
and U13562 (N_13562,N_12358,N_12149);
nand U13563 (N_13563,N_12881,N_12631);
or U13564 (N_13564,N_12663,N_12297);
xnor U13565 (N_13565,N_12543,N_12290);
nor U13566 (N_13566,N_12686,N_12416);
nor U13567 (N_13567,N_12021,N_12885);
nor U13568 (N_13568,N_12297,N_12314);
nand U13569 (N_13569,N_12137,N_12711);
xor U13570 (N_13570,N_12596,N_12556);
xor U13571 (N_13571,N_12971,N_12687);
nand U13572 (N_13572,N_12217,N_12846);
xor U13573 (N_13573,N_12437,N_12717);
or U13574 (N_13574,N_12690,N_12638);
or U13575 (N_13575,N_12354,N_12178);
or U13576 (N_13576,N_12405,N_12330);
and U13577 (N_13577,N_12913,N_12534);
or U13578 (N_13578,N_12124,N_12581);
nor U13579 (N_13579,N_12374,N_12523);
nor U13580 (N_13580,N_12577,N_12762);
xnor U13581 (N_13581,N_12243,N_12947);
or U13582 (N_13582,N_12765,N_12034);
nor U13583 (N_13583,N_12715,N_12728);
and U13584 (N_13584,N_12265,N_12307);
xnor U13585 (N_13585,N_12618,N_12962);
and U13586 (N_13586,N_12375,N_12185);
xnor U13587 (N_13587,N_12771,N_12409);
nand U13588 (N_13588,N_12134,N_12852);
nor U13589 (N_13589,N_12956,N_12851);
or U13590 (N_13590,N_12161,N_12875);
and U13591 (N_13591,N_12105,N_12816);
xnor U13592 (N_13592,N_12978,N_12385);
or U13593 (N_13593,N_12306,N_12223);
nor U13594 (N_13594,N_12282,N_12833);
nand U13595 (N_13595,N_12558,N_12291);
and U13596 (N_13596,N_12139,N_12359);
nor U13597 (N_13597,N_12257,N_12557);
or U13598 (N_13598,N_12498,N_12078);
and U13599 (N_13599,N_12868,N_12674);
xor U13600 (N_13600,N_12541,N_12276);
or U13601 (N_13601,N_12439,N_12257);
and U13602 (N_13602,N_12565,N_12209);
nand U13603 (N_13603,N_12925,N_12924);
nor U13604 (N_13604,N_12408,N_12542);
and U13605 (N_13605,N_12149,N_12627);
nand U13606 (N_13606,N_12893,N_12796);
xnor U13607 (N_13607,N_12963,N_12842);
or U13608 (N_13608,N_12178,N_12415);
or U13609 (N_13609,N_12131,N_12306);
nor U13610 (N_13610,N_12875,N_12634);
nor U13611 (N_13611,N_12242,N_12020);
xnor U13612 (N_13612,N_12212,N_12789);
nand U13613 (N_13613,N_12757,N_12012);
nor U13614 (N_13614,N_12714,N_12938);
or U13615 (N_13615,N_12264,N_12607);
and U13616 (N_13616,N_12888,N_12815);
xnor U13617 (N_13617,N_12555,N_12049);
and U13618 (N_13618,N_12960,N_12910);
nand U13619 (N_13619,N_12616,N_12261);
xor U13620 (N_13620,N_12612,N_12647);
or U13621 (N_13621,N_12395,N_12209);
nand U13622 (N_13622,N_12494,N_12187);
nor U13623 (N_13623,N_12509,N_12144);
nor U13624 (N_13624,N_12006,N_12869);
xor U13625 (N_13625,N_12553,N_12080);
and U13626 (N_13626,N_12340,N_12636);
and U13627 (N_13627,N_12727,N_12451);
and U13628 (N_13628,N_12471,N_12805);
and U13629 (N_13629,N_12610,N_12341);
nand U13630 (N_13630,N_12572,N_12493);
nand U13631 (N_13631,N_12186,N_12899);
nor U13632 (N_13632,N_12968,N_12867);
or U13633 (N_13633,N_12249,N_12451);
and U13634 (N_13634,N_12029,N_12729);
nand U13635 (N_13635,N_12199,N_12950);
and U13636 (N_13636,N_12967,N_12580);
xor U13637 (N_13637,N_12095,N_12301);
xor U13638 (N_13638,N_12574,N_12636);
nor U13639 (N_13639,N_12173,N_12042);
or U13640 (N_13640,N_12775,N_12350);
xnor U13641 (N_13641,N_12280,N_12715);
xor U13642 (N_13642,N_12893,N_12142);
or U13643 (N_13643,N_12416,N_12575);
or U13644 (N_13644,N_12208,N_12980);
nor U13645 (N_13645,N_12764,N_12306);
xnor U13646 (N_13646,N_12165,N_12781);
xor U13647 (N_13647,N_12981,N_12320);
or U13648 (N_13648,N_12208,N_12375);
and U13649 (N_13649,N_12837,N_12615);
nor U13650 (N_13650,N_12132,N_12521);
or U13651 (N_13651,N_12413,N_12755);
and U13652 (N_13652,N_12333,N_12436);
xor U13653 (N_13653,N_12760,N_12590);
xnor U13654 (N_13654,N_12522,N_12789);
or U13655 (N_13655,N_12908,N_12593);
and U13656 (N_13656,N_12804,N_12660);
nand U13657 (N_13657,N_12251,N_12498);
nand U13658 (N_13658,N_12078,N_12643);
and U13659 (N_13659,N_12272,N_12911);
and U13660 (N_13660,N_12135,N_12545);
nand U13661 (N_13661,N_12776,N_12242);
nand U13662 (N_13662,N_12784,N_12140);
nor U13663 (N_13663,N_12035,N_12890);
and U13664 (N_13664,N_12634,N_12713);
nand U13665 (N_13665,N_12826,N_12959);
xor U13666 (N_13666,N_12399,N_12476);
and U13667 (N_13667,N_12253,N_12576);
or U13668 (N_13668,N_12516,N_12354);
nand U13669 (N_13669,N_12238,N_12524);
xnor U13670 (N_13670,N_12694,N_12387);
and U13671 (N_13671,N_12299,N_12108);
nand U13672 (N_13672,N_12910,N_12804);
and U13673 (N_13673,N_12408,N_12527);
xnor U13674 (N_13674,N_12321,N_12076);
or U13675 (N_13675,N_12302,N_12370);
xor U13676 (N_13676,N_12033,N_12343);
nor U13677 (N_13677,N_12526,N_12890);
xnor U13678 (N_13678,N_12126,N_12953);
or U13679 (N_13679,N_12406,N_12807);
and U13680 (N_13680,N_12356,N_12248);
and U13681 (N_13681,N_12376,N_12972);
and U13682 (N_13682,N_12339,N_12657);
xor U13683 (N_13683,N_12669,N_12495);
and U13684 (N_13684,N_12144,N_12036);
and U13685 (N_13685,N_12208,N_12215);
xor U13686 (N_13686,N_12215,N_12806);
or U13687 (N_13687,N_12875,N_12246);
nand U13688 (N_13688,N_12168,N_12928);
and U13689 (N_13689,N_12618,N_12531);
nor U13690 (N_13690,N_12251,N_12163);
nand U13691 (N_13691,N_12725,N_12054);
xor U13692 (N_13692,N_12088,N_12253);
nor U13693 (N_13693,N_12791,N_12052);
and U13694 (N_13694,N_12241,N_12741);
and U13695 (N_13695,N_12405,N_12781);
nand U13696 (N_13696,N_12919,N_12434);
nand U13697 (N_13697,N_12786,N_12214);
or U13698 (N_13698,N_12305,N_12126);
and U13699 (N_13699,N_12130,N_12372);
nor U13700 (N_13700,N_12141,N_12609);
xor U13701 (N_13701,N_12880,N_12990);
or U13702 (N_13702,N_12321,N_12816);
xnor U13703 (N_13703,N_12621,N_12201);
nor U13704 (N_13704,N_12425,N_12002);
xor U13705 (N_13705,N_12512,N_12038);
nor U13706 (N_13706,N_12026,N_12319);
and U13707 (N_13707,N_12259,N_12709);
nor U13708 (N_13708,N_12513,N_12158);
nor U13709 (N_13709,N_12494,N_12420);
xor U13710 (N_13710,N_12843,N_12075);
nor U13711 (N_13711,N_12783,N_12836);
nand U13712 (N_13712,N_12792,N_12753);
nand U13713 (N_13713,N_12048,N_12403);
xnor U13714 (N_13714,N_12535,N_12673);
xnor U13715 (N_13715,N_12129,N_12850);
or U13716 (N_13716,N_12024,N_12174);
or U13717 (N_13717,N_12042,N_12655);
nor U13718 (N_13718,N_12720,N_12874);
nand U13719 (N_13719,N_12624,N_12144);
nor U13720 (N_13720,N_12535,N_12090);
nor U13721 (N_13721,N_12994,N_12244);
nand U13722 (N_13722,N_12513,N_12195);
and U13723 (N_13723,N_12574,N_12685);
xor U13724 (N_13724,N_12820,N_12460);
nand U13725 (N_13725,N_12552,N_12208);
nor U13726 (N_13726,N_12393,N_12817);
or U13727 (N_13727,N_12427,N_12161);
or U13728 (N_13728,N_12309,N_12998);
or U13729 (N_13729,N_12918,N_12143);
xnor U13730 (N_13730,N_12612,N_12867);
xor U13731 (N_13731,N_12064,N_12961);
nor U13732 (N_13732,N_12584,N_12599);
nand U13733 (N_13733,N_12956,N_12424);
or U13734 (N_13734,N_12431,N_12343);
nor U13735 (N_13735,N_12497,N_12070);
and U13736 (N_13736,N_12714,N_12944);
or U13737 (N_13737,N_12710,N_12861);
and U13738 (N_13738,N_12800,N_12842);
or U13739 (N_13739,N_12022,N_12792);
and U13740 (N_13740,N_12790,N_12487);
or U13741 (N_13741,N_12756,N_12929);
nor U13742 (N_13742,N_12485,N_12610);
xor U13743 (N_13743,N_12601,N_12228);
nand U13744 (N_13744,N_12329,N_12216);
xnor U13745 (N_13745,N_12445,N_12388);
or U13746 (N_13746,N_12185,N_12755);
and U13747 (N_13747,N_12376,N_12377);
nand U13748 (N_13748,N_12667,N_12448);
xnor U13749 (N_13749,N_12380,N_12916);
or U13750 (N_13750,N_12904,N_12695);
or U13751 (N_13751,N_12387,N_12440);
nor U13752 (N_13752,N_12575,N_12518);
xor U13753 (N_13753,N_12105,N_12154);
nand U13754 (N_13754,N_12700,N_12295);
nor U13755 (N_13755,N_12298,N_12384);
nand U13756 (N_13756,N_12167,N_12248);
nand U13757 (N_13757,N_12634,N_12484);
nand U13758 (N_13758,N_12786,N_12067);
xor U13759 (N_13759,N_12459,N_12604);
nor U13760 (N_13760,N_12049,N_12272);
and U13761 (N_13761,N_12358,N_12708);
nor U13762 (N_13762,N_12763,N_12966);
nand U13763 (N_13763,N_12121,N_12214);
nand U13764 (N_13764,N_12857,N_12988);
and U13765 (N_13765,N_12912,N_12739);
xnor U13766 (N_13766,N_12743,N_12511);
nand U13767 (N_13767,N_12869,N_12254);
and U13768 (N_13768,N_12480,N_12025);
nor U13769 (N_13769,N_12451,N_12546);
and U13770 (N_13770,N_12368,N_12177);
xnor U13771 (N_13771,N_12488,N_12474);
nor U13772 (N_13772,N_12749,N_12541);
nand U13773 (N_13773,N_12045,N_12651);
or U13774 (N_13774,N_12270,N_12712);
xor U13775 (N_13775,N_12889,N_12307);
nand U13776 (N_13776,N_12175,N_12694);
or U13777 (N_13777,N_12154,N_12869);
xnor U13778 (N_13778,N_12297,N_12486);
and U13779 (N_13779,N_12564,N_12745);
xnor U13780 (N_13780,N_12907,N_12804);
xor U13781 (N_13781,N_12658,N_12536);
and U13782 (N_13782,N_12323,N_12742);
nor U13783 (N_13783,N_12835,N_12842);
nor U13784 (N_13784,N_12670,N_12024);
or U13785 (N_13785,N_12067,N_12039);
nand U13786 (N_13786,N_12021,N_12121);
nor U13787 (N_13787,N_12547,N_12275);
or U13788 (N_13788,N_12196,N_12765);
or U13789 (N_13789,N_12900,N_12724);
and U13790 (N_13790,N_12713,N_12044);
nor U13791 (N_13791,N_12447,N_12303);
xnor U13792 (N_13792,N_12184,N_12481);
nor U13793 (N_13793,N_12083,N_12191);
xor U13794 (N_13794,N_12710,N_12264);
nand U13795 (N_13795,N_12376,N_12762);
nand U13796 (N_13796,N_12718,N_12502);
nor U13797 (N_13797,N_12432,N_12841);
or U13798 (N_13798,N_12298,N_12911);
or U13799 (N_13799,N_12590,N_12449);
nor U13800 (N_13800,N_12245,N_12477);
nand U13801 (N_13801,N_12501,N_12782);
nand U13802 (N_13802,N_12079,N_12127);
and U13803 (N_13803,N_12237,N_12004);
or U13804 (N_13804,N_12309,N_12423);
or U13805 (N_13805,N_12115,N_12880);
nor U13806 (N_13806,N_12836,N_12149);
and U13807 (N_13807,N_12577,N_12423);
and U13808 (N_13808,N_12819,N_12594);
and U13809 (N_13809,N_12491,N_12187);
or U13810 (N_13810,N_12946,N_12982);
and U13811 (N_13811,N_12915,N_12533);
nand U13812 (N_13812,N_12319,N_12822);
xor U13813 (N_13813,N_12183,N_12876);
nor U13814 (N_13814,N_12915,N_12901);
nor U13815 (N_13815,N_12680,N_12187);
nand U13816 (N_13816,N_12789,N_12376);
xor U13817 (N_13817,N_12879,N_12650);
nor U13818 (N_13818,N_12981,N_12710);
or U13819 (N_13819,N_12445,N_12711);
xnor U13820 (N_13820,N_12633,N_12210);
nor U13821 (N_13821,N_12320,N_12570);
and U13822 (N_13822,N_12710,N_12326);
or U13823 (N_13823,N_12094,N_12001);
and U13824 (N_13824,N_12968,N_12190);
nor U13825 (N_13825,N_12828,N_12001);
nand U13826 (N_13826,N_12413,N_12144);
or U13827 (N_13827,N_12273,N_12389);
xor U13828 (N_13828,N_12646,N_12972);
and U13829 (N_13829,N_12569,N_12520);
nand U13830 (N_13830,N_12282,N_12349);
or U13831 (N_13831,N_12485,N_12880);
nor U13832 (N_13832,N_12183,N_12076);
or U13833 (N_13833,N_12784,N_12947);
or U13834 (N_13834,N_12708,N_12717);
or U13835 (N_13835,N_12285,N_12511);
or U13836 (N_13836,N_12532,N_12141);
or U13837 (N_13837,N_12846,N_12295);
nor U13838 (N_13838,N_12499,N_12891);
and U13839 (N_13839,N_12122,N_12179);
or U13840 (N_13840,N_12619,N_12202);
or U13841 (N_13841,N_12065,N_12049);
and U13842 (N_13842,N_12820,N_12322);
nor U13843 (N_13843,N_12261,N_12305);
or U13844 (N_13844,N_12002,N_12649);
nand U13845 (N_13845,N_12883,N_12879);
nor U13846 (N_13846,N_12777,N_12305);
xnor U13847 (N_13847,N_12349,N_12159);
nand U13848 (N_13848,N_12163,N_12171);
nand U13849 (N_13849,N_12750,N_12424);
nor U13850 (N_13850,N_12338,N_12879);
and U13851 (N_13851,N_12277,N_12238);
nand U13852 (N_13852,N_12439,N_12820);
xnor U13853 (N_13853,N_12577,N_12476);
and U13854 (N_13854,N_12756,N_12921);
or U13855 (N_13855,N_12175,N_12283);
xor U13856 (N_13856,N_12035,N_12160);
and U13857 (N_13857,N_12240,N_12146);
or U13858 (N_13858,N_12308,N_12800);
nand U13859 (N_13859,N_12923,N_12991);
xnor U13860 (N_13860,N_12548,N_12442);
nor U13861 (N_13861,N_12048,N_12345);
nand U13862 (N_13862,N_12538,N_12215);
nand U13863 (N_13863,N_12829,N_12126);
nor U13864 (N_13864,N_12180,N_12999);
nor U13865 (N_13865,N_12557,N_12337);
nand U13866 (N_13866,N_12291,N_12629);
xnor U13867 (N_13867,N_12766,N_12001);
xor U13868 (N_13868,N_12517,N_12416);
or U13869 (N_13869,N_12221,N_12236);
nor U13870 (N_13870,N_12612,N_12753);
nand U13871 (N_13871,N_12331,N_12507);
or U13872 (N_13872,N_12702,N_12309);
xor U13873 (N_13873,N_12615,N_12456);
and U13874 (N_13874,N_12554,N_12692);
nor U13875 (N_13875,N_12048,N_12280);
xor U13876 (N_13876,N_12360,N_12434);
xnor U13877 (N_13877,N_12073,N_12572);
xnor U13878 (N_13878,N_12822,N_12434);
xor U13879 (N_13879,N_12615,N_12177);
and U13880 (N_13880,N_12871,N_12984);
or U13881 (N_13881,N_12820,N_12112);
xor U13882 (N_13882,N_12736,N_12535);
xor U13883 (N_13883,N_12432,N_12701);
xor U13884 (N_13884,N_12841,N_12317);
or U13885 (N_13885,N_12810,N_12681);
nor U13886 (N_13886,N_12876,N_12190);
nor U13887 (N_13887,N_12734,N_12092);
and U13888 (N_13888,N_12262,N_12019);
and U13889 (N_13889,N_12559,N_12910);
and U13890 (N_13890,N_12768,N_12590);
nor U13891 (N_13891,N_12665,N_12629);
xor U13892 (N_13892,N_12564,N_12773);
nor U13893 (N_13893,N_12935,N_12471);
or U13894 (N_13894,N_12337,N_12370);
nor U13895 (N_13895,N_12660,N_12323);
or U13896 (N_13896,N_12301,N_12583);
nor U13897 (N_13897,N_12821,N_12456);
nor U13898 (N_13898,N_12111,N_12346);
nor U13899 (N_13899,N_12503,N_12614);
and U13900 (N_13900,N_12912,N_12623);
nand U13901 (N_13901,N_12414,N_12184);
and U13902 (N_13902,N_12218,N_12610);
nand U13903 (N_13903,N_12880,N_12747);
xor U13904 (N_13904,N_12350,N_12351);
xnor U13905 (N_13905,N_12833,N_12831);
nor U13906 (N_13906,N_12115,N_12328);
nand U13907 (N_13907,N_12001,N_12501);
nor U13908 (N_13908,N_12847,N_12347);
xor U13909 (N_13909,N_12536,N_12057);
nor U13910 (N_13910,N_12586,N_12485);
xnor U13911 (N_13911,N_12634,N_12105);
xor U13912 (N_13912,N_12397,N_12514);
xnor U13913 (N_13913,N_12690,N_12930);
xnor U13914 (N_13914,N_12953,N_12622);
or U13915 (N_13915,N_12081,N_12924);
or U13916 (N_13916,N_12483,N_12942);
or U13917 (N_13917,N_12365,N_12674);
xnor U13918 (N_13918,N_12217,N_12148);
xnor U13919 (N_13919,N_12381,N_12424);
xnor U13920 (N_13920,N_12799,N_12183);
or U13921 (N_13921,N_12455,N_12852);
nor U13922 (N_13922,N_12895,N_12211);
nand U13923 (N_13923,N_12509,N_12006);
xor U13924 (N_13924,N_12348,N_12913);
or U13925 (N_13925,N_12153,N_12743);
nand U13926 (N_13926,N_12477,N_12868);
or U13927 (N_13927,N_12762,N_12880);
nor U13928 (N_13928,N_12453,N_12408);
and U13929 (N_13929,N_12822,N_12064);
and U13930 (N_13930,N_12172,N_12638);
or U13931 (N_13931,N_12337,N_12085);
and U13932 (N_13932,N_12555,N_12065);
or U13933 (N_13933,N_12946,N_12252);
nor U13934 (N_13934,N_12769,N_12762);
nand U13935 (N_13935,N_12139,N_12505);
nand U13936 (N_13936,N_12164,N_12464);
and U13937 (N_13937,N_12867,N_12644);
and U13938 (N_13938,N_12765,N_12239);
nor U13939 (N_13939,N_12562,N_12466);
xnor U13940 (N_13940,N_12183,N_12975);
xor U13941 (N_13941,N_12165,N_12022);
or U13942 (N_13942,N_12495,N_12334);
and U13943 (N_13943,N_12692,N_12365);
or U13944 (N_13944,N_12819,N_12951);
xor U13945 (N_13945,N_12759,N_12103);
nor U13946 (N_13946,N_12426,N_12871);
nor U13947 (N_13947,N_12559,N_12821);
xnor U13948 (N_13948,N_12415,N_12713);
and U13949 (N_13949,N_12662,N_12823);
nand U13950 (N_13950,N_12818,N_12780);
nor U13951 (N_13951,N_12605,N_12990);
nor U13952 (N_13952,N_12231,N_12744);
and U13953 (N_13953,N_12851,N_12139);
and U13954 (N_13954,N_12763,N_12874);
xor U13955 (N_13955,N_12952,N_12558);
xor U13956 (N_13956,N_12259,N_12091);
or U13957 (N_13957,N_12075,N_12998);
or U13958 (N_13958,N_12903,N_12265);
or U13959 (N_13959,N_12346,N_12753);
and U13960 (N_13960,N_12410,N_12444);
xnor U13961 (N_13961,N_12800,N_12244);
xnor U13962 (N_13962,N_12198,N_12174);
or U13963 (N_13963,N_12470,N_12493);
nand U13964 (N_13964,N_12603,N_12643);
nor U13965 (N_13965,N_12192,N_12761);
nand U13966 (N_13966,N_12282,N_12358);
xor U13967 (N_13967,N_12433,N_12003);
and U13968 (N_13968,N_12823,N_12738);
nand U13969 (N_13969,N_12845,N_12947);
xor U13970 (N_13970,N_12467,N_12984);
xnor U13971 (N_13971,N_12660,N_12902);
nand U13972 (N_13972,N_12205,N_12014);
nor U13973 (N_13973,N_12649,N_12012);
or U13974 (N_13974,N_12550,N_12398);
and U13975 (N_13975,N_12731,N_12987);
xor U13976 (N_13976,N_12683,N_12881);
or U13977 (N_13977,N_12995,N_12318);
and U13978 (N_13978,N_12715,N_12938);
and U13979 (N_13979,N_12774,N_12910);
nand U13980 (N_13980,N_12484,N_12533);
xnor U13981 (N_13981,N_12086,N_12676);
xor U13982 (N_13982,N_12226,N_12268);
nand U13983 (N_13983,N_12488,N_12754);
nor U13984 (N_13984,N_12742,N_12575);
xor U13985 (N_13985,N_12641,N_12465);
or U13986 (N_13986,N_12897,N_12266);
nor U13987 (N_13987,N_12337,N_12131);
or U13988 (N_13988,N_12067,N_12409);
xnor U13989 (N_13989,N_12663,N_12769);
xnor U13990 (N_13990,N_12211,N_12144);
and U13991 (N_13991,N_12812,N_12718);
and U13992 (N_13992,N_12692,N_12396);
nand U13993 (N_13993,N_12015,N_12121);
xor U13994 (N_13994,N_12308,N_12530);
or U13995 (N_13995,N_12774,N_12527);
and U13996 (N_13996,N_12945,N_12437);
nor U13997 (N_13997,N_12958,N_12870);
and U13998 (N_13998,N_12345,N_12732);
nand U13999 (N_13999,N_12153,N_12347);
nand U14000 (N_14000,N_13192,N_13259);
nor U14001 (N_14001,N_13733,N_13829);
nor U14002 (N_14002,N_13134,N_13734);
and U14003 (N_14003,N_13926,N_13881);
xor U14004 (N_14004,N_13189,N_13276);
or U14005 (N_14005,N_13530,N_13987);
xor U14006 (N_14006,N_13222,N_13549);
nand U14007 (N_14007,N_13520,N_13487);
nand U14008 (N_14008,N_13363,N_13080);
nor U14009 (N_14009,N_13162,N_13137);
xnor U14010 (N_14010,N_13203,N_13003);
or U14011 (N_14011,N_13286,N_13728);
and U14012 (N_14012,N_13191,N_13806);
and U14013 (N_14013,N_13117,N_13090);
or U14014 (N_14014,N_13506,N_13047);
nand U14015 (N_14015,N_13012,N_13198);
nor U14016 (N_14016,N_13292,N_13480);
and U14017 (N_14017,N_13788,N_13233);
xnor U14018 (N_14018,N_13284,N_13903);
nor U14019 (N_14019,N_13024,N_13679);
xnor U14020 (N_14020,N_13830,N_13209);
and U14021 (N_14021,N_13727,N_13256);
or U14022 (N_14022,N_13528,N_13540);
and U14023 (N_14023,N_13296,N_13025);
and U14024 (N_14024,N_13831,N_13544);
xor U14025 (N_14025,N_13581,N_13997);
nor U14026 (N_14026,N_13852,N_13768);
or U14027 (N_14027,N_13782,N_13389);
and U14028 (N_14028,N_13805,N_13247);
and U14029 (N_14029,N_13401,N_13312);
and U14030 (N_14030,N_13844,N_13622);
xor U14031 (N_14031,N_13394,N_13940);
and U14032 (N_14032,N_13238,N_13840);
or U14033 (N_14033,N_13927,N_13750);
nor U14034 (N_14034,N_13948,N_13364);
nor U14035 (N_14035,N_13217,N_13571);
nand U14036 (N_14036,N_13695,N_13241);
nand U14037 (N_14037,N_13596,N_13367);
xor U14038 (N_14038,N_13361,N_13639);
and U14039 (N_14039,N_13404,N_13803);
or U14040 (N_14040,N_13348,N_13907);
nor U14041 (N_14041,N_13490,N_13659);
nor U14042 (N_14042,N_13454,N_13166);
and U14043 (N_14043,N_13489,N_13471);
xor U14044 (N_14044,N_13475,N_13066);
nor U14045 (N_14045,N_13658,N_13625);
and U14046 (N_14046,N_13876,N_13780);
xor U14047 (N_14047,N_13666,N_13682);
nand U14048 (N_14048,N_13349,N_13763);
or U14049 (N_14049,N_13671,N_13204);
and U14050 (N_14050,N_13228,N_13350);
and U14051 (N_14051,N_13937,N_13947);
xnor U14052 (N_14052,N_13613,N_13373);
and U14053 (N_14053,N_13594,N_13512);
nor U14054 (N_14054,N_13657,N_13325);
or U14055 (N_14055,N_13163,N_13215);
nor U14056 (N_14056,N_13181,N_13150);
and U14057 (N_14057,N_13789,N_13176);
nor U14058 (N_14058,N_13158,N_13849);
nand U14059 (N_14059,N_13656,N_13774);
xnor U14060 (N_14060,N_13959,N_13161);
xnor U14061 (N_14061,N_13991,N_13764);
nor U14062 (N_14062,N_13107,N_13016);
nor U14063 (N_14063,N_13132,N_13171);
or U14064 (N_14064,N_13802,N_13328);
nand U14065 (N_14065,N_13297,N_13062);
nor U14066 (N_14066,N_13063,N_13887);
xor U14067 (N_14067,N_13989,N_13136);
and U14068 (N_14068,N_13633,N_13718);
and U14069 (N_14069,N_13413,N_13558);
and U14070 (N_14070,N_13731,N_13672);
or U14071 (N_14071,N_13023,N_13365);
and U14072 (N_14072,N_13555,N_13202);
nor U14073 (N_14073,N_13305,N_13368);
and U14074 (N_14074,N_13979,N_13482);
nor U14075 (N_14075,N_13048,N_13052);
nor U14076 (N_14076,N_13885,N_13850);
and U14077 (N_14077,N_13681,N_13152);
or U14078 (N_14078,N_13491,N_13393);
xor U14079 (N_14079,N_13443,N_13618);
and U14080 (N_14080,N_13953,N_13875);
xnor U14081 (N_14081,N_13965,N_13324);
xor U14082 (N_14082,N_13543,N_13600);
nand U14083 (N_14083,N_13472,N_13548);
nand U14084 (N_14084,N_13804,N_13356);
nand U14085 (N_14085,N_13399,N_13847);
xor U14086 (N_14086,N_13408,N_13021);
nor U14087 (N_14087,N_13624,N_13033);
and U14088 (N_14088,N_13603,N_13971);
nand U14089 (N_14089,N_13244,N_13466);
and U14090 (N_14090,N_13479,N_13485);
nor U14091 (N_14091,N_13042,N_13415);
nand U14092 (N_14092,N_13252,N_13705);
nor U14093 (N_14093,N_13470,N_13546);
nand U14094 (N_14094,N_13516,N_13142);
or U14095 (N_14095,N_13920,N_13978);
xor U14096 (N_14096,N_13535,N_13498);
nand U14097 (N_14097,N_13044,N_13330);
nand U14098 (N_14098,N_13605,N_13148);
nor U14099 (N_14099,N_13507,N_13067);
xor U14100 (N_14100,N_13901,N_13458);
or U14101 (N_14101,N_13041,N_13861);
and U14102 (N_14102,N_13029,N_13013);
or U14103 (N_14103,N_13968,N_13056);
or U14104 (N_14104,N_13468,N_13058);
xor U14105 (N_14105,N_13827,N_13122);
nand U14106 (N_14106,N_13684,N_13576);
nor U14107 (N_14107,N_13057,N_13007);
nand U14108 (N_14108,N_13869,N_13880);
and U14109 (N_14109,N_13912,N_13846);
xor U14110 (N_14110,N_13303,N_13634);
nor U14111 (N_14111,N_13429,N_13858);
nor U14112 (N_14112,N_13786,N_13329);
nand U14113 (N_14113,N_13623,N_13344);
nand U14114 (N_14114,N_13533,N_13074);
nor U14115 (N_14115,N_13434,N_13242);
xor U14116 (N_14116,N_13351,N_13323);
nor U14117 (N_14117,N_13868,N_13001);
and U14118 (N_14118,N_13385,N_13724);
nor U14119 (N_14119,N_13495,N_13065);
xor U14120 (N_14120,N_13500,N_13723);
xnor U14121 (N_14121,N_13165,N_13416);
and U14122 (N_14122,N_13983,N_13522);
nand U14123 (N_14123,N_13857,N_13932);
xnor U14124 (N_14124,N_13662,N_13197);
nor U14125 (N_14125,N_13248,N_13481);
nor U14126 (N_14126,N_13011,N_13419);
xor U14127 (N_14127,N_13668,N_13220);
or U14128 (N_14128,N_13336,N_13444);
nand U14129 (N_14129,N_13616,N_13414);
xnor U14130 (N_14130,N_13290,N_13263);
nor U14131 (N_14131,N_13588,N_13219);
nor U14132 (N_14132,N_13210,N_13697);
xor U14133 (N_14133,N_13144,N_13565);
or U14134 (N_14134,N_13924,N_13606);
or U14135 (N_14135,N_13638,N_13146);
xor U14136 (N_14136,N_13867,N_13964);
nor U14137 (N_14137,N_13039,N_13922);
xnor U14138 (N_14138,N_13185,N_13908);
nor U14139 (N_14139,N_13407,N_13494);
or U14140 (N_14140,N_13143,N_13645);
nand U14141 (N_14141,N_13539,N_13738);
xor U14142 (N_14142,N_13334,N_13730);
xnor U14143 (N_14143,N_13599,N_13164);
xnor U14144 (N_14144,N_13814,N_13227);
xor U14145 (N_14145,N_13655,N_13736);
xnor U14146 (N_14146,N_13116,N_13714);
and U14147 (N_14147,N_13905,N_13569);
nor U14148 (N_14148,N_13282,N_13902);
and U14149 (N_14149,N_13000,N_13442);
xor U14150 (N_14150,N_13870,N_13126);
xnor U14151 (N_14151,N_13726,N_13099);
nor U14152 (N_14152,N_13587,N_13376);
xor U14153 (N_14153,N_13918,N_13098);
nand U14154 (N_14154,N_13792,N_13871);
or U14155 (N_14155,N_13398,N_13196);
or U14156 (N_14156,N_13279,N_13421);
or U14157 (N_14157,N_13280,N_13317);
or U14158 (N_14158,N_13017,N_13194);
and U14159 (N_14159,N_13298,N_13936);
nor U14160 (N_14160,N_13557,N_13383);
nand U14161 (N_14161,N_13994,N_13759);
xor U14162 (N_14162,N_13627,N_13302);
xor U14163 (N_14163,N_13271,N_13182);
and U14164 (N_14164,N_13631,N_13299);
xnor U14165 (N_14165,N_13249,N_13526);
and U14166 (N_14166,N_13706,N_13583);
nand U14167 (N_14167,N_13307,N_13514);
nand U14168 (N_14168,N_13845,N_13930);
or U14169 (N_14169,N_13424,N_13493);
and U14170 (N_14170,N_13440,N_13542);
xor U14171 (N_14171,N_13878,N_13568);
or U14172 (N_14172,N_13332,N_13200);
or U14173 (N_14173,N_13295,N_13909);
and U14174 (N_14174,N_13430,N_13269);
nand U14175 (N_14175,N_13866,N_13888);
nand U14176 (N_14176,N_13151,N_13891);
xnor U14177 (N_14177,N_13283,N_13133);
and U14178 (N_14178,N_13689,N_13739);
and U14179 (N_14179,N_13545,N_13577);
xor U14180 (N_14180,N_13832,N_13050);
xor U14181 (N_14181,N_13128,N_13996);
xnor U14182 (N_14182,N_13747,N_13617);
or U14183 (N_14183,N_13713,N_13253);
xor U14184 (N_14184,N_13168,N_13221);
nand U14185 (N_14185,N_13641,N_13138);
xnor U14186 (N_14186,N_13669,N_13776);
nand U14187 (N_14187,N_13851,N_13818);
or U14188 (N_14188,N_13584,N_13499);
nor U14189 (N_14189,N_13529,N_13663);
and U14190 (N_14190,N_13860,N_13913);
xnor U14191 (N_14191,N_13127,N_13580);
or U14192 (N_14192,N_13834,N_13608);
and U14193 (N_14193,N_13147,N_13809);
xnor U14194 (N_14194,N_13826,N_13635);
or U14195 (N_14195,N_13766,N_13552);
or U14196 (N_14196,N_13790,N_13274);
nand U14197 (N_14197,N_13992,N_13883);
or U14198 (N_14198,N_13825,N_13308);
nand U14199 (N_14199,N_13748,N_13026);
xnor U14200 (N_14200,N_13962,N_13205);
xnor U14201 (N_14201,N_13423,N_13420);
or U14202 (N_14202,N_13855,N_13496);
nand U14203 (N_14203,N_13687,N_13187);
nor U14204 (N_14204,N_13793,N_13683);
nor U14205 (N_14205,N_13916,N_13534);
nor U14206 (N_14206,N_13167,N_13273);
nand U14207 (N_14207,N_13986,N_13173);
nand U14208 (N_14208,N_13155,N_13379);
xnor U14209 (N_14209,N_13245,N_13709);
and U14210 (N_14210,N_13092,N_13801);
nor U14211 (N_14211,N_13371,N_13060);
nor U14212 (N_14212,N_13783,N_13797);
and U14213 (N_14213,N_13100,N_13981);
nor U14214 (N_14214,N_13115,N_13836);
or U14215 (N_14215,N_13183,N_13536);
and U14216 (N_14216,N_13258,N_13553);
or U14217 (N_14217,N_13333,N_13833);
nor U14218 (N_14218,N_13644,N_13816);
or U14219 (N_14219,N_13114,N_13153);
and U14220 (N_14220,N_13813,N_13863);
nor U14221 (N_14221,N_13946,N_13914);
nor U14222 (N_14222,N_13751,N_13453);
nor U14223 (N_14223,N_13812,N_13199);
and U14224 (N_14224,N_13357,N_13206);
nand U14225 (N_14225,N_13717,N_13246);
nor U14226 (N_14226,N_13230,N_13752);
xnor U14227 (N_14227,N_13463,N_13770);
and U14228 (N_14228,N_13935,N_13111);
and U14229 (N_14229,N_13906,N_13340);
or U14230 (N_14230,N_13982,N_13059);
nand U14231 (N_14231,N_13360,N_13674);
or U14232 (N_14232,N_13574,N_13096);
nor U14233 (N_14233,N_13130,N_13201);
or U14234 (N_14234,N_13108,N_13642);
xnor U14235 (N_14235,N_13943,N_13698);
and U14236 (N_14236,N_13963,N_13281);
nor U14237 (N_14237,N_13769,N_13240);
xor U14238 (N_14238,N_13573,N_13208);
nand U14239 (N_14239,N_13339,N_13403);
xor U14240 (N_14240,N_13095,N_13711);
nor U14241 (N_14241,N_13380,N_13974);
xnor U14242 (N_14242,N_13139,N_13892);
and U14243 (N_14243,N_13084,N_13673);
nand U14244 (N_14244,N_13715,N_13649);
and U14245 (N_14245,N_13372,N_13076);
xnor U14246 (N_14246,N_13753,N_13945);
xnor U14247 (N_14247,N_13554,N_13452);
xnor U14248 (N_14248,N_13010,N_13938);
or U14249 (N_14249,N_13501,N_13505);
nor U14250 (N_14250,N_13619,N_13353);
or U14251 (N_14251,N_13678,N_13473);
nand U14252 (N_14252,N_13615,N_13523);
nor U14253 (N_14253,N_13400,N_13977);
and U14254 (N_14254,N_13054,N_13417);
nand U14255 (N_14255,N_13700,N_13765);
nor U14256 (N_14256,N_13510,N_13455);
and U14257 (N_14257,N_13886,N_13839);
nand U14258 (N_14258,N_13800,N_13180);
xnor U14259 (N_14259,N_13254,N_13216);
nor U14260 (N_14260,N_13664,N_13955);
or U14261 (N_14261,N_13999,N_13969);
and U14262 (N_14262,N_13218,N_13823);
nor U14263 (N_14263,N_13375,N_13984);
or U14264 (N_14264,N_13431,N_13502);
nand U14265 (N_14265,N_13951,N_13784);
nand U14266 (N_14266,N_13897,N_13118);
nor U14267 (N_14267,N_13464,N_13186);
and U14268 (N_14268,N_13824,N_13980);
nor U14269 (N_14269,N_13521,N_13022);
and U14270 (N_14270,N_13087,N_13019);
nand U14271 (N_14271,N_13449,N_13975);
and U14272 (N_14272,N_13125,N_13620);
xnor U14273 (N_14273,N_13266,N_13477);
nand U14274 (N_14274,N_13051,N_13184);
nand U14275 (N_14275,N_13676,N_13015);
and U14276 (N_14276,N_13145,N_13778);
xor U14277 (N_14277,N_13097,N_13973);
nand U14278 (N_14278,N_13355,N_13710);
or U14279 (N_14279,N_13229,N_13262);
nand U14280 (N_14280,N_13794,N_13952);
nand U14281 (N_14281,N_13175,N_13777);
or U14282 (N_14282,N_13636,N_13212);
nand U14283 (N_14283,N_13917,N_13459);
nand U14284 (N_14284,N_13313,N_13648);
nand U14285 (N_14285,N_13190,N_13395);
xor U14286 (N_14286,N_13315,N_13564);
or U14287 (N_14287,N_13411,N_13773);
nand U14288 (N_14288,N_13967,N_13749);
or U14289 (N_14289,N_13795,N_13856);
nand U14290 (N_14290,N_13094,N_13828);
nor U14291 (N_14291,N_13686,N_13582);
nand U14292 (N_14292,N_13032,N_13255);
xnor U14293 (N_14293,N_13745,N_13646);
and U14294 (N_14294,N_13744,N_13703);
nand U14295 (N_14295,N_13865,N_13559);
nor U14296 (N_14296,N_13159,N_13988);
xor U14297 (N_14297,N_13154,N_13251);
xor U14298 (N_14298,N_13289,N_13300);
or U14299 (N_14299,N_13310,N_13088);
nor U14300 (N_14300,N_13397,N_13278);
or U14301 (N_14301,N_13046,N_13425);
nand U14302 (N_14302,N_13654,N_13141);
and U14303 (N_14303,N_13838,N_13589);
nor U14304 (N_14304,N_13719,N_13607);
and U14305 (N_14305,N_13121,N_13680);
xnor U14306 (N_14306,N_13837,N_13716);
or U14307 (N_14307,N_13779,N_13864);
and U14308 (N_14308,N_13381,N_13028);
xnor U14309 (N_14309,N_13597,N_13985);
and U14310 (N_14310,N_13772,N_13515);
xor U14311 (N_14311,N_13235,N_13998);
nand U14312 (N_14312,N_13447,N_13265);
nand U14313 (N_14313,N_13223,N_13665);
nor U14314 (N_14314,N_13055,N_13661);
or U14315 (N_14315,N_13899,N_13527);
and U14316 (N_14316,N_13086,N_13882);
and U14317 (N_14317,N_13093,N_13775);
and U14318 (N_14318,N_13519,N_13586);
and U14319 (N_14319,N_13821,N_13231);
xor U14320 (N_14320,N_13049,N_13677);
nor U14321 (N_14321,N_13957,N_13848);
or U14322 (N_14322,N_13031,N_13933);
nand U14323 (N_14323,N_13740,N_13089);
xnor U14324 (N_14324,N_13105,N_13610);
nand U14325 (N_14325,N_13862,N_13091);
and U14326 (N_14326,N_13822,N_13517);
and U14327 (N_14327,N_13614,N_13072);
nand U14328 (N_14328,N_13083,N_13556);
nand U14329 (N_14329,N_13338,N_13598);
nand U14330 (N_14330,N_13541,N_13326);
nand U14331 (N_14331,N_13629,N_13359);
nand U14332 (N_14332,N_13288,N_13309);
nand U14333 (N_14333,N_13910,N_13002);
and U14334 (N_14334,N_13177,N_13889);
xnor U14335 (N_14335,N_13436,N_13810);
and U14336 (N_14336,N_13157,N_13193);
nor U14337 (N_14337,N_13304,N_13621);
nand U14338 (N_14338,N_13630,N_13369);
nand U14339 (N_14339,N_13213,N_13694);
nor U14340 (N_14340,N_13437,N_13239);
or U14341 (N_14341,N_13243,N_13040);
nor U14342 (N_14342,N_13123,N_13435);
nor U14343 (N_14343,N_13702,N_13799);
and U14344 (N_14344,N_13503,N_13699);
or U14345 (N_14345,N_13509,N_13504);
nor U14346 (N_14346,N_13426,N_13272);
nand U14347 (N_14347,N_13156,N_13101);
and U14348 (N_14348,N_13525,N_13073);
and U14349 (N_14349,N_13441,N_13585);
and U14350 (N_14350,N_13712,N_13874);
xnor U14351 (N_14351,N_13675,N_13322);
nand U14352 (N_14352,N_13064,N_13647);
xor U14353 (N_14353,N_13409,N_13257);
and U14354 (N_14354,N_13563,N_13224);
nand U14355 (N_14355,N_13035,N_13460);
nand U14356 (N_14356,N_13815,N_13593);
and U14357 (N_14357,N_13270,N_13037);
and U14358 (N_14358,N_13754,N_13391);
xnor U14359 (N_14359,N_13352,N_13537);
or U14360 (N_14360,N_13767,N_13808);
or U14361 (N_14361,N_13291,N_13082);
xnor U14362 (N_14362,N_13104,N_13457);
xnor U14363 (N_14363,N_13653,N_13928);
nor U14364 (N_14364,N_13179,N_13990);
nor U14365 (N_14365,N_13427,N_13277);
xnor U14366 (N_14366,N_13931,N_13550);
xnor U14367 (N_14367,N_13508,N_13561);
nand U14368 (N_14368,N_13894,N_13692);
and U14369 (N_14369,N_13188,N_13835);
and U14370 (N_14370,N_13112,N_13342);
nor U14371 (N_14371,N_13760,N_13318);
and U14372 (N_14372,N_13285,N_13958);
and U14373 (N_14373,N_13476,N_13070);
xor U14374 (N_14374,N_13611,N_13319);
and U14375 (N_14375,N_13178,N_13628);
xnor U14376 (N_14376,N_13036,N_13250);
nand U14377 (N_14377,N_13225,N_13428);
xor U14378 (N_14378,N_13879,N_13722);
nand U14379 (N_14379,N_13637,N_13451);
nand U14380 (N_14380,N_13884,N_13382);
or U14381 (N_14381,N_13172,N_13972);
or U14382 (N_14382,N_13562,N_13538);
nor U14383 (N_14383,N_13995,N_13798);
nand U14384 (N_14384,N_13796,N_13872);
and U14385 (N_14385,N_13954,N_13232);
and U14386 (N_14386,N_13904,N_13412);
xor U14387 (N_14387,N_13592,N_13853);
or U14388 (N_14388,N_13939,N_13018);
nand U14389 (N_14389,N_13316,N_13547);
xor U14390 (N_14390,N_13690,N_13004);
xnor U14391 (N_14391,N_13422,N_13966);
and U14392 (N_14392,N_13531,N_13729);
nand U14393 (N_14393,N_13532,N_13732);
nor U14394 (N_14394,N_13604,N_13446);
nand U14395 (N_14395,N_13120,N_13944);
xor U14396 (N_14396,N_13929,N_13014);
nor U14397 (N_14397,N_13234,N_13103);
and U14398 (N_14398,N_13934,N_13432);
or U14399 (N_14399,N_13721,N_13448);
xor U14400 (N_14400,N_13811,N_13735);
or U14401 (N_14401,N_13061,N_13077);
xor U14402 (N_14402,N_13742,N_13331);
or U14403 (N_14403,N_13819,N_13043);
xnor U14404 (N_14404,N_13691,N_13358);
and U14405 (N_14405,N_13027,N_13069);
nand U14406 (N_14406,N_13214,N_13129);
nand U14407 (N_14407,N_13685,N_13895);
xnor U14408 (N_14408,N_13113,N_13787);
xnor U14409 (N_14409,N_13950,N_13820);
nand U14410 (N_14410,N_13570,N_13439);
nor U14411 (N_14411,N_13462,N_13169);
nand U14412 (N_14412,N_13575,N_13488);
or U14413 (N_14413,N_13791,N_13890);
nor U14414 (N_14414,N_13237,N_13758);
or U14415 (N_14415,N_13260,N_13106);
nor U14416 (N_14416,N_13923,N_13696);
xnor U14417 (N_14417,N_13746,N_13942);
nor U14418 (N_14418,N_13921,N_13461);
nor U14419 (N_14419,N_13068,N_13651);
xnor U14420 (N_14420,N_13993,N_13211);
or U14421 (N_14421,N_13075,N_13560);
nor U14422 (N_14422,N_13785,N_13078);
and U14423 (N_14423,N_13377,N_13079);
nand U14424 (N_14424,N_13807,N_13226);
nor U14425 (N_14425,N_13327,N_13725);
nand U14426 (N_14426,N_13626,N_13402);
and U14427 (N_14427,N_13045,N_13406);
nand U14428 (N_14428,N_13660,N_13919);
nor U14429 (N_14429,N_13337,N_13275);
nand U14430 (N_14430,N_13781,N_13701);
xnor U14431 (N_14431,N_13707,N_13261);
xnor U14432 (N_14432,N_13450,N_13467);
nor U14433 (N_14433,N_13392,N_13590);
and U14434 (N_14434,N_13071,N_13135);
nor U14435 (N_14435,N_13433,N_13465);
xor U14436 (N_14436,N_13124,N_13484);
nor U14437 (N_14437,N_13038,N_13320);
nand U14438 (N_14438,N_13817,N_13602);
nand U14439 (N_14439,N_13418,N_13268);
and U14440 (N_14440,N_13008,N_13911);
xor U14441 (N_14441,N_13737,N_13756);
and U14442 (N_14442,N_13841,N_13497);
nand U14443 (N_14443,N_13670,N_13643);
and U14444 (N_14444,N_13362,N_13761);
nor U14445 (N_14445,N_13877,N_13961);
and U14446 (N_14446,N_13492,N_13970);
or U14447 (N_14447,N_13445,N_13843);
xor U14448 (N_14448,N_13511,N_13264);
or U14449 (N_14449,N_13667,N_13578);
nor U14450 (N_14450,N_13110,N_13306);
or U14451 (N_14451,N_13609,N_13898);
or U14452 (N_14452,N_13854,N_13207);
nand U14453 (N_14453,N_13925,N_13612);
nor U14454 (N_14454,N_13160,N_13119);
nand U14455 (N_14455,N_13566,N_13640);
or U14456 (N_14456,N_13595,N_13976);
nand U14457 (N_14457,N_13893,N_13474);
and U14458 (N_14458,N_13601,N_13354);
and U14459 (N_14459,N_13053,N_13771);
or U14460 (N_14460,N_13311,N_13518);
nand U14461 (N_14461,N_13006,N_13708);
xnor U14462 (N_14462,N_13387,N_13370);
or U14463 (N_14463,N_13301,N_13438);
and U14464 (N_14464,N_13900,N_13384);
and U14465 (N_14465,N_13693,N_13591);
nor U14466 (N_14466,N_13632,N_13567);
or U14467 (N_14467,N_13386,N_13030);
nand U14468 (N_14468,N_13650,N_13314);
xnor U14469 (N_14469,N_13949,N_13345);
nand U14470 (N_14470,N_13085,N_13896);
and U14471 (N_14471,N_13005,N_13743);
xor U14472 (N_14472,N_13346,N_13294);
nor U14473 (N_14473,N_13405,N_13149);
nor U14474 (N_14474,N_13456,N_13267);
xor U14475 (N_14475,N_13170,N_13572);
xor U14476 (N_14476,N_13688,N_13388);
nand U14477 (N_14477,N_13960,N_13335);
and U14478 (N_14478,N_13343,N_13859);
nand U14479 (N_14479,N_13741,N_13195);
nand U14480 (N_14480,N_13652,N_13321);
xnor U14481 (N_14481,N_13081,N_13410);
nor U14482 (N_14482,N_13378,N_13762);
and U14483 (N_14483,N_13524,N_13551);
nor U14484 (N_14484,N_13842,N_13131);
nor U14485 (N_14485,N_13956,N_13396);
nand U14486 (N_14486,N_13236,N_13757);
xor U14487 (N_14487,N_13720,N_13941);
nor U14488 (N_14488,N_13009,N_13755);
nor U14489 (N_14489,N_13102,N_13513);
nor U14490 (N_14490,N_13341,N_13287);
xor U14491 (N_14491,N_13478,N_13034);
xor U14492 (N_14492,N_13347,N_13109);
nand U14493 (N_14493,N_13704,N_13366);
nand U14494 (N_14494,N_13469,N_13293);
nand U14495 (N_14495,N_13486,N_13374);
nor U14496 (N_14496,N_13390,N_13174);
xnor U14497 (N_14497,N_13483,N_13140);
nor U14498 (N_14498,N_13579,N_13020);
or U14499 (N_14499,N_13873,N_13915);
nand U14500 (N_14500,N_13263,N_13166);
nor U14501 (N_14501,N_13136,N_13045);
xnor U14502 (N_14502,N_13547,N_13000);
xnor U14503 (N_14503,N_13388,N_13402);
and U14504 (N_14504,N_13368,N_13362);
or U14505 (N_14505,N_13820,N_13361);
xor U14506 (N_14506,N_13776,N_13475);
xor U14507 (N_14507,N_13150,N_13177);
and U14508 (N_14508,N_13630,N_13197);
or U14509 (N_14509,N_13057,N_13774);
nor U14510 (N_14510,N_13608,N_13585);
and U14511 (N_14511,N_13457,N_13514);
nor U14512 (N_14512,N_13154,N_13811);
xnor U14513 (N_14513,N_13708,N_13403);
nand U14514 (N_14514,N_13953,N_13446);
xnor U14515 (N_14515,N_13148,N_13640);
or U14516 (N_14516,N_13690,N_13839);
and U14517 (N_14517,N_13692,N_13707);
nand U14518 (N_14518,N_13095,N_13169);
xor U14519 (N_14519,N_13092,N_13496);
and U14520 (N_14520,N_13840,N_13695);
nand U14521 (N_14521,N_13872,N_13807);
nor U14522 (N_14522,N_13481,N_13866);
or U14523 (N_14523,N_13241,N_13570);
nand U14524 (N_14524,N_13513,N_13871);
nor U14525 (N_14525,N_13218,N_13099);
nor U14526 (N_14526,N_13577,N_13930);
and U14527 (N_14527,N_13321,N_13198);
or U14528 (N_14528,N_13250,N_13593);
xnor U14529 (N_14529,N_13659,N_13162);
nand U14530 (N_14530,N_13420,N_13826);
xnor U14531 (N_14531,N_13189,N_13412);
or U14532 (N_14532,N_13059,N_13137);
or U14533 (N_14533,N_13054,N_13194);
nand U14534 (N_14534,N_13756,N_13709);
nor U14535 (N_14535,N_13897,N_13328);
nand U14536 (N_14536,N_13973,N_13848);
xnor U14537 (N_14537,N_13517,N_13783);
nor U14538 (N_14538,N_13425,N_13833);
and U14539 (N_14539,N_13543,N_13081);
xnor U14540 (N_14540,N_13493,N_13859);
xnor U14541 (N_14541,N_13714,N_13091);
or U14542 (N_14542,N_13735,N_13509);
nand U14543 (N_14543,N_13300,N_13238);
nor U14544 (N_14544,N_13241,N_13411);
xnor U14545 (N_14545,N_13653,N_13170);
xnor U14546 (N_14546,N_13784,N_13519);
nand U14547 (N_14547,N_13757,N_13186);
and U14548 (N_14548,N_13068,N_13123);
nand U14549 (N_14549,N_13527,N_13268);
and U14550 (N_14550,N_13508,N_13960);
nand U14551 (N_14551,N_13180,N_13237);
or U14552 (N_14552,N_13054,N_13404);
xnor U14553 (N_14553,N_13437,N_13878);
and U14554 (N_14554,N_13463,N_13992);
xnor U14555 (N_14555,N_13603,N_13165);
and U14556 (N_14556,N_13672,N_13708);
nor U14557 (N_14557,N_13669,N_13903);
nand U14558 (N_14558,N_13975,N_13173);
or U14559 (N_14559,N_13468,N_13360);
or U14560 (N_14560,N_13180,N_13799);
nand U14561 (N_14561,N_13938,N_13078);
or U14562 (N_14562,N_13291,N_13585);
or U14563 (N_14563,N_13958,N_13537);
nand U14564 (N_14564,N_13637,N_13107);
xnor U14565 (N_14565,N_13267,N_13685);
and U14566 (N_14566,N_13587,N_13562);
nand U14567 (N_14567,N_13667,N_13230);
nor U14568 (N_14568,N_13865,N_13339);
and U14569 (N_14569,N_13575,N_13459);
nand U14570 (N_14570,N_13210,N_13158);
xnor U14571 (N_14571,N_13795,N_13594);
xnor U14572 (N_14572,N_13539,N_13922);
nand U14573 (N_14573,N_13262,N_13666);
nand U14574 (N_14574,N_13272,N_13799);
and U14575 (N_14575,N_13225,N_13224);
xnor U14576 (N_14576,N_13474,N_13662);
nand U14577 (N_14577,N_13535,N_13560);
nand U14578 (N_14578,N_13209,N_13338);
nor U14579 (N_14579,N_13144,N_13333);
nor U14580 (N_14580,N_13395,N_13375);
xor U14581 (N_14581,N_13307,N_13658);
nand U14582 (N_14582,N_13815,N_13211);
xnor U14583 (N_14583,N_13371,N_13839);
or U14584 (N_14584,N_13234,N_13743);
or U14585 (N_14585,N_13862,N_13626);
nand U14586 (N_14586,N_13528,N_13278);
nand U14587 (N_14587,N_13692,N_13913);
and U14588 (N_14588,N_13609,N_13764);
and U14589 (N_14589,N_13694,N_13462);
and U14590 (N_14590,N_13820,N_13390);
nand U14591 (N_14591,N_13709,N_13020);
and U14592 (N_14592,N_13267,N_13634);
nand U14593 (N_14593,N_13137,N_13851);
xor U14594 (N_14594,N_13269,N_13517);
nor U14595 (N_14595,N_13553,N_13452);
and U14596 (N_14596,N_13846,N_13847);
xnor U14597 (N_14597,N_13463,N_13587);
and U14598 (N_14598,N_13045,N_13884);
nand U14599 (N_14599,N_13101,N_13222);
xnor U14600 (N_14600,N_13902,N_13941);
nand U14601 (N_14601,N_13356,N_13940);
nor U14602 (N_14602,N_13049,N_13284);
and U14603 (N_14603,N_13589,N_13829);
or U14604 (N_14604,N_13424,N_13736);
xor U14605 (N_14605,N_13845,N_13352);
nor U14606 (N_14606,N_13834,N_13027);
or U14607 (N_14607,N_13529,N_13104);
xnor U14608 (N_14608,N_13031,N_13284);
or U14609 (N_14609,N_13005,N_13380);
and U14610 (N_14610,N_13336,N_13756);
nand U14611 (N_14611,N_13886,N_13378);
nand U14612 (N_14612,N_13831,N_13405);
and U14613 (N_14613,N_13694,N_13018);
or U14614 (N_14614,N_13804,N_13023);
xnor U14615 (N_14615,N_13416,N_13197);
nor U14616 (N_14616,N_13046,N_13952);
or U14617 (N_14617,N_13256,N_13925);
nor U14618 (N_14618,N_13232,N_13070);
nand U14619 (N_14619,N_13110,N_13388);
nor U14620 (N_14620,N_13874,N_13585);
or U14621 (N_14621,N_13724,N_13985);
nor U14622 (N_14622,N_13994,N_13724);
xnor U14623 (N_14623,N_13512,N_13206);
and U14624 (N_14624,N_13790,N_13533);
or U14625 (N_14625,N_13247,N_13674);
or U14626 (N_14626,N_13488,N_13519);
and U14627 (N_14627,N_13906,N_13495);
nand U14628 (N_14628,N_13188,N_13941);
nor U14629 (N_14629,N_13947,N_13457);
or U14630 (N_14630,N_13706,N_13279);
nand U14631 (N_14631,N_13444,N_13909);
xnor U14632 (N_14632,N_13833,N_13329);
and U14633 (N_14633,N_13235,N_13767);
nand U14634 (N_14634,N_13105,N_13363);
nand U14635 (N_14635,N_13594,N_13471);
nor U14636 (N_14636,N_13043,N_13101);
or U14637 (N_14637,N_13279,N_13366);
or U14638 (N_14638,N_13084,N_13117);
nand U14639 (N_14639,N_13938,N_13378);
nor U14640 (N_14640,N_13028,N_13810);
nand U14641 (N_14641,N_13141,N_13914);
xor U14642 (N_14642,N_13387,N_13999);
or U14643 (N_14643,N_13713,N_13197);
nor U14644 (N_14644,N_13269,N_13237);
nand U14645 (N_14645,N_13539,N_13943);
nand U14646 (N_14646,N_13810,N_13043);
and U14647 (N_14647,N_13212,N_13046);
nor U14648 (N_14648,N_13364,N_13774);
xor U14649 (N_14649,N_13015,N_13929);
xor U14650 (N_14650,N_13081,N_13225);
nor U14651 (N_14651,N_13089,N_13819);
nand U14652 (N_14652,N_13080,N_13082);
xnor U14653 (N_14653,N_13511,N_13049);
xnor U14654 (N_14654,N_13680,N_13151);
or U14655 (N_14655,N_13550,N_13967);
or U14656 (N_14656,N_13828,N_13822);
nor U14657 (N_14657,N_13787,N_13910);
and U14658 (N_14658,N_13119,N_13599);
nand U14659 (N_14659,N_13455,N_13810);
or U14660 (N_14660,N_13865,N_13806);
nor U14661 (N_14661,N_13689,N_13348);
and U14662 (N_14662,N_13818,N_13428);
xor U14663 (N_14663,N_13276,N_13469);
xnor U14664 (N_14664,N_13417,N_13135);
and U14665 (N_14665,N_13980,N_13784);
nand U14666 (N_14666,N_13700,N_13432);
or U14667 (N_14667,N_13823,N_13160);
xor U14668 (N_14668,N_13776,N_13193);
xnor U14669 (N_14669,N_13833,N_13089);
and U14670 (N_14670,N_13151,N_13911);
xor U14671 (N_14671,N_13536,N_13035);
xor U14672 (N_14672,N_13529,N_13102);
nand U14673 (N_14673,N_13779,N_13562);
xor U14674 (N_14674,N_13213,N_13207);
nor U14675 (N_14675,N_13139,N_13571);
nor U14676 (N_14676,N_13871,N_13446);
or U14677 (N_14677,N_13561,N_13165);
and U14678 (N_14678,N_13270,N_13432);
xnor U14679 (N_14679,N_13701,N_13078);
nand U14680 (N_14680,N_13000,N_13401);
nand U14681 (N_14681,N_13107,N_13112);
or U14682 (N_14682,N_13465,N_13200);
nor U14683 (N_14683,N_13644,N_13009);
nand U14684 (N_14684,N_13293,N_13235);
nor U14685 (N_14685,N_13704,N_13805);
and U14686 (N_14686,N_13828,N_13272);
and U14687 (N_14687,N_13336,N_13872);
nor U14688 (N_14688,N_13743,N_13077);
nand U14689 (N_14689,N_13318,N_13981);
or U14690 (N_14690,N_13335,N_13397);
nand U14691 (N_14691,N_13086,N_13838);
nand U14692 (N_14692,N_13455,N_13492);
nand U14693 (N_14693,N_13712,N_13658);
and U14694 (N_14694,N_13964,N_13256);
nor U14695 (N_14695,N_13495,N_13452);
and U14696 (N_14696,N_13133,N_13743);
nand U14697 (N_14697,N_13055,N_13925);
xnor U14698 (N_14698,N_13004,N_13694);
or U14699 (N_14699,N_13911,N_13761);
nor U14700 (N_14700,N_13512,N_13722);
nor U14701 (N_14701,N_13950,N_13217);
and U14702 (N_14702,N_13824,N_13973);
xnor U14703 (N_14703,N_13629,N_13845);
or U14704 (N_14704,N_13727,N_13408);
nand U14705 (N_14705,N_13813,N_13508);
xor U14706 (N_14706,N_13713,N_13171);
and U14707 (N_14707,N_13061,N_13149);
or U14708 (N_14708,N_13896,N_13004);
and U14709 (N_14709,N_13891,N_13356);
nand U14710 (N_14710,N_13065,N_13564);
or U14711 (N_14711,N_13910,N_13781);
or U14712 (N_14712,N_13390,N_13254);
nand U14713 (N_14713,N_13182,N_13934);
xor U14714 (N_14714,N_13671,N_13534);
and U14715 (N_14715,N_13429,N_13771);
and U14716 (N_14716,N_13474,N_13366);
and U14717 (N_14717,N_13736,N_13919);
nor U14718 (N_14718,N_13444,N_13250);
or U14719 (N_14719,N_13967,N_13994);
nor U14720 (N_14720,N_13934,N_13913);
nand U14721 (N_14721,N_13536,N_13595);
xnor U14722 (N_14722,N_13555,N_13913);
xor U14723 (N_14723,N_13747,N_13984);
and U14724 (N_14724,N_13598,N_13110);
xor U14725 (N_14725,N_13113,N_13954);
nand U14726 (N_14726,N_13350,N_13780);
nor U14727 (N_14727,N_13584,N_13207);
nand U14728 (N_14728,N_13288,N_13793);
and U14729 (N_14729,N_13999,N_13214);
and U14730 (N_14730,N_13155,N_13969);
and U14731 (N_14731,N_13109,N_13623);
and U14732 (N_14732,N_13261,N_13957);
nand U14733 (N_14733,N_13188,N_13552);
nand U14734 (N_14734,N_13068,N_13212);
and U14735 (N_14735,N_13022,N_13224);
xor U14736 (N_14736,N_13063,N_13694);
nor U14737 (N_14737,N_13197,N_13101);
nand U14738 (N_14738,N_13733,N_13209);
nor U14739 (N_14739,N_13621,N_13348);
and U14740 (N_14740,N_13807,N_13248);
nor U14741 (N_14741,N_13195,N_13177);
xnor U14742 (N_14742,N_13096,N_13430);
nand U14743 (N_14743,N_13103,N_13354);
xor U14744 (N_14744,N_13610,N_13391);
nor U14745 (N_14745,N_13634,N_13779);
xnor U14746 (N_14746,N_13949,N_13720);
nor U14747 (N_14747,N_13535,N_13582);
and U14748 (N_14748,N_13440,N_13482);
nand U14749 (N_14749,N_13594,N_13830);
xor U14750 (N_14750,N_13622,N_13046);
nand U14751 (N_14751,N_13965,N_13498);
nand U14752 (N_14752,N_13348,N_13664);
or U14753 (N_14753,N_13112,N_13569);
or U14754 (N_14754,N_13208,N_13912);
nand U14755 (N_14755,N_13543,N_13838);
nor U14756 (N_14756,N_13109,N_13801);
xor U14757 (N_14757,N_13318,N_13464);
or U14758 (N_14758,N_13082,N_13195);
or U14759 (N_14759,N_13151,N_13428);
or U14760 (N_14760,N_13577,N_13257);
or U14761 (N_14761,N_13989,N_13105);
nor U14762 (N_14762,N_13529,N_13300);
nor U14763 (N_14763,N_13839,N_13298);
and U14764 (N_14764,N_13089,N_13463);
or U14765 (N_14765,N_13184,N_13428);
nand U14766 (N_14766,N_13807,N_13405);
nor U14767 (N_14767,N_13852,N_13453);
or U14768 (N_14768,N_13661,N_13063);
or U14769 (N_14769,N_13778,N_13618);
xnor U14770 (N_14770,N_13258,N_13161);
nand U14771 (N_14771,N_13059,N_13761);
nand U14772 (N_14772,N_13100,N_13932);
and U14773 (N_14773,N_13517,N_13970);
nand U14774 (N_14774,N_13880,N_13457);
nand U14775 (N_14775,N_13833,N_13151);
nor U14776 (N_14776,N_13743,N_13764);
and U14777 (N_14777,N_13068,N_13735);
nand U14778 (N_14778,N_13423,N_13337);
xor U14779 (N_14779,N_13263,N_13311);
and U14780 (N_14780,N_13801,N_13071);
nor U14781 (N_14781,N_13719,N_13785);
nor U14782 (N_14782,N_13629,N_13689);
xnor U14783 (N_14783,N_13234,N_13502);
xnor U14784 (N_14784,N_13251,N_13613);
or U14785 (N_14785,N_13184,N_13797);
xnor U14786 (N_14786,N_13234,N_13246);
xnor U14787 (N_14787,N_13925,N_13854);
and U14788 (N_14788,N_13731,N_13598);
xor U14789 (N_14789,N_13265,N_13365);
or U14790 (N_14790,N_13557,N_13433);
nand U14791 (N_14791,N_13742,N_13374);
nor U14792 (N_14792,N_13210,N_13815);
and U14793 (N_14793,N_13104,N_13666);
nand U14794 (N_14794,N_13897,N_13531);
and U14795 (N_14795,N_13204,N_13520);
or U14796 (N_14796,N_13829,N_13451);
or U14797 (N_14797,N_13694,N_13674);
or U14798 (N_14798,N_13282,N_13105);
and U14799 (N_14799,N_13600,N_13590);
or U14800 (N_14800,N_13183,N_13210);
and U14801 (N_14801,N_13155,N_13913);
nand U14802 (N_14802,N_13746,N_13930);
and U14803 (N_14803,N_13308,N_13335);
and U14804 (N_14804,N_13211,N_13060);
xor U14805 (N_14805,N_13205,N_13141);
nor U14806 (N_14806,N_13634,N_13025);
nand U14807 (N_14807,N_13008,N_13669);
xor U14808 (N_14808,N_13495,N_13026);
nand U14809 (N_14809,N_13607,N_13008);
and U14810 (N_14810,N_13493,N_13029);
xor U14811 (N_14811,N_13942,N_13107);
and U14812 (N_14812,N_13856,N_13782);
nand U14813 (N_14813,N_13473,N_13581);
xnor U14814 (N_14814,N_13877,N_13641);
xnor U14815 (N_14815,N_13167,N_13691);
nor U14816 (N_14816,N_13553,N_13948);
nand U14817 (N_14817,N_13985,N_13519);
nor U14818 (N_14818,N_13909,N_13553);
or U14819 (N_14819,N_13346,N_13577);
or U14820 (N_14820,N_13998,N_13912);
or U14821 (N_14821,N_13158,N_13775);
xor U14822 (N_14822,N_13594,N_13402);
xor U14823 (N_14823,N_13500,N_13391);
xor U14824 (N_14824,N_13698,N_13272);
xnor U14825 (N_14825,N_13498,N_13608);
xnor U14826 (N_14826,N_13773,N_13093);
nor U14827 (N_14827,N_13263,N_13559);
xnor U14828 (N_14828,N_13602,N_13273);
and U14829 (N_14829,N_13122,N_13066);
nand U14830 (N_14830,N_13840,N_13000);
xor U14831 (N_14831,N_13330,N_13291);
and U14832 (N_14832,N_13920,N_13873);
nand U14833 (N_14833,N_13018,N_13626);
xor U14834 (N_14834,N_13721,N_13510);
nor U14835 (N_14835,N_13028,N_13370);
or U14836 (N_14836,N_13541,N_13282);
and U14837 (N_14837,N_13513,N_13466);
nand U14838 (N_14838,N_13002,N_13095);
and U14839 (N_14839,N_13684,N_13612);
nor U14840 (N_14840,N_13501,N_13688);
or U14841 (N_14841,N_13997,N_13360);
and U14842 (N_14842,N_13469,N_13010);
xor U14843 (N_14843,N_13836,N_13322);
and U14844 (N_14844,N_13126,N_13525);
or U14845 (N_14845,N_13400,N_13678);
xnor U14846 (N_14846,N_13653,N_13572);
xor U14847 (N_14847,N_13431,N_13707);
xnor U14848 (N_14848,N_13845,N_13541);
nor U14849 (N_14849,N_13381,N_13940);
and U14850 (N_14850,N_13822,N_13292);
nor U14851 (N_14851,N_13257,N_13160);
nor U14852 (N_14852,N_13464,N_13980);
xor U14853 (N_14853,N_13339,N_13927);
and U14854 (N_14854,N_13251,N_13253);
nor U14855 (N_14855,N_13256,N_13149);
nand U14856 (N_14856,N_13469,N_13782);
xnor U14857 (N_14857,N_13431,N_13814);
xor U14858 (N_14858,N_13581,N_13102);
nor U14859 (N_14859,N_13917,N_13259);
and U14860 (N_14860,N_13905,N_13980);
nand U14861 (N_14861,N_13280,N_13546);
or U14862 (N_14862,N_13181,N_13533);
xor U14863 (N_14863,N_13272,N_13031);
and U14864 (N_14864,N_13623,N_13892);
nand U14865 (N_14865,N_13704,N_13614);
xnor U14866 (N_14866,N_13895,N_13686);
or U14867 (N_14867,N_13013,N_13425);
nand U14868 (N_14868,N_13082,N_13394);
nand U14869 (N_14869,N_13164,N_13404);
and U14870 (N_14870,N_13066,N_13847);
nand U14871 (N_14871,N_13487,N_13491);
nor U14872 (N_14872,N_13287,N_13822);
nor U14873 (N_14873,N_13279,N_13077);
xnor U14874 (N_14874,N_13458,N_13983);
or U14875 (N_14875,N_13477,N_13816);
nand U14876 (N_14876,N_13518,N_13420);
and U14877 (N_14877,N_13719,N_13998);
xnor U14878 (N_14878,N_13696,N_13787);
and U14879 (N_14879,N_13932,N_13501);
nor U14880 (N_14880,N_13806,N_13388);
nand U14881 (N_14881,N_13700,N_13526);
and U14882 (N_14882,N_13228,N_13977);
nand U14883 (N_14883,N_13419,N_13835);
or U14884 (N_14884,N_13898,N_13983);
nand U14885 (N_14885,N_13997,N_13795);
and U14886 (N_14886,N_13944,N_13704);
xnor U14887 (N_14887,N_13809,N_13982);
or U14888 (N_14888,N_13760,N_13116);
nand U14889 (N_14889,N_13857,N_13828);
and U14890 (N_14890,N_13034,N_13538);
nor U14891 (N_14891,N_13048,N_13977);
nand U14892 (N_14892,N_13775,N_13254);
nor U14893 (N_14893,N_13579,N_13278);
or U14894 (N_14894,N_13150,N_13029);
or U14895 (N_14895,N_13604,N_13650);
or U14896 (N_14896,N_13396,N_13167);
xnor U14897 (N_14897,N_13802,N_13442);
xnor U14898 (N_14898,N_13539,N_13292);
nand U14899 (N_14899,N_13047,N_13873);
nor U14900 (N_14900,N_13488,N_13219);
nor U14901 (N_14901,N_13596,N_13666);
or U14902 (N_14902,N_13845,N_13967);
or U14903 (N_14903,N_13797,N_13212);
xor U14904 (N_14904,N_13271,N_13236);
nor U14905 (N_14905,N_13366,N_13840);
nand U14906 (N_14906,N_13237,N_13118);
or U14907 (N_14907,N_13926,N_13247);
nor U14908 (N_14908,N_13629,N_13928);
nor U14909 (N_14909,N_13419,N_13844);
and U14910 (N_14910,N_13312,N_13580);
and U14911 (N_14911,N_13313,N_13337);
and U14912 (N_14912,N_13083,N_13724);
and U14913 (N_14913,N_13379,N_13344);
nor U14914 (N_14914,N_13559,N_13386);
or U14915 (N_14915,N_13837,N_13619);
or U14916 (N_14916,N_13583,N_13350);
nand U14917 (N_14917,N_13928,N_13241);
or U14918 (N_14918,N_13434,N_13970);
nor U14919 (N_14919,N_13133,N_13576);
or U14920 (N_14920,N_13497,N_13007);
nand U14921 (N_14921,N_13085,N_13564);
and U14922 (N_14922,N_13275,N_13397);
or U14923 (N_14923,N_13541,N_13504);
nor U14924 (N_14924,N_13312,N_13170);
nand U14925 (N_14925,N_13244,N_13030);
nand U14926 (N_14926,N_13453,N_13033);
nor U14927 (N_14927,N_13307,N_13212);
xnor U14928 (N_14928,N_13265,N_13768);
or U14929 (N_14929,N_13089,N_13469);
nand U14930 (N_14930,N_13251,N_13816);
nand U14931 (N_14931,N_13852,N_13359);
nand U14932 (N_14932,N_13374,N_13510);
xor U14933 (N_14933,N_13073,N_13405);
and U14934 (N_14934,N_13120,N_13288);
nor U14935 (N_14935,N_13518,N_13885);
nand U14936 (N_14936,N_13916,N_13316);
nor U14937 (N_14937,N_13525,N_13832);
nor U14938 (N_14938,N_13658,N_13147);
xnor U14939 (N_14939,N_13678,N_13770);
and U14940 (N_14940,N_13391,N_13000);
nor U14941 (N_14941,N_13492,N_13522);
xor U14942 (N_14942,N_13599,N_13474);
and U14943 (N_14943,N_13064,N_13584);
and U14944 (N_14944,N_13782,N_13487);
or U14945 (N_14945,N_13194,N_13725);
nand U14946 (N_14946,N_13745,N_13882);
or U14947 (N_14947,N_13774,N_13273);
or U14948 (N_14948,N_13657,N_13733);
xnor U14949 (N_14949,N_13067,N_13241);
or U14950 (N_14950,N_13197,N_13423);
nor U14951 (N_14951,N_13173,N_13378);
or U14952 (N_14952,N_13627,N_13296);
or U14953 (N_14953,N_13798,N_13689);
or U14954 (N_14954,N_13638,N_13980);
nand U14955 (N_14955,N_13763,N_13941);
xor U14956 (N_14956,N_13501,N_13888);
nor U14957 (N_14957,N_13605,N_13129);
and U14958 (N_14958,N_13823,N_13441);
nor U14959 (N_14959,N_13131,N_13240);
and U14960 (N_14960,N_13009,N_13289);
nand U14961 (N_14961,N_13412,N_13259);
and U14962 (N_14962,N_13323,N_13913);
nand U14963 (N_14963,N_13462,N_13470);
xnor U14964 (N_14964,N_13068,N_13994);
xor U14965 (N_14965,N_13871,N_13239);
and U14966 (N_14966,N_13605,N_13444);
or U14967 (N_14967,N_13117,N_13402);
xor U14968 (N_14968,N_13924,N_13255);
or U14969 (N_14969,N_13159,N_13901);
xnor U14970 (N_14970,N_13727,N_13964);
or U14971 (N_14971,N_13983,N_13313);
nand U14972 (N_14972,N_13603,N_13955);
or U14973 (N_14973,N_13903,N_13423);
or U14974 (N_14974,N_13805,N_13107);
nor U14975 (N_14975,N_13110,N_13669);
nor U14976 (N_14976,N_13168,N_13072);
nor U14977 (N_14977,N_13811,N_13393);
or U14978 (N_14978,N_13314,N_13304);
nor U14979 (N_14979,N_13196,N_13844);
xnor U14980 (N_14980,N_13260,N_13991);
nand U14981 (N_14981,N_13957,N_13256);
nor U14982 (N_14982,N_13554,N_13081);
nor U14983 (N_14983,N_13635,N_13119);
nor U14984 (N_14984,N_13532,N_13849);
and U14985 (N_14985,N_13617,N_13931);
or U14986 (N_14986,N_13635,N_13005);
xnor U14987 (N_14987,N_13958,N_13128);
and U14988 (N_14988,N_13608,N_13614);
xnor U14989 (N_14989,N_13168,N_13487);
nor U14990 (N_14990,N_13303,N_13704);
and U14991 (N_14991,N_13840,N_13404);
and U14992 (N_14992,N_13096,N_13008);
or U14993 (N_14993,N_13411,N_13669);
xor U14994 (N_14994,N_13488,N_13762);
nand U14995 (N_14995,N_13104,N_13389);
nand U14996 (N_14996,N_13982,N_13390);
and U14997 (N_14997,N_13121,N_13673);
and U14998 (N_14998,N_13748,N_13738);
nor U14999 (N_14999,N_13146,N_13940);
and UO_0 (O_0,N_14902,N_14673);
and UO_1 (O_1,N_14017,N_14433);
xnor UO_2 (O_2,N_14863,N_14552);
nor UO_3 (O_3,N_14899,N_14698);
nor UO_4 (O_4,N_14199,N_14313);
or UO_5 (O_5,N_14892,N_14827);
nand UO_6 (O_6,N_14461,N_14364);
nor UO_7 (O_7,N_14343,N_14327);
and UO_8 (O_8,N_14918,N_14039);
xnor UO_9 (O_9,N_14751,N_14384);
nand UO_10 (O_10,N_14911,N_14415);
or UO_11 (O_11,N_14425,N_14897);
and UO_12 (O_12,N_14663,N_14968);
or UO_13 (O_13,N_14450,N_14641);
xnor UO_14 (O_14,N_14607,N_14989);
nor UO_15 (O_15,N_14920,N_14851);
or UO_16 (O_16,N_14981,N_14729);
and UO_17 (O_17,N_14620,N_14515);
or UO_18 (O_18,N_14967,N_14001);
xor UO_19 (O_19,N_14361,N_14690);
and UO_20 (O_20,N_14516,N_14168);
nand UO_21 (O_21,N_14209,N_14134);
and UO_22 (O_22,N_14426,N_14443);
nor UO_23 (O_23,N_14606,N_14195);
nor UO_24 (O_24,N_14359,N_14446);
and UO_25 (O_25,N_14308,N_14869);
nand UO_26 (O_26,N_14024,N_14783);
xnor UO_27 (O_27,N_14182,N_14662);
nand UO_28 (O_28,N_14848,N_14362);
and UO_29 (O_29,N_14575,N_14177);
or UO_30 (O_30,N_14345,N_14850);
xnor UO_31 (O_31,N_14337,N_14153);
nor UO_32 (O_32,N_14772,N_14432);
nor UO_33 (O_33,N_14538,N_14975);
nand UO_34 (O_34,N_14984,N_14581);
xnor UO_35 (O_35,N_14256,N_14929);
or UO_36 (O_36,N_14739,N_14665);
or UO_37 (O_37,N_14298,N_14315);
xor UO_38 (O_38,N_14936,N_14037);
and UO_39 (O_39,N_14189,N_14015);
and UO_40 (O_40,N_14213,N_14716);
or UO_41 (O_41,N_14499,N_14473);
or UO_42 (O_42,N_14556,N_14097);
nand UO_43 (O_43,N_14992,N_14796);
and UO_44 (O_44,N_14595,N_14890);
xnor UO_45 (O_45,N_14070,N_14903);
nand UO_46 (O_46,N_14533,N_14616);
or UO_47 (O_47,N_14314,N_14676);
xor UO_48 (O_48,N_14323,N_14059);
xor UO_49 (O_49,N_14321,N_14420);
nor UO_50 (O_50,N_14789,N_14760);
nor UO_51 (O_51,N_14683,N_14378);
nor UO_52 (O_52,N_14646,N_14471);
xor UO_53 (O_53,N_14476,N_14181);
and UO_54 (O_54,N_14470,N_14974);
nor UO_55 (O_55,N_14843,N_14222);
or UO_56 (O_56,N_14639,N_14108);
or UO_57 (O_57,N_14293,N_14688);
nand UO_58 (O_58,N_14464,N_14336);
nor UO_59 (O_59,N_14174,N_14221);
nand UO_60 (O_60,N_14808,N_14083);
xor UO_61 (O_61,N_14139,N_14949);
nand UO_62 (O_62,N_14160,N_14413);
nor UO_63 (O_63,N_14368,N_14834);
nor UO_64 (O_64,N_14236,N_14370);
nor UO_65 (O_65,N_14363,N_14303);
and UO_66 (O_66,N_14854,N_14360);
nor UO_67 (O_67,N_14574,N_14089);
or UO_68 (O_68,N_14332,N_14561);
xnor UO_69 (O_69,N_14594,N_14410);
nand UO_70 (O_70,N_14468,N_14535);
nor UO_71 (O_71,N_14232,N_14794);
xnor UO_72 (O_72,N_14054,N_14955);
or UO_73 (O_73,N_14365,N_14034);
xor UO_74 (O_74,N_14756,N_14735);
and UO_75 (O_75,N_14478,N_14479);
and UO_76 (O_76,N_14144,N_14304);
nand UO_77 (O_77,N_14094,N_14996);
nand UO_78 (O_78,N_14073,N_14386);
and UO_79 (O_79,N_14769,N_14529);
nor UO_80 (O_80,N_14489,N_14084);
xnor UO_81 (O_81,N_14583,N_14826);
nand UO_82 (O_82,N_14009,N_14693);
or UO_83 (O_83,N_14328,N_14914);
nor UO_84 (O_84,N_14238,N_14734);
nor UO_85 (O_85,N_14400,N_14109);
xor UO_86 (O_86,N_14008,N_14709);
and UO_87 (O_87,N_14483,N_14422);
nand UO_88 (O_88,N_14078,N_14952);
nor UO_89 (O_89,N_14490,N_14625);
nor UO_90 (O_90,N_14654,N_14119);
nor UO_91 (O_91,N_14136,N_14496);
nor UO_92 (O_92,N_14130,N_14966);
nor UO_93 (O_93,N_14995,N_14273);
or UO_94 (O_94,N_14985,N_14255);
nand UO_95 (O_95,N_14823,N_14220);
xnor UO_96 (O_96,N_14312,N_14960);
xnor UO_97 (O_97,N_14014,N_14669);
xor UO_98 (O_98,N_14055,N_14069);
xnor UO_99 (O_99,N_14656,N_14212);
xnor UO_100 (O_100,N_14472,N_14586);
nor UO_101 (O_101,N_14598,N_14839);
nand UO_102 (O_102,N_14736,N_14539);
or UO_103 (O_103,N_14604,N_14987);
and UO_104 (O_104,N_14747,N_14117);
and UO_105 (O_105,N_14243,N_14133);
or UO_106 (O_106,N_14605,N_14185);
or UO_107 (O_107,N_14068,N_14947);
or UO_108 (O_108,N_14946,N_14439);
nor UO_109 (O_109,N_14274,N_14610);
nor UO_110 (O_110,N_14513,N_14237);
nand UO_111 (O_111,N_14146,N_14272);
and UO_112 (O_112,N_14804,N_14099);
and UO_113 (O_113,N_14079,N_14532);
xor UO_114 (O_114,N_14460,N_14910);
or UO_115 (O_115,N_14506,N_14307);
nand UO_116 (O_116,N_14397,N_14294);
nand UO_117 (O_117,N_14667,N_14445);
or UO_118 (O_118,N_14487,N_14994);
nor UO_119 (O_119,N_14281,N_14093);
or UO_120 (O_120,N_14201,N_14339);
nor UO_121 (O_121,N_14208,N_14251);
or UO_122 (O_122,N_14018,N_14585);
xor UO_123 (O_123,N_14699,N_14777);
or UO_124 (O_124,N_14558,N_14706);
nor UO_125 (O_125,N_14036,N_14951);
nand UO_126 (O_126,N_14191,N_14675);
nand UO_127 (O_127,N_14424,N_14806);
xnor UO_128 (O_128,N_14141,N_14940);
and UO_129 (O_129,N_14879,N_14052);
nor UO_130 (O_130,N_14697,N_14395);
or UO_131 (O_131,N_14020,N_14053);
xor UO_132 (O_132,N_14098,N_14818);
xnor UO_133 (O_133,N_14322,N_14309);
or UO_134 (O_134,N_14265,N_14239);
xor UO_135 (O_135,N_14335,N_14188);
or UO_136 (O_136,N_14531,N_14548);
and UO_137 (O_137,N_14354,N_14534);
nor UO_138 (O_138,N_14569,N_14252);
xnor UO_139 (O_139,N_14026,N_14393);
and UO_140 (O_140,N_14830,N_14846);
xor UO_141 (O_141,N_14775,N_14124);
or UO_142 (O_142,N_14738,N_14280);
or UO_143 (O_143,N_14891,N_14922);
nor UO_144 (O_144,N_14787,N_14670);
and UO_145 (O_145,N_14025,N_14888);
nand UO_146 (O_146,N_14447,N_14927);
nor UO_147 (O_147,N_14710,N_14958);
nor UO_148 (O_148,N_14862,N_14828);
nor UO_149 (O_149,N_14455,N_14442);
nor UO_150 (O_150,N_14833,N_14044);
nor UO_151 (O_151,N_14745,N_14644);
nand UO_152 (O_152,N_14712,N_14061);
and UO_153 (O_153,N_14835,N_14492);
nand UO_154 (O_154,N_14408,N_14629);
nor UO_155 (O_155,N_14123,N_14715);
nand UO_156 (O_156,N_14825,N_14022);
or UO_157 (O_157,N_14887,N_14138);
nand UO_158 (O_158,N_14921,N_14633);
or UO_159 (O_159,N_14596,N_14795);
or UO_160 (O_160,N_14250,N_14925);
or UO_161 (O_161,N_14728,N_14986);
and UO_162 (O_162,N_14101,N_14741);
and UO_163 (O_163,N_14650,N_14873);
nand UO_164 (O_164,N_14132,N_14349);
and UO_165 (O_165,N_14584,N_14111);
and UO_166 (O_166,N_14474,N_14112);
nor UO_167 (O_167,N_14456,N_14901);
nor UO_168 (O_168,N_14032,N_14771);
nand UO_169 (O_169,N_14567,N_14626);
nand UO_170 (O_170,N_14029,N_14628);
xor UO_171 (O_171,N_14469,N_14190);
or UO_172 (O_172,N_14800,N_14198);
or UO_173 (O_173,N_14245,N_14963);
nor UO_174 (O_174,N_14493,N_14329);
xnor UO_175 (O_175,N_14216,N_14497);
xor UO_176 (O_176,N_14878,N_14318);
or UO_177 (O_177,N_14856,N_14341);
nand UO_178 (O_178,N_14935,N_14276);
xnor UO_179 (O_179,N_14217,N_14137);
xor UO_180 (O_180,N_14151,N_14350);
nand UO_181 (O_181,N_14021,N_14707);
xnor UO_182 (O_182,N_14344,N_14288);
and UO_183 (O_183,N_14708,N_14803);
xor UO_184 (O_184,N_14353,N_14161);
nor UO_185 (O_185,N_14486,N_14525);
nand UO_186 (O_186,N_14352,N_14689);
nand UO_187 (O_187,N_14781,N_14809);
nand UO_188 (O_188,N_14271,N_14300);
and UO_189 (O_189,N_14617,N_14430);
nor UO_190 (O_190,N_14909,N_14466);
nand UO_191 (O_191,N_14356,N_14224);
nor UO_192 (O_192,N_14778,N_14319);
nand UO_193 (O_193,N_14202,N_14253);
or UO_194 (O_194,N_14701,N_14045);
and UO_195 (O_195,N_14748,N_14269);
or UO_196 (O_196,N_14228,N_14553);
nor UO_197 (O_197,N_14085,N_14559);
nand UO_198 (O_198,N_14358,N_14006);
nor UO_199 (O_199,N_14346,N_14609);
nor UO_200 (O_200,N_14286,N_14964);
nor UO_201 (O_201,N_14999,N_14126);
xor UO_202 (O_202,N_14743,N_14782);
nor UO_203 (O_203,N_14776,N_14714);
nand UO_204 (O_204,N_14376,N_14155);
xnor UO_205 (O_205,N_14417,N_14591);
nor UO_206 (O_206,N_14284,N_14991);
nand UO_207 (O_207,N_14260,N_14159);
nand UO_208 (O_208,N_14779,N_14150);
or UO_209 (O_209,N_14234,N_14171);
or UO_210 (O_210,N_14791,N_14204);
nor UO_211 (O_211,N_14719,N_14064);
and UO_212 (O_212,N_14580,N_14379);
and UO_213 (O_213,N_14692,N_14816);
and UO_214 (O_214,N_14900,N_14545);
nand UO_215 (O_215,N_14416,N_14720);
xnor UO_216 (O_216,N_14162,N_14399);
or UO_217 (O_217,N_14428,N_14458);
nand UO_218 (O_218,N_14577,N_14687);
nand UO_219 (O_219,N_14454,N_14128);
or UO_220 (O_220,N_14564,N_14419);
or UO_221 (O_221,N_14223,N_14576);
or UO_222 (O_222,N_14131,N_14904);
nand UO_223 (O_223,N_14792,N_14031);
nor UO_224 (O_224,N_14305,N_14810);
nand UO_225 (O_225,N_14934,N_14167);
or UO_226 (O_226,N_14761,N_14510);
nand UO_227 (O_227,N_14722,N_14965);
and UO_228 (O_228,N_14297,N_14630);
xor UO_229 (O_229,N_14401,N_14624);
and UO_230 (O_230,N_14407,N_14435);
xnor UO_231 (O_231,N_14140,N_14868);
and UO_232 (O_232,N_14763,N_14842);
nor UO_233 (O_233,N_14819,N_14019);
or UO_234 (O_234,N_14291,N_14523);
or UO_235 (O_235,N_14330,N_14671);
nand UO_236 (O_236,N_14342,N_14048);
and UO_237 (O_237,N_14896,N_14512);
or UO_238 (O_238,N_14257,N_14311);
nor UO_239 (O_239,N_14495,N_14480);
or UO_240 (O_240,N_14773,N_14095);
xor UO_241 (O_241,N_14589,N_14638);
nor UO_242 (O_242,N_14814,N_14731);
or UO_243 (O_243,N_14649,N_14831);
or UO_244 (O_244,N_14742,N_14861);
xnor UO_245 (O_245,N_14369,N_14917);
nor UO_246 (O_246,N_14829,N_14732);
nand UO_247 (O_247,N_14081,N_14973);
nand UO_248 (O_248,N_14259,N_14355);
xor UO_249 (O_249,N_14267,N_14895);
or UO_250 (O_250,N_14954,N_14175);
nor UO_251 (O_251,N_14622,N_14103);
and UO_252 (O_252,N_14824,N_14429);
nor UO_253 (O_253,N_14923,N_14270);
nor UO_254 (O_254,N_14755,N_14075);
nand UO_255 (O_255,N_14858,N_14972);
or UO_256 (O_256,N_14404,N_14956);
and UO_257 (O_257,N_14587,N_14263);
xor UO_258 (O_258,N_14682,N_14549);
or UO_259 (O_259,N_14522,N_14411);
xnor UO_260 (O_260,N_14579,N_14340);
xnor UO_261 (O_261,N_14333,N_14551);
nor UO_262 (O_262,N_14813,N_14431);
nand UO_263 (O_263,N_14718,N_14636);
xnor UO_264 (O_264,N_14864,N_14046);
nand UO_265 (O_265,N_14684,N_14441);
xor UO_266 (O_266,N_14027,N_14105);
or UO_267 (O_267,N_14939,N_14158);
nand UO_268 (O_268,N_14012,N_14334);
nand UO_269 (O_269,N_14528,N_14004);
nor UO_270 (O_270,N_14893,N_14645);
xnor UO_271 (O_271,N_14647,N_14325);
and UO_272 (O_272,N_14268,N_14932);
xor UO_273 (O_273,N_14801,N_14230);
and UO_274 (O_274,N_14127,N_14142);
and UO_275 (O_275,N_14717,N_14740);
nor UO_276 (O_276,N_14184,N_14180);
xor UO_277 (O_277,N_14049,N_14320);
xnor UO_278 (O_278,N_14383,N_14568);
nor UO_279 (O_279,N_14302,N_14953);
xor UO_280 (O_280,N_14933,N_14076);
nand UO_281 (O_281,N_14603,N_14744);
and UO_282 (O_282,N_14519,N_14860);
or UO_283 (O_283,N_14685,N_14853);
nand UO_284 (O_284,N_14143,N_14948);
or UO_285 (O_285,N_14874,N_14241);
nand UO_286 (O_286,N_14149,N_14266);
nor UO_287 (O_287,N_14723,N_14950);
and UO_288 (O_288,N_14657,N_14894);
nand UO_289 (O_289,N_14942,N_14324);
xor UO_290 (O_290,N_14530,N_14058);
xnor UO_291 (O_291,N_14477,N_14805);
or UO_292 (O_292,N_14821,N_14348);
and UO_293 (O_293,N_14387,N_14372);
nor UO_294 (O_294,N_14043,N_14926);
and UO_295 (O_295,N_14962,N_14106);
nor UO_296 (O_296,N_14852,N_14375);
or UO_297 (O_297,N_14406,N_14067);
and UO_298 (O_298,N_14766,N_14060);
nor UO_299 (O_299,N_14409,N_14283);
nor UO_300 (O_300,N_14380,N_14357);
or UO_301 (O_301,N_14062,N_14886);
and UO_302 (O_302,N_14700,N_14543);
and UO_303 (O_303,N_14997,N_14453);
nand UO_304 (O_304,N_14659,N_14176);
and UO_305 (O_305,N_14215,N_14640);
nand UO_306 (O_306,N_14865,N_14990);
nor UO_307 (O_307,N_14203,N_14437);
nand UO_308 (O_308,N_14871,N_14817);
nor UO_309 (O_309,N_14005,N_14277);
and UO_310 (O_310,N_14642,N_14347);
or UO_311 (O_311,N_14086,N_14767);
xor UO_312 (O_312,N_14571,N_14292);
xnor UO_313 (O_313,N_14811,N_14163);
nand UO_314 (O_314,N_14310,N_14050);
or UO_315 (O_315,N_14841,N_14233);
nor UO_316 (O_316,N_14679,N_14517);
nor UO_317 (O_317,N_14875,N_14883);
nor UO_318 (O_318,N_14979,N_14110);
nand UO_319 (O_319,N_14275,N_14438);
or UO_320 (O_320,N_14573,N_14915);
and UO_321 (O_321,N_14768,N_14096);
or UO_322 (O_322,N_14674,N_14660);
nand UO_323 (O_323,N_14961,N_14544);
or UO_324 (O_324,N_14254,N_14091);
and UO_325 (O_325,N_14619,N_14002);
xnor UO_326 (O_326,N_14316,N_14173);
or UO_327 (O_327,N_14421,N_14762);
xor UO_328 (O_328,N_14423,N_14635);
and UO_329 (O_329,N_14080,N_14152);
or UO_330 (O_330,N_14377,N_14788);
and UO_331 (O_331,N_14798,N_14290);
and UO_332 (O_332,N_14371,N_14226);
nor UO_333 (O_333,N_14505,N_14385);
or UO_334 (O_334,N_14881,N_14116);
nor UO_335 (O_335,N_14481,N_14007);
or UO_336 (O_336,N_14113,N_14295);
nor UO_337 (O_337,N_14475,N_14547);
and UO_338 (O_338,N_14867,N_14634);
or UO_339 (O_339,N_14261,N_14655);
and UO_340 (O_340,N_14678,N_14691);
and UO_341 (O_341,N_14405,N_14389);
xor UO_342 (O_342,N_14695,N_14010);
nor UO_343 (O_343,N_14102,N_14518);
nor UO_344 (O_344,N_14192,N_14855);
nor UO_345 (O_345,N_14196,N_14351);
nor UO_346 (O_346,N_14702,N_14120);
nand UO_347 (O_347,N_14178,N_14976);
xnor UO_348 (O_348,N_14746,N_14554);
xor UO_349 (O_349,N_14597,N_14082);
nand UO_350 (O_350,N_14023,N_14057);
or UO_351 (O_351,N_14797,N_14187);
or UO_352 (O_352,N_14998,N_14289);
nor UO_353 (O_353,N_14374,N_14500);
xor UO_354 (O_354,N_14838,N_14562);
nor UO_355 (O_355,N_14392,N_14612);
xor UO_356 (O_356,N_14928,N_14770);
nor UO_357 (O_357,N_14793,N_14799);
or UO_358 (O_358,N_14566,N_14993);
xor UO_359 (O_359,N_14668,N_14231);
or UO_360 (O_360,N_14866,N_14135);
nand UO_361 (O_361,N_14414,N_14279);
nand UO_362 (O_362,N_14156,N_14394);
xnor UO_363 (O_363,N_14000,N_14367);
xor UO_364 (O_364,N_14730,N_14752);
or UO_365 (O_365,N_14959,N_14508);
or UO_366 (O_366,N_14227,N_14713);
xnor UO_367 (O_367,N_14711,N_14197);
or UO_368 (O_368,N_14072,N_14462);
xor UO_369 (O_369,N_14436,N_14885);
and UO_370 (O_370,N_14207,N_14877);
or UO_371 (O_371,N_14210,N_14524);
and UO_372 (O_372,N_14550,N_14672);
nand UO_373 (O_373,N_14246,N_14448);
nor UO_374 (O_374,N_14509,N_14172);
and UO_375 (O_375,N_14977,N_14844);
xor UO_376 (O_376,N_14186,N_14780);
and UO_377 (O_377,N_14593,N_14541);
nand UO_378 (O_378,N_14427,N_14115);
nor UO_379 (O_379,N_14278,N_14440);
or UO_380 (O_380,N_14122,N_14621);
and UO_381 (O_381,N_14398,N_14686);
or UO_382 (O_382,N_14287,N_14643);
or UO_383 (O_383,N_14724,N_14632);
xor UO_384 (O_384,N_14590,N_14907);
and UO_385 (O_385,N_14822,N_14077);
nand UO_386 (O_386,N_14484,N_14494);
xnor UO_387 (O_387,N_14179,N_14066);
xor UO_388 (O_388,N_14572,N_14857);
nor UO_389 (O_389,N_14882,N_14063);
or UO_390 (O_390,N_14941,N_14542);
and UO_391 (O_391,N_14412,N_14898);
and UO_392 (O_392,N_14983,N_14491);
nand UO_393 (O_393,N_14240,N_14944);
nor UO_394 (O_394,N_14264,N_14764);
and UO_395 (O_395,N_14498,N_14705);
and UO_396 (O_396,N_14402,N_14601);
and UO_397 (O_397,N_14872,N_14503);
nand UO_398 (O_398,N_14107,N_14390);
nor UO_399 (O_399,N_14118,N_14978);
nand UO_400 (O_400,N_14592,N_14721);
and UO_401 (O_401,N_14033,N_14611);
nand UO_402 (O_402,N_14038,N_14482);
or UO_403 (O_403,N_14666,N_14041);
nor UO_404 (O_404,N_14366,N_14047);
nor UO_405 (O_405,N_14681,N_14504);
and UO_406 (O_406,N_14459,N_14870);
xnor UO_407 (O_407,N_14758,N_14754);
nand UO_408 (O_408,N_14725,N_14849);
and UO_409 (O_409,N_14296,N_14880);
xor UO_410 (O_410,N_14065,N_14653);
nand UO_411 (O_411,N_14536,N_14520);
or UO_412 (O_412,N_14164,N_14090);
or UO_413 (O_413,N_14916,N_14757);
xnor UO_414 (O_414,N_14677,N_14765);
or UO_415 (O_415,N_14889,N_14444);
or UO_416 (O_416,N_14930,N_14812);
and UO_417 (O_417,N_14840,N_14836);
or UO_418 (O_418,N_14802,N_14557);
and UO_419 (O_419,N_14847,N_14147);
or UO_420 (O_420,N_14832,N_14457);
nor UO_421 (O_421,N_14449,N_14242);
nor UO_422 (O_422,N_14028,N_14815);
nor UO_423 (O_423,N_14924,N_14194);
xor UO_424 (O_424,N_14750,N_14884);
and UO_425 (O_425,N_14003,N_14627);
and UO_426 (O_426,N_14614,N_14249);
xnor UO_427 (O_427,N_14912,N_14467);
or UO_428 (O_428,N_14382,N_14051);
nand UO_429 (O_429,N_14971,N_14074);
nand UO_430 (O_430,N_14235,N_14943);
nor UO_431 (O_431,N_14527,N_14154);
nand UO_432 (O_432,N_14229,N_14514);
xor UO_433 (O_433,N_14526,N_14381);
and UO_434 (O_434,N_14905,N_14285);
nor UO_435 (O_435,N_14338,N_14919);
xor UO_436 (O_436,N_14183,N_14913);
xnor UO_437 (O_437,N_14373,N_14664);
nand UO_438 (O_438,N_14631,N_14403);
nor UO_439 (O_439,N_14011,N_14121);
nand UO_440 (O_440,N_14166,N_14726);
xor UO_441 (O_441,N_14391,N_14727);
or UO_442 (O_442,N_14326,N_14071);
and UO_443 (O_443,N_14248,N_14306);
and UO_444 (O_444,N_14970,N_14845);
and UO_445 (O_445,N_14651,N_14582);
or UO_446 (O_446,N_14957,N_14200);
or UO_447 (O_447,N_14488,N_14418);
and UO_448 (O_448,N_14148,N_14114);
or UO_449 (O_449,N_14661,N_14157);
xor UO_450 (O_450,N_14931,N_14637);
or UO_451 (O_451,N_14145,N_14088);
xnor UO_452 (O_452,N_14599,N_14753);
nor UO_453 (O_453,N_14104,N_14737);
and UO_454 (O_454,N_14615,N_14563);
nor UO_455 (O_455,N_14906,N_14694);
nor UO_456 (O_456,N_14170,N_14749);
nor UO_457 (O_457,N_14774,N_14451);
and UO_458 (O_458,N_14211,N_14035);
or UO_459 (O_459,N_14100,N_14560);
and UO_460 (O_460,N_14570,N_14206);
nor UO_461 (O_461,N_14502,N_14218);
and UO_462 (O_462,N_14969,N_14623);
xnor UO_463 (O_463,N_14785,N_14092);
and UO_464 (O_464,N_14317,N_14876);
nor UO_465 (O_465,N_14982,N_14784);
nor UO_466 (O_466,N_14938,N_14485);
xor UO_467 (O_467,N_14299,N_14837);
xor UO_468 (O_468,N_14247,N_14565);
xor UO_469 (O_469,N_14511,N_14613);
xor UO_470 (O_470,N_14225,N_14859);
nand UO_471 (O_471,N_14578,N_14608);
nor UO_472 (O_472,N_14129,N_14030);
nand UO_473 (O_473,N_14331,N_14988);
and UO_474 (O_474,N_14980,N_14521);
nand UO_475 (O_475,N_14658,N_14652);
nand UO_476 (O_476,N_14680,N_14258);
and UO_477 (O_477,N_14434,N_14540);
xor UO_478 (O_478,N_14452,N_14013);
nand UO_479 (O_479,N_14945,N_14040);
xnor UO_480 (O_480,N_14733,N_14219);
or UO_481 (O_481,N_14546,N_14696);
xor UO_482 (O_482,N_14588,N_14125);
and UO_483 (O_483,N_14648,N_14396);
nor UO_484 (O_484,N_14537,N_14388);
xor UO_485 (O_485,N_14087,N_14042);
xnor UO_486 (O_486,N_14205,N_14618);
nand UO_487 (O_487,N_14169,N_14282);
and UO_488 (O_488,N_14908,N_14759);
xnor UO_489 (O_489,N_14555,N_14602);
nand UO_490 (O_490,N_14501,N_14016);
nor UO_491 (O_491,N_14262,N_14704);
nand UO_492 (O_492,N_14244,N_14301);
or UO_493 (O_493,N_14703,N_14465);
nor UO_494 (O_494,N_14600,N_14463);
xnor UO_495 (O_495,N_14056,N_14820);
xnor UO_496 (O_496,N_14790,N_14786);
or UO_497 (O_497,N_14193,N_14165);
nand UO_498 (O_498,N_14937,N_14507);
and UO_499 (O_499,N_14214,N_14807);
and UO_500 (O_500,N_14223,N_14793);
or UO_501 (O_501,N_14231,N_14576);
nand UO_502 (O_502,N_14940,N_14333);
nor UO_503 (O_503,N_14776,N_14751);
and UO_504 (O_504,N_14456,N_14292);
xor UO_505 (O_505,N_14198,N_14575);
xnor UO_506 (O_506,N_14914,N_14863);
and UO_507 (O_507,N_14833,N_14187);
or UO_508 (O_508,N_14873,N_14936);
xnor UO_509 (O_509,N_14127,N_14211);
and UO_510 (O_510,N_14995,N_14878);
xnor UO_511 (O_511,N_14056,N_14265);
or UO_512 (O_512,N_14639,N_14466);
or UO_513 (O_513,N_14360,N_14691);
nand UO_514 (O_514,N_14047,N_14169);
nor UO_515 (O_515,N_14787,N_14173);
xnor UO_516 (O_516,N_14593,N_14904);
nor UO_517 (O_517,N_14395,N_14625);
nand UO_518 (O_518,N_14534,N_14401);
nor UO_519 (O_519,N_14253,N_14250);
nand UO_520 (O_520,N_14609,N_14555);
and UO_521 (O_521,N_14231,N_14800);
xnor UO_522 (O_522,N_14315,N_14187);
xor UO_523 (O_523,N_14576,N_14934);
nor UO_524 (O_524,N_14887,N_14285);
nand UO_525 (O_525,N_14673,N_14150);
nor UO_526 (O_526,N_14739,N_14758);
nand UO_527 (O_527,N_14986,N_14784);
and UO_528 (O_528,N_14178,N_14850);
nor UO_529 (O_529,N_14806,N_14813);
xor UO_530 (O_530,N_14420,N_14774);
or UO_531 (O_531,N_14631,N_14796);
nor UO_532 (O_532,N_14950,N_14022);
nand UO_533 (O_533,N_14533,N_14865);
nor UO_534 (O_534,N_14690,N_14420);
nand UO_535 (O_535,N_14343,N_14483);
or UO_536 (O_536,N_14946,N_14790);
nor UO_537 (O_537,N_14192,N_14195);
nor UO_538 (O_538,N_14618,N_14520);
nand UO_539 (O_539,N_14519,N_14776);
nand UO_540 (O_540,N_14043,N_14144);
nand UO_541 (O_541,N_14068,N_14704);
nor UO_542 (O_542,N_14996,N_14413);
xor UO_543 (O_543,N_14432,N_14070);
or UO_544 (O_544,N_14921,N_14212);
nand UO_545 (O_545,N_14625,N_14064);
xnor UO_546 (O_546,N_14390,N_14848);
and UO_547 (O_547,N_14396,N_14855);
and UO_548 (O_548,N_14430,N_14665);
xnor UO_549 (O_549,N_14672,N_14129);
nand UO_550 (O_550,N_14844,N_14593);
nand UO_551 (O_551,N_14895,N_14401);
or UO_552 (O_552,N_14455,N_14162);
nand UO_553 (O_553,N_14085,N_14793);
nor UO_554 (O_554,N_14060,N_14337);
nand UO_555 (O_555,N_14677,N_14474);
xor UO_556 (O_556,N_14087,N_14444);
nor UO_557 (O_557,N_14732,N_14008);
nand UO_558 (O_558,N_14810,N_14528);
nand UO_559 (O_559,N_14830,N_14828);
and UO_560 (O_560,N_14780,N_14907);
or UO_561 (O_561,N_14976,N_14880);
or UO_562 (O_562,N_14790,N_14168);
xor UO_563 (O_563,N_14860,N_14431);
and UO_564 (O_564,N_14223,N_14908);
or UO_565 (O_565,N_14301,N_14877);
and UO_566 (O_566,N_14799,N_14603);
or UO_567 (O_567,N_14452,N_14482);
and UO_568 (O_568,N_14101,N_14748);
nor UO_569 (O_569,N_14750,N_14758);
nor UO_570 (O_570,N_14396,N_14977);
and UO_571 (O_571,N_14798,N_14591);
nand UO_572 (O_572,N_14800,N_14509);
nand UO_573 (O_573,N_14604,N_14573);
nor UO_574 (O_574,N_14326,N_14875);
or UO_575 (O_575,N_14040,N_14777);
and UO_576 (O_576,N_14068,N_14538);
and UO_577 (O_577,N_14939,N_14072);
or UO_578 (O_578,N_14095,N_14622);
nor UO_579 (O_579,N_14148,N_14071);
nor UO_580 (O_580,N_14338,N_14818);
nor UO_581 (O_581,N_14869,N_14380);
xnor UO_582 (O_582,N_14616,N_14344);
nand UO_583 (O_583,N_14751,N_14836);
nand UO_584 (O_584,N_14494,N_14193);
or UO_585 (O_585,N_14007,N_14158);
xnor UO_586 (O_586,N_14490,N_14626);
nor UO_587 (O_587,N_14110,N_14579);
nand UO_588 (O_588,N_14477,N_14432);
nor UO_589 (O_589,N_14580,N_14419);
or UO_590 (O_590,N_14610,N_14090);
nor UO_591 (O_591,N_14175,N_14474);
nor UO_592 (O_592,N_14117,N_14014);
nor UO_593 (O_593,N_14808,N_14716);
xor UO_594 (O_594,N_14954,N_14930);
nand UO_595 (O_595,N_14046,N_14327);
and UO_596 (O_596,N_14361,N_14451);
xnor UO_597 (O_597,N_14500,N_14513);
or UO_598 (O_598,N_14006,N_14106);
or UO_599 (O_599,N_14444,N_14484);
or UO_600 (O_600,N_14696,N_14298);
or UO_601 (O_601,N_14678,N_14115);
nor UO_602 (O_602,N_14148,N_14665);
nand UO_603 (O_603,N_14860,N_14766);
nand UO_604 (O_604,N_14503,N_14722);
or UO_605 (O_605,N_14523,N_14253);
nand UO_606 (O_606,N_14087,N_14620);
xnor UO_607 (O_607,N_14231,N_14947);
nor UO_608 (O_608,N_14112,N_14978);
nor UO_609 (O_609,N_14128,N_14061);
nor UO_610 (O_610,N_14583,N_14164);
nand UO_611 (O_611,N_14686,N_14783);
or UO_612 (O_612,N_14108,N_14953);
xnor UO_613 (O_613,N_14178,N_14712);
xor UO_614 (O_614,N_14299,N_14365);
nand UO_615 (O_615,N_14539,N_14559);
nand UO_616 (O_616,N_14888,N_14225);
and UO_617 (O_617,N_14502,N_14340);
nor UO_618 (O_618,N_14907,N_14970);
or UO_619 (O_619,N_14963,N_14232);
and UO_620 (O_620,N_14965,N_14559);
nor UO_621 (O_621,N_14295,N_14375);
or UO_622 (O_622,N_14636,N_14604);
nand UO_623 (O_623,N_14707,N_14355);
or UO_624 (O_624,N_14545,N_14394);
xnor UO_625 (O_625,N_14142,N_14761);
nor UO_626 (O_626,N_14193,N_14613);
and UO_627 (O_627,N_14403,N_14064);
nand UO_628 (O_628,N_14323,N_14365);
or UO_629 (O_629,N_14784,N_14234);
nor UO_630 (O_630,N_14240,N_14185);
and UO_631 (O_631,N_14595,N_14988);
nor UO_632 (O_632,N_14641,N_14934);
and UO_633 (O_633,N_14596,N_14100);
nand UO_634 (O_634,N_14210,N_14909);
nand UO_635 (O_635,N_14279,N_14893);
or UO_636 (O_636,N_14014,N_14164);
nand UO_637 (O_637,N_14734,N_14719);
nor UO_638 (O_638,N_14289,N_14623);
xnor UO_639 (O_639,N_14411,N_14973);
nand UO_640 (O_640,N_14187,N_14611);
and UO_641 (O_641,N_14903,N_14911);
or UO_642 (O_642,N_14271,N_14138);
xnor UO_643 (O_643,N_14042,N_14835);
xnor UO_644 (O_644,N_14013,N_14098);
nor UO_645 (O_645,N_14572,N_14350);
and UO_646 (O_646,N_14309,N_14867);
xnor UO_647 (O_647,N_14298,N_14744);
xnor UO_648 (O_648,N_14835,N_14365);
or UO_649 (O_649,N_14754,N_14082);
nor UO_650 (O_650,N_14538,N_14122);
nand UO_651 (O_651,N_14457,N_14799);
or UO_652 (O_652,N_14987,N_14760);
and UO_653 (O_653,N_14769,N_14715);
nand UO_654 (O_654,N_14454,N_14424);
nand UO_655 (O_655,N_14992,N_14470);
or UO_656 (O_656,N_14963,N_14892);
nor UO_657 (O_657,N_14469,N_14533);
nand UO_658 (O_658,N_14469,N_14773);
nor UO_659 (O_659,N_14906,N_14992);
or UO_660 (O_660,N_14052,N_14443);
or UO_661 (O_661,N_14317,N_14336);
xor UO_662 (O_662,N_14416,N_14340);
and UO_663 (O_663,N_14426,N_14580);
and UO_664 (O_664,N_14804,N_14426);
nand UO_665 (O_665,N_14670,N_14009);
nor UO_666 (O_666,N_14358,N_14213);
xor UO_667 (O_667,N_14816,N_14754);
nand UO_668 (O_668,N_14811,N_14617);
xnor UO_669 (O_669,N_14757,N_14612);
xor UO_670 (O_670,N_14364,N_14899);
and UO_671 (O_671,N_14156,N_14845);
and UO_672 (O_672,N_14352,N_14177);
or UO_673 (O_673,N_14110,N_14312);
and UO_674 (O_674,N_14367,N_14621);
and UO_675 (O_675,N_14438,N_14648);
nand UO_676 (O_676,N_14653,N_14736);
or UO_677 (O_677,N_14913,N_14794);
xor UO_678 (O_678,N_14236,N_14986);
or UO_679 (O_679,N_14771,N_14527);
nand UO_680 (O_680,N_14345,N_14419);
or UO_681 (O_681,N_14026,N_14033);
nand UO_682 (O_682,N_14990,N_14004);
xor UO_683 (O_683,N_14053,N_14844);
nor UO_684 (O_684,N_14738,N_14214);
nand UO_685 (O_685,N_14000,N_14832);
or UO_686 (O_686,N_14139,N_14680);
xnor UO_687 (O_687,N_14608,N_14205);
nor UO_688 (O_688,N_14367,N_14343);
and UO_689 (O_689,N_14326,N_14363);
or UO_690 (O_690,N_14509,N_14803);
or UO_691 (O_691,N_14020,N_14496);
xor UO_692 (O_692,N_14466,N_14061);
xnor UO_693 (O_693,N_14640,N_14530);
or UO_694 (O_694,N_14760,N_14166);
nand UO_695 (O_695,N_14682,N_14688);
or UO_696 (O_696,N_14045,N_14421);
nand UO_697 (O_697,N_14233,N_14503);
nor UO_698 (O_698,N_14734,N_14980);
nand UO_699 (O_699,N_14139,N_14041);
or UO_700 (O_700,N_14708,N_14966);
nand UO_701 (O_701,N_14815,N_14730);
xnor UO_702 (O_702,N_14544,N_14561);
and UO_703 (O_703,N_14316,N_14806);
xor UO_704 (O_704,N_14781,N_14801);
and UO_705 (O_705,N_14346,N_14970);
or UO_706 (O_706,N_14503,N_14797);
and UO_707 (O_707,N_14157,N_14748);
nor UO_708 (O_708,N_14354,N_14735);
nand UO_709 (O_709,N_14906,N_14343);
and UO_710 (O_710,N_14891,N_14259);
xnor UO_711 (O_711,N_14963,N_14986);
nand UO_712 (O_712,N_14480,N_14035);
nor UO_713 (O_713,N_14825,N_14008);
and UO_714 (O_714,N_14995,N_14740);
nand UO_715 (O_715,N_14295,N_14276);
nor UO_716 (O_716,N_14591,N_14250);
nand UO_717 (O_717,N_14181,N_14381);
nand UO_718 (O_718,N_14295,N_14081);
and UO_719 (O_719,N_14295,N_14142);
nor UO_720 (O_720,N_14927,N_14011);
and UO_721 (O_721,N_14357,N_14316);
nand UO_722 (O_722,N_14338,N_14775);
nand UO_723 (O_723,N_14604,N_14596);
xnor UO_724 (O_724,N_14349,N_14721);
nand UO_725 (O_725,N_14952,N_14070);
and UO_726 (O_726,N_14605,N_14232);
xor UO_727 (O_727,N_14073,N_14650);
and UO_728 (O_728,N_14937,N_14150);
nand UO_729 (O_729,N_14517,N_14564);
nor UO_730 (O_730,N_14877,N_14385);
xor UO_731 (O_731,N_14395,N_14601);
and UO_732 (O_732,N_14269,N_14938);
xor UO_733 (O_733,N_14388,N_14795);
or UO_734 (O_734,N_14050,N_14357);
and UO_735 (O_735,N_14920,N_14643);
nand UO_736 (O_736,N_14412,N_14229);
and UO_737 (O_737,N_14622,N_14882);
xnor UO_738 (O_738,N_14546,N_14222);
xor UO_739 (O_739,N_14285,N_14720);
nor UO_740 (O_740,N_14958,N_14161);
or UO_741 (O_741,N_14161,N_14951);
or UO_742 (O_742,N_14438,N_14622);
xnor UO_743 (O_743,N_14821,N_14793);
and UO_744 (O_744,N_14447,N_14717);
nand UO_745 (O_745,N_14256,N_14066);
nand UO_746 (O_746,N_14725,N_14925);
and UO_747 (O_747,N_14429,N_14952);
xnor UO_748 (O_748,N_14153,N_14315);
or UO_749 (O_749,N_14648,N_14499);
xnor UO_750 (O_750,N_14663,N_14715);
nand UO_751 (O_751,N_14226,N_14603);
or UO_752 (O_752,N_14339,N_14053);
and UO_753 (O_753,N_14026,N_14637);
nor UO_754 (O_754,N_14161,N_14835);
xnor UO_755 (O_755,N_14559,N_14932);
xnor UO_756 (O_756,N_14362,N_14855);
nand UO_757 (O_757,N_14003,N_14712);
or UO_758 (O_758,N_14770,N_14844);
and UO_759 (O_759,N_14392,N_14285);
and UO_760 (O_760,N_14881,N_14683);
nor UO_761 (O_761,N_14688,N_14686);
or UO_762 (O_762,N_14297,N_14061);
and UO_763 (O_763,N_14631,N_14513);
xnor UO_764 (O_764,N_14154,N_14687);
and UO_765 (O_765,N_14608,N_14006);
nor UO_766 (O_766,N_14483,N_14897);
nor UO_767 (O_767,N_14296,N_14722);
xnor UO_768 (O_768,N_14237,N_14698);
nand UO_769 (O_769,N_14426,N_14197);
and UO_770 (O_770,N_14214,N_14350);
or UO_771 (O_771,N_14190,N_14835);
or UO_772 (O_772,N_14136,N_14300);
and UO_773 (O_773,N_14880,N_14451);
or UO_774 (O_774,N_14088,N_14826);
nand UO_775 (O_775,N_14133,N_14712);
nor UO_776 (O_776,N_14672,N_14468);
xor UO_777 (O_777,N_14217,N_14396);
and UO_778 (O_778,N_14304,N_14666);
and UO_779 (O_779,N_14450,N_14133);
xor UO_780 (O_780,N_14655,N_14078);
nand UO_781 (O_781,N_14461,N_14154);
nand UO_782 (O_782,N_14765,N_14042);
nand UO_783 (O_783,N_14587,N_14039);
xor UO_784 (O_784,N_14745,N_14498);
nand UO_785 (O_785,N_14659,N_14579);
and UO_786 (O_786,N_14679,N_14187);
xnor UO_787 (O_787,N_14130,N_14977);
or UO_788 (O_788,N_14342,N_14175);
nand UO_789 (O_789,N_14851,N_14691);
nand UO_790 (O_790,N_14466,N_14710);
xor UO_791 (O_791,N_14548,N_14300);
xnor UO_792 (O_792,N_14290,N_14113);
nand UO_793 (O_793,N_14252,N_14311);
nor UO_794 (O_794,N_14620,N_14991);
xor UO_795 (O_795,N_14290,N_14446);
and UO_796 (O_796,N_14346,N_14080);
xnor UO_797 (O_797,N_14635,N_14788);
nor UO_798 (O_798,N_14755,N_14504);
xor UO_799 (O_799,N_14015,N_14120);
and UO_800 (O_800,N_14809,N_14479);
nor UO_801 (O_801,N_14531,N_14743);
nand UO_802 (O_802,N_14683,N_14307);
and UO_803 (O_803,N_14230,N_14343);
nand UO_804 (O_804,N_14370,N_14778);
and UO_805 (O_805,N_14200,N_14786);
nor UO_806 (O_806,N_14022,N_14223);
nand UO_807 (O_807,N_14951,N_14330);
nand UO_808 (O_808,N_14330,N_14980);
xnor UO_809 (O_809,N_14112,N_14359);
nor UO_810 (O_810,N_14177,N_14532);
or UO_811 (O_811,N_14583,N_14602);
xor UO_812 (O_812,N_14971,N_14927);
nor UO_813 (O_813,N_14214,N_14024);
or UO_814 (O_814,N_14616,N_14653);
nand UO_815 (O_815,N_14514,N_14324);
nand UO_816 (O_816,N_14756,N_14033);
nand UO_817 (O_817,N_14461,N_14707);
and UO_818 (O_818,N_14152,N_14677);
and UO_819 (O_819,N_14468,N_14493);
or UO_820 (O_820,N_14865,N_14762);
and UO_821 (O_821,N_14362,N_14314);
xor UO_822 (O_822,N_14195,N_14605);
nor UO_823 (O_823,N_14652,N_14601);
xor UO_824 (O_824,N_14390,N_14809);
xor UO_825 (O_825,N_14991,N_14229);
and UO_826 (O_826,N_14722,N_14111);
xnor UO_827 (O_827,N_14248,N_14020);
or UO_828 (O_828,N_14640,N_14186);
nor UO_829 (O_829,N_14528,N_14158);
nand UO_830 (O_830,N_14221,N_14805);
or UO_831 (O_831,N_14013,N_14315);
xor UO_832 (O_832,N_14684,N_14217);
nor UO_833 (O_833,N_14188,N_14426);
and UO_834 (O_834,N_14613,N_14261);
nand UO_835 (O_835,N_14636,N_14252);
xnor UO_836 (O_836,N_14370,N_14697);
and UO_837 (O_837,N_14044,N_14656);
xor UO_838 (O_838,N_14706,N_14204);
xnor UO_839 (O_839,N_14231,N_14295);
nor UO_840 (O_840,N_14839,N_14880);
nand UO_841 (O_841,N_14331,N_14801);
nand UO_842 (O_842,N_14232,N_14175);
xor UO_843 (O_843,N_14662,N_14786);
nor UO_844 (O_844,N_14869,N_14272);
and UO_845 (O_845,N_14122,N_14956);
or UO_846 (O_846,N_14255,N_14349);
xor UO_847 (O_847,N_14580,N_14872);
nor UO_848 (O_848,N_14185,N_14862);
nor UO_849 (O_849,N_14950,N_14252);
nor UO_850 (O_850,N_14860,N_14522);
or UO_851 (O_851,N_14630,N_14506);
xor UO_852 (O_852,N_14715,N_14196);
nor UO_853 (O_853,N_14970,N_14424);
nand UO_854 (O_854,N_14272,N_14716);
nand UO_855 (O_855,N_14558,N_14287);
or UO_856 (O_856,N_14390,N_14617);
nor UO_857 (O_857,N_14971,N_14401);
or UO_858 (O_858,N_14717,N_14932);
or UO_859 (O_859,N_14855,N_14068);
nor UO_860 (O_860,N_14171,N_14973);
or UO_861 (O_861,N_14459,N_14036);
nand UO_862 (O_862,N_14688,N_14855);
nor UO_863 (O_863,N_14428,N_14929);
or UO_864 (O_864,N_14526,N_14365);
nand UO_865 (O_865,N_14470,N_14286);
xor UO_866 (O_866,N_14450,N_14417);
xor UO_867 (O_867,N_14704,N_14434);
or UO_868 (O_868,N_14986,N_14216);
xor UO_869 (O_869,N_14883,N_14115);
and UO_870 (O_870,N_14348,N_14865);
xnor UO_871 (O_871,N_14116,N_14509);
and UO_872 (O_872,N_14181,N_14697);
nor UO_873 (O_873,N_14893,N_14866);
nor UO_874 (O_874,N_14169,N_14170);
nand UO_875 (O_875,N_14720,N_14183);
xnor UO_876 (O_876,N_14418,N_14043);
nand UO_877 (O_877,N_14304,N_14943);
nor UO_878 (O_878,N_14026,N_14214);
and UO_879 (O_879,N_14880,N_14223);
and UO_880 (O_880,N_14159,N_14258);
nor UO_881 (O_881,N_14692,N_14489);
and UO_882 (O_882,N_14045,N_14408);
and UO_883 (O_883,N_14930,N_14276);
nor UO_884 (O_884,N_14387,N_14533);
and UO_885 (O_885,N_14302,N_14307);
and UO_886 (O_886,N_14570,N_14280);
or UO_887 (O_887,N_14332,N_14499);
xor UO_888 (O_888,N_14293,N_14050);
xnor UO_889 (O_889,N_14651,N_14969);
xnor UO_890 (O_890,N_14395,N_14877);
and UO_891 (O_891,N_14279,N_14485);
xnor UO_892 (O_892,N_14815,N_14252);
nand UO_893 (O_893,N_14041,N_14910);
nor UO_894 (O_894,N_14404,N_14897);
xor UO_895 (O_895,N_14539,N_14179);
or UO_896 (O_896,N_14007,N_14341);
nand UO_897 (O_897,N_14297,N_14175);
or UO_898 (O_898,N_14021,N_14051);
nand UO_899 (O_899,N_14451,N_14546);
nand UO_900 (O_900,N_14607,N_14588);
nor UO_901 (O_901,N_14583,N_14502);
nor UO_902 (O_902,N_14664,N_14285);
nand UO_903 (O_903,N_14168,N_14123);
nand UO_904 (O_904,N_14512,N_14383);
and UO_905 (O_905,N_14572,N_14822);
xnor UO_906 (O_906,N_14090,N_14993);
and UO_907 (O_907,N_14924,N_14215);
xor UO_908 (O_908,N_14774,N_14781);
or UO_909 (O_909,N_14429,N_14094);
nor UO_910 (O_910,N_14901,N_14788);
nor UO_911 (O_911,N_14929,N_14414);
xnor UO_912 (O_912,N_14110,N_14170);
and UO_913 (O_913,N_14444,N_14703);
nor UO_914 (O_914,N_14321,N_14565);
nor UO_915 (O_915,N_14332,N_14414);
and UO_916 (O_916,N_14474,N_14236);
or UO_917 (O_917,N_14968,N_14287);
nor UO_918 (O_918,N_14488,N_14842);
or UO_919 (O_919,N_14520,N_14924);
xnor UO_920 (O_920,N_14418,N_14022);
nand UO_921 (O_921,N_14965,N_14479);
or UO_922 (O_922,N_14074,N_14228);
nor UO_923 (O_923,N_14317,N_14207);
xnor UO_924 (O_924,N_14806,N_14523);
nand UO_925 (O_925,N_14522,N_14083);
nand UO_926 (O_926,N_14398,N_14084);
nor UO_927 (O_927,N_14763,N_14188);
and UO_928 (O_928,N_14864,N_14207);
nand UO_929 (O_929,N_14638,N_14944);
and UO_930 (O_930,N_14585,N_14157);
xnor UO_931 (O_931,N_14094,N_14184);
nand UO_932 (O_932,N_14999,N_14704);
or UO_933 (O_933,N_14922,N_14021);
xnor UO_934 (O_934,N_14426,N_14091);
and UO_935 (O_935,N_14987,N_14578);
nor UO_936 (O_936,N_14632,N_14134);
nor UO_937 (O_937,N_14841,N_14547);
and UO_938 (O_938,N_14420,N_14419);
or UO_939 (O_939,N_14064,N_14534);
and UO_940 (O_940,N_14398,N_14143);
nand UO_941 (O_941,N_14986,N_14763);
and UO_942 (O_942,N_14218,N_14550);
and UO_943 (O_943,N_14367,N_14552);
nand UO_944 (O_944,N_14965,N_14180);
xor UO_945 (O_945,N_14252,N_14427);
and UO_946 (O_946,N_14311,N_14423);
and UO_947 (O_947,N_14502,N_14796);
nor UO_948 (O_948,N_14476,N_14134);
nor UO_949 (O_949,N_14311,N_14022);
or UO_950 (O_950,N_14283,N_14702);
xor UO_951 (O_951,N_14104,N_14173);
and UO_952 (O_952,N_14657,N_14914);
xor UO_953 (O_953,N_14943,N_14818);
nor UO_954 (O_954,N_14325,N_14158);
and UO_955 (O_955,N_14169,N_14237);
xor UO_956 (O_956,N_14795,N_14719);
xor UO_957 (O_957,N_14506,N_14619);
or UO_958 (O_958,N_14559,N_14631);
nor UO_959 (O_959,N_14221,N_14612);
xor UO_960 (O_960,N_14960,N_14121);
nand UO_961 (O_961,N_14682,N_14555);
xnor UO_962 (O_962,N_14602,N_14404);
xor UO_963 (O_963,N_14740,N_14149);
xnor UO_964 (O_964,N_14898,N_14029);
nand UO_965 (O_965,N_14390,N_14616);
xor UO_966 (O_966,N_14097,N_14832);
nand UO_967 (O_967,N_14941,N_14594);
nor UO_968 (O_968,N_14208,N_14584);
or UO_969 (O_969,N_14430,N_14408);
nand UO_970 (O_970,N_14259,N_14161);
nand UO_971 (O_971,N_14967,N_14814);
nand UO_972 (O_972,N_14167,N_14499);
xor UO_973 (O_973,N_14848,N_14701);
nand UO_974 (O_974,N_14913,N_14637);
nand UO_975 (O_975,N_14673,N_14301);
nor UO_976 (O_976,N_14944,N_14800);
xor UO_977 (O_977,N_14817,N_14256);
xnor UO_978 (O_978,N_14989,N_14513);
or UO_979 (O_979,N_14955,N_14075);
and UO_980 (O_980,N_14285,N_14524);
and UO_981 (O_981,N_14764,N_14488);
xnor UO_982 (O_982,N_14085,N_14175);
and UO_983 (O_983,N_14321,N_14880);
and UO_984 (O_984,N_14948,N_14204);
nand UO_985 (O_985,N_14665,N_14137);
or UO_986 (O_986,N_14562,N_14887);
and UO_987 (O_987,N_14736,N_14402);
nor UO_988 (O_988,N_14270,N_14751);
or UO_989 (O_989,N_14533,N_14402);
nand UO_990 (O_990,N_14455,N_14219);
or UO_991 (O_991,N_14739,N_14043);
xnor UO_992 (O_992,N_14926,N_14243);
and UO_993 (O_993,N_14487,N_14240);
xnor UO_994 (O_994,N_14919,N_14678);
nor UO_995 (O_995,N_14058,N_14254);
or UO_996 (O_996,N_14959,N_14810);
nor UO_997 (O_997,N_14983,N_14678);
and UO_998 (O_998,N_14166,N_14470);
and UO_999 (O_999,N_14755,N_14431);
nand UO_1000 (O_1000,N_14626,N_14183);
nor UO_1001 (O_1001,N_14132,N_14684);
or UO_1002 (O_1002,N_14658,N_14044);
nor UO_1003 (O_1003,N_14182,N_14332);
nor UO_1004 (O_1004,N_14867,N_14545);
and UO_1005 (O_1005,N_14973,N_14624);
nor UO_1006 (O_1006,N_14280,N_14674);
nand UO_1007 (O_1007,N_14805,N_14617);
and UO_1008 (O_1008,N_14350,N_14224);
xnor UO_1009 (O_1009,N_14051,N_14365);
or UO_1010 (O_1010,N_14691,N_14363);
nand UO_1011 (O_1011,N_14769,N_14815);
nand UO_1012 (O_1012,N_14398,N_14678);
and UO_1013 (O_1013,N_14307,N_14754);
nand UO_1014 (O_1014,N_14311,N_14597);
nand UO_1015 (O_1015,N_14447,N_14399);
nand UO_1016 (O_1016,N_14404,N_14015);
and UO_1017 (O_1017,N_14302,N_14599);
and UO_1018 (O_1018,N_14130,N_14443);
xor UO_1019 (O_1019,N_14741,N_14894);
nand UO_1020 (O_1020,N_14656,N_14156);
and UO_1021 (O_1021,N_14718,N_14316);
nand UO_1022 (O_1022,N_14236,N_14083);
xor UO_1023 (O_1023,N_14462,N_14329);
xor UO_1024 (O_1024,N_14205,N_14634);
or UO_1025 (O_1025,N_14626,N_14048);
xor UO_1026 (O_1026,N_14285,N_14025);
nand UO_1027 (O_1027,N_14389,N_14268);
and UO_1028 (O_1028,N_14668,N_14767);
nand UO_1029 (O_1029,N_14981,N_14587);
nor UO_1030 (O_1030,N_14827,N_14875);
and UO_1031 (O_1031,N_14019,N_14803);
or UO_1032 (O_1032,N_14934,N_14818);
xor UO_1033 (O_1033,N_14966,N_14717);
xnor UO_1034 (O_1034,N_14078,N_14981);
nor UO_1035 (O_1035,N_14070,N_14180);
or UO_1036 (O_1036,N_14730,N_14957);
and UO_1037 (O_1037,N_14015,N_14377);
xnor UO_1038 (O_1038,N_14748,N_14076);
or UO_1039 (O_1039,N_14069,N_14960);
nor UO_1040 (O_1040,N_14598,N_14317);
or UO_1041 (O_1041,N_14279,N_14572);
xnor UO_1042 (O_1042,N_14221,N_14580);
nor UO_1043 (O_1043,N_14549,N_14389);
or UO_1044 (O_1044,N_14391,N_14345);
nand UO_1045 (O_1045,N_14684,N_14903);
or UO_1046 (O_1046,N_14543,N_14810);
or UO_1047 (O_1047,N_14791,N_14357);
nor UO_1048 (O_1048,N_14186,N_14817);
or UO_1049 (O_1049,N_14052,N_14523);
nor UO_1050 (O_1050,N_14501,N_14734);
nor UO_1051 (O_1051,N_14801,N_14010);
nor UO_1052 (O_1052,N_14144,N_14075);
or UO_1053 (O_1053,N_14697,N_14374);
nor UO_1054 (O_1054,N_14344,N_14519);
nand UO_1055 (O_1055,N_14001,N_14873);
nand UO_1056 (O_1056,N_14409,N_14095);
nand UO_1057 (O_1057,N_14184,N_14252);
and UO_1058 (O_1058,N_14976,N_14052);
nor UO_1059 (O_1059,N_14554,N_14822);
xor UO_1060 (O_1060,N_14675,N_14443);
xor UO_1061 (O_1061,N_14934,N_14152);
xnor UO_1062 (O_1062,N_14013,N_14904);
xnor UO_1063 (O_1063,N_14476,N_14563);
xnor UO_1064 (O_1064,N_14883,N_14632);
or UO_1065 (O_1065,N_14472,N_14395);
nor UO_1066 (O_1066,N_14527,N_14263);
nor UO_1067 (O_1067,N_14123,N_14308);
nand UO_1068 (O_1068,N_14219,N_14576);
and UO_1069 (O_1069,N_14871,N_14022);
nand UO_1070 (O_1070,N_14902,N_14268);
or UO_1071 (O_1071,N_14921,N_14538);
or UO_1072 (O_1072,N_14611,N_14684);
and UO_1073 (O_1073,N_14771,N_14232);
nor UO_1074 (O_1074,N_14318,N_14390);
xor UO_1075 (O_1075,N_14840,N_14827);
xor UO_1076 (O_1076,N_14163,N_14293);
xnor UO_1077 (O_1077,N_14098,N_14359);
xor UO_1078 (O_1078,N_14467,N_14997);
xnor UO_1079 (O_1079,N_14659,N_14222);
and UO_1080 (O_1080,N_14298,N_14911);
or UO_1081 (O_1081,N_14140,N_14703);
nand UO_1082 (O_1082,N_14791,N_14128);
nand UO_1083 (O_1083,N_14693,N_14666);
and UO_1084 (O_1084,N_14499,N_14817);
nand UO_1085 (O_1085,N_14599,N_14488);
nor UO_1086 (O_1086,N_14873,N_14482);
or UO_1087 (O_1087,N_14909,N_14460);
or UO_1088 (O_1088,N_14480,N_14622);
or UO_1089 (O_1089,N_14544,N_14261);
nand UO_1090 (O_1090,N_14105,N_14810);
and UO_1091 (O_1091,N_14890,N_14038);
nor UO_1092 (O_1092,N_14145,N_14730);
and UO_1093 (O_1093,N_14504,N_14448);
nand UO_1094 (O_1094,N_14853,N_14616);
nor UO_1095 (O_1095,N_14409,N_14499);
xnor UO_1096 (O_1096,N_14214,N_14422);
or UO_1097 (O_1097,N_14739,N_14625);
or UO_1098 (O_1098,N_14239,N_14247);
or UO_1099 (O_1099,N_14735,N_14544);
nand UO_1100 (O_1100,N_14528,N_14264);
nand UO_1101 (O_1101,N_14773,N_14100);
nand UO_1102 (O_1102,N_14472,N_14014);
or UO_1103 (O_1103,N_14267,N_14098);
nand UO_1104 (O_1104,N_14225,N_14251);
nand UO_1105 (O_1105,N_14316,N_14367);
or UO_1106 (O_1106,N_14823,N_14743);
nor UO_1107 (O_1107,N_14226,N_14065);
nand UO_1108 (O_1108,N_14617,N_14050);
nor UO_1109 (O_1109,N_14337,N_14281);
nand UO_1110 (O_1110,N_14542,N_14161);
and UO_1111 (O_1111,N_14114,N_14450);
nand UO_1112 (O_1112,N_14970,N_14095);
and UO_1113 (O_1113,N_14031,N_14931);
xor UO_1114 (O_1114,N_14657,N_14819);
and UO_1115 (O_1115,N_14120,N_14583);
nor UO_1116 (O_1116,N_14830,N_14110);
or UO_1117 (O_1117,N_14444,N_14046);
nand UO_1118 (O_1118,N_14243,N_14853);
and UO_1119 (O_1119,N_14157,N_14249);
or UO_1120 (O_1120,N_14535,N_14135);
nand UO_1121 (O_1121,N_14179,N_14588);
xnor UO_1122 (O_1122,N_14715,N_14685);
nand UO_1123 (O_1123,N_14117,N_14889);
nor UO_1124 (O_1124,N_14869,N_14877);
or UO_1125 (O_1125,N_14673,N_14827);
xor UO_1126 (O_1126,N_14365,N_14346);
nor UO_1127 (O_1127,N_14331,N_14588);
xor UO_1128 (O_1128,N_14464,N_14653);
xnor UO_1129 (O_1129,N_14434,N_14839);
nor UO_1130 (O_1130,N_14683,N_14702);
or UO_1131 (O_1131,N_14839,N_14287);
nor UO_1132 (O_1132,N_14623,N_14886);
xor UO_1133 (O_1133,N_14773,N_14855);
nand UO_1134 (O_1134,N_14453,N_14166);
nand UO_1135 (O_1135,N_14645,N_14459);
nor UO_1136 (O_1136,N_14567,N_14447);
or UO_1137 (O_1137,N_14299,N_14142);
or UO_1138 (O_1138,N_14068,N_14874);
and UO_1139 (O_1139,N_14184,N_14189);
nand UO_1140 (O_1140,N_14312,N_14073);
nand UO_1141 (O_1141,N_14045,N_14637);
xnor UO_1142 (O_1142,N_14703,N_14009);
nor UO_1143 (O_1143,N_14204,N_14835);
nor UO_1144 (O_1144,N_14020,N_14837);
xor UO_1145 (O_1145,N_14843,N_14720);
nand UO_1146 (O_1146,N_14878,N_14387);
nand UO_1147 (O_1147,N_14426,N_14512);
xor UO_1148 (O_1148,N_14029,N_14309);
nor UO_1149 (O_1149,N_14834,N_14903);
nand UO_1150 (O_1150,N_14184,N_14624);
nand UO_1151 (O_1151,N_14546,N_14631);
and UO_1152 (O_1152,N_14059,N_14156);
xor UO_1153 (O_1153,N_14841,N_14464);
xnor UO_1154 (O_1154,N_14622,N_14795);
or UO_1155 (O_1155,N_14854,N_14536);
and UO_1156 (O_1156,N_14162,N_14401);
xor UO_1157 (O_1157,N_14948,N_14697);
nand UO_1158 (O_1158,N_14927,N_14226);
nand UO_1159 (O_1159,N_14144,N_14538);
or UO_1160 (O_1160,N_14405,N_14579);
nor UO_1161 (O_1161,N_14184,N_14279);
nor UO_1162 (O_1162,N_14852,N_14105);
nor UO_1163 (O_1163,N_14892,N_14843);
and UO_1164 (O_1164,N_14120,N_14608);
nor UO_1165 (O_1165,N_14573,N_14649);
nand UO_1166 (O_1166,N_14052,N_14951);
xnor UO_1167 (O_1167,N_14450,N_14689);
nor UO_1168 (O_1168,N_14717,N_14327);
xnor UO_1169 (O_1169,N_14462,N_14851);
or UO_1170 (O_1170,N_14813,N_14577);
or UO_1171 (O_1171,N_14596,N_14087);
nand UO_1172 (O_1172,N_14708,N_14694);
and UO_1173 (O_1173,N_14212,N_14399);
nand UO_1174 (O_1174,N_14853,N_14226);
nor UO_1175 (O_1175,N_14880,N_14189);
xnor UO_1176 (O_1176,N_14068,N_14267);
nor UO_1177 (O_1177,N_14214,N_14432);
xor UO_1178 (O_1178,N_14620,N_14757);
nand UO_1179 (O_1179,N_14915,N_14487);
nor UO_1180 (O_1180,N_14630,N_14728);
xnor UO_1181 (O_1181,N_14848,N_14860);
or UO_1182 (O_1182,N_14446,N_14604);
nor UO_1183 (O_1183,N_14453,N_14749);
and UO_1184 (O_1184,N_14188,N_14933);
or UO_1185 (O_1185,N_14722,N_14760);
nor UO_1186 (O_1186,N_14992,N_14620);
or UO_1187 (O_1187,N_14522,N_14163);
xnor UO_1188 (O_1188,N_14690,N_14801);
nand UO_1189 (O_1189,N_14108,N_14961);
and UO_1190 (O_1190,N_14246,N_14243);
nor UO_1191 (O_1191,N_14711,N_14597);
xnor UO_1192 (O_1192,N_14321,N_14302);
nor UO_1193 (O_1193,N_14192,N_14298);
or UO_1194 (O_1194,N_14921,N_14355);
nor UO_1195 (O_1195,N_14467,N_14472);
and UO_1196 (O_1196,N_14444,N_14683);
or UO_1197 (O_1197,N_14752,N_14017);
nand UO_1198 (O_1198,N_14509,N_14204);
and UO_1199 (O_1199,N_14278,N_14269);
or UO_1200 (O_1200,N_14456,N_14223);
nand UO_1201 (O_1201,N_14355,N_14618);
xor UO_1202 (O_1202,N_14462,N_14696);
xor UO_1203 (O_1203,N_14860,N_14641);
nand UO_1204 (O_1204,N_14067,N_14031);
and UO_1205 (O_1205,N_14165,N_14776);
or UO_1206 (O_1206,N_14411,N_14958);
and UO_1207 (O_1207,N_14173,N_14222);
nand UO_1208 (O_1208,N_14964,N_14206);
nor UO_1209 (O_1209,N_14415,N_14698);
or UO_1210 (O_1210,N_14955,N_14001);
and UO_1211 (O_1211,N_14347,N_14816);
or UO_1212 (O_1212,N_14842,N_14168);
or UO_1213 (O_1213,N_14821,N_14210);
nand UO_1214 (O_1214,N_14798,N_14884);
nand UO_1215 (O_1215,N_14180,N_14991);
or UO_1216 (O_1216,N_14878,N_14296);
and UO_1217 (O_1217,N_14450,N_14797);
and UO_1218 (O_1218,N_14725,N_14127);
nor UO_1219 (O_1219,N_14046,N_14785);
nor UO_1220 (O_1220,N_14580,N_14688);
and UO_1221 (O_1221,N_14524,N_14048);
nor UO_1222 (O_1222,N_14160,N_14224);
xnor UO_1223 (O_1223,N_14335,N_14180);
nor UO_1224 (O_1224,N_14586,N_14192);
and UO_1225 (O_1225,N_14860,N_14170);
nor UO_1226 (O_1226,N_14693,N_14136);
or UO_1227 (O_1227,N_14463,N_14012);
or UO_1228 (O_1228,N_14939,N_14317);
and UO_1229 (O_1229,N_14201,N_14915);
and UO_1230 (O_1230,N_14403,N_14081);
nand UO_1231 (O_1231,N_14302,N_14138);
nor UO_1232 (O_1232,N_14400,N_14695);
or UO_1233 (O_1233,N_14179,N_14025);
and UO_1234 (O_1234,N_14303,N_14560);
and UO_1235 (O_1235,N_14039,N_14682);
and UO_1236 (O_1236,N_14838,N_14671);
or UO_1237 (O_1237,N_14903,N_14107);
and UO_1238 (O_1238,N_14144,N_14305);
nor UO_1239 (O_1239,N_14360,N_14262);
nand UO_1240 (O_1240,N_14760,N_14336);
and UO_1241 (O_1241,N_14284,N_14562);
nor UO_1242 (O_1242,N_14208,N_14279);
and UO_1243 (O_1243,N_14551,N_14590);
nand UO_1244 (O_1244,N_14742,N_14547);
nand UO_1245 (O_1245,N_14512,N_14754);
and UO_1246 (O_1246,N_14941,N_14848);
nor UO_1247 (O_1247,N_14651,N_14687);
nand UO_1248 (O_1248,N_14510,N_14397);
or UO_1249 (O_1249,N_14183,N_14737);
and UO_1250 (O_1250,N_14770,N_14196);
and UO_1251 (O_1251,N_14888,N_14995);
or UO_1252 (O_1252,N_14876,N_14971);
and UO_1253 (O_1253,N_14858,N_14277);
nand UO_1254 (O_1254,N_14232,N_14070);
and UO_1255 (O_1255,N_14901,N_14155);
and UO_1256 (O_1256,N_14536,N_14624);
nor UO_1257 (O_1257,N_14660,N_14950);
and UO_1258 (O_1258,N_14871,N_14530);
and UO_1259 (O_1259,N_14747,N_14431);
nor UO_1260 (O_1260,N_14055,N_14536);
xnor UO_1261 (O_1261,N_14937,N_14320);
and UO_1262 (O_1262,N_14301,N_14887);
nand UO_1263 (O_1263,N_14992,N_14017);
and UO_1264 (O_1264,N_14373,N_14984);
nor UO_1265 (O_1265,N_14058,N_14257);
nand UO_1266 (O_1266,N_14925,N_14051);
and UO_1267 (O_1267,N_14728,N_14284);
nor UO_1268 (O_1268,N_14746,N_14344);
nand UO_1269 (O_1269,N_14583,N_14846);
and UO_1270 (O_1270,N_14608,N_14869);
or UO_1271 (O_1271,N_14783,N_14782);
or UO_1272 (O_1272,N_14039,N_14736);
xor UO_1273 (O_1273,N_14709,N_14928);
nor UO_1274 (O_1274,N_14922,N_14934);
or UO_1275 (O_1275,N_14949,N_14088);
xor UO_1276 (O_1276,N_14548,N_14444);
or UO_1277 (O_1277,N_14408,N_14498);
xor UO_1278 (O_1278,N_14694,N_14165);
or UO_1279 (O_1279,N_14261,N_14418);
and UO_1280 (O_1280,N_14129,N_14836);
nand UO_1281 (O_1281,N_14569,N_14539);
xor UO_1282 (O_1282,N_14549,N_14785);
nand UO_1283 (O_1283,N_14778,N_14941);
nand UO_1284 (O_1284,N_14743,N_14676);
or UO_1285 (O_1285,N_14086,N_14177);
nor UO_1286 (O_1286,N_14906,N_14508);
nand UO_1287 (O_1287,N_14193,N_14722);
nand UO_1288 (O_1288,N_14929,N_14733);
nand UO_1289 (O_1289,N_14209,N_14529);
and UO_1290 (O_1290,N_14152,N_14269);
xor UO_1291 (O_1291,N_14414,N_14722);
xor UO_1292 (O_1292,N_14244,N_14091);
nor UO_1293 (O_1293,N_14127,N_14052);
xor UO_1294 (O_1294,N_14208,N_14680);
nand UO_1295 (O_1295,N_14892,N_14397);
xnor UO_1296 (O_1296,N_14576,N_14265);
nand UO_1297 (O_1297,N_14454,N_14280);
and UO_1298 (O_1298,N_14051,N_14705);
and UO_1299 (O_1299,N_14910,N_14030);
nand UO_1300 (O_1300,N_14059,N_14158);
and UO_1301 (O_1301,N_14862,N_14040);
nand UO_1302 (O_1302,N_14188,N_14526);
xor UO_1303 (O_1303,N_14253,N_14198);
xnor UO_1304 (O_1304,N_14713,N_14360);
nand UO_1305 (O_1305,N_14932,N_14056);
and UO_1306 (O_1306,N_14079,N_14917);
xnor UO_1307 (O_1307,N_14758,N_14846);
or UO_1308 (O_1308,N_14263,N_14892);
and UO_1309 (O_1309,N_14174,N_14014);
nand UO_1310 (O_1310,N_14327,N_14205);
and UO_1311 (O_1311,N_14464,N_14080);
xor UO_1312 (O_1312,N_14498,N_14737);
nand UO_1313 (O_1313,N_14897,N_14409);
nand UO_1314 (O_1314,N_14281,N_14388);
xor UO_1315 (O_1315,N_14823,N_14830);
or UO_1316 (O_1316,N_14382,N_14920);
nor UO_1317 (O_1317,N_14496,N_14267);
nor UO_1318 (O_1318,N_14711,N_14590);
xnor UO_1319 (O_1319,N_14155,N_14733);
and UO_1320 (O_1320,N_14169,N_14869);
or UO_1321 (O_1321,N_14185,N_14544);
nor UO_1322 (O_1322,N_14911,N_14074);
and UO_1323 (O_1323,N_14106,N_14596);
xnor UO_1324 (O_1324,N_14871,N_14396);
or UO_1325 (O_1325,N_14647,N_14121);
xor UO_1326 (O_1326,N_14212,N_14824);
nor UO_1327 (O_1327,N_14382,N_14554);
nor UO_1328 (O_1328,N_14394,N_14275);
and UO_1329 (O_1329,N_14369,N_14112);
xor UO_1330 (O_1330,N_14354,N_14844);
nor UO_1331 (O_1331,N_14508,N_14883);
or UO_1332 (O_1332,N_14514,N_14204);
and UO_1333 (O_1333,N_14844,N_14973);
xnor UO_1334 (O_1334,N_14253,N_14461);
xor UO_1335 (O_1335,N_14101,N_14164);
and UO_1336 (O_1336,N_14503,N_14593);
or UO_1337 (O_1337,N_14435,N_14999);
and UO_1338 (O_1338,N_14003,N_14861);
or UO_1339 (O_1339,N_14749,N_14516);
and UO_1340 (O_1340,N_14680,N_14927);
and UO_1341 (O_1341,N_14599,N_14412);
and UO_1342 (O_1342,N_14258,N_14841);
nor UO_1343 (O_1343,N_14789,N_14152);
and UO_1344 (O_1344,N_14509,N_14228);
and UO_1345 (O_1345,N_14833,N_14764);
xnor UO_1346 (O_1346,N_14631,N_14652);
nand UO_1347 (O_1347,N_14962,N_14249);
xor UO_1348 (O_1348,N_14909,N_14935);
nor UO_1349 (O_1349,N_14603,N_14691);
or UO_1350 (O_1350,N_14187,N_14266);
nand UO_1351 (O_1351,N_14369,N_14683);
nor UO_1352 (O_1352,N_14381,N_14750);
and UO_1353 (O_1353,N_14035,N_14874);
xor UO_1354 (O_1354,N_14308,N_14206);
nand UO_1355 (O_1355,N_14543,N_14811);
nand UO_1356 (O_1356,N_14384,N_14278);
or UO_1357 (O_1357,N_14482,N_14030);
nand UO_1358 (O_1358,N_14644,N_14659);
or UO_1359 (O_1359,N_14842,N_14704);
and UO_1360 (O_1360,N_14894,N_14475);
or UO_1361 (O_1361,N_14972,N_14451);
or UO_1362 (O_1362,N_14983,N_14464);
nand UO_1363 (O_1363,N_14858,N_14957);
or UO_1364 (O_1364,N_14592,N_14968);
nor UO_1365 (O_1365,N_14844,N_14345);
xor UO_1366 (O_1366,N_14243,N_14651);
and UO_1367 (O_1367,N_14514,N_14926);
xor UO_1368 (O_1368,N_14102,N_14551);
xnor UO_1369 (O_1369,N_14936,N_14327);
or UO_1370 (O_1370,N_14790,N_14989);
nor UO_1371 (O_1371,N_14132,N_14853);
nor UO_1372 (O_1372,N_14116,N_14194);
or UO_1373 (O_1373,N_14431,N_14940);
and UO_1374 (O_1374,N_14155,N_14800);
xor UO_1375 (O_1375,N_14738,N_14113);
nand UO_1376 (O_1376,N_14276,N_14639);
nor UO_1377 (O_1377,N_14097,N_14361);
nand UO_1378 (O_1378,N_14186,N_14422);
xor UO_1379 (O_1379,N_14416,N_14178);
and UO_1380 (O_1380,N_14692,N_14437);
nand UO_1381 (O_1381,N_14082,N_14167);
nand UO_1382 (O_1382,N_14041,N_14677);
nand UO_1383 (O_1383,N_14500,N_14940);
xnor UO_1384 (O_1384,N_14985,N_14554);
nor UO_1385 (O_1385,N_14109,N_14981);
or UO_1386 (O_1386,N_14109,N_14745);
xor UO_1387 (O_1387,N_14688,N_14391);
nand UO_1388 (O_1388,N_14804,N_14973);
nor UO_1389 (O_1389,N_14811,N_14988);
nor UO_1390 (O_1390,N_14324,N_14669);
and UO_1391 (O_1391,N_14712,N_14383);
nand UO_1392 (O_1392,N_14297,N_14307);
nor UO_1393 (O_1393,N_14822,N_14547);
and UO_1394 (O_1394,N_14092,N_14196);
xor UO_1395 (O_1395,N_14409,N_14107);
and UO_1396 (O_1396,N_14621,N_14022);
and UO_1397 (O_1397,N_14491,N_14795);
xnor UO_1398 (O_1398,N_14449,N_14873);
or UO_1399 (O_1399,N_14039,N_14430);
nor UO_1400 (O_1400,N_14752,N_14167);
and UO_1401 (O_1401,N_14523,N_14957);
and UO_1402 (O_1402,N_14533,N_14027);
and UO_1403 (O_1403,N_14896,N_14956);
nand UO_1404 (O_1404,N_14698,N_14329);
or UO_1405 (O_1405,N_14620,N_14530);
and UO_1406 (O_1406,N_14634,N_14798);
xnor UO_1407 (O_1407,N_14921,N_14662);
xor UO_1408 (O_1408,N_14730,N_14293);
nor UO_1409 (O_1409,N_14055,N_14078);
and UO_1410 (O_1410,N_14251,N_14631);
nand UO_1411 (O_1411,N_14223,N_14892);
and UO_1412 (O_1412,N_14194,N_14129);
nand UO_1413 (O_1413,N_14500,N_14181);
nand UO_1414 (O_1414,N_14645,N_14411);
xnor UO_1415 (O_1415,N_14331,N_14477);
nand UO_1416 (O_1416,N_14692,N_14379);
xnor UO_1417 (O_1417,N_14231,N_14984);
nand UO_1418 (O_1418,N_14861,N_14496);
nand UO_1419 (O_1419,N_14907,N_14718);
nand UO_1420 (O_1420,N_14904,N_14633);
nor UO_1421 (O_1421,N_14161,N_14384);
nor UO_1422 (O_1422,N_14258,N_14112);
or UO_1423 (O_1423,N_14648,N_14014);
and UO_1424 (O_1424,N_14465,N_14140);
and UO_1425 (O_1425,N_14635,N_14154);
nand UO_1426 (O_1426,N_14588,N_14803);
and UO_1427 (O_1427,N_14445,N_14385);
and UO_1428 (O_1428,N_14852,N_14934);
nor UO_1429 (O_1429,N_14564,N_14398);
or UO_1430 (O_1430,N_14308,N_14377);
and UO_1431 (O_1431,N_14564,N_14150);
nor UO_1432 (O_1432,N_14105,N_14081);
nor UO_1433 (O_1433,N_14521,N_14376);
or UO_1434 (O_1434,N_14583,N_14987);
nand UO_1435 (O_1435,N_14736,N_14106);
or UO_1436 (O_1436,N_14528,N_14725);
or UO_1437 (O_1437,N_14149,N_14048);
or UO_1438 (O_1438,N_14064,N_14215);
nand UO_1439 (O_1439,N_14545,N_14831);
or UO_1440 (O_1440,N_14219,N_14251);
nand UO_1441 (O_1441,N_14328,N_14263);
xor UO_1442 (O_1442,N_14092,N_14706);
nor UO_1443 (O_1443,N_14488,N_14092);
or UO_1444 (O_1444,N_14311,N_14678);
xnor UO_1445 (O_1445,N_14994,N_14234);
xnor UO_1446 (O_1446,N_14714,N_14565);
xnor UO_1447 (O_1447,N_14212,N_14957);
xnor UO_1448 (O_1448,N_14230,N_14865);
xor UO_1449 (O_1449,N_14195,N_14262);
nand UO_1450 (O_1450,N_14453,N_14290);
xor UO_1451 (O_1451,N_14124,N_14751);
nand UO_1452 (O_1452,N_14449,N_14152);
and UO_1453 (O_1453,N_14925,N_14857);
nand UO_1454 (O_1454,N_14791,N_14972);
nor UO_1455 (O_1455,N_14625,N_14900);
or UO_1456 (O_1456,N_14998,N_14686);
nor UO_1457 (O_1457,N_14989,N_14720);
and UO_1458 (O_1458,N_14029,N_14048);
xnor UO_1459 (O_1459,N_14770,N_14556);
xor UO_1460 (O_1460,N_14747,N_14946);
and UO_1461 (O_1461,N_14923,N_14177);
nor UO_1462 (O_1462,N_14038,N_14454);
and UO_1463 (O_1463,N_14585,N_14400);
nor UO_1464 (O_1464,N_14933,N_14113);
nand UO_1465 (O_1465,N_14228,N_14889);
and UO_1466 (O_1466,N_14236,N_14209);
nand UO_1467 (O_1467,N_14907,N_14454);
and UO_1468 (O_1468,N_14638,N_14414);
xnor UO_1469 (O_1469,N_14539,N_14115);
and UO_1470 (O_1470,N_14207,N_14644);
nor UO_1471 (O_1471,N_14150,N_14628);
or UO_1472 (O_1472,N_14936,N_14870);
or UO_1473 (O_1473,N_14723,N_14977);
nand UO_1474 (O_1474,N_14868,N_14413);
and UO_1475 (O_1475,N_14833,N_14082);
or UO_1476 (O_1476,N_14103,N_14633);
xor UO_1477 (O_1477,N_14253,N_14740);
nand UO_1478 (O_1478,N_14960,N_14239);
nor UO_1479 (O_1479,N_14426,N_14029);
nor UO_1480 (O_1480,N_14877,N_14052);
and UO_1481 (O_1481,N_14529,N_14595);
nor UO_1482 (O_1482,N_14407,N_14837);
nor UO_1483 (O_1483,N_14918,N_14671);
and UO_1484 (O_1484,N_14863,N_14033);
nor UO_1485 (O_1485,N_14887,N_14810);
nand UO_1486 (O_1486,N_14758,N_14788);
nor UO_1487 (O_1487,N_14474,N_14243);
xor UO_1488 (O_1488,N_14715,N_14488);
xor UO_1489 (O_1489,N_14972,N_14604);
nand UO_1490 (O_1490,N_14546,N_14973);
xor UO_1491 (O_1491,N_14842,N_14170);
nor UO_1492 (O_1492,N_14645,N_14989);
nor UO_1493 (O_1493,N_14239,N_14783);
and UO_1494 (O_1494,N_14022,N_14599);
xor UO_1495 (O_1495,N_14830,N_14711);
nand UO_1496 (O_1496,N_14604,N_14298);
nand UO_1497 (O_1497,N_14157,N_14045);
nor UO_1498 (O_1498,N_14038,N_14845);
xnor UO_1499 (O_1499,N_14651,N_14973);
xnor UO_1500 (O_1500,N_14841,N_14967);
and UO_1501 (O_1501,N_14382,N_14891);
nand UO_1502 (O_1502,N_14460,N_14617);
nand UO_1503 (O_1503,N_14624,N_14141);
and UO_1504 (O_1504,N_14565,N_14513);
nor UO_1505 (O_1505,N_14480,N_14371);
and UO_1506 (O_1506,N_14165,N_14702);
or UO_1507 (O_1507,N_14399,N_14382);
xor UO_1508 (O_1508,N_14336,N_14870);
or UO_1509 (O_1509,N_14052,N_14349);
nor UO_1510 (O_1510,N_14565,N_14137);
or UO_1511 (O_1511,N_14765,N_14084);
xor UO_1512 (O_1512,N_14192,N_14809);
xor UO_1513 (O_1513,N_14648,N_14751);
or UO_1514 (O_1514,N_14976,N_14977);
xor UO_1515 (O_1515,N_14690,N_14639);
xor UO_1516 (O_1516,N_14046,N_14840);
xnor UO_1517 (O_1517,N_14961,N_14927);
xnor UO_1518 (O_1518,N_14236,N_14840);
nor UO_1519 (O_1519,N_14936,N_14903);
or UO_1520 (O_1520,N_14613,N_14114);
nor UO_1521 (O_1521,N_14694,N_14916);
and UO_1522 (O_1522,N_14901,N_14411);
xnor UO_1523 (O_1523,N_14649,N_14572);
and UO_1524 (O_1524,N_14250,N_14954);
xnor UO_1525 (O_1525,N_14939,N_14689);
and UO_1526 (O_1526,N_14585,N_14370);
xor UO_1527 (O_1527,N_14823,N_14132);
and UO_1528 (O_1528,N_14848,N_14503);
or UO_1529 (O_1529,N_14057,N_14908);
nor UO_1530 (O_1530,N_14532,N_14710);
nor UO_1531 (O_1531,N_14294,N_14509);
xnor UO_1532 (O_1532,N_14588,N_14282);
xor UO_1533 (O_1533,N_14928,N_14989);
nor UO_1534 (O_1534,N_14888,N_14972);
nor UO_1535 (O_1535,N_14284,N_14278);
xnor UO_1536 (O_1536,N_14574,N_14872);
xor UO_1537 (O_1537,N_14391,N_14948);
nand UO_1538 (O_1538,N_14624,N_14419);
nand UO_1539 (O_1539,N_14983,N_14554);
xnor UO_1540 (O_1540,N_14391,N_14213);
xnor UO_1541 (O_1541,N_14813,N_14866);
xor UO_1542 (O_1542,N_14355,N_14496);
xor UO_1543 (O_1543,N_14775,N_14376);
or UO_1544 (O_1544,N_14485,N_14272);
nand UO_1545 (O_1545,N_14937,N_14764);
and UO_1546 (O_1546,N_14361,N_14110);
or UO_1547 (O_1547,N_14587,N_14320);
xor UO_1548 (O_1548,N_14035,N_14961);
xor UO_1549 (O_1549,N_14244,N_14331);
nand UO_1550 (O_1550,N_14363,N_14231);
or UO_1551 (O_1551,N_14096,N_14371);
and UO_1552 (O_1552,N_14120,N_14901);
nand UO_1553 (O_1553,N_14781,N_14714);
xor UO_1554 (O_1554,N_14241,N_14677);
xor UO_1555 (O_1555,N_14614,N_14211);
nor UO_1556 (O_1556,N_14998,N_14258);
xor UO_1557 (O_1557,N_14040,N_14300);
and UO_1558 (O_1558,N_14848,N_14994);
nand UO_1559 (O_1559,N_14693,N_14656);
xnor UO_1560 (O_1560,N_14761,N_14806);
and UO_1561 (O_1561,N_14247,N_14062);
xnor UO_1562 (O_1562,N_14854,N_14980);
xor UO_1563 (O_1563,N_14536,N_14177);
nand UO_1564 (O_1564,N_14814,N_14175);
nor UO_1565 (O_1565,N_14635,N_14640);
nand UO_1566 (O_1566,N_14527,N_14739);
nor UO_1567 (O_1567,N_14889,N_14276);
xor UO_1568 (O_1568,N_14253,N_14566);
nand UO_1569 (O_1569,N_14342,N_14728);
or UO_1570 (O_1570,N_14392,N_14739);
nor UO_1571 (O_1571,N_14241,N_14803);
nor UO_1572 (O_1572,N_14227,N_14790);
and UO_1573 (O_1573,N_14927,N_14048);
and UO_1574 (O_1574,N_14512,N_14587);
or UO_1575 (O_1575,N_14368,N_14723);
nand UO_1576 (O_1576,N_14793,N_14319);
xor UO_1577 (O_1577,N_14874,N_14685);
or UO_1578 (O_1578,N_14757,N_14574);
nor UO_1579 (O_1579,N_14343,N_14709);
or UO_1580 (O_1580,N_14645,N_14655);
xor UO_1581 (O_1581,N_14227,N_14753);
or UO_1582 (O_1582,N_14227,N_14861);
or UO_1583 (O_1583,N_14936,N_14309);
nor UO_1584 (O_1584,N_14537,N_14520);
or UO_1585 (O_1585,N_14696,N_14472);
xnor UO_1586 (O_1586,N_14766,N_14574);
or UO_1587 (O_1587,N_14546,N_14757);
xor UO_1588 (O_1588,N_14036,N_14531);
nand UO_1589 (O_1589,N_14346,N_14464);
and UO_1590 (O_1590,N_14589,N_14627);
nor UO_1591 (O_1591,N_14466,N_14132);
nor UO_1592 (O_1592,N_14183,N_14533);
or UO_1593 (O_1593,N_14860,N_14448);
and UO_1594 (O_1594,N_14816,N_14872);
xor UO_1595 (O_1595,N_14758,N_14205);
or UO_1596 (O_1596,N_14431,N_14899);
or UO_1597 (O_1597,N_14728,N_14787);
and UO_1598 (O_1598,N_14518,N_14951);
nand UO_1599 (O_1599,N_14253,N_14456);
xor UO_1600 (O_1600,N_14502,N_14658);
and UO_1601 (O_1601,N_14577,N_14132);
xor UO_1602 (O_1602,N_14112,N_14277);
or UO_1603 (O_1603,N_14181,N_14456);
and UO_1604 (O_1604,N_14152,N_14974);
nand UO_1605 (O_1605,N_14717,N_14254);
nor UO_1606 (O_1606,N_14301,N_14288);
and UO_1607 (O_1607,N_14633,N_14021);
nand UO_1608 (O_1608,N_14723,N_14369);
or UO_1609 (O_1609,N_14959,N_14574);
or UO_1610 (O_1610,N_14641,N_14620);
and UO_1611 (O_1611,N_14411,N_14095);
nand UO_1612 (O_1612,N_14444,N_14150);
nor UO_1613 (O_1613,N_14947,N_14639);
and UO_1614 (O_1614,N_14630,N_14890);
nand UO_1615 (O_1615,N_14259,N_14737);
and UO_1616 (O_1616,N_14122,N_14472);
xnor UO_1617 (O_1617,N_14587,N_14354);
xnor UO_1618 (O_1618,N_14247,N_14148);
nor UO_1619 (O_1619,N_14050,N_14987);
xor UO_1620 (O_1620,N_14572,N_14863);
nand UO_1621 (O_1621,N_14078,N_14545);
nand UO_1622 (O_1622,N_14121,N_14018);
nor UO_1623 (O_1623,N_14189,N_14989);
or UO_1624 (O_1624,N_14670,N_14148);
or UO_1625 (O_1625,N_14933,N_14255);
xor UO_1626 (O_1626,N_14987,N_14764);
nor UO_1627 (O_1627,N_14845,N_14570);
or UO_1628 (O_1628,N_14095,N_14606);
or UO_1629 (O_1629,N_14877,N_14405);
nand UO_1630 (O_1630,N_14347,N_14691);
xor UO_1631 (O_1631,N_14561,N_14720);
nand UO_1632 (O_1632,N_14029,N_14965);
or UO_1633 (O_1633,N_14866,N_14760);
or UO_1634 (O_1634,N_14537,N_14982);
nor UO_1635 (O_1635,N_14012,N_14308);
xnor UO_1636 (O_1636,N_14838,N_14347);
or UO_1637 (O_1637,N_14706,N_14227);
nand UO_1638 (O_1638,N_14871,N_14965);
nand UO_1639 (O_1639,N_14106,N_14782);
and UO_1640 (O_1640,N_14357,N_14264);
or UO_1641 (O_1641,N_14671,N_14230);
or UO_1642 (O_1642,N_14836,N_14307);
and UO_1643 (O_1643,N_14891,N_14760);
xor UO_1644 (O_1644,N_14943,N_14014);
nor UO_1645 (O_1645,N_14619,N_14987);
nor UO_1646 (O_1646,N_14427,N_14539);
and UO_1647 (O_1647,N_14418,N_14308);
or UO_1648 (O_1648,N_14433,N_14311);
nand UO_1649 (O_1649,N_14884,N_14672);
xor UO_1650 (O_1650,N_14569,N_14677);
and UO_1651 (O_1651,N_14525,N_14459);
nand UO_1652 (O_1652,N_14969,N_14929);
nand UO_1653 (O_1653,N_14924,N_14498);
nand UO_1654 (O_1654,N_14560,N_14520);
nor UO_1655 (O_1655,N_14294,N_14731);
or UO_1656 (O_1656,N_14409,N_14334);
and UO_1657 (O_1657,N_14393,N_14396);
nand UO_1658 (O_1658,N_14822,N_14465);
xor UO_1659 (O_1659,N_14588,N_14009);
nand UO_1660 (O_1660,N_14657,N_14826);
and UO_1661 (O_1661,N_14253,N_14800);
and UO_1662 (O_1662,N_14301,N_14845);
xor UO_1663 (O_1663,N_14526,N_14936);
and UO_1664 (O_1664,N_14111,N_14060);
or UO_1665 (O_1665,N_14475,N_14705);
or UO_1666 (O_1666,N_14454,N_14782);
nor UO_1667 (O_1667,N_14293,N_14900);
or UO_1668 (O_1668,N_14724,N_14170);
nor UO_1669 (O_1669,N_14616,N_14636);
xnor UO_1670 (O_1670,N_14292,N_14233);
xnor UO_1671 (O_1671,N_14410,N_14694);
or UO_1672 (O_1672,N_14472,N_14798);
nand UO_1673 (O_1673,N_14578,N_14082);
xor UO_1674 (O_1674,N_14322,N_14520);
nand UO_1675 (O_1675,N_14304,N_14534);
nor UO_1676 (O_1676,N_14908,N_14396);
or UO_1677 (O_1677,N_14682,N_14146);
nand UO_1678 (O_1678,N_14167,N_14169);
nor UO_1679 (O_1679,N_14809,N_14372);
or UO_1680 (O_1680,N_14876,N_14858);
or UO_1681 (O_1681,N_14418,N_14405);
or UO_1682 (O_1682,N_14968,N_14505);
nor UO_1683 (O_1683,N_14778,N_14186);
xnor UO_1684 (O_1684,N_14916,N_14000);
nor UO_1685 (O_1685,N_14246,N_14831);
xnor UO_1686 (O_1686,N_14395,N_14592);
nor UO_1687 (O_1687,N_14314,N_14458);
nand UO_1688 (O_1688,N_14648,N_14053);
nand UO_1689 (O_1689,N_14943,N_14342);
nor UO_1690 (O_1690,N_14968,N_14175);
nand UO_1691 (O_1691,N_14952,N_14806);
nor UO_1692 (O_1692,N_14405,N_14716);
or UO_1693 (O_1693,N_14323,N_14640);
and UO_1694 (O_1694,N_14627,N_14557);
or UO_1695 (O_1695,N_14234,N_14376);
or UO_1696 (O_1696,N_14719,N_14968);
and UO_1697 (O_1697,N_14400,N_14927);
xor UO_1698 (O_1698,N_14367,N_14922);
nand UO_1699 (O_1699,N_14142,N_14790);
or UO_1700 (O_1700,N_14478,N_14813);
nand UO_1701 (O_1701,N_14226,N_14892);
nor UO_1702 (O_1702,N_14344,N_14593);
or UO_1703 (O_1703,N_14049,N_14361);
and UO_1704 (O_1704,N_14641,N_14578);
nor UO_1705 (O_1705,N_14930,N_14134);
nor UO_1706 (O_1706,N_14322,N_14094);
or UO_1707 (O_1707,N_14707,N_14810);
or UO_1708 (O_1708,N_14214,N_14849);
nor UO_1709 (O_1709,N_14809,N_14245);
nand UO_1710 (O_1710,N_14739,N_14661);
and UO_1711 (O_1711,N_14421,N_14070);
nor UO_1712 (O_1712,N_14245,N_14546);
or UO_1713 (O_1713,N_14504,N_14385);
or UO_1714 (O_1714,N_14854,N_14607);
nor UO_1715 (O_1715,N_14788,N_14958);
nor UO_1716 (O_1716,N_14708,N_14565);
nand UO_1717 (O_1717,N_14482,N_14969);
nand UO_1718 (O_1718,N_14395,N_14566);
nor UO_1719 (O_1719,N_14977,N_14442);
or UO_1720 (O_1720,N_14417,N_14442);
nand UO_1721 (O_1721,N_14736,N_14011);
nand UO_1722 (O_1722,N_14645,N_14574);
nand UO_1723 (O_1723,N_14958,N_14678);
or UO_1724 (O_1724,N_14724,N_14719);
nand UO_1725 (O_1725,N_14821,N_14536);
xor UO_1726 (O_1726,N_14904,N_14500);
or UO_1727 (O_1727,N_14463,N_14195);
or UO_1728 (O_1728,N_14184,N_14362);
nand UO_1729 (O_1729,N_14175,N_14560);
xnor UO_1730 (O_1730,N_14327,N_14798);
nand UO_1731 (O_1731,N_14787,N_14329);
nand UO_1732 (O_1732,N_14296,N_14363);
xor UO_1733 (O_1733,N_14729,N_14524);
nand UO_1734 (O_1734,N_14215,N_14509);
or UO_1735 (O_1735,N_14854,N_14487);
nand UO_1736 (O_1736,N_14520,N_14067);
xnor UO_1737 (O_1737,N_14754,N_14822);
and UO_1738 (O_1738,N_14926,N_14924);
nor UO_1739 (O_1739,N_14211,N_14044);
xnor UO_1740 (O_1740,N_14492,N_14977);
and UO_1741 (O_1741,N_14412,N_14741);
nor UO_1742 (O_1742,N_14629,N_14504);
or UO_1743 (O_1743,N_14146,N_14359);
nand UO_1744 (O_1744,N_14686,N_14250);
or UO_1745 (O_1745,N_14916,N_14440);
nand UO_1746 (O_1746,N_14952,N_14600);
xor UO_1747 (O_1747,N_14924,N_14781);
nor UO_1748 (O_1748,N_14244,N_14177);
nor UO_1749 (O_1749,N_14774,N_14228);
and UO_1750 (O_1750,N_14657,N_14165);
nand UO_1751 (O_1751,N_14070,N_14271);
nand UO_1752 (O_1752,N_14681,N_14189);
nor UO_1753 (O_1753,N_14339,N_14748);
and UO_1754 (O_1754,N_14305,N_14504);
and UO_1755 (O_1755,N_14994,N_14598);
nor UO_1756 (O_1756,N_14863,N_14347);
nor UO_1757 (O_1757,N_14671,N_14201);
xnor UO_1758 (O_1758,N_14866,N_14218);
nor UO_1759 (O_1759,N_14652,N_14641);
nand UO_1760 (O_1760,N_14490,N_14718);
nor UO_1761 (O_1761,N_14712,N_14824);
or UO_1762 (O_1762,N_14444,N_14544);
and UO_1763 (O_1763,N_14677,N_14162);
or UO_1764 (O_1764,N_14315,N_14226);
or UO_1765 (O_1765,N_14004,N_14071);
and UO_1766 (O_1766,N_14960,N_14146);
nor UO_1767 (O_1767,N_14631,N_14055);
nor UO_1768 (O_1768,N_14530,N_14459);
nand UO_1769 (O_1769,N_14385,N_14471);
xnor UO_1770 (O_1770,N_14805,N_14078);
nor UO_1771 (O_1771,N_14846,N_14474);
and UO_1772 (O_1772,N_14183,N_14724);
xor UO_1773 (O_1773,N_14438,N_14520);
nor UO_1774 (O_1774,N_14565,N_14860);
nand UO_1775 (O_1775,N_14349,N_14771);
nand UO_1776 (O_1776,N_14719,N_14784);
nor UO_1777 (O_1777,N_14593,N_14293);
xnor UO_1778 (O_1778,N_14632,N_14782);
and UO_1779 (O_1779,N_14912,N_14917);
and UO_1780 (O_1780,N_14827,N_14525);
xnor UO_1781 (O_1781,N_14060,N_14274);
or UO_1782 (O_1782,N_14660,N_14038);
or UO_1783 (O_1783,N_14216,N_14969);
or UO_1784 (O_1784,N_14611,N_14882);
or UO_1785 (O_1785,N_14818,N_14110);
or UO_1786 (O_1786,N_14733,N_14381);
xnor UO_1787 (O_1787,N_14612,N_14206);
nand UO_1788 (O_1788,N_14927,N_14954);
nor UO_1789 (O_1789,N_14085,N_14478);
or UO_1790 (O_1790,N_14062,N_14173);
or UO_1791 (O_1791,N_14207,N_14918);
or UO_1792 (O_1792,N_14704,N_14751);
nor UO_1793 (O_1793,N_14591,N_14277);
nor UO_1794 (O_1794,N_14399,N_14950);
and UO_1795 (O_1795,N_14628,N_14248);
and UO_1796 (O_1796,N_14071,N_14036);
or UO_1797 (O_1797,N_14931,N_14104);
or UO_1798 (O_1798,N_14624,N_14066);
nor UO_1799 (O_1799,N_14162,N_14684);
xor UO_1800 (O_1800,N_14246,N_14899);
and UO_1801 (O_1801,N_14466,N_14833);
and UO_1802 (O_1802,N_14000,N_14361);
or UO_1803 (O_1803,N_14098,N_14721);
xnor UO_1804 (O_1804,N_14199,N_14694);
nor UO_1805 (O_1805,N_14938,N_14462);
nand UO_1806 (O_1806,N_14630,N_14856);
or UO_1807 (O_1807,N_14246,N_14149);
nand UO_1808 (O_1808,N_14607,N_14428);
nor UO_1809 (O_1809,N_14835,N_14189);
and UO_1810 (O_1810,N_14821,N_14204);
xnor UO_1811 (O_1811,N_14261,N_14649);
xor UO_1812 (O_1812,N_14542,N_14672);
or UO_1813 (O_1813,N_14824,N_14106);
or UO_1814 (O_1814,N_14795,N_14822);
or UO_1815 (O_1815,N_14156,N_14271);
or UO_1816 (O_1816,N_14113,N_14792);
xnor UO_1817 (O_1817,N_14289,N_14175);
nand UO_1818 (O_1818,N_14166,N_14074);
nor UO_1819 (O_1819,N_14853,N_14636);
nand UO_1820 (O_1820,N_14254,N_14870);
or UO_1821 (O_1821,N_14877,N_14323);
and UO_1822 (O_1822,N_14216,N_14470);
and UO_1823 (O_1823,N_14255,N_14812);
xnor UO_1824 (O_1824,N_14823,N_14921);
nand UO_1825 (O_1825,N_14600,N_14941);
nor UO_1826 (O_1826,N_14238,N_14256);
and UO_1827 (O_1827,N_14714,N_14518);
nor UO_1828 (O_1828,N_14265,N_14080);
or UO_1829 (O_1829,N_14773,N_14211);
or UO_1830 (O_1830,N_14004,N_14353);
xor UO_1831 (O_1831,N_14802,N_14614);
xor UO_1832 (O_1832,N_14102,N_14380);
and UO_1833 (O_1833,N_14245,N_14191);
xnor UO_1834 (O_1834,N_14020,N_14545);
and UO_1835 (O_1835,N_14295,N_14490);
xor UO_1836 (O_1836,N_14946,N_14028);
nand UO_1837 (O_1837,N_14335,N_14834);
nor UO_1838 (O_1838,N_14642,N_14179);
and UO_1839 (O_1839,N_14338,N_14302);
nand UO_1840 (O_1840,N_14232,N_14980);
or UO_1841 (O_1841,N_14058,N_14916);
and UO_1842 (O_1842,N_14910,N_14554);
nor UO_1843 (O_1843,N_14782,N_14729);
and UO_1844 (O_1844,N_14890,N_14182);
or UO_1845 (O_1845,N_14419,N_14764);
or UO_1846 (O_1846,N_14391,N_14905);
nand UO_1847 (O_1847,N_14673,N_14223);
nor UO_1848 (O_1848,N_14230,N_14272);
and UO_1849 (O_1849,N_14799,N_14220);
nand UO_1850 (O_1850,N_14054,N_14249);
nand UO_1851 (O_1851,N_14656,N_14521);
nor UO_1852 (O_1852,N_14181,N_14096);
or UO_1853 (O_1853,N_14598,N_14447);
nand UO_1854 (O_1854,N_14775,N_14748);
and UO_1855 (O_1855,N_14974,N_14536);
and UO_1856 (O_1856,N_14225,N_14911);
nand UO_1857 (O_1857,N_14680,N_14427);
and UO_1858 (O_1858,N_14981,N_14757);
xor UO_1859 (O_1859,N_14042,N_14737);
xnor UO_1860 (O_1860,N_14655,N_14124);
nor UO_1861 (O_1861,N_14748,N_14417);
xor UO_1862 (O_1862,N_14156,N_14340);
nand UO_1863 (O_1863,N_14283,N_14375);
nand UO_1864 (O_1864,N_14735,N_14347);
xnor UO_1865 (O_1865,N_14148,N_14561);
nor UO_1866 (O_1866,N_14342,N_14983);
nand UO_1867 (O_1867,N_14560,N_14592);
nor UO_1868 (O_1868,N_14250,N_14182);
and UO_1869 (O_1869,N_14688,N_14675);
and UO_1870 (O_1870,N_14005,N_14897);
xnor UO_1871 (O_1871,N_14099,N_14659);
or UO_1872 (O_1872,N_14662,N_14616);
and UO_1873 (O_1873,N_14416,N_14603);
xnor UO_1874 (O_1874,N_14115,N_14299);
xnor UO_1875 (O_1875,N_14359,N_14171);
nand UO_1876 (O_1876,N_14161,N_14601);
or UO_1877 (O_1877,N_14369,N_14003);
nand UO_1878 (O_1878,N_14112,N_14403);
xnor UO_1879 (O_1879,N_14603,N_14106);
and UO_1880 (O_1880,N_14488,N_14048);
nand UO_1881 (O_1881,N_14100,N_14594);
nor UO_1882 (O_1882,N_14428,N_14898);
nand UO_1883 (O_1883,N_14356,N_14412);
and UO_1884 (O_1884,N_14193,N_14366);
and UO_1885 (O_1885,N_14912,N_14734);
or UO_1886 (O_1886,N_14968,N_14694);
nor UO_1887 (O_1887,N_14488,N_14464);
xnor UO_1888 (O_1888,N_14375,N_14486);
or UO_1889 (O_1889,N_14128,N_14236);
nand UO_1890 (O_1890,N_14929,N_14562);
nor UO_1891 (O_1891,N_14368,N_14638);
xor UO_1892 (O_1892,N_14156,N_14284);
xnor UO_1893 (O_1893,N_14352,N_14233);
or UO_1894 (O_1894,N_14327,N_14027);
xor UO_1895 (O_1895,N_14589,N_14357);
or UO_1896 (O_1896,N_14695,N_14637);
nor UO_1897 (O_1897,N_14091,N_14892);
nor UO_1898 (O_1898,N_14715,N_14541);
nand UO_1899 (O_1899,N_14534,N_14456);
or UO_1900 (O_1900,N_14430,N_14127);
xor UO_1901 (O_1901,N_14285,N_14024);
and UO_1902 (O_1902,N_14293,N_14625);
and UO_1903 (O_1903,N_14412,N_14635);
or UO_1904 (O_1904,N_14842,N_14463);
or UO_1905 (O_1905,N_14606,N_14784);
or UO_1906 (O_1906,N_14714,N_14972);
xor UO_1907 (O_1907,N_14327,N_14641);
nand UO_1908 (O_1908,N_14024,N_14883);
xor UO_1909 (O_1909,N_14584,N_14236);
and UO_1910 (O_1910,N_14980,N_14548);
or UO_1911 (O_1911,N_14852,N_14833);
nor UO_1912 (O_1912,N_14948,N_14884);
nor UO_1913 (O_1913,N_14522,N_14033);
xnor UO_1914 (O_1914,N_14003,N_14638);
xnor UO_1915 (O_1915,N_14209,N_14629);
and UO_1916 (O_1916,N_14768,N_14090);
xor UO_1917 (O_1917,N_14901,N_14725);
nand UO_1918 (O_1918,N_14343,N_14999);
and UO_1919 (O_1919,N_14074,N_14049);
xor UO_1920 (O_1920,N_14823,N_14249);
or UO_1921 (O_1921,N_14089,N_14810);
nand UO_1922 (O_1922,N_14553,N_14759);
xnor UO_1923 (O_1923,N_14889,N_14983);
xor UO_1924 (O_1924,N_14821,N_14260);
and UO_1925 (O_1925,N_14980,N_14393);
xnor UO_1926 (O_1926,N_14225,N_14714);
nor UO_1927 (O_1927,N_14566,N_14951);
nand UO_1928 (O_1928,N_14035,N_14884);
nor UO_1929 (O_1929,N_14511,N_14065);
nor UO_1930 (O_1930,N_14936,N_14882);
nand UO_1931 (O_1931,N_14389,N_14126);
and UO_1932 (O_1932,N_14003,N_14252);
nor UO_1933 (O_1933,N_14378,N_14929);
nor UO_1934 (O_1934,N_14463,N_14037);
xor UO_1935 (O_1935,N_14756,N_14057);
nor UO_1936 (O_1936,N_14355,N_14133);
xor UO_1937 (O_1937,N_14135,N_14459);
or UO_1938 (O_1938,N_14154,N_14663);
xor UO_1939 (O_1939,N_14678,N_14071);
and UO_1940 (O_1940,N_14726,N_14401);
xnor UO_1941 (O_1941,N_14667,N_14258);
and UO_1942 (O_1942,N_14178,N_14077);
nor UO_1943 (O_1943,N_14560,N_14373);
xor UO_1944 (O_1944,N_14687,N_14554);
and UO_1945 (O_1945,N_14827,N_14615);
nor UO_1946 (O_1946,N_14070,N_14904);
and UO_1947 (O_1947,N_14006,N_14885);
and UO_1948 (O_1948,N_14187,N_14688);
nand UO_1949 (O_1949,N_14127,N_14921);
xnor UO_1950 (O_1950,N_14705,N_14601);
nor UO_1951 (O_1951,N_14525,N_14196);
or UO_1952 (O_1952,N_14112,N_14559);
or UO_1953 (O_1953,N_14447,N_14137);
nor UO_1954 (O_1954,N_14210,N_14261);
nand UO_1955 (O_1955,N_14816,N_14378);
and UO_1956 (O_1956,N_14123,N_14863);
nor UO_1957 (O_1957,N_14972,N_14655);
nor UO_1958 (O_1958,N_14018,N_14867);
or UO_1959 (O_1959,N_14128,N_14108);
nor UO_1960 (O_1960,N_14180,N_14638);
nand UO_1961 (O_1961,N_14668,N_14889);
nand UO_1962 (O_1962,N_14253,N_14294);
nand UO_1963 (O_1963,N_14290,N_14273);
nor UO_1964 (O_1964,N_14769,N_14148);
and UO_1965 (O_1965,N_14200,N_14153);
and UO_1966 (O_1966,N_14662,N_14156);
nor UO_1967 (O_1967,N_14431,N_14478);
nand UO_1968 (O_1968,N_14873,N_14818);
nor UO_1969 (O_1969,N_14059,N_14393);
or UO_1970 (O_1970,N_14526,N_14660);
xor UO_1971 (O_1971,N_14032,N_14268);
nand UO_1972 (O_1972,N_14956,N_14156);
or UO_1973 (O_1973,N_14469,N_14183);
and UO_1974 (O_1974,N_14587,N_14749);
or UO_1975 (O_1975,N_14396,N_14598);
nand UO_1976 (O_1976,N_14635,N_14093);
nor UO_1977 (O_1977,N_14351,N_14242);
or UO_1978 (O_1978,N_14756,N_14451);
and UO_1979 (O_1979,N_14804,N_14521);
and UO_1980 (O_1980,N_14072,N_14638);
nand UO_1981 (O_1981,N_14572,N_14529);
xnor UO_1982 (O_1982,N_14636,N_14852);
and UO_1983 (O_1983,N_14360,N_14914);
nand UO_1984 (O_1984,N_14098,N_14608);
or UO_1985 (O_1985,N_14818,N_14016);
or UO_1986 (O_1986,N_14004,N_14070);
nor UO_1987 (O_1987,N_14211,N_14787);
nand UO_1988 (O_1988,N_14865,N_14538);
nand UO_1989 (O_1989,N_14380,N_14633);
and UO_1990 (O_1990,N_14303,N_14961);
nor UO_1991 (O_1991,N_14498,N_14788);
xnor UO_1992 (O_1992,N_14809,N_14652);
nand UO_1993 (O_1993,N_14560,N_14504);
or UO_1994 (O_1994,N_14244,N_14600);
nor UO_1995 (O_1995,N_14474,N_14615);
nand UO_1996 (O_1996,N_14222,N_14489);
or UO_1997 (O_1997,N_14241,N_14777);
or UO_1998 (O_1998,N_14382,N_14409);
xor UO_1999 (O_1999,N_14630,N_14707);
endmodule