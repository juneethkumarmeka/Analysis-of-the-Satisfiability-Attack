module basic_2000_20000_2500_100_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nand U0 (N_0,In_12,In_906);
xnor U1 (N_1,In_274,In_345);
nand U2 (N_2,In_103,In_326);
or U3 (N_3,In_634,In_1596);
nand U4 (N_4,In_370,In_1968);
nand U5 (N_5,In_921,In_329);
xnor U6 (N_6,In_1957,In_1213);
or U7 (N_7,In_629,In_500);
and U8 (N_8,In_1222,In_1660);
and U9 (N_9,In_1007,In_1654);
xor U10 (N_10,In_243,In_963);
and U11 (N_11,In_427,In_491);
or U12 (N_12,In_1127,In_418);
nand U13 (N_13,In_1062,In_76);
or U14 (N_14,In_211,In_1652);
nand U15 (N_15,In_167,In_1872);
or U16 (N_16,In_1363,In_225);
nand U17 (N_17,In_907,In_1891);
and U18 (N_18,In_831,In_1029);
xnor U19 (N_19,In_1651,In_368);
or U20 (N_20,In_1734,In_1852);
and U21 (N_21,In_65,In_461);
nor U22 (N_22,In_842,In_1430);
nand U23 (N_23,In_861,In_1815);
and U24 (N_24,In_312,In_880);
nor U25 (N_25,In_955,In_388);
nor U26 (N_26,In_1884,In_510);
nand U27 (N_27,In_760,In_337);
nand U28 (N_28,In_235,In_1955);
xnor U29 (N_29,In_622,In_1827);
nand U30 (N_30,In_625,In_1328);
xor U31 (N_31,In_1105,In_1542);
or U32 (N_32,In_1488,In_245);
xnor U33 (N_33,In_1672,In_297);
nor U34 (N_34,In_507,In_177);
nand U35 (N_35,In_1706,In_1440);
and U36 (N_36,In_1677,In_636);
or U37 (N_37,In_1124,In_269);
xnor U38 (N_38,In_1251,In_1317);
and U39 (N_39,In_1063,In_346);
nand U40 (N_40,In_737,In_8);
xor U41 (N_41,In_1560,In_1113);
and U42 (N_42,In_209,In_1163);
nand U43 (N_43,In_202,In_778);
and U44 (N_44,In_795,In_1004);
and U45 (N_45,In_813,In_695);
nor U46 (N_46,In_1885,In_1749);
nor U47 (N_47,In_1189,In_335);
xnor U48 (N_48,In_435,In_1271);
or U49 (N_49,In_118,In_414);
and U50 (N_50,In_1368,In_1559);
and U51 (N_51,In_837,In_811);
nand U52 (N_52,In_1716,In_536);
nor U53 (N_53,In_1412,In_988);
or U54 (N_54,In_254,In_561);
xor U55 (N_55,In_1682,In_1835);
xnor U56 (N_56,In_1080,In_678);
nand U57 (N_57,In_1620,In_1057);
nand U58 (N_58,In_1042,In_242);
xor U59 (N_59,In_1608,In_293);
xor U60 (N_60,In_1226,In_1595);
nor U61 (N_61,In_727,In_1110);
nor U62 (N_62,In_1856,In_983);
xor U63 (N_63,In_431,In_1896);
or U64 (N_64,In_1438,In_303);
nor U65 (N_65,In_1107,In_24);
or U66 (N_66,In_71,In_94);
or U67 (N_67,In_1050,In_1990);
or U68 (N_68,In_1805,In_815);
or U69 (N_69,In_640,In_492);
and U70 (N_70,In_1209,In_1300);
nand U71 (N_71,In_1250,In_1703);
nand U72 (N_72,In_630,In_1155);
nor U73 (N_73,In_908,In_1808);
xor U74 (N_74,In_573,In_29);
nor U75 (N_75,In_321,In_1619);
nor U76 (N_76,In_1294,In_1958);
xor U77 (N_77,In_125,In_393);
nand U78 (N_78,In_1413,In_1941);
or U79 (N_79,In_358,In_708);
and U80 (N_80,In_474,In_133);
or U81 (N_81,In_115,In_1859);
or U82 (N_82,In_1159,In_1888);
and U83 (N_83,In_542,In_472);
or U84 (N_84,In_408,In_1252);
nor U85 (N_85,In_978,In_657);
xnor U86 (N_86,In_1332,In_598);
xor U87 (N_87,In_1244,In_193);
nand U88 (N_88,In_1006,In_1115);
and U89 (N_89,In_462,In_1579);
nor U90 (N_90,In_1870,In_54);
nand U91 (N_91,In_1366,In_1290);
and U92 (N_92,In_1178,In_1594);
xnor U93 (N_93,In_1785,In_620);
and U94 (N_94,In_1587,In_974);
nand U95 (N_95,In_199,In_1425);
nor U96 (N_96,In_399,In_338);
or U97 (N_97,In_612,In_247);
and U98 (N_98,In_713,In_1642);
nor U99 (N_99,In_1784,In_445);
nor U100 (N_100,In_1517,In_336);
or U101 (N_101,In_1765,In_1934);
or U102 (N_102,In_1347,In_529);
nand U103 (N_103,In_1128,In_1617);
nor U104 (N_104,In_330,In_1303);
and U105 (N_105,In_1218,In_1174);
nor U106 (N_106,In_1378,In_503);
xnor U107 (N_107,In_1699,In_188);
or U108 (N_108,In_628,In_1370);
nor U109 (N_109,In_1771,In_1612);
and U110 (N_110,In_1479,In_1101);
nor U111 (N_111,In_1460,In_1588);
or U112 (N_112,In_949,In_859);
and U113 (N_113,In_1089,In_944);
nand U114 (N_114,In_531,In_410);
nor U115 (N_115,In_17,In_1287);
nor U116 (N_116,In_201,In_555);
and U117 (N_117,In_191,In_1148);
nor U118 (N_118,In_1286,In_1814);
nor U119 (N_119,In_705,In_1622);
nand U120 (N_120,In_1025,In_960);
or U121 (N_121,In_977,In_796);
xor U122 (N_122,In_1601,In_1624);
or U123 (N_123,In_68,In_1635);
nor U124 (N_124,In_315,In_1014);
nand U125 (N_125,In_590,In_1);
or U126 (N_126,In_271,In_463);
xor U127 (N_127,In_846,In_1139);
nand U128 (N_128,In_877,In_1708);
or U129 (N_129,In_1843,In_878);
nand U130 (N_130,In_642,In_1506);
xnor U131 (N_131,In_1343,In_1758);
nand U132 (N_132,In_353,In_22);
nand U133 (N_133,In_1834,In_549);
xor U134 (N_134,In_728,In_925);
and U135 (N_135,In_350,In_646);
and U136 (N_136,In_751,In_1613);
xnor U137 (N_137,In_1680,In_1496);
or U138 (N_138,In_4,In_902);
xor U139 (N_139,In_1992,In_654);
or U140 (N_140,In_46,In_1033);
xnor U141 (N_141,In_25,In_311);
and U142 (N_142,In_1600,In_1787);
nor U143 (N_143,In_92,In_1298);
nand U144 (N_144,In_993,In_164);
nand U145 (N_145,In_1136,In_422);
nand U146 (N_146,In_145,In_119);
and U147 (N_147,In_1848,In_306);
nand U148 (N_148,In_524,In_1515);
or U149 (N_149,In_79,In_73);
and U150 (N_150,In_707,In_97);
and U151 (N_151,In_1340,In_539);
and U152 (N_152,In_954,In_107);
nand U153 (N_153,In_364,In_1272);
nor U154 (N_154,In_912,In_1754);
nor U155 (N_155,In_231,In_540);
and U156 (N_156,In_100,In_319);
xnor U157 (N_157,In_765,In_1694);
and U158 (N_158,In_722,In_547);
or U159 (N_159,In_1362,In_515);
nand U160 (N_160,In_658,In_819);
xor U161 (N_161,In_631,In_1054);
xnor U162 (N_162,In_1149,In_351);
and U163 (N_163,In_697,In_1395);
and U164 (N_164,In_270,In_317);
and U165 (N_165,In_369,In_348);
or U166 (N_166,In_522,In_1830);
or U167 (N_167,In_26,In_273);
or U168 (N_168,In_1727,In_1043);
nor U169 (N_169,In_1273,In_1188);
nor U170 (N_170,In_893,In_1507);
or U171 (N_171,In_31,In_126);
or U172 (N_172,In_742,In_123);
nand U173 (N_173,In_1925,In_1372);
nor U174 (N_174,In_1943,In_23);
nand U175 (N_175,In_101,In_1659);
or U176 (N_176,In_1932,In_1711);
and U177 (N_177,In_721,In_0);
nor U178 (N_178,In_1569,In_1772);
and U179 (N_179,In_232,In_953);
and U180 (N_180,In_817,In_552);
and U181 (N_181,In_733,In_537);
xnor U182 (N_182,In_1602,In_1324);
and U183 (N_183,In_930,In_998);
nand U184 (N_184,In_1307,In_980);
nand U185 (N_185,In_1192,In_1609);
nor U186 (N_186,In_714,In_415);
nor U187 (N_187,In_279,In_804);
and U188 (N_188,In_425,In_1768);
nand U189 (N_189,In_1079,In_1500);
nor U190 (N_190,In_989,In_436);
nand U191 (N_191,In_286,In_716);
nand U192 (N_192,In_1072,In_1093);
nand U193 (N_193,In_739,In_1942);
and U194 (N_194,In_217,In_400);
xor U195 (N_195,In_1863,In_992);
nand U196 (N_196,In_1633,In_1094);
and U197 (N_197,In_1590,In_216);
nor U198 (N_198,In_314,In_236);
nand U199 (N_199,In_502,In_1897);
nand U200 (N_200,In_858,In_806);
nand U201 (N_201,N_101,In_210);
and U202 (N_202,In_1810,In_1952);
nor U203 (N_203,In_782,In_1837);
and U204 (N_204,In_580,In_1933);
nor U205 (N_205,In_535,In_610);
nand U206 (N_206,N_3,In_121);
nand U207 (N_207,In_1184,In_1426);
nand U208 (N_208,In_1923,In_1543);
or U209 (N_209,In_1466,In_111);
nor U210 (N_210,In_1759,In_936);
or U211 (N_211,In_1051,In_173);
xor U212 (N_212,N_57,In_152);
nor U213 (N_213,In_1972,In_854);
and U214 (N_214,In_1230,In_1349);
nand U215 (N_215,In_868,In_1867);
xnor U216 (N_216,In_413,In_1741);
nand U217 (N_217,In_1945,In_1431);
or U218 (N_218,In_1257,In_768);
nor U219 (N_219,In_1966,In_391);
nor U220 (N_220,In_812,In_3);
nand U221 (N_221,In_885,In_791);
and U222 (N_222,In_407,N_41);
nand U223 (N_223,In_770,In_698);
xnor U224 (N_224,In_1570,In_1540);
or U225 (N_225,In_440,In_816);
nor U226 (N_226,In_1895,In_790);
nor U227 (N_227,N_81,In_282);
and U228 (N_228,In_1150,In_1535);
or U229 (N_229,In_1212,In_1820);
xor U230 (N_230,In_1593,In_5);
nor U231 (N_231,In_385,In_1670);
or U232 (N_232,In_141,In_807);
or U233 (N_233,In_1887,In_1384);
nand U234 (N_234,In_1935,In_471);
nor U235 (N_235,In_339,In_300);
and U236 (N_236,In_426,In_758);
and U237 (N_237,In_151,In_11);
and U238 (N_238,In_1009,In_1224);
nor U239 (N_239,N_30,In_122);
and U240 (N_240,In_839,In_693);
and U241 (N_241,In_389,In_834);
nand U242 (N_242,In_624,N_20);
nor U243 (N_243,In_449,In_475);
or U244 (N_244,N_168,In_477);
or U245 (N_245,N_129,In_1817);
nand U246 (N_246,N_159,In_1165);
and U247 (N_247,In_1164,In_77);
nor U248 (N_248,N_87,In_281);
or U249 (N_249,In_1434,In_898);
xnor U250 (N_250,In_551,In_1971);
and U251 (N_251,In_1160,In_1797);
or U252 (N_252,In_918,In_1446);
nand U253 (N_253,In_1770,In_143);
nand U254 (N_254,In_1187,In_672);
xnor U255 (N_255,In_1898,In_1112);
nand U256 (N_256,In_725,In_1854);
nor U257 (N_257,In_711,In_1437);
or U258 (N_258,In_589,In_1208);
and U259 (N_259,In_567,In_40);
nor U260 (N_260,In_1875,In_224);
nand U261 (N_261,N_74,In_1649);
or U262 (N_262,N_122,In_576);
and U263 (N_263,In_301,In_582);
xnor U264 (N_264,In_377,In_588);
nand U265 (N_265,In_1979,In_1147);
or U266 (N_266,In_565,In_1166);
and U267 (N_267,In_586,In_1376);
or U268 (N_268,In_1056,In_548);
nand U269 (N_269,N_147,In_1319);
nor U270 (N_270,N_26,In_1665);
xnor U271 (N_271,In_439,In_95);
xor U272 (N_272,In_578,In_1508);
nor U273 (N_273,In_1533,In_952);
and U274 (N_274,In_1389,In_69);
nor U275 (N_275,In_1402,N_75);
or U276 (N_276,In_1240,In_1428);
and U277 (N_277,In_1909,In_1120);
nand U278 (N_278,In_700,In_771);
nand U279 (N_279,N_136,In_1678);
or U280 (N_280,In_1641,N_175);
nand U281 (N_281,In_996,N_5);
and U282 (N_282,In_757,In_596);
or U283 (N_283,In_1838,In_1599);
xor U284 (N_284,In_207,In_682);
nor U285 (N_285,In_176,In_1211);
xor U286 (N_286,In_847,In_1233);
or U287 (N_287,In_1845,In_1297);
xor U288 (N_288,In_1791,In_1198);
or U289 (N_289,In_1499,In_1695);
xnor U290 (N_290,N_16,In_1354);
and U291 (N_291,In_99,In_438);
or U292 (N_292,In_1219,In_140);
nor U293 (N_293,In_387,In_1400);
nor U294 (N_294,In_189,In_1513);
nor U295 (N_295,In_512,In_546);
xnor U296 (N_296,In_593,In_1778);
nor U297 (N_297,In_911,In_994);
nor U298 (N_298,In_699,In_361);
or U299 (N_299,In_1186,In_1138);
nor U300 (N_300,In_67,In_1194);
xor U301 (N_301,In_999,N_47);
nand U302 (N_302,In_1227,In_1255);
or U303 (N_303,In_1877,In_493);
or U304 (N_304,In_609,In_1322);
nor U305 (N_305,In_1393,In_1397);
and U306 (N_306,In_844,In_653);
or U307 (N_307,In_356,In_163);
and U308 (N_308,In_1295,In_1637);
nor U309 (N_309,In_75,In_1950);
and U310 (N_310,In_1723,In_947);
or U311 (N_311,N_148,In_1926);
nor U312 (N_312,In_937,In_290);
nand U313 (N_313,In_1145,In_1643);
and U314 (N_314,In_941,In_1067);
nand U315 (N_315,N_111,In_1804);
nor U316 (N_316,In_206,In_730);
and U317 (N_317,In_16,In_1457);
nor U318 (N_318,In_327,In_1454);
xor U319 (N_319,In_845,In_135);
or U320 (N_320,In_919,In_940);
and U321 (N_321,In_55,N_141);
nand U322 (N_322,In_867,N_116);
nand U323 (N_323,In_649,N_82);
nand U324 (N_324,In_1792,In_694);
nor U325 (N_325,In_1752,In_1162);
xnor U326 (N_326,In_1279,N_162);
or U327 (N_327,In_1490,In_875);
nand U328 (N_328,In_848,In_1308);
nor U329 (N_329,In_241,In_935);
or U330 (N_330,In_1179,In_1365);
or U331 (N_331,In_1125,In_951);
or U332 (N_332,In_1246,In_1141);
nand U333 (N_333,In_1175,N_151);
and U334 (N_334,N_135,In_1475);
nor U335 (N_335,In_486,In_1688);
xnor U336 (N_336,In_1869,In_456);
xnor U337 (N_337,In_566,N_163);
nand U338 (N_338,In_675,In_909);
and U339 (N_339,In_230,In_1415);
xor U340 (N_340,In_736,In_931);
nand U341 (N_341,In_1653,In_248);
xor U342 (N_342,In_1028,In_1323);
and U343 (N_343,In_1704,N_23);
and U344 (N_344,In_1301,In_1524);
or U345 (N_345,N_8,In_913);
xnor U346 (N_346,In_1756,In_406);
xor U347 (N_347,N_43,In_1698);
or U348 (N_348,In_1152,In_1554);
nand U349 (N_349,In_63,In_1451);
nand U350 (N_350,In_647,In_1256);
nand U351 (N_351,In_1767,In_84);
nand U352 (N_352,In_442,In_1060);
and U353 (N_353,In_1202,In_1161);
and U354 (N_354,In_805,In_1455);
xnor U355 (N_355,In_1310,In_1630);
nand U356 (N_356,In_1098,In_444);
xnor U357 (N_357,In_1151,In_779);
or U358 (N_358,In_538,In_1879);
xnor U359 (N_359,In_213,In_1861);
and U360 (N_360,In_1581,In_772);
and U361 (N_361,In_1463,In_448);
xor U362 (N_362,In_743,In_533);
xnor U363 (N_363,In_394,In_1077);
nand U364 (N_364,In_1799,In_1625);
nor U365 (N_365,In_61,N_72);
xnor U366 (N_366,In_1065,N_67);
xnor U367 (N_367,In_1846,In_969);
or U368 (N_368,In_1763,In_840);
nand U369 (N_369,In_1385,In_1833);
xor U370 (N_370,In_1731,In_405);
and U371 (N_371,In_223,In_1561);
nor U372 (N_372,N_139,In_873);
and U373 (N_373,In_464,In_632);
and U374 (N_374,In_291,In_1865);
or U375 (N_375,In_172,In_467);
and U376 (N_376,N_51,In_49);
or U377 (N_377,In_1712,In_520);
xor U378 (N_378,In_1911,In_659);
nand U379 (N_379,In_1505,In_190);
or U380 (N_380,In_554,In_1087);
nor U381 (N_381,In_280,In_354);
nor U382 (N_382,In_1527,In_1074);
and U383 (N_383,In_1276,In_975);
nand U384 (N_384,N_54,In_1487);
nand U385 (N_385,In_1265,In_1871);
or U386 (N_386,In_729,In_1410);
xnor U387 (N_387,In_979,In_403);
nand U388 (N_388,In_1274,In_1564);
and U389 (N_389,In_1858,In_789);
nand U390 (N_390,In_473,In_1521);
nor U391 (N_391,In_1586,In_948);
or U392 (N_392,In_1225,In_1951);
nor U393 (N_393,N_45,N_113);
nand U394 (N_394,In_530,In_1509);
nor U395 (N_395,In_1022,In_1900);
and U396 (N_396,N_83,In_1070);
xor U397 (N_397,N_104,In_1580);
or U398 (N_398,In_1041,In_1055);
xnor U399 (N_399,In_1657,In_479);
and U400 (N_400,N_374,In_543);
or U401 (N_401,In_78,In_1850);
and U402 (N_402,In_1377,In_1461);
and U403 (N_403,In_1631,In_964);
and U404 (N_404,In_108,In_27);
nor U405 (N_405,In_1371,In_1260);
nor U406 (N_406,In_268,N_367);
or U407 (N_407,In_171,N_256);
nor U408 (N_408,In_583,In_341);
nand U409 (N_409,In_1730,In_295);
and U410 (N_410,In_641,N_36);
xnor U411 (N_411,In_342,N_250);
or U412 (N_412,In_1242,N_290);
nor U413 (N_413,In_967,In_334);
nor U414 (N_414,In_830,In_869);
nor U415 (N_415,In_1243,N_262);
xnor U416 (N_416,In_1550,In_1545);
xor U417 (N_417,In_1082,In_1855);
or U418 (N_418,In_1414,In_703);
and U419 (N_419,N_114,In_1266);
xnor U420 (N_420,N_259,In_525);
and U421 (N_421,N_121,In_1221);
nand U422 (N_422,In_965,In_1190);
and U423 (N_423,In_876,In_1497);
and U424 (N_424,N_146,In_508);
and U425 (N_425,In_560,In_1283);
nand U426 (N_426,N_124,In_20);
or U427 (N_427,In_1849,N_382);
nand U428 (N_428,N_119,In_1241);
nor U429 (N_429,N_272,In_841);
nor U430 (N_430,N_98,In_1563);
and U431 (N_431,In_797,In_1489);
nand U432 (N_432,In_52,In_1961);
xor U433 (N_433,N_219,In_1525);
nand U434 (N_434,In_749,In_597);
nand U435 (N_435,In_1938,In_212);
nand U436 (N_436,In_1292,In_1424);
nor U437 (N_437,In_755,In_252);
xnor U438 (N_438,N_69,In_1367);
or U439 (N_439,N_246,In_1956);
nor U440 (N_440,In_1318,In_506);
nor U441 (N_441,In_203,In_267);
nor U442 (N_442,N_34,N_49);
nand U443 (N_443,In_763,In_411);
nand U444 (N_444,N_126,In_1526);
and U445 (N_445,In_1516,In_824);
nor U446 (N_446,In_1477,In_1953);
xor U447 (N_447,N_318,In_170);
xor U448 (N_448,N_174,In_910);
xnor U449 (N_449,In_623,In_409);
and U450 (N_450,In_90,In_655);
nand U451 (N_451,In_357,In_1391);
or U452 (N_452,In_1793,In_60);
nor U453 (N_453,N_302,In_518);
nor U454 (N_454,In_1929,In_459);
and U455 (N_455,In_835,N_360);
nor U456 (N_456,In_572,N_120);
or U457 (N_457,In_829,In_1568);
nor U458 (N_458,In_1114,In_93);
xor U459 (N_459,In_1789,In_159);
or U460 (N_460,In_434,In_1628);
nor U461 (N_461,In_249,In_1713);
or U462 (N_462,In_924,In_278);
nor U463 (N_463,In_1201,In_1049);
nor U464 (N_464,N_153,In_1905);
and U465 (N_465,In_1960,N_252);
or U466 (N_466,In_1553,In_169);
nor U467 (N_467,In_1036,In_401);
and U468 (N_468,In_1034,In_1313);
nand U469 (N_469,N_388,In_162);
and U470 (N_470,In_1685,In_723);
and U471 (N_471,In_820,In_575);
nor U472 (N_472,In_136,In_1404);
or U473 (N_473,In_420,N_39);
or U474 (N_474,In_220,N_398);
nand U475 (N_475,In_792,N_276);
nand U476 (N_476,In_117,In_1725);
or U477 (N_477,In_1614,In_1997);
xnor U478 (N_478,N_229,In_1504);
and U479 (N_479,In_1656,In_810);
or U480 (N_480,N_341,In_366);
and U481 (N_481,In_1335,In_375);
or U482 (N_482,In_945,In_1142);
xor U483 (N_483,In_686,In_1269);
or U484 (N_484,In_987,N_257);
and U485 (N_485,In_1616,In_1206);
nor U486 (N_486,In_296,In_1995);
nand U487 (N_487,In_1133,N_233);
nand U488 (N_488,In_392,In_6);
nor U489 (N_489,N_220,In_1172);
xnor U490 (N_490,In_718,In_240);
nor U491 (N_491,In_1937,In_865);
nor U492 (N_492,In_1118,In_1751);
or U493 (N_493,In_1405,In_1345);
or U494 (N_494,N_183,In_1005);
and U495 (N_495,In_1156,In_1693);
or U496 (N_496,In_1248,In_1618);
xnor U497 (N_497,In_21,In_1796);
xnor U498 (N_498,In_638,N_210);
nor U499 (N_499,In_1886,In_997);
xor U500 (N_500,In_670,In_1531);
nand U501 (N_501,In_1959,In_19);
xor U502 (N_502,In_36,In_1573);
xnor U503 (N_503,In_1032,In_82);
and U504 (N_504,In_432,In_325);
nor U505 (N_505,In_1176,In_956);
and U506 (N_506,In_922,In_251);
xor U507 (N_507,In_1182,In_1111);
nand U508 (N_508,In_1673,In_1541);
and U509 (N_509,In_644,In_149);
or U510 (N_510,N_95,In_679);
and U511 (N_511,N_66,In_476);
nor U512 (N_512,N_369,In_1718);
nor U513 (N_513,N_53,In_1824);
nand U514 (N_514,N_191,In_904);
xnor U515 (N_515,N_325,N_64);
or U516 (N_516,In_1249,In_1889);
or U517 (N_517,In_1916,In_112);
and U518 (N_518,In_1289,N_306);
nand U519 (N_519,In_1291,N_312);
and U520 (N_520,N_371,In_1928);
and U521 (N_521,In_787,In_1530);
nand U522 (N_522,N_32,In_1583);
xnor U523 (N_523,In_1510,In_441);
xor U524 (N_524,In_1433,In_1629);
nor U525 (N_525,In_663,In_1816);
xnor U526 (N_526,In_139,In_1728);
nor U527 (N_527,In_1261,N_389);
or U528 (N_528,N_133,In_929);
xnor U529 (N_529,In_1383,N_329);
nor U530 (N_530,In_595,In_1103);
nor U531 (N_531,In_1904,In_1126);
nor U532 (N_532,In_1514,N_173);
nor U533 (N_533,In_1337,N_157);
nor U534 (N_534,In_304,N_377);
and U535 (N_535,N_327,In_1623);
nor U536 (N_536,In_600,N_283);
and U537 (N_537,In_692,N_364);
and U538 (N_538,In_900,In_219);
xnor U539 (N_539,In_1267,N_6);
xor U540 (N_540,N_340,In_526);
nand U541 (N_541,In_1908,In_1134);
nand U542 (N_542,In_1010,In_131);
nand U543 (N_543,In_1394,In_1692);
nand U544 (N_544,In_1566,N_260);
xor U545 (N_545,In_1474,In_1203);
and U546 (N_546,In_1476,N_131);
and U547 (N_547,N_339,N_76);
nand U548 (N_548,In_962,N_336);
and U549 (N_549,In_1851,In_1982);
or U550 (N_550,N_170,In_302);
nand U551 (N_551,In_155,N_237);
nand U552 (N_552,In_1102,In_1326);
nand U553 (N_553,In_259,In_1131);
and U554 (N_554,In_244,In_1572);
and U555 (N_555,In_1684,N_305);
and U556 (N_556,In_423,N_228);
xor U557 (N_557,In_195,In_397);
nand U558 (N_558,In_246,In_1023);
or U559 (N_559,In_50,In_550);
or U560 (N_560,In_1092,In_619);
nand U561 (N_561,In_1907,N_285);
xor U562 (N_562,In_671,In_1903);
or U563 (N_563,N_60,In_1320);
xnor U564 (N_564,In_914,In_1470);
nand U565 (N_565,N_94,In_1024);
and U566 (N_566,In_1597,N_282);
or U567 (N_567,In_995,In_299);
nor U568 (N_568,N_197,In_233);
nand U569 (N_569,N_11,In_1661);
and U570 (N_570,N_299,In_454);
nand U571 (N_571,In_1465,In_1046);
xor U572 (N_572,N_314,N_212);
and U573 (N_573,In_1336,In_976);
xnor U574 (N_574,In_466,N_373);
or U575 (N_575,N_99,In_1450);
nor U576 (N_576,In_1204,In_1726);
or U577 (N_577,In_556,In_926);
or U578 (N_578,In_1610,In_1001);
or U579 (N_579,In_1798,In_871);
and U580 (N_580,In_607,In_1775);
nand U581 (N_581,In_183,In_1293);
nand U582 (N_582,In_972,In_1228);
nor U583 (N_583,In_437,In_1485);
xor U584 (N_584,In_895,In_1494);
xnor U585 (N_585,In_1117,In_381);
nand U586 (N_586,In_365,In_1441);
xor U587 (N_587,In_581,In_1710);
nand U588 (N_588,In_1574,In_1978);
or U589 (N_589,In_544,In_1146);
xnor U590 (N_590,In_1122,N_397);
nand U591 (N_591,N_350,In_1697);
nand U592 (N_592,In_1795,In_1216);
and U593 (N_593,In_1640,In_618);
and U594 (N_594,In_1381,In_1235);
or U595 (N_595,In_534,In_1408);
nand U596 (N_596,In_850,In_1472);
xnor U597 (N_597,In_1449,N_203);
and U598 (N_598,In_1757,In_484);
nor U599 (N_599,In_1552,In_887);
or U600 (N_600,In_1936,N_442);
nor U601 (N_601,N_491,In_320);
and U602 (N_602,In_181,N_546);
or U603 (N_603,In_28,In_982);
or U604 (N_604,In_1922,N_19);
and U605 (N_605,In_1671,In_541);
xor U606 (N_606,N_239,In_1750);
xor U607 (N_607,N_355,In_1947);
xor U608 (N_608,N_561,In_1679);
and U609 (N_609,N_278,N_15);
or U610 (N_610,In_1732,In_1674);
nor U611 (N_611,In_1471,In_775);
nand U612 (N_612,In_1921,N_536);
nor U613 (N_613,N_255,In_416);
and U614 (N_614,In_604,In_934);
nand U615 (N_615,In_174,N_198);
and U616 (N_616,In_114,N_96);
and U617 (N_617,In_331,In_1129);
and U618 (N_618,N_380,N_310);
xor U619 (N_619,In_643,In_182);
and U620 (N_620,In_1215,In_1358);
or U621 (N_621,N_24,In_380);
or U622 (N_622,N_164,In_417);
or U623 (N_623,In_932,N_109);
or U624 (N_624,In_1802,In_684);
or U625 (N_625,In_1720,N_292);
nor U626 (N_626,In_1914,In_185);
nor U627 (N_627,In_214,N_460);
nor U628 (N_628,In_1003,In_793);
nor U629 (N_629,N_184,In_1829);
xnor U630 (N_630,N_161,In_158);
nor U631 (N_631,In_545,In_1881);
nor U632 (N_632,In_148,N_416);
xor U633 (N_633,N_345,In_1964);
nor U634 (N_634,N_531,N_232);
nand U635 (N_635,In_1761,In_1719);
nor U636 (N_636,In_1589,In_823);
and U637 (N_637,N_488,In_1137);
xnor U638 (N_638,In_731,N_293);
nor U639 (N_639,In_650,N_65);
nor U640 (N_640,In_1234,N_456);
nand U641 (N_641,N_200,N_202);
nand U642 (N_642,In_1305,N_201);
xor U643 (N_643,N_171,In_180);
and U644 (N_644,In_1567,In_234);
nand U645 (N_645,In_1205,N_527);
or U646 (N_646,In_1075,N_273);
and U647 (N_647,In_1037,N_245);
nand U648 (N_648,In_1350,In_1090);
nor U649 (N_649,In_986,In_1396);
xnor U650 (N_650,In_568,In_1724);
nor U651 (N_651,In_1747,In_352);
or U652 (N_652,In_1740,N_489);
nand U653 (N_653,In_87,In_886);
nand U654 (N_654,In_1207,In_184);
nor U655 (N_655,In_1549,N_482);
nand U656 (N_656,N_401,N_529);
nand U657 (N_657,In_1577,In_1379);
nor U658 (N_658,In_1058,N_266);
and U659 (N_659,In_1876,In_1946);
and U660 (N_660,In_724,N_549);
nand U661 (N_661,In_1168,N_169);
nand U662 (N_662,In_127,N_180);
or U663 (N_663,In_1443,In_372);
nand U664 (N_664,In_1066,N_408);
xor U665 (N_665,N_461,N_18);
and U666 (N_666,In_1558,In_1502);
or U667 (N_667,N_365,N_97);
nor U668 (N_668,In_1154,In_198);
xor U669 (N_669,N_132,In_1666);
xor U670 (N_670,In_1737,In_1664);
and U671 (N_671,In_1974,N_46);
xnor U672 (N_672,In_744,In_1311);
or U673 (N_673,N_386,In_784);
nor U674 (N_674,In_621,In_599);
or U675 (N_675,N_21,N_300);
and U676 (N_676,In_1325,In_637);
and U677 (N_677,In_794,In_1140);
and U678 (N_678,In_376,N_196);
and U679 (N_679,N_118,In_635);
or U680 (N_680,In_1994,In_1417);
or U681 (N_681,In_1773,N_117);
and U682 (N_682,In_1786,In_1860);
xor U683 (N_683,N_79,In_1456);
nand U684 (N_684,In_450,In_667);
nand U685 (N_685,N_486,N_599);
or U686 (N_686,In_1764,In_1327);
nor U687 (N_687,In_288,In_1444);
nand U688 (N_688,In_1467,N_458);
nand U689 (N_689,In_9,In_1644);
xor U690 (N_690,N_275,In_124);
nor U691 (N_691,In_1333,In_1555);
or U692 (N_692,In_879,In_1076);
xor U693 (N_693,In_957,N_213);
xnor U694 (N_694,In_1421,N_361);
or U695 (N_695,N_195,In_832);
or U696 (N_696,N_414,In_1984);
nor U697 (N_697,In_1442,N_501);
xnor U698 (N_698,In_990,In_1018);
and U699 (N_699,In_404,N_223);
nand U700 (N_700,In_1086,N_315);
and U701 (N_701,In_1464,In_310);
xnor U702 (N_702,N_512,In_496);
xor U703 (N_703,In_83,N_466);
nand U704 (N_704,In_1766,In_1386);
xor U705 (N_705,N_281,N_391);
or U706 (N_706,N_483,N_515);
nor U707 (N_707,N_485,In_1647);
or U708 (N_708,In_367,In_1388);
nand U709 (N_709,N_346,N_286);
nand U710 (N_710,N_14,N_586);
nor U711 (N_711,N_565,In_51);
and U712 (N_712,N_418,In_883);
nand U713 (N_713,N_500,N_592);
or U714 (N_714,In_516,In_1375);
and U715 (N_715,In_318,In_1011);
and U716 (N_716,In_1498,In_1401);
and U717 (N_717,N_574,N_384);
and U718 (N_718,In_89,N_73);
or U719 (N_719,In_1068,N_436);
and U720 (N_720,N_509,In_165);
nor U721 (N_721,N_199,In_1296);
and U722 (N_722,In_1681,N_508);
or U723 (N_723,N_226,In_460);
or U724 (N_724,In_594,In_706);
xnor U725 (N_725,In_371,N_392);
xnor U726 (N_726,In_1015,N_63);
nand U727 (N_727,In_892,N_569);
xor U728 (N_728,In_1236,In_305);
or U729 (N_729,In_1217,In_1536);
xnor U730 (N_730,In_255,In_1432);
and U731 (N_731,In_1170,In_685);
xor U732 (N_732,In_673,In_1998);
or U733 (N_733,In_197,N_28);
nor U734 (N_734,In_1299,In_558);
and U735 (N_735,In_452,In_487);
or U736 (N_736,In_258,In_1344);
xor U737 (N_737,N_143,In_591);
xnor U738 (N_738,In_396,In_144);
xor U739 (N_739,N_449,In_262);
and U740 (N_740,In_579,N_425);
nor U741 (N_741,N_152,In_1548);
xnor U742 (N_742,In_966,N_274);
nand U743 (N_743,In_943,In_1701);
nand U744 (N_744,In_1989,In_1883);
nor U745 (N_745,In_480,In_584);
nor U746 (N_746,N_231,N_59);
xnor U747 (N_747,In_1314,In_453);
xor U748 (N_748,In_767,N_597);
nand U749 (N_749,N_484,N_535);
or U750 (N_750,In_469,In_294);
and U751 (N_751,In_433,In_150);
xnor U752 (N_752,In_1715,N_593);
and U753 (N_753,In_704,In_881);
nand U754 (N_754,In_1705,In_362);
nor U755 (N_755,In_1714,In_1357);
nor U756 (N_756,In_627,In_421);
or U757 (N_757,In_1760,N_379);
or U758 (N_758,In_81,In_1270);
nand U759 (N_759,N_473,N_333);
xor U760 (N_760,In_18,In_1987);
or U761 (N_761,In_802,N_303);
xnor U762 (N_762,In_1650,In_1576);
nand U763 (N_763,In_373,In_1912);
xor U764 (N_764,In_1537,In_187);
nand U765 (N_765,In_1668,In_803);
or U766 (N_766,In_674,N_313);
nor U767 (N_767,N_61,N_230);
or U768 (N_768,N_440,N_1);
or U769 (N_769,In_991,In_639);
and U770 (N_770,In_7,In_1059);
and U771 (N_771,In_1944,In_1030);
and U772 (N_772,In_783,In_323);
nor U773 (N_773,N_410,N_538);
nand U774 (N_774,In_1790,In_98);
nor U775 (N_775,In_1480,In_1983);
or U776 (N_776,In_156,N_324);
nand U777 (N_777,N_514,N_428);
nor U778 (N_778,In_128,In_1707);
and U779 (N_779,In_499,In_1407);
nand U780 (N_780,N_296,In_1171);
xnor U781 (N_781,In_1940,In_1069);
nand U782 (N_782,In_1210,In_710);
or U783 (N_783,N_585,In_1181);
nand U784 (N_784,In_161,In_483);
nand U785 (N_785,N_172,In_1986);
xnor U786 (N_786,In_57,In_324);
nor U787 (N_787,N_205,In_1615);
xnor U788 (N_788,N_443,N_552);
nand U789 (N_789,In_1334,In_1655);
and U790 (N_790,N_258,N_511);
nand U791 (N_791,In_1061,In_1985);
and U792 (N_792,In_1478,N_497);
and U793 (N_793,N_309,In_1116);
xor U794 (N_794,N_142,N_447);
and U795 (N_795,In_66,In_1780);
or U796 (N_796,In_1083,In_289);
nor U797 (N_797,In_1556,In_1862);
and U798 (N_798,In_916,N_470);
nor U799 (N_799,N_331,N_513);
nor U800 (N_800,N_603,In_656);
or U801 (N_801,In_857,In_1965);
xnor U802 (N_802,In_322,In_1064);
nor U803 (N_803,In_961,N_187);
nand U804 (N_804,In_1777,In_1264);
nor U805 (N_805,In_424,In_1607);
and U806 (N_806,N_799,In_613);
xor U807 (N_807,In_308,N_754);
xnor U808 (N_808,In_1021,In_37);
nor U809 (N_809,In_1220,N_682);
xor U810 (N_810,In_606,N_643);
xnor U811 (N_811,In_836,N_780);
xnor U812 (N_812,N_718,In_843);
nand U813 (N_813,N_317,N_158);
nor U814 (N_814,In_1369,In_1153);
or U815 (N_815,In_501,In_1520);
or U816 (N_816,N_641,In_1084);
or U817 (N_817,N_323,In_1452);
nor U818 (N_818,In_1339,N_676);
nand U819 (N_819,In_738,In_513);
xor U820 (N_820,N_459,In_928);
xor U821 (N_821,In_1284,N_58);
nand U822 (N_822,In_1027,N_782);
nand U823 (N_823,N_798,In_664);
and U824 (N_824,In_1702,In_455);
nand U825 (N_825,In_1330,In_611);
nand U826 (N_826,In_1809,In_39);
or U827 (N_827,In_874,In_1831);
xor U828 (N_828,In_833,In_227);
xor U829 (N_829,N_745,N_400);
and U830 (N_830,In_1254,In_1980);
and U831 (N_831,In_1981,In_1528);
nor U832 (N_832,In_10,N_249);
or U833 (N_833,In_276,In_1917);
and U834 (N_834,In_1196,N_144);
xnor U835 (N_835,In_398,In_1636);
nor U836 (N_836,In_42,N_269);
and U837 (N_837,In_1351,In_355);
nor U838 (N_838,N_337,In_1360);
and U839 (N_839,In_798,In_616);
or U840 (N_840,N_759,In_862);
nor U841 (N_841,N_4,N_127);
nor U842 (N_842,In_1237,In_1419);
nand U843 (N_843,In_661,N_771);
or U844 (N_844,N_476,N_85);
xor U845 (N_845,N_478,In_984);
nor U846 (N_846,In_1519,N_580);
nand U847 (N_847,In_1557,In_1309);
and U848 (N_848,In_1169,In_14);
nor U849 (N_849,In_1547,In_1387);
and U850 (N_850,N_698,In_226);
or U851 (N_851,In_1748,N_541);
nor U852 (N_852,N_446,N_721);
nand U853 (N_853,In_681,In_468);
or U854 (N_854,In_72,In_1263);
xor U855 (N_855,N_645,N_222);
nand U856 (N_856,In_1949,In_602);
nor U857 (N_857,N_432,In_1648);
or U858 (N_858,In_866,In_923);
and U859 (N_859,N_110,N_368);
xnor U860 (N_860,N_362,N_669);
xor U861 (N_861,In_1807,N_668);
nor U862 (N_862,N_50,N_722);
and U863 (N_863,In_363,In_1495);
nor U864 (N_864,In_378,N_507);
nand U865 (N_865,In_1755,N_777);
xnor U866 (N_866,N_680,N_247);
xnor U867 (N_867,In_985,In_1238);
xor U868 (N_868,In_1331,In_1275);
nor U869 (N_869,N_685,N_767);
nor U870 (N_870,N_494,N_701);
and U871 (N_871,N_402,N_215);
xor U872 (N_872,In_1409,In_1893);
xnor U873 (N_873,N_291,In_1611);
and U874 (N_874,In_884,N_618);
nand U875 (N_875,In_1302,In_382);
nor U876 (N_876,In_1031,In_429);
nand U877 (N_877,In_614,N_123);
nand U878 (N_878,N_248,In_838);
nor U879 (N_879,N_559,In_113);
or U880 (N_880,N_467,In_179);
or U881 (N_881,N_630,In_1352);
xnor U882 (N_882,N_613,N_308);
xor U883 (N_883,N_797,In_1801);
nor U884 (N_884,In_1321,N_453);
or U885 (N_885,N_385,In_933);
xnor U886 (N_886,N_638,In_1539);
nand U887 (N_887,In_851,In_1993);
xor U888 (N_888,N_720,In_759);
or U889 (N_889,In_43,In_773);
and U890 (N_890,N_40,N_394);
xor U891 (N_891,In_1448,In_1411);
xor U892 (N_892,In_1735,In_1769);
and U893 (N_893,In_1342,N_294);
or U894 (N_894,In_585,N_156);
nand U895 (N_895,In_292,N_241);
nor U896 (N_896,N_335,N_567);
nor U897 (N_897,In_1035,In_1420);
nand U898 (N_898,In_776,N_37);
and U899 (N_899,In_1753,N_715);
or U900 (N_900,N_526,In_1012);
and U901 (N_901,In_1973,N_713);
and U902 (N_902,N_737,In_668);
nor U903 (N_903,In_264,In_1627);
and U904 (N_904,In_1008,N_457);
xnor U905 (N_905,N_739,In_1288);
nor U906 (N_906,N_522,In_263);
and U907 (N_907,N_700,N_288);
nor U908 (N_908,In_1828,N_752);
nand U909 (N_909,In_80,N_743);
nor U910 (N_910,N_594,N_562);
or U911 (N_911,N_463,In_1085);
xnor U912 (N_912,N_105,N_22);
and U913 (N_913,N_93,In_56);
or U914 (N_914,N_675,N_591);
nand U915 (N_915,N_776,In_1931);
nor U916 (N_916,In_864,In_1736);
nor U917 (N_917,N_650,N_581);
nand U918 (N_918,N_640,N_542);
and U919 (N_919,In_1468,In_1841);
or U920 (N_920,N_658,In_1106);
xor U921 (N_921,In_959,In_1304);
and U922 (N_922,In_1806,In_504);
nand U923 (N_923,N_644,N_639);
and U924 (N_924,N_705,N_710);
or U925 (N_925,N_35,In_1638);
nor U926 (N_926,N_176,In_1306);
xnor U927 (N_927,In_1459,In_1717);
nand U928 (N_928,N_381,N_423);
nand U929 (N_929,N_55,In_1239);
xnor U930 (N_930,In_497,N_793);
nand U931 (N_931,In_1683,In_1913);
nand U932 (N_932,In_443,In_514);
or U933 (N_933,In_1052,N_84);
nor U934 (N_934,In_250,In_132);
and U935 (N_935,N_42,In_1177);
xor U936 (N_936,In_896,In_349);
and U937 (N_937,N_717,In_359);
and U938 (N_938,In_1890,N_544);
nand U939 (N_939,N_86,N_518);
or U940 (N_940,In_285,In_517);
nor U941 (N_941,N_528,N_207);
or U942 (N_942,In_328,In_489);
or U943 (N_943,In_45,In_1632);
xnor U944 (N_944,N_600,In_96);
nor U945 (N_945,In_196,In_690);
xor U946 (N_946,In_971,N_421);
or U947 (N_947,N_383,In_374);
or U948 (N_948,N_90,N_179);
nand U949 (N_949,N_188,N_738);
nand U950 (N_950,In_13,N_697);
nor U951 (N_951,In_32,N_712);
and U952 (N_952,N_563,In_1930);
xor U953 (N_953,In_528,In_574);
nor U954 (N_954,In_1842,In_34);
nand U955 (N_955,N_696,In_307);
xnor U956 (N_956,In_1919,In_715);
or U957 (N_957,N_411,N_289);
and U958 (N_958,In_1822,In_1047);
nand U959 (N_959,In_1779,N_240);
and U960 (N_960,In_822,N_277);
nor U961 (N_961,N_503,N_548);
xor U962 (N_962,In_1097,In_801);
or U963 (N_963,N_224,In_1130);
xor U964 (N_964,In_175,N_612);
xor U965 (N_965,N_674,N_455);
nand U966 (N_966,In_277,In_1902);
xnor U967 (N_967,N_468,N_637);
or U968 (N_968,N_590,N_615);
nor U969 (N_969,In_178,N_130);
and U970 (N_970,N_322,In_687);
or U971 (N_971,In_1645,In_465);
nand U972 (N_972,N_298,N_417);
and U973 (N_973,In_1812,In_1873);
xnor U974 (N_974,N_504,In_1639);
xnor U975 (N_975,In_215,N_753);
nand U976 (N_976,In_298,N_452);
or U977 (N_977,In_1948,N_564);
or U978 (N_978,In_1696,N_741);
and U979 (N_979,In_1017,N_795);
or U980 (N_980,N_787,In_1927);
xnor U981 (N_981,N_573,N_422);
or U982 (N_982,N_242,In_1746);
nand U983 (N_983,N_655,In_142);
xor U984 (N_984,In_333,In_47);
nor U985 (N_985,In_1231,In_137);
xor U986 (N_986,N_347,N_631);
nor U987 (N_987,N_372,N_311);
or U988 (N_988,In_1634,N_642);
xor U989 (N_989,In_1346,N_540);
or U990 (N_990,N_789,In_1348);
nand U991 (N_991,N_791,In_677);
and U992 (N_992,N_464,In_970);
nor U993 (N_993,In_192,N_44);
nand U994 (N_994,N_543,N_7);
nand U995 (N_995,N_693,In_603);
xor U996 (N_996,In_719,In_917);
and U997 (N_997,N_0,N_607);
nand U998 (N_998,N_667,N_684);
and U999 (N_999,N_583,N_724);
nand U1000 (N_1000,In_726,In_283);
nor U1001 (N_1001,N_971,In_1423);
and U1002 (N_1002,N_778,N_490);
or U1003 (N_1003,In_688,N_946);
or U1004 (N_1004,N_927,N_999);
and U1005 (N_1005,N_403,In_1800);
nor U1006 (N_1006,In_1048,N_125);
or U1007 (N_1007,N_608,In_428);
xnor U1008 (N_1008,N_566,N_280);
nor U1009 (N_1009,N_906,N_595);
nor U1010 (N_1010,In_1262,N_839);
and U1011 (N_1011,N_634,In_1095);
nor U1012 (N_1012,In_592,In_1598);
and U1013 (N_1013,In_70,In_626);
and U1014 (N_1014,N_936,N_610);
nor U1015 (N_1015,N_375,N_321);
xnor U1016 (N_1016,N_959,N_395);
xnor U1017 (N_1017,N_284,In_1258);
and U1018 (N_1018,In_272,N_659);
nor U1019 (N_1019,In_1044,N_251);
nor U1020 (N_1020,In_30,N_378);
nand U1021 (N_1021,N_728,In_1781);
nor U1022 (N_1022,N_941,N_429);
and U1023 (N_1023,In_1584,In_882);
xor U1024 (N_1024,N_108,N_965);
and U1025 (N_1025,In_863,In_481);
nand U1026 (N_1026,N_472,In_652);
xnor U1027 (N_1027,In_1691,In_505);
and U1028 (N_1028,In_64,In_261);
xor U1029 (N_1029,In_257,In_752);
xnor U1030 (N_1030,N_227,N_89);
and U1031 (N_1031,N_649,In_58);
or U1032 (N_1032,N_523,N_405);
and U1033 (N_1033,N_920,N_896);
xor U1034 (N_1034,N_584,In_1016);
or U1035 (N_1035,N_194,In_1104);
nor U1036 (N_1036,In_59,In_1285);
xnor U1037 (N_1037,N_942,N_989);
nor U1038 (N_1038,N_923,N_493);
xnor U1039 (N_1039,In_1690,N_596);
nand U1040 (N_1040,In_200,In_1874);
and U1041 (N_1041,N_881,In_570);
nor U1042 (N_1042,N_679,N_747);
xor U1043 (N_1043,N_702,N_623);
xnor U1044 (N_1044,N_761,In_1722);
nand U1045 (N_1045,In_157,In_853);
nor U1046 (N_1046,N_800,In_559);
nor U1047 (N_1047,In_1374,In_1783);
and U1048 (N_1048,N_426,In_601);
nor U1049 (N_1049,In_237,In_1676);
or U1050 (N_1050,N_621,N_474);
nand U1051 (N_1051,In_696,N_268);
nor U1052 (N_1052,In_1143,In_1836);
nor U1053 (N_1053,In_1429,N_860);
nand U1054 (N_1054,N_824,N_577);
or U1055 (N_1055,N_960,N_666);
or U1056 (N_1056,In_747,N_814);
xor U1057 (N_1057,In_1546,N_208);
or U1058 (N_1058,N_415,N_817);
nand U1059 (N_1059,In_1020,In_265);
or U1060 (N_1060,In_62,In_1825);
nand U1061 (N_1061,In_1406,In_239);
and U1062 (N_1062,In_332,In_1493);
or U1063 (N_1063,N_393,In_110);
nand U1064 (N_1064,In_808,In_946);
xnor U1065 (N_1065,In_1045,N_576);
nor U1066 (N_1066,N_165,In_735);
xor U1067 (N_1067,In_1963,In_569);
nand U1068 (N_1068,N_598,In_1899);
or U1069 (N_1069,In_1832,In_1435);
nor U1070 (N_1070,N_626,N_775);
and U1071 (N_1071,N_193,In_1416);
or U1072 (N_1072,N_808,N_844);
nand U1073 (N_1073,N_349,In_1967);
or U1074 (N_1074,In_1214,N_178);
nor U1075 (N_1075,N_270,N_332);
nand U1076 (N_1076,In_1646,N_316);
xnor U1077 (N_1077,In_458,In_1977);
nor U1078 (N_1078,N_972,In_899);
nand U1079 (N_1079,N_980,N_823);
nor U1080 (N_1080,In_482,N_891);
nand U1081 (N_1081,N_636,N_962);
nand U1082 (N_1082,In_105,N_773);
xnor U1083 (N_1083,N_431,In_260);
and U1084 (N_1084,In_1709,In_1868);
nor U1085 (N_1085,N_764,In_973);
or U1086 (N_1086,In_780,N_916);
or U1087 (N_1087,N_547,N_177);
nand U1088 (N_1088,N_751,In_764);
xnor U1089 (N_1089,N_886,In_1088);
nand U1090 (N_1090,N_462,In_1403);
nor U1091 (N_1091,N_516,N_672);
and U1092 (N_1092,N_909,In_557);
xnor U1093 (N_1093,In_938,N_128);
xnor U1094 (N_1094,N_951,In_1253);
and U1095 (N_1095,N_663,N_88);
nor U1096 (N_1096,In_897,In_1039);
nor U1097 (N_1097,In_1819,In_1364);
xor U1098 (N_1098,In_1157,N_520);
or U1099 (N_1099,In_218,N_818);
and U1100 (N_1100,N_678,N_396);
nand U1101 (N_1101,N_654,N_475);
and U1102 (N_1102,N_204,N_708);
nand U1103 (N_1103,N_768,N_847);
or U1104 (N_1104,In_981,N_903);
nand U1105 (N_1105,N_304,In_669);
nor U1106 (N_1106,In_1939,In_494);
or U1107 (N_1107,N_857,N_149);
or U1108 (N_1108,N_870,N_992);
or U1109 (N_1109,In_1604,N_56);
xnor U1110 (N_1110,In_1744,In_48);
and U1111 (N_1111,In_1380,N_52);
and U1112 (N_1112,N_115,N_211);
and U1113 (N_1113,In_701,N_632);
and U1114 (N_1114,In_1534,N_838);
nand U1115 (N_1115,In_147,N_794);
or U1116 (N_1116,In_1338,In_1312);
nor U1117 (N_1117,In_1091,N_216);
nand U1118 (N_1118,In_800,In_35);
nand U1119 (N_1119,N_863,In_523);
nand U1120 (N_1120,N_694,N_225);
and U1121 (N_1121,N_625,In_691);
or U1122 (N_1122,N_167,In_1571);
nor U1123 (N_1123,N_238,N_609);
nor U1124 (N_1124,In_1281,N_709);
nor U1125 (N_1125,In_1469,In_1924);
or U1126 (N_1126,N_107,In_85);
or U1127 (N_1127,N_582,N_970);
or U1128 (N_1128,N_681,In_1882);
nand U1129 (N_1129,In_53,N_555);
or U1130 (N_1130,In_1538,In_1910);
or U1131 (N_1131,N_517,In_1491);
xnor U1132 (N_1132,In_888,N_947);
and U1133 (N_1133,N_888,N_236);
nand U1134 (N_1134,In_1606,In_1511);
or U1135 (N_1135,N_664,N_855);
nand U1136 (N_1136,In_1341,N_894);
and U1137 (N_1137,N_703,N_465);
nor U1138 (N_1138,In_1458,N_840);
nand U1139 (N_1139,N_661,N_437);
and U1140 (N_1140,N_545,N_78);
or U1141 (N_1141,N_723,N_804);
nor U1142 (N_1142,N_802,In_153);
nand U1143 (N_1143,In_134,In_605);
nand U1144 (N_1144,N_487,N_606);
nor U1145 (N_1145,In_1847,In_1901);
and U1146 (N_1146,N_334,N_907);
or U1147 (N_1147,N_558,N_913);
nor U1148 (N_1148,In_1864,N_945);
or U1149 (N_1149,N_189,In_1144);
nor U1150 (N_1150,In_1135,N_779);
and U1151 (N_1151,N_735,In_430);
or U1152 (N_1152,In_1197,In_446);
or U1153 (N_1153,N_77,N_939);
xnor U1154 (N_1154,In_490,In_818);
and U1155 (N_1155,N_969,N_788);
and U1156 (N_1156,N_662,In_562);
and U1157 (N_1157,N_948,N_792);
nor U1158 (N_1158,N_897,In_2);
nor U1159 (N_1159,N_326,In_38);
xnor U1160 (N_1160,N_140,In_1532);
nor U1161 (N_1161,N_689,N_898);
nand U1162 (N_1162,In_1970,In_1195);
nand U1163 (N_1163,N_554,N_448);
xor U1164 (N_1164,In_1811,N_656);
nand U1165 (N_1165,N_351,In_769);
and U1166 (N_1166,N_803,In_1669);
or U1167 (N_1167,N_706,N_390);
xnor U1168 (N_1168,N_235,N_887);
or U1169 (N_1169,N_9,N_961);
nor U1170 (N_1170,In_1575,N_677);
and U1171 (N_1171,N_409,In_1663);
nand U1172 (N_1172,In_1512,In_683);
nor U1173 (N_1173,N_964,In_717);
nor U1174 (N_1174,N_495,N_774);
xor U1175 (N_1175,N_427,N_412);
and U1176 (N_1176,N_27,In_1894);
nor U1177 (N_1177,N_430,In_745);
nor U1178 (N_1178,N_192,N_433);
or U1179 (N_1179,In_379,In_1123);
nand U1180 (N_1180,In_958,N_931);
or U1181 (N_1181,In_1399,N_699);
xnor U1182 (N_1182,In_222,In_1818);
nor U1183 (N_1183,N_805,In_1962);
or U1184 (N_1184,N_810,N_568);
xor U1185 (N_1185,In_732,In_645);
or U1186 (N_1186,N_750,N_653);
and U1187 (N_1187,N_873,N_950);
and U1188 (N_1188,In_1729,In_1745);
or U1189 (N_1189,N_879,N_660);
or U1190 (N_1190,N_704,N_815);
nor U1191 (N_1191,In_221,In_238);
nor U1192 (N_1192,In_894,In_1689);
nor U1193 (N_1193,N_843,N_100);
xor U1194 (N_1194,In_116,In_1483);
nor U1195 (N_1195,N_155,N_762);
nor U1196 (N_1196,In_412,N_628);
nand U1197 (N_1197,In_1099,N_740);
or U1198 (N_1198,In_1918,N_825);
nand U1199 (N_1199,In_316,In_309);
xnor U1200 (N_1200,In_662,N_716);
xnor U1201 (N_1201,N_1142,N_983);
or U1202 (N_1202,N_973,In_386);
nand U1203 (N_1203,N_786,N_530);
nand U1204 (N_1204,In_146,N_892);
nor U1205 (N_1205,N_1032,N_1163);
or U1206 (N_1206,In_266,N_1158);
or U1207 (N_1207,N_1041,N_1164);
and U1208 (N_1208,N_1151,N_861);
nand U1209 (N_1209,N_714,N_866);
nand U1210 (N_1210,N_790,In_1121);
and U1211 (N_1211,N_871,N_1094);
nor U1212 (N_1212,N_1025,N_614);
or U1213 (N_1213,N_243,In_1840);
and U1214 (N_1214,In_1439,N_829);
or U1215 (N_1215,N_998,In_1794);
and U1216 (N_1216,In_1920,N_925);
xor U1217 (N_1217,In_208,N_506);
and U1218 (N_1218,N_890,In_1427);
and U1219 (N_1219,In_74,In_1100);
xnor U1220 (N_1220,N_930,In_1282);
xor U1221 (N_1221,N_244,In_1782);
nor U1222 (N_1222,In_1687,In_872);
nor U1223 (N_1223,In_253,In_1667);
nand U1224 (N_1224,N_985,In_712);
xnor U1225 (N_1225,In_1000,In_1742);
or U1226 (N_1226,N_910,N_917);
nand U1227 (N_1227,N_560,N_1130);
nand U1228 (N_1228,N_1161,N_185);
xor U1229 (N_1229,N_469,N_1181);
or U1230 (N_1230,In_1823,N_885);
xnor U1231 (N_1231,In_870,N_477);
xnor U1232 (N_1232,In_1482,In_1565);
or U1233 (N_1233,N_533,In_33);
nand U1234 (N_1234,N_781,N_982);
xnor U1235 (N_1235,In_761,N_875);
xor U1236 (N_1236,In_571,In_665);
nor U1237 (N_1237,N_977,In_154);
nand U1238 (N_1238,N_218,N_1039);
nand U1239 (N_1239,N_154,In_553);
and U1240 (N_1240,N_1013,N_1004);
and U1241 (N_1241,N_1027,In_905);
and U1242 (N_1242,In_1501,N_749);
or U1243 (N_1243,N_832,In_1373);
or U1244 (N_1244,In_519,N_354);
or U1245 (N_1245,In_720,N_952);
or U1246 (N_1246,In_228,N_624);
xor U1247 (N_1247,N_858,N_765);
nor U1248 (N_1248,N_1033,N_1074);
nand U1249 (N_1249,N_376,N_845);
and U1250 (N_1250,In_1975,N_1186);
nor U1251 (N_1251,N_1005,N_471);
xnor U1252 (N_1252,N_519,In_1167);
nand U1253 (N_1253,N_363,In_1259);
nor U1254 (N_1254,N_1016,N_1169);
xor U1255 (N_1255,N_1185,N_1167);
nor U1256 (N_1256,In_1392,N_611);
and U1257 (N_1257,N_731,N_997);
or U1258 (N_1258,N_1168,N_1179);
or U1259 (N_1259,In_313,In_608);
nor U1260 (N_1260,In_814,N_865);
and U1261 (N_1261,In_102,In_88);
xnor U1262 (N_1262,In_1522,N_1018);
nor U1263 (N_1263,In_86,N_1145);
nor U1264 (N_1264,N_1056,N_550);
or U1265 (N_1265,In_799,In_676);
nor U1266 (N_1266,In_1738,N_880);
nor U1267 (N_1267,N_424,N_719);
nor U1268 (N_1268,N_1117,N_806);
nand U1269 (N_1269,N_994,In_511);
nor U1270 (N_1270,N_134,In_1355);
nand U1271 (N_1271,N_1189,N_1035);
and U1272 (N_1272,N_1177,In_786);
or U1273 (N_1273,N_1159,In_1247);
and U1274 (N_1274,In_532,N_957);
xor U1275 (N_1275,N_1114,N_1007);
xnor U1276 (N_1276,In_1484,N_1196);
nand U1277 (N_1277,N_1090,N_966);
nor U1278 (N_1278,N_1190,In_1019);
nand U1279 (N_1279,N_1023,N_841);
and U1280 (N_1280,In_1108,In_1592);
and U1281 (N_1281,N_1193,In_15);
nand U1282 (N_1282,N_1028,N_1086);
or U1283 (N_1283,In_1109,N_622);
nor U1284 (N_1284,In_615,N_1137);
nand U1285 (N_1285,In_1529,In_746);
xnor U1286 (N_1286,N_1110,N_510);
nor U1287 (N_1287,In_577,N_1104);
nor U1288 (N_1288,In_229,In_109);
nor U1289 (N_1289,In_1158,N_534);
nor U1290 (N_1290,N_1069,N_1132);
and U1291 (N_1291,N_651,N_254);
nand U1292 (N_1292,N_1009,N_103);
or U1293 (N_1293,N_911,N_816);
nand U1294 (N_1294,In_855,N_922);
xor U1295 (N_1295,N_849,N_1043);
and U1296 (N_1296,N_953,In_120);
and U1297 (N_1297,N_974,N_137);
nor U1298 (N_1298,N_859,In_186);
or U1299 (N_1299,N_1065,N_670);
or U1300 (N_1300,N_1107,N_1029);
and U1301 (N_1301,In_1675,N_1122);
or U1302 (N_1302,In_390,In_1361);
xor U1303 (N_1303,In_498,N_297);
and U1304 (N_1304,In_1743,N_968);
nand U1305 (N_1305,N_1140,N_1178);
nor U1306 (N_1306,In_1976,In_1826);
and U1307 (N_1307,In_1562,N_683);
xor U1308 (N_1308,N_29,N_499);
and U1309 (N_1309,N_617,N_742);
nand U1310 (N_1310,In_762,N_665);
nor U1311 (N_1311,N_736,N_1123);
nand U1312 (N_1312,N_963,N_214);
nor U1313 (N_1313,N_579,N_1089);
or U1314 (N_1314,N_206,N_1141);
nor U1315 (N_1315,In_1200,N_353);
nor U1316 (N_1316,N_505,N_1026);
and U1317 (N_1317,N_872,N_406);
xor U1318 (N_1318,N_571,N_221);
nand U1319 (N_1319,N_1152,N_842);
nand U1320 (N_1320,In_942,N_846);
nor U1321 (N_1321,In_1954,In_1582);
nand U1322 (N_1322,N_1172,N_1047);
nand U1323 (N_1323,N_1108,N_833);
and U1324 (N_1324,N_801,In_1813);
or U1325 (N_1325,N_1034,N_958);
and U1326 (N_1326,N_1073,In_1906);
and U1327 (N_1327,N_933,N_1098);
nand U1328 (N_1328,In_809,In_849);
nor U1329 (N_1329,N_1036,N_532);
and U1330 (N_1330,N_904,N_1080);
and U1331 (N_1331,N_1052,N_267);
nor U1332 (N_1332,N_342,N_1100);
nor U1333 (N_1333,In_495,In_1398);
or U1334 (N_1334,N_1129,N_856);
and U1335 (N_1335,N_627,In_740);
nor U1336 (N_1336,N_589,In_1418);
nor U1337 (N_1337,N_1156,In_470);
nand U1338 (N_1338,N_435,N_444);
or U1339 (N_1339,N_940,N_852);
nor U1340 (N_1340,In_44,In_106);
and U1341 (N_1341,In_194,In_781);
nand U1342 (N_1342,In_1481,N_1097);
nand U1343 (N_1343,N_1050,N_348);
and U1344 (N_1344,In_856,N_835);
nand U1345 (N_1345,N_732,In_383);
and U1346 (N_1346,N_33,N_1001);
or U1347 (N_1347,N_343,N_160);
xnor U1348 (N_1348,In_1988,N_279);
nand U1349 (N_1349,N_330,N_785);
and U1350 (N_1350,N_979,N_729);
xnor U1351 (N_1351,N_692,N_1139);
nand U1352 (N_1352,In_1788,N_1017);
nor U1353 (N_1353,N_1070,In_927);
and U1354 (N_1354,N_450,In_347);
xor U1355 (N_1355,In_1436,In_950);
nor U1356 (N_1356,N_633,In_1486);
nand U1357 (N_1357,N_868,N_502);
nand U1358 (N_1358,N_1053,N_1081);
or U1359 (N_1359,N_938,In_1268);
nor U1360 (N_1360,In_1821,In_1422);
or U1361 (N_1361,N_1162,N_1084);
nor U1362 (N_1362,In_785,N_1046);
nand U1363 (N_1363,N_265,N_934);
and U1364 (N_1364,N_900,N_1015);
or U1365 (N_1365,N_1113,N_1077);
xor U1366 (N_1366,N_851,N_102);
nor U1367 (N_1367,N_217,N_819);
nor U1368 (N_1368,N_1037,In_91);
xnor U1369 (N_1369,In_395,N_1199);
nor U1370 (N_1370,N_895,In_748);
or U1371 (N_1371,N_914,N_434);
and U1372 (N_1372,In_1191,In_1390);
xor U1373 (N_1373,N_1191,N_1067);
or U1374 (N_1374,N_1180,N_1055);
or U1375 (N_1375,In_204,N_1143);
and U1376 (N_1376,N_525,N_687);
nor U1377 (N_1377,N_1131,In_915);
nor U1378 (N_1378,N_867,In_1658);
nor U1379 (N_1379,In_1544,N_48);
xor U1380 (N_1380,In_1223,In_1193);
or U1381 (N_1381,N_830,N_263);
nor U1382 (N_1382,N_1149,N_834);
or U1383 (N_1383,In_1626,N_1144);
nor U1384 (N_1384,N_1008,N_604);
xor U1385 (N_1385,N_1030,In_1277);
and U1386 (N_1386,In_527,In_1999);
xor U1387 (N_1387,N_1060,In_1762);
xor U1388 (N_1388,In_1621,N_587);
xnor U1389 (N_1389,N_80,N_287);
or U1390 (N_1390,In_1096,In_1329);
and U1391 (N_1391,N_921,N_441);
xor U1392 (N_1392,In_1445,N_17);
and U1393 (N_1393,N_578,N_1072);
nor U1394 (N_1394,N_812,N_1126);
nand U1395 (N_1395,N_370,N_990);
xnor U1396 (N_1396,N_344,N_1135);
nand U1397 (N_1397,N_1155,In_1229);
and U1398 (N_1398,N_1059,N_912);
xor U1399 (N_1399,In_1969,In_741);
or U1400 (N_1400,N_1068,N_1268);
xnor U1401 (N_1401,N_1254,N_1203);
xnor U1402 (N_1402,N_807,N_1188);
xnor U1403 (N_1403,In_168,N_438);
and U1404 (N_1404,N_1317,N_38);
nand U1405 (N_1405,N_31,N_1300);
nor U1406 (N_1406,N_92,In_1185);
and U1407 (N_1407,N_539,N_551);
nand U1408 (N_1408,N_1044,In_1447);
nand U1409 (N_1409,N_1224,In_1733);
xor U1410 (N_1410,N_1194,N_190);
and U1411 (N_1411,In_828,N_1192);
or U1412 (N_1412,N_1337,N_407);
or U1413 (N_1413,N_261,N_1157);
xnor U1414 (N_1414,In_1183,N_1301);
nand U1415 (N_1415,N_1346,In_104);
nand U1416 (N_1416,N_1356,N_616);
and U1417 (N_1417,N_755,N_1253);
and U1418 (N_1418,N_733,N_1236);
nor U1419 (N_1419,N_602,N_1166);
nor U1420 (N_1420,N_646,N_648);
nor U1421 (N_1421,N_1058,N_1221);
and U1422 (N_1422,In_1603,N_820);
and U1423 (N_1423,N_1214,N_556);
nor U1424 (N_1424,N_1358,N_1024);
xor U1425 (N_1425,In_734,N_1133);
and U1426 (N_1426,N_1256,N_1210);
or U1427 (N_1427,N_629,N_572);
nor U1428 (N_1428,N_328,N_1136);
nand U1429 (N_1429,N_783,N_1120);
or U1430 (N_1430,N_1386,N_1264);
nand U1431 (N_1431,In_256,N_1088);
or U1432 (N_1432,N_915,N_1388);
nand U1433 (N_1433,N_356,N_1252);
nor U1434 (N_1434,N_727,N_822);
and U1435 (N_1435,N_1334,N_1344);
or U1436 (N_1436,N_848,N_1223);
or U1437 (N_1437,N_1380,N_1319);
nand U1438 (N_1438,N_766,N_1295);
xor U1439 (N_1439,N_821,In_777);
or U1440 (N_1440,N_1175,N_1019);
nor U1441 (N_1441,N_1218,N_1318);
xnor U1442 (N_1442,In_766,N_445);
xor U1443 (N_1443,N_1324,N_869);
xnor U1444 (N_1444,In_754,In_1081);
or U1445 (N_1445,N_1119,N_1370);
nand U1446 (N_1446,N_1345,N_1375);
nand U1447 (N_1447,In_1803,N_1297);
xnor U1448 (N_1448,N_1079,N_182);
xnor U1449 (N_1449,N_1357,N_757);
or U1450 (N_1450,In_485,N_1305);
xor U1451 (N_1451,N_1219,N_1082);
and U1452 (N_1452,N_657,N_671);
or U1453 (N_1453,N_1112,In_1774);
nor U1454 (N_1454,N_1381,N_1174);
and U1455 (N_1455,N_1266,N_836);
nor U1456 (N_1456,N_1298,N_976);
and U1457 (N_1457,N_605,N_1061);
nand U1458 (N_1458,N_1206,In_1523);
nand U1459 (N_1459,N_70,N_1115);
nor U1460 (N_1460,N_1078,In_617);
and U1461 (N_1461,In_343,N_784);
nand U1462 (N_1462,N_1204,N_1237);
and U1463 (N_1463,N_1327,N_588);
and U1464 (N_1464,N_1280,N_1313);
and U1465 (N_1465,N_1362,In_825);
nand U1466 (N_1466,N_1257,N_1125);
and U1467 (N_1467,N_1038,N_647);
xnor U1468 (N_1468,N_1202,N_1250);
nand U1469 (N_1469,In_478,N_112);
xor U1470 (N_1470,N_301,N_1306);
and U1471 (N_1471,N_619,N_884);
nand U1472 (N_1472,N_673,In_360);
nor U1473 (N_1473,N_889,N_479);
or U1474 (N_1474,In_1071,N_496);
nand U1475 (N_1475,N_1283,N_1121);
nand U1476 (N_1476,N_935,N_1217);
xor U1477 (N_1477,In_1173,N_271);
xnor U1478 (N_1478,N_883,N_521);
and U1479 (N_1479,N_1312,N_932);
or U1480 (N_1480,N_1014,N_1103);
and U1481 (N_1481,N_995,In_709);
xor U1482 (N_1482,N_1349,N_1012);
and U1483 (N_1483,In_1078,N_1385);
nand U1484 (N_1484,N_1310,N_12);
or U1485 (N_1485,In_166,N_320);
nor U1486 (N_1486,In_340,N_295);
nand U1487 (N_1487,N_1292,N_831);
nor U1488 (N_1488,In_680,N_1377);
xor U1489 (N_1489,N_1296,In_753);
or U1490 (N_1490,N_1261,N_690);
xnor U1491 (N_1491,In_756,In_1382);
xor U1492 (N_1492,N_1275,N_991);
nor U1493 (N_1493,N_772,In_1013);
and U1494 (N_1494,N_1109,N_1234);
nand U1495 (N_1495,N_358,N_1154);
and U1496 (N_1496,N_481,N_1057);
nor U1497 (N_1497,N_138,N_954);
nand U1498 (N_1498,N_1170,N_1063);
nand U1499 (N_1499,N_746,N_1229);
nand U1500 (N_1500,In_344,N_1321);
or U1501 (N_1501,In_1662,N_996);
or U1502 (N_1502,N_234,N_1289);
and U1503 (N_1503,N_1282,N_1201);
or U1504 (N_1504,N_1006,In_284);
nor U1505 (N_1505,N_987,In_750);
nor U1506 (N_1506,N_498,N_809);
and U1507 (N_1507,N_553,N_1369);
nand U1508 (N_1508,N_1000,In_1180);
and U1509 (N_1509,N_899,N_1397);
nand U1510 (N_1510,N_454,N_1308);
nand U1511 (N_1511,In_774,N_924);
nand U1512 (N_1512,N_181,N_944);
xnor U1513 (N_1513,N_1307,N_2);
nor U1514 (N_1514,N_726,In_903);
or U1515 (N_1515,N_730,In_890);
or U1516 (N_1516,N_1365,In_402);
and U1517 (N_1517,N_1398,N_1054);
nor U1518 (N_1518,N_413,In_457);
xnor U1519 (N_1519,N_71,N_1251);
and U1520 (N_1520,In_826,In_1853);
nor U1521 (N_1521,N_926,In_1053);
or U1522 (N_1522,N_1002,N_1071);
nand U1523 (N_1523,N_1316,N_480);
or U1524 (N_1524,N_928,In_509);
xnor U1525 (N_1525,N_1355,N_688);
xor U1526 (N_1526,N_10,In_1503);
nor U1527 (N_1527,N_1208,In_651);
or U1528 (N_1528,N_1290,N_352);
nand U1529 (N_1529,N_1062,N_366);
or U1530 (N_1530,N_319,N_1212);
nand U1531 (N_1531,N_1291,N_1273);
nor U1532 (N_1532,In_860,N_209);
xor U1533 (N_1533,N_1245,N_1372);
nand U1534 (N_1534,N_338,N_1124);
and U1535 (N_1535,N_1148,In_447);
nand U1536 (N_1536,N_1333,N_902);
xor U1537 (N_1537,N_826,N_601);
nor U1538 (N_1538,N_1272,N_357);
xnor U1539 (N_1539,N_1286,In_1991);
or U1540 (N_1540,N_399,N_1363);
or U1541 (N_1541,N_1220,N_760);
nor U1542 (N_1542,N_956,In_633);
nand U1543 (N_1543,N_769,N_691);
nor U1544 (N_1544,N_1209,N_1106);
and U1545 (N_1545,In_1700,N_1083);
and U1546 (N_1546,In_821,N_949);
nor U1547 (N_1547,N_1389,N_905);
or U1548 (N_1548,N_1347,In_1002);
and U1549 (N_1549,N_1138,In_666);
nor U1550 (N_1550,N_893,N_91);
nor U1551 (N_1551,In_1844,N_1049);
nand U1552 (N_1552,In_564,N_876);
nor U1553 (N_1553,In_1132,In_1073);
nand U1554 (N_1554,In_384,N_1197);
nor U1555 (N_1555,In_205,N_874);
nor U1556 (N_1556,N_1315,N_1281);
xor U1557 (N_1557,N_1330,N_1215);
nor U1558 (N_1558,In_1739,N_264);
or U1559 (N_1559,N_1101,N_1075);
nor U1560 (N_1560,N_1269,N_1226);
nand U1561 (N_1561,N_1332,N_1182);
xnor U1562 (N_1562,N_25,N_734);
or U1563 (N_1563,In_1315,In_1721);
or U1564 (N_1564,N_813,N_1353);
nor U1565 (N_1565,N_1093,N_1207);
and U1566 (N_1566,N_1311,In_1356);
nor U1567 (N_1567,In_968,N_1392);
and U1568 (N_1568,N_1118,N_1225);
xnor U1569 (N_1569,N_796,N_1395);
or U1570 (N_1570,N_758,In_1245);
or U1571 (N_1571,N_1134,In_1551);
xnor U1572 (N_1572,N_451,In_689);
nand U1573 (N_1573,N_1359,N_1288);
nor U1574 (N_1574,N_1354,In_1492);
xor U1575 (N_1575,In_1232,N_359);
and U1576 (N_1576,N_1248,N_1200);
xor U1577 (N_1577,N_1331,N_1339);
xnor U1578 (N_1578,N_1368,In_901);
or U1579 (N_1579,N_1325,N_1116);
or U1580 (N_1580,N_1294,N_1176);
nand U1581 (N_1581,N_1235,In_451);
nor U1582 (N_1582,In_1839,N_853);
or U1583 (N_1583,N_1045,N_307);
and U1584 (N_1584,N_850,N_1271);
and U1585 (N_1585,N_1099,N_1287);
xnor U1586 (N_1586,N_1003,N_1246);
and U1587 (N_1587,N_420,N_1378);
xor U1588 (N_1588,N_1096,N_1040);
and U1589 (N_1589,N_1393,In_1026);
xor U1590 (N_1590,In_660,N_1205);
and U1591 (N_1591,N_419,In_287);
and U1592 (N_1592,N_1092,N_1277);
and U1593 (N_1593,N_1146,N_1020);
nor U1594 (N_1594,N_1399,N_1304);
xnor U1595 (N_1595,In_1280,N_877);
nand U1596 (N_1596,N_1263,N_1394);
or U1597 (N_1597,In_1880,In_1776);
nor U1598 (N_1598,N_1384,N_1128);
and U1599 (N_1599,In_488,N_770);
nor U1600 (N_1600,N_1549,N_1249);
or U1601 (N_1601,N_1262,N_955);
xor U1602 (N_1602,In_1453,N_1242);
nor U1603 (N_1603,N_1391,N_1580);
or U1604 (N_1604,N_1402,In_1915);
xor U1605 (N_1605,N_1446,N_1342);
nor U1606 (N_1606,In_275,N_1441);
and U1607 (N_1607,N_1478,N_1450);
xnor U1608 (N_1608,N_1410,N_937);
nand U1609 (N_1609,N_1556,N_1076);
and U1610 (N_1610,N_1463,N_1567);
nor U1611 (N_1611,N_1547,N_1559);
or U1612 (N_1612,N_1476,N_1581);
or U1613 (N_1613,In_1878,In_1578);
or U1614 (N_1614,N_1526,In_702);
nor U1615 (N_1615,In_648,In_1605);
or U1616 (N_1616,N_1494,N_1534);
xnor U1617 (N_1617,N_439,N_1198);
xor U1618 (N_1618,N_1484,N_1533);
and U1619 (N_1619,N_1340,N_1195);
or U1620 (N_1620,N_1258,N_1461);
and U1621 (N_1621,N_1470,N_1265);
nor U1622 (N_1622,N_1416,N_1299);
and U1623 (N_1623,N_1360,N_1383);
nor U1624 (N_1624,N_1531,N_1507);
nor U1625 (N_1625,N_1558,N_1537);
nand U1626 (N_1626,In_1686,N_1569);
and U1627 (N_1627,N_1594,N_1405);
nor U1628 (N_1628,N_620,N_1477);
nor U1629 (N_1629,N_1560,In_827);
nor U1630 (N_1630,N_166,N_1588);
or U1631 (N_1631,N_570,N_1302);
nand U1632 (N_1632,N_711,N_1599);
and U1633 (N_1633,N_1485,N_827);
xnor U1634 (N_1634,N_1432,N_862);
or U1635 (N_1635,N_1467,N_1512);
xor U1636 (N_1636,N_1434,N_1335);
and U1637 (N_1637,N_744,N_1453);
or U1638 (N_1638,N_1230,In_1359);
or U1639 (N_1639,N_1173,N_1511);
xnor U1640 (N_1640,N_1452,N_878);
and U1641 (N_1641,N_1482,N_652);
nor U1642 (N_1642,N_557,N_1211);
or U1643 (N_1643,N_1472,N_1105);
nand U1644 (N_1644,N_1576,N_68);
xnor U1645 (N_1645,N_1241,In_1591);
nor U1646 (N_1646,N_1473,N_707);
nand U1647 (N_1647,N_1171,N_1525);
nand U1648 (N_1648,N_1048,N_811);
nand U1649 (N_1649,N_106,N_1425);
and U1650 (N_1650,N_1095,N_1573);
xnor U1651 (N_1651,N_1498,N_1343);
xnor U1652 (N_1652,N_1532,N_145);
or U1653 (N_1653,N_1309,N_492);
xnor U1654 (N_1654,N_837,N_1419);
nor U1655 (N_1655,N_763,N_1326);
nor U1656 (N_1656,N_1323,In_1278);
or U1657 (N_1657,N_1091,N_1587);
xor U1658 (N_1658,N_1506,N_1431);
nor U1659 (N_1659,N_1127,N_1457);
and U1660 (N_1660,N_1238,N_1426);
xor U1661 (N_1661,N_1553,N_1490);
or U1662 (N_1662,N_1403,N_1445);
xnor U1663 (N_1663,N_1400,N_1279);
nand U1664 (N_1664,N_1247,N_1285);
or U1665 (N_1665,N_1367,In_1199);
xnor U1666 (N_1666,N_1348,In_138);
or U1667 (N_1667,N_1462,N_1510);
nor U1668 (N_1668,N_975,N_1469);
nand U1669 (N_1669,In_920,N_943);
or U1670 (N_1670,N_1488,N_1437);
or U1671 (N_1671,N_981,N_1487);
nand U1672 (N_1672,N_1418,N_1352);
nand U1673 (N_1673,N_253,N_1379);
nand U1674 (N_1674,N_1538,N_1429);
nand U1675 (N_1675,N_1341,N_986);
or U1676 (N_1676,N_1486,N_1447);
nor U1677 (N_1677,N_1259,N_1565);
or U1678 (N_1678,In_419,N_1545);
xnor U1679 (N_1679,N_1535,N_1539);
and U1680 (N_1680,N_1278,N_1592);
nand U1681 (N_1681,N_1550,N_854);
nand U1682 (N_1682,N_1501,N_62);
nand U1683 (N_1683,In_41,N_828);
xor U1684 (N_1684,N_1564,N_1240);
nand U1685 (N_1685,N_1184,N_908);
xnor U1686 (N_1686,N_1584,N_1085);
or U1687 (N_1687,N_1213,N_575);
nor U1688 (N_1688,N_1427,N_1577);
or U1689 (N_1689,N_1540,N_1293);
nand U1690 (N_1690,N_1303,N_1586);
or U1691 (N_1691,N_1031,N_524);
and U1692 (N_1692,N_1433,N_1390);
nor U1693 (N_1693,N_1366,N_1422);
nand U1694 (N_1694,N_1481,N_1459);
xnor U1695 (N_1695,N_1582,N_1376);
xor U1696 (N_1696,N_1442,N_1598);
nor U1697 (N_1697,In_1316,N_1555);
nand U1698 (N_1698,N_1523,N_1471);
nand U1699 (N_1699,N_1243,N_1516);
nor U1700 (N_1700,N_1228,N_1500);
xor U1701 (N_1701,N_1066,N_1464);
xor U1702 (N_1702,N_1160,N_1585);
xor U1703 (N_1703,N_1458,N_1492);
nor U1704 (N_1704,In_587,N_1449);
xnor U1705 (N_1705,N_1042,N_1570);
nand U1706 (N_1706,N_1527,N_1274);
xnor U1707 (N_1707,N_1373,N_1420);
xor U1708 (N_1708,N_1364,N_695);
nor U1709 (N_1709,N_1536,N_1480);
nor U1710 (N_1710,N_1489,N_1502);
nand U1711 (N_1711,N_1021,N_1524);
nor U1712 (N_1712,N_1374,N_1597);
and U1713 (N_1713,In_1119,N_1528);
or U1714 (N_1714,N_1232,In_889);
nor U1715 (N_1715,N_1231,N_1589);
nand U1716 (N_1716,N_988,N_1408);
and U1717 (N_1717,N_1406,N_1460);
xor U1718 (N_1718,N_1412,N_1415);
or U1719 (N_1719,N_1276,N_1505);
nor U1720 (N_1720,N_901,N_1474);
or U1721 (N_1721,In_521,N_1496);
xor U1722 (N_1722,N_1270,N_1595);
xor U1723 (N_1723,N_1351,N_1513);
nand U1724 (N_1724,N_1515,N_1411);
nand U1725 (N_1725,N_1561,N_1583);
nor U1726 (N_1726,N_1421,N_1010);
nor U1727 (N_1727,N_1591,N_1596);
and U1728 (N_1728,N_1451,N_1244);
nor U1729 (N_1729,N_1552,N_1409);
or U1730 (N_1730,N_1314,In_160);
nand U1731 (N_1731,N_1440,N_756);
nand U1732 (N_1732,N_1239,N_1465);
nor U1733 (N_1733,N_1284,N_1338);
nor U1734 (N_1734,N_1361,N_1435);
xnor U1735 (N_1735,In_130,N_1022);
nor U1736 (N_1736,N_1443,In_1462);
nor U1737 (N_1737,N_1227,N_1590);
xor U1738 (N_1738,N_1439,N_864);
xnor U1739 (N_1739,N_1216,N_1428);
xnor U1740 (N_1740,N_1520,N_1521);
nand U1741 (N_1741,N_1468,N_1530);
or U1742 (N_1742,N_1566,N_1544);
nand U1743 (N_1743,N_1497,N_387);
and U1744 (N_1744,N_882,N_1543);
xor U1745 (N_1745,N_1563,In_1038);
xor U1746 (N_1746,N_1479,N_1514);
and U1747 (N_1747,N_1183,In_1473);
or U1748 (N_1748,N_1499,N_1233);
nand U1749 (N_1749,N_1571,N_1424);
and U1750 (N_1750,N_1519,N_1541);
nand U1751 (N_1751,In_1866,N_1187);
and U1752 (N_1752,N_1222,N_929);
nor U1753 (N_1753,N_1051,N_1493);
xnor U1754 (N_1754,N_1087,N_1557);
xnor U1755 (N_1755,N_1396,N_1153);
xor U1756 (N_1756,N_1456,N_404);
and U1757 (N_1757,N_1371,In_1353);
or U1758 (N_1758,N_1504,N_1255);
nand U1759 (N_1759,N_1551,N_967);
xor U1760 (N_1760,N_1423,In_939);
nor U1761 (N_1761,N_1417,N_1267);
or U1762 (N_1762,N_1448,N_1562);
or U1763 (N_1763,N_13,N_1554);
nand U1764 (N_1764,N_1579,In_1585);
xnor U1765 (N_1765,N_1466,N_919);
xnor U1766 (N_1766,N_1483,N_1491);
and U1767 (N_1767,N_1438,N_1322);
or U1768 (N_1768,N_1548,N_1436);
or U1769 (N_1769,N_1147,N_1455);
nand U1770 (N_1770,N_1328,N_1413);
xnor U1771 (N_1771,N_1509,N_1546);
and U1772 (N_1772,N_537,In_852);
and U1773 (N_1773,N_1064,N_1568);
nor U1774 (N_1774,N_150,In_563);
and U1775 (N_1775,In_1040,N_1165);
nand U1776 (N_1776,In_1518,N_1495);
nand U1777 (N_1777,N_1111,N_1542);
nor U1778 (N_1778,In_129,In_1996);
nand U1779 (N_1779,N_1518,N_1336);
xor U1780 (N_1780,N_1517,N_984);
nand U1781 (N_1781,N_1572,N_635);
and U1782 (N_1782,N_1329,N_1350);
nor U1783 (N_1783,N_1575,N_1414);
nand U1784 (N_1784,N_978,N_1102);
xor U1785 (N_1785,N_1404,N_725);
xor U1786 (N_1786,N_686,N_1475);
nand U1787 (N_1787,N_1150,N_748);
nor U1788 (N_1788,In_891,N_1387);
nand U1789 (N_1789,N_1011,In_788);
and U1790 (N_1790,N_993,N_186);
nor U1791 (N_1791,N_1578,N_1407);
nand U1792 (N_1792,N_1593,N_1508);
or U1793 (N_1793,N_1444,N_1401);
nand U1794 (N_1794,N_1522,N_1382);
xor U1795 (N_1795,N_1529,N_1320);
and U1796 (N_1796,N_1430,In_1857);
xnor U1797 (N_1797,N_1503,N_1260);
nand U1798 (N_1798,N_918,N_1574);
nor U1799 (N_1799,In_1892,N_1454);
nor U1800 (N_1800,N_1706,N_1691);
xnor U1801 (N_1801,N_1759,N_1737);
xnor U1802 (N_1802,N_1628,N_1669);
and U1803 (N_1803,N_1623,N_1696);
xnor U1804 (N_1804,N_1752,N_1638);
and U1805 (N_1805,N_1749,N_1796);
nand U1806 (N_1806,N_1660,N_1797);
xor U1807 (N_1807,N_1659,N_1719);
nor U1808 (N_1808,N_1729,N_1777);
nor U1809 (N_1809,N_1773,N_1699);
and U1810 (N_1810,N_1634,N_1666);
or U1811 (N_1811,N_1661,N_1671);
and U1812 (N_1812,N_1781,N_1686);
nor U1813 (N_1813,N_1609,N_1718);
or U1814 (N_1814,N_1757,N_1748);
nor U1815 (N_1815,N_1791,N_1769);
or U1816 (N_1816,N_1619,N_1701);
and U1817 (N_1817,N_1716,N_1709);
nand U1818 (N_1818,N_1707,N_1667);
or U1819 (N_1819,N_1606,N_1690);
and U1820 (N_1820,N_1687,N_1766);
nor U1821 (N_1821,N_1656,N_1767);
nand U1822 (N_1822,N_1613,N_1778);
and U1823 (N_1823,N_1650,N_1625);
nor U1824 (N_1824,N_1604,N_1772);
nand U1825 (N_1825,N_1714,N_1768);
xor U1826 (N_1826,N_1751,N_1636);
nor U1827 (N_1827,N_1668,N_1639);
or U1828 (N_1828,N_1703,N_1723);
or U1829 (N_1829,N_1754,N_1645);
nor U1830 (N_1830,N_1787,N_1774);
nand U1831 (N_1831,N_1731,N_1655);
nand U1832 (N_1832,N_1607,N_1775);
nand U1833 (N_1833,N_1713,N_1700);
nand U1834 (N_1834,N_1711,N_1653);
or U1835 (N_1835,N_1732,N_1637);
nand U1836 (N_1836,N_1758,N_1761);
nor U1837 (N_1837,N_1600,N_1727);
or U1838 (N_1838,N_1735,N_1741);
and U1839 (N_1839,N_1684,N_1601);
xor U1840 (N_1840,N_1692,N_1631);
nor U1841 (N_1841,N_1683,N_1730);
or U1842 (N_1842,N_1780,N_1770);
and U1843 (N_1843,N_1657,N_1618);
nand U1844 (N_1844,N_1695,N_1624);
nor U1845 (N_1845,N_1743,N_1633);
xor U1846 (N_1846,N_1764,N_1611);
and U1847 (N_1847,N_1726,N_1708);
and U1848 (N_1848,N_1664,N_1682);
or U1849 (N_1849,N_1693,N_1629);
xnor U1850 (N_1850,N_1675,N_1779);
or U1851 (N_1851,N_1649,N_1680);
or U1852 (N_1852,N_1760,N_1673);
nor U1853 (N_1853,N_1755,N_1753);
nor U1854 (N_1854,N_1670,N_1790);
nand U1855 (N_1855,N_1728,N_1792);
nor U1856 (N_1856,N_1662,N_1722);
and U1857 (N_1857,N_1632,N_1725);
and U1858 (N_1858,N_1622,N_1799);
and U1859 (N_1859,N_1626,N_1798);
xnor U1860 (N_1860,N_1608,N_1785);
nor U1861 (N_1861,N_1776,N_1724);
nand U1862 (N_1862,N_1747,N_1617);
nor U1863 (N_1863,N_1615,N_1702);
nor U1864 (N_1864,N_1652,N_1642);
xor U1865 (N_1865,N_1614,N_1721);
and U1866 (N_1866,N_1665,N_1771);
and U1867 (N_1867,N_1676,N_1745);
nor U1868 (N_1868,N_1750,N_1782);
xor U1869 (N_1869,N_1789,N_1697);
and U1870 (N_1870,N_1762,N_1744);
or U1871 (N_1871,N_1715,N_1679);
xor U1872 (N_1872,N_1663,N_1612);
nor U1873 (N_1873,N_1694,N_1742);
or U1874 (N_1874,N_1620,N_1704);
xnor U1875 (N_1875,N_1641,N_1765);
xnor U1876 (N_1876,N_1736,N_1644);
nand U1877 (N_1877,N_1678,N_1672);
xnor U1878 (N_1878,N_1734,N_1677);
and U1879 (N_1879,N_1648,N_1688);
nor U1880 (N_1880,N_1783,N_1739);
nand U1881 (N_1881,N_1793,N_1784);
nor U1882 (N_1882,N_1740,N_1786);
or U1883 (N_1883,N_1605,N_1705);
or U1884 (N_1884,N_1643,N_1746);
nand U1885 (N_1885,N_1685,N_1640);
and U1886 (N_1886,N_1674,N_1698);
nor U1887 (N_1887,N_1651,N_1720);
and U1888 (N_1888,N_1630,N_1658);
or U1889 (N_1889,N_1627,N_1689);
nor U1890 (N_1890,N_1712,N_1654);
xnor U1891 (N_1891,N_1621,N_1616);
or U1892 (N_1892,N_1602,N_1646);
and U1893 (N_1893,N_1763,N_1756);
nand U1894 (N_1894,N_1794,N_1603);
or U1895 (N_1895,N_1733,N_1647);
or U1896 (N_1896,N_1681,N_1710);
nor U1897 (N_1897,N_1788,N_1635);
xnor U1898 (N_1898,N_1795,N_1717);
and U1899 (N_1899,N_1738,N_1610);
nor U1900 (N_1900,N_1705,N_1619);
nand U1901 (N_1901,N_1626,N_1629);
nor U1902 (N_1902,N_1625,N_1722);
nor U1903 (N_1903,N_1632,N_1688);
nor U1904 (N_1904,N_1691,N_1793);
nor U1905 (N_1905,N_1768,N_1791);
or U1906 (N_1906,N_1758,N_1696);
nand U1907 (N_1907,N_1730,N_1704);
or U1908 (N_1908,N_1689,N_1680);
and U1909 (N_1909,N_1705,N_1779);
and U1910 (N_1910,N_1687,N_1636);
nor U1911 (N_1911,N_1619,N_1790);
and U1912 (N_1912,N_1712,N_1791);
and U1913 (N_1913,N_1629,N_1716);
nor U1914 (N_1914,N_1697,N_1632);
and U1915 (N_1915,N_1775,N_1683);
nor U1916 (N_1916,N_1799,N_1659);
or U1917 (N_1917,N_1786,N_1711);
nor U1918 (N_1918,N_1746,N_1673);
nor U1919 (N_1919,N_1719,N_1721);
nand U1920 (N_1920,N_1778,N_1648);
nor U1921 (N_1921,N_1660,N_1769);
or U1922 (N_1922,N_1768,N_1716);
nand U1923 (N_1923,N_1737,N_1787);
xnor U1924 (N_1924,N_1697,N_1680);
xnor U1925 (N_1925,N_1688,N_1708);
and U1926 (N_1926,N_1648,N_1628);
nor U1927 (N_1927,N_1645,N_1664);
nor U1928 (N_1928,N_1619,N_1797);
nand U1929 (N_1929,N_1704,N_1733);
nand U1930 (N_1930,N_1667,N_1757);
and U1931 (N_1931,N_1792,N_1697);
or U1932 (N_1932,N_1775,N_1701);
and U1933 (N_1933,N_1682,N_1708);
nand U1934 (N_1934,N_1763,N_1603);
or U1935 (N_1935,N_1678,N_1628);
nand U1936 (N_1936,N_1722,N_1795);
xnor U1937 (N_1937,N_1761,N_1688);
or U1938 (N_1938,N_1619,N_1788);
nand U1939 (N_1939,N_1731,N_1747);
and U1940 (N_1940,N_1614,N_1628);
nand U1941 (N_1941,N_1612,N_1745);
or U1942 (N_1942,N_1614,N_1712);
nand U1943 (N_1943,N_1632,N_1638);
and U1944 (N_1944,N_1602,N_1736);
and U1945 (N_1945,N_1626,N_1733);
or U1946 (N_1946,N_1611,N_1655);
xor U1947 (N_1947,N_1772,N_1706);
nor U1948 (N_1948,N_1676,N_1740);
or U1949 (N_1949,N_1789,N_1751);
and U1950 (N_1950,N_1771,N_1634);
nor U1951 (N_1951,N_1740,N_1623);
xor U1952 (N_1952,N_1700,N_1618);
xnor U1953 (N_1953,N_1660,N_1696);
and U1954 (N_1954,N_1757,N_1730);
nor U1955 (N_1955,N_1720,N_1739);
nand U1956 (N_1956,N_1687,N_1612);
or U1957 (N_1957,N_1748,N_1714);
xor U1958 (N_1958,N_1670,N_1717);
and U1959 (N_1959,N_1621,N_1781);
nand U1960 (N_1960,N_1768,N_1655);
and U1961 (N_1961,N_1705,N_1744);
nor U1962 (N_1962,N_1757,N_1648);
nor U1963 (N_1963,N_1741,N_1663);
or U1964 (N_1964,N_1639,N_1709);
nor U1965 (N_1965,N_1690,N_1623);
nand U1966 (N_1966,N_1718,N_1686);
xor U1967 (N_1967,N_1784,N_1623);
nor U1968 (N_1968,N_1641,N_1603);
nand U1969 (N_1969,N_1732,N_1654);
and U1970 (N_1970,N_1628,N_1616);
nor U1971 (N_1971,N_1730,N_1707);
xor U1972 (N_1972,N_1621,N_1653);
and U1973 (N_1973,N_1620,N_1671);
xnor U1974 (N_1974,N_1649,N_1625);
and U1975 (N_1975,N_1654,N_1697);
nand U1976 (N_1976,N_1768,N_1636);
nor U1977 (N_1977,N_1642,N_1686);
or U1978 (N_1978,N_1782,N_1762);
nor U1979 (N_1979,N_1623,N_1622);
nand U1980 (N_1980,N_1610,N_1780);
and U1981 (N_1981,N_1752,N_1602);
or U1982 (N_1982,N_1780,N_1686);
or U1983 (N_1983,N_1703,N_1686);
nand U1984 (N_1984,N_1686,N_1648);
nor U1985 (N_1985,N_1730,N_1766);
and U1986 (N_1986,N_1647,N_1655);
and U1987 (N_1987,N_1708,N_1747);
nor U1988 (N_1988,N_1640,N_1769);
or U1989 (N_1989,N_1762,N_1775);
or U1990 (N_1990,N_1697,N_1696);
or U1991 (N_1991,N_1602,N_1741);
nor U1992 (N_1992,N_1702,N_1664);
and U1993 (N_1993,N_1683,N_1644);
xor U1994 (N_1994,N_1616,N_1636);
and U1995 (N_1995,N_1790,N_1754);
xnor U1996 (N_1996,N_1631,N_1707);
and U1997 (N_1997,N_1603,N_1608);
or U1998 (N_1998,N_1766,N_1715);
nand U1999 (N_1999,N_1784,N_1684);
xnor U2000 (N_2000,N_1838,N_1856);
nand U2001 (N_2001,N_1835,N_1870);
nand U2002 (N_2002,N_1941,N_1923);
or U2003 (N_2003,N_1948,N_1827);
and U2004 (N_2004,N_1860,N_1983);
and U2005 (N_2005,N_1879,N_1848);
nor U2006 (N_2006,N_1821,N_1896);
nor U2007 (N_2007,N_1818,N_1992);
and U2008 (N_2008,N_1850,N_1857);
xor U2009 (N_2009,N_1822,N_1898);
xnor U2010 (N_2010,N_1981,N_1846);
and U2011 (N_2011,N_1905,N_1951);
and U2012 (N_2012,N_1874,N_1834);
xnor U2013 (N_2013,N_1969,N_1816);
or U2014 (N_2014,N_1864,N_1970);
or U2015 (N_2015,N_1807,N_1967);
or U2016 (N_2016,N_1899,N_1868);
nor U2017 (N_2017,N_1962,N_1993);
nand U2018 (N_2018,N_1825,N_1830);
and U2019 (N_2019,N_1893,N_1833);
nand U2020 (N_2020,N_1926,N_1862);
nand U2021 (N_2021,N_1980,N_1932);
and U2022 (N_2022,N_1804,N_1984);
and U2023 (N_2023,N_1933,N_1851);
nand U2024 (N_2024,N_1875,N_1885);
and U2025 (N_2025,N_1972,N_1853);
xor U2026 (N_2026,N_1936,N_1910);
xor U2027 (N_2027,N_1802,N_1881);
nand U2028 (N_2028,N_1858,N_1909);
nor U2029 (N_2029,N_1842,N_1968);
xor U2030 (N_2030,N_1872,N_1889);
xor U2031 (N_2031,N_1883,N_1894);
and U2032 (N_2032,N_1918,N_1954);
xor U2033 (N_2033,N_1852,N_1952);
or U2034 (N_2034,N_1963,N_1955);
nand U2035 (N_2035,N_1934,N_1888);
nand U2036 (N_2036,N_1903,N_1908);
nand U2037 (N_2037,N_1829,N_1998);
nand U2038 (N_2038,N_1817,N_1878);
nor U2039 (N_2039,N_1849,N_1895);
and U2040 (N_2040,N_1940,N_1997);
xor U2041 (N_2041,N_1866,N_1994);
nor U2042 (N_2042,N_1841,N_1813);
or U2043 (N_2043,N_1925,N_1924);
or U2044 (N_2044,N_1826,N_1901);
or U2045 (N_2045,N_1815,N_1904);
nand U2046 (N_2046,N_1880,N_1950);
xnor U2047 (N_2047,N_1946,N_1978);
and U2048 (N_2048,N_1808,N_1854);
or U2049 (N_2049,N_1986,N_1844);
nor U2050 (N_2050,N_1930,N_1911);
nor U2051 (N_2051,N_1996,N_1811);
nand U2052 (N_2052,N_1990,N_1902);
xnor U2053 (N_2053,N_1974,N_1945);
nor U2054 (N_2054,N_1979,N_1964);
nand U2055 (N_2055,N_1912,N_1931);
xnor U2056 (N_2056,N_1832,N_1922);
xor U2057 (N_2057,N_1855,N_1873);
and U2058 (N_2058,N_1919,N_1914);
nor U2059 (N_2059,N_1845,N_1812);
xor U2060 (N_2060,N_1892,N_1973);
and U2061 (N_2061,N_1991,N_1938);
or U2062 (N_2062,N_1928,N_1805);
nand U2063 (N_2063,N_1831,N_1820);
xnor U2064 (N_2064,N_1915,N_1837);
xnor U2065 (N_2065,N_1819,N_1877);
nor U2066 (N_2066,N_1966,N_1863);
xnor U2067 (N_2067,N_1987,N_1803);
nor U2068 (N_2068,N_1800,N_1989);
nor U2069 (N_2069,N_1927,N_1935);
and U2070 (N_2070,N_1810,N_1859);
xnor U2071 (N_2071,N_1887,N_1999);
and U2072 (N_2072,N_1801,N_1839);
or U2073 (N_2073,N_1977,N_1884);
and U2074 (N_2074,N_1906,N_1995);
and U2075 (N_2075,N_1942,N_1917);
nand U2076 (N_2076,N_1886,N_1869);
and U2077 (N_2077,N_1882,N_1985);
or U2078 (N_2078,N_1823,N_1947);
nor U2079 (N_2079,N_1976,N_1913);
xor U2080 (N_2080,N_1982,N_1867);
xnor U2081 (N_2081,N_1971,N_1959);
and U2082 (N_2082,N_1956,N_1916);
nand U2083 (N_2083,N_1824,N_1891);
xor U2084 (N_2084,N_1900,N_1949);
nor U2085 (N_2085,N_1809,N_1876);
nor U2086 (N_2086,N_1897,N_1961);
xnor U2087 (N_2087,N_1943,N_1944);
nor U2088 (N_2088,N_1960,N_1957);
or U2089 (N_2089,N_1937,N_1965);
xor U2090 (N_2090,N_1890,N_1988);
nand U2091 (N_2091,N_1920,N_1828);
or U2092 (N_2092,N_1953,N_1865);
nand U2093 (N_2093,N_1847,N_1843);
nand U2094 (N_2094,N_1907,N_1836);
nand U2095 (N_2095,N_1861,N_1806);
xor U2096 (N_2096,N_1921,N_1840);
nand U2097 (N_2097,N_1939,N_1814);
and U2098 (N_2098,N_1871,N_1929);
nand U2099 (N_2099,N_1975,N_1958);
nor U2100 (N_2100,N_1958,N_1897);
and U2101 (N_2101,N_1803,N_1865);
nand U2102 (N_2102,N_1990,N_1983);
and U2103 (N_2103,N_1912,N_1836);
or U2104 (N_2104,N_1831,N_1862);
and U2105 (N_2105,N_1915,N_1923);
nand U2106 (N_2106,N_1831,N_1982);
xnor U2107 (N_2107,N_1976,N_1806);
and U2108 (N_2108,N_1856,N_1948);
nor U2109 (N_2109,N_1986,N_1801);
nand U2110 (N_2110,N_1975,N_1913);
nand U2111 (N_2111,N_1913,N_1916);
or U2112 (N_2112,N_1819,N_1808);
nor U2113 (N_2113,N_1898,N_1978);
nor U2114 (N_2114,N_1873,N_1823);
nand U2115 (N_2115,N_1932,N_1825);
nor U2116 (N_2116,N_1921,N_1980);
nand U2117 (N_2117,N_1994,N_1988);
nor U2118 (N_2118,N_1823,N_1818);
nor U2119 (N_2119,N_1969,N_1995);
nor U2120 (N_2120,N_1825,N_1913);
nand U2121 (N_2121,N_1859,N_1967);
or U2122 (N_2122,N_1920,N_1858);
nand U2123 (N_2123,N_1907,N_1810);
and U2124 (N_2124,N_1870,N_1874);
and U2125 (N_2125,N_1886,N_1815);
nand U2126 (N_2126,N_1902,N_1869);
nand U2127 (N_2127,N_1801,N_1874);
xnor U2128 (N_2128,N_1800,N_1976);
and U2129 (N_2129,N_1868,N_1911);
nor U2130 (N_2130,N_1960,N_1873);
xor U2131 (N_2131,N_1925,N_1949);
nand U2132 (N_2132,N_1931,N_1939);
nand U2133 (N_2133,N_1982,N_1920);
nor U2134 (N_2134,N_1805,N_1848);
or U2135 (N_2135,N_1993,N_1887);
nor U2136 (N_2136,N_1881,N_1904);
nor U2137 (N_2137,N_1925,N_1997);
nor U2138 (N_2138,N_1888,N_1895);
or U2139 (N_2139,N_1975,N_1812);
and U2140 (N_2140,N_1918,N_1876);
and U2141 (N_2141,N_1854,N_1981);
xor U2142 (N_2142,N_1806,N_1915);
nor U2143 (N_2143,N_1884,N_1968);
and U2144 (N_2144,N_1870,N_1979);
nand U2145 (N_2145,N_1880,N_1808);
nor U2146 (N_2146,N_1831,N_1834);
and U2147 (N_2147,N_1830,N_1882);
xor U2148 (N_2148,N_1976,N_1993);
or U2149 (N_2149,N_1859,N_1864);
nand U2150 (N_2150,N_1933,N_1956);
nor U2151 (N_2151,N_1995,N_1813);
nand U2152 (N_2152,N_1948,N_1873);
or U2153 (N_2153,N_1969,N_1991);
or U2154 (N_2154,N_1845,N_1851);
nor U2155 (N_2155,N_1836,N_1966);
nor U2156 (N_2156,N_1982,N_1905);
xnor U2157 (N_2157,N_1914,N_1868);
and U2158 (N_2158,N_1892,N_1961);
or U2159 (N_2159,N_1958,N_1947);
xnor U2160 (N_2160,N_1837,N_1933);
xnor U2161 (N_2161,N_1941,N_1964);
nor U2162 (N_2162,N_1927,N_1899);
and U2163 (N_2163,N_1934,N_1979);
nor U2164 (N_2164,N_1936,N_1921);
nand U2165 (N_2165,N_1924,N_1897);
and U2166 (N_2166,N_1976,N_1801);
nand U2167 (N_2167,N_1876,N_1937);
nand U2168 (N_2168,N_1815,N_1923);
or U2169 (N_2169,N_1846,N_1805);
nor U2170 (N_2170,N_1852,N_1945);
nor U2171 (N_2171,N_1980,N_1801);
nand U2172 (N_2172,N_1843,N_1844);
and U2173 (N_2173,N_1888,N_1955);
nor U2174 (N_2174,N_1872,N_1917);
or U2175 (N_2175,N_1851,N_1929);
nor U2176 (N_2176,N_1972,N_1844);
xnor U2177 (N_2177,N_1921,N_1955);
or U2178 (N_2178,N_1834,N_1813);
xnor U2179 (N_2179,N_1846,N_1898);
nor U2180 (N_2180,N_1913,N_1971);
and U2181 (N_2181,N_1918,N_1937);
nor U2182 (N_2182,N_1960,N_1916);
nor U2183 (N_2183,N_1929,N_1905);
nor U2184 (N_2184,N_1835,N_1926);
xnor U2185 (N_2185,N_1968,N_1887);
xor U2186 (N_2186,N_1928,N_1931);
nor U2187 (N_2187,N_1921,N_1807);
nor U2188 (N_2188,N_1839,N_1946);
xnor U2189 (N_2189,N_1817,N_1844);
and U2190 (N_2190,N_1887,N_1981);
and U2191 (N_2191,N_1882,N_1874);
nor U2192 (N_2192,N_1947,N_1991);
nor U2193 (N_2193,N_1886,N_1981);
or U2194 (N_2194,N_1940,N_1924);
nand U2195 (N_2195,N_1895,N_1970);
nor U2196 (N_2196,N_1963,N_1867);
nor U2197 (N_2197,N_1923,N_1940);
xor U2198 (N_2198,N_1936,N_1937);
nor U2199 (N_2199,N_1948,N_1876);
nand U2200 (N_2200,N_2168,N_2158);
nor U2201 (N_2201,N_2193,N_2174);
or U2202 (N_2202,N_2150,N_2058);
and U2203 (N_2203,N_2087,N_2126);
xor U2204 (N_2204,N_2063,N_2179);
xor U2205 (N_2205,N_2022,N_2133);
nand U2206 (N_2206,N_2131,N_2147);
or U2207 (N_2207,N_2161,N_2002);
nand U2208 (N_2208,N_2138,N_2082);
xnor U2209 (N_2209,N_2127,N_2144);
and U2210 (N_2210,N_2057,N_2109);
and U2211 (N_2211,N_2044,N_2180);
xor U2212 (N_2212,N_2125,N_2021);
nand U2213 (N_2213,N_2198,N_2190);
or U2214 (N_2214,N_2078,N_2005);
nand U2215 (N_2215,N_2196,N_2037);
xor U2216 (N_2216,N_2080,N_2006);
nor U2217 (N_2217,N_2017,N_2154);
xor U2218 (N_2218,N_2072,N_2136);
xnor U2219 (N_2219,N_2088,N_2012);
or U2220 (N_2220,N_2159,N_2110);
and U2221 (N_2221,N_2007,N_2011);
xnor U2222 (N_2222,N_2020,N_2143);
or U2223 (N_2223,N_2079,N_2041);
nor U2224 (N_2224,N_2075,N_2128);
xor U2225 (N_2225,N_2048,N_2083);
and U2226 (N_2226,N_2081,N_2001);
xnor U2227 (N_2227,N_2070,N_2184);
nand U2228 (N_2228,N_2106,N_2027);
and U2229 (N_2229,N_2163,N_2175);
nand U2230 (N_2230,N_2003,N_2123);
nand U2231 (N_2231,N_2124,N_2118);
xor U2232 (N_2232,N_2113,N_2121);
nor U2233 (N_2233,N_2065,N_2149);
and U2234 (N_2234,N_2129,N_2046);
nand U2235 (N_2235,N_2115,N_2039);
nand U2236 (N_2236,N_2191,N_2137);
xor U2237 (N_2237,N_2117,N_2162);
and U2238 (N_2238,N_2086,N_2074);
nand U2239 (N_2239,N_2160,N_2103);
and U2240 (N_2240,N_2004,N_2024);
nor U2241 (N_2241,N_2192,N_2178);
nor U2242 (N_2242,N_2114,N_2064);
nand U2243 (N_2243,N_2187,N_2102);
and U2244 (N_2244,N_2016,N_2139);
xor U2245 (N_2245,N_2153,N_2120);
nor U2246 (N_2246,N_2052,N_2067);
nor U2247 (N_2247,N_2093,N_2073);
or U2248 (N_2248,N_2076,N_2181);
or U2249 (N_2249,N_2098,N_2099);
nor U2250 (N_2250,N_2151,N_2104);
nand U2251 (N_2251,N_2023,N_2148);
or U2252 (N_2252,N_2028,N_2172);
and U2253 (N_2253,N_2042,N_2056);
and U2254 (N_2254,N_2013,N_2155);
and U2255 (N_2255,N_2059,N_2108);
xnor U2256 (N_2256,N_2036,N_2055);
nor U2257 (N_2257,N_2197,N_2182);
and U2258 (N_2258,N_2119,N_2188);
nor U2259 (N_2259,N_2101,N_2040);
nand U2260 (N_2260,N_2060,N_2043);
and U2261 (N_2261,N_2066,N_2009);
and U2262 (N_2262,N_2164,N_2169);
nor U2263 (N_2263,N_2031,N_2030);
or U2264 (N_2264,N_2025,N_2096);
nand U2265 (N_2265,N_2105,N_2142);
or U2266 (N_2266,N_2047,N_2152);
or U2267 (N_2267,N_2156,N_2195);
or U2268 (N_2268,N_2092,N_2018);
and U2269 (N_2269,N_2089,N_2185);
and U2270 (N_2270,N_2167,N_2032);
nor U2271 (N_2271,N_2170,N_2186);
nor U2272 (N_2272,N_2122,N_2029);
xnor U2273 (N_2273,N_2014,N_2100);
and U2274 (N_2274,N_2084,N_2183);
or U2275 (N_2275,N_2095,N_2008);
and U2276 (N_2276,N_2068,N_2157);
or U2277 (N_2277,N_2034,N_2061);
xnor U2278 (N_2278,N_2140,N_2111);
nor U2279 (N_2279,N_2146,N_2090);
or U2280 (N_2280,N_2165,N_2141);
and U2281 (N_2281,N_2000,N_2097);
or U2282 (N_2282,N_2177,N_2053);
nor U2283 (N_2283,N_2019,N_2134);
or U2284 (N_2284,N_2077,N_2026);
nand U2285 (N_2285,N_2069,N_2199);
nand U2286 (N_2286,N_2116,N_2107);
nand U2287 (N_2287,N_2189,N_2194);
nand U2288 (N_2288,N_2051,N_2176);
and U2289 (N_2289,N_2045,N_2071);
or U2290 (N_2290,N_2112,N_2038);
nand U2291 (N_2291,N_2171,N_2054);
xor U2292 (N_2292,N_2132,N_2135);
nand U2293 (N_2293,N_2049,N_2145);
xnor U2294 (N_2294,N_2050,N_2091);
and U2295 (N_2295,N_2010,N_2130);
nand U2296 (N_2296,N_2015,N_2035);
nand U2297 (N_2297,N_2166,N_2085);
or U2298 (N_2298,N_2094,N_2173);
or U2299 (N_2299,N_2062,N_2033);
nor U2300 (N_2300,N_2142,N_2148);
nor U2301 (N_2301,N_2112,N_2125);
and U2302 (N_2302,N_2195,N_2148);
nor U2303 (N_2303,N_2085,N_2004);
or U2304 (N_2304,N_2018,N_2143);
or U2305 (N_2305,N_2097,N_2046);
and U2306 (N_2306,N_2145,N_2077);
and U2307 (N_2307,N_2151,N_2187);
or U2308 (N_2308,N_2028,N_2043);
xor U2309 (N_2309,N_2118,N_2140);
nor U2310 (N_2310,N_2103,N_2001);
nand U2311 (N_2311,N_2086,N_2165);
nor U2312 (N_2312,N_2059,N_2136);
nand U2313 (N_2313,N_2067,N_2093);
nor U2314 (N_2314,N_2041,N_2082);
xnor U2315 (N_2315,N_2095,N_2170);
nand U2316 (N_2316,N_2005,N_2034);
or U2317 (N_2317,N_2096,N_2037);
nand U2318 (N_2318,N_2028,N_2151);
xnor U2319 (N_2319,N_2097,N_2081);
nand U2320 (N_2320,N_2065,N_2093);
xor U2321 (N_2321,N_2190,N_2169);
and U2322 (N_2322,N_2145,N_2074);
nand U2323 (N_2323,N_2058,N_2107);
nand U2324 (N_2324,N_2015,N_2091);
and U2325 (N_2325,N_2100,N_2108);
xor U2326 (N_2326,N_2007,N_2019);
xnor U2327 (N_2327,N_2041,N_2003);
nor U2328 (N_2328,N_2173,N_2193);
xnor U2329 (N_2329,N_2145,N_2020);
and U2330 (N_2330,N_2004,N_2053);
nand U2331 (N_2331,N_2079,N_2091);
nand U2332 (N_2332,N_2139,N_2090);
xor U2333 (N_2333,N_2037,N_2178);
xnor U2334 (N_2334,N_2155,N_2142);
and U2335 (N_2335,N_2115,N_2102);
xnor U2336 (N_2336,N_2104,N_2184);
xnor U2337 (N_2337,N_2132,N_2123);
or U2338 (N_2338,N_2137,N_2158);
nand U2339 (N_2339,N_2039,N_2111);
and U2340 (N_2340,N_2160,N_2099);
and U2341 (N_2341,N_2004,N_2029);
nor U2342 (N_2342,N_2140,N_2066);
or U2343 (N_2343,N_2132,N_2042);
nand U2344 (N_2344,N_2062,N_2199);
xnor U2345 (N_2345,N_2056,N_2107);
or U2346 (N_2346,N_2060,N_2174);
nor U2347 (N_2347,N_2100,N_2171);
xnor U2348 (N_2348,N_2183,N_2108);
and U2349 (N_2349,N_2045,N_2118);
xnor U2350 (N_2350,N_2178,N_2121);
or U2351 (N_2351,N_2152,N_2175);
xor U2352 (N_2352,N_2068,N_2010);
and U2353 (N_2353,N_2144,N_2090);
nand U2354 (N_2354,N_2064,N_2055);
and U2355 (N_2355,N_2107,N_2015);
xnor U2356 (N_2356,N_2107,N_2105);
and U2357 (N_2357,N_2126,N_2052);
or U2358 (N_2358,N_2140,N_2152);
nand U2359 (N_2359,N_2070,N_2138);
nor U2360 (N_2360,N_2199,N_2103);
xor U2361 (N_2361,N_2088,N_2121);
nand U2362 (N_2362,N_2061,N_2003);
nand U2363 (N_2363,N_2108,N_2001);
or U2364 (N_2364,N_2133,N_2158);
nand U2365 (N_2365,N_2190,N_2020);
xor U2366 (N_2366,N_2177,N_2146);
nor U2367 (N_2367,N_2030,N_2134);
nand U2368 (N_2368,N_2066,N_2149);
xnor U2369 (N_2369,N_2045,N_2155);
or U2370 (N_2370,N_2186,N_2064);
nor U2371 (N_2371,N_2019,N_2173);
xor U2372 (N_2372,N_2117,N_2099);
nand U2373 (N_2373,N_2079,N_2153);
nor U2374 (N_2374,N_2088,N_2165);
or U2375 (N_2375,N_2163,N_2008);
xor U2376 (N_2376,N_2129,N_2123);
xnor U2377 (N_2377,N_2186,N_2130);
or U2378 (N_2378,N_2166,N_2154);
nor U2379 (N_2379,N_2155,N_2012);
nand U2380 (N_2380,N_2001,N_2138);
and U2381 (N_2381,N_2104,N_2001);
or U2382 (N_2382,N_2184,N_2002);
or U2383 (N_2383,N_2035,N_2171);
or U2384 (N_2384,N_2069,N_2080);
nand U2385 (N_2385,N_2023,N_2147);
and U2386 (N_2386,N_2160,N_2026);
nor U2387 (N_2387,N_2112,N_2168);
or U2388 (N_2388,N_2016,N_2058);
nand U2389 (N_2389,N_2198,N_2115);
nand U2390 (N_2390,N_2031,N_2187);
xnor U2391 (N_2391,N_2010,N_2069);
and U2392 (N_2392,N_2079,N_2178);
or U2393 (N_2393,N_2057,N_2149);
xor U2394 (N_2394,N_2018,N_2181);
nor U2395 (N_2395,N_2193,N_2035);
nand U2396 (N_2396,N_2098,N_2145);
nand U2397 (N_2397,N_2112,N_2105);
nor U2398 (N_2398,N_2183,N_2035);
nand U2399 (N_2399,N_2093,N_2112);
nand U2400 (N_2400,N_2293,N_2200);
xor U2401 (N_2401,N_2317,N_2385);
nand U2402 (N_2402,N_2361,N_2360);
or U2403 (N_2403,N_2233,N_2289);
or U2404 (N_2404,N_2377,N_2291);
xor U2405 (N_2405,N_2217,N_2335);
nand U2406 (N_2406,N_2374,N_2231);
nand U2407 (N_2407,N_2322,N_2255);
and U2408 (N_2408,N_2222,N_2206);
or U2409 (N_2409,N_2354,N_2333);
nor U2410 (N_2410,N_2353,N_2367);
or U2411 (N_2411,N_2337,N_2388);
xor U2412 (N_2412,N_2273,N_2286);
nand U2413 (N_2413,N_2307,N_2274);
xnor U2414 (N_2414,N_2323,N_2284);
or U2415 (N_2415,N_2341,N_2327);
nor U2416 (N_2416,N_2304,N_2209);
and U2417 (N_2417,N_2380,N_2292);
and U2418 (N_2418,N_2271,N_2305);
nor U2419 (N_2419,N_2275,N_2347);
or U2420 (N_2420,N_2202,N_2205);
nand U2421 (N_2421,N_2203,N_2296);
and U2422 (N_2422,N_2393,N_2373);
nand U2423 (N_2423,N_2269,N_2342);
nor U2424 (N_2424,N_2262,N_2207);
and U2425 (N_2425,N_2243,N_2316);
and U2426 (N_2426,N_2366,N_2257);
or U2427 (N_2427,N_2265,N_2208);
and U2428 (N_2428,N_2339,N_2219);
nand U2429 (N_2429,N_2364,N_2266);
nor U2430 (N_2430,N_2379,N_2301);
nor U2431 (N_2431,N_2389,N_2329);
and U2432 (N_2432,N_2378,N_2306);
or U2433 (N_2433,N_2370,N_2324);
nand U2434 (N_2434,N_2280,N_2282);
nor U2435 (N_2435,N_2314,N_2210);
xnor U2436 (N_2436,N_2214,N_2350);
or U2437 (N_2437,N_2254,N_2352);
nor U2438 (N_2438,N_2325,N_2259);
nor U2439 (N_2439,N_2235,N_2315);
nand U2440 (N_2440,N_2253,N_2295);
or U2441 (N_2441,N_2326,N_2264);
and U2442 (N_2442,N_2237,N_2281);
or U2443 (N_2443,N_2239,N_2220);
nand U2444 (N_2444,N_2270,N_2396);
nand U2445 (N_2445,N_2224,N_2363);
nand U2446 (N_2446,N_2319,N_2236);
nand U2447 (N_2447,N_2225,N_2228);
and U2448 (N_2448,N_2397,N_2332);
xnor U2449 (N_2449,N_2287,N_2276);
nand U2450 (N_2450,N_2371,N_2355);
or U2451 (N_2451,N_2362,N_2290);
nand U2452 (N_2452,N_2356,N_2232);
or U2453 (N_2453,N_2204,N_2390);
or U2454 (N_2454,N_2384,N_2376);
nor U2455 (N_2455,N_2343,N_2261);
nor U2456 (N_2456,N_2250,N_2387);
nand U2457 (N_2457,N_2391,N_2213);
nand U2458 (N_2458,N_2216,N_2234);
and U2459 (N_2459,N_2375,N_2212);
nand U2460 (N_2460,N_2398,N_2399);
and U2461 (N_2461,N_2340,N_2348);
nor U2462 (N_2462,N_2338,N_2382);
or U2463 (N_2463,N_2218,N_2300);
xnor U2464 (N_2464,N_2223,N_2369);
nand U2465 (N_2465,N_2331,N_2240);
and U2466 (N_2466,N_2238,N_2244);
and U2467 (N_2467,N_2365,N_2381);
nor U2468 (N_2468,N_2312,N_2351);
and U2469 (N_2469,N_2394,N_2395);
and U2470 (N_2470,N_2248,N_2349);
nor U2471 (N_2471,N_2318,N_2247);
and U2472 (N_2472,N_2260,N_2242);
nand U2473 (N_2473,N_2299,N_2336);
nand U2474 (N_2474,N_2368,N_2346);
nor U2475 (N_2475,N_2241,N_2201);
xor U2476 (N_2476,N_2230,N_2211);
or U2477 (N_2477,N_2256,N_2263);
or U2478 (N_2478,N_2311,N_2303);
xnor U2479 (N_2479,N_2258,N_2279);
and U2480 (N_2480,N_2267,N_2386);
xor U2481 (N_2481,N_2392,N_2345);
nor U2482 (N_2482,N_2229,N_2334);
and U2483 (N_2483,N_2320,N_2372);
nor U2484 (N_2484,N_2321,N_2283);
or U2485 (N_2485,N_2288,N_2294);
nor U2486 (N_2486,N_2226,N_2252);
or U2487 (N_2487,N_2251,N_2297);
or U2488 (N_2488,N_2215,N_2246);
or U2489 (N_2489,N_2227,N_2358);
nor U2490 (N_2490,N_2328,N_2298);
nand U2491 (N_2491,N_2383,N_2357);
and U2492 (N_2492,N_2268,N_2309);
and U2493 (N_2493,N_2278,N_2330);
xor U2494 (N_2494,N_2249,N_2313);
nand U2495 (N_2495,N_2221,N_2308);
xor U2496 (N_2496,N_2285,N_2359);
nand U2497 (N_2497,N_2310,N_2344);
xnor U2498 (N_2498,N_2272,N_2277);
xnor U2499 (N_2499,N_2302,N_2245);
and U2500 (N_2500,N_2347,N_2376);
xor U2501 (N_2501,N_2269,N_2267);
and U2502 (N_2502,N_2364,N_2240);
nand U2503 (N_2503,N_2282,N_2395);
nand U2504 (N_2504,N_2355,N_2236);
and U2505 (N_2505,N_2235,N_2363);
xnor U2506 (N_2506,N_2389,N_2264);
and U2507 (N_2507,N_2331,N_2302);
or U2508 (N_2508,N_2216,N_2350);
nand U2509 (N_2509,N_2333,N_2219);
or U2510 (N_2510,N_2301,N_2334);
nand U2511 (N_2511,N_2349,N_2391);
and U2512 (N_2512,N_2232,N_2345);
or U2513 (N_2513,N_2295,N_2390);
nand U2514 (N_2514,N_2202,N_2384);
and U2515 (N_2515,N_2250,N_2270);
nor U2516 (N_2516,N_2243,N_2235);
xor U2517 (N_2517,N_2285,N_2257);
xor U2518 (N_2518,N_2366,N_2275);
and U2519 (N_2519,N_2360,N_2288);
or U2520 (N_2520,N_2220,N_2234);
xnor U2521 (N_2521,N_2217,N_2314);
xor U2522 (N_2522,N_2313,N_2284);
nand U2523 (N_2523,N_2393,N_2350);
nor U2524 (N_2524,N_2327,N_2338);
or U2525 (N_2525,N_2200,N_2372);
xnor U2526 (N_2526,N_2319,N_2294);
or U2527 (N_2527,N_2383,N_2280);
and U2528 (N_2528,N_2280,N_2375);
xnor U2529 (N_2529,N_2379,N_2274);
or U2530 (N_2530,N_2302,N_2394);
or U2531 (N_2531,N_2377,N_2304);
nor U2532 (N_2532,N_2295,N_2209);
xor U2533 (N_2533,N_2281,N_2284);
and U2534 (N_2534,N_2320,N_2200);
and U2535 (N_2535,N_2281,N_2294);
or U2536 (N_2536,N_2396,N_2315);
or U2537 (N_2537,N_2339,N_2234);
nor U2538 (N_2538,N_2246,N_2306);
nand U2539 (N_2539,N_2221,N_2325);
nand U2540 (N_2540,N_2269,N_2380);
and U2541 (N_2541,N_2318,N_2336);
xnor U2542 (N_2542,N_2364,N_2330);
and U2543 (N_2543,N_2340,N_2343);
nor U2544 (N_2544,N_2279,N_2206);
xor U2545 (N_2545,N_2296,N_2220);
or U2546 (N_2546,N_2270,N_2214);
or U2547 (N_2547,N_2273,N_2217);
or U2548 (N_2548,N_2221,N_2306);
xnor U2549 (N_2549,N_2352,N_2274);
or U2550 (N_2550,N_2208,N_2324);
nand U2551 (N_2551,N_2276,N_2254);
or U2552 (N_2552,N_2377,N_2228);
nand U2553 (N_2553,N_2330,N_2381);
and U2554 (N_2554,N_2252,N_2329);
xnor U2555 (N_2555,N_2232,N_2201);
or U2556 (N_2556,N_2363,N_2339);
or U2557 (N_2557,N_2289,N_2320);
nor U2558 (N_2558,N_2332,N_2220);
xor U2559 (N_2559,N_2365,N_2379);
xnor U2560 (N_2560,N_2335,N_2307);
or U2561 (N_2561,N_2205,N_2259);
xnor U2562 (N_2562,N_2353,N_2204);
nor U2563 (N_2563,N_2382,N_2218);
xor U2564 (N_2564,N_2249,N_2326);
or U2565 (N_2565,N_2323,N_2290);
nor U2566 (N_2566,N_2385,N_2235);
or U2567 (N_2567,N_2336,N_2315);
xor U2568 (N_2568,N_2393,N_2225);
and U2569 (N_2569,N_2368,N_2388);
xor U2570 (N_2570,N_2211,N_2265);
and U2571 (N_2571,N_2386,N_2243);
nor U2572 (N_2572,N_2235,N_2278);
or U2573 (N_2573,N_2396,N_2285);
xor U2574 (N_2574,N_2238,N_2282);
nor U2575 (N_2575,N_2313,N_2282);
nor U2576 (N_2576,N_2381,N_2333);
and U2577 (N_2577,N_2341,N_2251);
and U2578 (N_2578,N_2205,N_2356);
and U2579 (N_2579,N_2394,N_2319);
xor U2580 (N_2580,N_2270,N_2254);
and U2581 (N_2581,N_2238,N_2268);
or U2582 (N_2582,N_2260,N_2222);
or U2583 (N_2583,N_2203,N_2293);
or U2584 (N_2584,N_2398,N_2357);
xnor U2585 (N_2585,N_2349,N_2290);
nand U2586 (N_2586,N_2390,N_2213);
or U2587 (N_2587,N_2275,N_2205);
nor U2588 (N_2588,N_2214,N_2297);
and U2589 (N_2589,N_2335,N_2237);
or U2590 (N_2590,N_2269,N_2207);
or U2591 (N_2591,N_2257,N_2215);
nor U2592 (N_2592,N_2356,N_2260);
or U2593 (N_2593,N_2202,N_2370);
nor U2594 (N_2594,N_2332,N_2340);
and U2595 (N_2595,N_2375,N_2309);
or U2596 (N_2596,N_2326,N_2391);
nand U2597 (N_2597,N_2382,N_2316);
or U2598 (N_2598,N_2261,N_2218);
nor U2599 (N_2599,N_2228,N_2260);
xnor U2600 (N_2600,N_2522,N_2561);
nor U2601 (N_2601,N_2415,N_2504);
and U2602 (N_2602,N_2462,N_2482);
xor U2603 (N_2603,N_2496,N_2527);
or U2604 (N_2604,N_2451,N_2525);
xnor U2605 (N_2605,N_2400,N_2446);
nand U2606 (N_2606,N_2480,N_2530);
or U2607 (N_2607,N_2521,N_2563);
nor U2608 (N_2608,N_2401,N_2539);
nor U2609 (N_2609,N_2403,N_2544);
or U2610 (N_2610,N_2487,N_2404);
nor U2611 (N_2611,N_2586,N_2590);
nand U2612 (N_2612,N_2442,N_2471);
nor U2613 (N_2613,N_2440,N_2558);
or U2614 (N_2614,N_2470,N_2531);
nand U2615 (N_2615,N_2536,N_2515);
xnor U2616 (N_2616,N_2594,N_2540);
nand U2617 (N_2617,N_2421,N_2479);
and U2618 (N_2618,N_2455,N_2503);
xnor U2619 (N_2619,N_2551,N_2562);
and U2620 (N_2620,N_2587,N_2464);
and U2621 (N_2621,N_2565,N_2460);
or U2622 (N_2622,N_2444,N_2494);
xnor U2623 (N_2623,N_2454,N_2488);
or U2624 (N_2624,N_2474,N_2567);
or U2625 (N_2625,N_2578,N_2445);
or U2626 (N_2626,N_2513,N_2577);
and U2627 (N_2627,N_2437,N_2493);
nand U2628 (N_2628,N_2484,N_2598);
xnor U2629 (N_2629,N_2417,N_2433);
or U2630 (N_2630,N_2461,N_2523);
or U2631 (N_2631,N_2599,N_2507);
xor U2632 (N_2632,N_2436,N_2429);
and U2633 (N_2633,N_2495,N_2447);
nor U2634 (N_2634,N_2456,N_2423);
xor U2635 (N_2635,N_2508,N_2443);
nand U2636 (N_2636,N_2512,N_2579);
nand U2637 (N_2637,N_2505,N_2549);
and U2638 (N_2638,N_2427,N_2426);
nor U2639 (N_2639,N_2407,N_2477);
nor U2640 (N_2640,N_2490,N_2459);
nand U2641 (N_2641,N_2431,N_2564);
and U2642 (N_2642,N_2492,N_2408);
or U2643 (N_2643,N_2411,N_2518);
or U2644 (N_2644,N_2458,N_2406);
nor U2645 (N_2645,N_2405,N_2448);
xor U2646 (N_2646,N_2580,N_2542);
nor U2647 (N_2647,N_2535,N_2498);
or U2648 (N_2648,N_2468,N_2418);
nand U2649 (N_2649,N_2425,N_2597);
xnor U2650 (N_2650,N_2574,N_2571);
nand U2651 (N_2651,N_2424,N_2478);
and U2652 (N_2652,N_2572,N_2420);
nor U2653 (N_2653,N_2560,N_2452);
or U2654 (N_2654,N_2547,N_2486);
and U2655 (N_2655,N_2559,N_2534);
and U2656 (N_2656,N_2416,N_2485);
and U2657 (N_2657,N_2491,N_2595);
nand U2658 (N_2658,N_2533,N_2457);
and U2659 (N_2659,N_2581,N_2463);
nand U2660 (N_2660,N_2538,N_2435);
nand U2661 (N_2661,N_2532,N_2541);
xor U2662 (N_2662,N_2556,N_2511);
nor U2663 (N_2663,N_2501,N_2410);
or U2664 (N_2664,N_2509,N_2517);
nor U2665 (N_2665,N_2412,N_2575);
xnor U2666 (N_2666,N_2514,N_2573);
nor U2667 (N_2667,N_2550,N_2537);
xnor U2668 (N_2668,N_2466,N_2584);
nand U2669 (N_2669,N_2543,N_2510);
nor U2670 (N_2670,N_2583,N_2545);
nor U2671 (N_2671,N_2481,N_2409);
nand U2672 (N_2672,N_2566,N_2570);
nand U2673 (N_2673,N_2472,N_2502);
xnor U2674 (N_2674,N_2500,N_2546);
xor U2675 (N_2675,N_2438,N_2473);
nand U2676 (N_2676,N_2548,N_2589);
or U2677 (N_2677,N_2419,N_2476);
and U2678 (N_2678,N_2467,N_2439);
and U2679 (N_2679,N_2520,N_2569);
xor U2680 (N_2680,N_2434,N_2576);
and U2681 (N_2681,N_2428,N_2402);
xnor U2682 (N_2682,N_2475,N_2588);
or U2683 (N_2683,N_2552,N_2568);
nor U2684 (N_2684,N_2489,N_2483);
xor U2685 (N_2685,N_2593,N_2554);
nor U2686 (N_2686,N_2582,N_2506);
nor U2687 (N_2687,N_2592,N_2453);
nor U2688 (N_2688,N_2469,N_2524);
and U2689 (N_2689,N_2499,N_2465);
xnor U2690 (N_2690,N_2413,N_2555);
nand U2691 (N_2691,N_2432,N_2528);
nand U2692 (N_2692,N_2553,N_2591);
or U2693 (N_2693,N_2449,N_2422);
nor U2694 (N_2694,N_2450,N_2526);
and U2695 (N_2695,N_2497,N_2516);
and U2696 (N_2696,N_2596,N_2430);
nand U2697 (N_2697,N_2519,N_2557);
xor U2698 (N_2698,N_2414,N_2529);
xor U2699 (N_2699,N_2441,N_2585);
or U2700 (N_2700,N_2400,N_2437);
xnor U2701 (N_2701,N_2571,N_2573);
xor U2702 (N_2702,N_2504,N_2470);
nor U2703 (N_2703,N_2533,N_2523);
nand U2704 (N_2704,N_2535,N_2428);
and U2705 (N_2705,N_2575,N_2595);
or U2706 (N_2706,N_2570,N_2409);
or U2707 (N_2707,N_2455,N_2450);
nor U2708 (N_2708,N_2426,N_2592);
nand U2709 (N_2709,N_2408,N_2581);
nor U2710 (N_2710,N_2522,N_2433);
nor U2711 (N_2711,N_2428,N_2404);
nor U2712 (N_2712,N_2491,N_2486);
or U2713 (N_2713,N_2563,N_2568);
nor U2714 (N_2714,N_2495,N_2411);
and U2715 (N_2715,N_2420,N_2596);
and U2716 (N_2716,N_2494,N_2511);
nor U2717 (N_2717,N_2462,N_2503);
xnor U2718 (N_2718,N_2461,N_2418);
nand U2719 (N_2719,N_2432,N_2409);
nand U2720 (N_2720,N_2480,N_2427);
or U2721 (N_2721,N_2526,N_2595);
or U2722 (N_2722,N_2565,N_2478);
nor U2723 (N_2723,N_2441,N_2502);
or U2724 (N_2724,N_2515,N_2444);
nand U2725 (N_2725,N_2593,N_2599);
xnor U2726 (N_2726,N_2455,N_2562);
nand U2727 (N_2727,N_2454,N_2485);
or U2728 (N_2728,N_2586,N_2550);
nor U2729 (N_2729,N_2424,N_2488);
nand U2730 (N_2730,N_2464,N_2535);
nor U2731 (N_2731,N_2505,N_2437);
nor U2732 (N_2732,N_2568,N_2553);
and U2733 (N_2733,N_2426,N_2522);
nor U2734 (N_2734,N_2575,N_2513);
and U2735 (N_2735,N_2513,N_2550);
or U2736 (N_2736,N_2421,N_2461);
or U2737 (N_2737,N_2469,N_2422);
and U2738 (N_2738,N_2450,N_2469);
nand U2739 (N_2739,N_2408,N_2570);
nand U2740 (N_2740,N_2508,N_2402);
or U2741 (N_2741,N_2567,N_2448);
or U2742 (N_2742,N_2492,N_2404);
or U2743 (N_2743,N_2467,N_2426);
xor U2744 (N_2744,N_2459,N_2516);
nand U2745 (N_2745,N_2596,N_2478);
nand U2746 (N_2746,N_2589,N_2435);
xor U2747 (N_2747,N_2515,N_2428);
nor U2748 (N_2748,N_2568,N_2572);
nor U2749 (N_2749,N_2516,N_2455);
and U2750 (N_2750,N_2498,N_2450);
or U2751 (N_2751,N_2430,N_2433);
nor U2752 (N_2752,N_2549,N_2513);
xor U2753 (N_2753,N_2443,N_2493);
or U2754 (N_2754,N_2412,N_2450);
and U2755 (N_2755,N_2531,N_2435);
or U2756 (N_2756,N_2475,N_2459);
nand U2757 (N_2757,N_2575,N_2564);
and U2758 (N_2758,N_2532,N_2578);
and U2759 (N_2759,N_2496,N_2567);
xor U2760 (N_2760,N_2407,N_2481);
xnor U2761 (N_2761,N_2523,N_2517);
xor U2762 (N_2762,N_2502,N_2544);
nand U2763 (N_2763,N_2522,N_2437);
nor U2764 (N_2764,N_2450,N_2417);
xor U2765 (N_2765,N_2582,N_2547);
or U2766 (N_2766,N_2540,N_2419);
and U2767 (N_2767,N_2489,N_2554);
xor U2768 (N_2768,N_2519,N_2585);
nor U2769 (N_2769,N_2485,N_2497);
and U2770 (N_2770,N_2480,N_2505);
nor U2771 (N_2771,N_2463,N_2570);
xnor U2772 (N_2772,N_2534,N_2572);
nand U2773 (N_2773,N_2566,N_2446);
nor U2774 (N_2774,N_2454,N_2564);
and U2775 (N_2775,N_2587,N_2407);
xnor U2776 (N_2776,N_2490,N_2403);
or U2777 (N_2777,N_2554,N_2482);
xnor U2778 (N_2778,N_2431,N_2497);
nor U2779 (N_2779,N_2401,N_2523);
and U2780 (N_2780,N_2468,N_2524);
xor U2781 (N_2781,N_2460,N_2543);
and U2782 (N_2782,N_2473,N_2417);
nand U2783 (N_2783,N_2488,N_2451);
nand U2784 (N_2784,N_2476,N_2575);
nand U2785 (N_2785,N_2403,N_2482);
nand U2786 (N_2786,N_2494,N_2505);
or U2787 (N_2787,N_2570,N_2429);
and U2788 (N_2788,N_2523,N_2464);
nand U2789 (N_2789,N_2413,N_2462);
or U2790 (N_2790,N_2566,N_2448);
xnor U2791 (N_2791,N_2513,N_2492);
or U2792 (N_2792,N_2565,N_2528);
or U2793 (N_2793,N_2420,N_2483);
or U2794 (N_2794,N_2582,N_2445);
nor U2795 (N_2795,N_2547,N_2545);
and U2796 (N_2796,N_2592,N_2553);
or U2797 (N_2797,N_2447,N_2411);
xor U2798 (N_2798,N_2452,N_2463);
nor U2799 (N_2799,N_2415,N_2436);
or U2800 (N_2800,N_2611,N_2712);
or U2801 (N_2801,N_2795,N_2670);
nor U2802 (N_2802,N_2605,N_2706);
nor U2803 (N_2803,N_2661,N_2627);
nand U2804 (N_2804,N_2601,N_2690);
xnor U2805 (N_2805,N_2681,N_2776);
xor U2806 (N_2806,N_2651,N_2607);
or U2807 (N_2807,N_2756,N_2677);
nand U2808 (N_2808,N_2784,N_2610);
and U2809 (N_2809,N_2672,N_2727);
xnor U2810 (N_2810,N_2632,N_2780);
nand U2811 (N_2811,N_2694,N_2705);
nor U2812 (N_2812,N_2680,N_2768);
nand U2813 (N_2813,N_2732,N_2631);
xnor U2814 (N_2814,N_2799,N_2783);
or U2815 (N_2815,N_2613,N_2642);
nor U2816 (N_2816,N_2709,N_2778);
nand U2817 (N_2817,N_2774,N_2621);
nor U2818 (N_2818,N_2630,N_2603);
nand U2819 (N_2819,N_2798,N_2794);
or U2820 (N_2820,N_2618,N_2796);
xnor U2821 (N_2821,N_2793,N_2791);
nand U2822 (N_2822,N_2788,N_2708);
or U2823 (N_2823,N_2753,N_2655);
nand U2824 (N_2824,N_2759,N_2702);
nand U2825 (N_2825,N_2781,N_2682);
nand U2826 (N_2826,N_2638,N_2609);
or U2827 (N_2827,N_2634,N_2792);
or U2828 (N_2828,N_2738,N_2723);
nor U2829 (N_2829,N_2637,N_2782);
or U2830 (N_2830,N_2648,N_2724);
or U2831 (N_2831,N_2664,N_2710);
and U2832 (N_2832,N_2720,N_2676);
nor U2833 (N_2833,N_2692,N_2742);
xnor U2834 (N_2834,N_2764,N_2711);
nand U2835 (N_2835,N_2766,N_2612);
or U2836 (N_2836,N_2743,N_2725);
and U2837 (N_2837,N_2622,N_2674);
nand U2838 (N_2838,N_2721,N_2750);
nor U2839 (N_2839,N_2739,N_2729);
nor U2840 (N_2840,N_2640,N_2633);
and U2841 (N_2841,N_2666,N_2704);
nor U2842 (N_2842,N_2624,N_2779);
or U2843 (N_2843,N_2737,N_2652);
or U2844 (N_2844,N_2660,N_2735);
or U2845 (N_2845,N_2647,N_2669);
or U2846 (N_2846,N_2718,N_2678);
or U2847 (N_2847,N_2726,N_2656);
and U2848 (N_2848,N_2626,N_2697);
xnor U2849 (N_2849,N_2635,N_2758);
nand U2850 (N_2850,N_2698,N_2604);
nor U2851 (N_2851,N_2600,N_2688);
xor U2852 (N_2852,N_2675,N_2608);
nor U2853 (N_2853,N_2749,N_2645);
or U2854 (N_2854,N_2773,N_2644);
nand U2855 (N_2855,N_2614,N_2696);
nor U2856 (N_2856,N_2734,N_2789);
and U2857 (N_2857,N_2767,N_2747);
or U2858 (N_2858,N_2728,N_2763);
or U2859 (N_2859,N_2667,N_2719);
or U2860 (N_2860,N_2636,N_2639);
xor U2861 (N_2861,N_2701,N_2699);
nor U2862 (N_2862,N_2746,N_2716);
and U2863 (N_2863,N_2751,N_2785);
xor U2864 (N_2864,N_2663,N_2748);
and U2865 (N_2865,N_2684,N_2700);
nand U2866 (N_2866,N_2760,N_2730);
or U2867 (N_2867,N_2685,N_2617);
or U2868 (N_2868,N_2679,N_2703);
or U2869 (N_2869,N_2770,N_2687);
and U2870 (N_2870,N_2659,N_2755);
xnor U2871 (N_2871,N_2654,N_2722);
nand U2872 (N_2872,N_2736,N_2741);
nor U2873 (N_2873,N_2745,N_2715);
xnor U2874 (N_2874,N_2673,N_2713);
xnor U2875 (N_2875,N_2740,N_2797);
xor U2876 (N_2876,N_2683,N_2641);
nand U2877 (N_2877,N_2744,N_2646);
or U2878 (N_2878,N_2620,N_2777);
xor U2879 (N_2879,N_2762,N_2765);
nand U2880 (N_2880,N_2790,N_2689);
and U2881 (N_2881,N_2733,N_2619);
xor U2882 (N_2882,N_2769,N_2658);
or U2883 (N_2883,N_2629,N_2714);
and U2884 (N_2884,N_2771,N_2668);
xor U2885 (N_2885,N_2649,N_2671);
xnor U2886 (N_2886,N_2625,N_2693);
xnor U2887 (N_2887,N_2691,N_2623);
xnor U2888 (N_2888,N_2628,N_2752);
nand U2889 (N_2889,N_2787,N_2657);
or U2890 (N_2890,N_2731,N_2653);
and U2891 (N_2891,N_2786,N_2615);
nand U2892 (N_2892,N_2662,N_2754);
and U2893 (N_2893,N_2602,N_2757);
or U2894 (N_2894,N_2775,N_2643);
or U2895 (N_2895,N_2686,N_2695);
nand U2896 (N_2896,N_2717,N_2707);
or U2897 (N_2897,N_2761,N_2606);
xor U2898 (N_2898,N_2772,N_2665);
or U2899 (N_2899,N_2650,N_2616);
nand U2900 (N_2900,N_2723,N_2660);
and U2901 (N_2901,N_2632,N_2704);
xor U2902 (N_2902,N_2652,N_2739);
or U2903 (N_2903,N_2713,N_2781);
xnor U2904 (N_2904,N_2758,N_2741);
nor U2905 (N_2905,N_2636,N_2642);
xor U2906 (N_2906,N_2782,N_2609);
and U2907 (N_2907,N_2736,N_2717);
nor U2908 (N_2908,N_2767,N_2718);
nor U2909 (N_2909,N_2608,N_2761);
nand U2910 (N_2910,N_2708,N_2737);
nor U2911 (N_2911,N_2605,N_2717);
nand U2912 (N_2912,N_2682,N_2641);
and U2913 (N_2913,N_2719,N_2771);
nand U2914 (N_2914,N_2629,N_2774);
or U2915 (N_2915,N_2668,N_2794);
xnor U2916 (N_2916,N_2723,N_2748);
or U2917 (N_2917,N_2757,N_2691);
nor U2918 (N_2918,N_2795,N_2766);
nand U2919 (N_2919,N_2630,N_2771);
nand U2920 (N_2920,N_2760,N_2676);
xnor U2921 (N_2921,N_2733,N_2618);
nand U2922 (N_2922,N_2697,N_2682);
xor U2923 (N_2923,N_2765,N_2794);
or U2924 (N_2924,N_2721,N_2751);
nor U2925 (N_2925,N_2727,N_2779);
nor U2926 (N_2926,N_2774,N_2733);
nor U2927 (N_2927,N_2666,N_2744);
xnor U2928 (N_2928,N_2682,N_2618);
nand U2929 (N_2929,N_2684,N_2760);
or U2930 (N_2930,N_2786,N_2678);
and U2931 (N_2931,N_2625,N_2632);
or U2932 (N_2932,N_2608,N_2747);
xnor U2933 (N_2933,N_2725,N_2689);
nand U2934 (N_2934,N_2793,N_2755);
nand U2935 (N_2935,N_2648,N_2695);
and U2936 (N_2936,N_2693,N_2627);
nor U2937 (N_2937,N_2780,N_2706);
xnor U2938 (N_2938,N_2632,N_2786);
xnor U2939 (N_2939,N_2779,N_2692);
nor U2940 (N_2940,N_2735,N_2640);
and U2941 (N_2941,N_2679,N_2618);
nor U2942 (N_2942,N_2614,N_2693);
or U2943 (N_2943,N_2657,N_2778);
nor U2944 (N_2944,N_2741,N_2699);
or U2945 (N_2945,N_2788,N_2743);
or U2946 (N_2946,N_2777,N_2701);
nand U2947 (N_2947,N_2643,N_2687);
xor U2948 (N_2948,N_2784,N_2794);
or U2949 (N_2949,N_2770,N_2670);
nand U2950 (N_2950,N_2731,N_2671);
xnor U2951 (N_2951,N_2636,N_2653);
xnor U2952 (N_2952,N_2685,N_2603);
and U2953 (N_2953,N_2719,N_2689);
nor U2954 (N_2954,N_2711,N_2718);
and U2955 (N_2955,N_2725,N_2733);
xnor U2956 (N_2956,N_2657,N_2607);
nand U2957 (N_2957,N_2751,N_2675);
nor U2958 (N_2958,N_2685,N_2735);
xor U2959 (N_2959,N_2661,N_2607);
and U2960 (N_2960,N_2718,N_2731);
or U2961 (N_2961,N_2645,N_2626);
or U2962 (N_2962,N_2690,N_2647);
nand U2963 (N_2963,N_2704,N_2780);
xnor U2964 (N_2964,N_2772,N_2743);
or U2965 (N_2965,N_2788,N_2707);
and U2966 (N_2966,N_2636,N_2798);
nor U2967 (N_2967,N_2746,N_2675);
or U2968 (N_2968,N_2650,N_2720);
xnor U2969 (N_2969,N_2669,N_2639);
and U2970 (N_2970,N_2669,N_2792);
nor U2971 (N_2971,N_2744,N_2796);
xor U2972 (N_2972,N_2683,N_2662);
nor U2973 (N_2973,N_2744,N_2709);
nand U2974 (N_2974,N_2646,N_2628);
nand U2975 (N_2975,N_2652,N_2673);
or U2976 (N_2976,N_2716,N_2690);
nand U2977 (N_2977,N_2691,N_2743);
and U2978 (N_2978,N_2754,N_2671);
xnor U2979 (N_2979,N_2701,N_2760);
or U2980 (N_2980,N_2639,N_2702);
xor U2981 (N_2981,N_2665,N_2661);
nand U2982 (N_2982,N_2721,N_2701);
nand U2983 (N_2983,N_2743,N_2606);
xnor U2984 (N_2984,N_2771,N_2700);
xnor U2985 (N_2985,N_2738,N_2626);
or U2986 (N_2986,N_2707,N_2756);
xor U2987 (N_2987,N_2725,N_2760);
and U2988 (N_2988,N_2682,N_2723);
or U2989 (N_2989,N_2678,N_2743);
or U2990 (N_2990,N_2715,N_2724);
and U2991 (N_2991,N_2669,N_2675);
and U2992 (N_2992,N_2625,N_2600);
xnor U2993 (N_2993,N_2649,N_2700);
nand U2994 (N_2994,N_2641,N_2735);
nor U2995 (N_2995,N_2628,N_2660);
nor U2996 (N_2996,N_2676,N_2728);
or U2997 (N_2997,N_2695,N_2631);
xnor U2998 (N_2998,N_2706,N_2711);
nor U2999 (N_2999,N_2620,N_2642);
nand U3000 (N_3000,N_2894,N_2853);
nand U3001 (N_3001,N_2833,N_2839);
or U3002 (N_3002,N_2913,N_2859);
xor U3003 (N_3003,N_2994,N_2960);
or U3004 (N_3004,N_2841,N_2980);
nor U3005 (N_3005,N_2826,N_2945);
xor U3006 (N_3006,N_2879,N_2831);
xor U3007 (N_3007,N_2969,N_2810);
nand U3008 (N_3008,N_2992,N_2849);
xnor U3009 (N_3009,N_2857,N_2896);
or U3010 (N_3010,N_2961,N_2889);
and U3011 (N_3011,N_2997,N_2865);
xnor U3012 (N_3012,N_2972,N_2918);
and U3013 (N_3013,N_2866,N_2931);
or U3014 (N_3014,N_2912,N_2802);
nor U3015 (N_3015,N_2953,N_2858);
xnor U3016 (N_3016,N_2883,N_2902);
or U3017 (N_3017,N_2814,N_2808);
nand U3018 (N_3018,N_2964,N_2806);
xnor U3019 (N_3019,N_2856,N_2996);
nand U3020 (N_3020,N_2904,N_2929);
xor U3021 (N_3021,N_2962,N_2899);
and U3022 (N_3022,N_2967,N_2932);
nand U3023 (N_3023,N_2876,N_2936);
and U3024 (N_3024,N_2812,N_2872);
or U3025 (N_3025,N_2923,N_2877);
or U3026 (N_3026,N_2917,N_2854);
xnor U3027 (N_3027,N_2978,N_2875);
nand U3028 (N_3028,N_2966,N_2855);
nand U3029 (N_3029,N_2890,N_2801);
nor U3030 (N_3030,N_2867,N_2942);
or U3031 (N_3031,N_2829,N_2914);
and U3032 (N_3032,N_2934,N_2959);
or U3033 (N_3033,N_2830,N_2882);
nor U3034 (N_3034,N_2800,N_2916);
and U3035 (N_3035,N_2892,N_2989);
or U3036 (N_3036,N_2821,N_2956);
nor U3037 (N_3037,N_2911,N_2958);
nand U3038 (N_3038,N_2925,N_2905);
and U3039 (N_3039,N_2847,N_2926);
xnor U3040 (N_3040,N_2817,N_2982);
nor U3041 (N_3041,N_2888,N_2837);
xor U3042 (N_3042,N_2868,N_2840);
or U3043 (N_3043,N_2822,N_2921);
or U3044 (N_3044,N_2977,N_2907);
nand U3045 (N_3045,N_2878,N_2993);
nand U3046 (N_3046,N_2995,N_2954);
and U3047 (N_3047,N_2842,N_2844);
or U3048 (N_3048,N_2825,N_2971);
or U3049 (N_3049,N_2818,N_2940);
and U3050 (N_3050,N_2968,N_2887);
nor U3051 (N_3051,N_2986,N_2828);
xor U3052 (N_3052,N_2909,N_2947);
or U3053 (N_3053,N_2815,N_2943);
nand U3054 (N_3054,N_2860,N_2846);
nor U3055 (N_3055,N_2852,N_2937);
xnor U3056 (N_3056,N_2990,N_2924);
and U3057 (N_3057,N_2948,N_2927);
nor U3058 (N_3058,N_2938,N_2803);
nand U3059 (N_3059,N_2957,N_2933);
xor U3060 (N_3060,N_2979,N_2949);
xnor U3061 (N_3061,N_2900,N_2898);
or U3062 (N_3062,N_2998,N_2885);
and U3063 (N_3063,N_2819,N_2910);
nand U3064 (N_3064,N_2871,N_2955);
nor U3065 (N_3065,N_2893,N_2862);
or U3066 (N_3066,N_2824,N_2809);
nor U3067 (N_3067,N_2816,N_2930);
and U3068 (N_3068,N_2811,N_2988);
nor U3069 (N_3069,N_2906,N_2946);
nand U3070 (N_3070,N_2935,N_2981);
and U3071 (N_3071,N_2835,N_2970);
nor U3072 (N_3072,N_2908,N_2991);
xor U3073 (N_3073,N_2845,N_2919);
nand U3074 (N_3074,N_2832,N_2928);
nand U3075 (N_3075,N_2941,N_2874);
xor U3076 (N_3076,N_2880,N_2950);
nand U3077 (N_3077,N_2965,N_2985);
and U3078 (N_3078,N_2861,N_2983);
and U3079 (N_3079,N_2820,N_2975);
nand U3080 (N_3080,N_2886,N_2895);
and U3081 (N_3081,N_2813,N_2974);
and U3082 (N_3082,N_2884,N_2963);
nor U3083 (N_3083,N_2897,N_2987);
xnor U3084 (N_3084,N_2863,N_2976);
nor U3085 (N_3085,N_2891,N_2851);
nand U3086 (N_3086,N_2807,N_2901);
xnor U3087 (N_3087,N_2903,N_2834);
xor U3088 (N_3088,N_2973,N_2939);
xnor U3089 (N_3089,N_2920,N_2869);
and U3090 (N_3090,N_2999,N_2843);
xnor U3091 (N_3091,N_2915,N_2870);
xnor U3092 (N_3092,N_2864,N_2823);
or U3093 (N_3093,N_2836,N_2838);
nor U3094 (N_3094,N_2827,N_2944);
or U3095 (N_3095,N_2984,N_2804);
and U3096 (N_3096,N_2848,N_2881);
nand U3097 (N_3097,N_2952,N_2951);
and U3098 (N_3098,N_2922,N_2873);
xor U3099 (N_3099,N_2850,N_2805);
and U3100 (N_3100,N_2924,N_2956);
xor U3101 (N_3101,N_2907,N_2962);
nor U3102 (N_3102,N_2934,N_2873);
or U3103 (N_3103,N_2896,N_2898);
nor U3104 (N_3104,N_2816,N_2983);
and U3105 (N_3105,N_2911,N_2821);
nor U3106 (N_3106,N_2832,N_2883);
nand U3107 (N_3107,N_2844,N_2982);
and U3108 (N_3108,N_2928,N_2823);
xor U3109 (N_3109,N_2888,N_2804);
nor U3110 (N_3110,N_2818,N_2809);
or U3111 (N_3111,N_2944,N_2885);
nor U3112 (N_3112,N_2845,N_2882);
nor U3113 (N_3113,N_2995,N_2884);
xor U3114 (N_3114,N_2904,N_2890);
nor U3115 (N_3115,N_2936,N_2832);
nor U3116 (N_3116,N_2804,N_2811);
nand U3117 (N_3117,N_2832,N_2994);
nor U3118 (N_3118,N_2938,N_2944);
nand U3119 (N_3119,N_2853,N_2998);
xor U3120 (N_3120,N_2911,N_2868);
and U3121 (N_3121,N_2973,N_2875);
xnor U3122 (N_3122,N_2981,N_2952);
or U3123 (N_3123,N_2938,N_2987);
or U3124 (N_3124,N_2932,N_2943);
and U3125 (N_3125,N_2817,N_2845);
xor U3126 (N_3126,N_2839,N_2956);
nand U3127 (N_3127,N_2863,N_2887);
nor U3128 (N_3128,N_2879,N_2886);
and U3129 (N_3129,N_2937,N_2917);
xnor U3130 (N_3130,N_2893,N_2953);
nor U3131 (N_3131,N_2937,N_2835);
or U3132 (N_3132,N_2907,N_2827);
or U3133 (N_3133,N_2845,N_2956);
nand U3134 (N_3134,N_2918,N_2860);
nor U3135 (N_3135,N_2996,N_2843);
or U3136 (N_3136,N_2873,N_2930);
or U3137 (N_3137,N_2831,N_2800);
xnor U3138 (N_3138,N_2997,N_2849);
and U3139 (N_3139,N_2999,N_2955);
xor U3140 (N_3140,N_2806,N_2997);
or U3141 (N_3141,N_2853,N_2905);
and U3142 (N_3142,N_2857,N_2922);
nor U3143 (N_3143,N_2862,N_2869);
xnor U3144 (N_3144,N_2925,N_2822);
nor U3145 (N_3145,N_2851,N_2854);
xor U3146 (N_3146,N_2970,N_2918);
nor U3147 (N_3147,N_2939,N_2909);
or U3148 (N_3148,N_2854,N_2963);
nand U3149 (N_3149,N_2876,N_2923);
nand U3150 (N_3150,N_2824,N_2818);
nand U3151 (N_3151,N_2966,N_2939);
or U3152 (N_3152,N_2858,N_2906);
or U3153 (N_3153,N_2896,N_2946);
xor U3154 (N_3154,N_2862,N_2952);
xor U3155 (N_3155,N_2827,N_2982);
nand U3156 (N_3156,N_2810,N_2908);
and U3157 (N_3157,N_2920,N_2842);
xor U3158 (N_3158,N_2932,N_2869);
and U3159 (N_3159,N_2885,N_2928);
xnor U3160 (N_3160,N_2944,N_2932);
xor U3161 (N_3161,N_2890,N_2883);
nor U3162 (N_3162,N_2847,N_2870);
nand U3163 (N_3163,N_2840,N_2804);
nand U3164 (N_3164,N_2980,N_2847);
or U3165 (N_3165,N_2830,N_2958);
nand U3166 (N_3166,N_2963,N_2908);
nor U3167 (N_3167,N_2810,N_2824);
or U3168 (N_3168,N_2991,N_2813);
or U3169 (N_3169,N_2858,N_2984);
xor U3170 (N_3170,N_2844,N_2938);
xnor U3171 (N_3171,N_2875,N_2815);
or U3172 (N_3172,N_2851,N_2950);
xor U3173 (N_3173,N_2833,N_2899);
xor U3174 (N_3174,N_2949,N_2919);
or U3175 (N_3175,N_2847,N_2819);
and U3176 (N_3176,N_2884,N_2924);
nand U3177 (N_3177,N_2908,N_2986);
nand U3178 (N_3178,N_2976,N_2907);
nor U3179 (N_3179,N_2997,N_2903);
or U3180 (N_3180,N_2994,N_2993);
xor U3181 (N_3181,N_2933,N_2825);
and U3182 (N_3182,N_2824,N_2933);
nor U3183 (N_3183,N_2992,N_2969);
or U3184 (N_3184,N_2846,N_2978);
or U3185 (N_3185,N_2988,N_2928);
nand U3186 (N_3186,N_2925,N_2848);
or U3187 (N_3187,N_2830,N_2881);
or U3188 (N_3188,N_2843,N_2910);
or U3189 (N_3189,N_2888,N_2897);
and U3190 (N_3190,N_2915,N_2814);
or U3191 (N_3191,N_2938,N_2830);
nor U3192 (N_3192,N_2864,N_2964);
nand U3193 (N_3193,N_2882,N_2907);
nor U3194 (N_3194,N_2805,N_2881);
nand U3195 (N_3195,N_2809,N_2916);
nor U3196 (N_3196,N_2839,N_2868);
and U3197 (N_3197,N_2928,N_2883);
xnor U3198 (N_3198,N_2945,N_2948);
and U3199 (N_3199,N_2964,N_2871);
nand U3200 (N_3200,N_3098,N_3052);
nand U3201 (N_3201,N_3038,N_3110);
nand U3202 (N_3202,N_3127,N_3049);
xnor U3203 (N_3203,N_3036,N_3149);
nand U3204 (N_3204,N_3175,N_3022);
and U3205 (N_3205,N_3160,N_3062);
and U3206 (N_3206,N_3164,N_3088);
nand U3207 (N_3207,N_3042,N_3179);
nor U3208 (N_3208,N_3124,N_3167);
xor U3209 (N_3209,N_3025,N_3172);
nand U3210 (N_3210,N_3067,N_3093);
nor U3211 (N_3211,N_3058,N_3123);
xor U3212 (N_3212,N_3059,N_3181);
nor U3213 (N_3213,N_3078,N_3010);
xnor U3214 (N_3214,N_3112,N_3156);
nor U3215 (N_3215,N_3136,N_3171);
nor U3216 (N_3216,N_3084,N_3008);
nand U3217 (N_3217,N_3105,N_3162);
nand U3218 (N_3218,N_3044,N_3122);
or U3219 (N_3219,N_3026,N_3033);
and U3220 (N_3220,N_3125,N_3054);
xor U3221 (N_3221,N_3007,N_3050);
or U3222 (N_3222,N_3144,N_3103);
nand U3223 (N_3223,N_3109,N_3192);
and U3224 (N_3224,N_3090,N_3170);
xor U3225 (N_3225,N_3014,N_3154);
nor U3226 (N_3226,N_3047,N_3186);
and U3227 (N_3227,N_3194,N_3151);
xor U3228 (N_3228,N_3002,N_3064);
nor U3229 (N_3229,N_3121,N_3094);
and U3230 (N_3230,N_3030,N_3005);
and U3231 (N_3231,N_3120,N_3161);
and U3232 (N_3232,N_3029,N_3081);
and U3233 (N_3233,N_3043,N_3079);
xor U3234 (N_3234,N_3126,N_3015);
and U3235 (N_3235,N_3101,N_3066);
and U3236 (N_3236,N_3119,N_3063);
or U3237 (N_3237,N_3150,N_3017);
and U3238 (N_3238,N_3193,N_3184);
and U3239 (N_3239,N_3074,N_3100);
nand U3240 (N_3240,N_3189,N_3028);
xor U3241 (N_3241,N_3020,N_3113);
or U3242 (N_3242,N_3152,N_3096);
xor U3243 (N_3243,N_3041,N_3141);
and U3244 (N_3244,N_3140,N_3039);
or U3245 (N_3245,N_3155,N_3012);
or U3246 (N_3246,N_3177,N_3048);
or U3247 (N_3247,N_3013,N_3191);
or U3248 (N_3248,N_3190,N_3024);
or U3249 (N_3249,N_3000,N_3114);
xnor U3250 (N_3250,N_3023,N_3130);
xor U3251 (N_3251,N_3053,N_3055);
xor U3252 (N_3252,N_3158,N_3045);
xnor U3253 (N_3253,N_3021,N_3056);
or U3254 (N_3254,N_3085,N_3137);
xnor U3255 (N_3255,N_3115,N_3142);
xnor U3256 (N_3256,N_3009,N_3143);
nand U3257 (N_3257,N_3135,N_3068);
or U3258 (N_3258,N_3146,N_3180);
nor U3259 (N_3259,N_3071,N_3197);
or U3260 (N_3260,N_3006,N_3003);
or U3261 (N_3261,N_3060,N_3116);
xor U3262 (N_3262,N_3195,N_3131);
xor U3263 (N_3263,N_3083,N_3089);
nor U3264 (N_3264,N_3032,N_3165);
nand U3265 (N_3265,N_3106,N_3173);
nand U3266 (N_3266,N_3051,N_3134);
xor U3267 (N_3267,N_3091,N_3095);
xor U3268 (N_3268,N_3027,N_3086);
xnor U3269 (N_3269,N_3108,N_3040);
and U3270 (N_3270,N_3163,N_3196);
and U3271 (N_3271,N_3057,N_3148);
xor U3272 (N_3272,N_3178,N_3185);
nand U3273 (N_3273,N_3099,N_3061);
nor U3274 (N_3274,N_3198,N_3166);
xor U3275 (N_3275,N_3129,N_3169);
nand U3276 (N_3276,N_3102,N_3082);
nand U3277 (N_3277,N_3073,N_3069);
xnor U3278 (N_3278,N_3138,N_3188);
or U3279 (N_3279,N_3174,N_3097);
and U3280 (N_3280,N_3139,N_3087);
nor U3281 (N_3281,N_3147,N_3080);
and U3282 (N_3282,N_3183,N_3019);
nor U3283 (N_3283,N_3104,N_3168);
xor U3284 (N_3284,N_3182,N_3046);
and U3285 (N_3285,N_3199,N_3037);
nor U3286 (N_3286,N_3001,N_3153);
nor U3287 (N_3287,N_3159,N_3117);
nor U3288 (N_3288,N_3016,N_3075);
nand U3289 (N_3289,N_3065,N_3004);
and U3290 (N_3290,N_3132,N_3133);
nor U3291 (N_3291,N_3031,N_3111);
or U3292 (N_3292,N_3077,N_3107);
and U3293 (N_3293,N_3034,N_3035);
nand U3294 (N_3294,N_3076,N_3187);
xnor U3295 (N_3295,N_3092,N_3128);
nor U3296 (N_3296,N_3011,N_3072);
nand U3297 (N_3297,N_3118,N_3145);
and U3298 (N_3298,N_3176,N_3018);
or U3299 (N_3299,N_3157,N_3070);
or U3300 (N_3300,N_3029,N_3122);
nor U3301 (N_3301,N_3075,N_3005);
and U3302 (N_3302,N_3020,N_3088);
and U3303 (N_3303,N_3119,N_3091);
or U3304 (N_3304,N_3047,N_3057);
nand U3305 (N_3305,N_3049,N_3199);
xnor U3306 (N_3306,N_3193,N_3148);
xnor U3307 (N_3307,N_3110,N_3033);
or U3308 (N_3308,N_3150,N_3180);
xor U3309 (N_3309,N_3198,N_3148);
nand U3310 (N_3310,N_3163,N_3128);
nand U3311 (N_3311,N_3180,N_3073);
nor U3312 (N_3312,N_3019,N_3161);
or U3313 (N_3313,N_3188,N_3004);
nor U3314 (N_3314,N_3069,N_3055);
nor U3315 (N_3315,N_3076,N_3138);
xnor U3316 (N_3316,N_3058,N_3078);
nor U3317 (N_3317,N_3007,N_3100);
and U3318 (N_3318,N_3188,N_3104);
xnor U3319 (N_3319,N_3094,N_3008);
xnor U3320 (N_3320,N_3060,N_3163);
nor U3321 (N_3321,N_3142,N_3110);
xnor U3322 (N_3322,N_3132,N_3058);
nor U3323 (N_3323,N_3195,N_3094);
nor U3324 (N_3324,N_3137,N_3111);
nor U3325 (N_3325,N_3124,N_3049);
nor U3326 (N_3326,N_3155,N_3094);
nor U3327 (N_3327,N_3055,N_3133);
or U3328 (N_3328,N_3093,N_3035);
and U3329 (N_3329,N_3026,N_3036);
and U3330 (N_3330,N_3083,N_3064);
or U3331 (N_3331,N_3134,N_3050);
xnor U3332 (N_3332,N_3073,N_3015);
or U3333 (N_3333,N_3078,N_3112);
nand U3334 (N_3334,N_3045,N_3075);
or U3335 (N_3335,N_3094,N_3078);
nand U3336 (N_3336,N_3034,N_3170);
nand U3337 (N_3337,N_3169,N_3003);
nand U3338 (N_3338,N_3062,N_3067);
nor U3339 (N_3339,N_3075,N_3040);
or U3340 (N_3340,N_3041,N_3180);
nand U3341 (N_3341,N_3118,N_3061);
or U3342 (N_3342,N_3022,N_3045);
and U3343 (N_3343,N_3065,N_3106);
nor U3344 (N_3344,N_3180,N_3108);
and U3345 (N_3345,N_3166,N_3084);
xnor U3346 (N_3346,N_3116,N_3080);
or U3347 (N_3347,N_3147,N_3101);
or U3348 (N_3348,N_3055,N_3089);
and U3349 (N_3349,N_3102,N_3081);
xor U3350 (N_3350,N_3094,N_3009);
or U3351 (N_3351,N_3024,N_3065);
and U3352 (N_3352,N_3175,N_3123);
and U3353 (N_3353,N_3178,N_3164);
nand U3354 (N_3354,N_3111,N_3015);
xor U3355 (N_3355,N_3011,N_3027);
or U3356 (N_3356,N_3059,N_3071);
or U3357 (N_3357,N_3153,N_3004);
nand U3358 (N_3358,N_3041,N_3003);
xor U3359 (N_3359,N_3132,N_3086);
nand U3360 (N_3360,N_3168,N_3130);
xnor U3361 (N_3361,N_3001,N_3026);
and U3362 (N_3362,N_3159,N_3017);
and U3363 (N_3363,N_3187,N_3020);
or U3364 (N_3364,N_3009,N_3131);
nand U3365 (N_3365,N_3173,N_3009);
or U3366 (N_3366,N_3045,N_3068);
or U3367 (N_3367,N_3017,N_3131);
or U3368 (N_3368,N_3062,N_3048);
and U3369 (N_3369,N_3080,N_3032);
and U3370 (N_3370,N_3106,N_3092);
nor U3371 (N_3371,N_3167,N_3016);
xor U3372 (N_3372,N_3154,N_3180);
xnor U3373 (N_3373,N_3088,N_3148);
nor U3374 (N_3374,N_3097,N_3127);
xnor U3375 (N_3375,N_3055,N_3098);
or U3376 (N_3376,N_3140,N_3105);
or U3377 (N_3377,N_3137,N_3115);
nand U3378 (N_3378,N_3101,N_3102);
and U3379 (N_3379,N_3040,N_3076);
xor U3380 (N_3380,N_3195,N_3190);
xor U3381 (N_3381,N_3000,N_3171);
xor U3382 (N_3382,N_3127,N_3079);
and U3383 (N_3383,N_3083,N_3106);
nand U3384 (N_3384,N_3156,N_3179);
and U3385 (N_3385,N_3190,N_3097);
and U3386 (N_3386,N_3031,N_3148);
and U3387 (N_3387,N_3070,N_3169);
xor U3388 (N_3388,N_3034,N_3114);
and U3389 (N_3389,N_3190,N_3038);
and U3390 (N_3390,N_3068,N_3024);
nor U3391 (N_3391,N_3176,N_3113);
nand U3392 (N_3392,N_3020,N_3060);
nand U3393 (N_3393,N_3080,N_3057);
or U3394 (N_3394,N_3028,N_3183);
nor U3395 (N_3395,N_3111,N_3037);
nand U3396 (N_3396,N_3033,N_3170);
nand U3397 (N_3397,N_3076,N_3060);
nor U3398 (N_3398,N_3155,N_3181);
or U3399 (N_3399,N_3092,N_3107);
nor U3400 (N_3400,N_3336,N_3208);
xnor U3401 (N_3401,N_3323,N_3234);
and U3402 (N_3402,N_3247,N_3345);
or U3403 (N_3403,N_3305,N_3287);
and U3404 (N_3404,N_3245,N_3335);
xor U3405 (N_3405,N_3375,N_3388);
and U3406 (N_3406,N_3332,N_3258);
nand U3407 (N_3407,N_3390,N_3356);
nand U3408 (N_3408,N_3257,N_3278);
xor U3409 (N_3409,N_3200,N_3296);
and U3410 (N_3410,N_3286,N_3374);
or U3411 (N_3411,N_3297,N_3294);
or U3412 (N_3412,N_3307,N_3264);
xnor U3413 (N_3413,N_3276,N_3254);
nand U3414 (N_3414,N_3367,N_3275);
xor U3415 (N_3415,N_3211,N_3221);
and U3416 (N_3416,N_3277,N_3365);
and U3417 (N_3417,N_3225,N_3273);
or U3418 (N_3418,N_3291,N_3338);
or U3419 (N_3419,N_3330,N_3314);
and U3420 (N_3420,N_3353,N_3212);
or U3421 (N_3421,N_3238,N_3327);
or U3422 (N_3422,N_3393,N_3331);
nand U3423 (N_3423,N_3267,N_3298);
and U3424 (N_3424,N_3230,N_3381);
or U3425 (N_3425,N_3363,N_3265);
or U3426 (N_3426,N_3289,N_3309);
nor U3427 (N_3427,N_3359,N_3360);
xor U3428 (N_3428,N_3308,N_3269);
nand U3429 (N_3429,N_3285,N_3246);
nor U3430 (N_3430,N_3223,N_3394);
xnor U3431 (N_3431,N_3358,N_3292);
xor U3432 (N_3432,N_3318,N_3213);
nand U3433 (N_3433,N_3239,N_3214);
xnor U3434 (N_3434,N_3397,N_3255);
nor U3435 (N_3435,N_3312,N_3355);
nand U3436 (N_3436,N_3343,N_3272);
nor U3437 (N_3437,N_3281,N_3399);
and U3438 (N_3438,N_3271,N_3299);
xor U3439 (N_3439,N_3340,N_3380);
nor U3440 (N_3440,N_3203,N_3266);
nor U3441 (N_3441,N_3389,N_3372);
or U3442 (N_3442,N_3382,N_3224);
and U3443 (N_3443,N_3316,N_3209);
nor U3444 (N_3444,N_3352,N_3373);
xor U3445 (N_3445,N_3231,N_3354);
or U3446 (N_3446,N_3325,N_3282);
xnor U3447 (N_3447,N_3369,N_3398);
nand U3448 (N_3448,N_3201,N_3319);
nor U3449 (N_3449,N_3216,N_3283);
or U3450 (N_3450,N_3205,N_3290);
or U3451 (N_3451,N_3301,N_3253);
or U3452 (N_3452,N_3302,N_3341);
or U3453 (N_3453,N_3321,N_3279);
xor U3454 (N_3454,N_3317,N_3322);
xnor U3455 (N_3455,N_3385,N_3241);
nor U3456 (N_3456,N_3344,N_3249);
nor U3457 (N_3457,N_3243,N_3364);
nor U3458 (N_3458,N_3348,N_3370);
nor U3459 (N_3459,N_3242,N_3260);
or U3460 (N_3460,N_3329,N_3326);
nand U3461 (N_3461,N_3217,N_3215);
or U3462 (N_3462,N_3248,N_3251);
and U3463 (N_3463,N_3220,N_3207);
and U3464 (N_3464,N_3280,N_3263);
xnor U3465 (N_3465,N_3218,N_3284);
nor U3466 (N_3466,N_3386,N_3244);
or U3467 (N_3467,N_3304,N_3293);
xor U3468 (N_3468,N_3379,N_3270);
or U3469 (N_3469,N_3378,N_3262);
nand U3470 (N_3470,N_3303,N_3311);
and U3471 (N_3471,N_3222,N_3250);
nor U3472 (N_3472,N_3371,N_3315);
xor U3473 (N_3473,N_3261,N_3202);
and U3474 (N_3474,N_3320,N_3339);
xnor U3475 (N_3475,N_3235,N_3350);
xor U3476 (N_3476,N_3368,N_3342);
nand U3477 (N_3477,N_3383,N_3384);
nand U3478 (N_3478,N_3337,N_3300);
or U3479 (N_3479,N_3233,N_3206);
nand U3480 (N_3480,N_3347,N_3232);
xor U3481 (N_3481,N_3256,N_3236);
nand U3482 (N_3482,N_3391,N_3295);
nand U3483 (N_3483,N_3306,N_3366);
xnor U3484 (N_3484,N_3228,N_3210);
nor U3485 (N_3485,N_3334,N_3376);
xor U3486 (N_3486,N_3328,N_3313);
or U3487 (N_3487,N_3357,N_3268);
or U3488 (N_3488,N_3252,N_3349);
xor U3489 (N_3489,N_3288,N_3229);
nor U3490 (N_3490,N_3392,N_3274);
xnor U3491 (N_3491,N_3310,N_3361);
or U3492 (N_3492,N_3226,N_3333);
and U3493 (N_3493,N_3219,N_3395);
or U3494 (N_3494,N_3351,N_3237);
xnor U3495 (N_3495,N_3362,N_3259);
nand U3496 (N_3496,N_3387,N_3346);
nand U3497 (N_3497,N_3204,N_3377);
and U3498 (N_3498,N_3396,N_3227);
xor U3499 (N_3499,N_3324,N_3240);
or U3500 (N_3500,N_3248,N_3202);
nand U3501 (N_3501,N_3280,N_3322);
nand U3502 (N_3502,N_3227,N_3266);
and U3503 (N_3503,N_3360,N_3260);
or U3504 (N_3504,N_3302,N_3231);
xor U3505 (N_3505,N_3259,N_3246);
or U3506 (N_3506,N_3313,N_3202);
or U3507 (N_3507,N_3321,N_3289);
nor U3508 (N_3508,N_3236,N_3390);
nand U3509 (N_3509,N_3314,N_3365);
xor U3510 (N_3510,N_3340,N_3293);
or U3511 (N_3511,N_3203,N_3282);
and U3512 (N_3512,N_3351,N_3319);
nand U3513 (N_3513,N_3270,N_3392);
nand U3514 (N_3514,N_3398,N_3302);
nor U3515 (N_3515,N_3257,N_3253);
nand U3516 (N_3516,N_3323,N_3363);
xnor U3517 (N_3517,N_3346,N_3321);
nand U3518 (N_3518,N_3304,N_3398);
and U3519 (N_3519,N_3227,N_3365);
and U3520 (N_3520,N_3381,N_3207);
and U3521 (N_3521,N_3279,N_3275);
xnor U3522 (N_3522,N_3318,N_3217);
xor U3523 (N_3523,N_3359,N_3295);
xor U3524 (N_3524,N_3390,N_3357);
and U3525 (N_3525,N_3251,N_3393);
xnor U3526 (N_3526,N_3321,N_3219);
xor U3527 (N_3527,N_3261,N_3200);
nand U3528 (N_3528,N_3336,N_3232);
or U3529 (N_3529,N_3274,N_3356);
nand U3530 (N_3530,N_3364,N_3241);
nor U3531 (N_3531,N_3230,N_3376);
or U3532 (N_3532,N_3305,N_3216);
nor U3533 (N_3533,N_3226,N_3286);
xor U3534 (N_3534,N_3278,N_3255);
nor U3535 (N_3535,N_3386,N_3259);
nor U3536 (N_3536,N_3222,N_3242);
nand U3537 (N_3537,N_3323,N_3307);
or U3538 (N_3538,N_3296,N_3279);
xor U3539 (N_3539,N_3387,N_3269);
xor U3540 (N_3540,N_3383,N_3289);
xor U3541 (N_3541,N_3279,N_3329);
nand U3542 (N_3542,N_3222,N_3213);
nand U3543 (N_3543,N_3256,N_3277);
nand U3544 (N_3544,N_3388,N_3315);
and U3545 (N_3545,N_3348,N_3336);
or U3546 (N_3546,N_3341,N_3233);
nor U3547 (N_3547,N_3383,N_3296);
nor U3548 (N_3548,N_3396,N_3224);
nor U3549 (N_3549,N_3294,N_3212);
and U3550 (N_3550,N_3254,N_3258);
and U3551 (N_3551,N_3330,N_3321);
nand U3552 (N_3552,N_3278,N_3248);
or U3553 (N_3553,N_3383,N_3369);
nand U3554 (N_3554,N_3376,N_3273);
nand U3555 (N_3555,N_3387,N_3329);
and U3556 (N_3556,N_3379,N_3393);
or U3557 (N_3557,N_3386,N_3223);
nor U3558 (N_3558,N_3333,N_3373);
xnor U3559 (N_3559,N_3393,N_3285);
xor U3560 (N_3560,N_3259,N_3387);
xnor U3561 (N_3561,N_3229,N_3205);
or U3562 (N_3562,N_3307,N_3309);
or U3563 (N_3563,N_3235,N_3278);
nand U3564 (N_3564,N_3366,N_3218);
xnor U3565 (N_3565,N_3347,N_3393);
nor U3566 (N_3566,N_3242,N_3356);
and U3567 (N_3567,N_3255,N_3318);
and U3568 (N_3568,N_3249,N_3291);
nor U3569 (N_3569,N_3370,N_3241);
nor U3570 (N_3570,N_3370,N_3279);
xor U3571 (N_3571,N_3213,N_3210);
and U3572 (N_3572,N_3369,N_3308);
nor U3573 (N_3573,N_3300,N_3282);
xnor U3574 (N_3574,N_3312,N_3238);
or U3575 (N_3575,N_3305,N_3265);
or U3576 (N_3576,N_3314,N_3236);
xnor U3577 (N_3577,N_3389,N_3305);
or U3578 (N_3578,N_3279,N_3262);
or U3579 (N_3579,N_3221,N_3290);
or U3580 (N_3580,N_3327,N_3368);
nor U3581 (N_3581,N_3342,N_3206);
or U3582 (N_3582,N_3384,N_3316);
or U3583 (N_3583,N_3228,N_3324);
nor U3584 (N_3584,N_3336,N_3341);
xor U3585 (N_3585,N_3225,N_3247);
nand U3586 (N_3586,N_3206,N_3387);
nor U3587 (N_3587,N_3394,N_3338);
nand U3588 (N_3588,N_3332,N_3306);
nor U3589 (N_3589,N_3299,N_3282);
nand U3590 (N_3590,N_3320,N_3244);
nand U3591 (N_3591,N_3225,N_3244);
xor U3592 (N_3592,N_3266,N_3307);
or U3593 (N_3593,N_3237,N_3211);
nor U3594 (N_3594,N_3271,N_3215);
or U3595 (N_3595,N_3372,N_3270);
or U3596 (N_3596,N_3315,N_3297);
and U3597 (N_3597,N_3267,N_3225);
nor U3598 (N_3598,N_3278,N_3243);
nand U3599 (N_3599,N_3298,N_3259);
or U3600 (N_3600,N_3529,N_3501);
xnor U3601 (N_3601,N_3585,N_3486);
xor U3602 (N_3602,N_3411,N_3586);
xnor U3603 (N_3603,N_3400,N_3565);
and U3604 (N_3604,N_3554,N_3582);
and U3605 (N_3605,N_3598,N_3461);
xnor U3606 (N_3606,N_3511,N_3551);
nor U3607 (N_3607,N_3405,N_3469);
xor U3608 (N_3608,N_3449,N_3481);
nor U3609 (N_3609,N_3430,N_3516);
and U3610 (N_3610,N_3443,N_3476);
and U3611 (N_3611,N_3555,N_3504);
and U3612 (N_3612,N_3572,N_3523);
or U3613 (N_3613,N_3425,N_3442);
xor U3614 (N_3614,N_3513,N_3571);
and U3615 (N_3615,N_3521,N_3455);
and U3616 (N_3616,N_3459,N_3491);
xnor U3617 (N_3617,N_3496,N_3512);
nor U3618 (N_3618,N_3557,N_3418);
xor U3619 (N_3619,N_3517,N_3440);
nand U3620 (N_3620,N_3537,N_3489);
or U3621 (N_3621,N_3505,N_3460);
xor U3622 (N_3622,N_3577,N_3478);
nand U3623 (N_3623,N_3527,N_3497);
nand U3624 (N_3624,N_3434,N_3483);
and U3625 (N_3625,N_3433,N_3453);
xor U3626 (N_3626,N_3406,N_3592);
or U3627 (N_3627,N_3539,N_3414);
nand U3628 (N_3628,N_3589,N_3508);
or U3629 (N_3629,N_3468,N_3561);
nand U3630 (N_3630,N_3412,N_3550);
xnor U3631 (N_3631,N_3543,N_3439);
nand U3632 (N_3632,N_3428,N_3456);
nor U3633 (N_3633,N_3526,N_3426);
nand U3634 (N_3634,N_3482,N_3503);
xnor U3635 (N_3635,N_3590,N_3553);
and U3636 (N_3636,N_3588,N_3444);
xor U3637 (N_3637,N_3474,N_3534);
or U3638 (N_3638,N_3532,N_3424);
or U3639 (N_3639,N_3432,N_3558);
xnor U3640 (N_3640,N_3587,N_3579);
nand U3641 (N_3641,N_3542,N_3573);
nand U3642 (N_3642,N_3450,N_3436);
nor U3643 (N_3643,N_3580,N_3420);
nor U3644 (N_3644,N_3519,N_3536);
or U3645 (N_3645,N_3502,N_3591);
nand U3646 (N_3646,N_3528,N_3574);
or U3647 (N_3647,N_3566,N_3413);
nand U3648 (N_3648,N_3494,N_3416);
or U3649 (N_3649,N_3463,N_3510);
and U3650 (N_3650,N_3467,N_3531);
nor U3651 (N_3651,N_3583,N_3417);
nand U3652 (N_3652,N_3475,N_3593);
nand U3653 (N_3653,N_3547,N_3599);
nor U3654 (N_3654,N_3484,N_3451);
and U3655 (N_3655,N_3530,N_3562);
and U3656 (N_3656,N_3429,N_3470);
or U3657 (N_3657,N_3454,N_3437);
nor U3658 (N_3658,N_3471,N_3404);
xnor U3659 (N_3659,N_3560,N_3490);
or U3660 (N_3660,N_3544,N_3488);
and U3661 (N_3661,N_3500,N_3438);
and U3662 (N_3662,N_3457,N_3446);
xor U3663 (N_3663,N_3584,N_3518);
nor U3664 (N_3664,N_3552,N_3545);
nor U3665 (N_3665,N_3465,N_3458);
nor U3666 (N_3666,N_3415,N_3431);
and U3667 (N_3667,N_3515,N_3403);
nand U3668 (N_3668,N_3448,N_3548);
or U3669 (N_3669,N_3533,N_3506);
nor U3670 (N_3670,N_3423,N_3472);
xor U3671 (N_3671,N_3578,N_3538);
and U3672 (N_3672,N_3597,N_3575);
nand U3673 (N_3673,N_3568,N_3441);
xor U3674 (N_3674,N_3556,N_3408);
or U3675 (N_3675,N_3410,N_3581);
nor U3676 (N_3676,N_3464,N_3522);
nand U3677 (N_3677,N_3487,N_3564);
nor U3678 (N_3678,N_3419,N_3447);
xnor U3679 (N_3679,N_3479,N_3514);
xor U3680 (N_3680,N_3401,N_3594);
xnor U3681 (N_3681,N_3549,N_3492);
nand U3682 (N_3682,N_3546,N_3495);
nand U3683 (N_3683,N_3485,N_3520);
nor U3684 (N_3684,N_3407,N_3427);
xor U3685 (N_3685,N_3570,N_3493);
xor U3686 (N_3686,N_3445,N_3473);
and U3687 (N_3687,N_3525,N_3409);
or U3688 (N_3688,N_3480,N_3535);
nand U3689 (N_3689,N_3477,N_3595);
or U3690 (N_3690,N_3422,N_3498);
xor U3691 (N_3691,N_3421,N_3402);
or U3692 (N_3692,N_3559,N_3541);
and U3693 (N_3693,N_3569,N_3596);
xor U3694 (N_3694,N_3524,N_3452);
nor U3695 (N_3695,N_3576,N_3567);
or U3696 (N_3696,N_3462,N_3499);
xnor U3697 (N_3697,N_3507,N_3509);
xnor U3698 (N_3698,N_3540,N_3435);
xnor U3699 (N_3699,N_3466,N_3563);
or U3700 (N_3700,N_3423,N_3490);
or U3701 (N_3701,N_3427,N_3594);
xnor U3702 (N_3702,N_3434,N_3421);
nand U3703 (N_3703,N_3422,N_3567);
nand U3704 (N_3704,N_3405,N_3535);
or U3705 (N_3705,N_3511,N_3554);
and U3706 (N_3706,N_3461,N_3436);
and U3707 (N_3707,N_3459,N_3567);
nor U3708 (N_3708,N_3544,N_3481);
or U3709 (N_3709,N_3488,N_3499);
or U3710 (N_3710,N_3586,N_3550);
nor U3711 (N_3711,N_3502,N_3442);
nand U3712 (N_3712,N_3532,N_3455);
nand U3713 (N_3713,N_3455,N_3433);
nand U3714 (N_3714,N_3478,N_3436);
nor U3715 (N_3715,N_3579,N_3563);
xor U3716 (N_3716,N_3489,N_3596);
and U3717 (N_3717,N_3408,N_3486);
xor U3718 (N_3718,N_3456,N_3544);
nor U3719 (N_3719,N_3456,N_3401);
nor U3720 (N_3720,N_3439,N_3550);
xnor U3721 (N_3721,N_3590,N_3495);
nand U3722 (N_3722,N_3509,N_3534);
nor U3723 (N_3723,N_3579,N_3582);
and U3724 (N_3724,N_3523,N_3500);
xor U3725 (N_3725,N_3472,N_3451);
or U3726 (N_3726,N_3552,N_3465);
or U3727 (N_3727,N_3580,N_3402);
nor U3728 (N_3728,N_3561,N_3421);
or U3729 (N_3729,N_3591,N_3535);
nor U3730 (N_3730,N_3545,N_3578);
or U3731 (N_3731,N_3560,N_3479);
xnor U3732 (N_3732,N_3517,N_3438);
nand U3733 (N_3733,N_3401,N_3505);
nand U3734 (N_3734,N_3443,N_3575);
nor U3735 (N_3735,N_3546,N_3564);
xor U3736 (N_3736,N_3406,N_3458);
nor U3737 (N_3737,N_3415,N_3434);
xnor U3738 (N_3738,N_3424,N_3521);
nor U3739 (N_3739,N_3459,N_3582);
and U3740 (N_3740,N_3416,N_3471);
xor U3741 (N_3741,N_3406,N_3553);
nand U3742 (N_3742,N_3577,N_3503);
and U3743 (N_3743,N_3420,N_3561);
and U3744 (N_3744,N_3575,N_3586);
and U3745 (N_3745,N_3484,N_3438);
or U3746 (N_3746,N_3434,N_3468);
or U3747 (N_3747,N_3493,N_3448);
nor U3748 (N_3748,N_3490,N_3506);
nand U3749 (N_3749,N_3558,N_3409);
xnor U3750 (N_3750,N_3473,N_3459);
nand U3751 (N_3751,N_3513,N_3449);
or U3752 (N_3752,N_3430,N_3459);
nor U3753 (N_3753,N_3589,N_3514);
nand U3754 (N_3754,N_3415,N_3549);
nor U3755 (N_3755,N_3570,N_3500);
and U3756 (N_3756,N_3537,N_3544);
nand U3757 (N_3757,N_3480,N_3509);
nand U3758 (N_3758,N_3495,N_3593);
and U3759 (N_3759,N_3454,N_3577);
xor U3760 (N_3760,N_3556,N_3502);
nand U3761 (N_3761,N_3589,N_3495);
xnor U3762 (N_3762,N_3434,N_3593);
and U3763 (N_3763,N_3524,N_3545);
nand U3764 (N_3764,N_3591,N_3417);
nand U3765 (N_3765,N_3482,N_3517);
xor U3766 (N_3766,N_3528,N_3558);
xnor U3767 (N_3767,N_3552,N_3442);
nand U3768 (N_3768,N_3536,N_3544);
nand U3769 (N_3769,N_3526,N_3468);
xnor U3770 (N_3770,N_3527,N_3441);
nand U3771 (N_3771,N_3584,N_3429);
or U3772 (N_3772,N_3495,N_3540);
or U3773 (N_3773,N_3405,N_3476);
nand U3774 (N_3774,N_3501,N_3438);
nand U3775 (N_3775,N_3495,N_3531);
or U3776 (N_3776,N_3508,N_3457);
nor U3777 (N_3777,N_3426,N_3414);
nand U3778 (N_3778,N_3534,N_3560);
and U3779 (N_3779,N_3585,N_3456);
xnor U3780 (N_3780,N_3510,N_3583);
nand U3781 (N_3781,N_3527,N_3509);
or U3782 (N_3782,N_3561,N_3511);
nand U3783 (N_3783,N_3476,N_3560);
or U3784 (N_3784,N_3438,N_3572);
xnor U3785 (N_3785,N_3458,N_3444);
nand U3786 (N_3786,N_3490,N_3513);
or U3787 (N_3787,N_3537,N_3404);
nor U3788 (N_3788,N_3410,N_3407);
nand U3789 (N_3789,N_3446,N_3520);
nand U3790 (N_3790,N_3459,N_3523);
nand U3791 (N_3791,N_3457,N_3527);
nor U3792 (N_3792,N_3440,N_3553);
nand U3793 (N_3793,N_3480,N_3573);
nand U3794 (N_3794,N_3498,N_3472);
xnor U3795 (N_3795,N_3536,N_3405);
or U3796 (N_3796,N_3434,N_3479);
and U3797 (N_3797,N_3529,N_3531);
and U3798 (N_3798,N_3462,N_3559);
nand U3799 (N_3799,N_3480,N_3502);
nand U3800 (N_3800,N_3636,N_3711);
nor U3801 (N_3801,N_3671,N_3610);
and U3802 (N_3802,N_3720,N_3784);
and U3803 (N_3803,N_3786,N_3764);
and U3804 (N_3804,N_3656,N_3747);
and U3805 (N_3805,N_3777,N_3664);
or U3806 (N_3806,N_3738,N_3614);
nor U3807 (N_3807,N_3702,N_3616);
nand U3808 (N_3808,N_3739,N_3727);
nand U3809 (N_3809,N_3686,N_3635);
nand U3810 (N_3810,N_3743,N_3698);
and U3811 (N_3811,N_3795,N_3700);
xnor U3812 (N_3812,N_3628,N_3678);
xor U3813 (N_3813,N_3737,N_3696);
xor U3814 (N_3814,N_3687,N_3751);
and U3815 (N_3815,N_3620,N_3679);
and U3816 (N_3816,N_3745,N_3680);
xor U3817 (N_3817,N_3746,N_3668);
and U3818 (N_3818,N_3607,N_3730);
or U3819 (N_3819,N_3728,N_3638);
xnor U3820 (N_3820,N_3783,N_3761);
nor U3821 (N_3821,N_3781,N_3753);
and U3822 (N_3822,N_3689,N_3622);
or U3823 (N_3823,N_3791,N_3758);
nand U3824 (N_3824,N_3787,N_3632);
xnor U3825 (N_3825,N_3693,N_3677);
nand U3826 (N_3826,N_3667,N_3619);
and U3827 (N_3827,N_3782,N_3708);
xnor U3828 (N_3828,N_3659,N_3719);
xor U3829 (N_3829,N_3756,N_3731);
and U3830 (N_3830,N_3754,N_3609);
nand U3831 (N_3831,N_3769,N_3654);
nor U3832 (N_3832,N_3774,N_3740);
nand U3833 (N_3833,N_3767,N_3716);
and U3834 (N_3834,N_3666,N_3613);
xor U3835 (N_3835,N_3732,N_3631);
and U3836 (N_3836,N_3721,N_3658);
xnor U3837 (N_3837,N_3776,N_3752);
nor U3838 (N_3838,N_3771,N_3624);
nor U3839 (N_3839,N_3629,N_3697);
xnor U3840 (N_3840,N_3744,N_3797);
or U3841 (N_3841,N_3798,N_3643);
nand U3842 (N_3842,N_3652,N_3703);
nor U3843 (N_3843,N_3644,N_3625);
xnor U3844 (N_3844,N_3646,N_3692);
and U3845 (N_3845,N_3605,N_3749);
and U3846 (N_3846,N_3729,N_3755);
or U3847 (N_3847,N_3639,N_3640);
nand U3848 (N_3848,N_3688,N_3672);
nand U3849 (N_3849,N_3669,N_3760);
and U3850 (N_3850,N_3675,N_3765);
nand U3851 (N_3851,N_3701,N_3681);
nand U3852 (N_3852,N_3655,N_3673);
xor U3853 (N_3853,N_3723,N_3726);
or U3854 (N_3854,N_3617,N_3789);
xor U3855 (N_3855,N_3651,N_3772);
nor U3856 (N_3856,N_3603,N_3691);
or U3857 (N_3857,N_3601,N_3653);
nand U3858 (N_3858,N_3750,N_3630);
nor U3859 (N_3859,N_3790,N_3799);
nor U3860 (N_3860,N_3796,N_3741);
and U3861 (N_3861,N_3633,N_3634);
and U3862 (N_3862,N_3676,N_3706);
and U3863 (N_3863,N_3733,N_3611);
xnor U3864 (N_3864,N_3661,N_3712);
xnor U3865 (N_3865,N_3621,N_3649);
nor U3866 (N_3866,N_3718,N_3788);
nor U3867 (N_3867,N_3742,N_3725);
and U3868 (N_3868,N_3773,N_3785);
nor U3869 (N_3869,N_3627,N_3674);
or U3870 (N_3870,N_3606,N_3780);
and U3871 (N_3871,N_3734,N_3647);
nor U3872 (N_3872,N_3735,N_3717);
or U3873 (N_3873,N_3748,N_3618);
and U3874 (N_3874,N_3615,N_3608);
and U3875 (N_3875,N_3637,N_3736);
and U3876 (N_3876,N_3690,N_3670);
xor U3877 (N_3877,N_3763,N_3657);
xnor U3878 (N_3878,N_3695,N_3683);
or U3879 (N_3879,N_3768,N_3770);
or U3880 (N_3880,N_3641,N_3626);
nand U3881 (N_3881,N_3648,N_3705);
or U3882 (N_3882,N_3707,N_3757);
or U3883 (N_3883,N_3694,N_3665);
nand U3884 (N_3884,N_3604,N_3759);
xnor U3885 (N_3885,N_3775,N_3722);
or U3886 (N_3886,N_3662,N_3663);
nor U3887 (N_3887,N_3684,N_3623);
xor U3888 (N_3888,N_3779,N_3778);
and U3889 (N_3889,N_3600,N_3762);
nor U3890 (N_3890,N_3766,N_3642);
xnor U3891 (N_3891,N_3650,N_3602);
nor U3892 (N_3892,N_3682,N_3612);
xnor U3893 (N_3893,N_3645,N_3710);
and U3894 (N_3894,N_3713,N_3699);
nand U3895 (N_3895,N_3660,N_3709);
or U3896 (N_3896,N_3793,N_3704);
or U3897 (N_3897,N_3724,N_3714);
xnor U3898 (N_3898,N_3685,N_3792);
or U3899 (N_3899,N_3715,N_3794);
xnor U3900 (N_3900,N_3711,N_3666);
nor U3901 (N_3901,N_3636,N_3690);
or U3902 (N_3902,N_3667,N_3782);
nor U3903 (N_3903,N_3783,N_3649);
xor U3904 (N_3904,N_3676,N_3705);
nor U3905 (N_3905,N_3623,N_3656);
or U3906 (N_3906,N_3713,N_3789);
nor U3907 (N_3907,N_3737,N_3613);
nor U3908 (N_3908,N_3739,N_3696);
nor U3909 (N_3909,N_3674,N_3665);
nor U3910 (N_3910,N_3667,N_3662);
or U3911 (N_3911,N_3730,N_3602);
xor U3912 (N_3912,N_3743,N_3609);
and U3913 (N_3913,N_3780,N_3714);
xnor U3914 (N_3914,N_3759,N_3771);
nand U3915 (N_3915,N_3762,N_3648);
and U3916 (N_3916,N_3732,N_3678);
or U3917 (N_3917,N_3711,N_3685);
or U3918 (N_3918,N_3620,N_3762);
or U3919 (N_3919,N_3656,N_3649);
nor U3920 (N_3920,N_3663,N_3758);
nor U3921 (N_3921,N_3768,N_3653);
nor U3922 (N_3922,N_3743,N_3751);
and U3923 (N_3923,N_3729,N_3739);
nand U3924 (N_3924,N_3760,N_3737);
or U3925 (N_3925,N_3769,N_3618);
xor U3926 (N_3926,N_3682,N_3676);
nand U3927 (N_3927,N_3793,N_3715);
xnor U3928 (N_3928,N_3728,N_3699);
or U3929 (N_3929,N_3745,N_3721);
nand U3930 (N_3930,N_3727,N_3661);
and U3931 (N_3931,N_3666,N_3639);
and U3932 (N_3932,N_3691,N_3630);
and U3933 (N_3933,N_3750,N_3765);
and U3934 (N_3934,N_3785,N_3714);
nand U3935 (N_3935,N_3611,N_3681);
nand U3936 (N_3936,N_3760,N_3795);
xnor U3937 (N_3937,N_3788,N_3771);
xor U3938 (N_3938,N_3701,N_3650);
xnor U3939 (N_3939,N_3643,N_3695);
nor U3940 (N_3940,N_3767,N_3682);
nand U3941 (N_3941,N_3792,N_3733);
xnor U3942 (N_3942,N_3757,N_3652);
xor U3943 (N_3943,N_3761,N_3663);
or U3944 (N_3944,N_3614,N_3703);
nor U3945 (N_3945,N_3704,N_3763);
or U3946 (N_3946,N_3655,N_3748);
or U3947 (N_3947,N_3793,N_3780);
nand U3948 (N_3948,N_3711,N_3640);
and U3949 (N_3949,N_3688,N_3733);
or U3950 (N_3950,N_3663,N_3748);
xnor U3951 (N_3951,N_3767,N_3731);
nor U3952 (N_3952,N_3715,N_3655);
and U3953 (N_3953,N_3661,N_3794);
and U3954 (N_3954,N_3730,N_3702);
nor U3955 (N_3955,N_3730,N_3681);
nor U3956 (N_3956,N_3784,N_3649);
and U3957 (N_3957,N_3668,N_3734);
nand U3958 (N_3958,N_3671,N_3735);
or U3959 (N_3959,N_3641,N_3632);
and U3960 (N_3960,N_3613,N_3695);
and U3961 (N_3961,N_3719,N_3768);
or U3962 (N_3962,N_3675,N_3744);
or U3963 (N_3963,N_3776,N_3730);
and U3964 (N_3964,N_3717,N_3681);
nand U3965 (N_3965,N_3632,N_3781);
xnor U3966 (N_3966,N_3620,N_3751);
nor U3967 (N_3967,N_3717,N_3790);
and U3968 (N_3968,N_3601,N_3652);
nand U3969 (N_3969,N_3759,N_3690);
xnor U3970 (N_3970,N_3654,N_3697);
nor U3971 (N_3971,N_3735,N_3623);
nand U3972 (N_3972,N_3640,N_3685);
and U3973 (N_3973,N_3728,N_3636);
or U3974 (N_3974,N_3716,N_3649);
nor U3975 (N_3975,N_3611,N_3634);
nor U3976 (N_3976,N_3714,N_3626);
nand U3977 (N_3977,N_3782,N_3759);
xnor U3978 (N_3978,N_3650,N_3677);
xor U3979 (N_3979,N_3714,N_3645);
nand U3980 (N_3980,N_3712,N_3664);
nor U3981 (N_3981,N_3639,N_3759);
nor U3982 (N_3982,N_3745,N_3780);
and U3983 (N_3983,N_3784,N_3787);
xor U3984 (N_3984,N_3679,N_3600);
xnor U3985 (N_3985,N_3761,N_3774);
nor U3986 (N_3986,N_3797,N_3647);
or U3987 (N_3987,N_3771,N_3608);
or U3988 (N_3988,N_3636,N_3676);
or U3989 (N_3989,N_3630,N_3701);
and U3990 (N_3990,N_3611,N_3753);
and U3991 (N_3991,N_3671,N_3631);
and U3992 (N_3992,N_3710,N_3614);
nand U3993 (N_3993,N_3702,N_3698);
or U3994 (N_3994,N_3662,N_3741);
xor U3995 (N_3995,N_3760,N_3705);
and U3996 (N_3996,N_3721,N_3648);
nor U3997 (N_3997,N_3644,N_3748);
or U3998 (N_3998,N_3645,N_3778);
xor U3999 (N_3999,N_3667,N_3795);
and U4000 (N_4000,N_3945,N_3918);
or U4001 (N_4001,N_3812,N_3862);
xnor U4002 (N_4002,N_3907,N_3870);
and U4003 (N_4003,N_3974,N_3874);
and U4004 (N_4004,N_3970,N_3980);
and U4005 (N_4005,N_3882,N_3818);
and U4006 (N_4006,N_3892,N_3982);
xnor U4007 (N_4007,N_3959,N_3823);
xnor U4008 (N_4008,N_3849,N_3951);
and U4009 (N_4009,N_3966,N_3856);
nand U4010 (N_4010,N_3865,N_3926);
nand U4011 (N_4011,N_3869,N_3928);
and U4012 (N_4012,N_3954,N_3977);
xnor U4013 (N_4013,N_3805,N_3851);
xnor U4014 (N_4014,N_3871,N_3934);
xnor U4015 (N_4015,N_3930,N_3993);
and U4016 (N_4016,N_3842,N_3990);
and U4017 (N_4017,N_3912,N_3820);
xor U4018 (N_4018,N_3833,N_3913);
nand U4019 (N_4019,N_3873,N_3979);
and U4020 (N_4020,N_3888,N_3824);
or U4021 (N_4021,N_3855,N_3887);
and U4022 (N_4022,N_3973,N_3878);
xor U4023 (N_4023,N_3910,N_3829);
xor U4024 (N_4024,N_3802,N_3859);
nor U4025 (N_4025,N_3936,N_3801);
nor U4026 (N_4026,N_3999,N_3898);
xnor U4027 (N_4027,N_3969,N_3964);
xor U4028 (N_4028,N_3872,N_3958);
and U4029 (N_4029,N_3989,N_3809);
and U4030 (N_4030,N_3877,N_3944);
nand U4031 (N_4031,N_3831,N_3889);
nand U4032 (N_4032,N_3995,N_3950);
and U4033 (N_4033,N_3868,N_3853);
xnor U4034 (N_4034,N_3858,N_3976);
or U4035 (N_4035,N_3899,N_3937);
and U4036 (N_4036,N_3992,N_3939);
and U4037 (N_4037,N_3943,N_3813);
nor U4038 (N_4038,N_3965,N_3956);
nand U4039 (N_4039,N_3848,N_3963);
and U4040 (N_4040,N_3875,N_3920);
nor U4041 (N_4041,N_3808,N_3938);
nor U4042 (N_4042,N_3884,N_3852);
or U4043 (N_4043,N_3925,N_3984);
nor U4044 (N_4044,N_3861,N_3886);
xnor U4045 (N_4045,N_3857,N_3840);
and U4046 (N_4046,N_3916,N_3987);
xor U4047 (N_4047,N_3828,N_3998);
and U4048 (N_4048,N_3835,N_3978);
nand U4049 (N_4049,N_3983,N_3915);
nor U4050 (N_4050,N_3864,N_3827);
and U4051 (N_4051,N_3814,N_3923);
nor U4052 (N_4052,N_3948,N_3909);
nor U4053 (N_4053,N_3949,N_3906);
or U4054 (N_4054,N_3891,N_3815);
nand U4055 (N_4055,N_3847,N_3932);
nand U4056 (N_4056,N_3894,N_3843);
nor U4057 (N_4057,N_3924,N_3896);
and U4058 (N_4058,N_3839,N_3957);
and U4059 (N_4059,N_3991,N_3961);
nor U4060 (N_4060,N_3986,N_3806);
or U4061 (N_4061,N_3914,N_3940);
xnor U4062 (N_4062,N_3921,N_3952);
nor U4063 (N_4063,N_3935,N_3819);
or U4064 (N_4064,N_3854,N_3846);
nor U4065 (N_4065,N_3947,N_3962);
and U4066 (N_4066,N_3931,N_3900);
nand U4067 (N_4067,N_3845,N_3841);
xnor U4068 (N_4068,N_3879,N_3933);
and U4069 (N_4069,N_3942,N_3883);
nand U4070 (N_4070,N_3803,N_3972);
or U4071 (N_4071,N_3844,N_3804);
nor U4072 (N_4072,N_3971,N_3895);
nor U4073 (N_4073,N_3985,N_3941);
xor U4074 (N_4074,N_3880,N_3890);
or U4075 (N_4075,N_3968,N_3975);
nand U4076 (N_4076,N_3967,N_3822);
nor U4077 (N_4077,N_3994,N_3919);
or U4078 (N_4078,N_3903,N_3917);
nand U4079 (N_4079,N_3946,N_3902);
nand U4080 (N_4080,N_3893,N_3927);
xnor U4081 (N_4081,N_3834,N_3838);
xor U4082 (N_4082,N_3816,N_3897);
nand U4083 (N_4083,N_3810,N_3929);
nor U4084 (N_4084,N_3825,N_3953);
nor U4085 (N_4085,N_3876,N_3863);
nand U4086 (N_4086,N_3866,N_3826);
nor U4087 (N_4087,N_3821,N_3908);
nand U4088 (N_4088,N_3988,N_3860);
nand U4089 (N_4089,N_3885,N_3960);
nand U4090 (N_4090,N_3850,N_3832);
nand U4091 (N_4091,N_3811,N_3901);
or U4092 (N_4092,N_3867,N_3881);
or U4093 (N_4093,N_3905,N_3836);
xnor U4094 (N_4094,N_3830,N_3922);
xnor U4095 (N_4095,N_3911,N_3800);
xnor U4096 (N_4096,N_3996,N_3904);
or U4097 (N_4097,N_3997,N_3817);
xnor U4098 (N_4098,N_3955,N_3981);
and U4099 (N_4099,N_3837,N_3807);
or U4100 (N_4100,N_3944,N_3963);
nor U4101 (N_4101,N_3810,N_3960);
nor U4102 (N_4102,N_3837,N_3959);
xor U4103 (N_4103,N_3899,N_3998);
or U4104 (N_4104,N_3896,N_3972);
nor U4105 (N_4105,N_3947,N_3838);
and U4106 (N_4106,N_3910,N_3801);
and U4107 (N_4107,N_3900,N_3809);
nor U4108 (N_4108,N_3928,N_3874);
nor U4109 (N_4109,N_3981,N_3925);
and U4110 (N_4110,N_3860,N_3858);
nor U4111 (N_4111,N_3873,N_3828);
xor U4112 (N_4112,N_3908,N_3891);
nor U4113 (N_4113,N_3916,N_3947);
and U4114 (N_4114,N_3972,N_3883);
nand U4115 (N_4115,N_3910,N_3819);
or U4116 (N_4116,N_3812,N_3923);
and U4117 (N_4117,N_3826,N_3812);
nand U4118 (N_4118,N_3808,N_3809);
xor U4119 (N_4119,N_3948,N_3862);
xnor U4120 (N_4120,N_3953,N_3925);
and U4121 (N_4121,N_3986,N_3994);
or U4122 (N_4122,N_3894,N_3815);
xor U4123 (N_4123,N_3984,N_3835);
nand U4124 (N_4124,N_3978,N_3940);
nor U4125 (N_4125,N_3857,N_3811);
nand U4126 (N_4126,N_3849,N_3856);
or U4127 (N_4127,N_3815,N_3917);
nand U4128 (N_4128,N_3937,N_3980);
xor U4129 (N_4129,N_3853,N_3957);
nor U4130 (N_4130,N_3811,N_3996);
nor U4131 (N_4131,N_3917,N_3887);
and U4132 (N_4132,N_3958,N_3836);
and U4133 (N_4133,N_3843,N_3946);
or U4134 (N_4134,N_3921,N_3856);
or U4135 (N_4135,N_3945,N_3833);
nor U4136 (N_4136,N_3891,N_3848);
or U4137 (N_4137,N_3877,N_3826);
nor U4138 (N_4138,N_3990,N_3863);
nor U4139 (N_4139,N_3910,N_3912);
xnor U4140 (N_4140,N_3851,N_3986);
or U4141 (N_4141,N_3878,N_3985);
xor U4142 (N_4142,N_3965,N_3944);
xor U4143 (N_4143,N_3965,N_3821);
and U4144 (N_4144,N_3991,N_3975);
nand U4145 (N_4145,N_3930,N_3861);
or U4146 (N_4146,N_3958,N_3870);
xnor U4147 (N_4147,N_3880,N_3998);
and U4148 (N_4148,N_3816,N_3800);
and U4149 (N_4149,N_3894,N_3848);
xnor U4150 (N_4150,N_3849,N_3890);
nand U4151 (N_4151,N_3829,N_3888);
and U4152 (N_4152,N_3982,N_3965);
xnor U4153 (N_4153,N_3809,N_3896);
and U4154 (N_4154,N_3833,N_3812);
or U4155 (N_4155,N_3805,N_3946);
or U4156 (N_4156,N_3823,N_3849);
and U4157 (N_4157,N_3963,N_3857);
xnor U4158 (N_4158,N_3930,N_3914);
and U4159 (N_4159,N_3845,N_3880);
nand U4160 (N_4160,N_3906,N_3993);
nor U4161 (N_4161,N_3878,N_3958);
nand U4162 (N_4162,N_3873,N_3892);
nor U4163 (N_4163,N_3816,N_3912);
nor U4164 (N_4164,N_3994,N_3921);
or U4165 (N_4165,N_3988,N_3970);
nand U4166 (N_4166,N_3830,N_3855);
and U4167 (N_4167,N_3822,N_3862);
and U4168 (N_4168,N_3879,N_3958);
nor U4169 (N_4169,N_3832,N_3957);
or U4170 (N_4170,N_3986,N_3823);
xnor U4171 (N_4171,N_3993,N_3820);
xor U4172 (N_4172,N_3955,N_3980);
xnor U4173 (N_4173,N_3919,N_3957);
nor U4174 (N_4174,N_3989,N_3937);
and U4175 (N_4175,N_3987,N_3943);
nand U4176 (N_4176,N_3851,N_3997);
nand U4177 (N_4177,N_3922,N_3984);
nor U4178 (N_4178,N_3874,N_3806);
nor U4179 (N_4179,N_3809,N_3822);
nor U4180 (N_4180,N_3903,N_3944);
nand U4181 (N_4181,N_3885,N_3818);
nor U4182 (N_4182,N_3956,N_3841);
nor U4183 (N_4183,N_3955,N_3801);
or U4184 (N_4184,N_3914,N_3842);
or U4185 (N_4185,N_3938,N_3937);
nor U4186 (N_4186,N_3983,N_3822);
xor U4187 (N_4187,N_3924,N_3887);
and U4188 (N_4188,N_3974,N_3982);
and U4189 (N_4189,N_3847,N_3806);
nor U4190 (N_4190,N_3810,N_3900);
xnor U4191 (N_4191,N_3840,N_3864);
or U4192 (N_4192,N_3808,N_3954);
nand U4193 (N_4193,N_3994,N_3802);
xor U4194 (N_4194,N_3861,N_3909);
or U4195 (N_4195,N_3982,N_3895);
nor U4196 (N_4196,N_3852,N_3982);
nand U4197 (N_4197,N_3855,N_3910);
xnor U4198 (N_4198,N_3896,N_3999);
xnor U4199 (N_4199,N_3901,N_3996);
nand U4200 (N_4200,N_4057,N_4115);
and U4201 (N_4201,N_4103,N_4097);
nand U4202 (N_4202,N_4063,N_4032);
and U4203 (N_4203,N_4102,N_4141);
or U4204 (N_4204,N_4125,N_4154);
and U4205 (N_4205,N_4126,N_4164);
nand U4206 (N_4206,N_4199,N_4105);
nor U4207 (N_4207,N_4124,N_4040);
or U4208 (N_4208,N_4116,N_4119);
or U4209 (N_4209,N_4118,N_4023);
nor U4210 (N_4210,N_4046,N_4019);
xnor U4211 (N_4211,N_4198,N_4131);
or U4212 (N_4212,N_4050,N_4184);
and U4213 (N_4213,N_4088,N_4128);
xor U4214 (N_4214,N_4052,N_4015);
or U4215 (N_4215,N_4082,N_4086);
nor U4216 (N_4216,N_4087,N_4129);
and U4217 (N_4217,N_4009,N_4068);
xnor U4218 (N_4218,N_4186,N_4172);
or U4219 (N_4219,N_4000,N_4005);
nand U4220 (N_4220,N_4085,N_4021);
or U4221 (N_4221,N_4193,N_4147);
xor U4222 (N_4222,N_4190,N_4002);
and U4223 (N_4223,N_4142,N_4001);
and U4224 (N_4224,N_4048,N_4170);
nor U4225 (N_4225,N_4174,N_4194);
nor U4226 (N_4226,N_4155,N_4010);
xor U4227 (N_4227,N_4197,N_4069);
nand U4228 (N_4228,N_4030,N_4123);
or U4229 (N_4229,N_4045,N_4058);
or U4230 (N_4230,N_4064,N_4031);
xnor U4231 (N_4231,N_4027,N_4127);
or U4232 (N_4232,N_4113,N_4067);
and U4233 (N_4233,N_4008,N_4051);
nand U4234 (N_4234,N_4036,N_4077);
or U4235 (N_4235,N_4081,N_4042);
xnor U4236 (N_4236,N_4162,N_4017);
nor U4237 (N_4237,N_4156,N_4028);
or U4238 (N_4238,N_4062,N_4139);
nor U4239 (N_4239,N_4054,N_4151);
xor U4240 (N_4240,N_4003,N_4158);
and U4241 (N_4241,N_4065,N_4178);
and U4242 (N_4242,N_4099,N_4132);
or U4243 (N_4243,N_4181,N_4034);
xnor U4244 (N_4244,N_4183,N_4080);
or U4245 (N_4245,N_4144,N_4136);
nand U4246 (N_4246,N_4177,N_4020);
nand U4247 (N_4247,N_4145,N_4029);
xnor U4248 (N_4248,N_4006,N_4189);
or U4249 (N_4249,N_4038,N_4195);
nand U4250 (N_4250,N_4133,N_4075);
xor U4251 (N_4251,N_4161,N_4140);
xnor U4252 (N_4252,N_4166,N_4153);
nor U4253 (N_4253,N_4121,N_4060);
and U4254 (N_4254,N_4025,N_4175);
or U4255 (N_4255,N_4150,N_4106);
nand U4256 (N_4256,N_4092,N_4047);
nor U4257 (N_4257,N_4059,N_4196);
nand U4258 (N_4258,N_4111,N_4188);
nor U4259 (N_4259,N_4096,N_4192);
nand U4260 (N_4260,N_4110,N_4101);
and U4261 (N_4261,N_4041,N_4169);
and U4262 (N_4262,N_4095,N_4146);
or U4263 (N_4263,N_4130,N_4039);
and U4264 (N_4264,N_4149,N_4182);
and U4265 (N_4265,N_4070,N_4035);
or U4266 (N_4266,N_4013,N_4094);
and U4267 (N_4267,N_4044,N_4104);
or U4268 (N_4268,N_4168,N_4076);
xnor U4269 (N_4269,N_4083,N_4163);
nor U4270 (N_4270,N_4148,N_4157);
nand U4271 (N_4271,N_4091,N_4066);
or U4272 (N_4272,N_4138,N_4143);
nand U4273 (N_4273,N_4072,N_4179);
nand U4274 (N_4274,N_4185,N_4098);
xor U4275 (N_4275,N_4089,N_4078);
nand U4276 (N_4276,N_4159,N_4090);
xor U4277 (N_4277,N_4016,N_4173);
and U4278 (N_4278,N_4037,N_4167);
and U4279 (N_4279,N_4117,N_4043);
and U4280 (N_4280,N_4176,N_4120);
and U4281 (N_4281,N_4093,N_4109);
xnor U4282 (N_4282,N_4053,N_4112);
xor U4283 (N_4283,N_4160,N_4011);
nand U4284 (N_4284,N_4122,N_4107);
and U4285 (N_4285,N_4171,N_4055);
and U4286 (N_4286,N_4187,N_4071);
or U4287 (N_4287,N_4018,N_4022);
xnor U4288 (N_4288,N_4014,N_4061);
xnor U4289 (N_4289,N_4007,N_4073);
or U4290 (N_4290,N_4165,N_4152);
nor U4291 (N_4291,N_4024,N_4114);
or U4292 (N_4292,N_4100,N_4135);
or U4293 (N_4293,N_4079,N_4033);
or U4294 (N_4294,N_4012,N_4074);
xor U4295 (N_4295,N_4191,N_4049);
nor U4296 (N_4296,N_4180,N_4137);
and U4297 (N_4297,N_4056,N_4004);
and U4298 (N_4298,N_4026,N_4084);
nand U4299 (N_4299,N_4134,N_4108);
xor U4300 (N_4300,N_4099,N_4055);
nand U4301 (N_4301,N_4150,N_4194);
and U4302 (N_4302,N_4098,N_4065);
nor U4303 (N_4303,N_4106,N_4135);
nand U4304 (N_4304,N_4189,N_4030);
and U4305 (N_4305,N_4066,N_4051);
nand U4306 (N_4306,N_4143,N_4001);
or U4307 (N_4307,N_4168,N_4088);
or U4308 (N_4308,N_4089,N_4190);
nor U4309 (N_4309,N_4018,N_4065);
xnor U4310 (N_4310,N_4165,N_4002);
xnor U4311 (N_4311,N_4111,N_4198);
and U4312 (N_4312,N_4096,N_4064);
xnor U4313 (N_4313,N_4095,N_4021);
xnor U4314 (N_4314,N_4143,N_4044);
xnor U4315 (N_4315,N_4145,N_4179);
xnor U4316 (N_4316,N_4085,N_4032);
or U4317 (N_4317,N_4007,N_4114);
nand U4318 (N_4318,N_4044,N_4156);
or U4319 (N_4319,N_4042,N_4176);
or U4320 (N_4320,N_4042,N_4044);
nand U4321 (N_4321,N_4191,N_4107);
and U4322 (N_4322,N_4084,N_4193);
xnor U4323 (N_4323,N_4102,N_4086);
or U4324 (N_4324,N_4194,N_4187);
and U4325 (N_4325,N_4039,N_4075);
xnor U4326 (N_4326,N_4138,N_4137);
nand U4327 (N_4327,N_4088,N_4176);
nand U4328 (N_4328,N_4000,N_4082);
or U4329 (N_4329,N_4077,N_4017);
xnor U4330 (N_4330,N_4135,N_4147);
or U4331 (N_4331,N_4074,N_4106);
nor U4332 (N_4332,N_4071,N_4138);
or U4333 (N_4333,N_4160,N_4134);
nor U4334 (N_4334,N_4125,N_4177);
nor U4335 (N_4335,N_4139,N_4137);
or U4336 (N_4336,N_4123,N_4062);
nand U4337 (N_4337,N_4199,N_4116);
and U4338 (N_4338,N_4037,N_4152);
or U4339 (N_4339,N_4006,N_4149);
nor U4340 (N_4340,N_4181,N_4185);
nor U4341 (N_4341,N_4137,N_4090);
or U4342 (N_4342,N_4171,N_4159);
nand U4343 (N_4343,N_4084,N_4036);
nor U4344 (N_4344,N_4197,N_4122);
nor U4345 (N_4345,N_4059,N_4042);
or U4346 (N_4346,N_4122,N_4044);
nand U4347 (N_4347,N_4189,N_4167);
and U4348 (N_4348,N_4150,N_4079);
and U4349 (N_4349,N_4022,N_4033);
or U4350 (N_4350,N_4064,N_4154);
nor U4351 (N_4351,N_4003,N_4129);
and U4352 (N_4352,N_4172,N_4161);
nor U4353 (N_4353,N_4106,N_4039);
and U4354 (N_4354,N_4036,N_4025);
nand U4355 (N_4355,N_4133,N_4084);
nor U4356 (N_4356,N_4135,N_4159);
nand U4357 (N_4357,N_4189,N_4024);
nand U4358 (N_4358,N_4028,N_4092);
and U4359 (N_4359,N_4168,N_4053);
nand U4360 (N_4360,N_4033,N_4068);
and U4361 (N_4361,N_4001,N_4153);
and U4362 (N_4362,N_4170,N_4111);
xnor U4363 (N_4363,N_4018,N_4109);
nand U4364 (N_4364,N_4096,N_4015);
nand U4365 (N_4365,N_4026,N_4193);
nor U4366 (N_4366,N_4141,N_4034);
nor U4367 (N_4367,N_4027,N_4094);
xnor U4368 (N_4368,N_4143,N_4160);
and U4369 (N_4369,N_4060,N_4016);
and U4370 (N_4370,N_4102,N_4094);
nor U4371 (N_4371,N_4054,N_4128);
and U4372 (N_4372,N_4113,N_4017);
nor U4373 (N_4373,N_4178,N_4103);
nand U4374 (N_4374,N_4012,N_4191);
and U4375 (N_4375,N_4126,N_4185);
nand U4376 (N_4376,N_4193,N_4081);
nand U4377 (N_4377,N_4005,N_4076);
and U4378 (N_4378,N_4064,N_4177);
nand U4379 (N_4379,N_4071,N_4121);
nor U4380 (N_4380,N_4168,N_4073);
xnor U4381 (N_4381,N_4104,N_4145);
or U4382 (N_4382,N_4036,N_4038);
nor U4383 (N_4383,N_4094,N_4106);
nand U4384 (N_4384,N_4197,N_4113);
and U4385 (N_4385,N_4018,N_4195);
nand U4386 (N_4386,N_4042,N_4188);
and U4387 (N_4387,N_4057,N_4150);
nand U4388 (N_4388,N_4113,N_4014);
xor U4389 (N_4389,N_4194,N_4075);
and U4390 (N_4390,N_4122,N_4170);
or U4391 (N_4391,N_4199,N_4146);
xnor U4392 (N_4392,N_4049,N_4066);
and U4393 (N_4393,N_4172,N_4134);
xnor U4394 (N_4394,N_4184,N_4081);
xor U4395 (N_4395,N_4003,N_4047);
and U4396 (N_4396,N_4178,N_4185);
nand U4397 (N_4397,N_4121,N_4127);
xor U4398 (N_4398,N_4178,N_4116);
xor U4399 (N_4399,N_4072,N_4013);
xnor U4400 (N_4400,N_4389,N_4206);
nor U4401 (N_4401,N_4249,N_4364);
xor U4402 (N_4402,N_4202,N_4338);
or U4403 (N_4403,N_4361,N_4241);
nand U4404 (N_4404,N_4284,N_4300);
and U4405 (N_4405,N_4237,N_4355);
and U4406 (N_4406,N_4230,N_4332);
xor U4407 (N_4407,N_4330,N_4367);
nand U4408 (N_4408,N_4275,N_4253);
and U4409 (N_4409,N_4339,N_4220);
nand U4410 (N_4410,N_4320,N_4281);
and U4411 (N_4411,N_4377,N_4278);
or U4412 (N_4412,N_4395,N_4285);
nor U4413 (N_4413,N_4293,N_4274);
and U4414 (N_4414,N_4263,N_4387);
nor U4415 (N_4415,N_4318,N_4336);
xor U4416 (N_4416,N_4295,N_4335);
nor U4417 (N_4417,N_4282,N_4371);
or U4418 (N_4418,N_4217,N_4375);
xnor U4419 (N_4419,N_4399,N_4218);
or U4420 (N_4420,N_4311,N_4214);
nand U4421 (N_4421,N_4260,N_4248);
or U4422 (N_4422,N_4257,N_4326);
nand U4423 (N_4423,N_4236,N_4269);
xor U4424 (N_4424,N_4298,N_4290);
or U4425 (N_4425,N_4201,N_4359);
and U4426 (N_4426,N_4267,N_4209);
nor U4427 (N_4427,N_4229,N_4323);
and U4428 (N_4428,N_4234,N_4208);
nand U4429 (N_4429,N_4243,N_4327);
nand U4430 (N_4430,N_4291,N_4264);
nor U4431 (N_4431,N_4319,N_4381);
nand U4432 (N_4432,N_4216,N_4345);
and U4433 (N_4433,N_4391,N_4343);
xor U4434 (N_4434,N_4242,N_4346);
and U4435 (N_4435,N_4277,N_4366);
and U4436 (N_4436,N_4272,N_4350);
nand U4437 (N_4437,N_4251,N_4266);
or U4438 (N_4438,N_4380,N_4255);
nor U4439 (N_4439,N_4265,N_4382);
xor U4440 (N_4440,N_4289,N_4261);
and U4441 (N_4441,N_4205,N_4279);
nor U4442 (N_4442,N_4360,N_4273);
nand U4443 (N_4443,N_4200,N_4369);
nor U4444 (N_4444,N_4348,N_4344);
xor U4445 (N_4445,N_4259,N_4365);
and U4446 (N_4446,N_4254,N_4307);
and U4447 (N_4447,N_4398,N_4204);
and U4448 (N_4448,N_4235,N_4325);
nand U4449 (N_4449,N_4294,N_4341);
nand U4450 (N_4450,N_4283,N_4390);
xor U4451 (N_4451,N_4231,N_4312);
xnor U4452 (N_4452,N_4368,N_4340);
nand U4453 (N_4453,N_4397,N_4213);
xor U4454 (N_4454,N_4313,N_4379);
nor U4455 (N_4455,N_4219,N_4393);
xnor U4456 (N_4456,N_4386,N_4337);
nor U4457 (N_4457,N_4392,N_4210);
nand U4458 (N_4458,N_4317,N_4256);
nor U4459 (N_4459,N_4226,N_4315);
nor U4460 (N_4460,N_4252,N_4280);
xor U4461 (N_4461,N_4342,N_4246);
or U4462 (N_4462,N_4353,N_4247);
or U4463 (N_4463,N_4358,N_4357);
xnor U4464 (N_4464,N_4227,N_4212);
nand U4465 (N_4465,N_4370,N_4232);
nand U4466 (N_4466,N_4372,N_4304);
and U4467 (N_4467,N_4314,N_4238);
nand U4468 (N_4468,N_4301,N_4207);
nor U4469 (N_4469,N_4292,N_4310);
nor U4470 (N_4470,N_4245,N_4384);
and U4471 (N_4471,N_4287,N_4306);
nor U4472 (N_4472,N_4258,N_4221);
nor U4473 (N_4473,N_4268,N_4286);
xor U4474 (N_4474,N_4250,N_4303);
and U4475 (N_4475,N_4396,N_4328);
xor U4476 (N_4476,N_4374,N_4305);
and U4477 (N_4477,N_4334,N_4321);
nand U4478 (N_4478,N_4362,N_4299);
nor U4479 (N_4479,N_4352,N_4324);
and U4480 (N_4480,N_4222,N_4276);
and U4481 (N_4481,N_4233,N_4308);
or U4482 (N_4482,N_4228,N_4356);
nor U4483 (N_4483,N_4211,N_4331);
nand U4484 (N_4484,N_4316,N_4271);
xnor U4485 (N_4485,N_4224,N_4309);
or U4486 (N_4486,N_4394,N_4373);
nand U4487 (N_4487,N_4223,N_4322);
nand U4488 (N_4488,N_4385,N_4302);
and U4489 (N_4489,N_4351,N_4296);
or U4490 (N_4490,N_4225,N_4329);
nor U4491 (N_4491,N_4363,N_4297);
or U4492 (N_4492,N_4354,N_4347);
and U4493 (N_4493,N_4244,N_4378);
nor U4494 (N_4494,N_4262,N_4203);
nand U4495 (N_4495,N_4215,N_4288);
nor U4496 (N_4496,N_4376,N_4333);
and U4497 (N_4497,N_4349,N_4240);
nand U4498 (N_4498,N_4270,N_4383);
or U4499 (N_4499,N_4388,N_4239);
or U4500 (N_4500,N_4378,N_4361);
and U4501 (N_4501,N_4325,N_4392);
nand U4502 (N_4502,N_4366,N_4367);
nor U4503 (N_4503,N_4313,N_4209);
nor U4504 (N_4504,N_4217,N_4278);
xor U4505 (N_4505,N_4374,N_4330);
nor U4506 (N_4506,N_4222,N_4218);
or U4507 (N_4507,N_4354,N_4286);
nor U4508 (N_4508,N_4334,N_4293);
nand U4509 (N_4509,N_4388,N_4269);
nor U4510 (N_4510,N_4306,N_4334);
or U4511 (N_4511,N_4309,N_4249);
and U4512 (N_4512,N_4378,N_4299);
nor U4513 (N_4513,N_4383,N_4334);
nor U4514 (N_4514,N_4233,N_4343);
or U4515 (N_4515,N_4390,N_4321);
nor U4516 (N_4516,N_4205,N_4359);
nor U4517 (N_4517,N_4278,N_4233);
nand U4518 (N_4518,N_4232,N_4383);
and U4519 (N_4519,N_4242,N_4324);
xor U4520 (N_4520,N_4357,N_4229);
xor U4521 (N_4521,N_4385,N_4250);
or U4522 (N_4522,N_4232,N_4348);
and U4523 (N_4523,N_4359,N_4304);
and U4524 (N_4524,N_4381,N_4252);
nor U4525 (N_4525,N_4306,N_4302);
nor U4526 (N_4526,N_4383,N_4242);
nand U4527 (N_4527,N_4343,N_4236);
nand U4528 (N_4528,N_4361,N_4221);
or U4529 (N_4529,N_4306,N_4314);
nand U4530 (N_4530,N_4318,N_4207);
and U4531 (N_4531,N_4224,N_4228);
nor U4532 (N_4532,N_4384,N_4204);
nand U4533 (N_4533,N_4306,N_4283);
nor U4534 (N_4534,N_4207,N_4367);
and U4535 (N_4535,N_4340,N_4247);
or U4536 (N_4536,N_4372,N_4300);
and U4537 (N_4537,N_4213,N_4313);
nand U4538 (N_4538,N_4323,N_4224);
xnor U4539 (N_4539,N_4200,N_4327);
nand U4540 (N_4540,N_4323,N_4257);
nor U4541 (N_4541,N_4368,N_4208);
xnor U4542 (N_4542,N_4256,N_4282);
and U4543 (N_4543,N_4334,N_4240);
or U4544 (N_4544,N_4311,N_4227);
nand U4545 (N_4545,N_4216,N_4306);
nor U4546 (N_4546,N_4224,N_4258);
xor U4547 (N_4547,N_4308,N_4212);
xnor U4548 (N_4548,N_4341,N_4303);
xnor U4549 (N_4549,N_4210,N_4273);
nor U4550 (N_4550,N_4262,N_4334);
nand U4551 (N_4551,N_4205,N_4310);
and U4552 (N_4552,N_4373,N_4284);
or U4553 (N_4553,N_4204,N_4317);
nor U4554 (N_4554,N_4240,N_4375);
or U4555 (N_4555,N_4357,N_4362);
nand U4556 (N_4556,N_4374,N_4388);
xnor U4557 (N_4557,N_4290,N_4385);
nand U4558 (N_4558,N_4268,N_4245);
nand U4559 (N_4559,N_4308,N_4276);
and U4560 (N_4560,N_4355,N_4375);
xnor U4561 (N_4561,N_4294,N_4264);
and U4562 (N_4562,N_4366,N_4293);
xnor U4563 (N_4563,N_4308,N_4307);
nand U4564 (N_4564,N_4321,N_4335);
nand U4565 (N_4565,N_4234,N_4332);
or U4566 (N_4566,N_4253,N_4363);
and U4567 (N_4567,N_4311,N_4348);
and U4568 (N_4568,N_4328,N_4242);
nand U4569 (N_4569,N_4309,N_4208);
xnor U4570 (N_4570,N_4335,N_4239);
xor U4571 (N_4571,N_4331,N_4216);
nand U4572 (N_4572,N_4264,N_4393);
or U4573 (N_4573,N_4254,N_4322);
nor U4574 (N_4574,N_4386,N_4303);
and U4575 (N_4575,N_4347,N_4245);
nor U4576 (N_4576,N_4331,N_4321);
nor U4577 (N_4577,N_4396,N_4309);
and U4578 (N_4578,N_4273,N_4229);
and U4579 (N_4579,N_4228,N_4395);
xnor U4580 (N_4580,N_4218,N_4359);
nand U4581 (N_4581,N_4391,N_4233);
nand U4582 (N_4582,N_4371,N_4276);
nand U4583 (N_4583,N_4225,N_4366);
nor U4584 (N_4584,N_4235,N_4200);
and U4585 (N_4585,N_4365,N_4276);
and U4586 (N_4586,N_4316,N_4294);
nand U4587 (N_4587,N_4245,N_4200);
nor U4588 (N_4588,N_4351,N_4393);
nor U4589 (N_4589,N_4265,N_4366);
nor U4590 (N_4590,N_4327,N_4233);
nand U4591 (N_4591,N_4229,N_4212);
xor U4592 (N_4592,N_4372,N_4275);
nand U4593 (N_4593,N_4217,N_4238);
and U4594 (N_4594,N_4347,N_4207);
and U4595 (N_4595,N_4214,N_4383);
nor U4596 (N_4596,N_4369,N_4310);
nand U4597 (N_4597,N_4326,N_4349);
xor U4598 (N_4598,N_4273,N_4301);
nand U4599 (N_4599,N_4206,N_4351);
and U4600 (N_4600,N_4469,N_4517);
or U4601 (N_4601,N_4461,N_4552);
or U4602 (N_4602,N_4411,N_4428);
nand U4603 (N_4603,N_4454,N_4465);
or U4604 (N_4604,N_4570,N_4442);
xnor U4605 (N_4605,N_4475,N_4486);
nor U4606 (N_4606,N_4481,N_4560);
and U4607 (N_4607,N_4426,N_4439);
or U4608 (N_4608,N_4586,N_4488);
or U4609 (N_4609,N_4514,N_4527);
or U4610 (N_4610,N_4403,N_4484);
xor U4611 (N_4611,N_4513,N_4590);
and U4612 (N_4612,N_4482,N_4412);
nand U4613 (N_4613,N_4492,N_4537);
or U4614 (N_4614,N_4538,N_4447);
and U4615 (N_4615,N_4578,N_4496);
xor U4616 (N_4616,N_4456,N_4564);
or U4617 (N_4617,N_4522,N_4432);
nand U4618 (N_4618,N_4577,N_4529);
nand U4619 (N_4619,N_4446,N_4540);
or U4620 (N_4620,N_4563,N_4452);
nand U4621 (N_4621,N_4558,N_4430);
nor U4622 (N_4622,N_4471,N_4479);
or U4623 (N_4623,N_4499,N_4406);
or U4624 (N_4624,N_4501,N_4541);
or U4625 (N_4625,N_4476,N_4450);
nor U4626 (N_4626,N_4434,N_4528);
nor U4627 (N_4627,N_4555,N_4497);
and U4628 (N_4628,N_4585,N_4425);
or U4629 (N_4629,N_4444,N_4561);
nand U4630 (N_4630,N_4419,N_4485);
and U4631 (N_4631,N_4420,N_4477);
nand U4632 (N_4632,N_4505,N_4421);
nor U4633 (N_4633,N_4402,N_4569);
or U4634 (N_4634,N_4562,N_4591);
nor U4635 (N_4635,N_4531,N_4451);
nor U4636 (N_4636,N_4422,N_4512);
xor U4637 (N_4637,N_4437,N_4459);
and U4638 (N_4638,N_4427,N_4441);
and U4639 (N_4639,N_4511,N_4583);
nor U4640 (N_4640,N_4539,N_4559);
and U4641 (N_4641,N_4523,N_4519);
and U4642 (N_4642,N_4460,N_4556);
and U4643 (N_4643,N_4545,N_4515);
nand U4644 (N_4644,N_4478,N_4438);
xnor U4645 (N_4645,N_4580,N_4551);
xnor U4646 (N_4646,N_4500,N_4423);
nand U4647 (N_4647,N_4417,N_4453);
or U4648 (N_4648,N_4581,N_4468);
xnor U4649 (N_4649,N_4400,N_4494);
or U4650 (N_4650,N_4553,N_4463);
xnor U4651 (N_4651,N_4487,N_4470);
or U4652 (N_4652,N_4436,N_4507);
xor U4653 (N_4653,N_4582,N_4567);
xor U4654 (N_4654,N_4464,N_4589);
or U4655 (N_4655,N_4588,N_4592);
and U4656 (N_4656,N_4415,N_4466);
nor U4657 (N_4657,N_4440,N_4554);
nand U4658 (N_4658,N_4533,N_4435);
nand U4659 (N_4659,N_4579,N_4546);
nand U4660 (N_4660,N_4472,N_4535);
or U4661 (N_4661,N_4498,N_4491);
xnor U4662 (N_4662,N_4408,N_4424);
nand U4663 (N_4663,N_4532,N_4599);
or U4664 (N_4664,N_4508,N_4502);
nor U4665 (N_4665,N_4429,N_4473);
and U4666 (N_4666,N_4548,N_4509);
nor U4667 (N_4667,N_4542,N_4516);
and U4668 (N_4668,N_4587,N_4534);
nor U4669 (N_4669,N_4490,N_4445);
and U4670 (N_4670,N_4565,N_4489);
nand U4671 (N_4671,N_4433,N_4594);
xnor U4672 (N_4672,N_4449,N_4404);
or U4673 (N_4673,N_4536,N_4524);
nor U4674 (N_4674,N_4480,N_4547);
and U4675 (N_4675,N_4566,N_4557);
or U4676 (N_4676,N_4530,N_4503);
xnor U4677 (N_4677,N_4483,N_4455);
and U4678 (N_4678,N_4584,N_4598);
and U4679 (N_4679,N_4593,N_4574);
or U4680 (N_4680,N_4568,N_4504);
nand U4681 (N_4681,N_4443,N_4595);
nand U4682 (N_4682,N_4543,N_4576);
nand U4683 (N_4683,N_4495,N_4413);
nor U4684 (N_4684,N_4571,N_4418);
and U4685 (N_4685,N_4573,N_4474);
nand U4686 (N_4686,N_4462,N_4405);
xnor U4687 (N_4687,N_4521,N_4410);
xor U4688 (N_4688,N_4448,N_4575);
or U4689 (N_4689,N_4457,N_4549);
and U4690 (N_4690,N_4431,N_4525);
nand U4691 (N_4691,N_4544,N_4550);
nor U4692 (N_4692,N_4493,N_4597);
or U4693 (N_4693,N_4416,N_4510);
xor U4694 (N_4694,N_4467,N_4518);
nand U4695 (N_4695,N_4407,N_4401);
nor U4696 (N_4696,N_4520,N_4596);
nand U4697 (N_4697,N_4506,N_4458);
nand U4698 (N_4698,N_4572,N_4526);
or U4699 (N_4699,N_4409,N_4414);
xnor U4700 (N_4700,N_4568,N_4501);
nand U4701 (N_4701,N_4439,N_4498);
nor U4702 (N_4702,N_4463,N_4485);
nor U4703 (N_4703,N_4512,N_4545);
and U4704 (N_4704,N_4501,N_4580);
and U4705 (N_4705,N_4468,N_4414);
xnor U4706 (N_4706,N_4479,N_4508);
xor U4707 (N_4707,N_4473,N_4513);
nand U4708 (N_4708,N_4418,N_4537);
and U4709 (N_4709,N_4538,N_4461);
nor U4710 (N_4710,N_4521,N_4564);
and U4711 (N_4711,N_4457,N_4423);
nor U4712 (N_4712,N_4506,N_4580);
nor U4713 (N_4713,N_4466,N_4506);
xnor U4714 (N_4714,N_4557,N_4404);
nor U4715 (N_4715,N_4514,N_4491);
xnor U4716 (N_4716,N_4420,N_4508);
and U4717 (N_4717,N_4467,N_4403);
and U4718 (N_4718,N_4466,N_4535);
nor U4719 (N_4719,N_4407,N_4560);
nand U4720 (N_4720,N_4462,N_4551);
nand U4721 (N_4721,N_4438,N_4550);
nand U4722 (N_4722,N_4483,N_4465);
xnor U4723 (N_4723,N_4548,N_4491);
and U4724 (N_4724,N_4491,N_4540);
or U4725 (N_4725,N_4474,N_4558);
and U4726 (N_4726,N_4567,N_4442);
nor U4727 (N_4727,N_4450,N_4527);
nand U4728 (N_4728,N_4459,N_4420);
or U4729 (N_4729,N_4589,N_4592);
xnor U4730 (N_4730,N_4427,N_4414);
xor U4731 (N_4731,N_4599,N_4492);
or U4732 (N_4732,N_4400,N_4596);
and U4733 (N_4733,N_4589,N_4408);
nor U4734 (N_4734,N_4406,N_4435);
nand U4735 (N_4735,N_4524,N_4486);
and U4736 (N_4736,N_4473,N_4447);
or U4737 (N_4737,N_4512,N_4572);
or U4738 (N_4738,N_4486,N_4496);
nor U4739 (N_4739,N_4428,N_4432);
or U4740 (N_4740,N_4569,N_4589);
nor U4741 (N_4741,N_4581,N_4452);
and U4742 (N_4742,N_4401,N_4436);
xor U4743 (N_4743,N_4458,N_4550);
xor U4744 (N_4744,N_4594,N_4457);
or U4745 (N_4745,N_4570,N_4414);
xor U4746 (N_4746,N_4545,N_4514);
xnor U4747 (N_4747,N_4588,N_4457);
xnor U4748 (N_4748,N_4456,N_4411);
xnor U4749 (N_4749,N_4456,N_4578);
xnor U4750 (N_4750,N_4474,N_4513);
xor U4751 (N_4751,N_4420,N_4530);
xnor U4752 (N_4752,N_4413,N_4554);
nand U4753 (N_4753,N_4414,N_4459);
nand U4754 (N_4754,N_4591,N_4447);
nand U4755 (N_4755,N_4585,N_4482);
xnor U4756 (N_4756,N_4450,N_4434);
or U4757 (N_4757,N_4434,N_4584);
xor U4758 (N_4758,N_4410,N_4561);
or U4759 (N_4759,N_4403,N_4415);
xor U4760 (N_4760,N_4470,N_4570);
xnor U4761 (N_4761,N_4473,N_4482);
nor U4762 (N_4762,N_4498,N_4422);
nand U4763 (N_4763,N_4432,N_4493);
nor U4764 (N_4764,N_4401,N_4517);
xor U4765 (N_4765,N_4538,N_4419);
xnor U4766 (N_4766,N_4541,N_4469);
nand U4767 (N_4767,N_4408,N_4597);
or U4768 (N_4768,N_4598,N_4543);
or U4769 (N_4769,N_4547,N_4404);
nand U4770 (N_4770,N_4515,N_4500);
xnor U4771 (N_4771,N_4434,N_4508);
nand U4772 (N_4772,N_4555,N_4400);
nor U4773 (N_4773,N_4574,N_4473);
or U4774 (N_4774,N_4434,N_4497);
or U4775 (N_4775,N_4576,N_4415);
and U4776 (N_4776,N_4537,N_4577);
and U4777 (N_4777,N_4571,N_4598);
xor U4778 (N_4778,N_4406,N_4460);
nand U4779 (N_4779,N_4486,N_4489);
nand U4780 (N_4780,N_4525,N_4529);
nand U4781 (N_4781,N_4536,N_4529);
and U4782 (N_4782,N_4473,N_4492);
xor U4783 (N_4783,N_4519,N_4514);
and U4784 (N_4784,N_4414,N_4509);
and U4785 (N_4785,N_4402,N_4560);
nor U4786 (N_4786,N_4531,N_4447);
nand U4787 (N_4787,N_4465,N_4416);
and U4788 (N_4788,N_4577,N_4430);
and U4789 (N_4789,N_4478,N_4589);
or U4790 (N_4790,N_4538,N_4597);
xnor U4791 (N_4791,N_4564,N_4443);
xnor U4792 (N_4792,N_4592,N_4584);
nand U4793 (N_4793,N_4458,N_4472);
nor U4794 (N_4794,N_4401,N_4557);
and U4795 (N_4795,N_4421,N_4480);
or U4796 (N_4796,N_4443,N_4466);
and U4797 (N_4797,N_4466,N_4578);
xnor U4798 (N_4798,N_4406,N_4554);
or U4799 (N_4799,N_4414,N_4540);
nand U4800 (N_4800,N_4722,N_4777);
and U4801 (N_4801,N_4702,N_4798);
and U4802 (N_4802,N_4757,N_4713);
nor U4803 (N_4803,N_4678,N_4668);
nand U4804 (N_4804,N_4635,N_4696);
nand U4805 (N_4805,N_4746,N_4624);
xnor U4806 (N_4806,N_4787,N_4791);
nor U4807 (N_4807,N_4756,N_4754);
nor U4808 (N_4808,N_4701,N_4730);
nor U4809 (N_4809,N_4737,N_4627);
xnor U4810 (N_4810,N_4688,N_4751);
nand U4811 (N_4811,N_4610,N_4645);
xor U4812 (N_4812,N_4646,N_4775);
xor U4813 (N_4813,N_4729,N_4774);
nand U4814 (N_4814,N_4733,N_4652);
nand U4815 (N_4815,N_4738,N_4602);
xnor U4816 (N_4816,N_4622,N_4643);
nor U4817 (N_4817,N_4683,N_4648);
nand U4818 (N_4818,N_4640,N_4694);
nand U4819 (N_4819,N_4749,N_4785);
nor U4820 (N_4820,N_4634,N_4747);
nand U4821 (N_4821,N_4772,N_4623);
and U4822 (N_4822,N_4709,N_4795);
or U4823 (N_4823,N_4677,N_4669);
and U4824 (N_4824,N_4748,N_4676);
or U4825 (N_4825,N_4674,N_4614);
or U4826 (N_4826,N_4673,N_4761);
and U4827 (N_4827,N_4712,N_4717);
nand U4828 (N_4828,N_4734,N_4707);
and U4829 (N_4829,N_4641,N_4788);
nor U4830 (N_4830,N_4708,N_4609);
or U4831 (N_4831,N_4690,N_4784);
or U4832 (N_4832,N_4631,N_4719);
or U4833 (N_4833,N_4799,N_4782);
or U4834 (N_4834,N_4778,N_4618);
or U4835 (N_4835,N_4762,N_4685);
and U4836 (N_4836,N_4693,N_4695);
nand U4837 (N_4837,N_4796,N_4632);
xnor U4838 (N_4838,N_4764,N_4759);
nor U4839 (N_4839,N_4604,N_4611);
nand U4840 (N_4840,N_4682,N_4692);
and U4841 (N_4841,N_4630,N_4792);
nor U4842 (N_4842,N_4689,N_4658);
or U4843 (N_4843,N_4654,N_4686);
nor U4844 (N_4844,N_4711,N_4663);
or U4845 (N_4845,N_4731,N_4606);
nand U4846 (N_4846,N_4664,N_4650);
or U4847 (N_4847,N_4714,N_4638);
xnor U4848 (N_4848,N_4727,N_4655);
and U4849 (N_4849,N_4710,N_4681);
or U4850 (N_4850,N_4769,N_4703);
and U4851 (N_4851,N_4720,N_4662);
or U4852 (N_4852,N_4705,N_4755);
xor U4853 (N_4853,N_4697,N_4607);
and U4854 (N_4854,N_4716,N_4753);
or U4855 (N_4855,N_4653,N_4789);
nand U4856 (N_4856,N_4626,N_4691);
or U4857 (N_4857,N_4671,N_4770);
xor U4858 (N_4858,N_4642,N_4615);
or U4859 (N_4859,N_4699,N_4732);
xnor U4860 (N_4860,N_4659,N_4735);
xnor U4861 (N_4861,N_4667,N_4752);
nand U4862 (N_4862,N_4763,N_4780);
or U4863 (N_4863,N_4684,N_4715);
and U4864 (N_4864,N_4700,N_4793);
xnor U4865 (N_4865,N_4726,N_4600);
xnor U4866 (N_4866,N_4625,N_4629);
or U4867 (N_4867,N_4612,N_4617);
xnor U4868 (N_4868,N_4794,N_4698);
xnor U4869 (N_4869,N_4644,N_4790);
nand U4870 (N_4870,N_4721,N_4706);
nor U4871 (N_4871,N_4783,N_4767);
nor U4872 (N_4872,N_4724,N_4637);
xnor U4873 (N_4873,N_4741,N_4776);
xor U4874 (N_4874,N_4744,N_4639);
xnor U4875 (N_4875,N_4723,N_4661);
and U4876 (N_4876,N_4675,N_4740);
nand U4877 (N_4877,N_4743,N_4768);
nand U4878 (N_4878,N_4771,N_4704);
nor U4879 (N_4879,N_4670,N_4725);
nand U4880 (N_4880,N_4613,N_4633);
nor U4881 (N_4881,N_4773,N_4601);
nand U4882 (N_4882,N_4750,N_4728);
xor U4883 (N_4883,N_4758,N_4636);
or U4884 (N_4884,N_4742,N_4781);
nor U4885 (N_4885,N_4603,N_4679);
and U4886 (N_4886,N_4628,N_4665);
nand U4887 (N_4887,N_4620,N_4760);
and U4888 (N_4888,N_4786,N_4765);
or U4889 (N_4889,N_4797,N_4739);
nor U4890 (N_4890,N_4657,N_4660);
and U4891 (N_4891,N_4672,N_4766);
and U4892 (N_4892,N_4619,N_4649);
nand U4893 (N_4893,N_4680,N_4651);
and U4894 (N_4894,N_4718,N_4779);
xor U4895 (N_4895,N_4745,N_4605);
xor U4896 (N_4896,N_4608,N_4687);
nand U4897 (N_4897,N_4736,N_4647);
nand U4898 (N_4898,N_4621,N_4616);
xor U4899 (N_4899,N_4666,N_4656);
or U4900 (N_4900,N_4758,N_4674);
xnor U4901 (N_4901,N_4731,N_4730);
and U4902 (N_4902,N_4703,N_4733);
xnor U4903 (N_4903,N_4683,N_4716);
and U4904 (N_4904,N_4629,N_4692);
nand U4905 (N_4905,N_4600,N_4724);
and U4906 (N_4906,N_4788,N_4677);
or U4907 (N_4907,N_4678,N_4655);
or U4908 (N_4908,N_4797,N_4704);
or U4909 (N_4909,N_4636,N_4694);
or U4910 (N_4910,N_4630,N_4784);
xnor U4911 (N_4911,N_4711,N_4797);
or U4912 (N_4912,N_4675,N_4707);
nor U4913 (N_4913,N_4636,N_4627);
nor U4914 (N_4914,N_4693,N_4678);
or U4915 (N_4915,N_4642,N_4714);
nand U4916 (N_4916,N_4669,N_4707);
xnor U4917 (N_4917,N_4755,N_4731);
xor U4918 (N_4918,N_4708,N_4635);
or U4919 (N_4919,N_4692,N_4711);
or U4920 (N_4920,N_4707,N_4697);
xnor U4921 (N_4921,N_4660,N_4738);
nor U4922 (N_4922,N_4762,N_4681);
nor U4923 (N_4923,N_4709,N_4652);
nor U4924 (N_4924,N_4782,N_4769);
and U4925 (N_4925,N_4779,N_4618);
and U4926 (N_4926,N_4781,N_4620);
and U4927 (N_4927,N_4633,N_4761);
xnor U4928 (N_4928,N_4621,N_4678);
or U4929 (N_4929,N_4676,N_4700);
xnor U4930 (N_4930,N_4606,N_4658);
or U4931 (N_4931,N_4643,N_4764);
xor U4932 (N_4932,N_4741,N_4785);
xor U4933 (N_4933,N_4610,N_4695);
or U4934 (N_4934,N_4780,N_4681);
and U4935 (N_4935,N_4608,N_4626);
and U4936 (N_4936,N_4768,N_4713);
and U4937 (N_4937,N_4712,N_4766);
and U4938 (N_4938,N_4692,N_4683);
nand U4939 (N_4939,N_4790,N_4729);
and U4940 (N_4940,N_4608,N_4681);
or U4941 (N_4941,N_4667,N_4643);
nand U4942 (N_4942,N_4672,N_4669);
nand U4943 (N_4943,N_4669,N_4663);
or U4944 (N_4944,N_4682,N_4716);
and U4945 (N_4945,N_4624,N_4644);
nor U4946 (N_4946,N_4604,N_4654);
nor U4947 (N_4947,N_4715,N_4658);
xnor U4948 (N_4948,N_4696,N_4764);
nand U4949 (N_4949,N_4776,N_4609);
nor U4950 (N_4950,N_4681,N_4627);
or U4951 (N_4951,N_4681,N_4701);
and U4952 (N_4952,N_4682,N_4617);
xnor U4953 (N_4953,N_4614,N_4708);
nand U4954 (N_4954,N_4663,N_4665);
nand U4955 (N_4955,N_4626,N_4614);
or U4956 (N_4956,N_4633,N_4739);
and U4957 (N_4957,N_4673,N_4764);
nand U4958 (N_4958,N_4684,N_4644);
or U4959 (N_4959,N_4612,N_4701);
nor U4960 (N_4960,N_4725,N_4637);
nor U4961 (N_4961,N_4639,N_4749);
nor U4962 (N_4962,N_4684,N_4630);
nor U4963 (N_4963,N_4656,N_4714);
or U4964 (N_4964,N_4738,N_4784);
nor U4965 (N_4965,N_4687,N_4703);
nand U4966 (N_4966,N_4757,N_4676);
or U4967 (N_4967,N_4777,N_4728);
nor U4968 (N_4968,N_4695,N_4788);
or U4969 (N_4969,N_4682,N_4641);
xor U4970 (N_4970,N_4696,N_4624);
nand U4971 (N_4971,N_4710,N_4738);
and U4972 (N_4972,N_4750,N_4665);
nand U4973 (N_4973,N_4796,N_4608);
and U4974 (N_4974,N_4659,N_4631);
xnor U4975 (N_4975,N_4784,N_4620);
and U4976 (N_4976,N_4718,N_4678);
nand U4977 (N_4977,N_4600,N_4681);
nor U4978 (N_4978,N_4652,N_4796);
or U4979 (N_4979,N_4688,N_4632);
nand U4980 (N_4980,N_4789,N_4703);
nor U4981 (N_4981,N_4721,N_4677);
nor U4982 (N_4982,N_4663,N_4612);
or U4983 (N_4983,N_4655,N_4638);
nor U4984 (N_4984,N_4738,N_4765);
nor U4985 (N_4985,N_4765,N_4684);
nand U4986 (N_4986,N_4720,N_4799);
or U4987 (N_4987,N_4649,N_4713);
or U4988 (N_4988,N_4601,N_4609);
nand U4989 (N_4989,N_4655,N_4725);
nand U4990 (N_4990,N_4718,N_4666);
xnor U4991 (N_4991,N_4731,N_4610);
and U4992 (N_4992,N_4743,N_4733);
nor U4993 (N_4993,N_4743,N_4742);
or U4994 (N_4994,N_4618,N_4741);
xor U4995 (N_4995,N_4615,N_4602);
or U4996 (N_4996,N_4701,N_4700);
or U4997 (N_4997,N_4676,N_4607);
xor U4998 (N_4998,N_4636,N_4794);
and U4999 (N_4999,N_4613,N_4790);
and U5000 (N_5000,N_4962,N_4808);
xnor U5001 (N_5001,N_4975,N_4848);
nand U5002 (N_5002,N_4915,N_4911);
xnor U5003 (N_5003,N_4822,N_4994);
or U5004 (N_5004,N_4931,N_4857);
nand U5005 (N_5005,N_4886,N_4988);
and U5006 (N_5006,N_4819,N_4809);
or U5007 (N_5007,N_4800,N_4982);
nor U5008 (N_5008,N_4804,N_4969);
nor U5009 (N_5009,N_4906,N_4901);
or U5010 (N_5010,N_4999,N_4944);
and U5011 (N_5011,N_4806,N_4871);
nor U5012 (N_5012,N_4889,N_4813);
or U5013 (N_5013,N_4948,N_4960);
nor U5014 (N_5014,N_4971,N_4963);
nand U5015 (N_5015,N_4966,N_4843);
or U5016 (N_5016,N_4900,N_4974);
and U5017 (N_5017,N_4905,N_4981);
nor U5018 (N_5018,N_4851,N_4841);
and U5019 (N_5019,N_4883,N_4874);
xnor U5020 (N_5020,N_4842,N_4965);
nand U5021 (N_5021,N_4818,N_4876);
or U5022 (N_5022,N_4890,N_4908);
nand U5023 (N_5023,N_4891,N_4961);
xor U5024 (N_5024,N_4922,N_4924);
and U5025 (N_5025,N_4898,N_4847);
nand U5026 (N_5026,N_4882,N_4985);
xor U5027 (N_5027,N_4826,N_4836);
nor U5028 (N_5028,N_4941,N_4954);
and U5029 (N_5029,N_4824,N_4881);
nor U5030 (N_5030,N_4863,N_4921);
or U5031 (N_5031,N_4932,N_4872);
nand U5032 (N_5032,N_4927,N_4946);
or U5033 (N_5033,N_4992,N_4828);
and U5034 (N_5034,N_4861,N_4839);
nor U5035 (N_5035,N_4814,N_4856);
nand U5036 (N_5036,N_4973,N_4917);
xnor U5037 (N_5037,N_4895,N_4972);
or U5038 (N_5038,N_4850,N_4949);
or U5039 (N_5039,N_4940,N_4964);
and U5040 (N_5040,N_4860,N_4945);
xor U5041 (N_5041,N_4928,N_4845);
and U5042 (N_5042,N_4866,N_4957);
or U5043 (N_5043,N_4884,N_4996);
or U5044 (N_5044,N_4914,N_4879);
xnor U5045 (N_5045,N_4993,N_4936);
nand U5046 (N_5046,N_4862,N_4838);
xnor U5047 (N_5047,N_4849,N_4893);
and U5048 (N_5048,N_4978,N_4892);
and U5049 (N_5049,N_4919,N_4875);
xnor U5050 (N_5050,N_4833,N_4991);
and U5051 (N_5051,N_4853,N_4858);
or U5052 (N_5052,N_4897,N_4997);
xor U5053 (N_5053,N_4854,N_4986);
or U5054 (N_5054,N_4953,N_4868);
or U5055 (N_5055,N_4916,N_4930);
xor U5056 (N_5056,N_4955,N_4820);
nor U5057 (N_5057,N_4811,N_4980);
and U5058 (N_5058,N_4888,N_4837);
and U5059 (N_5059,N_4815,N_4933);
and U5060 (N_5060,N_4816,N_4947);
xor U5061 (N_5061,N_4937,N_4817);
or U5062 (N_5062,N_4958,N_4977);
nor U5063 (N_5063,N_4967,N_4987);
and U5064 (N_5064,N_4878,N_4976);
nand U5065 (N_5065,N_4925,N_4865);
xnor U5066 (N_5066,N_4912,N_4909);
nand U5067 (N_5067,N_4802,N_4807);
xnor U5068 (N_5068,N_4835,N_4867);
or U5069 (N_5069,N_4801,N_4942);
nand U5070 (N_5070,N_4823,N_4864);
nor U5071 (N_5071,N_4840,N_4952);
nor U5072 (N_5072,N_4873,N_4910);
or U5073 (N_5073,N_4810,N_4812);
nor U5074 (N_5074,N_4984,N_4877);
and U5075 (N_5075,N_4929,N_4903);
and U5076 (N_5076,N_4998,N_4902);
xnor U5077 (N_5077,N_4913,N_4956);
xnor U5078 (N_5078,N_4894,N_4899);
nor U5079 (N_5079,N_4803,N_4904);
nor U5080 (N_5080,N_4943,N_4995);
and U5081 (N_5081,N_4844,N_4968);
xor U5082 (N_5082,N_4870,N_4859);
nand U5083 (N_5083,N_4869,N_4830);
or U5084 (N_5084,N_4983,N_4950);
nor U5085 (N_5085,N_4880,N_4938);
and U5086 (N_5086,N_4935,N_4923);
nor U5087 (N_5087,N_4887,N_4907);
nor U5088 (N_5088,N_4827,N_4852);
or U5089 (N_5089,N_4959,N_4834);
or U5090 (N_5090,N_4829,N_4920);
or U5091 (N_5091,N_4855,N_4821);
or U5092 (N_5092,N_4832,N_4970);
xor U5093 (N_5093,N_4951,N_4918);
nor U5094 (N_5094,N_4979,N_4846);
and U5095 (N_5095,N_4825,N_4885);
or U5096 (N_5096,N_4990,N_4805);
and U5097 (N_5097,N_4934,N_4926);
nand U5098 (N_5098,N_4831,N_4989);
nor U5099 (N_5099,N_4939,N_4896);
nor U5100 (N_5100,N_4807,N_4855);
xnor U5101 (N_5101,N_4896,N_4827);
xnor U5102 (N_5102,N_4932,N_4924);
or U5103 (N_5103,N_4851,N_4961);
nand U5104 (N_5104,N_4873,N_4930);
nor U5105 (N_5105,N_4859,N_4839);
xor U5106 (N_5106,N_4888,N_4962);
and U5107 (N_5107,N_4901,N_4911);
or U5108 (N_5108,N_4816,N_4885);
nor U5109 (N_5109,N_4857,N_4898);
and U5110 (N_5110,N_4951,N_4931);
xnor U5111 (N_5111,N_4943,N_4938);
or U5112 (N_5112,N_4886,N_4827);
and U5113 (N_5113,N_4862,N_4873);
and U5114 (N_5114,N_4847,N_4985);
or U5115 (N_5115,N_4946,N_4823);
and U5116 (N_5116,N_4911,N_4858);
nand U5117 (N_5117,N_4808,N_4887);
nand U5118 (N_5118,N_4802,N_4859);
xnor U5119 (N_5119,N_4873,N_4922);
nand U5120 (N_5120,N_4886,N_4945);
or U5121 (N_5121,N_4873,N_4944);
nand U5122 (N_5122,N_4992,N_4835);
nand U5123 (N_5123,N_4898,N_4929);
or U5124 (N_5124,N_4919,N_4998);
nand U5125 (N_5125,N_4925,N_4967);
nand U5126 (N_5126,N_4985,N_4820);
or U5127 (N_5127,N_4889,N_4999);
and U5128 (N_5128,N_4801,N_4805);
and U5129 (N_5129,N_4976,N_4867);
and U5130 (N_5130,N_4813,N_4969);
nor U5131 (N_5131,N_4996,N_4845);
nor U5132 (N_5132,N_4974,N_4919);
xnor U5133 (N_5133,N_4853,N_4861);
or U5134 (N_5134,N_4970,N_4999);
xor U5135 (N_5135,N_4907,N_4889);
or U5136 (N_5136,N_4968,N_4838);
nor U5137 (N_5137,N_4815,N_4806);
xnor U5138 (N_5138,N_4896,N_4986);
or U5139 (N_5139,N_4871,N_4991);
xor U5140 (N_5140,N_4837,N_4864);
or U5141 (N_5141,N_4835,N_4981);
or U5142 (N_5142,N_4976,N_4954);
xnor U5143 (N_5143,N_4998,N_4841);
xnor U5144 (N_5144,N_4818,N_4815);
xor U5145 (N_5145,N_4883,N_4895);
nand U5146 (N_5146,N_4996,N_4869);
nand U5147 (N_5147,N_4884,N_4973);
nand U5148 (N_5148,N_4948,N_4801);
nand U5149 (N_5149,N_4859,N_4985);
and U5150 (N_5150,N_4902,N_4871);
nor U5151 (N_5151,N_4820,N_4944);
or U5152 (N_5152,N_4961,N_4988);
nor U5153 (N_5153,N_4957,N_4922);
nand U5154 (N_5154,N_4973,N_4974);
nand U5155 (N_5155,N_4813,N_4861);
or U5156 (N_5156,N_4977,N_4949);
nand U5157 (N_5157,N_4982,N_4930);
nor U5158 (N_5158,N_4835,N_4991);
nand U5159 (N_5159,N_4923,N_4998);
and U5160 (N_5160,N_4867,N_4987);
nand U5161 (N_5161,N_4908,N_4919);
nand U5162 (N_5162,N_4844,N_4824);
or U5163 (N_5163,N_4938,N_4820);
and U5164 (N_5164,N_4967,N_4971);
and U5165 (N_5165,N_4975,N_4913);
xnor U5166 (N_5166,N_4982,N_4808);
or U5167 (N_5167,N_4910,N_4902);
xnor U5168 (N_5168,N_4975,N_4963);
nor U5169 (N_5169,N_4941,N_4928);
nand U5170 (N_5170,N_4832,N_4941);
nand U5171 (N_5171,N_4951,N_4873);
and U5172 (N_5172,N_4969,N_4983);
nand U5173 (N_5173,N_4945,N_4931);
xnor U5174 (N_5174,N_4958,N_4852);
nand U5175 (N_5175,N_4839,N_4971);
or U5176 (N_5176,N_4886,N_4912);
nand U5177 (N_5177,N_4809,N_4988);
nand U5178 (N_5178,N_4957,N_4967);
nor U5179 (N_5179,N_4865,N_4944);
or U5180 (N_5180,N_4828,N_4930);
and U5181 (N_5181,N_4922,N_4989);
xnor U5182 (N_5182,N_4805,N_4985);
nand U5183 (N_5183,N_4909,N_4942);
nor U5184 (N_5184,N_4854,N_4884);
and U5185 (N_5185,N_4830,N_4978);
nand U5186 (N_5186,N_4825,N_4992);
or U5187 (N_5187,N_4900,N_4805);
or U5188 (N_5188,N_4885,N_4812);
and U5189 (N_5189,N_4809,N_4966);
xor U5190 (N_5190,N_4861,N_4811);
xor U5191 (N_5191,N_4808,N_4995);
and U5192 (N_5192,N_4978,N_4960);
or U5193 (N_5193,N_4994,N_4900);
and U5194 (N_5194,N_4982,N_4825);
or U5195 (N_5195,N_4868,N_4996);
xnor U5196 (N_5196,N_4864,N_4913);
or U5197 (N_5197,N_4823,N_4933);
nand U5198 (N_5198,N_4987,N_4881);
nor U5199 (N_5199,N_4861,N_4956);
and U5200 (N_5200,N_5121,N_5057);
and U5201 (N_5201,N_5117,N_5089);
or U5202 (N_5202,N_5036,N_5079);
nand U5203 (N_5203,N_5052,N_5120);
xnor U5204 (N_5204,N_5174,N_5014);
nand U5205 (N_5205,N_5069,N_5012);
nand U5206 (N_5206,N_5158,N_5171);
nor U5207 (N_5207,N_5104,N_5035);
nor U5208 (N_5208,N_5172,N_5097);
xnor U5209 (N_5209,N_5017,N_5094);
or U5210 (N_5210,N_5123,N_5063);
and U5211 (N_5211,N_5144,N_5165);
nand U5212 (N_5212,N_5160,N_5133);
xor U5213 (N_5213,N_5076,N_5066);
nor U5214 (N_5214,N_5000,N_5167);
nor U5215 (N_5215,N_5013,N_5003);
xor U5216 (N_5216,N_5010,N_5064);
or U5217 (N_5217,N_5053,N_5109);
xnor U5218 (N_5218,N_5149,N_5148);
nand U5219 (N_5219,N_5038,N_5159);
or U5220 (N_5220,N_5002,N_5033);
nor U5221 (N_5221,N_5018,N_5182);
and U5222 (N_5222,N_5152,N_5068);
or U5223 (N_5223,N_5001,N_5091);
and U5224 (N_5224,N_5138,N_5082);
nor U5225 (N_5225,N_5112,N_5118);
and U5226 (N_5226,N_5119,N_5029);
nand U5227 (N_5227,N_5045,N_5039);
nand U5228 (N_5228,N_5073,N_5176);
nor U5229 (N_5229,N_5188,N_5040);
xor U5230 (N_5230,N_5048,N_5187);
nor U5231 (N_5231,N_5043,N_5166);
or U5232 (N_5232,N_5026,N_5179);
or U5233 (N_5233,N_5080,N_5192);
and U5234 (N_5234,N_5044,N_5011);
and U5235 (N_5235,N_5086,N_5085);
or U5236 (N_5236,N_5190,N_5020);
and U5237 (N_5237,N_5074,N_5132);
or U5238 (N_5238,N_5071,N_5092);
or U5239 (N_5239,N_5024,N_5046);
and U5240 (N_5240,N_5164,N_5193);
or U5241 (N_5241,N_5126,N_5054);
and U5242 (N_5242,N_5183,N_5141);
nand U5243 (N_5243,N_5031,N_5191);
nand U5244 (N_5244,N_5198,N_5095);
nand U5245 (N_5245,N_5041,N_5116);
or U5246 (N_5246,N_5162,N_5108);
nor U5247 (N_5247,N_5090,N_5113);
xnor U5248 (N_5248,N_5047,N_5099);
nand U5249 (N_5249,N_5019,N_5096);
and U5250 (N_5250,N_5147,N_5065);
xor U5251 (N_5251,N_5131,N_5168);
and U5252 (N_5252,N_5125,N_5137);
and U5253 (N_5253,N_5084,N_5136);
nand U5254 (N_5254,N_5060,N_5197);
nor U5255 (N_5255,N_5122,N_5103);
and U5256 (N_5256,N_5111,N_5083);
xnor U5257 (N_5257,N_5184,N_5189);
nor U5258 (N_5258,N_5161,N_5185);
nor U5259 (N_5259,N_5127,N_5142);
or U5260 (N_5260,N_5087,N_5006);
xnor U5261 (N_5261,N_5173,N_5021);
or U5262 (N_5262,N_5051,N_5163);
nor U5263 (N_5263,N_5134,N_5107);
nand U5264 (N_5264,N_5081,N_5049);
nor U5265 (N_5265,N_5129,N_5151);
nor U5266 (N_5266,N_5030,N_5156);
nand U5267 (N_5267,N_5088,N_5032);
nor U5268 (N_5268,N_5143,N_5027);
and U5269 (N_5269,N_5135,N_5175);
nor U5270 (N_5270,N_5194,N_5196);
xnor U5271 (N_5271,N_5075,N_5004);
nand U5272 (N_5272,N_5056,N_5124);
nand U5273 (N_5273,N_5062,N_5145);
xnor U5274 (N_5274,N_5146,N_5110);
and U5275 (N_5275,N_5101,N_5115);
or U5276 (N_5276,N_5130,N_5177);
nor U5277 (N_5277,N_5169,N_5050);
or U5278 (N_5278,N_5180,N_5061);
nor U5279 (N_5279,N_5154,N_5022);
xor U5280 (N_5280,N_5195,N_5093);
nand U5281 (N_5281,N_5005,N_5015);
or U5282 (N_5282,N_5009,N_5058);
or U5283 (N_5283,N_5106,N_5028);
and U5284 (N_5284,N_5139,N_5037);
nor U5285 (N_5285,N_5181,N_5025);
xnor U5286 (N_5286,N_5023,N_5150);
xnor U5287 (N_5287,N_5128,N_5042);
and U5288 (N_5288,N_5034,N_5102);
nor U5289 (N_5289,N_5105,N_5100);
and U5290 (N_5290,N_5157,N_5008);
xor U5291 (N_5291,N_5072,N_5155);
nand U5292 (N_5292,N_5186,N_5070);
and U5293 (N_5293,N_5016,N_5140);
nand U5294 (N_5294,N_5007,N_5077);
nand U5295 (N_5295,N_5170,N_5153);
and U5296 (N_5296,N_5098,N_5199);
nand U5297 (N_5297,N_5059,N_5078);
or U5298 (N_5298,N_5055,N_5114);
and U5299 (N_5299,N_5067,N_5178);
or U5300 (N_5300,N_5103,N_5174);
and U5301 (N_5301,N_5186,N_5159);
or U5302 (N_5302,N_5090,N_5197);
and U5303 (N_5303,N_5164,N_5067);
nor U5304 (N_5304,N_5089,N_5112);
and U5305 (N_5305,N_5005,N_5147);
xnor U5306 (N_5306,N_5056,N_5134);
or U5307 (N_5307,N_5137,N_5017);
xor U5308 (N_5308,N_5046,N_5174);
xor U5309 (N_5309,N_5182,N_5199);
xor U5310 (N_5310,N_5041,N_5011);
nor U5311 (N_5311,N_5179,N_5102);
and U5312 (N_5312,N_5174,N_5022);
or U5313 (N_5313,N_5085,N_5068);
nand U5314 (N_5314,N_5134,N_5020);
or U5315 (N_5315,N_5089,N_5009);
and U5316 (N_5316,N_5051,N_5156);
or U5317 (N_5317,N_5181,N_5107);
and U5318 (N_5318,N_5185,N_5197);
xor U5319 (N_5319,N_5153,N_5161);
and U5320 (N_5320,N_5061,N_5108);
and U5321 (N_5321,N_5132,N_5003);
nand U5322 (N_5322,N_5052,N_5197);
xnor U5323 (N_5323,N_5110,N_5017);
nand U5324 (N_5324,N_5005,N_5152);
xnor U5325 (N_5325,N_5161,N_5087);
and U5326 (N_5326,N_5159,N_5139);
and U5327 (N_5327,N_5194,N_5039);
or U5328 (N_5328,N_5122,N_5121);
and U5329 (N_5329,N_5007,N_5084);
and U5330 (N_5330,N_5143,N_5051);
or U5331 (N_5331,N_5071,N_5024);
or U5332 (N_5332,N_5033,N_5059);
or U5333 (N_5333,N_5006,N_5160);
and U5334 (N_5334,N_5137,N_5104);
and U5335 (N_5335,N_5173,N_5075);
xnor U5336 (N_5336,N_5001,N_5173);
or U5337 (N_5337,N_5184,N_5170);
or U5338 (N_5338,N_5076,N_5089);
and U5339 (N_5339,N_5081,N_5064);
xnor U5340 (N_5340,N_5024,N_5155);
nor U5341 (N_5341,N_5129,N_5076);
and U5342 (N_5342,N_5072,N_5190);
xnor U5343 (N_5343,N_5085,N_5043);
and U5344 (N_5344,N_5155,N_5174);
or U5345 (N_5345,N_5171,N_5176);
xnor U5346 (N_5346,N_5001,N_5050);
nand U5347 (N_5347,N_5063,N_5196);
nor U5348 (N_5348,N_5182,N_5185);
or U5349 (N_5349,N_5052,N_5179);
nor U5350 (N_5350,N_5009,N_5103);
nand U5351 (N_5351,N_5119,N_5068);
or U5352 (N_5352,N_5104,N_5011);
nor U5353 (N_5353,N_5053,N_5170);
nand U5354 (N_5354,N_5194,N_5089);
nor U5355 (N_5355,N_5063,N_5014);
xor U5356 (N_5356,N_5047,N_5153);
xnor U5357 (N_5357,N_5055,N_5150);
and U5358 (N_5358,N_5134,N_5042);
xnor U5359 (N_5359,N_5143,N_5124);
nor U5360 (N_5360,N_5071,N_5097);
xor U5361 (N_5361,N_5036,N_5097);
xor U5362 (N_5362,N_5138,N_5149);
or U5363 (N_5363,N_5114,N_5133);
xor U5364 (N_5364,N_5094,N_5045);
nand U5365 (N_5365,N_5155,N_5016);
nand U5366 (N_5366,N_5020,N_5040);
or U5367 (N_5367,N_5180,N_5002);
and U5368 (N_5368,N_5193,N_5032);
and U5369 (N_5369,N_5148,N_5167);
and U5370 (N_5370,N_5000,N_5142);
xnor U5371 (N_5371,N_5042,N_5187);
or U5372 (N_5372,N_5199,N_5118);
nand U5373 (N_5373,N_5022,N_5168);
and U5374 (N_5374,N_5039,N_5043);
nor U5375 (N_5375,N_5175,N_5100);
nand U5376 (N_5376,N_5136,N_5021);
nor U5377 (N_5377,N_5170,N_5174);
or U5378 (N_5378,N_5118,N_5012);
xnor U5379 (N_5379,N_5035,N_5016);
and U5380 (N_5380,N_5031,N_5179);
nor U5381 (N_5381,N_5164,N_5101);
nor U5382 (N_5382,N_5053,N_5134);
xor U5383 (N_5383,N_5045,N_5130);
xor U5384 (N_5384,N_5092,N_5187);
or U5385 (N_5385,N_5017,N_5000);
nor U5386 (N_5386,N_5037,N_5133);
nand U5387 (N_5387,N_5181,N_5089);
nand U5388 (N_5388,N_5039,N_5164);
and U5389 (N_5389,N_5100,N_5189);
or U5390 (N_5390,N_5171,N_5073);
nand U5391 (N_5391,N_5156,N_5044);
nor U5392 (N_5392,N_5166,N_5134);
xnor U5393 (N_5393,N_5176,N_5001);
xnor U5394 (N_5394,N_5106,N_5053);
xnor U5395 (N_5395,N_5027,N_5022);
xnor U5396 (N_5396,N_5116,N_5119);
nor U5397 (N_5397,N_5134,N_5175);
xnor U5398 (N_5398,N_5024,N_5030);
and U5399 (N_5399,N_5099,N_5154);
and U5400 (N_5400,N_5345,N_5387);
nor U5401 (N_5401,N_5307,N_5324);
or U5402 (N_5402,N_5241,N_5247);
nand U5403 (N_5403,N_5254,N_5310);
or U5404 (N_5404,N_5383,N_5312);
and U5405 (N_5405,N_5202,N_5371);
nand U5406 (N_5406,N_5344,N_5259);
nor U5407 (N_5407,N_5349,N_5331);
nor U5408 (N_5408,N_5242,N_5299);
nand U5409 (N_5409,N_5365,N_5257);
xor U5410 (N_5410,N_5201,N_5263);
or U5411 (N_5411,N_5360,N_5226);
nand U5412 (N_5412,N_5322,N_5253);
and U5413 (N_5413,N_5320,N_5295);
nand U5414 (N_5414,N_5222,N_5316);
nand U5415 (N_5415,N_5231,N_5352);
and U5416 (N_5416,N_5279,N_5364);
and U5417 (N_5417,N_5298,N_5378);
xor U5418 (N_5418,N_5338,N_5300);
or U5419 (N_5419,N_5292,N_5392);
nor U5420 (N_5420,N_5379,N_5200);
or U5421 (N_5421,N_5272,N_5373);
or U5422 (N_5422,N_5280,N_5369);
or U5423 (N_5423,N_5216,N_5311);
xor U5424 (N_5424,N_5240,N_5225);
nand U5425 (N_5425,N_5335,N_5206);
nor U5426 (N_5426,N_5207,N_5395);
or U5427 (N_5427,N_5326,N_5277);
nor U5428 (N_5428,N_5313,N_5288);
or U5429 (N_5429,N_5382,N_5346);
xor U5430 (N_5430,N_5212,N_5256);
nor U5431 (N_5431,N_5397,N_5325);
xnor U5432 (N_5432,N_5381,N_5329);
xor U5433 (N_5433,N_5367,N_5319);
nand U5434 (N_5434,N_5223,N_5374);
and U5435 (N_5435,N_5293,N_5362);
or U5436 (N_5436,N_5215,N_5399);
xnor U5437 (N_5437,N_5332,N_5281);
nand U5438 (N_5438,N_5353,N_5328);
nor U5439 (N_5439,N_5237,N_5363);
or U5440 (N_5440,N_5270,N_5219);
or U5441 (N_5441,N_5283,N_5239);
and U5442 (N_5442,N_5230,N_5385);
nor U5443 (N_5443,N_5214,N_5296);
xor U5444 (N_5444,N_5209,N_5236);
nor U5445 (N_5445,N_5389,N_5302);
or U5446 (N_5446,N_5267,N_5251);
or U5447 (N_5447,N_5341,N_5258);
nor U5448 (N_5448,N_5261,N_5252);
nand U5449 (N_5449,N_5356,N_5264);
and U5450 (N_5450,N_5334,N_5327);
or U5451 (N_5451,N_5249,N_5229);
or U5452 (N_5452,N_5211,N_5210);
nand U5453 (N_5453,N_5351,N_5318);
xor U5454 (N_5454,N_5217,N_5243);
or U5455 (N_5455,N_5330,N_5282);
xor U5456 (N_5456,N_5358,N_5278);
and U5457 (N_5457,N_5244,N_5317);
nand U5458 (N_5458,N_5393,N_5386);
nor U5459 (N_5459,N_5359,N_5245);
nor U5460 (N_5460,N_5314,N_5275);
xor U5461 (N_5461,N_5366,N_5290);
nor U5462 (N_5462,N_5342,N_5355);
xnor U5463 (N_5463,N_5232,N_5213);
and U5464 (N_5464,N_5372,N_5390);
or U5465 (N_5465,N_5291,N_5269);
or U5466 (N_5466,N_5233,N_5321);
or U5467 (N_5467,N_5304,N_5250);
xor U5468 (N_5468,N_5333,N_5361);
nand U5469 (N_5469,N_5271,N_5340);
nand U5470 (N_5470,N_5375,N_5274);
and U5471 (N_5471,N_5376,N_5357);
nor U5472 (N_5472,N_5203,N_5266);
xor U5473 (N_5473,N_5221,N_5323);
nor U5474 (N_5474,N_5396,N_5308);
xor U5475 (N_5475,N_5370,N_5246);
xnor U5476 (N_5476,N_5208,N_5220);
xor U5477 (N_5477,N_5368,N_5384);
nand U5478 (N_5478,N_5227,N_5204);
xor U5479 (N_5479,N_5394,N_5306);
nand U5480 (N_5480,N_5248,N_5380);
or U5481 (N_5481,N_5268,N_5294);
and U5482 (N_5482,N_5315,N_5309);
xnor U5483 (N_5483,N_5289,N_5285);
xor U5484 (N_5484,N_5343,N_5297);
xnor U5485 (N_5485,N_5305,N_5228);
nand U5486 (N_5486,N_5377,N_5339);
and U5487 (N_5487,N_5336,N_5234);
xnor U5488 (N_5488,N_5337,N_5265);
nor U5489 (N_5489,N_5354,N_5255);
nor U5490 (N_5490,N_5218,N_5301);
xnor U5491 (N_5491,N_5238,N_5347);
or U5492 (N_5492,N_5348,N_5287);
and U5493 (N_5493,N_5391,N_5205);
xnor U5494 (N_5494,N_5260,N_5224);
nor U5495 (N_5495,N_5235,N_5262);
nor U5496 (N_5496,N_5284,N_5350);
xnor U5497 (N_5497,N_5388,N_5273);
nor U5498 (N_5498,N_5398,N_5286);
and U5499 (N_5499,N_5303,N_5276);
nor U5500 (N_5500,N_5297,N_5313);
nand U5501 (N_5501,N_5278,N_5292);
xnor U5502 (N_5502,N_5323,N_5207);
and U5503 (N_5503,N_5278,N_5213);
xor U5504 (N_5504,N_5273,N_5256);
or U5505 (N_5505,N_5279,N_5220);
or U5506 (N_5506,N_5249,N_5210);
nand U5507 (N_5507,N_5243,N_5345);
nor U5508 (N_5508,N_5378,N_5303);
nor U5509 (N_5509,N_5201,N_5235);
xnor U5510 (N_5510,N_5270,N_5271);
nor U5511 (N_5511,N_5283,N_5207);
and U5512 (N_5512,N_5218,N_5398);
or U5513 (N_5513,N_5384,N_5202);
and U5514 (N_5514,N_5313,N_5382);
or U5515 (N_5515,N_5290,N_5236);
nand U5516 (N_5516,N_5288,N_5233);
nand U5517 (N_5517,N_5366,N_5389);
xnor U5518 (N_5518,N_5381,N_5318);
and U5519 (N_5519,N_5285,N_5266);
and U5520 (N_5520,N_5316,N_5233);
and U5521 (N_5521,N_5238,N_5372);
nor U5522 (N_5522,N_5332,N_5381);
and U5523 (N_5523,N_5268,N_5329);
or U5524 (N_5524,N_5384,N_5399);
nand U5525 (N_5525,N_5300,N_5262);
and U5526 (N_5526,N_5389,N_5322);
and U5527 (N_5527,N_5350,N_5253);
or U5528 (N_5528,N_5200,N_5314);
or U5529 (N_5529,N_5360,N_5346);
nor U5530 (N_5530,N_5334,N_5382);
and U5531 (N_5531,N_5371,N_5229);
or U5532 (N_5532,N_5374,N_5285);
xor U5533 (N_5533,N_5344,N_5339);
and U5534 (N_5534,N_5261,N_5272);
and U5535 (N_5535,N_5352,N_5333);
and U5536 (N_5536,N_5209,N_5370);
xor U5537 (N_5537,N_5301,N_5257);
xnor U5538 (N_5538,N_5299,N_5225);
or U5539 (N_5539,N_5277,N_5255);
nand U5540 (N_5540,N_5221,N_5364);
and U5541 (N_5541,N_5305,N_5318);
or U5542 (N_5542,N_5342,N_5294);
or U5543 (N_5543,N_5281,N_5316);
or U5544 (N_5544,N_5284,N_5263);
xor U5545 (N_5545,N_5295,N_5312);
or U5546 (N_5546,N_5292,N_5334);
xnor U5547 (N_5547,N_5215,N_5354);
and U5548 (N_5548,N_5394,N_5324);
nand U5549 (N_5549,N_5229,N_5268);
xor U5550 (N_5550,N_5279,N_5222);
xor U5551 (N_5551,N_5375,N_5290);
or U5552 (N_5552,N_5281,N_5358);
nand U5553 (N_5553,N_5358,N_5234);
and U5554 (N_5554,N_5282,N_5306);
and U5555 (N_5555,N_5336,N_5370);
or U5556 (N_5556,N_5344,N_5388);
nand U5557 (N_5557,N_5371,N_5215);
nand U5558 (N_5558,N_5263,N_5289);
nand U5559 (N_5559,N_5397,N_5248);
xnor U5560 (N_5560,N_5239,N_5369);
xor U5561 (N_5561,N_5216,N_5233);
and U5562 (N_5562,N_5387,N_5277);
or U5563 (N_5563,N_5296,N_5248);
xnor U5564 (N_5564,N_5299,N_5219);
nand U5565 (N_5565,N_5367,N_5304);
nor U5566 (N_5566,N_5373,N_5251);
xor U5567 (N_5567,N_5334,N_5343);
and U5568 (N_5568,N_5216,N_5265);
and U5569 (N_5569,N_5273,N_5210);
nand U5570 (N_5570,N_5367,N_5323);
or U5571 (N_5571,N_5326,N_5293);
and U5572 (N_5572,N_5297,N_5312);
nand U5573 (N_5573,N_5346,N_5388);
nand U5574 (N_5574,N_5218,N_5340);
and U5575 (N_5575,N_5396,N_5254);
nand U5576 (N_5576,N_5324,N_5378);
xnor U5577 (N_5577,N_5250,N_5342);
and U5578 (N_5578,N_5314,N_5396);
and U5579 (N_5579,N_5295,N_5211);
xor U5580 (N_5580,N_5376,N_5346);
nor U5581 (N_5581,N_5242,N_5384);
xor U5582 (N_5582,N_5297,N_5296);
and U5583 (N_5583,N_5203,N_5248);
nand U5584 (N_5584,N_5329,N_5337);
nor U5585 (N_5585,N_5355,N_5357);
nor U5586 (N_5586,N_5371,N_5230);
or U5587 (N_5587,N_5383,N_5381);
xor U5588 (N_5588,N_5247,N_5254);
or U5589 (N_5589,N_5319,N_5343);
xor U5590 (N_5590,N_5269,N_5354);
or U5591 (N_5591,N_5370,N_5328);
nor U5592 (N_5592,N_5374,N_5373);
and U5593 (N_5593,N_5219,N_5391);
or U5594 (N_5594,N_5261,N_5330);
xor U5595 (N_5595,N_5386,N_5330);
or U5596 (N_5596,N_5289,N_5375);
xor U5597 (N_5597,N_5358,N_5375);
and U5598 (N_5598,N_5319,N_5355);
or U5599 (N_5599,N_5393,N_5347);
nand U5600 (N_5600,N_5569,N_5448);
nand U5601 (N_5601,N_5593,N_5451);
xor U5602 (N_5602,N_5468,N_5463);
nand U5603 (N_5603,N_5425,N_5411);
xnor U5604 (N_5604,N_5464,N_5502);
and U5605 (N_5605,N_5592,N_5548);
and U5606 (N_5606,N_5554,N_5429);
xnor U5607 (N_5607,N_5493,N_5573);
nor U5608 (N_5608,N_5431,N_5599);
xnor U5609 (N_5609,N_5405,N_5585);
and U5610 (N_5610,N_5562,N_5506);
and U5611 (N_5611,N_5420,N_5469);
nor U5612 (N_5612,N_5514,N_5461);
nand U5613 (N_5613,N_5535,N_5570);
xor U5614 (N_5614,N_5483,N_5576);
xor U5615 (N_5615,N_5565,N_5440);
xnor U5616 (N_5616,N_5523,N_5516);
or U5617 (N_5617,N_5471,N_5433);
or U5618 (N_5618,N_5567,N_5503);
nand U5619 (N_5619,N_5434,N_5481);
or U5620 (N_5620,N_5494,N_5445);
nor U5621 (N_5621,N_5563,N_5582);
nand U5622 (N_5622,N_5515,N_5487);
nand U5623 (N_5623,N_5595,N_5438);
or U5624 (N_5624,N_5552,N_5476);
nor U5625 (N_5625,N_5591,N_5534);
nand U5626 (N_5626,N_5526,N_5550);
nor U5627 (N_5627,N_5501,N_5581);
nand U5628 (N_5628,N_5512,N_5557);
or U5629 (N_5629,N_5568,N_5407);
or U5630 (N_5630,N_5524,N_5492);
or U5631 (N_5631,N_5456,N_5488);
xnor U5632 (N_5632,N_5478,N_5466);
xnor U5633 (N_5633,N_5482,N_5453);
nor U5634 (N_5634,N_5528,N_5589);
nand U5635 (N_5635,N_5426,N_5556);
or U5636 (N_5636,N_5546,N_5491);
or U5637 (N_5637,N_5537,N_5467);
nor U5638 (N_5638,N_5419,N_5564);
nor U5639 (N_5639,N_5490,N_5413);
xor U5640 (N_5640,N_5495,N_5480);
nor U5641 (N_5641,N_5415,N_5455);
and U5642 (N_5642,N_5549,N_5509);
and U5643 (N_5643,N_5470,N_5561);
and U5644 (N_5644,N_5500,N_5409);
xor U5645 (N_5645,N_5566,N_5498);
or U5646 (N_5646,N_5408,N_5541);
nand U5647 (N_5647,N_5532,N_5410);
or U5648 (N_5648,N_5544,N_5439);
or U5649 (N_5649,N_5450,N_5530);
nand U5650 (N_5650,N_5597,N_5449);
nor U5651 (N_5651,N_5477,N_5437);
nand U5652 (N_5652,N_5525,N_5527);
and U5653 (N_5653,N_5584,N_5558);
xor U5654 (N_5654,N_5596,N_5533);
or U5655 (N_5655,N_5517,N_5522);
nand U5656 (N_5656,N_5594,N_5519);
or U5657 (N_5657,N_5575,N_5578);
nor U5658 (N_5658,N_5472,N_5432);
or U5659 (N_5659,N_5574,N_5587);
xor U5660 (N_5660,N_5430,N_5580);
and U5661 (N_5661,N_5436,N_5401);
or U5662 (N_5662,N_5560,N_5559);
and U5663 (N_5663,N_5486,N_5442);
or U5664 (N_5664,N_5414,N_5518);
and U5665 (N_5665,N_5520,N_5507);
or U5666 (N_5666,N_5427,N_5499);
xor U5667 (N_5667,N_5402,N_5435);
and U5668 (N_5668,N_5540,N_5510);
and U5669 (N_5669,N_5571,N_5475);
nor U5670 (N_5670,N_5479,N_5497);
xnor U5671 (N_5671,N_5484,N_5416);
or U5672 (N_5672,N_5577,N_5441);
nand U5673 (N_5673,N_5536,N_5588);
nor U5674 (N_5674,N_5531,N_5572);
or U5675 (N_5675,N_5454,N_5446);
xnor U5676 (N_5676,N_5598,N_5418);
or U5677 (N_5677,N_5457,N_5508);
nand U5678 (N_5678,N_5542,N_5547);
nand U5679 (N_5679,N_5422,N_5529);
or U5680 (N_5680,N_5538,N_5404);
or U5681 (N_5681,N_5590,N_5424);
and U5682 (N_5682,N_5504,N_5474);
and U5683 (N_5683,N_5417,N_5452);
nor U5684 (N_5684,N_5459,N_5489);
and U5685 (N_5685,N_5473,N_5539);
and U5686 (N_5686,N_5586,N_5513);
and U5687 (N_5687,N_5447,N_5428);
xnor U5688 (N_5688,N_5412,N_5444);
and U5689 (N_5689,N_5458,N_5583);
nand U5690 (N_5690,N_5579,N_5543);
xor U5691 (N_5691,N_5545,N_5551);
xor U5692 (N_5692,N_5553,N_5421);
and U5693 (N_5693,N_5403,N_5462);
or U5694 (N_5694,N_5505,N_5496);
nand U5695 (N_5695,N_5521,N_5400);
nor U5696 (N_5696,N_5485,N_5460);
nor U5697 (N_5697,N_5406,N_5423);
xnor U5698 (N_5698,N_5443,N_5555);
nor U5699 (N_5699,N_5465,N_5511);
nor U5700 (N_5700,N_5598,N_5408);
nand U5701 (N_5701,N_5497,N_5449);
and U5702 (N_5702,N_5589,N_5587);
xor U5703 (N_5703,N_5521,N_5499);
or U5704 (N_5704,N_5457,N_5445);
nor U5705 (N_5705,N_5508,N_5435);
and U5706 (N_5706,N_5468,N_5590);
or U5707 (N_5707,N_5470,N_5531);
and U5708 (N_5708,N_5434,N_5452);
nor U5709 (N_5709,N_5451,N_5484);
xnor U5710 (N_5710,N_5565,N_5496);
nor U5711 (N_5711,N_5597,N_5413);
nor U5712 (N_5712,N_5587,N_5575);
or U5713 (N_5713,N_5402,N_5411);
xnor U5714 (N_5714,N_5422,N_5456);
and U5715 (N_5715,N_5416,N_5528);
nand U5716 (N_5716,N_5584,N_5565);
nor U5717 (N_5717,N_5591,N_5405);
xor U5718 (N_5718,N_5460,N_5406);
or U5719 (N_5719,N_5490,N_5445);
and U5720 (N_5720,N_5505,N_5425);
or U5721 (N_5721,N_5410,N_5486);
or U5722 (N_5722,N_5488,N_5513);
and U5723 (N_5723,N_5568,N_5519);
nor U5724 (N_5724,N_5434,N_5503);
and U5725 (N_5725,N_5591,N_5555);
nor U5726 (N_5726,N_5456,N_5583);
nor U5727 (N_5727,N_5421,N_5432);
nor U5728 (N_5728,N_5515,N_5503);
xor U5729 (N_5729,N_5436,N_5451);
xnor U5730 (N_5730,N_5432,N_5599);
xnor U5731 (N_5731,N_5507,N_5430);
xor U5732 (N_5732,N_5418,N_5457);
nand U5733 (N_5733,N_5403,N_5416);
nand U5734 (N_5734,N_5487,N_5522);
or U5735 (N_5735,N_5590,N_5531);
nor U5736 (N_5736,N_5476,N_5517);
nand U5737 (N_5737,N_5510,N_5538);
or U5738 (N_5738,N_5519,N_5585);
xnor U5739 (N_5739,N_5576,N_5455);
and U5740 (N_5740,N_5410,N_5495);
and U5741 (N_5741,N_5595,N_5523);
or U5742 (N_5742,N_5466,N_5425);
nor U5743 (N_5743,N_5409,N_5467);
nand U5744 (N_5744,N_5411,N_5527);
xor U5745 (N_5745,N_5452,N_5557);
and U5746 (N_5746,N_5457,N_5494);
nor U5747 (N_5747,N_5591,N_5402);
nand U5748 (N_5748,N_5565,N_5572);
nor U5749 (N_5749,N_5457,N_5554);
xnor U5750 (N_5750,N_5556,N_5510);
or U5751 (N_5751,N_5459,N_5433);
xnor U5752 (N_5752,N_5417,N_5557);
or U5753 (N_5753,N_5557,N_5550);
xor U5754 (N_5754,N_5533,N_5463);
nand U5755 (N_5755,N_5486,N_5589);
xnor U5756 (N_5756,N_5469,N_5463);
or U5757 (N_5757,N_5569,N_5490);
nand U5758 (N_5758,N_5427,N_5560);
nand U5759 (N_5759,N_5439,N_5443);
nand U5760 (N_5760,N_5594,N_5582);
nor U5761 (N_5761,N_5457,N_5597);
nand U5762 (N_5762,N_5482,N_5489);
and U5763 (N_5763,N_5426,N_5416);
nor U5764 (N_5764,N_5444,N_5464);
xor U5765 (N_5765,N_5552,N_5570);
or U5766 (N_5766,N_5480,N_5404);
and U5767 (N_5767,N_5562,N_5593);
xnor U5768 (N_5768,N_5459,N_5527);
and U5769 (N_5769,N_5414,N_5413);
or U5770 (N_5770,N_5585,N_5471);
nor U5771 (N_5771,N_5452,N_5545);
or U5772 (N_5772,N_5501,N_5437);
or U5773 (N_5773,N_5569,N_5562);
nor U5774 (N_5774,N_5594,N_5474);
or U5775 (N_5775,N_5422,N_5583);
and U5776 (N_5776,N_5545,N_5460);
and U5777 (N_5777,N_5588,N_5534);
nor U5778 (N_5778,N_5501,N_5489);
nand U5779 (N_5779,N_5428,N_5437);
nor U5780 (N_5780,N_5597,N_5431);
or U5781 (N_5781,N_5482,N_5518);
nor U5782 (N_5782,N_5450,N_5582);
nor U5783 (N_5783,N_5472,N_5483);
or U5784 (N_5784,N_5440,N_5413);
and U5785 (N_5785,N_5599,N_5519);
nand U5786 (N_5786,N_5570,N_5575);
or U5787 (N_5787,N_5562,N_5411);
xnor U5788 (N_5788,N_5565,N_5413);
nor U5789 (N_5789,N_5400,N_5481);
or U5790 (N_5790,N_5591,N_5511);
nand U5791 (N_5791,N_5592,N_5439);
and U5792 (N_5792,N_5500,N_5517);
nand U5793 (N_5793,N_5487,N_5557);
or U5794 (N_5794,N_5563,N_5578);
nor U5795 (N_5795,N_5417,N_5599);
nand U5796 (N_5796,N_5455,N_5408);
and U5797 (N_5797,N_5491,N_5571);
nor U5798 (N_5798,N_5466,N_5460);
or U5799 (N_5799,N_5505,N_5401);
or U5800 (N_5800,N_5625,N_5791);
nand U5801 (N_5801,N_5748,N_5696);
nand U5802 (N_5802,N_5669,N_5759);
xor U5803 (N_5803,N_5666,N_5652);
nand U5804 (N_5804,N_5660,N_5747);
nor U5805 (N_5805,N_5796,N_5776);
or U5806 (N_5806,N_5603,N_5657);
nor U5807 (N_5807,N_5771,N_5644);
nor U5808 (N_5808,N_5631,N_5690);
or U5809 (N_5809,N_5600,N_5757);
nor U5810 (N_5810,N_5694,N_5756);
and U5811 (N_5811,N_5650,N_5686);
nor U5812 (N_5812,N_5676,N_5613);
or U5813 (N_5813,N_5705,N_5674);
or U5814 (N_5814,N_5645,N_5717);
nor U5815 (N_5815,N_5668,N_5628);
xor U5816 (N_5816,N_5708,N_5607);
nor U5817 (N_5817,N_5742,N_5688);
and U5818 (N_5818,N_5699,N_5678);
xnor U5819 (N_5819,N_5719,N_5712);
nor U5820 (N_5820,N_5639,N_5627);
xnor U5821 (N_5821,N_5697,N_5663);
and U5822 (N_5822,N_5745,N_5715);
nand U5823 (N_5823,N_5623,N_5703);
and U5824 (N_5824,N_5762,N_5718);
or U5825 (N_5825,N_5685,N_5615);
and U5826 (N_5826,N_5659,N_5637);
nand U5827 (N_5827,N_5610,N_5729);
xnor U5828 (N_5828,N_5734,N_5721);
nand U5829 (N_5829,N_5709,N_5790);
nor U5830 (N_5830,N_5682,N_5723);
nor U5831 (N_5831,N_5653,N_5784);
xor U5832 (N_5832,N_5716,N_5750);
nand U5833 (N_5833,N_5728,N_5642);
and U5834 (N_5834,N_5722,N_5604);
nor U5835 (N_5835,N_5638,N_5741);
and U5836 (N_5836,N_5780,N_5793);
xnor U5837 (N_5837,N_5763,N_5661);
and U5838 (N_5838,N_5778,N_5664);
nand U5839 (N_5839,N_5612,N_5755);
nand U5840 (N_5840,N_5680,N_5693);
xnor U5841 (N_5841,N_5622,N_5772);
xor U5842 (N_5842,N_5632,N_5629);
nand U5843 (N_5843,N_5633,N_5683);
xor U5844 (N_5844,N_5770,N_5797);
nor U5845 (N_5845,N_5601,N_5752);
nor U5846 (N_5846,N_5635,N_5731);
nand U5847 (N_5847,N_5704,N_5630);
or U5848 (N_5848,N_5798,N_5611);
nor U5849 (N_5849,N_5651,N_5617);
and U5850 (N_5850,N_5605,N_5788);
xor U5851 (N_5851,N_5746,N_5673);
nor U5852 (N_5852,N_5667,N_5769);
nor U5853 (N_5853,N_5754,N_5794);
or U5854 (N_5854,N_5781,N_5691);
nor U5855 (N_5855,N_5765,N_5649);
xor U5856 (N_5856,N_5737,N_5736);
or U5857 (N_5857,N_5618,N_5783);
or U5858 (N_5858,N_5626,N_5760);
or U5859 (N_5859,N_5753,N_5743);
and U5860 (N_5860,N_5656,N_5725);
and U5861 (N_5861,N_5738,N_5641);
or U5862 (N_5862,N_5616,N_5710);
xnor U5863 (N_5863,N_5662,N_5679);
nor U5864 (N_5864,N_5799,N_5782);
and U5865 (N_5865,N_5672,N_5675);
xnor U5866 (N_5866,N_5711,N_5789);
nor U5867 (N_5867,N_5634,N_5749);
nand U5868 (N_5868,N_5740,N_5609);
and U5869 (N_5869,N_5692,N_5640);
and U5870 (N_5870,N_5695,N_5665);
xor U5871 (N_5871,N_5785,N_5655);
and U5872 (N_5872,N_5726,N_5687);
xnor U5873 (N_5873,N_5621,N_5773);
nand U5874 (N_5874,N_5764,N_5670);
and U5875 (N_5875,N_5608,N_5646);
nand U5876 (N_5876,N_5766,N_5767);
or U5877 (N_5877,N_5702,N_5671);
nand U5878 (N_5878,N_5751,N_5698);
nand U5879 (N_5879,N_5720,N_5624);
nor U5880 (N_5880,N_5602,N_5744);
nor U5881 (N_5881,N_5654,N_5606);
nand U5882 (N_5882,N_5619,N_5707);
or U5883 (N_5883,N_5643,N_5792);
nand U5884 (N_5884,N_5787,N_5701);
nor U5885 (N_5885,N_5735,N_5758);
or U5886 (N_5886,N_5779,N_5714);
and U5887 (N_5887,N_5647,N_5786);
xnor U5888 (N_5888,N_5636,N_5620);
xnor U5889 (N_5889,N_5768,N_5658);
or U5890 (N_5890,N_5684,N_5732);
xor U5891 (N_5891,N_5677,N_5724);
and U5892 (N_5892,N_5774,N_5700);
and U5893 (N_5893,N_5795,N_5761);
xnor U5894 (N_5894,N_5689,N_5713);
xnor U5895 (N_5895,N_5739,N_5727);
or U5896 (N_5896,N_5775,N_5648);
and U5897 (N_5897,N_5614,N_5730);
or U5898 (N_5898,N_5706,N_5777);
or U5899 (N_5899,N_5733,N_5681);
xor U5900 (N_5900,N_5790,N_5641);
nor U5901 (N_5901,N_5627,N_5601);
xnor U5902 (N_5902,N_5693,N_5672);
nor U5903 (N_5903,N_5752,N_5714);
nor U5904 (N_5904,N_5609,N_5793);
nand U5905 (N_5905,N_5656,N_5613);
or U5906 (N_5906,N_5630,N_5786);
nand U5907 (N_5907,N_5702,N_5716);
nor U5908 (N_5908,N_5622,N_5615);
nor U5909 (N_5909,N_5712,N_5742);
or U5910 (N_5910,N_5754,N_5763);
nand U5911 (N_5911,N_5649,N_5664);
xnor U5912 (N_5912,N_5759,N_5785);
xor U5913 (N_5913,N_5783,N_5687);
or U5914 (N_5914,N_5658,N_5714);
nor U5915 (N_5915,N_5615,N_5652);
nand U5916 (N_5916,N_5632,N_5714);
and U5917 (N_5917,N_5673,N_5764);
xnor U5918 (N_5918,N_5773,N_5625);
xor U5919 (N_5919,N_5746,N_5616);
and U5920 (N_5920,N_5785,N_5776);
and U5921 (N_5921,N_5600,N_5789);
and U5922 (N_5922,N_5672,N_5794);
or U5923 (N_5923,N_5614,N_5727);
nor U5924 (N_5924,N_5627,N_5613);
or U5925 (N_5925,N_5617,N_5742);
or U5926 (N_5926,N_5731,N_5652);
nor U5927 (N_5927,N_5616,N_5663);
nand U5928 (N_5928,N_5679,N_5758);
nor U5929 (N_5929,N_5697,N_5687);
nand U5930 (N_5930,N_5794,N_5659);
and U5931 (N_5931,N_5658,N_5759);
and U5932 (N_5932,N_5631,N_5788);
nand U5933 (N_5933,N_5751,N_5776);
nand U5934 (N_5934,N_5652,N_5655);
and U5935 (N_5935,N_5754,N_5652);
nor U5936 (N_5936,N_5780,N_5738);
nand U5937 (N_5937,N_5714,N_5789);
or U5938 (N_5938,N_5631,N_5628);
xor U5939 (N_5939,N_5631,N_5771);
and U5940 (N_5940,N_5602,N_5673);
xnor U5941 (N_5941,N_5634,N_5748);
or U5942 (N_5942,N_5619,N_5608);
nor U5943 (N_5943,N_5688,N_5730);
xor U5944 (N_5944,N_5685,N_5676);
xnor U5945 (N_5945,N_5674,N_5794);
and U5946 (N_5946,N_5785,N_5659);
nand U5947 (N_5947,N_5648,N_5728);
and U5948 (N_5948,N_5716,N_5754);
xnor U5949 (N_5949,N_5798,N_5651);
nor U5950 (N_5950,N_5656,N_5658);
nand U5951 (N_5951,N_5795,N_5727);
xor U5952 (N_5952,N_5764,N_5787);
nor U5953 (N_5953,N_5787,N_5674);
xnor U5954 (N_5954,N_5662,N_5794);
xnor U5955 (N_5955,N_5604,N_5688);
nor U5956 (N_5956,N_5767,N_5737);
nor U5957 (N_5957,N_5659,N_5662);
nand U5958 (N_5958,N_5634,N_5656);
and U5959 (N_5959,N_5680,N_5603);
and U5960 (N_5960,N_5776,N_5610);
xnor U5961 (N_5961,N_5682,N_5643);
xor U5962 (N_5962,N_5779,N_5610);
or U5963 (N_5963,N_5742,N_5725);
and U5964 (N_5964,N_5617,N_5787);
nand U5965 (N_5965,N_5785,N_5765);
xnor U5966 (N_5966,N_5791,N_5718);
and U5967 (N_5967,N_5615,N_5654);
xnor U5968 (N_5968,N_5761,N_5679);
xor U5969 (N_5969,N_5792,N_5681);
and U5970 (N_5970,N_5637,N_5670);
or U5971 (N_5971,N_5646,N_5654);
or U5972 (N_5972,N_5626,N_5726);
and U5973 (N_5973,N_5796,N_5742);
nand U5974 (N_5974,N_5698,N_5766);
xor U5975 (N_5975,N_5626,N_5649);
or U5976 (N_5976,N_5699,N_5626);
nand U5977 (N_5977,N_5743,N_5781);
and U5978 (N_5978,N_5747,N_5633);
xor U5979 (N_5979,N_5685,N_5629);
nand U5980 (N_5980,N_5626,N_5713);
nand U5981 (N_5981,N_5797,N_5690);
nor U5982 (N_5982,N_5634,N_5693);
nand U5983 (N_5983,N_5683,N_5636);
xor U5984 (N_5984,N_5620,N_5767);
nor U5985 (N_5985,N_5630,N_5763);
and U5986 (N_5986,N_5638,N_5641);
nand U5987 (N_5987,N_5791,N_5774);
or U5988 (N_5988,N_5753,N_5710);
or U5989 (N_5989,N_5683,N_5743);
xnor U5990 (N_5990,N_5708,N_5642);
and U5991 (N_5991,N_5795,N_5768);
nor U5992 (N_5992,N_5731,N_5615);
nor U5993 (N_5993,N_5728,N_5620);
nor U5994 (N_5994,N_5792,N_5646);
nor U5995 (N_5995,N_5791,N_5762);
or U5996 (N_5996,N_5686,N_5784);
or U5997 (N_5997,N_5602,N_5708);
xnor U5998 (N_5998,N_5785,N_5700);
nand U5999 (N_5999,N_5747,N_5755);
and U6000 (N_6000,N_5977,N_5892);
nor U6001 (N_6001,N_5939,N_5959);
xor U6002 (N_6002,N_5981,N_5813);
nor U6003 (N_6003,N_5951,N_5874);
and U6004 (N_6004,N_5801,N_5960);
and U6005 (N_6005,N_5965,N_5912);
nand U6006 (N_6006,N_5873,N_5923);
xor U6007 (N_6007,N_5887,N_5896);
nand U6008 (N_6008,N_5839,N_5867);
nor U6009 (N_6009,N_5847,N_5921);
and U6010 (N_6010,N_5995,N_5868);
nand U6011 (N_6011,N_5953,N_5930);
and U6012 (N_6012,N_5831,N_5902);
nand U6013 (N_6013,N_5865,N_5856);
and U6014 (N_6014,N_5889,N_5956);
and U6015 (N_6015,N_5904,N_5980);
xor U6016 (N_6016,N_5840,N_5970);
and U6017 (N_6017,N_5944,N_5881);
or U6018 (N_6018,N_5973,N_5994);
xnor U6019 (N_6019,N_5803,N_5907);
nor U6020 (N_6020,N_5999,N_5946);
nor U6021 (N_6021,N_5911,N_5835);
nor U6022 (N_6022,N_5807,N_5945);
or U6023 (N_6023,N_5919,N_5816);
xor U6024 (N_6024,N_5957,N_5824);
xnor U6025 (N_6025,N_5858,N_5998);
or U6026 (N_6026,N_5948,N_5933);
or U6027 (N_6027,N_5844,N_5810);
xnor U6028 (N_6028,N_5978,N_5993);
or U6029 (N_6029,N_5954,N_5802);
nor U6030 (N_6030,N_5888,N_5818);
and U6031 (N_6031,N_5845,N_5860);
and U6032 (N_6032,N_5806,N_5812);
xnor U6033 (N_6033,N_5950,N_5986);
xnor U6034 (N_6034,N_5894,N_5822);
or U6035 (N_6035,N_5832,N_5964);
or U6036 (N_6036,N_5877,N_5997);
nor U6037 (N_6037,N_5851,N_5857);
nor U6038 (N_6038,N_5931,N_5885);
and U6039 (N_6039,N_5938,N_5967);
nand U6040 (N_6040,N_5870,N_5804);
nand U6041 (N_6041,N_5826,N_5855);
xor U6042 (N_6042,N_5983,N_5922);
nor U6043 (N_6043,N_5859,N_5833);
and U6044 (N_6044,N_5836,N_5971);
xor U6045 (N_6045,N_5992,N_5949);
and U6046 (N_6046,N_5958,N_5811);
and U6047 (N_6047,N_5815,N_5838);
or U6048 (N_6048,N_5864,N_5926);
and U6049 (N_6049,N_5982,N_5900);
or U6050 (N_6050,N_5935,N_5884);
xnor U6051 (N_6051,N_5937,N_5985);
xnor U6052 (N_6052,N_5925,N_5843);
and U6053 (N_6053,N_5863,N_5910);
nand U6054 (N_6054,N_5901,N_5823);
xnor U6055 (N_6055,N_5987,N_5962);
xnor U6056 (N_6056,N_5830,N_5890);
nor U6057 (N_6057,N_5903,N_5862);
and U6058 (N_6058,N_5852,N_5842);
nor U6059 (N_6059,N_5990,N_5891);
or U6060 (N_6060,N_5879,N_5996);
nor U6061 (N_6061,N_5886,N_5866);
xnor U6062 (N_6062,N_5947,N_5934);
nor U6063 (N_6063,N_5976,N_5849);
or U6064 (N_6064,N_5899,N_5928);
nand U6065 (N_6065,N_5809,N_5827);
or U6066 (N_6066,N_5952,N_5975);
nand U6067 (N_6067,N_5968,N_5837);
and U6068 (N_6068,N_5821,N_5854);
and U6069 (N_6069,N_5800,N_5808);
nor U6070 (N_6070,N_5909,N_5989);
nor U6071 (N_6071,N_5820,N_5966);
or U6072 (N_6072,N_5991,N_5914);
and U6073 (N_6073,N_5805,N_5915);
xnor U6074 (N_6074,N_5955,N_5908);
xnor U6075 (N_6075,N_5876,N_5875);
and U6076 (N_6076,N_5906,N_5924);
xor U6077 (N_6077,N_5841,N_5882);
and U6078 (N_6078,N_5829,N_5817);
xnor U6079 (N_6079,N_5941,N_5905);
or U6080 (N_6080,N_5918,N_5972);
nor U6081 (N_6081,N_5848,N_5979);
or U6082 (N_6082,N_5880,N_5988);
or U6083 (N_6083,N_5895,N_5961);
or U6084 (N_6084,N_5872,N_5853);
and U6085 (N_6085,N_5819,N_5929);
nor U6086 (N_6086,N_5893,N_5828);
and U6087 (N_6087,N_5897,N_5846);
nor U6088 (N_6088,N_5984,N_5878);
or U6089 (N_6089,N_5883,N_5898);
nand U6090 (N_6090,N_5943,N_5940);
and U6091 (N_6091,N_5920,N_5917);
nor U6092 (N_6092,N_5834,N_5927);
and U6093 (N_6093,N_5916,N_5942);
xor U6094 (N_6094,N_5861,N_5871);
and U6095 (N_6095,N_5974,N_5869);
nor U6096 (N_6096,N_5814,N_5932);
xor U6097 (N_6097,N_5969,N_5913);
and U6098 (N_6098,N_5963,N_5825);
or U6099 (N_6099,N_5850,N_5936);
or U6100 (N_6100,N_5938,N_5842);
xnor U6101 (N_6101,N_5804,N_5999);
nor U6102 (N_6102,N_5871,N_5857);
nor U6103 (N_6103,N_5852,N_5874);
and U6104 (N_6104,N_5898,N_5891);
nor U6105 (N_6105,N_5925,N_5841);
or U6106 (N_6106,N_5804,N_5857);
or U6107 (N_6107,N_5930,N_5894);
or U6108 (N_6108,N_5958,N_5843);
or U6109 (N_6109,N_5863,N_5993);
nand U6110 (N_6110,N_5838,N_5876);
and U6111 (N_6111,N_5985,N_5924);
and U6112 (N_6112,N_5953,N_5884);
nand U6113 (N_6113,N_5853,N_5976);
nand U6114 (N_6114,N_5889,N_5867);
xor U6115 (N_6115,N_5929,N_5972);
or U6116 (N_6116,N_5941,N_5976);
nand U6117 (N_6117,N_5878,N_5820);
or U6118 (N_6118,N_5826,N_5835);
or U6119 (N_6119,N_5888,N_5984);
and U6120 (N_6120,N_5861,N_5991);
nor U6121 (N_6121,N_5856,N_5837);
xnor U6122 (N_6122,N_5835,N_5937);
and U6123 (N_6123,N_5915,N_5806);
or U6124 (N_6124,N_5844,N_5874);
nand U6125 (N_6125,N_5874,N_5948);
nand U6126 (N_6126,N_5825,N_5892);
xor U6127 (N_6127,N_5982,N_5852);
nand U6128 (N_6128,N_5856,N_5924);
and U6129 (N_6129,N_5930,N_5887);
and U6130 (N_6130,N_5949,N_5822);
nand U6131 (N_6131,N_5968,N_5861);
or U6132 (N_6132,N_5865,N_5855);
nand U6133 (N_6133,N_5967,N_5879);
nand U6134 (N_6134,N_5925,N_5907);
nor U6135 (N_6135,N_5938,N_5933);
or U6136 (N_6136,N_5807,N_5895);
or U6137 (N_6137,N_5959,N_5872);
xnor U6138 (N_6138,N_5903,N_5920);
nor U6139 (N_6139,N_5884,N_5980);
nand U6140 (N_6140,N_5844,N_5993);
xnor U6141 (N_6141,N_5842,N_5820);
and U6142 (N_6142,N_5896,N_5967);
xor U6143 (N_6143,N_5920,N_5954);
and U6144 (N_6144,N_5838,N_5902);
and U6145 (N_6145,N_5962,N_5945);
xor U6146 (N_6146,N_5992,N_5974);
nor U6147 (N_6147,N_5952,N_5841);
nor U6148 (N_6148,N_5892,N_5915);
and U6149 (N_6149,N_5849,N_5958);
or U6150 (N_6150,N_5968,N_5819);
nor U6151 (N_6151,N_5982,N_5906);
nand U6152 (N_6152,N_5994,N_5992);
xnor U6153 (N_6153,N_5864,N_5971);
nand U6154 (N_6154,N_5843,N_5800);
and U6155 (N_6155,N_5875,N_5869);
nand U6156 (N_6156,N_5955,N_5823);
xor U6157 (N_6157,N_5928,N_5966);
or U6158 (N_6158,N_5850,N_5826);
nor U6159 (N_6159,N_5965,N_5934);
nand U6160 (N_6160,N_5800,N_5851);
nand U6161 (N_6161,N_5817,N_5896);
xnor U6162 (N_6162,N_5909,N_5885);
and U6163 (N_6163,N_5980,N_5850);
or U6164 (N_6164,N_5894,N_5838);
or U6165 (N_6165,N_5992,N_5966);
or U6166 (N_6166,N_5904,N_5966);
xor U6167 (N_6167,N_5857,N_5951);
nor U6168 (N_6168,N_5942,N_5810);
and U6169 (N_6169,N_5833,N_5880);
xor U6170 (N_6170,N_5836,N_5991);
nor U6171 (N_6171,N_5881,N_5924);
and U6172 (N_6172,N_5880,N_5954);
xor U6173 (N_6173,N_5885,N_5877);
nand U6174 (N_6174,N_5977,N_5993);
xor U6175 (N_6175,N_5809,N_5807);
or U6176 (N_6176,N_5879,N_5962);
nor U6177 (N_6177,N_5868,N_5936);
or U6178 (N_6178,N_5999,N_5871);
and U6179 (N_6179,N_5917,N_5965);
nor U6180 (N_6180,N_5814,N_5998);
nor U6181 (N_6181,N_5805,N_5874);
nand U6182 (N_6182,N_5879,N_5815);
nor U6183 (N_6183,N_5900,N_5908);
nor U6184 (N_6184,N_5991,N_5941);
xor U6185 (N_6185,N_5901,N_5825);
nor U6186 (N_6186,N_5981,N_5871);
nand U6187 (N_6187,N_5857,N_5982);
and U6188 (N_6188,N_5951,N_5920);
xnor U6189 (N_6189,N_5866,N_5826);
and U6190 (N_6190,N_5900,N_5925);
and U6191 (N_6191,N_5959,N_5998);
nand U6192 (N_6192,N_5903,N_5805);
nand U6193 (N_6193,N_5999,N_5929);
or U6194 (N_6194,N_5892,N_5922);
or U6195 (N_6195,N_5929,N_5894);
nand U6196 (N_6196,N_5838,N_5870);
nor U6197 (N_6197,N_5917,N_5973);
nand U6198 (N_6198,N_5818,N_5986);
nand U6199 (N_6199,N_5971,N_5956);
nand U6200 (N_6200,N_6169,N_6105);
nor U6201 (N_6201,N_6155,N_6127);
nand U6202 (N_6202,N_6100,N_6102);
nor U6203 (N_6203,N_6171,N_6154);
nand U6204 (N_6204,N_6173,N_6037);
nand U6205 (N_6205,N_6012,N_6092);
xor U6206 (N_6206,N_6055,N_6160);
nand U6207 (N_6207,N_6096,N_6043);
and U6208 (N_6208,N_6073,N_6177);
xnor U6209 (N_6209,N_6195,N_6056);
xor U6210 (N_6210,N_6054,N_6159);
or U6211 (N_6211,N_6072,N_6052);
nand U6212 (N_6212,N_6185,N_6106);
and U6213 (N_6213,N_6027,N_6199);
xnor U6214 (N_6214,N_6198,N_6080);
nor U6215 (N_6215,N_6121,N_6086);
and U6216 (N_6216,N_6040,N_6175);
nor U6217 (N_6217,N_6015,N_6089);
or U6218 (N_6218,N_6031,N_6001);
xnor U6219 (N_6219,N_6062,N_6134);
and U6220 (N_6220,N_6085,N_6178);
nand U6221 (N_6221,N_6104,N_6066);
xnor U6222 (N_6222,N_6194,N_6125);
nor U6223 (N_6223,N_6141,N_6025);
xnor U6224 (N_6224,N_6146,N_6186);
and U6225 (N_6225,N_6192,N_6165);
or U6226 (N_6226,N_6189,N_6065);
nand U6227 (N_6227,N_6046,N_6011);
nor U6228 (N_6228,N_6020,N_6183);
and U6229 (N_6229,N_6042,N_6135);
nor U6230 (N_6230,N_6111,N_6017);
and U6231 (N_6231,N_6190,N_6068);
xnor U6232 (N_6232,N_6019,N_6117);
xor U6233 (N_6233,N_6147,N_6132);
and U6234 (N_6234,N_6197,N_6188);
or U6235 (N_6235,N_6145,N_6083);
nor U6236 (N_6236,N_6079,N_6182);
and U6237 (N_6237,N_6029,N_6174);
and U6238 (N_6238,N_6051,N_6059);
nor U6239 (N_6239,N_6170,N_6166);
nor U6240 (N_6240,N_6007,N_6140);
xnor U6241 (N_6241,N_6163,N_6181);
or U6242 (N_6242,N_6047,N_6143);
nor U6243 (N_6243,N_6149,N_6032);
or U6244 (N_6244,N_6036,N_6152);
or U6245 (N_6245,N_6024,N_6108);
and U6246 (N_6246,N_6058,N_6044);
nor U6247 (N_6247,N_6126,N_6022);
xnor U6248 (N_6248,N_6120,N_6028);
nand U6249 (N_6249,N_6090,N_6006);
xor U6250 (N_6250,N_6045,N_6093);
xnor U6251 (N_6251,N_6167,N_6041);
xor U6252 (N_6252,N_6076,N_6196);
nand U6253 (N_6253,N_6142,N_6081);
or U6254 (N_6254,N_6033,N_6087);
nand U6255 (N_6255,N_6023,N_6158);
xor U6256 (N_6256,N_6103,N_6018);
nor U6257 (N_6257,N_6187,N_6053);
xor U6258 (N_6258,N_6074,N_6097);
xnor U6259 (N_6259,N_6131,N_6164);
and U6260 (N_6260,N_6000,N_6168);
xor U6261 (N_6261,N_6057,N_6161);
and U6262 (N_6262,N_6050,N_6049);
nor U6263 (N_6263,N_6109,N_6156);
xor U6264 (N_6264,N_6150,N_6136);
nand U6265 (N_6265,N_6030,N_6077);
and U6266 (N_6266,N_6021,N_6180);
nand U6267 (N_6267,N_6075,N_6115);
nand U6268 (N_6268,N_6069,N_6008);
nand U6269 (N_6269,N_6067,N_6113);
nand U6270 (N_6270,N_6091,N_6088);
and U6271 (N_6271,N_6157,N_6039);
or U6272 (N_6272,N_6016,N_6179);
or U6273 (N_6273,N_6014,N_6002);
nor U6274 (N_6274,N_6184,N_6144);
and U6275 (N_6275,N_6009,N_6094);
and U6276 (N_6276,N_6133,N_6035);
and U6277 (N_6277,N_6193,N_6139);
nand U6278 (N_6278,N_6122,N_6010);
nor U6279 (N_6279,N_6004,N_6005);
or U6280 (N_6280,N_6095,N_6070);
or U6281 (N_6281,N_6060,N_6112);
or U6282 (N_6282,N_6013,N_6123);
nand U6283 (N_6283,N_6130,N_6078);
xor U6284 (N_6284,N_6151,N_6082);
nor U6285 (N_6285,N_6172,N_6129);
or U6286 (N_6286,N_6114,N_6148);
or U6287 (N_6287,N_6101,N_6116);
nand U6288 (N_6288,N_6071,N_6098);
xnor U6289 (N_6289,N_6162,N_6153);
nand U6290 (N_6290,N_6119,N_6107);
nand U6291 (N_6291,N_6110,N_6038);
nor U6292 (N_6292,N_6061,N_6034);
xnor U6293 (N_6293,N_6118,N_6138);
or U6294 (N_6294,N_6003,N_6063);
or U6295 (N_6295,N_6191,N_6176);
or U6296 (N_6296,N_6026,N_6099);
nand U6297 (N_6297,N_6124,N_6137);
or U6298 (N_6298,N_6128,N_6084);
nor U6299 (N_6299,N_6048,N_6064);
or U6300 (N_6300,N_6159,N_6087);
and U6301 (N_6301,N_6123,N_6149);
nand U6302 (N_6302,N_6080,N_6144);
nor U6303 (N_6303,N_6180,N_6026);
and U6304 (N_6304,N_6082,N_6057);
or U6305 (N_6305,N_6011,N_6174);
xnor U6306 (N_6306,N_6064,N_6128);
nand U6307 (N_6307,N_6084,N_6092);
nand U6308 (N_6308,N_6103,N_6096);
and U6309 (N_6309,N_6068,N_6195);
nand U6310 (N_6310,N_6043,N_6188);
nor U6311 (N_6311,N_6135,N_6072);
and U6312 (N_6312,N_6099,N_6041);
nand U6313 (N_6313,N_6154,N_6117);
and U6314 (N_6314,N_6033,N_6043);
xor U6315 (N_6315,N_6187,N_6178);
nand U6316 (N_6316,N_6084,N_6001);
and U6317 (N_6317,N_6035,N_6093);
or U6318 (N_6318,N_6134,N_6031);
and U6319 (N_6319,N_6136,N_6165);
and U6320 (N_6320,N_6004,N_6074);
nand U6321 (N_6321,N_6182,N_6090);
and U6322 (N_6322,N_6152,N_6060);
and U6323 (N_6323,N_6078,N_6108);
and U6324 (N_6324,N_6066,N_6113);
xnor U6325 (N_6325,N_6093,N_6132);
and U6326 (N_6326,N_6112,N_6002);
or U6327 (N_6327,N_6197,N_6199);
nand U6328 (N_6328,N_6078,N_6090);
nand U6329 (N_6329,N_6104,N_6195);
and U6330 (N_6330,N_6069,N_6067);
xnor U6331 (N_6331,N_6100,N_6148);
and U6332 (N_6332,N_6075,N_6163);
nor U6333 (N_6333,N_6031,N_6143);
nor U6334 (N_6334,N_6044,N_6086);
and U6335 (N_6335,N_6011,N_6097);
xor U6336 (N_6336,N_6150,N_6172);
and U6337 (N_6337,N_6121,N_6117);
and U6338 (N_6338,N_6082,N_6068);
nor U6339 (N_6339,N_6162,N_6121);
nand U6340 (N_6340,N_6179,N_6027);
and U6341 (N_6341,N_6181,N_6111);
nor U6342 (N_6342,N_6129,N_6118);
nor U6343 (N_6343,N_6082,N_6060);
nor U6344 (N_6344,N_6071,N_6174);
xor U6345 (N_6345,N_6015,N_6141);
xnor U6346 (N_6346,N_6168,N_6041);
nor U6347 (N_6347,N_6044,N_6191);
nor U6348 (N_6348,N_6100,N_6036);
nor U6349 (N_6349,N_6024,N_6169);
or U6350 (N_6350,N_6170,N_6145);
or U6351 (N_6351,N_6045,N_6152);
and U6352 (N_6352,N_6005,N_6196);
and U6353 (N_6353,N_6186,N_6066);
and U6354 (N_6354,N_6075,N_6013);
xor U6355 (N_6355,N_6127,N_6165);
nor U6356 (N_6356,N_6026,N_6165);
and U6357 (N_6357,N_6045,N_6156);
and U6358 (N_6358,N_6194,N_6118);
or U6359 (N_6359,N_6072,N_6018);
xnor U6360 (N_6360,N_6138,N_6100);
and U6361 (N_6361,N_6035,N_6187);
or U6362 (N_6362,N_6131,N_6003);
and U6363 (N_6363,N_6005,N_6009);
nor U6364 (N_6364,N_6019,N_6002);
nand U6365 (N_6365,N_6018,N_6078);
xor U6366 (N_6366,N_6040,N_6095);
xnor U6367 (N_6367,N_6072,N_6024);
nor U6368 (N_6368,N_6122,N_6040);
or U6369 (N_6369,N_6133,N_6052);
and U6370 (N_6370,N_6158,N_6185);
nor U6371 (N_6371,N_6169,N_6021);
or U6372 (N_6372,N_6107,N_6134);
or U6373 (N_6373,N_6031,N_6187);
xnor U6374 (N_6374,N_6164,N_6058);
xor U6375 (N_6375,N_6001,N_6180);
or U6376 (N_6376,N_6048,N_6095);
and U6377 (N_6377,N_6018,N_6025);
xnor U6378 (N_6378,N_6102,N_6045);
nand U6379 (N_6379,N_6185,N_6076);
or U6380 (N_6380,N_6034,N_6109);
nor U6381 (N_6381,N_6190,N_6006);
nor U6382 (N_6382,N_6106,N_6043);
or U6383 (N_6383,N_6042,N_6097);
nor U6384 (N_6384,N_6125,N_6059);
nor U6385 (N_6385,N_6091,N_6125);
nor U6386 (N_6386,N_6193,N_6092);
nand U6387 (N_6387,N_6151,N_6000);
nand U6388 (N_6388,N_6110,N_6030);
nand U6389 (N_6389,N_6046,N_6133);
and U6390 (N_6390,N_6013,N_6176);
xnor U6391 (N_6391,N_6148,N_6019);
and U6392 (N_6392,N_6108,N_6157);
xnor U6393 (N_6393,N_6096,N_6172);
and U6394 (N_6394,N_6023,N_6116);
nor U6395 (N_6395,N_6023,N_6014);
xor U6396 (N_6396,N_6071,N_6137);
nand U6397 (N_6397,N_6182,N_6027);
or U6398 (N_6398,N_6172,N_6020);
or U6399 (N_6399,N_6183,N_6147);
xor U6400 (N_6400,N_6257,N_6296);
or U6401 (N_6401,N_6289,N_6376);
nor U6402 (N_6402,N_6205,N_6390);
nor U6403 (N_6403,N_6388,N_6303);
xnor U6404 (N_6404,N_6355,N_6395);
nand U6405 (N_6405,N_6278,N_6258);
nor U6406 (N_6406,N_6383,N_6329);
or U6407 (N_6407,N_6262,N_6269);
nand U6408 (N_6408,N_6304,N_6350);
and U6409 (N_6409,N_6327,N_6239);
xor U6410 (N_6410,N_6307,N_6325);
nand U6411 (N_6411,N_6337,N_6276);
xor U6412 (N_6412,N_6288,N_6221);
xnor U6413 (N_6413,N_6238,N_6213);
nand U6414 (N_6414,N_6268,N_6387);
nor U6415 (N_6415,N_6243,N_6374);
and U6416 (N_6416,N_6373,N_6361);
or U6417 (N_6417,N_6246,N_6314);
nand U6418 (N_6418,N_6399,N_6302);
nand U6419 (N_6419,N_6287,N_6209);
or U6420 (N_6420,N_6280,N_6294);
nor U6421 (N_6421,N_6382,N_6323);
xnor U6422 (N_6422,N_6375,N_6384);
and U6423 (N_6423,N_6250,N_6217);
nand U6424 (N_6424,N_6347,N_6311);
and U6425 (N_6425,N_6206,N_6378);
nand U6426 (N_6426,N_6398,N_6356);
or U6427 (N_6427,N_6233,N_6218);
nor U6428 (N_6428,N_6219,N_6393);
or U6429 (N_6429,N_6254,N_6333);
nand U6430 (N_6430,N_6208,N_6335);
and U6431 (N_6431,N_6271,N_6253);
xnor U6432 (N_6432,N_6312,N_6348);
or U6433 (N_6433,N_6214,N_6277);
nand U6434 (N_6434,N_6203,N_6386);
xor U6435 (N_6435,N_6265,N_6344);
xnor U6436 (N_6436,N_6308,N_6310);
nor U6437 (N_6437,N_6305,N_6232);
and U6438 (N_6438,N_6245,N_6379);
xnor U6439 (N_6439,N_6227,N_6255);
xor U6440 (N_6440,N_6229,N_6292);
nor U6441 (N_6441,N_6334,N_6241);
or U6442 (N_6442,N_6352,N_6363);
xnor U6443 (N_6443,N_6298,N_6364);
xnor U6444 (N_6444,N_6264,N_6207);
and U6445 (N_6445,N_6313,N_6336);
xnor U6446 (N_6446,N_6358,N_6392);
or U6447 (N_6447,N_6222,N_6346);
xor U6448 (N_6448,N_6234,N_6366);
xor U6449 (N_6449,N_6370,N_6372);
xor U6450 (N_6450,N_6275,N_6223);
xnor U6451 (N_6451,N_6319,N_6212);
or U6452 (N_6452,N_6283,N_6291);
and U6453 (N_6453,N_6357,N_6306);
nor U6454 (N_6454,N_6349,N_6354);
nand U6455 (N_6455,N_6318,N_6389);
nor U6456 (N_6456,N_6228,N_6396);
or U6457 (N_6457,N_6252,N_6377);
or U6458 (N_6458,N_6381,N_6261);
xor U6459 (N_6459,N_6320,N_6345);
nand U6460 (N_6460,N_6247,N_6328);
xnor U6461 (N_6461,N_6279,N_6249);
and U6462 (N_6462,N_6281,N_6297);
nor U6463 (N_6463,N_6362,N_6341);
nor U6464 (N_6464,N_6359,N_6266);
xnor U6465 (N_6465,N_6235,N_6295);
or U6466 (N_6466,N_6263,N_6340);
and U6467 (N_6467,N_6201,N_6394);
and U6468 (N_6468,N_6244,N_6368);
nand U6469 (N_6469,N_6200,N_6270);
nand U6470 (N_6470,N_6342,N_6286);
or U6471 (N_6471,N_6339,N_6224);
nand U6472 (N_6472,N_6365,N_6237);
and U6473 (N_6473,N_6282,N_6316);
nand U6474 (N_6474,N_6315,N_6301);
nand U6475 (N_6475,N_6299,N_6371);
nand U6476 (N_6476,N_6317,N_6240);
or U6477 (N_6477,N_6220,N_6215);
or U6478 (N_6478,N_6360,N_6369);
nand U6479 (N_6479,N_6300,N_6202);
and U6480 (N_6480,N_6332,N_6211);
xor U6481 (N_6481,N_6338,N_6290);
and U6482 (N_6482,N_6330,N_6248);
nand U6483 (N_6483,N_6331,N_6267);
nand U6484 (N_6484,N_6260,N_6226);
nand U6485 (N_6485,N_6259,N_6322);
xor U6486 (N_6486,N_6343,N_6216);
xnor U6487 (N_6487,N_6293,N_6251);
xor U6488 (N_6488,N_6242,N_6324);
and U6489 (N_6489,N_6225,N_6351);
or U6490 (N_6490,N_6273,N_6353);
or U6491 (N_6491,N_6367,N_6397);
or U6492 (N_6492,N_6284,N_6210);
nor U6493 (N_6493,N_6321,N_6385);
xor U6494 (N_6494,N_6230,N_6391);
nand U6495 (N_6495,N_6204,N_6274);
and U6496 (N_6496,N_6256,N_6380);
or U6497 (N_6497,N_6285,N_6272);
nor U6498 (N_6498,N_6231,N_6309);
xor U6499 (N_6499,N_6236,N_6326);
nand U6500 (N_6500,N_6280,N_6345);
xor U6501 (N_6501,N_6375,N_6220);
nor U6502 (N_6502,N_6307,N_6216);
or U6503 (N_6503,N_6339,N_6384);
xnor U6504 (N_6504,N_6349,N_6219);
nor U6505 (N_6505,N_6363,N_6252);
xnor U6506 (N_6506,N_6307,N_6221);
nand U6507 (N_6507,N_6350,N_6290);
nor U6508 (N_6508,N_6271,N_6272);
xor U6509 (N_6509,N_6235,N_6337);
xnor U6510 (N_6510,N_6326,N_6394);
xor U6511 (N_6511,N_6395,N_6228);
and U6512 (N_6512,N_6213,N_6212);
or U6513 (N_6513,N_6301,N_6340);
nor U6514 (N_6514,N_6324,N_6251);
nor U6515 (N_6515,N_6303,N_6365);
xnor U6516 (N_6516,N_6316,N_6286);
xor U6517 (N_6517,N_6274,N_6357);
nor U6518 (N_6518,N_6365,N_6233);
nor U6519 (N_6519,N_6224,N_6281);
nor U6520 (N_6520,N_6362,N_6378);
xnor U6521 (N_6521,N_6360,N_6370);
and U6522 (N_6522,N_6202,N_6258);
and U6523 (N_6523,N_6375,N_6247);
or U6524 (N_6524,N_6312,N_6232);
xor U6525 (N_6525,N_6371,N_6333);
nand U6526 (N_6526,N_6231,N_6272);
and U6527 (N_6527,N_6207,N_6209);
or U6528 (N_6528,N_6236,N_6200);
xor U6529 (N_6529,N_6235,N_6264);
nand U6530 (N_6530,N_6271,N_6226);
or U6531 (N_6531,N_6378,N_6333);
nand U6532 (N_6532,N_6212,N_6382);
and U6533 (N_6533,N_6399,N_6294);
nor U6534 (N_6534,N_6385,N_6358);
and U6535 (N_6535,N_6229,N_6394);
xor U6536 (N_6536,N_6234,N_6303);
nor U6537 (N_6537,N_6281,N_6360);
or U6538 (N_6538,N_6219,N_6285);
nor U6539 (N_6539,N_6380,N_6278);
and U6540 (N_6540,N_6357,N_6348);
nand U6541 (N_6541,N_6220,N_6203);
or U6542 (N_6542,N_6378,N_6248);
nor U6543 (N_6543,N_6343,N_6345);
xor U6544 (N_6544,N_6369,N_6303);
or U6545 (N_6545,N_6381,N_6266);
nor U6546 (N_6546,N_6379,N_6315);
nor U6547 (N_6547,N_6309,N_6326);
nor U6548 (N_6548,N_6289,N_6226);
nor U6549 (N_6549,N_6264,N_6321);
or U6550 (N_6550,N_6294,N_6220);
and U6551 (N_6551,N_6278,N_6397);
nand U6552 (N_6552,N_6308,N_6302);
and U6553 (N_6553,N_6208,N_6328);
and U6554 (N_6554,N_6296,N_6357);
or U6555 (N_6555,N_6200,N_6386);
xnor U6556 (N_6556,N_6368,N_6255);
nor U6557 (N_6557,N_6378,N_6200);
or U6558 (N_6558,N_6399,N_6336);
nor U6559 (N_6559,N_6226,N_6380);
xor U6560 (N_6560,N_6379,N_6293);
or U6561 (N_6561,N_6308,N_6266);
nand U6562 (N_6562,N_6303,N_6286);
xor U6563 (N_6563,N_6347,N_6250);
or U6564 (N_6564,N_6274,N_6343);
nand U6565 (N_6565,N_6331,N_6252);
or U6566 (N_6566,N_6214,N_6283);
nand U6567 (N_6567,N_6264,N_6239);
xnor U6568 (N_6568,N_6203,N_6371);
and U6569 (N_6569,N_6333,N_6219);
nand U6570 (N_6570,N_6377,N_6222);
xnor U6571 (N_6571,N_6227,N_6220);
and U6572 (N_6572,N_6285,N_6224);
xor U6573 (N_6573,N_6271,N_6308);
nand U6574 (N_6574,N_6346,N_6304);
xnor U6575 (N_6575,N_6342,N_6364);
xor U6576 (N_6576,N_6239,N_6277);
and U6577 (N_6577,N_6300,N_6204);
xnor U6578 (N_6578,N_6260,N_6268);
nor U6579 (N_6579,N_6291,N_6246);
xor U6580 (N_6580,N_6323,N_6355);
and U6581 (N_6581,N_6248,N_6266);
nor U6582 (N_6582,N_6217,N_6232);
nor U6583 (N_6583,N_6230,N_6221);
xor U6584 (N_6584,N_6378,N_6205);
xnor U6585 (N_6585,N_6321,N_6392);
nor U6586 (N_6586,N_6229,N_6212);
nor U6587 (N_6587,N_6340,N_6339);
xor U6588 (N_6588,N_6291,N_6275);
or U6589 (N_6589,N_6245,N_6227);
nor U6590 (N_6590,N_6241,N_6269);
and U6591 (N_6591,N_6234,N_6328);
xnor U6592 (N_6592,N_6281,N_6356);
or U6593 (N_6593,N_6278,N_6215);
nand U6594 (N_6594,N_6361,N_6229);
or U6595 (N_6595,N_6351,N_6243);
and U6596 (N_6596,N_6396,N_6307);
nor U6597 (N_6597,N_6378,N_6246);
xor U6598 (N_6598,N_6346,N_6317);
and U6599 (N_6599,N_6253,N_6378);
xnor U6600 (N_6600,N_6505,N_6599);
xor U6601 (N_6601,N_6557,N_6465);
xnor U6602 (N_6602,N_6534,N_6506);
and U6603 (N_6603,N_6484,N_6524);
xor U6604 (N_6604,N_6452,N_6574);
xnor U6605 (N_6605,N_6543,N_6434);
or U6606 (N_6606,N_6538,N_6542);
and U6607 (N_6607,N_6489,N_6576);
nand U6608 (N_6608,N_6436,N_6537);
or U6609 (N_6609,N_6412,N_6588);
nand U6610 (N_6610,N_6570,N_6456);
nand U6611 (N_6611,N_6491,N_6450);
nor U6612 (N_6612,N_6468,N_6567);
and U6613 (N_6613,N_6454,N_6558);
xnor U6614 (N_6614,N_6500,N_6470);
xnor U6615 (N_6615,N_6564,N_6415);
or U6616 (N_6616,N_6529,N_6428);
and U6617 (N_6617,N_6481,N_6582);
nor U6618 (N_6618,N_6403,N_6493);
nand U6619 (N_6619,N_6466,N_6523);
and U6620 (N_6620,N_6424,N_6482);
nor U6621 (N_6621,N_6515,N_6581);
xor U6622 (N_6622,N_6535,N_6411);
or U6623 (N_6623,N_6420,N_6573);
and U6624 (N_6624,N_6565,N_6519);
or U6625 (N_6625,N_6554,N_6553);
and U6626 (N_6626,N_6541,N_6591);
nand U6627 (N_6627,N_6414,N_6563);
or U6628 (N_6628,N_6475,N_6413);
and U6629 (N_6629,N_6511,N_6528);
or U6630 (N_6630,N_6516,N_6406);
nor U6631 (N_6631,N_6510,N_6501);
and U6632 (N_6632,N_6400,N_6552);
or U6633 (N_6633,N_6546,N_6592);
xnor U6634 (N_6634,N_6458,N_6539);
or U6635 (N_6635,N_6462,N_6597);
nand U6636 (N_6636,N_6522,N_6585);
and U6637 (N_6637,N_6547,N_6596);
xor U6638 (N_6638,N_6512,N_6430);
xnor U6639 (N_6639,N_6531,N_6401);
xor U6640 (N_6640,N_6410,N_6440);
xnor U6641 (N_6641,N_6459,N_6530);
or U6642 (N_6642,N_6532,N_6409);
or U6643 (N_6643,N_6548,N_6425);
xnor U6644 (N_6644,N_6569,N_6568);
nand U6645 (N_6645,N_6432,N_6586);
xnor U6646 (N_6646,N_6504,N_6513);
and U6647 (N_6647,N_6476,N_6584);
nand U6648 (N_6648,N_6453,N_6488);
or U6649 (N_6649,N_6487,N_6408);
xnor U6650 (N_6650,N_6467,N_6480);
or U6651 (N_6651,N_6473,N_6499);
and U6652 (N_6652,N_6580,N_6445);
nor U6653 (N_6653,N_6517,N_6478);
nor U6654 (N_6654,N_6544,N_6433);
and U6655 (N_6655,N_6422,N_6598);
nor U6656 (N_6656,N_6579,N_6427);
or U6657 (N_6657,N_6578,N_6561);
or U6658 (N_6658,N_6404,N_6438);
xnor U6659 (N_6659,N_6559,N_6560);
nand U6660 (N_6660,N_6502,N_6521);
nor U6661 (N_6661,N_6464,N_6572);
xor U6662 (N_6662,N_6441,N_6485);
xor U6663 (N_6663,N_6405,N_6429);
and U6664 (N_6664,N_6447,N_6518);
or U6665 (N_6665,N_6494,N_6419);
and U6666 (N_6666,N_6444,N_6469);
and U6667 (N_6667,N_6439,N_6437);
nand U6668 (N_6668,N_6446,N_6471);
nand U6669 (N_6669,N_6562,N_6508);
nor U6670 (N_6670,N_6503,N_6555);
nand U6671 (N_6671,N_6577,N_6556);
and U6672 (N_6672,N_6590,N_6497);
or U6673 (N_6673,N_6431,N_6455);
nand U6674 (N_6674,N_6477,N_6461);
or U6675 (N_6675,N_6421,N_6495);
or U6676 (N_6676,N_6566,N_6595);
or U6677 (N_6677,N_6575,N_6426);
nor U6678 (N_6678,N_6418,N_6571);
xnor U6679 (N_6679,N_6448,N_6540);
nor U6680 (N_6680,N_6463,N_6549);
nand U6681 (N_6681,N_6460,N_6509);
xnor U6682 (N_6682,N_6435,N_6490);
nand U6683 (N_6683,N_6423,N_6583);
nor U6684 (N_6684,N_6593,N_6474);
xnor U6685 (N_6685,N_6527,N_6449);
nor U6686 (N_6686,N_6496,N_6443);
nand U6687 (N_6687,N_6407,N_6498);
nand U6688 (N_6688,N_6514,N_6402);
nand U6689 (N_6689,N_6536,N_6416);
xnor U6690 (N_6690,N_6442,N_6417);
or U6691 (N_6691,N_6479,N_6533);
xnor U6692 (N_6692,N_6545,N_6472);
and U6693 (N_6693,N_6550,N_6525);
nor U6694 (N_6694,N_6526,N_6551);
nor U6695 (N_6695,N_6594,N_6507);
nand U6696 (N_6696,N_6589,N_6483);
nor U6697 (N_6697,N_6492,N_6520);
and U6698 (N_6698,N_6587,N_6486);
nand U6699 (N_6699,N_6457,N_6451);
xnor U6700 (N_6700,N_6528,N_6476);
xor U6701 (N_6701,N_6480,N_6534);
or U6702 (N_6702,N_6531,N_6598);
xor U6703 (N_6703,N_6507,N_6526);
nor U6704 (N_6704,N_6478,N_6516);
xnor U6705 (N_6705,N_6404,N_6481);
and U6706 (N_6706,N_6529,N_6579);
nor U6707 (N_6707,N_6422,N_6413);
and U6708 (N_6708,N_6456,N_6554);
and U6709 (N_6709,N_6411,N_6420);
xor U6710 (N_6710,N_6520,N_6570);
or U6711 (N_6711,N_6534,N_6453);
nor U6712 (N_6712,N_6450,N_6490);
nand U6713 (N_6713,N_6422,N_6466);
or U6714 (N_6714,N_6545,N_6453);
and U6715 (N_6715,N_6462,N_6424);
nor U6716 (N_6716,N_6580,N_6511);
nor U6717 (N_6717,N_6504,N_6566);
and U6718 (N_6718,N_6461,N_6408);
nor U6719 (N_6719,N_6423,N_6558);
or U6720 (N_6720,N_6484,N_6593);
or U6721 (N_6721,N_6528,N_6461);
and U6722 (N_6722,N_6553,N_6435);
or U6723 (N_6723,N_6433,N_6498);
xnor U6724 (N_6724,N_6566,N_6551);
nor U6725 (N_6725,N_6424,N_6457);
or U6726 (N_6726,N_6464,N_6423);
xor U6727 (N_6727,N_6429,N_6422);
and U6728 (N_6728,N_6531,N_6556);
xnor U6729 (N_6729,N_6428,N_6554);
or U6730 (N_6730,N_6464,N_6568);
or U6731 (N_6731,N_6550,N_6436);
nor U6732 (N_6732,N_6453,N_6409);
nor U6733 (N_6733,N_6465,N_6536);
nand U6734 (N_6734,N_6513,N_6563);
or U6735 (N_6735,N_6489,N_6596);
nor U6736 (N_6736,N_6519,N_6468);
nor U6737 (N_6737,N_6526,N_6564);
xnor U6738 (N_6738,N_6576,N_6429);
nand U6739 (N_6739,N_6401,N_6444);
xnor U6740 (N_6740,N_6451,N_6472);
nor U6741 (N_6741,N_6540,N_6516);
xnor U6742 (N_6742,N_6543,N_6521);
and U6743 (N_6743,N_6499,N_6464);
and U6744 (N_6744,N_6505,N_6400);
nand U6745 (N_6745,N_6597,N_6450);
nand U6746 (N_6746,N_6484,N_6596);
and U6747 (N_6747,N_6490,N_6434);
and U6748 (N_6748,N_6515,N_6418);
nor U6749 (N_6749,N_6456,N_6496);
nand U6750 (N_6750,N_6407,N_6514);
or U6751 (N_6751,N_6560,N_6448);
nor U6752 (N_6752,N_6532,N_6557);
nand U6753 (N_6753,N_6513,N_6452);
xor U6754 (N_6754,N_6404,N_6472);
nand U6755 (N_6755,N_6423,N_6596);
and U6756 (N_6756,N_6435,N_6475);
or U6757 (N_6757,N_6404,N_6423);
or U6758 (N_6758,N_6404,N_6445);
nor U6759 (N_6759,N_6568,N_6421);
nand U6760 (N_6760,N_6462,N_6463);
nand U6761 (N_6761,N_6493,N_6569);
and U6762 (N_6762,N_6526,N_6588);
and U6763 (N_6763,N_6533,N_6447);
nor U6764 (N_6764,N_6585,N_6496);
and U6765 (N_6765,N_6529,N_6500);
xor U6766 (N_6766,N_6513,N_6449);
xor U6767 (N_6767,N_6425,N_6420);
and U6768 (N_6768,N_6536,N_6405);
xor U6769 (N_6769,N_6505,N_6535);
nand U6770 (N_6770,N_6515,N_6555);
or U6771 (N_6771,N_6425,N_6597);
or U6772 (N_6772,N_6502,N_6410);
xor U6773 (N_6773,N_6520,N_6405);
nand U6774 (N_6774,N_6401,N_6560);
or U6775 (N_6775,N_6573,N_6416);
nand U6776 (N_6776,N_6412,N_6480);
and U6777 (N_6777,N_6467,N_6513);
xor U6778 (N_6778,N_6472,N_6473);
or U6779 (N_6779,N_6552,N_6526);
nand U6780 (N_6780,N_6552,N_6519);
and U6781 (N_6781,N_6487,N_6418);
and U6782 (N_6782,N_6535,N_6551);
or U6783 (N_6783,N_6566,N_6454);
and U6784 (N_6784,N_6539,N_6556);
xnor U6785 (N_6785,N_6527,N_6579);
nand U6786 (N_6786,N_6562,N_6457);
and U6787 (N_6787,N_6498,N_6466);
xor U6788 (N_6788,N_6400,N_6589);
and U6789 (N_6789,N_6524,N_6544);
and U6790 (N_6790,N_6465,N_6479);
or U6791 (N_6791,N_6422,N_6475);
or U6792 (N_6792,N_6488,N_6557);
and U6793 (N_6793,N_6437,N_6463);
nand U6794 (N_6794,N_6580,N_6512);
and U6795 (N_6795,N_6523,N_6452);
xnor U6796 (N_6796,N_6422,N_6426);
and U6797 (N_6797,N_6419,N_6517);
xor U6798 (N_6798,N_6596,N_6448);
nor U6799 (N_6799,N_6401,N_6562);
nand U6800 (N_6800,N_6668,N_6776);
or U6801 (N_6801,N_6688,N_6730);
and U6802 (N_6802,N_6789,N_6694);
nand U6803 (N_6803,N_6722,N_6637);
or U6804 (N_6804,N_6727,N_6713);
nor U6805 (N_6805,N_6720,N_6621);
or U6806 (N_6806,N_6653,N_6699);
or U6807 (N_6807,N_6746,N_6629);
xor U6808 (N_6808,N_6604,N_6648);
nand U6809 (N_6809,N_6601,N_6704);
xor U6810 (N_6810,N_6770,N_6673);
nor U6811 (N_6811,N_6618,N_6641);
nand U6812 (N_6812,N_6771,N_6686);
or U6813 (N_6813,N_6785,N_6797);
or U6814 (N_6814,N_6775,N_6600);
xnor U6815 (N_6815,N_6607,N_6687);
nand U6816 (N_6816,N_6658,N_6700);
or U6817 (N_6817,N_6761,N_6677);
or U6818 (N_6818,N_6634,N_6769);
nor U6819 (N_6819,N_6630,N_6717);
nor U6820 (N_6820,N_6609,N_6611);
xor U6821 (N_6821,N_6643,N_6794);
or U6822 (N_6822,N_6685,N_6735);
xnor U6823 (N_6823,N_6627,N_6610);
nor U6824 (N_6824,N_6777,N_6636);
xor U6825 (N_6825,N_6613,N_6721);
or U6826 (N_6826,N_6750,N_6795);
or U6827 (N_6827,N_6614,N_6663);
nand U6828 (N_6828,N_6726,N_6645);
xnor U6829 (N_6829,N_6734,N_6741);
and U6830 (N_6830,N_6620,N_6683);
or U6831 (N_6831,N_6796,N_6725);
and U6832 (N_6832,N_6684,N_6605);
and U6833 (N_6833,N_6774,N_6642);
and U6834 (N_6834,N_6657,N_6754);
xor U6835 (N_6835,N_6651,N_6612);
xnor U6836 (N_6836,N_6788,N_6772);
nand U6837 (N_6837,N_6675,N_6639);
or U6838 (N_6838,N_6757,N_6659);
nor U6839 (N_6839,N_6792,N_6631);
and U6840 (N_6840,N_6758,N_6670);
and U6841 (N_6841,N_6692,N_6752);
and U6842 (N_6842,N_6678,N_6695);
or U6843 (N_6843,N_6703,N_6705);
xor U6844 (N_6844,N_6737,N_6674);
or U6845 (N_6845,N_6664,N_6728);
or U6846 (N_6846,N_6667,N_6766);
nand U6847 (N_6847,N_6743,N_6778);
or U6848 (N_6848,N_6798,N_6644);
xor U6849 (N_6849,N_6744,N_6784);
xor U6850 (N_6850,N_6635,N_6606);
nand U6851 (N_6851,N_6655,N_6628);
xnor U6852 (N_6852,N_6619,N_6764);
xor U6853 (N_6853,N_6665,N_6747);
or U6854 (N_6854,N_6765,N_6768);
and U6855 (N_6855,N_6696,N_6753);
or U6856 (N_6856,N_6679,N_6603);
xor U6857 (N_6857,N_6723,N_6739);
nor U6858 (N_6858,N_6779,N_6740);
nor U6859 (N_6859,N_6652,N_6762);
nand U6860 (N_6860,N_6671,N_6697);
nor U6861 (N_6861,N_6650,N_6759);
nand U6862 (N_6862,N_6669,N_6693);
nand U6863 (N_6863,N_6712,N_6625);
nand U6864 (N_6864,N_6742,N_6719);
nor U6865 (N_6865,N_6654,N_6672);
nand U6866 (N_6866,N_6714,N_6680);
and U6867 (N_6867,N_6640,N_6755);
and U6868 (N_6868,N_6733,N_6701);
xnor U6869 (N_6869,N_6790,N_6660);
nor U6870 (N_6870,N_6690,N_6689);
or U6871 (N_6871,N_6745,N_6738);
nand U6872 (N_6872,N_6646,N_6763);
xnor U6873 (N_6873,N_6780,N_6787);
nor U6874 (N_6874,N_6602,N_6767);
or U6875 (N_6875,N_6661,N_6782);
xor U6876 (N_6876,N_6793,N_6633);
nand U6877 (N_6877,N_6702,N_6624);
nor U6878 (N_6878,N_6691,N_6608);
xnor U6879 (N_6879,N_6791,N_6666);
or U6880 (N_6880,N_6724,N_6732);
and U6881 (N_6881,N_6783,N_6707);
xnor U6882 (N_6882,N_6656,N_6626);
nor U6883 (N_6883,N_6756,N_6706);
xnor U6884 (N_6884,N_6749,N_6632);
nand U6885 (N_6885,N_6682,N_6781);
nor U6886 (N_6886,N_6799,N_6715);
nor U6887 (N_6887,N_6760,N_6649);
or U6888 (N_6888,N_6638,N_6617);
xnor U6889 (N_6889,N_6716,N_6615);
and U6890 (N_6890,N_6709,N_6698);
or U6891 (N_6891,N_6718,N_6748);
nand U6892 (N_6892,N_6616,N_6731);
nand U6893 (N_6893,N_6623,N_6710);
nand U6894 (N_6894,N_6711,N_6708);
xnor U6895 (N_6895,N_6676,N_6681);
and U6896 (N_6896,N_6622,N_6751);
nand U6897 (N_6897,N_6773,N_6662);
and U6898 (N_6898,N_6729,N_6736);
or U6899 (N_6899,N_6786,N_6647);
xor U6900 (N_6900,N_6623,N_6634);
nand U6901 (N_6901,N_6699,N_6742);
xor U6902 (N_6902,N_6668,N_6718);
nor U6903 (N_6903,N_6626,N_6788);
xnor U6904 (N_6904,N_6782,N_6761);
xnor U6905 (N_6905,N_6605,N_6722);
nand U6906 (N_6906,N_6668,N_6749);
or U6907 (N_6907,N_6796,N_6662);
nand U6908 (N_6908,N_6626,N_6727);
and U6909 (N_6909,N_6771,N_6727);
nand U6910 (N_6910,N_6789,N_6737);
or U6911 (N_6911,N_6609,N_6796);
nor U6912 (N_6912,N_6724,N_6642);
and U6913 (N_6913,N_6721,N_6772);
nand U6914 (N_6914,N_6732,N_6609);
or U6915 (N_6915,N_6739,N_6649);
or U6916 (N_6916,N_6636,N_6600);
nand U6917 (N_6917,N_6670,N_6788);
nor U6918 (N_6918,N_6788,N_6760);
and U6919 (N_6919,N_6685,N_6771);
and U6920 (N_6920,N_6614,N_6777);
and U6921 (N_6921,N_6685,N_6649);
nor U6922 (N_6922,N_6734,N_6733);
and U6923 (N_6923,N_6725,N_6723);
and U6924 (N_6924,N_6603,N_6667);
xor U6925 (N_6925,N_6740,N_6799);
and U6926 (N_6926,N_6719,N_6645);
or U6927 (N_6927,N_6605,N_6661);
and U6928 (N_6928,N_6798,N_6795);
and U6929 (N_6929,N_6753,N_6792);
nor U6930 (N_6930,N_6732,N_6654);
nand U6931 (N_6931,N_6650,N_6790);
or U6932 (N_6932,N_6643,N_6697);
and U6933 (N_6933,N_6654,N_6782);
or U6934 (N_6934,N_6723,N_6786);
or U6935 (N_6935,N_6627,N_6743);
nand U6936 (N_6936,N_6764,N_6704);
nand U6937 (N_6937,N_6719,N_6643);
or U6938 (N_6938,N_6697,N_6674);
or U6939 (N_6939,N_6729,N_6621);
nand U6940 (N_6940,N_6697,N_6771);
nand U6941 (N_6941,N_6671,N_6700);
nor U6942 (N_6942,N_6628,N_6615);
nand U6943 (N_6943,N_6623,N_6600);
or U6944 (N_6944,N_6620,N_6758);
nor U6945 (N_6945,N_6697,N_6607);
and U6946 (N_6946,N_6732,N_6766);
and U6947 (N_6947,N_6645,N_6616);
and U6948 (N_6948,N_6647,N_6751);
xor U6949 (N_6949,N_6644,N_6618);
or U6950 (N_6950,N_6607,N_6678);
nor U6951 (N_6951,N_6624,N_6759);
or U6952 (N_6952,N_6606,N_6708);
and U6953 (N_6953,N_6770,N_6734);
nor U6954 (N_6954,N_6620,N_6669);
xor U6955 (N_6955,N_6636,N_6684);
or U6956 (N_6956,N_6719,N_6793);
nand U6957 (N_6957,N_6674,N_6652);
xor U6958 (N_6958,N_6690,N_6625);
and U6959 (N_6959,N_6702,N_6629);
and U6960 (N_6960,N_6785,N_6786);
xor U6961 (N_6961,N_6778,N_6610);
and U6962 (N_6962,N_6744,N_6749);
nand U6963 (N_6963,N_6772,N_6621);
nand U6964 (N_6964,N_6711,N_6687);
or U6965 (N_6965,N_6734,N_6777);
xnor U6966 (N_6966,N_6679,N_6651);
xor U6967 (N_6967,N_6624,N_6697);
or U6968 (N_6968,N_6790,N_6674);
nor U6969 (N_6969,N_6767,N_6789);
or U6970 (N_6970,N_6684,N_6719);
xnor U6971 (N_6971,N_6797,N_6740);
nor U6972 (N_6972,N_6783,N_6789);
nor U6973 (N_6973,N_6759,N_6774);
nand U6974 (N_6974,N_6739,N_6677);
nand U6975 (N_6975,N_6755,N_6734);
and U6976 (N_6976,N_6758,N_6769);
or U6977 (N_6977,N_6635,N_6734);
nor U6978 (N_6978,N_6710,N_6721);
nand U6979 (N_6979,N_6656,N_6613);
nor U6980 (N_6980,N_6676,N_6693);
nand U6981 (N_6981,N_6636,N_6608);
nand U6982 (N_6982,N_6785,N_6601);
xnor U6983 (N_6983,N_6767,N_6650);
or U6984 (N_6984,N_6748,N_6668);
nor U6985 (N_6985,N_6719,N_6761);
or U6986 (N_6986,N_6738,N_6733);
and U6987 (N_6987,N_6710,N_6699);
xnor U6988 (N_6988,N_6715,N_6726);
nor U6989 (N_6989,N_6738,N_6774);
nor U6990 (N_6990,N_6685,N_6658);
nand U6991 (N_6991,N_6601,N_6782);
and U6992 (N_6992,N_6653,N_6687);
or U6993 (N_6993,N_6625,N_6787);
nor U6994 (N_6994,N_6630,N_6793);
nor U6995 (N_6995,N_6775,N_6642);
nand U6996 (N_6996,N_6603,N_6647);
or U6997 (N_6997,N_6647,N_6641);
or U6998 (N_6998,N_6689,N_6719);
nor U6999 (N_6999,N_6629,N_6767);
nand U7000 (N_7000,N_6845,N_6909);
xnor U7001 (N_7001,N_6832,N_6842);
or U7002 (N_7002,N_6982,N_6872);
or U7003 (N_7003,N_6859,N_6864);
or U7004 (N_7004,N_6956,N_6938);
nor U7005 (N_7005,N_6904,N_6967);
or U7006 (N_7006,N_6894,N_6840);
or U7007 (N_7007,N_6922,N_6829);
or U7008 (N_7008,N_6930,N_6957);
nand U7009 (N_7009,N_6821,N_6825);
xnor U7010 (N_7010,N_6906,N_6849);
nand U7011 (N_7011,N_6885,N_6943);
nand U7012 (N_7012,N_6847,N_6959);
nand U7013 (N_7013,N_6927,N_6932);
or U7014 (N_7014,N_6946,N_6955);
nand U7015 (N_7015,N_6879,N_6949);
nand U7016 (N_7016,N_6812,N_6852);
nand U7017 (N_7017,N_6935,N_6841);
and U7018 (N_7018,N_6884,N_6961);
nor U7019 (N_7019,N_6858,N_6816);
nor U7020 (N_7020,N_6933,N_6918);
nor U7021 (N_7021,N_6815,N_6972);
nor U7022 (N_7022,N_6837,N_6910);
xor U7023 (N_7023,N_6846,N_6986);
or U7024 (N_7024,N_6834,N_6948);
xnor U7025 (N_7025,N_6907,N_6952);
xnor U7026 (N_7026,N_6809,N_6874);
or U7027 (N_7027,N_6999,N_6934);
xnor U7028 (N_7028,N_6871,N_6800);
xor U7029 (N_7029,N_6960,N_6882);
nand U7030 (N_7030,N_6903,N_6898);
xor U7031 (N_7031,N_6851,N_6855);
nand U7032 (N_7032,N_6878,N_6835);
or U7033 (N_7033,N_6875,N_6912);
or U7034 (N_7034,N_6870,N_6876);
xnor U7035 (N_7035,N_6822,N_6997);
and U7036 (N_7036,N_6813,N_6941);
or U7037 (N_7037,N_6890,N_6966);
xnor U7038 (N_7038,N_6865,N_6838);
or U7039 (N_7039,N_6989,N_6908);
nor U7040 (N_7040,N_6970,N_6839);
nor U7041 (N_7041,N_6820,N_6977);
or U7042 (N_7042,N_6811,N_6945);
nor U7043 (N_7043,N_6856,N_6901);
and U7044 (N_7044,N_6940,N_6976);
and U7045 (N_7045,N_6973,N_6857);
nor U7046 (N_7046,N_6996,N_6833);
xnor U7047 (N_7047,N_6891,N_6917);
nand U7048 (N_7048,N_6862,N_6817);
or U7049 (N_7049,N_6892,N_6867);
and U7050 (N_7050,N_6863,N_6873);
xnor U7051 (N_7051,N_6936,N_6810);
nand U7052 (N_7052,N_6896,N_6889);
nand U7053 (N_7053,N_6881,N_6861);
nor U7054 (N_7054,N_6854,N_6853);
nand U7055 (N_7055,N_6942,N_6804);
nand U7056 (N_7056,N_6803,N_6968);
or U7057 (N_7057,N_6931,N_6831);
nor U7058 (N_7058,N_6805,N_6830);
and U7059 (N_7059,N_6823,N_6979);
xor U7060 (N_7060,N_6951,N_6819);
xnor U7061 (N_7061,N_6801,N_6923);
nand U7062 (N_7062,N_6806,N_6984);
or U7063 (N_7063,N_6915,N_6939);
xor U7064 (N_7064,N_6953,N_6900);
or U7065 (N_7065,N_6808,N_6868);
or U7066 (N_7066,N_6905,N_6985);
xor U7067 (N_7067,N_6993,N_6869);
xor U7068 (N_7068,N_6998,N_6911);
xor U7069 (N_7069,N_6929,N_6887);
or U7070 (N_7070,N_6964,N_6824);
and U7071 (N_7071,N_6828,N_6947);
xor U7072 (N_7072,N_6974,N_6848);
and U7073 (N_7073,N_6924,N_6843);
or U7074 (N_7074,N_6995,N_6850);
nand U7075 (N_7075,N_6994,N_6902);
xor U7076 (N_7076,N_6844,N_6991);
and U7077 (N_7077,N_6826,N_6880);
nor U7078 (N_7078,N_6971,N_6978);
xor U7079 (N_7079,N_6866,N_6990);
and U7080 (N_7080,N_6963,N_6992);
nor U7081 (N_7081,N_6883,N_6886);
or U7082 (N_7082,N_6962,N_6913);
and U7083 (N_7083,N_6836,N_6893);
nor U7084 (N_7084,N_6807,N_6877);
and U7085 (N_7085,N_6914,N_6969);
nor U7086 (N_7086,N_6965,N_6916);
nor U7087 (N_7087,N_6954,N_6921);
xnor U7088 (N_7088,N_6944,N_6818);
xor U7089 (N_7089,N_6981,N_6827);
nor U7090 (N_7090,N_6926,N_6980);
xnor U7091 (N_7091,N_6958,N_6895);
and U7092 (N_7092,N_6899,N_6950);
nand U7093 (N_7093,N_6988,N_6928);
or U7094 (N_7094,N_6925,N_6802);
xnor U7095 (N_7095,N_6920,N_6897);
or U7096 (N_7096,N_6987,N_6983);
xnor U7097 (N_7097,N_6888,N_6814);
nor U7098 (N_7098,N_6860,N_6975);
xnor U7099 (N_7099,N_6937,N_6919);
nor U7100 (N_7100,N_6820,N_6979);
nor U7101 (N_7101,N_6829,N_6930);
nor U7102 (N_7102,N_6919,N_6853);
nor U7103 (N_7103,N_6850,N_6819);
nor U7104 (N_7104,N_6870,N_6812);
and U7105 (N_7105,N_6895,N_6929);
xnor U7106 (N_7106,N_6935,N_6951);
nand U7107 (N_7107,N_6848,N_6909);
and U7108 (N_7108,N_6984,N_6951);
nand U7109 (N_7109,N_6915,N_6809);
nor U7110 (N_7110,N_6861,N_6970);
nor U7111 (N_7111,N_6860,N_6985);
nor U7112 (N_7112,N_6986,N_6963);
nor U7113 (N_7113,N_6988,N_6964);
or U7114 (N_7114,N_6963,N_6878);
nor U7115 (N_7115,N_6836,N_6821);
and U7116 (N_7116,N_6893,N_6875);
nand U7117 (N_7117,N_6877,N_6972);
and U7118 (N_7118,N_6983,N_6925);
xnor U7119 (N_7119,N_6841,N_6973);
nor U7120 (N_7120,N_6918,N_6809);
nand U7121 (N_7121,N_6854,N_6966);
nand U7122 (N_7122,N_6911,N_6811);
xor U7123 (N_7123,N_6956,N_6993);
and U7124 (N_7124,N_6983,N_6877);
nor U7125 (N_7125,N_6914,N_6992);
xor U7126 (N_7126,N_6932,N_6901);
xnor U7127 (N_7127,N_6856,N_6995);
or U7128 (N_7128,N_6952,N_6803);
and U7129 (N_7129,N_6972,N_6947);
nor U7130 (N_7130,N_6816,N_6909);
or U7131 (N_7131,N_6878,N_6974);
xnor U7132 (N_7132,N_6870,N_6885);
or U7133 (N_7133,N_6808,N_6891);
and U7134 (N_7134,N_6919,N_6940);
or U7135 (N_7135,N_6959,N_6944);
nand U7136 (N_7136,N_6862,N_6978);
or U7137 (N_7137,N_6967,N_6998);
nand U7138 (N_7138,N_6805,N_6955);
nor U7139 (N_7139,N_6944,N_6858);
nand U7140 (N_7140,N_6901,N_6850);
xor U7141 (N_7141,N_6968,N_6926);
or U7142 (N_7142,N_6884,N_6943);
xor U7143 (N_7143,N_6877,N_6918);
and U7144 (N_7144,N_6829,N_6936);
or U7145 (N_7145,N_6936,N_6811);
or U7146 (N_7146,N_6811,N_6940);
xnor U7147 (N_7147,N_6970,N_6811);
xor U7148 (N_7148,N_6931,N_6893);
or U7149 (N_7149,N_6854,N_6805);
and U7150 (N_7150,N_6960,N_6930);
and U7151 (N_7151,N_6962,N_6822);
and U7152 (N_7152,N_6972,N_6892);
nand U7153 (N_7153,N_6907,N_6831);
or U7154 (N_7154,N_6967,N_6835);
nand U7155 (N_7155,N_6802,N_6975);
and U7156 (N_7156,N_6933,N_6997);
or U7157 (N_7157,N_6903,N_6881);
and U7158 (N_7158,N_6984,N_6882);
xor U7159 (N_7159,N_6818,N_6975);
nand U7160 (N_7160,N_6954,N_6939);
or U7161 (N_7161,N_6901,N_6808);
nand U7162 (N_7162,N_6956,N_6887);
and U7163 (N_7163,N_6924,N_6895);
xnor U7164 (N_7164,N_6878,N_6973);
and U7165 (N_7165,N_6953,N_6843);
or U7166 (N_7166,N_6819,N_6847);
and U7167 (N_7167,N_6977,N_6807);
nand U7168 (N_7168,N_6827,N_6972);
and U7169 (N_7169,N_6885,N_6852);
nor U7170 (N_7170,N_6954,N_6912);
and U7171 (N_7171,N_6857,N_6836);
nor U7172 (N_7172,N_6978,N_6980);
and U7173 (N_7173,N_6895,N_6935);
nor U7174 (N_7174,N_6931,N_6995);
and U7175 (N_7175,N_6828,N_6918);
xnor U7176 (N_7176,N_6935,N_6843);
nor U7177 (N_7177,N_6836,N_6829);
nor U7178 (N_7178,N_6999,N_6907);
or U7179 (N_7179,N_6830,N_6862);
or U7180 (N_7180,N_6941,N_6927);
nor U7181 (N_7181,N_6958,N_6918);
nand U7182 (N_7182,N_6951,N_6870);
xor U7183 (N_7183,N_6818,N_6888);
or U7184 (N_7184,N_6926,N_6869);
nand U7185 (N_7185,N_6816,N_6998);
nor U7186 (N_7186,N_6971,N_6835);
or U7187 (N_7187,N_6943,N_6833);
and U7188 (N_7188,N_6962,N_6843);
nand U7189 (N_7189,N_6921,N_6950);
or U7190 (N_7190,N_6999,N_6901);
xor U7191 (N_7191,N_6899,N_6914);
xnor U7192 (N_7192,N_6953,N_6930);
and U7193 (N_7193,N_6992,N_6910);
or U7194 (N_7194,N_6895,N_6826);
or U7195 (N_7195,N_6945,N_6890);
or U7196 (N_7196,N_6984,N_6960);
nand U7197 (N_7197,N_6890,N_6918);
xnor U7198 (N_7198,N_6976,N_6804);
and U7199 (N_7199,N_6954,N_6845);
xor U7200 (N_7200,N_7035,N_7195);
or U7201 (N_7201,N_7047,N_7132);
xor U7202 (N_7202,N_7015,N_7151);
nand U7203 (N_7203,N_7192,N_7154);
and U7204 (N_7204,N_7032,N_7084);
nand U7205 (N_7205,N_7169,N_7105);
nor U7206 (N_7206,N_7116,N_7155);
nand U7207 (N_7207,N_7076,N_7070);
or U7208 (N_7208,N_7001,N_7189);
nand U7209 (N_7209,N_7174,N_7172);
nand U7210 (N_7210,N_7038,N_7009);
nand U7211 (N_7211,N_7100,N_7118);
nand U7212 (N_7212,N_7111,N_7078);
and U7213 (N_7213,N_7050,N_7115);
xor U7214 (N_7214,N_7020,N_7041);
or U7215 (N_7215,N_7058,N_7170);
nand U7216 (N_7216,N_7046,N_7109);
nand U7217 (N_7217,N_7194,N_7044);
nand U7218 (N_7218,N_7068,N_7081);
or U7219 (N_7219,N_7176,N_7030);
xor U7220 (N_7220,N_7167,N_7080);
nand U7221 (N_7221,N_7177,N_7075);
or U7222 (N_7222,N_7137,N_7086);
or U7223 (N_7223,N_7135,N_7171);
nand U7224 (N_7224,N_7114,N_7130);
xnor U7225 (N_7225,N_7049,N_7007);
nor U7226 (N_7226,N_7051,N_7102);
xor U7227 (N_7227,N_7011,N_7063);
xor U7228 (N_7228,N_7085,N_7064);
and U7229 (N_7229,N_7018,N_7168);
nor U7230 (N_7230,N_7042,N_7197);
xnor U7231 (N_7231,N_7184,N_7056);
nor U7232 (N_7232,N_7134,N_7092);
nand U7233 (N_7233,N_7074,N_7128);
xor U7234 (N_7234,N_7185,N_7125);
nor U7235 (N_7235,N_7048,N_7071);
and U7236 (N_7236,N_7065,N_7120);
and U7237 (N_7237,N_7196,N_7161);
and U7238 (N_7238,N_7014,N_7067);
and U7239 (N_7239,N_7026,N_7123);
and U7240 (N_7240,N_7158,N_7156);
or U7241 (N_7241,N_7052,N_7149);
nand U7242 (N_7242,N_7000,N_7082);
and U7243 (N_7243,N_7054,N_7037);
and U7244 (N_7244,N_7173,N_7140);
nand U7245 (N_7245,N_7033,N_7040);
xor U7246 (N_7246,N_7147,N_7142);
or U7247 (N_7247,N_7010,N_7098);
or U7248 (N_7248,N_7089,N_7164);
and U7249 (N_7249,N_7053,N_7160);
nand U7250 (N_7250,N_7097,N_7159);
and U7251 (N_7251,N_7126,N_7193);
and U7252 (N_7252,N_7023,N_7017);
and U7253 (N_7253,N_7028,N_7110);
and U7254 (N_7254,N_7066,N_7107);
nor U7255 (N_7255,N_7165,N_7183);
and U7256 (N_7256,N_7122,N_7162);
and U7257 (N_7257,N_7005,N_7153);
xnor U7258 (N_7258,N_7055,N_7104);
or U7259 (N_7259,N_7190,N_7036);
nor U7260 (N_7260,N_7141,N_7127);
or U7261 (N_7261,N_7124,N_7094);
xor U7262 (N_7262,N_7191,N_7131);
nor U7263 (N_7263,N_7088,N_7182);
nor U7264 (N_7264,N_7083,N_7166);
or U7265 (N_7265,N_7003,N_7025);
or U7266 (N_7266,N_7006,N_7039);
and U7267 (N_7267,N_7133,N_7199);
nor U7268 (N_7268,N_7146,N_7144);
or U7269 (N_7269,N_7060,N_7180);
nand U7270 (N_7270,N_7119,N_7057);
xnor U7271 (N_7271,N_7093,N_7101);
or U7272 (N_7272,N_7034,N_7077);
xnor U7273 (N_7273,N_7148,N_7016);
nor U7274 (N_7274,N_7113,N_7073);
nand U7275 (N_7275,N_7103,N_7008);
or U7276 (N_7276,N_7027,N_7029);
or U7277 (N_7277,N_7112,N_7198);
and U7278 (N_7278,N_7186,N_7062);
nand U7279 (N_7279,N_7150,N_7019);
or U7280 (N_7280,N_7002,N_7139);
or U7281 (N_7281,N_7045,N_7090);
xnor U7282 (N_7282,N_7072,N_7012);
xnor U7283 (N_7283,N_7099,N_7152);
nand U7284 (N_7284,N_7108,N_7059);
and U7285 (N_7285,N_7079,N_7031);
and U7286 (N_7286,N_7129,N_7138);
xor U7287 (N_7287,N_7022,N_7121);
xor U7288 (N_7288,N_7179,N_7024);
nor U7289 (N_7289,N_7021,N_7043);
xor U7290 (N_7290,N_7004,N_7091);
and U7291 (N_7291,N_7163,N_7136);
xor U7292 (N_7292,N_7178,N_7145);
and U7293 (N_7293,N_7143,N_7175);
nand U7294 (N_7294,N_7106,N_7117);
nor U7295 (N_7295,N_7181,N_7095);
xnor U7296 (N_7296,N_7157,N_7187);
xnor U7297 (N_7297,N_7188,N_7069);
and U7298 (N_7298,N_7013,N_7087);
or U7299 (N_7299,N_7096,N_7061);
or U7300 (N_7300,N_7104,N_7192);
nand U7301 (N_7301,N_7150,N_7170);
xor U7302 (N_7302,N_7180,N_7099);
and U7303 (N_7303,N_7087,N_7080);
xnor U7304 (N_7304,N_7079,N_7169);
and U7305 (N_7305,N_7109,N_7146);
nand U7306 (N_7306,N_7162,N_7002);
xnor U7307 (N_7307,N_7012,N_7167);
or U7308 (N_7308,N_7110,N_7128);
and U7309 (N_7309,N_7102,N_7002);
xor U7310 (N_7310,N_7092,N_7037);
and U7311 (N_7311,N_7142,N_7099);
nor U7312 (N_7312,N_7033,N_7106);
or U7313 (N_7313,N_7018,N_7176);
xnor U7314 (N_7314,N_7177,N_7108);
xnor U7315 (N_7315,N_7108,N_7094);
xor U7316 (N_7316,N_7093,N_7188);
and U7317 (N_7317,N_7090,N_7018);
nand U7318 (N_7318,N_7185,N_7176);
or U7319 (N_7319,N_7022,N_7014);
nor U7320 (N_7320,N_7074,N_7065);
xnor U7321 (N_7321,N_7025,N_7183);
and U7322 (N_7322,N_7153,N_7032);
nor U7323 (N_7323,N_7056,N_7169);
nand U7324 (N_7324,N_7027,N_7007);
nand U7325 (N_7325,N_7012,N_7009);
xor U7326 (N_7326,N_7178,N_7116);
or U7327 (N_7327,N_7072,N_7118);
or U7328 (N_7328,N_7136,N_7177);
xor U7329 (N_7329,N_7092,N_7094);
and U7330 (N_7330,N_7027,N_7041);
xor U7331 (N_7331,N_7180,N_7127);
or U7332 (N_7332,N_7122,N_7001);
xnor U7333 (N_7333,N_7065,N_7140);
nand U7334 (N_7334,N_7168,N_7114);
nor U7335 (N_7335,N_7147,N_7008);
nor U7336 (N_7336,N_7192,N_7064);
or U7337 (N_7337,N_7050,N_7056);
xnor U7338 (N_7338,N_7158,N_7014);
nand U7339 (N_7339,N_7180,N_7024);
and U7340 (N_7340,N_7110,N_7004);
xnor U7341 (N_7341,N_7118,N_7152);
nand U7342 (N_7342,N_7068,N_7190);
or U7343 (N_7343,N_7190,N_7183);
or U7344 (N_7344,N_7137,N_7185);
and U7345 (N_7345,N_7130,N_7066);
and U7346 (N_7346,N_7163,N_7151);
and U7347 (N_7347,N_7099,N_7041);
or U7348 (N_7348,N_7162,N_7103);
nand U7349 (N_7349,N_7055,N_7008);
nand U7350 (N_7350,N_7046,N_7176);
xnor U7351 (N_7351,N_7031,N_7083);
xor U7352 (N_7352,N_7031,N_7047);
nor U7353 (N_7353,N_7114,N_7188);
or U7354 (N_7354,N_7019,N_7049);
xnor U7355 (N_7355,N_7071,N_7189);
nor U7356 (N_7356,N_7187,N_7030);
and U7357 (N_7357,N_7067,N_7072);
nor U7358 (N_7358,N_7098,N_7146);
nor U7359 (N_7359,N_7082,N_7056);
or U7360 (N_7360,N_7089,N_7022);
nand U7361 (N_7361,N_7068,N_7182);
or U7362 (N_7362,N_7161,N_7088);
and U7363 (N_7363,N_7164,N_7172);
or U7364 (N_7364,N_7171,N_7154);
xor U7365 (N_7365,N_7196,N_7110);
or U7366 (N_7366,N_7113,N_7001);
nand U7367 (N_7367,N_7111,N_7048);
and U7368 (N_7368,N_7134,N_7048);
nor U7369 (N_7369,N_7133,N_7060);
nand U7370 (N_7370,N_7053,N_7033);
xnor U7371 (N_7371,N_7182,N_7091);
and U7372 (N_7372,N_7184,N_7072);
nor U7373 (N_7373,N_7146,N_7182);
and U7374 (N_7374,N_7031,N_7134);
and U7375 (N_7375,N_7124,N_7040);
nor U7376 (N_7376,N_7010,N_7142);
nor U7377 (N_7377,N_7055,N_7147);
and U7378 (N_7378,N_7122,N_7003);
or U7379 (N_7379,N_7180,N_7146);
nand U7380 (N_7380,N_7117,N_7161);
xnor U7381 (N_7381,N_7126,N_7107);
xor U7382 (N_7382,N_7112,N_7007);
xor U7383 (N_7383,N_7140,N_7181);
nand U7384 (N_7384,N_7199,N_7117);
or U7385 (N_7385,N_7062,N_7191);
and U7386 (N_7386,N_7013,N_7149);
nand U7387 (N_7387,N_7173,N_7167);
and U7388 (N_7388,N_7137,N_7089);
nand U7389 (N_7389,N_7007,N_7117);
xor U7390 (N_7390,N_7028,N_7019);
or U7391 (N_7391,N_7024,N_7195);
xnor U7392 (N_7392,N_7021,N_7186);
and U7393 (N_7393,N_7047,N_7089);
or U7394 (N_7394,N_7191,N_7156);
nand U7395 (N_7395,N_7077,N_7173);
nand U7396 (N_7396,N_7019,N_7094);
nand U7397 (N_7397,N_7158,N_7057);
nor U7398 (N_7398,N_7050,N_7183);
nor U7399 (N_7399,N_7000,N_7199);
or U7400 (N_7400,N_7269,N_7353);
nor U7401 (N_7401,N_7320,N_7387);
nand U7402 (N_7402,N_7367,N_7231);
nand U7403 (N_7403,N_7297,N_7270);
and U7404 (N_7404,N_7335,N_7207);
nand U7405 (N_7405,N_7379,N_7315);
xor U7406 (N_7406,N_7397,N_7252);
and U7407 (N_7407,N_7308,N_7212);
nor U7408 (N_7408,N_7238,N_7220);
and U7409 (N_7409,N_7321,N_7339);
nor U7410 (N_7410,N_7338,N_7386);
and U7411 (N_7411,N_7332,N_7323);
or U7412 (N_7412,N_7259,N_7377);
nand U7413 (N_7413,N_7368,N_7225);
nand U7414 (N_7414,N_7241,N_7245);
or U7415 (N_7415,N_7200,N_7262);
nand U7416 (N_7416,N_7279,N_7214);
nor U7417 (N_7417,N_7360,N_7283);
or U7418 (N_7418,N_7282,N_7322);
and U7419 (N_7419,N_7209,N_7345);
and U7420 (N_7420,N_7330,N_7389);
nand U7421 (N_7421,N_7233,N_7374);
nor U7422 (N_7422,N_7266,N_7364);
and U7423 (N_7423,N_7277,N_7268);
nand U7424 (N_7424,N_7357,N_7208);
and U7425 (N_7425,N_7300,N_7340);
nand U7426 (N_7426,N_7327,N_7329);
xor U7427 (N_7427,N_7358,N_7244);
nor U7428 (N_7428,N_7234,N_7254);
or U7429 (N_7429,N_7264,N_7346);
nor U7430 (N_7430,N_7230,N_7304);
nor U7431 (N_7431,N_7267,N_7210);
nor U7432 (N_7432,N_7363,N_7236);
and U7433 (N_7433,N_7394,N_7351);
or U7434 (N_7434,N_7355,N_7347);
nand U7435 (N_7435,N_7348,N_7301);
or U7436 (N_7436,N_7295,N_7365);
or U7437 (N_7437,N_7296,N_7224);
nand U7438 (N_7438,N_7393,N_7253);
nand U7439 (N_7439,N_7285,N_7219);
or U7440 (N_7440,N_7384,N_7328);
nor U7441 (N_7441,N_7293,N_7204);
nor U7442 (N_7442,N_7286,N_7292);
nand U7443 (N_7443,N_7284,N_7222);
nand U7444 (N_7444,N_7276,N_7337);
nor U7445 (N_7445,N_7336,N_7274);
xnor U7446 (N_7446,N_7318,N_7399);
and U7447 (N_7447,N_7309,N_7359);
nor U7448 (N_7448,N_7350,N_7215);
nand U7449 (N_7449,N_7344,N_7362);
nor U7450 (N_7450,N_7278,N_7202);
nor U7451 (N_7451,N_7246,N_7263);
and U7452 (N_7452,N_7343,N_7294);
nor U7453 (N_7453,N_7203,N_7319);
nor U7454 (N_7454,N_7361,N_7213);
xnor U7455 (N_7455,N_7395,N_7206);
xor U7456 (N_7456,N_7317,N_7272);
or U7457 (N_7457,N_7251,N_7299);
or U7458 (N_7458,N_7232,N_7242);
or U7459 (N_7459,N_7305,N_7229);
and U7460 (N_7460,N_7291,N_7260);
xnor U7461 (N_7461,N_7290,N_7227);
xnor U7462 (N_7462,N_7342,N_7324);
nand U7463 (N_7463,N_7280,N_7366);
or U7464 (N_7464,N_7221,N_7239);
nand U7465 (N_7465,N_7352,N_7275);
nor U7466 (N_7466,N_7311,N_7298);
or U7467 (N_7467,N_7256,N_7257);
xnor U7468 (N_7468,N_7211,N_7341);
and U7469 (N_7469,N_7381,N_7388);
nor U7470 (N_7470,N_7261,N_7314);
or U7471 (N_7471,N_7240,N_7372);
or U7472 (N_7472,N_7306,N_7334);
and U7473 (N_7473,N_7243,N_7307);
or U7474 (N_7474,N_7356,N_7250);
or U7475 (N_7475,N_7302,N_7325);
nor U7476 (N_7476,N_7380,N_7396);
or U7477 (N_7477,N_7287,N_7201);
nor U7478 (N_7478,N_7281,N_7235);
and U7479 (N_7479,N_7237,N_7216);
nor U7480 (N_7480,N_7369,N_7265);
xor U7481 (N_7481,N_7218,N_7312);
or U7482 (N_7482,N_7383,N_7392);
nand U7483 (N_7483,N_7313,N_7289);
nand U7484 (N_7484,N_7248,N_7217);
or U7485 (N_7485,N_7373,N_7273);
nand U7486 (N_7486,N_7316,N_7288);
or U7487 (N_7487,N_7391,N_7249);
xor U7488 (N_7488,N_7398,N_7228);
or U7489 (N_7489,N_7370,N_7371);
xor U7490 (N_7490,N_7258,N_7376);
or U7491 (N_7491,N_7205,N_7333);
nand U7492 (N_7492,N_7331,N_7271);
or U7493 (N_7493,N_7378,N_7247);
xnor U7494 (N_7494,N_7390,N_7226);
and U7495 (N_7495,N_7223,N_7385);
xnor U7496 (N_7496,N_7349,N_7375);
xnor U7497 (N_7497,N_7382,N_7255);
xnor U7498 (N_7498,N_7354,N_7326);
nor U7499 (N_7499,N_7310,N_7303);
xnor U7500 (N_7500,N_7365,N_7375);
nor U7501 (N_7501,N_7374,N_7217);
and U7502 (N_7502,N_7399,N_7276);
nor U7503 (N_7503,N_7294,N_7360);
nor U7504 (N_7504,N_7281,N_7317);
or U7505 (N_7505,N_7318,N_7204);
and U7506 (N_7506,N_7374,N_7230);
or U7507 (N_7507,N_7369,N_7384);
nor U7508 (N_7508,N_7319,N_7391);
nor U7509 (N_7509,N_7263,N_7378);
nor U7510 (N_7510,N_7267,N_7298);
and U7511 (N_7511,N_7250,N_7345);
or U7512 (N_7512,N_7269,N_7305);
xor U7513 (N_7513,N_7302,N_7318);
nor U7514 (N_7514,N_7241,N_7364);
nand U7515 (N_7515,N_7384,N_7262);
and U7516 (N_7516,N_7208,N_7314);
and U7517 (N_7517,N_7307,N_7368);
or U7518 (N_7518,N_7341,N_7363);
and U7519 (N_7519,N_7230,N_7285);
xnor U7520 (N_7520,N_7272,N_7220);
or U7521 (N_7521,N_7255,N_7296);
and U7522 (N_7522,N_7392,N_7324);
or U7523 (N_7523,N_7319,N_7220);
nand U7524 (N_7524,N_7286,N_7387);
and U7525 (N_7525,N_7275,N_7311);
or U7526 (N_7526,N_7214,N_7278);
xnor U7527 (N_7527,N_7288,N_7319);
xnor U7528 (N_7528,N_7326,N_7276);
xor U7529 (N_7529,N_7333,N_7387);
and U7530 (N_7530,N_7230,N_7332);
nor U7531 (N_7531,N_7274,N_7373);
or U7532 (N_7532,N_7375,N_7228);
and U7533 (N_7533,N_7397,N_7361);
xor U7534 (N_7534,N_7361,N_7277);
and U7535 (N_7535,N_7282,N_7326);
nor U7536 (N_7536,N_7215,N_7313);
nor U7537 (N_7537,N_7353,N_7241);
xor U7538 (N_7538,N_7272,N_7347);
or U7539 (N_7539,N_7358,N_7320);
or U7540 (N_7540,N_7378,N_7269);
xnor U7541 (N_7541,N_7295,N_7346);
nand U7542 (N_7542,N_7385,N_7269);
nand U7543 (N_7543,N_7290,N_7346);
and U7544 (N_7544,N_7348,N_7335);
nor U7545 (N_7545,N_7219,N_7261);
or U7546 (N_7546,N_7371,N_7395);
nand U7547 (N_7547,N_7303,N_7203);
and U7548 (N_7548,N_7399,N_7248);
nor U7549 (N_7549,N_7341,N_7290);
nand U7550 (N_7550,N_7306,N_7210);
nand U7551 (N_7551,N_7299,N_7303);
and U7552 (N_7552,N_7362,N_7363);
nand U7553 (N_7553,N_7360,N_7314);
xor U7554 (N_7554,N_7200,N_7359);
nand U7555 (N_7555,N_7241,N_7355);
and U7556 (N_7556,N_7238,N_7246);
nor U7557 (N_7557,N_7216,N_7309);
or U7558 (N_7558,N_7324,N_7207);
xnor U7559 (N_7559,N_7366,N_7371);
xor U7560 (N_7560,N_7298,N_7331);
or U7561 (N_7561,N_7254,N_7385);
nor U7562 (N_7562,N_7370,N_7292);
or U7563 (N_7563,N_7396,N_7264);
nor U7564 (N_7564,N_7223,N_7254);
nor U7565 (N_7565,N_7228,N_7283);
nand U7566 (N_7566,N_7206,N_7260);
nor U7567 (N_7567,N_7212,N_7238);
xor U7568 (N_7568,N_7394,N_7303);
and U7569 (N_7569,N_7309,N_7211);
and U7570 (N_7570,N_7256,N_7298);
xnor U7571 (N_7571,N_7351,N_7211);
xnor U7572 (N_7572,N_7326,N_7313);
and U7573 (N_7573,N_7232,N_7395);
and U7574 (N_7574,N_7314,N_7348);
and U7575 (N_7575,N_7209,N_7305);
nand U7576 (N_7576,N_7364,N_7382);
and U7577 (N_7577,N_7305,N_7376);
and U7578 (N_7578,N_7248,N_7323);
nor U7579 (N_7579,N_7216,N_7203);
xnor U7580 (N_7580,N_7216,N_7398);
nor U7581 (N_7581,N_7204,N_7241);
nor U7582 (N_7582,N_7323,N_7377);
and U7583 (N_7583,N_7351,N_7250);
nand U7584 (N_7584,N_7361,N_7239);
or U7585 (N_7585,N_7249,N_7321);
xnor U7586 (N_7586,N_7360,N_7370);
xor U7587 (N_7587,N_7372,N_7233);
xor U7588 (N_7588,N_7381,N_7277);
nand U7589 (N_7589,N_7314,N_7342);
and U7590 (N_7590,N_7397,N_7318);
and U7591 (N_7591,N_7273,N_7229);
nand U7592 (N_7592,N_7307,N_7316);
nor U7593 (N_7593,N_7314,N_7244);
nor U7594 (N_7594,N_7213,N_7230);
and U7595 (N_7595,N_7287,N_7327);
nand U7596 (N_7596,N_7344,N_7388);
and U7597 (N_7597,N_7253,N_7348);
or U7598 (N_7598,N_7254,N_7380);
or U7599 (N_7599,N_7265,N_7348);
nor U7600 (N_7600,N_7482,N_7539);
nor U7601 (N_7601,N_7407,N_7544);
and U7602 (N_7602,N_7439,N_7444);
and U7603 (N_7603,N_7453,N_7477);
xnor U7604 (N_7604,N_7467,N_7465);
or U7605 (N_7605,N_7584,N_7529);
or U7606 (N_7606,N_7469,N_7510);
xnor U7607 (N_7607,N_7526,N_7521);
or U7608 (N_7608,N_7530,N_7400);
and U7609 (N_7609,N_7590,N_7473);
nor U7610 (N_7610,N_7440,N_7492);
nand U7611 (N_7611,N_7426,N_7497);
nor U7612 (N_7612,N_7511,N_7423);
and U7613 (N_7613,N_7401,N_7564);
nor U7614 (N_7614,N_7577,N_7522);
nor U7615 (N_7615,N_7496,N_7468);
and U7616 (N_7616,N_7517,N_7456);
nand U7617 (N_7617,N_7498,N_7472);
xnor U7618 (N_7618,N_7520,N_7528);
nor U7619 (N_7619,N_7422,N_7459);
nor U7620 (N_7620,N_7514,N_7425);
nand U7621 (N_7621,N_7452,N_7420);
nand U7622 (N_7622,N_7479,N_7515);
nand U7623 (N_7623,N_7556,N_7489);
nor U7624 (N_7624,N_7484,N_7445);
or U7625 (N_7625,N_7437,N_7432);
or U7626 (N_7626,N_7527,N_7474);
nand U7627 (N_7627,N_7443,N_7536);
nor U7628 (N_7628,N_7503,N_7416);
or U7629 (N_7629,N_7586,N_7480);
nand U7630 (N_7630,N_7562,N_7413);
or U7631 (N_7631,N_7403,N_7500);
and U7632 (N_7632,N_7424,N_7570);
nand U7633 (N_7633,N_7419,N_7567);
xor U7634 (N_7634,N_7561,N_7417);
nand U7635 (N_7635,N_7523,N_7580);
or U7636 (N_7636,N_7576,N_7595);
nor U7637 (N_7637,N_7411,N_7588);
xnor U7638 (N_7638,N_7463,N_7441);
nand U7639 (N_7639,N_7585,N_7483);
and U7640 (N_7640,N_7534,N_7505);
or U7641 (N_7641,N_7504,N_7462);
and U7642 (N_7642,N_7475,N_7435);
nor U7643 (N_7643,N_7507,N_7540);
or U7644 (N_7644,N_7560,N_7518);
nor U7645 (N_7645,N_7438,N_7478);
and U7646 (N_7646,N_7458,N_7538);
or U7647 (N_7647,N_7555,N_7592);
and U7648 (N_7648,N_7583,N_7558);
and U7649 (N_7649,N_7549,N_7554);
and U7650 (N_7650,N_7430,N_7410);
and U7651 (N_7651,N_7559,N_7557);
nor U7652 (N_7652,N_7481,N_7446);
nand U7653 (N_7653,N_7545,N_7448);
nor U7654 (N_7654,N_7594,N_7541);
or U7655 (N_7655,N_7593,N_7499);
xnor U7656 (N_7656,N_7506,N_7442);
nand U7657 (N_7657,N_7551,N_7535);
nor U7658 (N_7658,N_7431,N_7404);
or U7659 (N_7659,N_7454,N_7508);
nor U7660 (N_7660,N_7524,N_7405);
nor U7661 (N_7661,N_7546,N_7563);
nand U7662 (N_7662,N_7485,N_7457);
nor U7663 (N_7663,N_7495,N_7414);
nor U7664 (N_7664,N_7493,N_7571);
and U7665 (N_7665,N_7532,N_7550);
nor U7666 (N_7666,N_7537,N_7449);
nor U7667 (N_7667,N_7525,N_7533);
nand U7668 (N_7668,N_7568,N_7409);
xnor U7669 (N_7669,N_7406,N_7589);
nor U7670 (N_7670,N_7450,N_7587);
nor U7671 (N_7671,N_7548,N_7408);
xor U7672 (N_7672,N_7569,N_7573);
nor U7673 (N_7673,N_7491,N_7470);
nor U7674 (N_7674,N_7427,N_7579);
or U7675 (N_7675,N_7466,N_7531);
nor U7676 (N_7676,N_7476,N_7494);
nand U7677 (N_7677,N_7565,N_7542);
xnor U7678 (N_7678,N_7421,N_7578);
xor U7679 (N_7679,N_7402,N_7460);
nand U7680 (N_7680,N_7487,N_7434);
and U7681 (N_7681,N_7433,N_7572);
nor U7682 (N_7682,N_7552,N_7581);
xor U7683 (N_7683,N_7464,N_7513);
or U7684 (N_7684,N_7543,N_7436);
xor U7685 (N_7685,N_7509,N_7566);
and U7686 (N_7686,N_7447,N_7461);
xor U7687 (N_7687,N_7501,N_7428);
xor U7688 (N_7688,N_7471,N_7429);
nand U7689 (N_7689,N_7553,N_7596);
nand U7690 (N_7690,N_7516,N_7490);
or U7691 (N_7691,N_7598,N_7519);
xnor U7692 (N_7692,N_7488,N_7591);
xor U7693 (N_7693,N_7415,N_7512);
xnor U7694 (N_7694,N_7575,N_7597);
xnor U7695 (N_7695,N_7486,N_7418);
nand U7696 (N_7696,N_7547,N_7599);
nand U7697 (N_7697,N_7455,N_7582);
xnor U7698 (N_7698,N_7412,N_7451);
and U7699 (N_7699,N_7574,N_7502);
xnor U7700 (N_7700,N_7498,N_7516);
xnor U7701 (N_7701,N_7597,N_7450);
xnor U7702 (N_7702,N_7455,N_7523);
or U7703 (N_7703,N_7427,N_7549);
nand U7704 (N_7704,N_7414,N_7405);
xor U7705 (N_7705,N_7490,N_7572);
nand U7706 (N_7706,N_7477,N_7406);
nor U7707 (N_7707,N_7472,N_7504);
or U7708 (N_7708,N_7409,N_7510);
and U7709 (N_7709,N_7599,N_7406);
and U7710 (N_7710,N_7502,N_7408);
nand U7711 (N_7711,N_7478,N_7401);
nand U7712 (N_7712,N_7412,N_7437);
xor U7713 (N_7713,N_7497,N_7492);
nor U7714 (N_7714,N_7403,N_7593);
xnor U7715 (N_7715,N_7530,N_7465);
nand U7716 (N_7716,N_7402,N_7475);
nor U7717 (N_7717,N_7590,N_7450);
xnor U7718 (N_7718,N_7425,N_7536);
and U7719 (N_7719,N_7429,N_7420);
nor U7720 (N_7720,N_7471,N_7510);
and U7721 (N_7721,N_7557,N_7466);
and U7722 (N_7722,N_7551,N_7426);
or U7723 (N_7723,N_7515,N_7586);
nand U7724 (N_7724,N_7487,N_7551);
nand U7725 (N_7725,N_7523,N_7546);
nor U7726 (N_7726,N_7425,N_7541);
and U7727 (N_7727,N_7436,N_7531);
or U7728 (N_7728,N_7448,N_7411);
and U7729 (N_7729,N_7406,N_7463);
or U7730 (N_7730,N_7555,N_7509);
xnor U7731 (N_7731,N_7479,N_7463);
nand U7732 (N_7732,N_7575,N_7429);
or U7733 (N_7733,N_7494,N_7507);
xnor U7734 (N_7734,N_7570,N_7404);
nor U7735 (N_7735,N_7403,N_7524);
xnor U7736 (N_7736,N_7421,N_7567);
or U7737 (N_7737,N_7438,N_7546);
nand U7738 (N_7738,N_7553,N_7489);
and U7739 (N_7739,N_7489,N_7485);
and U7740 (N_7740,N_7461,N_7460);
and U7741 (N_7741,N_7426,N_7562);
or U7742 (N_7742,N_7590,N_7583);
xor U7743 (N_7743,N_7580,N_7587);
nor U7744 (N_7744,N_7491,N_7502);
nand U7745 (N_7745,N_7439,N_7487);
nor U7746 (N_7746,N_7472,N_7494);
nand U7747 (N_7747,N_7593,N_7443);
nand U7748 (N_7748,N_7573,N_7483);
nand U7749 (N_7749,N_7460,N_7450);
xor U7750 (N_7750,N_7407,N_7417);
or U7751 (N_7751,N_7560,N_7410);
or U7752 (N_7752,N_7532,N_7409);
xnor U7753 (N_7753,N_7436,N_7549);
and U7754 (N_7754,N_7449,N_7457);
and U7755 (N_7755,N_7573,N_7442);
or U7756 (N_7756,N_7526,N_7466);
nor U7757 (N_7757,N_7525,N_7598);
xor U7758 (N_7758,N_7492,N_7571);
nand U7759 (N_7759,N_7404,N_7503);
xnor U7760 (N_7760,N_7460,N_7502);
xnor U7761 (N_7761,N_7476,N_7522);
xnor U7762 (N_7762,N_7515,N_7522);
nand U7763 (N_7763,N_7518,N_7429);
nand U7764 (N_7764,N_7557,N_7427);
nand U7765 (N_7765,N_7504,N_7522);
and U7766 (N_7766,N_7511,N_7515);
nor U7767 (N_7767,N_7495,N_7515);
nor U7768 (N_7768,N_7558,N_7425);
or U7769 (N_7769,N_7574,N_7504);
xor U7770 (N_7770,N_7508,N_7550);
or U7771 (N_7771,N_7562,N_7434);
nand U7772 (N_7772,N_7417,N_7501);
xnor U7773 (N_7773,N_7511,N_7594);
xnor U7774 (N_7774,N_7562,N_7469);
nand U7775 (N_7775,N_7492,N_7500);
nand U7776 (N_7776,N_7471,N_7591);
or U7777 (N_7777,N_7475,N_7443);
nor U7778 (N_7778,N_7405,N_7447);
nand U7779 (N_7779,N_7562,N_7527);
or U7780 (N_7780,N_7567,N_7474);
nor U7781 (N_7781,N_7553,N_7486);
or U7782 (N_7782,N_7537,N_7483);
and U7783 (N_7783,N_7413,N_7544);
or U7784 (N_7784,N_7557,N_7443);
nor U7785 (N_7785,N_7592,N_7421);
nor U7786 (N_7786,N_7556,N_7577);
and U7787 (N_7787,N_7587,N_7495);
or U7788 (N_7788,N_7413,N_7496);
xnor U7789 (N_7789,N_7584,N_7507);
xor U7790 (N_7790,N_7458,N_7485);
and U7791 (N_7791,N_7499,N_7559);
nor U7792 (N_7792,N_7463,N_7549);
xor U7793 (N_7793,N_7430,N_7536);
nand U7794 (N_7794,N_7542,N_7548);
xor U7795 (N_7795,N_7440,N_7493);
xnor U7796 (N_7796,N_7535,N_7532);
nor U7797 (N_7797,N_7525,N_7440);
nor U7798 (N_7798,N_7592,N_7414);
and U7799 (N_7799,N_7597,N_7487);
and U7800 (N_7800,N_7618,N_7760);
or U7801 (N_7801,N_7725,N_7780);
xor U7802 (N_7802,N_7674,N_7792);
and U7803 (N_7803,N_7765,N_7716);
or U7804 (N_7804,N_7676,N_7604);
nand U7805 (N_7805,N_7677,N_7634);
or U7806 (N_7806,N_7661,N_7663);
and U7807 (N_7807,N_7646,N_7686);
xor U7808 (N_7808,N_7684,N_7770);
or U7809 (N_7809,N_7789,N_7723);
nand U7810 (N_7810,N_7621,N_7795);
or U7811 (N_7811,N_7701,N_7797);
xor U7812 (N_7812,N_7679,N_7712);
xor U7813 (N_7813,N_7670,N_7731);
nor U7814 (N_7814,N_7707,N_7666);
nor U7815 (N_7815,N_7662,N_7703);
and U7816 (N_7816,N_7757,N_7654);
and U7817 (N_7817,N_7743,N_7776);
and U7818 (N_7818,N_7706,N_7798);
or U7819 (N_7819,N_7788,N_7733);
xnor U7820 (N_7820,N_7614,N_7779);
or U7821 (N_7821,N_7615,N_7715);
nand U7822 (N_7822,N_7741,N_7652);
xor U7823 (N_7823,N_7740,N_7695);
xnor U7824 (N_7824,N_7685,N_7632);
nor U7825 (N_7825,N_7708,N_7696);
and U7826 (N_7826,N_7787,N_7625);
nand U7827 (N_7827,N_7688,N_7600);
or U7828 (N_7828,N_7612,N_7642);
xnor U7829 (N_7829,N_7605,N_7705);
and U7830 (N_7830,N_7758,N_7766);
or U7831 (N_7831,N_7774,N_7735);
xnor U7832 (N_7832,N_7683,N_7637);
xor U7833 (N_7833,N_7647,N_7610);
nand U7834 (N_7834,N_7692,N_7781);
nor U7835 (N_7835,N_7636,N_7764);
nor U7836 (N_7836,N_7622,N_7665);
xnor U7837 (N_7837,N_7656,N_7777);
nor U7838 (N_7838,N_7775,N_7624);
nand U7839 (N_7839,N_7773,N_7623);
nor U7840 (N_7840,N_7672,N_7710);
nand U7841 (N_7841,N_7738,N_7671);
xnor U7842 (N_7842,N_7633,N_7609);
xor U7843 (N_7843,N_7724,N_7644);
nand U7844 (N_7844,N_7611,N_7606);
xor U7845 (N_7845,N_7627,N_7645);
and U7846 (N_7846,N_7713,N_7700);
or U7847 (N_7847,N_7745,N_7619);
nand U7848 (N_7848,N_7720,N_7796);
nor U7849 (N_7849,N_7640,N_7727);
xnor U7850 (N_7850,N_7754,N_7659);
and U7851 (N_7851,N_7709,N_7768);
or U7852 (N_7852,N_7783,N_7730);
and U7853 (N_7853,N_7699,N_7697);
or U7854 (N_7854,N_7772,N_7613);
nand U7855 (N_7855,N_7602,N_7739);
xnor U7856 (N_7856,N_7667,N_7680);
or U7857 (N_7857,N_7753,N_7687);
and U7858 (N_7858,N_7658,N_7689);
and U7859 (N_7859,N_7755,N_7722);
nor U7860 (N_7860,N_7762,N_7732);
and U7861 (N_7861,N_7601,N_7691);
xnor U7862 (N_7862,N_7750,N_7721);
xor U7863 (N_7863,N_7748,N_7734);
xnor U7864 (N_7864,N_7607,N_7669);
or U7865 (N_7865,N_7608,N_7698);
nand U7866 (N_7866,N_7648,N_7630);
nand U7867 (N_7867,N_7704,N_7769);
nand U7868 (N_7868,N_7714,N_7744);
nor U7869 (N_7869,N_7681,N_7759);
nand U7870 (N_7870,N_7690,N_7617);
xnor U7871 (N_7871,N_7719,N_7751);
nand U7872 (N_7872,N_7664,N_7767);
and U7873 (N_7873,N_7694,N_7702);
and U7874 (N_7874,N_7749,N_7717);
and U7875 (N_7875,N_7786,N_7657);
or U7876 (N_7876,N_7616,N_7675);
nor U7877 (N_7877,N_7660,N_7673);
and U7878 (N_7878,N_7643,N_7628);
and U7879 (N_7879,N_7631,N_7693);
nor U7880 (N_7880,N_7747,N_7639);
or U7881 (N_7881,N_7729,N_7799);
nor U7882 (N_7882,N_7668,N_7771);
or U7883 (N_7883,N_7782,N_7785);
or U7884 (N_7884,N_7784,N_7678);
and U7885 (N_7885,N_7737,N_7742);
nand U7886 (N_7886,N_7728,N_7794);
and U7887 (N_7887,N_7638,N_7711);
and U7888 (N_7888,N_7635,N_7790);
xor U7889 (N_7889,N_7653,N_7620);
or U7890 (N_7890,N_7793,N_7791);
nand U7891 (N_7891,N_7736,N_7682);
and U7892 (N_7892,N_7763,N_7641);
and U7893 (N_7893,N_7655,N_7649);
nor U7894 (N_7894,N_7752,N_7726);
and U7895 (N_7895,N_7778,N_7761);
or U7896 (N_7896,N_7603,N_7756);
and U7897 (N_7897,N_7629,N_7718);
or U7898 (N_7898,N_7651,N_7650);
xnor U7899 (N_7899,N_7746,N_7626);
and U7900 (N_7900,N_7635,N_7723);
nor U7901 (N_7901,N_7740,N_7620);
nand U7902 (N_7902,N_7607,N_7761);
xnor U7903 (N_7903,N_7635,N_7670);
xor U7904 (N_7904,N_7676,N_7788);
nand U7905 (N_7905,N_7723,N_7780);
nand U7906 (N_7906,N_7745,N_7717);
or U7907 (N_7907,N_7679,N_7663);
nor U7908 (N_7908,N_7630,N_7688);
nor U7909 (N_7909,N_7633,N_7629);
nor U7910 (N_7910,N_7603,N_7608);
xnor U7911 (N_7911,N_7786,N_7619);
or U7912 (N_7912,N_7770,N_7653);
nand U7913 (N_7913,N_7602,N_7644);
or U7914 (N_7914,N_7674,N_7676);
nor U7915 (N_7915,N_7631,N_7657);
xnor U7916 (N_7916,N_7668,N_7748);
and U7917 (N_7917,N_7741,N_7766);
xnor U7918 (N_7918,N_7766,N_7639);
and U7919 (N_7919,N_7650,N_7624);
nand U7920 (N_7920,N_7703,N_7784);
and U7921 (N_7921,N_7615,N_7659);
nand U7922 (N_7922,N_7781,N_7701);
and U7923 (N_7923,N_7727,N_7743);
nand U7924 (N_7924,N_7670,N_7763);
or U7925 (N_7925,N_7753,N_7715);
xor U7926 (N_7926,N_7727,N_7703);
nand U7927 (N_7927,N_7745,N_7657);
nand U7928 (N_7928,N_7774,N_7779);
or U7929 (N_7929,N_7638,N_7642);
nand U7930 (N_7930,N_7696,N_7781);
xor U7931 (N_7931,N_7769,N_7748);
nor U7932 (N_7932,N_7794,N_7707);
nor U7933 (N_7933,N_7788,N_7617);
xnor U7934 (N_7934,N_7637,N_7608);
nor U7935 (N_7935,N_7610,N_7714);
nand U7936 (N_7936,N_7622,N_7719);
nor U7937 (N_7937,N_7687,N_7714);
nand U7938 (N_7938,N_7679,N_7601);
and U7939 (N_7939,N_7718,N_7685);
xor U7940 (N_7940,N_7747,N_7799);
xor U7941 (N_7941,N_7771,N_7772);
nand U7942 (N_7942,N_7623,N_7757);
xor U7943 (N_7943,N_7704,N_7690);
xnor U7944 (N_7944,N_7776,N_7713);
and U7945 (N_7945,N_7762,N_7607);
nand U7946 (N_7946,N_7665,N_7638);
xor U7947 (N_7947,N_7675,N_7661);
nand U7948 (N_7948,N_7632,N_7735);
nor U7949 (N_7949,N_7691,N_7668);
xor U7950 (N_7950,N_7676,N_7784);
and U7951 (N_7951,N_7792,N_7762);
or U7952 (N_7952,N_7692,N_7766);
xor U7953 (N_7953,N_7674,N_7654);
or U7954 (N_7954,N_7792,N_7734);
nand U7955 (N_7955,N_7744,N_7627);
nor U7956 (N_7956,N_7657,N_7676);
or U7957 (N_7957,N_7668,N_7630);
xor U7958 (N_7958,N_7705,N_7718);
xor U7959 (N_7959,N_7759,N_7670);
xor U7960 (N_7960,N_7739,N_7635);
xor U7961 (N_7961,N_7667,N_7787);
and U7962 (N_7962,N_7641,N_7664);
xnor U7963 (N_7963,N_7734,N_7676);
and U7964 (N_7964,N_7725,N_7724);
nor U7965 (N_7965,N_7644,N_7622);
xnor U7966 (N_7966,N_7603,N_7772);
or U7967 (N_7967,N_7634,N_7644);
xnor U7968 (N_7968,N_7782,N_7603);
and U7969 (N_7969,N_7603,N_7683);
and U7970 (N_7970,N_7746,N_7662);
nor U7971 (N_7971,N_7731,N_7614);
nand U7972 (N_7972,N_7648,N_7742);
xnor U7973 (N_7973,N_7708,N_7682);
or U7974 (N_7974,N_7602,N_7746);
or U7975 (N_7975,N_7778,N_7694);
or U7976 (N_7976,N_7663,N_7718);
or U7977 (N_7977,N_7787,N_7652);
or U7978 (N_7978,N_7711,N_7669);
or U7979 (N_7979,N_7680,N_7640);
nand U7980 (N_7980,N_7744,N_7644);
or U7981 (N_7981,N_7675,N_7615);
nand U7982 (N_7982,N_7719,N_7630);
and U7983 (N_7983,N_7622,N_7733);
xor U7984 (N_7984,N_7688,N_7634);
and U7985 (N_7985,N_7678,N_7776);
or U7986 (N_7986,N_7629,N_7772);
or U7987 (N_7987,N_7706,N_7746);
xor U7988 (N_7988,N_7635,N_7689);
nor U7989 (N_7989,N_7665,N_7766);
or U7990 (N_7990,N_7765,N_7752);
nor U7991 (N_7991,N_7748,N_7742);
or U7992 (N_7992,N_7610,N_7665);
nand U7993 (N_7993,N_7785,N_7624);
xnor U7994 (N_7994,N_7634,N_7691);
nor U7995 (N_7995,N_7787,N_7762);
and U7996 (N_7996,N_7776,N_7685);
nor U7997 (N_7997,N_7711,N_7635);
or U7998 (N_7998,N_7689,N_7671);
xnor U7999 (N_7999,N_7765,N_7777);
nor U8000 (N_8000,N_7884,N_7951);
xnor U8001 (N_8001,N_7972,N_7971);
and U8002 (N_8002,N_7869,N_7851);
or U8003 (N_8003,N_7896,N_7802);
nor U8004 (N_8004,N_7942,N_7854);
or U8005 (N_8005,N_7840,N_7841);
nand U8006 (N_8006,N_7823,N_7830);
xnor U8007 (N_8007,N_7899,N_7989);
or U8008 (N_8008,N_7836,N_7986);
and U8009 (N_8009,N_7955,N_7937);
nor U8010 (N_8010,N_7890,N_7992);
nor U8011 (N_8011,N_7976,N_7885);
xor U8012 (N_8012,N_7868,N_7956);
or U8013 (N_8013,N_7891,N_7936);
nor U8014 (N_8014,N_7873,N_7912);
or U8015 (N_8015,N_7879,N_7934);
and U8016 (N_8016,N_7888,N_7943);
or U8017 (N_8017,N_7847,N_7866);
nor U8018 (N_8018,N_7893,N_7945);
nand U8019 (N_8019,N_7923,N_7975);
or U8020 (N_8020,N_7979,N_7982);
nor U8021 (N_8021,N_7878,N_7970);
and U8022 (N_8022,N_7861,N_7995);
or U8023 (N_8023,N_7931,N_7906);
or U8024 (N_8024,N_7875,N_7839);
nand U8025 (N_8025,N_7918,N_7870);
and U8026 (N_8026,N_7900,N_7926);
and U8027 (N_8027,N_7944,N_7867);
xor U8028 (N_8028,N_7813,N_7927);
and U8029 (N_8029,N_7973,N_7855);
and U8030 (N_8030,N_7957,N_7984);
and U8031 (N_8031,N_7871,N_7985);
nor U8032 (N_8032,N_7815,N_7922);
xor U8033 (N_8033,N_7826,N_7905);
nand U8034 (N_8034,N_7910,N_7880);
xor U8035 (N_8035,N_7860,N_7849);
nor U8036 (N_8036,N_7953,N_7962);
nor U8037 (N_8037,N_7814,N_7844);
or U8038 (N_8038,N_7949,N_7886);
and U8039 (N_8039,N_7938,N_7846);
or U8040 (N_8040,N_7822,N_7831);
nor U8041 (N_8041,N_7859,N_7974);
nand U8042 (N_8042,N_7825,N_7950);
or U8043 (N_8043,N_7835,N_7996);
xnor U8044 (N_8044,N_7816,N_7845);
nand U8045 (N_8045,N_7933,N_7865);
or U8046 (N_8046,N_7930,N_7817);
and U8047 (N_8047,N_7842,N_7964);
and U8048 (N_8048,N_7812,N_7853);
and U8049 (N_8049,N_7925,N_7991);
nand U8050 (N_8050,N_7808,N_7901);
xnor U8051 (N_8051,N_7852,N_7883);
or U8052 (N_8052,N_7876,N_7941);
xnor U8053 (N_8053,N_7821,N_7894);
nor U8054 (N_8054,N_7916,N_7837);
xor U8055 (N_8055,N_7902,N_7935);
nor U8056 (N_8056,N_7856,N_7833);
xnor U8057 (N_8057,N_7824,N_7832);
nand U8058 (N_8058,N_7993,N_7960);
or U8059 (N_8059,N_7978,N_7954);
and U8060 (N_8060,N_7872,N_7850);
and U8061 (N_8061,N_7908,N_7952);
xnor U8062 (N_8062,N_7999,N_7903);
nor U8063 (N_8063,N_7803,N_7966);
and U8064 (N_8064,N_7843,N_7801);
nor U8065 (N_8065,N_7997,N_7827);
and U8066 (N_8066,N_7983,N_7914);
nand U8067 (N_8067,N_7858,N_7963);
nand U8068 (N_8068,N_7887,N_7913);
nand U8069 (N_8069,N_7967,N_7877);
and U8070 (N_8070,N_7959,N_7881);
nand U8071 (N_8071,N_7898,N_7911);
and U8072 (N_8072,N_7921,N_7969);
xor U8073 (N_8073,N_7920,N_7882);
or U8074 (N_8074,N_7965,N_7804);
nand U8075 (N_8075,N_7980,N_7990);
or U8076 (N_8076,N_7915,N_7904);
nand U8077 (N_8077,N_7820,N_7828);
or U8078 (N_8078,N_7874,N_7819);
nor U8079 (N_8079,N_7863,N_7864);
xor U8080 (N_8080,N_7857,N_7988);
nor U8081 (N_8081,N_7862,N_7946);
xnor U8082 (N_8082,N_7968,N_7987);
nor U8083 (N_8083,N_7948,N_7929);
nor U8084 (N_8084,N_7917,N_7834);
xnor U8085 (N_8085,N_7895,N_7811);
nor U8086 (N_8086,N_7940,N_7994);
and U8087 (N_8087,N_7800,N_7807);
xnor U8088 (N_8088,N_7907,N_7818);
nand U8089 (N_8089,N_7829,N_7998);
and U8090 (N_8090,N_7897,N_7924);
nand U8091 (N_8091,N_7958,N_7928);
xor U8092 (N_8092,N_7947,N_7805);
nand U8093 (N_8093,N_7838,N_7892);
and U8094 (N_8094,N_7919,N_7809);
nand U8095 (N_8095,N_7909,N_7810);
or U8096 (N_8096,N_7981,N_7889);
or U8097 (N_8097,N_7806,N_7977);
nand U8098 (N_8098,N_7848,N_7961);
xor U8099 (N_8099,N_7932,N_7939);
nor U8100 (N_8100,N_7999,N_7973);
xor U8101 (N_8101,N_7851,N_7982);
or U8102 (N_8102,N_7902,N_7817);
nor U8103 (N_8103,N_7888,N_7893);
xnor U8104 (N_8104,N_7973,N_7899);
xnor U8105 (N_8105,N_7837,N_7924);
nand U8106 (N_8106,N_7842,N_7882);
nor U8107 (N_8107,N_7839,N_7859);
or U8108 (N_8108,N_7899,N_7908);
or U8109 (N_8109,N_7940,N_7933);
xnor U8110 (N_8110,N_7944,N_7989);
and U8111 (N_8111,N_7874,N_7857);
and U8112 (N_8112,N_7932,N_7849);
and U8113 (N_8113,N_7975,N_7908);
nor U8114 (N_8114,N_7907,N_7848);
or U8115 (N_8115,N_7939,N_7836);
or U8116 (N_8116,N_7866,N_7988);
and U8117 (N_8117,N_7869,N_7912);
or U8118 (N_8118,N_7961,N_7837);
or U8119 (N_8119,N_7847,N_7991);
nor U8120 (N_8120,N_7876,N_7989);
or U8121 (N_8121,N_7878,N_7967);
nor U8122 (N_8122,N_7811,N_7875);
nor U8123 (N_8123,N_7942,N_7903);
nor U8124 (N_8124,N_7883,N_7912);
nor U8125 (N_8125,N_7823,N_7859);
nor U8126 (N_8126,N_7845,N_7944);
or U8127 (N_8127,N_7862,N_7837);
nand U8128 (N_8128,N_7977,N_7993);
or U8129 (N_8129,N_7982,N_7966);
xor U8130 (N_8130,N_7867,N_7993);
xor U8131 (N_8131,N_7912,N_7831);
nand U8132 (N_8132,N_7943,N_7921);
nor U8133 (N_8133,N_7952,N_7984);
or U8134 (N_8134,N_7937,N_7830);
or U8135 (N_8135,N_7884,N_7876);
xnor U8136 (N_8136,N_7847,N_7808);
nor U8137 (N_8137,N_7813,N_7953);
nor U8138 (N_8138,N_7923,N_7960);
and U8139 (N_8139,N_7824,N_7890);
xnor U8140 (N_8140,N_7896,N_7991);
xnor U8141 (N_8141,N_7865,N_7885);
nor U8142 (N_8142,N_7910,N_7914);
nor U8143 (N_8143,N_7954,N_7811);
nor U8144 (N_8144,N_7949,N_7802);
or U8145 (N_8145,N_7968,N_7990);
and U8146 (N_8146,N_7942,N_7839);
or U8147 (N_8147,N_7941,N_7949);
or U8148 (N_8148,N_7879,N_7918);
or U8149 (N_8149,N_7970,N_7997);
nor U8150 (N_8150,N_7884,N_7817);
nand U8151 (N_8151,N_7960,N_7801);
or U8152 (N_8152,N_7996,N_7886);
or U8153 (N_8153,N_7980,N_7845);
or U8154 (N_8154,N_7853,N_7943);
xor U8155 (N_8155,N_7855,N_7852);
xor U8156 (N_8156,N_7867,N_7836);
and U8157 (N_8157,N_7960,N_7917);
or U8158 (N_8158,N_7896,N_7883);
xor U8159 (N_8159,N_7800,N_7923);
nand U8160 (N_8160,N_7952,N_7890);
xor U8161 (N_8161,N_7885,N_7950);
or U8162 (N_8162,N_7967,N_7826);
xnor U8163 (N_8163,N_7920,N_7814);
xor U8164 (N_8164,N_7937,N_7812);
nand U8165 (N_8165,N_7903,N_7994);
nor U8166 (N_8166,N_7974,N_7965);
nor U8167 (N_8167,N_7884,N_7992);
xnor U8168 (N_8168,N_7827,N_7925);
nand U8169 (N_8169,N_7945,N_7905);
or U8170 (N_8170,N_7917,N_7972);
or U8171 (N_8171,N_7903,N_7886);
and U8172 (N_8172,N_7997,N_7990);
or U8173 (N_8173,N_7805,N_7830);
nand U8174 (N_8174,N_7955,N_7830);
and U8175 (N_8175,N_7966,N_7955);
xnor U8176 (N_8176,N_7870,N_7805);
or U8177 (N_8177,N_7825,N_7885);
nor U8178 (N_8178,N_7912,N_7826);
nand U8179 (N_8179,N_7945,N_7884);
and U8180 (N_8180,N_7833,N_7923);
or U8181 (N_8181,N_7843,N_7888);
and U8182 (N_8182,N_7817,N_7849);
nand U8183 (N_8183,N_7840,N_7973);
or U8184 (N_8184,N_7814,N_7904);
or U8185 (N_8185,N_7867,N_7879);
nand U8186 (N_8186,N_7805,N_7954);
nand U8187 (N_8187,N_7945,N_7930);
or U8188 (N_8188,N_7952,N_7810);
nand U8189 (N_8189,N_7816,N_7808);
and U8190 (N_8190,N_7933,N_7849);
nand U8191 (N_8191,N_7846,N_7836);
and U8192 (N_8192,N_7956,N_7923);
or U8193 (N_8193,N_7861,N_7883);
xor U8194 (N_8194,N_7839,N_7877);
or U8195 (N_8195,N_7830,N_7843);
nor U8196 (N_8196,N_7838,N_7908);
or U8197 (N_8197,N_7907,N_7800);
nor U8198 (N_8198,N_7868,N_7912);
xor U8199 (N_8199,N_7933,N_7936);
or U8200 (N_8200,N_8071,N_8027);
xor U8201 (N_8201,N_8135,N_8128);
nand U8202 (N_8202,N_8030,N_8160);
and U8203 (N_8203,N_8155,N_8197);
xor U8204 (N_8204,N_8118,N_8061);
nand U8205 (N_8205,N_8068,N_8091);
nand U8206 (N_8206,N_8152,N_8072);
nand U8207 (N_8207,N_8020,N_8003);
or U8208 (N_8208,N_8015,N_8194);
and U8209 (N_8209,N_8076,N_8146);
or U8210 (N_8210,N_8059,N_8166);
or U8211 (N_8211,N_8131,N_8074);
xnor U8212 (N_8212,N_8114,N_8064);
nand U8213 (N_8213,N_8134,N_8028);
nand U8214 (N_8214,N_8161,N_8172);
nand U8215 (N_8215,N_8127,N_8024);
or U8216 (N_8216,N_8005,N_8139);
nand U8217 (N_8217,N_8056,N_8110);
or U8218 (N_8218,N_8007,N_8174);
xor U8219 (N_8219,N_8132,N_8122);
xnor U8220 (N_8220,N_8034,N_8108);
nand U8221 (N_8221,N_8001,N_8021);
and U8222 (N_8222,N_8189,N_8018);
or U8223 (N_8223,N_8058,N_8148);
nand U8224 (N_8224,N_8191,N_8125);
xnor U8225 (N_8225,N_8037,N_8186);
nand U8226 (N_8226,N_8060,N_8038);
and U8227 (N_8227,N_8078,N_8013);
xnor U8228 (N_8228,N_8102,N_8178);
xor U8229 (N_8229,N_8079,N_8065);
nand U8230 (N_8230,N_8039,N_8107);
xor U8231 (N_8231,N_8156,N_8004);
or U8232 (N_8232,N_8133,N_8130);
nand U8233 (N_8233,N_8142,N_8137);
and U8234 (N_8234,N_8096,N_8090);
or U8235 (N_8235,N_8116,N_8159);
xnor U8236 (N_8236,N_8040,N_8164);
nand U8237 (N_8237,N_8082,N_8149);
nor U8238 (N_8238,N_8106,N_8175);
xor U8239 (N_8239,N_8045,N_8181);
xnor U8240 (N_8240,N_8052,N_8077);
nand U8241 (N_8241,N_8073,N_8049);
or U8242 (N_8242,N_8173,N_8011);
nor U8243 (N_8243,N_8150,N_8033);
nor U8244 (N_8244,N_8136,N_8051);
and U8245 (N_8245,N_8067,N_8089);
nand U8246 (N_8246,N_8123,N_8098);
and U8247 (N_8247,N_8083,N_8048);
and U8248 (N_8248,N_8062,N_8145);
xnor U8249 (N_8249,N_8093,N_8121);
xor U8250 (N_8250,N_8109,N_8047);
xnor U8251 (N_8251,N_8036,N_8054);
nand U8252 (N_8252,N_8113,N_8000);
nor U8253 (N_8253,N_8171,N_8032);
nand U8254 (N_8254,N_8162,N_8100);
and U8255 (N_8255,N_8023,N_8140);
or U8256 (N_8256,N_8002,N_8179);
and U8257 (N_8257,N_8088,N_8193);
nor U8258 (N_8258,N_8012,N_8042);
nand U8259 (N_8259,N_8168,N_8025);
and U8260 (N_8260,N_8184,N_8099);
or U8261 (N_8261,N_8043,N_8111);
nor U8262 (N_8262,N_8177,N_8183);
nor U8263 (N_8263,N_8094,N_8080);
nand U8264 (N_8264,N_8017,N_8095);
xor U8265 (N_8265,N_8097,N_8087);
nor U8266 (N_8266,N_8063,N_8180);
and U8267 (N_8267,N_8112,N_8019);
xor U8268 (N_8268,N_8192,N_8016);
or U8269 (N_8269,N_8010,N_8143);
and U8270 (N_8270,N_8199,N_8029);
and U8271 (N_8271,N_8014,N_8129);
nand U8272 (N_8272,N_8101,N_8153);
and U8273 (N_8273,N_8041,N_8141);
or U8274 (N_8274,N_8176,N_8066);
nor U8275 (N_8275,N_8120,N_8103);
nand U8276 (N_8276,N_8055,N_8053);
nand U8277 (N_8277,N_8124,N_8198);
nor U8278 (N_8278,N_8169,N_8138);
xor U8279 (N_8279,N_8069,N_8157);
xnor U8280 (N_8280,N_8147,N_8163);
nor U8281 (N_8281,N_8085,N_8196);
nor U8282 (N_8282,N_8081,N_8044);
and U8283 (N_8283,N_8170,N_8046);
nor U8284 (N_8284,N_8031,N_8195);
xnor U8285 (N_8285,N_8117,N_8187);
and U8286 (N_8286,N_8165,N_8185);
or U8287 (N_8287,N_8154,N_8144);
nor U8288 (N_8288,N_8190,N_8158);
xor U8289 (N_8289,N_8115,N_8084);
nand U8290 (N_8290,N_8151,N_8070);
or U8291 (N_8291,N_8119,N_8188);
nor U8292 (N_8292,N_8008,N_8006);
nand U8293 (N_8293,N_8182,N_8026);
or U8294 (N_8294,N_8057,N_8022);
and U8295 (N_8295,N_8104,N_8050);
nor U8296 (N_8296,N_8092,N_8105);
or U8297 (N_8297,N_8075,N_8086);
xnor U8298 (N_8298,N_8167,N_8126);
nand U8299 (N_8299,N_8035,N_8009);
or U8300 (N_8300,N_8029,N_8190);
nor U8301 (N_8301,N_8079,N_8086);
or U8302 (N_8302,N_8067,N_8038);
and U8303 (N_8303,N_8154,N_8145);
nor U8304 (N_8304,N_8149,N_8107);
xnor U8305 (N_8305,N_8148,N_8009);
or U8306 (N_8306,N_8100,N_8026);
and U8307 (N_8307,N_8027,N_8053);
nor U8308 (N_8308,N_8099,N_8114);
and U8309 (N_8309,N_8121,N_8116);
nand U8310 (N_8310,N_8143,N_8157);
nand U8311 (N_8311,N_8028,N_8046);
nand U8312 (N_8312,N_8001,N_8047);
xnor U8313 (N_8313,N_8001,N_8107);
xnor U8314 (N_8314,N_8003,N_8012);
xnor U8315 (N_8315,N_8010,N_8055);
or U8316 (N_8316,N_8198,N_8180);
and U8317 (N_8317,N_8113,N_8138);
nand U8318 (N_8318,N_8173,N_8007);
and U8319 (N_8319,N_8147,N_8088);
xor U8320 (N_8320,N_8155,N_8087);
or U8321 (N_8321,N_8078,N_8025);
nor U8322 (N_8322,N_8107,N_8115);
nand U8323 (N_8323,N_8100,N_8016);
nor U8324 (N_8324,N_8069,N_8194);
xor U8325 (N_8325,N_8150,N_8128);
and U8326 (N_8326,N_8183,N_8051);
xnor U8327 (N_8327,N_8025,N_8059);
nor U8328 (N_8328,N_8177,N_8021);
nor U8329 (N_8329,N_8095,N_8166);
nor U8330 (N_8330,N_8126,N_8053);
nand U8331 (N_8331,N_8014,N_8010);
nand U8332 (N_8332,N_8097,N_8002);
nand U8333 (N_8333,N_8186,N_8076);
xnor U8334 (N_8334,N_8170,N_8172);
nor U8335 (N_8335,N_8126,N_8150);
and U8336 (N_8336,N_8184,N_8078);
nor U8337 (N_8337,N_8050,N_8039);
nand U8338 (N_8338,N_8043,N_8032);
or U8339 (N_8339,N_8027,N_8186);
xor U8340 (N_8340,N_8011,N_8019);
and U8341 (N_8341,N_8112,N_8196);
and U8342 (N_8342,N_8131,N_8123);
and U8343 (N_8343,N_8183,N_8128);
or U8344 (N_8344,N_8128,N_8184);
nor U8345 (N_8345,N_8016,N_8133);
and U8346 (N_8346,N_8156,N_8031);
or U8347 (N_8347,N_8150,N_8142);
xnor U8348 (N_8348,N_8094,N_8194);
nor U8349 (N_8349,N_8051,N_8154);
or U8350 (N_8350,N_8180,N_8006);
nand U8351 (N_8351,N_8140,N_8061);
nand U8352 (N_8352,N_8005,N_8101);
or U8353 (N_8353,N_8182,N_8159);
xnor U8354 (N_8354,N_8155,N_8154);
nor U8355 (N_8355,N_8095,N_8045);
and U8356 (N_8356,N_8099,N_8157);
nand U8357 (N_8357,N_8131,N_8046);
nand U8358 (N_8358,N_8115,N_8129);
xor U8359 (N_8359,N_8029,N_8013);
and U8360 (N_8360,N_8172,N_8060);
and U8361 (N_8361,N_8146,N_8073);
nor U8362 (N_8362,N_8068,N_8181);
nand U8363 (N_8363,N_8016,N_8078);
and U8364 (N_8364,N_8089,N_8126);
nor U8365 (N_8365,N_8110,N_8103);
nor U8366 (N_8366,N_8197,N_8152);
nor U8367 (N_8367,N_8151,N_8069);
and U8368 (N_8368,N_8112,N_8078);
xnor U8369 (N_8369,N_8175,N_8163);
and U8370 (N_8370,N_8183,N_8113);
and U8371 (N_8371,N_8078,N_8169);
nand U8372 (N_8372,N_8105,N_8099);
and U8373 (N_8373,N_8166,N_8140);
nand U8374 (N_8374,N_8048,N_8152);
nor U8375 (N_8375,N_8050,N_8052);
xnor U8376 (N_8376,N_8087,N_8060);
or U8377 (N_8377,N_8050,N_8187);
and U8378 (N_8378,N_8187,N_8053);
xnor U8379 (N_8379,N_8168,N_8036);
xor U8380 (N_8380,N_8001,N_8108);
xor U8381 (N_8381,N_8115,N_8092);
xnor U8382 (N_8382,N_8077,N_8072);
xnor U8383 (N_8383,N_8020,N_8022);
nand U8384 (N_8384,N_8105,N_8125);
or U8385 (N_8385,N_8049,N_8082);
nand U8386 (N_8386,N_8039,N_8146);
or U8387 (N_8387,N_8131,N_8169);
nor U8388 (N_8388,N_8188,N_8123);
nor U8389 (N_8389,N_8075,N_8089);
xor U8390 (N_8390,N_8062,N_8075);
xor U8391 (N_8391,N_8176,N_8101);
and U8392 (N_8392,N_8180,N_8024);
nor U8393 (N_8393,N_8164,N_8081);
or U8394 (N_8394,N_8092,N_8155);
or U8395 (N_8395,N_8052,N_8064);
and U8396 (N_8396,N_8159,N_8042);
and U8397 (N_8397,N_8142,N_8197);
or U8398 (N_8398,N_8058,N_8120);
and U8399 (N_8399,N_8083,N_8082);
xor U8400 (N_8400,N_8293,N_8331);
or U8401 (N_8401,N_8211,N_8213);
nand U8402 (N_8402,N_8220,N_8301);
or U8403 (N_8403,N_8330,N_8381);
nor U8404 (N_8404,N_8378,N_8355);
nor U8405 (N_8405,N_8310,N_8204);
and U8406 (N_8406,N_8373,N_8291);
xor U8407 (N_8407,N_8200,N_8268);
xnor U8408 (N_8408,N_8228,N_8274);
nand U8409 (N_8409,N_8322,N_8239);
xnor U8410 (N_8410,N_8234,N_8302);
or U8411 (N_8411,N_8385,N_8344);
and U8412 (N_8412,N_8246,N_8384);
and U8413 (N_8413,N_8313,N_8372);
nand U8414 (N_8414,N_8386,N_8252);
or U8415 (N_8415,N_8303,N_8299);
or U8416 (N_8416,N_8208,N_8203);
nor U8417 (N_8417,N_8223,N_8216);
xnor U8418 (N_8418,N_8327,N_8392);
or U8419 (N_8419,N_8332,N_8281);
nand U8420 (N_8420,N_8267,N_8219);
xnor U8421 (N_8421,N_8230,N_8316);
and U8422 (N_8422,N_8292,N_8306);
or U8423 (N_8423,N_8287,N_8340);
nor U8424 (N_8424,N_8202,N_8269);
xnor U8425 (N_8425,N_8398,N_8396);
nand U8426 (N_8426,N_8352,N_8311);
xor U8427 (N_8427,N_8377,N_8270);
xnor U8428 (N_8428,N_8248,N_8249);
xor U8429 (N_8429,N_8260,N_8298);
nand U8430 (N_8430,N_8368,N_8359);
nand U8431 (N_8431,N_8304,N_8285);
xnor U8432 (N_8432,N_8279,N_8337);
or U8433 (N_8433,N_8276,N_8362);
nor U8434 (N_8434,N_8387,N_8232);
xor U8435 (N_8435,N_8300,N_8379);
or U8436 (N_8436,N_8369,N_8382);
or U8437 (N_8437,N_8336,N_8214);
or U8438 (N_8438,N_8262,N_8238);
nor U8439 (N_8439,N_8370,N_8236);
nor U8440 (N_8440,N_8254,N_8317);
nand U8441 (N_8441,N_8391,N_8342);
and U8442 (N_8442,N_8264,N_8375);
xnor U8443 (N_8443,N_8272,N_8278);
nand U8444 (N_8444,N_8222,N_8329);
nor U8445 (N_8445,N_8324,N_8288);
or U8446 (N_8446,N_8393,N_8212);
nor U8447 (N_8447,N_8271,N_8314);
nand U8448 (N_8448,N_8245,N_8354);
nand U8449 (N_8449,N_8371,N_8207);
nand U8450 (N_8450,N_8265,N_8226);
xnor U8451 (N_8451,N_8389,N_8289);
xnor U8452 (N_8452,N_8383,N_8345);
xor U8453 (N_8453,N_8256,N_8357);
and U8454 (N_8454,N_8374,N_8255);
or U8455 (N_8455,N_8218,N_8356);
xor U8456 (N_8456,N_8326,N_8315);
xnor U8457 (N_8457,N_8358,N_8243);
nand U8458 (N_8458,N_8363,N_8305);
and U8459 (N_8459,N_8376,N_8233);
nor U8460 (N_8460,N_8210,N_8201);
nand U8461 (N_8461,N_8253,N_8250);
and U8462 (N_8462,N_8309,N_8297);
xnor U8463 (N_8463,N_8312,N_8390);
xor U8464 (N_8464,N_8294,N_8242);
or U8465 (N_8465,N_8296,N_8380);
nor U8466 (N_8466,N_8290,N_8320);
nand U8467 (N_8467,N_8240,N_8353);
and U8468 (N_8468,N_8215,N_8348);
or U8469 (N_8469,N_8244,N_8231);
nand U8470 (N_8470,N_8225,N_8338);
xor U8471 (N_8471,N_8227,N_8283);
or U8472 (N_8472,N_8328,N_8280);
nand U8473 (N_8473,N_8399,N_8394);
and U8474 (N_8474,N_8361,N_8360);
nor U8475 (N_8475,N_8282,N_8339);
nor U8476 (N_8476,N_8321,N_8263);
and U8477 (N_8477,N_8341,N_8366);
nand U8478 (N_8478,N_8333,N_8273);
or U8479 (N_8479,N_8325,N_8257);
or U8480 (N_8480,N_8334,N_8284);
nand U8481 (N_8481,N_8258,N_8277);
nor U8482 (N_8482,N_8318,N_8388);
nor U8483 (N_8483,N_8209,N_8266);
nand U8484 (N_8484,N_8235,N_8206);
xor U8485 (N_8485,N_8346,N_8349);
xor U8486 (N_8486,N_8335,N_8229);
and U8487 (N_8487,N_8365,N_8350);
and U8488 (N_8488,N_8295,N_8395);
nand U8489 (N_8489,N_8364,N_8367);
nand U8490 (N_8490,N_8247,N_8217);
nor U8491 (N_8491,N_8319,N_8307);
xor U8492 (N_8492,N_8205,N_8351);
and U8493 (N_8493,N_8251,N_8308);
xor U8494 (N_8494,N_8261,N_8323);
nor U8495 (N_8495,N_8221,N_8275);
nor U8496 (N_8496,N_8347,N_8241);
xor U8497 (N_8497,N_8237,N_8343);
and U8498 (N_8498,N_8259,N_8224);
or U8499 (N_8499,N_8286,N_8397);
nand U8500 (N_8500,N_8290,N_8273);
nand U8501 (N_8501,N_8300,N_8263);
and U8502 (N_8502,N_8279,N_8217);
nor U8503 (N_8503,N_8345,N_8244);
nand U8504 (N_8504,N_8339,N_8359);
or U8505 (N_8505,N_8232,N_8309);
and U8506 (N_8506,N_8344,N_8218);
or U8507 (N_8507,N_8368,N_8243);
xnor U8508 (N_8508,N_8273,N_8262);
and U8509 (N_8509,N_8208,N_8320);
xnor U8510 (N_8510,N_8323,N_8303);
nand U8511 (N_8511,N_8325,N_8256);
xnor U8512 (N_8512,N_8269,N_8354);
and U8513 (N_8513,N_8394,N_8252);
xnor U8514 (N_8514,N_8250,N_8364);
nor U8515 (N_8515,N_8359,N_8246);
and U8516 (N_8516,N_8294,N_8396);
nor U8517 (N_8517,N_8240,N_8259);
xor U8518 (N_8518,N_8337,N_8284);
nor U8519 (N_8519,N_8394,N_8259);
nor U8520 (N_8520,N_8373,N_8349);
and U8521 (N_8521,N_8398,N_8251);
nand U8522 (N_8522,N_8384,N_8269);
nor U8523 (N_8523,N_8373,N_8229);
xnor U8524 (N_8524,N_8245,N_8237);
nor U8525 (N_8525,N_8345,N_8382);
nor U8526 (N_8526,N_8341,N_8279);
xor U8527 (N_8527,N_8378,N_8312);
nand U8528 (N_8528,N_8220,N_8224);
and U8529 (N_8529,N_8261,N_8284);
xnor U8530 (N_8530,N_8324,N_8202);
and U8531 (N_8531,N_8299,N_8380);
xnor U8532 (N_8532,N_8216,N_8292);
and U8533 (N_8533,N_8294,N_8270);
xnor U8534 (N_8534,N_8381,N_8213);
xnor U8535 (N_8535,N_8220,N_8371);
nand U8536 (N_8536,N_8294,N_8247);
nand U8537 (N_8537,N_8239,N_8392);
and U8538 (N_8538,N_8321,N_8392);
and U8539 (N_8539,N_8219,N_8361);
xor U8540 (N_8540,N_8243,N_8202);
and U8541 (N_8541,N_8228,N_8390);
xnor U8542 (N_8542,N_8303,N_8384);
nand U8543 (N_8543,N_8389,N_8399);
nand U8544 (N_8544,N_8327,N_8222);
xor U8545 (N_8545,N_8300,N_8235);
nor U8546 (N_8546,N_8321,N_8378);
and U8547 (N_8547,N_8279,N_8330);
or U8548 (N_8548,N_8265,N_8238);
xnor U8549 (N_8549,N_8301,N_8369);
or U8550 (N_8550,N_8302,N_8379);
nand U8551 (N_8551,N_8270,N_8213);
or U8552 (N_8552,N_8349,N_8293);
or U8553 (N_8553,N_8317,N_8203);
xnor U8554 (N_8554,N_8300,N_8290);
and U8555 (N_8555,N_8200,N_8292);
or U8556 (N_8556,N_8391,N_8373);
nor U8557 (N_8557,N_8260,N_8208);
and U8558 (N_8558,N_8249,N_8298);
or U8559 (N_8559,N_8279,N_8321);
nor U8560 (N_8560,N_8334,N_8352);
or U8561 (N_8561,N_8248,N_8350);
or U8562 (N_8562,N_8293,N_8364);
nand U8563 (N_8563,N_8323,N_8255);
nor U8564 (N_8564,N_8393,N_8278);
or U8565 (N_8565,N_8362,N_8373);
xnor U8566 (N_8566,N_8369,N_8293);
xnor U8567 (N_8567,N_8209,N_8294);
nand U8568 (N_8568,N_8329,N_8279);
or U8569 (N_8569,N_8312,N_8323);
or U8570 (N_8570,N_8271,N_8295);
nand U8571 (N_8571,N_8200,N_8250);
and U8572 (N_8572,N_8262,N_8361);
xor U8573 (N_8573,N_8253,N_8278);
nand U8574 (N_8574,N_8359,N_8280);
nor U8575 (N_8575,N_8300,N_8351);
and U8576 (N_8576,N_8377,N_8391);
nand U8577 (N_8577,N_8383,N_8312);
or U8578 (N_8578,N_8295,N_8331);
nand U8579 (N_8579,N_8230,N_8312);
nand U8580 (N_8580,N_8285,N_8387);
xnor U8581 (N_8581,N_8269,N_8334);
and U8582 (N_8582,N_8284,N_8234);
and U8583 (N_8583,N_8276,N_8379);
xnor U8584 (N_8584,N_8202,N_8236);
xnor U8585 (N_8585,N_8375,N_8378);
nor U8586 (N_8586,N_8330,N_8385);
nor U8587 (N_8587,N_8231,N_8257);
nand U8588 (N_8588,N_8334,N_8398);
nand U8589 (N_8589,N_8204,N_8331);
nor U8590 (N_8590,N_8254,N_8270);
xnor U8591 (N_8591,N_8277,N_8296);
or U8592 (N_8592,N_8258,N_8260);
or U8593 (N_8593,N_8224,N_8300);
nand U8594 (N_8594,N_8376,N_8243);
nor U8595 (N_8595,N_8285,N_8300);
xnor U8596 (N_8596,N_8348,N_8217);
xor U8597 (N_8597,N_8224,N_8273);
xnor U8598 (N_8598,N_8351,N_8245);
and U8599 (N_8599,N_8263,N_8354);
and U8600 (N_8600,N_8453,N_8422);
nand U8601 (N_8601,N_8507,N_8468);
and U8602 (N_8602,N_8408,N_8493);
or U8603 (N_8603,N_8491,N_8536);
or U8604 (N_8604,N_8582,N_8470);
or U8605 (N_8605,N_8500,N_8532);
and U8606 (N_8606,N_8599,N_8591);
or U8607 (N_8607,N_8490,N_8561);
nand U8608 (N_8608,N_8511,N_8409);
xor U8609 (N_8609,N_8560,N_8423);
or U8610 (N_8610,N_8462,N_8598);
or U8611 (N_8611,N_8497,N_8530);
nand U8612 (N_8612,N_8501,N_8440);
nor U8613 (N_8613,N_8518,N_8526);
nand U8614 (N_8614,N_8412,N_8459);
nor U8615 (N_8615,N_8478,N_8419);
and U8616 (N_8616,N_8436,N_8428);
and U8617 (N_8617,N_8541,N_8448);
and U8618 (N_8618,N_8405,N_8458);
and U8619 (N_8619,N_8445,N_8472);
or U8620 (N_8620,N_8535,N_8502);
xor U8621 (N_8621,N_8517,N_8488);
nand U8622 (N_8622,N_8531,N_8442);
and U8623 (N_8623,N_8433,N_8452);
nor U8624 (N_8624,N_8588,N_8571);
nand U8625 (N_8625,N_8524,N_8569);
or U8626 (N_8626,N_8481,N_8596);
and U8627 (N_8627,N_8595,N_8558);
nor U8628 (N_8628,N_8523,N_8577);
nor U8629 (N_8629,N_8548,N_8441);
nor U8630 (N_8630,N_8461,N_8566);
or U8631 (N_8631,N_8544,N_8471);
nor U8632 (N_8632,N_8499,N_8403);
nand U8633 (N_8633,N_8549,N_8513);
xor U8634 (N_8634,N_8414,N_8555);
nand U8635 (N_8635,N_8584,N_8463);
xnor U8636 (N_8636,N_8533,N_8590);
xnor U8637 (N_8637,N_8456,N_8585);
or U8638 (N_8638,N_8537,N_8475);
or U8639 (N_8639,N_8427,N_8457);
nor U8640 (N_8640,N_8438,N_8514);
xnor U8641 (N_8641,N_8444,N_8416);
xor U8642 (N_8642,N_8477,N_8534);
and U8643 (N_8643,N_8552,N_8492);
or U8644 (N_8644,N_8402,N_8597);
xor U8645 (N_8645,N_8510,N_8543);
or U8646 (N_8646,N_8411,N_8574);
xnor U8647 (N_8647,N_8527,N_8447);
or U8648 (N_8648,N_8480,N_8464);
and U8649 (N_8649,N_8476,N_8521);
or U8650 (N_8650,N_8451,N_8525);
nand U8651 (N_8651,N_8406,N_8512);
nor U8652 (N_8652,N_8469,N_8455);
and U8653 (N_8653,N_8564,N_8439);
and U8654 (N_8654,N_8426,N_8494);
and U8655 (N_8655,N_8431,N_8509);
xnor U8656 (N_8656,N_8505,N_8429);
or U8657 (N_8657,N_8483,N_8553);
xnor U8658 (N_8658,N_8587,N_8454);
or U8659 (N_8659,N_8520,N_8487);
and U8660 (N_8660,N_8508,N_8506);
nor U8661 (N_8661,N_8413,N_8586);
xor U8662 (N_8662,N_8410,N_8593);
and U8663 (N_8663,N_8559,N_8562);
and U8664 (N_8664,N_8579,N_8539);
xnor U8665 (N_8665,N_8594,N_8400);
xnor U8666 (N_8666,N_8592,N_8576);
or U8667 (N_8667,N_8465,N_8565);
nand U8668 (N_8668,N_8479,N_8573);
and U8669 (N_8669,N_8546,N_8437);
nand U8670 (N_8670,N_8482,N_8449);
nor U8671 (N_8671,N_8460,N_8554);
and U8672 (N_8672,N_8415,N_8418);
nand U8673 (N_8673,N_8417,N_8515);
and U8674 (N_8674,N_8516,N_8556);
and U8675 (N_8675,N_8580,N_8450);
and U8676 (N_8676,N_8489,N_8401);
or U8677 (N_8677,N_8496,N_8432);
nand U8678 (N_8678,N_8583,N_8542);
and U8679 (N_8679,N_8519,N_8570);
nand U8680 (N_8680,N_8443,N_8495);
and U8681 (N_8681,N_8424,N_8446);
or U8682 (N_8682,N_8434,N_8522);
and U8683 (N_8683,N_8503,N_8484);
nand U8684 (N_8684,N_8467,N_8421);
nand U8685 (N_8685,N_8575,N_8430);
or U8686 (N_8686,N_8529,N_8474);
or U8687 (N_8687,N_8498,N_8407);
and U8688 (N_8688,N_8578,N_8557);
and U8689 (N_8689,N_8545,N_8551);
nand U8690 (N_8690,N_8581,N_8572);
and U8691 (N_8691,N_8563,N_8550);
xor U8692 (N_8692,N_8528,N_8473);
or U8693 (N_8693,N_8404,N_8466);
or U8694 (N_8694,N_8425,N_8420);
nand U8695 (N_8695,N_8567,N_8568);
xor U8696 (N_8696,N_8435,N_8485);
and U8697 (N_8697,N_8538,N_8540);
nor U8698 (N_8698,N_8486,N_8589);
and U8699 (N_8699,N_8504,N_8547);
nand U8700 (N_8700,N_8525,N_8459);
and U8701 (N_8701,N_8471,N_8510);
or U8702 (N_8702,N_8403,N_8449);
or U8703 (N_8703,N_8518,N_8408);
nand U8704 (N_8704,N_8565,N_8413);
or U8705 (N_8705,N_8585,N_8433);
nand U8706 (N_8706,N_8535,N_8526);
xnor U8707 (N_8707,N_8423,N_8434);
xnor U8708 (N_8708,N_8419,N_8508);
nor U8709 (N_8709,N_8401,N_8576);
xnor U8710 (N_8710,N_8430,N_8505);
nand U8711 (N_8711,N_8592,N_8588);
xor U8712 (N_8712,N_8570,N_8581);
nand U8713 (N_8713,N_8411,N_8552);
or U8714 (N_8714,N_8568,N_8573);
nor U8715 (N_8715,N_8592,N_8496);
nand U8716 (N_8716,N_8532,N_8568);
nand U8717 (N_8717,N_8428,N_8539);
xor U8718 (N_8718,N_8587,N_8473);
and U8719 (N_8719,N_8528,N_8558);
xor U8720 (N_8720,N_8588,N_8502);
nand U8721 (N_8721,N_8538,N_8529);
xor U8722 (N_8722,N_8446,N_8400);
nor U8723 (N_8723,N_8431,N_8453);
and U8724 (N_8724,N_8579,N_8488);
xnor U8725 (N_8725,N_8452,N_8499);
nor U8726 (N_8726,N_8425,N_8457);
nand U8727 (N_8727,N_8452,N_8577);
and U8728 (N_8728,N_8409,N_8420);
xor U8729 (N_8729,N_8485,N_8449);
xor U8730 (N_8730,N_8453,N_8417);
or U8731 (N_8731,N_8541,N_8418);
or U8732 (N_8732,N_8438,N_8548);
and U8733 (N_8733,N_8435,N_8594);
xnor U8734 (N_8734,N_8415,N_8547);
xor U8735 (N_8735,N_8548,N_8525);
nand U8736 (N_8736,N_8571,N_8402);
nand U8737 (N_8737,N_8498,N_8528);
nor U8738 (N_8738,N_8484,N_8403);
or U8739 (N_8739,N_8434,N_8549);
and U8740 (N_8740,N_8464,N_8434);
nor U8741 (N_8741,N_8531,N_8575);
nand U8742 (N_8742,N_8498,N_8593);
and U8743 (N_8743,N_8423,N_8424);
or U8744 (N_8744,N_8476,N_8583);
or U8745 (N_8745,N_8559,N_8479);
nand U8746 (N_8746,N_8580,N_8556);
and U8747 (N_8747,N_8459,N_8469);
nor U8748 (N_8748,N_8507,N_8531);
or U8749 (N_8749,N_8456,N_8465);
xnor U8750 (N_8750,N_8489,N_8403);
and U8751 (N_8751,N_8504,N_8566);
nand U8752 (N_8752,N_8483,N_8578);
or U8753 (N_8753,N_8528,N_8469);
or U8754 (N_8754,N_8434,N_8593);
xor U8755 (N_8755,N_8575,N_8571);
and U8756 (N_8756,N_8464,N_8472);
xnor U8757 (N_8757,N_8583,N_8539);
nor U8758 (N_8758,N_8464,N_8437);
or U8759 (N_8759,N_8569,N_8514);
nand U8760 (N_8760,N_8574,N_8454);
or U8761 (N_8761,N_8504,N_8415);
nand U8762 (N_8762,N_8586,N_8446);
or U8763 (N_8763,N_8429,N_8512);
and U8764 (N_8764,N_8566,N_8455);
and U8765 (N_8765,N_8424,N_8405);
and U8766 (N_8766,N_8490,N_8454);
nand U8767 (N_8767,N_8583,N_8405);
or U8768 (N_8768,N_8598,N_8526);
or U8769 (N_8769,N_8475,N_8528);
nor U8770 (N_8770,N_8454,N_8504);
nand U8771 (N_8771,N_8535,N_8445);
and U8772 (N_8772,N_8540,N_8556);
nor U8773 (N_8773,N_8402,N_8526);
and U8774 (N_8774,N_8462,N_8578);
or U8775 (N_8775,N_8591,N_8432);
xor U8776 (N_8776,N_8553,N_8534);
nor U8777 (N_8777,N_8425,N_8408);
nor U8778 (N_8778,N_8559,N_8437);
and U8779 (N_8779,N_8461,N_8472);
nor U8780 (N_8780,N_8598,N_8471);
xor U8781 (N_8781,N_8591,N_8550);
nand U8782 (N_8782,N_8576,N_8491);
or U8783 (N_8783,N_8511,N_8567);
nor U8784 (N_8784,N_8591,N_8553);
nor U8785 (N_8785,N_8427,N_8446);
and U8786 (N_8786,N_8505,N_8484);
xor U8787 (N_8787,N_8501,N_8428);
and U8788 (N_8788,N_8546,N_8519);
or U8789 (N_8789,N_8426,N_8488);
nor U8790 (N_8790,N_8525,N_8496);
nand U8791 (N_8791,N_8568,N_8428);
xor U8792 (N_8792,N_8595,N_8482);
nor U8793 (N_8793,N_8596,N_8576);
and U8794 (N_8794,N_8493,N_8501);
nand U8795 (N_8795,N_8567,N_8456);
nand U8796 (N_8796,N_8503,N_8460);
and U8797 (N_8797,N_8445,N_8572);
and U8798 (N_8798,N_8460,N_8413);
or U8799 (N_8799,N_8578,N_8427);
nor U8800 (N_8800,N_8703,N_8699);
or U8801 (N_8801,N_8733,N_8629);
xor U8802 (N_8802,N_8683,N_8730);
nand U8803 (N_8803,N_8622,N_8685);
and U8804 (N_8804,N_8799,N_8790);
nand U8805 (N_8805,N_8741,N_8749);
xor U8806 (N_8806,N_8704,N_8692);
nor U8807 (N_8807,N_8716,N_8772);
nor U8808 (N_8808,N_8708,N_8756);
and U8809 (N_8809,N_8725,N_8639);
xor U8810 (N_8810,N_8735,N_8760);
nor U8811 (N_8811,N_8675,N_8686);
nor U8812 (N_8812,N_8724,N_8705);
xnor U8813 (N_8813,N_8743,N_8626);
nand U8814 (N_8814,N_8712,N_8660);
and U8815 (N_8815,N_8765,N_8696);
and U8816 (N_8816,N_8621,N_8651);
nand U8817 (N_8817,N_8734,N_8628);
nor U8818 (N_8818,N_8640,N_8795);
xnor U8819 (N_8819,N_8690,N_8747);
and U8820 (N_8820,N_8611,N_8659);
and U8821 (N_8821,N_8737,N_8619);
nand U8822 (N_8822,N_8647,N_8606);
nor U8823 (N_8823,N_8755,N_8781);
and U8824 (N_8824,N_8676,N_8715);
and U8825 (N_8825,N_8697,N_8752);
or U8826 (N_8826,N_8631,N_8607);
nand U8827 (N_8827,N_8763,N_8608);
xnor U8828 (N_8828,N_8787,N_8648);
xor U8829 (N_8829,N_8713,N_8644);
xor U8830 (N_8830,N_8664,N_8646);
nor U8831 (N_8831,N_8707,N_8753);
or U8832 (N_8832,N_8636,N_8638);
nand U8833 (N_8833,N_8767,N_8630);
and U8834 (N_8834,N_8788,N_8662);
or U8835 (N_8835,N_8719,N_8625);
and U8836 (N_8836,N_8600,N_8612);
xor U8837 (N_8837,N_8601,N_8658);
and U8838 (N_8838,N_8736,N_8605);
xor U8839 (N_8839,N_8750,N_8602);
or U8840 (N_8840,N_8714,N_8711);
xnor U8841 (N_8841,N_8742,N_8776);
nand U8842 (N_8842,N_8794,N_8613);
and U8843 (N_8843,N_8635,N_8603);
xor U8844 (N_8844,N_8642,N_8627);
xnor U8845 (N_8845,N_8762,N_8678);
nor U8846 (N_8846,N_8780,N_8623);
or U8847 (N_8847,N_8693,N_8679);
nand U8848 (N_8848,N_8671,N_8669);
and U8849 (N_8849,N_8670,N_8744);
xnor U8850 (N_8850,N_8754,N_8777);
and U8851 (N_8851,N_8720,N_8641);
and U8852 (N_8852,N_8774,N_8637);
xnor U8853 (N_8853,N_8687,N_8773);
or U8854 (N_8854,N_8610,N_8666);
nor U8855 (N_8855,N_8791,N_8632);
nand U8856 (N_8856,N_8768,N_8778);
nor U8857 (N_8857,N_8657,N_8717);
nand U8858 (N_8858,N_8652,N_8695);
nor U8859 (N_8859,N_8618,N_8649);
or U8860 (N_8860,N_8633,N_8796);
xor U8861 (N_8861,N_8609,N_8779);
nor U8862 (N_8862,N_8723,N_8764);
xor U8863 (N_8863,N_8615,N_8604);
nand U8864 (N_8864,N_8745,N_8739);
nor U8865 (N_8865,N_8727,N_8698);
nand U8866 (N_8866,N_8757,N_8746);
and U8867 (N_8867,N_8655,N_8616);
nor U8868 (N_8868,N_8677,N_8709);
or U8869 (N_8869,N_8748,N_8689);
nor U8870 (N_8870,N_8761,N_8721);
xor U8871 (N_8871,N_8792,N_8706);
and U8872 (N_8872,N_8674,N_8653);
xnor U8873 (N_8873,N_8691,N_8654);
nand U8874 (N_8874,N_8751,N_8650);
and U8875 (N_8875,N_8663,N_8758);
xor U8876 (N_8876,N_8710,N_8797);
nand U8877 (N_8877,N_8786,N_8738);
nand U8878 (N_8878,N_8701,N_8785);
and U8879 (N_8879,N_8694,N_8729);
or U8880 (N_8880,N_8645,N_8766);
or U8881 (N_8881,N_8614,N_8688);
and U8882 (N_8882,N_8681,N_8656);
xor U8883 (N_8883,N_8617,N_8620);
and U8884 (N_8884,N_8634,N_8784);
xnor U8885 (N_8885,N_8722,N_8798);
and U8886 (N_8886,N_8665,N_8789);
nor U8887 (N_8887,N_8680,N_8775);
and U8888 (N_8888,N_8793,N_8682);
nor U8889 (N_8889,N_8770,N_8783);
nand U8890 (N_8890,N_8700,N_8732);
and U8891 (N_8891,N_8661,N_8782);
or U8892 (N_8892,N_8684,N_8718);
and U8893 (N_8893,N_8731,N_8740);
nor U8894 (N_8894,N_8668,N_8769);
xor U8895 (N_8895,N_8759,N_8643);
nand U8896 (N_8896,N_8726,N_8667);
nor U8897 (N_8897,N_8771,N_8702);
and U8898 (N_8898,N_8624,N_8672);
nor U8899 (N_8899,N_8673,N_8728);
or U8900 (N_8900,N_8718,N_8751);
and U8901 (N_8901,N_8711,N_8746);
or U8902 (N_8902,N_8709,N_8634);
and U8903 (N_8903,N_8661,N_8642);
xor U8904 (N_8904,N_8694,N_8673);
or U8905 (N_8905,N_8753,N_8613);
nor U8906 (N_8906,N_8677,N_8731);
nor U8907 (N_8907,N_8770,N_8746);
nor U8908 (N_8908,N_8744,N_8787);
xor U8909 (N_8909,N_8676,N_8773);
nor U8910 (N_8910,N_8769,N_8674);
nand U8911 (N_8911,N_8752,N_8702);
or U8912 (N_8912,N_8628,N_8669);
and U8913 (N_8913,N_8637,N_8690);
nor U8914 (N_8914,N_8737,N_8657);
or U8915 (N_8915,N_8618,N_8669);
and U8916 (N_8916,N_8752,N_8622);
or U8917 (N_8917,N_8700,N_8753);
and U8918 (N_8918,N_8723,N_8671);
or U8919 (N_8919,N_8717,N_8753);
nand U8920 (N_8920,N_8720,N_8655);
xor U8921 (N_8921,N_8603,N_8704);
and U8922 (N_8922,N_8708,N_8712);
nand U8923 (N_8923,N_8796,N_8644);
nand U8924 (N_8924,N_8788,N_8654);
or U8925 (N_8925,N_8742,N_8677);
nor U8926 (N_8926,N_8716,N_8789);
and U8927 (N_8927,N_8669,N_8690);
nor U8928 (N_8928,N_8736,N_8780);
nor U8929 (N_8929,N_8638,N_8785);
nand U8930 (N_8930,N_8797,N_8679);
or U8931 (N_8931,N_8779,N_8741);
nand U8932 (N_8932,N_8754,N_8610);
xor U8933 (N_8933,N_8756,N_8740);
nor U8934 (N_8934,N_8646,N_8730);
nand U8935 (N_8935,N_8742,N_8642);
xor U8936 (N_8936,N_8642,N_8704);
xnor U8937 (N_8937,N_8648,N_8732);
nor U8938 (N_8938,N_8630,N_8665);
xnor U8939 (N_8939,N_8756,N_8739);
and U8940 (N_8940,N_8755,N_8663);
or U8941 (N_8941,N_8625,N_8612);
xnor U8942 (N_8942,N_8628,N_8722);
nand U8943 (N_8943,N_8712,N_8682);
or U8944 (N_8944,N_8758,N_8612);
nand U8945 (N_8945,N_8677,N_8609);
nand U8946 (N_8946,N_8727,N_8670);
and U8947 (N_8947,N_8797,N_8620);
nand U8948 (N_8948,N_8608,N_8616);
nand U8949 (N_8949,N_8791,N_8639);
nand U8950 (N_8950,N_8787,N_8607);
nand U8951 (N_8951,N_8738,N_8790);
xnor U8952 (N_8952,N_8713,N_8684);
and U8953 (N_8953,N_8645,N_8735);
nand U8954 (N_8954,N_8691,N_8673);
xnor U8955 (N_8955,N_8625,N_8790);
or U8956 (N_8956,N_8755,N_8646);
xor U8957 (N_8957,N_8675,N_8660);
nand U8958 (N_8958,N_8693,N_8708);
and U8959 (N_8959,N_8671,N_8716);
xnor U8960 (N_8960,N_8673,N_8686);
and U8961 (N_8961,N_8606,N_8724);
or U8962 (N_8962,N_8628,N_8666);
nor U8963 (N_8963,N_8758,N_8625);
and U8964 (N_8964,N_8656,N_8646);
or U8965 (N_8965,N_8638,N_8731);
nor U8966 (N_8966,N_8683,N_8610);
nor U8967 (N_8967,N_8600,N_8710);
nor U8968 (N_8968,N_8627,N_8663);
nor U8969 (N_8969,N_8636,N_8712);
and U8970 (N_8970,N_8610,N_8698);
nor U8971 (N_8971,N_8630,N_8642);
nor U8972 (N_8972,N_8711,N_8724);
xnor U8973 (N_8973,N_8703,N_8632);
xor U8974 (N_8974,N_8794,N_8672);
and U8975 (N_8975,N_8737,N_8637);
nand U8976 (N_8976,N_8674,N_8627);
xor U8977 (N_8977,N_8606,N_8622);
xnor U8978 (N_8978,N_8648,N_8675);
xor U8979 (N_8979,N_8692,N_8762);
nor U8980 (N_8980,N_8648,N_8786);
nand U8981 (N_8981,N_8620,N_8734);
xnor U8982 (N_8982,N_8601,N_8778);
and U8983 (N_8983,N_8664,N_8683);
nor U8984 (N_8984,N_8642,N_8764);
or U8985 (N_8985,N_8773,N_8707);
or U8986 (N_8986,N_8710,N_8732);
nor U8987 (N_8987,N_8603,N_8612);
and U8988 (N_8988,N_8766,N_8647);
nor U8989 (N_8989,N_8717,N_8627);
or U8990 (N_8990,N_8756,N_8720);
or U8991 (N_8991,N_8770,N_8703);
and U8992 (N_8992,N_8796,N_8665);
or U8993 (N_8993,N_8782,N_8790);
nor U8994 (N_8994,N_8679,N_8716);
or U8995 (N_8995,N_8684,N_8609);
and U8996 (N_8996,N_8700,N_8781);
and U8997 (N_8997,N_8607,N_8647);
or U8998 (N_8998,N_8613,N_8630);
nor U8999 (N_8999,N_8777,N_8747);
or U9000 (N_9000,N_8870,N_8823);
nor U9001 (N_9001,N_8841,N_8869);
or U9002 (N_9002,N_8940,N_8983);
nor U9003 (N_9003,N_8881,N_8846);
nor U9004 (N_9004,N_8891,N_8812);
xor U9005 (N_9005,N_8908,N_8906);
and U9006 (N_9006,N_8897,N_8920);
nand U9007 (N_9007,N_8919,N_8883);
xnor U9008 (N_9008,N_8804,N_8921);
nor U9009 (N_9009,N_8987,N_8813);
nand U9010 (N_9010,N_8877,N_8917);
and U9011 (N_9011,N_8997,N_8829);
nand U9012 (N_9012,N_8949,N_8950);
nand U9013 (N_9013,N_8972,N_8857);
or U9014 (N_9014,N_8884,N_8901);
nand U9015 (N_9015,N_8975,N_8887);
nor U9016 (N_9016,N_8918,N_8827);
or U9017 (N_9017,N_8970,N_8900);
or U9018 (N_9018,N_8939,N_8902);
nand U9019 (N_9019,N_8895,N_8933);
xor U9020 (N_9020,N_8811,N_8926);
xor U9021 (N_9021,N_8816,N_8929);
xor U9022 (N_9022,N_8872,N_8814);
nand U9023 (N_9023,N_8968,N_8867);
nand U9024 (N_9024,N_8899,N_8953);
and U9025 (N_9025,N_8938,N_8892);
nor U9026 (N_9026,N_8992,N_8834);
and U9027 (N_9027,N_8858,N_8828);
xnor U9028 (N_9028,N_8805,N_8952);
and U9029 (N_9029,N_8890,N_8948);
or U9030 (N_9030,N_8954,N_8896);
or U9031 (N_9031,N_8982,N_8893);
nand U9032 (N_9032,N_8910,N_8862);
and U9033 (N_9033,N_8973,N_8946);
xnor U9034 (N_9034,N_8989,N_8830);
or U9035 (N_9035,N_8807,N_8980);
xnor U9036 (N_9036,N_8976,N_8889);
or U9037 (N_9037,N_8935,N_8836);
or U9038 (N_9038,N_8874,N_8961);
nand U9039 (N_9039,N_8923,N_8904);
or U9040 (N_9040,N_8821,N_8873);
or U9041 (N_9041,N_8863,N_8966);
nor U9042 (N_9042,N_8817,N_8964);
nand U9043 (N_9043,N_8850,N_8859);
nor U9044 (N_9044,N_8865,N_8969);
xnor U9045 (N_9045,N_8925,N_8951);
nand U9046 (N_9046,N_8916,N_8994);
xnor U9047 (N_9047,N_8839,N_8924);
nor U9048 (N_9048,N_8934,N_8922);
or U9049 (N_9049,N_8942,N_8871);
xnor U9050 (N_9050,N_8844,N_8837);
and U9051 (N_9051,N_8998,N_8803);
nand U9052 (N_9052,N_8988,N_8856);
xor U9053 (N_9053,N_8886,N_8944);
or U9054 (N_9054,N_8932,N_8941);
nand U9055 (N_9055,N_8984,N_8981);
nor U9056 (N_9056,N_8840,N_8815);
nand U9057 (N_9057,N_8928,N_8855);
nand U9058 (N_9058,N_8835,N_8957);
nor U9059 (N_9059,N_8956,N_8894);
nor U9060 (N_9060,N_8930,N_8931);
and U9061 (N_9061,N_8838,N_8854);
xor U9062 (N_9062,N_8878,N_8912);
nand U9063 (N_9063,N_8971,N_8801);
xor U9064 (N_9064,N_8945,N_8985);
and U9065 (N_9065,N_8875,N_8960);
and U9066 (N_9066,N_8962,N_8911);
and U9067 (N_9067,N_8955,N_8820);
nor U9068 (N_9068,N_8879,N_8866);
and U9069 (N_9069,N_8808,N_8907);
and U9070 (N_9070,N_8885,N_8991);
or U9071 (N_9071,N_8965,N_8888);
and U9072 (N_9072,N_8903,N_8963);
xor U9073 (N_9073,N_8826,N_8818);
and U9074 (N_9074,N_8979,N_8915);
or U9075 (N_9075,N_8898,N_8847);
xnor U9076 (N_9076,N_8882,N_8905);
nor U9077 (N_9077,N_8937,N_8851);
nor U9078 (N_9078,N_8832,N_8990);
and U9079 (N_9079,N_8876,N_8810);
nand U9080 (N_9080,N_8864,N_8802);
xnor U9081 (N_9081,N_8986,N_8978);
nand U9082 (N_9082,N_8947,N_8999);
xnor U9083 (N_9083,N_8861,N_8927);
xnor U9084 (N_9084,N_8800,N_8974);
nor U9085 (N_9085,N_8860,N_8809);
nor U9086 (N_9086,N_8868,N_8996);
nand U9087 (N_9087,N_8852,N_8959);
or U9088 (N_9088,N_8995,N_8806);
nor U9089 (N_9089,N_8842,N_8943);
nand U9090 (N_9090,N_8977,N_8845);
xnor U9091 (N_9091,N_8909,N_8848);
nor U9092 (N_9092,N_8936,N_8914);
or U9093 (N_9093,N_8822,N_8819);
xor U9094 (N_9094,N_8880,N_8833);
nor U9095 (N_9095,N_8913,N_8831);
xnor U9096 (N_9096,N_8958,N_8853);
or U9097 (N_9097,N_8843,N_8825);
nor U9098 (N_9098,N_8824,N_8993);
or U9099 (N_9099,N_8967,N_8849);
or U9100 (N_9100,N_8903,N_8962);
or U9101 (N_9101,N_8903,N_8893);
and U9102 (N_9102,N_8882,N_8952);
nand U9103 (N_9103,N_8808,N_8809);
or U9104 (N_9104,N_8940,N_8883);
nand U9105 (N_9105,N_8839,N_8865);
and U9106 (N_9106,N_8825,N_8891);
and U9107 (N_9107,N_8927,N_8988);
or U9108 (N_9108,N_8808,N_8948);
nor U9109 (N_9109,N_8958,N_8980);
nor U9110 (N_9110,N_8833,N_8967);
and U9111 (N_9111,N_8939,N_8819);
and U9112 (N_9112,N_8895,N_8988);
and U9113 (N_9113,N_8916,N_8889);
nand U9114 (N_9114,N_8926,N_8840);
or U9115 (N_9115,N_8983,N_8958);
nand U9116 (N_9116,N_8884,N_8886);
nand U9117 (N_9117,N_8953,N_8853);
xor U9118 (N_9118,N_8837,N_8891);
nand U9119 (N_9119,N_8934,N_8925);
xor U9120 (N_9120,N_8838,N_8933);
xnor U9121 (N_9121,N_8961,N_8992);
xnor U9122 (N_9122,N_8927,N_8835);
or U9123 (N_9123,N_8801,N_8998);
xor U9124 (N_9124,N_8890,N_8844);
xor U9125 (N_9125,N_8919,N_8999);
or U9126 (N_9126,N_8800,N_8841);
xnor U9127 (N_9127,N_8884,N_8816);
xnor U9128 (N_9128,N_8827,N_8968);
or U9129 (N_9129,N_8934,N_8979);
and U9130 (N_9130,N_8804,N_8858);
xor U9131 (N_9131,N_8882,N_8927);
nor U9132 (N_9132,N_8963,N_8916);
nand U9133 (N_9133,N_8984,N_8987);
nor U9134 (N_9134,N_8841,N_8805);
nand U9135 (N_9135,N_8949,N_8880);
and U9136 (N_9136,N_8867,N_8826);
nand U9137 (N_9137,N_8889,N_8913);
and U9138 (N_9138,N_8936,N_8991);
or U9139 (N_9139,N_8859,N_8867);
or U9140 (N_9140,N_8874,N_8963);
or U9141 (N_9141,N_8909,N_8829);
or U9142 (N_9142,N_8836,N_8927);
xnor U9143 (N_9143,N_8941,N_8827);
nor U9144 (N_9144,N_8872,N_8893);
or U9145 (N_9145,N_8996,N_8999);
nor U9146 (N_9146,N_8959,N_8855);
xnor U9147 (N_9147,N_8845,N_8889);
nand U9148 (N_9148,N_8850,N_8855);
nor U9149 (N_9149,N_8892,N_8887);
or U9150 (N_9150,N_8832,N_8989);
nor U9151 (N_9151,N_8977,N_8998);
nor U9152 (N_9152,N_8828,N_8995);
and U9153 (N_9153,N_8838,N_8986);
xnor U9154 (N_9154,N_8960,N_8872);
xor U9155 (N_9155,N_8805,N_8827);
xor U9156 (N_9156,N_8876,N_8806);
or U9157 (N_9157,N_8863,N_8923);
or U9158 (N_9158,N_8864,N_8987);
xnor U9159 (N_9159,N_8848,N_8857);
xnor U9160 (N_9160,N_8838,N_8966);
xnor U9161 (N_9161,N_8996,N_8802);
nor U9162 (N_9162,N_8992,N_8822);
or U9163 (N_9163,N_8869,N_8804);
and U9164 (N_9164,N_8811,N_8879);
and U9165 (N_9165,N_8968,N_8808);
xnor U9166 (N_9166,N_8860,N_8874);
nor U9167 (N_9167,N_8804,N_8814);
nand U9168 (N_9168,N_8931,N_8986);
or U9169 (N_9169,N_8940,N_8927);
or U9170 (N_9170,N_8919,N_8945);
nor U9171 (N_9171,N_8879,N_8818);
nand U9172 (N_9172,N_8834,N_8867);
nor U9173 (N_9173,N_8995,N_8983);
nand U9174 (N_9174,N_8853,N_8806);
and U9175 (N_9175,N_8878,N_8892);
or U9176 (N_9176,N_8801,N_8937);
or U9177 (N_9177,N_8902,N_8946);
or U9178 (N_9178,N_8972,N_8974);
nand U9179 (N_9179,N_8860,N_8892);
and U9180 (N_9180,N_8818,N_8903);
nand U9181 (N_9181,N_8948,N_8838);
nor U9182 (N_9182,N_8953,N_8837);
xnor U9183 (N_9183,N_8831,N_8820);
nor U9184 (N_9184,N_8970,N_8879);
and U9185 (N_9185,N_8802,N_8891);
or U9186 (N_9186,N_8827,N_8923);
and U9187 (N_9187,N_8938,N_8935);
xnor U9188 (N_9188,N_8834,N_8825);
xnor U9189 (N_9189,N_8817,N_8919);
and U9190 (N_9190,N_8846,N_8971);
nand U9191 (N_9191,N_8855,N_8938);
nand U9192 (N_9192,N_8974,N_8825);
nor U9193 (N_9193,N_8898,N_8901);
or U9194 (N_9194,N_8979,N_8960);
and U9195 (N_9195,N_8933,N_8815);
and U9196 (N_9196,N_8974,N_8952);
and U9197 (N_9197,N_8878,N_8984);
nand U9198 (N_9198,N_8985,N_8962);
or U9199 (N_9199,N_8839,N_8968);
xor U9200 (N_9200,N_9177,N_9119);
nand U9201 (N_9201,N_9058,N_9101);
and U9202 (N_9202,N_9013,N_9027);
xor U9203 (N_9203,N_9014,N_9114);
nor U9204 (N_9204,N_9034,N_9173);
xnor U9205 (N_9205,N_9070,N_9039);
nand U9206 (N_9206,N_9146,N_9126);
and U9207 (N_9207,N_9127,N_9011);
nor U9208 (N_9208,N_9064,N_9046);
xor U9209 (N_9209,N_9047,N_9091);
nand U9210 (N_9210,N_9017,N_9163);
xnor U9211 (N_9211,N_9158,N_9079);
nor U9212 (N_9212,N_9144,N_9107);
and U9213 (N_9213,N_9097,N_9065);
and U9214 (N_9214,N_9069,N_9080);
xor U9215 (N_9215,N_9197,N_9129);
xnor U9216 (N_9216,N_9136,N_9118);
nor U9217 (N_9217,N_9137,N_9054);
or U9218 (N_9218,N_9141,N_9196);
nor U9219 (N_9219,N_9010,N_9115);
nor U9220 (N_9220,N_9139,N_9074);
nand U9221 (N_9221,N_9019,N_9186);
or U9222 (N_9222,N_9135,N_9111);
nor U9223 (N_9223,N_9008,N_9155);
xnor U9224 (N_9224,N_9134,N_9169);
and U9225 (N_9225,N_9116,N_9153);
xnor U9226 (N_9226,N_9007,N_9143);
nand U9227 (N_9227,N_9145,N_9188);
nor U9228 (N_9228,N_9002,N_9084);
nor U9229 (N_9229,N_9168,N_9049);
nand U9230 (N_9230,N_9082,N_9176);
and U9231 (N_9231,N_9192,N_9181);
or U9232 (N_9232,N_9160,N_9006);
nor U9233 (N_9233,N_9040,N_9043);
xnor U9234 (N_9234,N_9128,N_9175);
nand U9235 (N_9235,N_9193,N_9122);
nor U9236 (N_9236,N_9053,N_9178);
or U9237 (N_9237,N_9104,N_9103);
nor U9238 (N_9238,N_9190,N_9105);
or U9239 (N_9239,N_9081,N_9066);
or U9240 (N_9240,N_9140,N_9045);
nand U9241 (N_9241,N_9033,N_9093);
xor U9242 (N_9242,N_9113,N_9121);
and U9243 (N_9243,N_9072,N_9162);
nand U9244 (N_9244,N_9003,N_9077);
nor U9245 (N_9245,N_9159,N_9183);
nand U9246 (N_9246,N_9021,N_9016);
and U9247 (N_9247,N_9094,N_9032);
or U9248 (N_9248,N_9063,N_9130);
nor U9249 (N_9249,N_9018,N_9059);
nor U9250 (N_9250,N_9012,N_9184);
nand U9251 (N_9251,N_9123,N_9044);
nor U9252 (N_9252,N_9075,N_9152);
xor U9253 (N_9253,N_9089,N_9071);
xnor U9254 (N_9254,N_9055,N_9038);
nand U9255 (N_9255,N_9004,N_9199);
nand U9256 (N_9256,N_9198,N_9023);
nor U9257 (N_9257,N_9087,N_9167);
nand U9258 (N_9258,N_9161,N_9078);
or U9259 (N_9259,N_9138,N_9106);
nor U9260 (N_9260,N_9048,N_9131);
or U9261 (N_9261,N_9124,N_9088);
and U9262 (N_9262,N_9024,N_9076);
and U9263 (N_9263,N_9157,N_9098);
nor U9264 (N_9264,N_9149,N_9100);
and U9265 (N_9265,N_9000,N_9099);
xnor U9266 (N_9266,N_9005,N_9051);
xor U9267 (N_9267,N_9185,N_9170);
and U9268 (N_9268,N_9147,N_9028);
and U9269 (N_9269,N_9179,N_9086);
or U9270 (N_9270,N_9110,N_9120);
nand U9271 (N_9271,N_9029,N_9022);
and U9272 (N_9272,N_9154,N_9117);
nor U9273 (N_9273,N_9165,N_9085);
nand U9274 (N_9274,N_9096,N_9057);
nand U9275 (N_9275,N_9194,N_9166);
and U9276 (N_9276,N_9025,N_9095);
and U9277 (N_9277,N_9102,N_9151);
xnor U9278 (N_9278,N_9150,N_9191);
and U9279 (N_9279,N_9171,N_9180);
nor U9280 (N_9280,N_9015,N_9068);
xnor U9281 (N_9281,N_9030,N_9037);
nand U9282 (N_9282,N_9035,N_9112);
or U9283 (N_9283,N_9187,N_9108);
and U9284 (N_9284,N_9182,N_9083);
nor U9285 (N_9285,N_9026,N_9092);
xor U9286 (N_9286,N_9132,N_9073);
and U9287 (N_9287,N_9142,N_9148);
or U9288 (N_9288,N_9125,N_9133);
nor U9289 (N_9289,N_9041,N_9164);
and U9290 (N_9290,N_9009,N_9020);
nor U9291 (N_9291,N_9036,N_9060);
or U9292 (N_9292,N_9172,N_9001);
xor U9293 (N_9293,N_9056,N_9174);
xor U9294 (N_9294,N_9050,N_9067);
or U9295 (N_9295,N_9031,N_9062);
xor U9296 (N_9296,N_9052,N_9156);
nand U9297 (N_9297,N_9090,N_9042);
nor U9298 (N_9298,N_9061,N_9109);
nor U9299 (N_9299,N_9195,N_9189);
or U9300 (N_9300,N_9068,N_9192);
or U9301 (N_9301,N_9140,N_9092);
xor U9302 (N_9302,N_9177,N_9105);
nor U9303 (N_9303,N_9102,N_9047);
nor U9304 (N_9304,N_9010,N_9002);
nand U9305 (N_9305,N_9122,N_9007);
nand U9306 (N_9306,N_9112,N_9078);
and U9307 (N_9307,N_9095,N_9188);
and U9308 (N_9308,N_9010,N_9111);
xnor U9309 (N_9309,N_9175,N_9035);
xor U9310 (N_9310,N_9066,N_9099);
nand U9311 (N_9311,N_9168,N_9172);
nand U9312 (N_9312,N_9001,N_9162);
xnor U9313 (N_9313,N_9056,N_9102);
or U9314 (N_9314,N_9113,N_9194);
and U9315 (N_9315,N_9003,N_9192);
nand U9316 (N_9316,N_9112,N_9184);
nor U9317 (N_9317,N_9125,N_9051);
or U9318 (N_9318,N_9009,N_9033);
or U9319 (N_9319,N_9064,N_9119);
and U9320 (N_9320,N_9086,N_9055);
xor U9321 (N_9321,N_9052,N_9149);
and U9322 (N_9322,N_9149,N_9058);
xor U9323 (N_9323,N_9009,N_9034);
nor U9324 (N_9324,N_9135,N_9126);
or U9325 (N_9325,N_9104,N_9131);
or U9326 (N_9326,N_9049,N_9137);
xor U9327 (N_9327,N_9102,N_9051);
or U9328 (N_9328,N_9190,N_9058);
nand U9329 (N_9329,N_9159,N_9107);
nand U9330 (N_9330,N_9044,N_9020);
xor U9331 (N_9331,N_9059,N_9171);
nor U9332 (N_9332,N_9059,N_9084);
xor U9333 (N_9333,N_9022,N_9153);
and U9334 (N_9334,N_9045,N_9127);
or U9335 (N_9335,N_9116,N_9007);
xor U9336 (N_9336,N_9113,N_9177);
xnor U9337 (N_9337,N_9092,N_9106);
nand U9338 (N_9338,N_9155,N_9003);
xor U9339 (N_9339,N_9100,N_9150);
nand U9340 (N_9340,N_9089,N_9054);
xnor U9341 (N_9341,N_9189,N_9115);
xor U9342 (N_9342,N_9113,N_9010);
or U9343 (N_9343,N_9153,N_9011);
nor U9344 (N_9344,N_9182,N_9043);
nor U9345 (N_9345,N_9118,N_9025);
nor U9346 (N_9346,N_9080,N_9136);
nand U9347 (N_9347,N_9140,N_9165);
or U9348 (N_9348,N_9083,N_9128);
and U9349 (N_9349,N_9184,N_9071);
nor U9350 (N_9350,N_9189,N_9136);
xor U9351 (N_9351,N_9014,N_9153);
nand U9352 (N_9352,N_9106,N_9032);
nand U9353 (N_9353,N_9108,N_9075);
nor U9354 (N_9354,N_9045,N_9189);
xnor U9355 (N_9355,N_9177,N_9037);
xor U9356 (N_9356,N_9197,N_9062);
nor U9357 (N_9357,N_9135,N_9092);
or U9358 (N_9358,N_9121,N_9093);
xor U9359 (N_9359,N_9167,N_9165);
and U9360 (N_9360,N_9009,N_9149);
nor U9361 (N_9361,N_9005,N_9189);
or U9362 (N_9362,N_9180,N_9076);
nor U9363 (N_9363,N_9166,N_9183);
xor U9364 (N_9364,N_9115,N_9020);
xnor U9365 (N_9365,N_9173,N_9116);
or U9366 (N_9366,N_9073,N_9003);
or U9367 (N_9367,N_9086,N_9085);
and U9368 (N_9368,N_9050,N_9087);
xor U9369 (N_9369,N_9063,N_9140);
nor U9370 (N_9370,N_9173,N_9198);
and U9371 (N_9371,N_9006,N_9116);
nand U9372 (N_9372,N_9169,N_9184);
nor U9373 (N_9373,N_9007,N_9040);
nand U9374 (N_9374,N_9069,N_9178);
or U9375 (N_9375,N_9104,N_9021);
nand U9376 (N_9376,N_9132,N_9037);
xnor U9377 (N_9377,N_9053,N_9145);
nor U9378 (N_9378,N_9166,N_9028);
xor U9379 (N_9379,N_9137,N_9091);
and U9380 (N_9380,N_9027,N_9076);
xnor U9381 (N_9381,N_9101,N_9193);
and U9382 (N_9382,N_9174,N_9018);
and U9383 (N_9383,N_9157,N_9017);
nand U9384 (N_9384,N_9156,N_9131);
xnor U9385 (N_9385,N_9176,N_9034);
and U9386 (N_9386,N_9110,N_9169);
nand U9387 (N_9387,N_9140,N_9154);
nor U9388 (N_9388,N_9128,N_9073);
or U9389 (N_9389,N_9154,N_9058);
nor U9390 (N_9390,N_9173,N_9057);
nand U9391 (N_9391,N_9062,N_9140);
xor U9392 (N_9392,N_9112,N_9070);
nor U9393 (N_9393,N_9135,N_9183);
nor U9394 (N_9394,N_9174,N_9012);
nand U9395 (N_9395,N_9159,N_9116);
and U9396 (N_9396,N_9067,N_9053);
or U9397 (N_9397,N_9145,N_9042);
or U9398 (N_9398,N_9187,N_9101);
and U9399 (N_9399,N_9117,N_9127);
and U9400 (N_9400,N_9216,N_9244);
nand U9401 (N_9401,N_9324,N_9349);
nand U9402 (N_9402,N_9284,N_9378);
or U9403 (N_9403,N_9297,N_9214);
and U9404 (N_9404,N_9335,N_9341);
nor U9405 (N_9405,N_9316,N_9203);
or U9406 (N_9406,N_9243,N_9328);
and U9407 (N_9407,N_9356,N_9289);
nor U9408 (N_9408,N_9217,N_9200);
and U9409 (N_9409,N_9248,N_9241);
nor U9410 (N_9410,N_9242,N_9322);
or U9411 (N_9411,N_9372,N_9210);
nand U9412 (N_9412,N_9206,N_9262);
nand U9413 (N_9413,N_9299,N_9336);
and U9414 (N_9414,N_9360,N_9279);
and U9415 (N_9415,N_9309,N_9268);
nor U9416 (N_9416,N_9264,N_9325);
and U9417 (N_9417,N_9307,N_9333);
or U9418 (N_9418,N_9290,N_9386);
and U9419 (N_9419,N_9301,N_9267);
and U9420 (N_9420,N_9375,N_9390);
nor U9421 (N_9421,N_9215,N_9276);
and U9422 (N_9422,N_9394,N_9338);
xor U9423 (N_9423,N_9293,N_9318);
nor U9424 (N_9424,N_9227,N_9342);
nand U9425 (N_9425,N_9205,N_9397);
nand U9426 (N_9426,N_9332,N_9339);
xnor U9427 (N_9427,N_9229,N_9317);
nor U9428 (N_9428,N_9347,N_9296);
and U9429 (N_9429,N_9234,N_9209);
and U9430 (N_9430,N_9388,N_9250);
nor U9431 (N_9431,N_9365,N_9272);
nand U9432 (N_9432,N_9269,N_9384);
or U9433 (N_9433,N_9399,N_9257);
nor U9434 (N_9434,N_9329,N_9270);
nor U9435 (N_9435,N_9396,N_9208);
nand U9436 (N_9436,N_9369,N_9213);
or U9437 (N_9437,N_9238,N_9260);
xnor U9438 (N_9438,N_9352,N_9358);
or U9439 (N_9439,N_9280,N_9344);
and U9440 (N_9440,N_9334,N_9246);
and U9441 (N_9441,N_9380,N_9298);
and U9442 (N_9442,N_9256,N_9273);
xor U9443 (N_9443,N_9259,N_9212);
nand U9444 (N_9444,N_9252,N_9258);
nor U9445 (N_9445,N_9359,N_9314);
and U9446 (N_9446,N_9211,N_9362);
xor U9447 (N_9447,N_9236,N_9286);
xor U9448 (N_9448,N_9337,N_9232);
and U9449 (N_9449,N_9207,N_9265);
nand U9450 (N_9450,N_9326,N_9278);
or U9451 (N_9451,N_9228,N_9249);
nor U9452 (N_9452,N_9308,N_9281);
and U9453 (N_9453,N_9225,N_9287);
xnor U9454 (N_9454,N_9222,N_9354);
nand U9455 (N_9455,N_9240,N_9391);
or U9456 (N_9456,N_9323,N_9368);
and U9457 (N_9457,N_9351,N_9366);
and U9458 (N_9458,N_9294,N_9320);
xor U9459 (N_9459,N_9377,N_9285);
nand U9460 (N_9460,N_9266,N_9305);
or U9461 (N_9461,N_9376,N_9319);
and U9462 (N_9462,N_9371,N_9271);
and U9463 (N_9463,N_9370,N_9304);
xnor U9464 (N_9464,N_9350,N_9306);
or U9465 (N_9465,N_9288,N_9361);
nand U9466 (N_9466,N_9364,N_9235);
xnor U9467 (N_9467,N_9311,N_9381);
nand U9468 (N_9468,N_9226,N_9389);
and U9469 (N_9469,N_9255,N_9395);
xor U9470 (N_9470,N_9313,N_9218);
or U9471 (N_9471,N_9254,N_9382);
nand U9472 (N_9472,N_9221,N_9363);
xnor U9473 (N_9473,N_9295,N_9330);
and U9474 (N_9474,N_9202,N_9204);
nand U9475 (N_9475,N_9223,N_9348);
or U9476 (N_9476,N_9321,N_9261);
or U9477 (N_9477,N_9275,N_9251);
xnor U9478 (N_9478,N_9282,N_9392);
nand U9479 (N_9479,N_9283,N_9303);
xnor U9480 (N_9480,N_9277,N_9233);
and U9481 (N_9481,N_9263,N_9230);
or U9482 (N_9482,N_9331,N_9292);
nand U9483 (N_9483,N_9387,N_9231);
and U9484 (N_9484,N_9355,N_9201);
or U9485 (N_9485,N_9239,N_9357);
and U9486 (N_9486,N_9302,N_9237);
nand U9487 (N_9487,N_9393,N_9373);
xnor U9488 (N_9488,N_9343,N_9310);
and U9489 (N_9489,N_9274,N_9253);
or U9490 (N_9490,N_9379,N_9398);
nand U9491 (N_9491,N_9300,N_9385);
and U9492 (N_9492,N_9345,N_9383);
xor U9493 (N_9493,N_9340,N_9224);
or U9494 (N_9494,N_9312,N_9220);
nor U9495 (N_9495,N_9219,N_9291);
xnor U9496 (N_9496,N_9247,N_9315);
and U9497 (N_9497,N_9346,N_9367);
xor U9498 (N_9498,N_9374,N_9327);
nor U9499 (N_9499,N_9353,N_9245);
nand U9500 (N_9500,N_9250,N_9340);
nand U9501 (N_9501,N_9347,N_9295);
nor U9502 (N_9502,N_9283,N_9216);
nand U9503 (N_9503,N_9393,N_9320);
and U9504 (N_9504,N_9263,N_9391);
or U9505 (N_9505,N_9373,N_9245);
xor U9506 (N_9506,N_9244,N_9345);
and U9507 (N_9507,N_9379,N_9364);
and U9508 (N_9508,N_9327,N_9324);
or U9509 (N_9509,N_9206,N_9387);
nor U9510 (N_9510,N_9201,N_9369);
xnor U9511 (N_9511,N_9239,N_9310);
nor U9512 (N_9512,N_9333,N_9253);
or U9513 (N_9513,N_9279,N_9213);
or U9514 (N_9514,N_9236,N_9215);
or U9515 (N_9515,N_9222,N_9320);
nor U9516 (N_9516,N_9283,N_9360);
and U9517 (N_9517,N_9322,N_9275);
and U9518 (N_9518,N_9303,N_9202);
nor U9519 (N_9519,N_9212,N_9382);
and U9520 (N_9520,N_9233,N_9267);
and U9521 (N_9521,N_9247,N_9251);
and U9522 (N_9522,N_9234,N_9228);
or U9523 (N_9523,N_9367,N_9386);
and U9524 (N_9524,N_9218,N_9242);
and U9525 (N_9525,N_9284,N_9380);
nor U9526 (N_9526,N_9295,N_9283);
xor U9527 (N_9527,N_9310,N_9313);
and U9528 (N_9528,N_9307,N_9226);
nand U9529 (N_9529,N_9346,N_9276);
nor U9530 (N_9530,N_9264,N_9224);
and U9531 (N_9531,N_9382,N_9349);
or U9532 (N_9532,N_9219,N_9321);
xnor U9533 (N_9533,N_9372,N_9245);
and U9534 (N_9534,N_9233,N_9228);
or U9535 (N_9535,N_9315,N_9242);
nor U9536 (N_9536,N_9226,N_9310);
or U9537 (N_9537,N_9209,N_9302);
xor U9538 (N_9538,N_9262,N_9204);
xnor U9539 (N_9539,N_9224,N_9267);
nor U9540 (N_9540,N_9344,N_9325);
or U9541 (N_9541,N_9377,N_9225);
and U9542 (N_9542,N_9341,N_9330);
nand U9543 (N_9543,N_9237,N_9256);
and U9544 (N_9544,N_9337,N_9295);
xnor U9545 (N_9545,N_9263,N_9397);
xnor U9546 (N_9546,N_9259,N_9298);
nor U9547 (N_9547,N_9316,N_9331);
or U9548 (N_9548,N_9207,N_9340);
xor U9549 (N_9549,N_9215,N_9390);
and U9550 (N_9550,N_9373,N_9312);
nor U9551 (N_9551,N_9382,N_9335);
and U9552 (N_9552,N_9396,N_9278);
and U9553 (N_9553,N_9287,N_9364);
nand U9554 (N_9554,N_9255,N_9307);
or U9555 (N_9555,N_9387,N_9318);
xnor U9556 (N_9556,N_9261,N_9207);
and U9557 (N_9557,N_9264,N_9398);
xor U9558 (N_9558,N_9352,N_9260);
or U9559 (N_9559,N_9245,N_9236);
xor U9560 (N_9560,N_9278,N_9376);
nand U9561 (N_9561,N_9278,N_9285);
or U9562 (N_9562,N_9382,N_9259);
or U9563 (N_9563,N_9251,N_9242);
nand U9564 (N_9564,N_9257,N_9302);
and U9565 (N_9565,N_9289,N_9337);
nand U9566 (N_9566,N_9323,N_9244);
or U9567 (N_9567,N_9376,N_9233);
and U9568 (N_9568,N_9304,N_9279);
xnor U9569 (N_9569,N_9274,N_9285);
and U9570 (N_9570,N_9245,N_9347);
and U9571 (N_9571,N_9357,N_9275);
nand U9572 (N_9572,N_9353,N_9220);
or U9573 (N_9573,N_9324,N_9388);
xor U9574 (N_9574,N_9220,N_9260);
xor U9575 (N_9575,N_9384,N_9279);
nand U9576 (N_9576,N_9378,N_9325);
xnor U9577 (N_9577,N_9311,N_9242);
and U9578 (N_9578,N_9342,N_9213);
nor U9579 (N_9579,N_9359,N_9338);
nor U9580 (N_9580,N_9302,N_9208);
and U9581 (N_9581,N_9265,N_9345);
xor U9582 (N_9582,N_9294,N_9289);
and U9583 (N_9583,N_9364,N_9384);
xnor U9584 (N_9584,N_9345,N_9302);
or U9585 (N_9585,N_9358,N_9380);
nand U9586 (N_9586,N_9329,N_9207);
and U9587 (N_9587,N_9319,N_9296);
nor U9588 (N_9588,N_9263,N_9211);
and U9589 (N_9589,N_9372,N_9381);
or U9590 (N_9590,N_9399,N_9270);
nor U9591 (N_9591,N_9387,N_9329);
and U9592 (N_9592,N_9365,N_9386);
xor U9593 (N_9593,N_9362,N_9304);
and U9594 (N_9594,N_9207,N_9334);
and U9595 (N_9595,N_9255,N_9209);
nand U9596 (N_9596,N_9245,N_9314);
xnor U9597 (N_9597,N_9240,N_9239);
or U9598 (N_9598,N_9293,N_9347);
nand U9599 (N_9599,N_9339,N_9279);
nor U9600 (N_9600,N_9551,N_9564);
or U9601 (N_9601,N_9456,N_9583);
or U9602 (N_9602,N_9473,N_9404);
nand U9603 (N_9603,N_9496,N_9453);
nand U9604 (N_9604,N_9421,N_9585);
nor U9605 (N_9605,N_9517,N_9470);
nor U9606 (N_9606,N_9490,N_9498);
nand U9607 (N_9607,N_9539,N_9546);
xnor U9608 (N_9608,N_9523,N_9464);
nand U9609 (N_9609,N_9543,N_9499);
xnor U9610 (N_9610,N_9485,N_9514);
or U9611 (N_9611,N_9589,N_9418);
and U9612 (N_9612,N_9483,N_9401);
or U9613 (N_9613,N_9491,N_9562);
or U9614 (N_9614,N_9519,N_9548);
nand U9615 (N_9615,N_9420,N_9451);
nand U9616 (N_9616,N_9422,N_9525);
nand U9617 (N_9617,N_9591,N_9441);
and U9618 (N_9618,N_9510,N_9426);
nor U9619 (N_9619,N_9482,N_9458);
nand U9620 (N_9620,N_9581,N_9481);
nand U9621 (N_9621,N_9433,N_9571);
nor U9622 (N_9622,N_9557,N_9552);
nand U9623 (N_9623,N_9414,N_9566);
xor U9624 (N_9624,N_9415,N_9430);
nand U9625 (N_9625,N_9461,N_9416);
xor U9626 (N_9626,N_9560,N_9572);
xnor U9627 (N_9627,N_9568,N_9595);
and U9628 (N_9628,N_9544,N_9493);
and U9629 (N_9629,N_9538,N_9501);
or U9630 (N_9630,N_9529,N_9584);
and U9631 (N_9631,N_9513,N_9489);
nand U9632 (N_9632,N_9593,N_9406);
xor U9633 (N_9633,N_9569,N_9575);
xnor U9634 (N_9634,N_9476,N_9556);
and U9635 (N_9635,N_9537,N_9509);
nor U9636 (N_9636,N_9446,N_9549);
or U9637 (N_9637,N_9452,N_9521);
nor U9638 (N_9638,N_9536,N_9553);
or U9639 (N_9639,N_9424,N_9515);
nor U9640 (N_9640,N_9455,N_9596);
xnor U9641 (N_9641,N_9504,N_9425);
or U9642 (N_9642,N_9474,N_9408);
and U9643 (N_9643,N_9547,N_9577);
and U9644 (N_9644,N_9419,N_9518);
and U9645 (N_9645,N_9508,N_9467);
nand U9646 (N_9646,N_9540,N_9402);
nand U9647 (N_9647,N_9417,N_9484);
nor U9648 (N_9648,N_9503,N_9559);
nand U9649 (N_9649,N_9405,N_9460);
nor U9650 (N_9650,N_9541,N_9495);
nor U9651 (N_9651,N_9492,N_9439);
xor U9652 (N_9652,N_9479,N_9459);
nor U9653 (N_9653,N_9478,N_9599);
nor U9654 (N_9654,N_9431,N_9486);
xnor U9655 (N_9655,N_9507,N_9555);
nand U9656 (N_9656,N_9527,N_9502);
nor U9657 (N_9657,N_9469,N_9454);
nand U9658 (N_9658,N_9444,N_9570);
nor U9659 (N_9659,N_9533,N_9477);
or U9660 (N_9660,N_9561,N_9465);
xor U9661 (N_9661,N_9472,N_9563);
xor U9662 (N_9662,N_9450,N_9443);
xor U9663 (N_9663,N_9594,N_9574);
nor U9664 (N_9664,N_9400,N_9497);
xnor U9665 (N_9665,N_9580,N_9597);
nor U9666 (N_9666,N_9442,N_9558);
and U9667 (N_9667,N_9598,N_9573);
nor U9668 (N_9668,N_9411,N_9466);
and U9669 (N_9669,N_9534,N_9542);
nor U9670 (N_9670,N_9506,N_9531);
or U9671 (N_9671,N_9480,N_9520);
or U9672 (N_9672,N_9423,N_9522);
and U9673 (N_9673,N_9407,N_9412);
and U9674 (N_9674,N_9530,N_9588);
nor U9675 (N_9675,N_9579,N_9592);
or U9676 (N_9676,N_9554,N_9449);
nor U9677 (N_9677,N_9410,N_9435);
xnor U9678 (N_9678,N_9565,N_9500);
nand U9679 (N_9679,N_9428,N_9512);
and U9680 (N_9680,N_9437,N_9409);
nand U9681 (N_9681,N_9494,N_9445);
nor U9682 (N_9682,N_9528,N_9462);
xor U9683 (N_9683,N_9545,N_9463);
and U9684 (N_9684,N_9403,N_9590);
nor U9685 (N_9685,N_9535,N_9448);
and U9686 (N_9686,N_9427,N_9576);
or U9687 (N_9687,N_9526,N_9440);
xnor U9688 (N_9688,N_9471,N_9550);
nand U9689 (N_9689,N_9434,N_9432);
xor U9690 (N_9690,N_9587,N_9582);
nand U9691 (N_9691,N_9475,N_9511);
and U9692 (N_9692,N_9524,N_9447);
xor U9693 (N_9693,N_9586,N_9487);
nand U9694 (N_9694,N_9578,N_9436);
nand U9695 (N_9695,N_9516,N_9505);
nor U9696 (N_9696,N_9567,N_9438);
or U9697 (N_9697,N_9468,N_9413);
nor U9698 (N_9698,N_9488,N_9429);
and U9699 (N_9699,N_9457,N_9532);
xnor U9700 (N_9700,N_9561,N_9482);
and U9701 (N_9701,N_9455,N_9519);
or U9702 (N_9702,N_9414,N_9564);
and U9703 (N_9703,N_9545,N_9520);
and U9704 (N_9704,N_9597,N_9502);
nor U9705 (N_9705,N_9484,N_9532);
nor U9706 (N_9706,N_9511,N_9591);
or U9707 (N_9707,N_9408,N_9428);
or U9708 (N_9708,N_9522,N_9407);
nor U9709 (N_9709,N_9423,N_9537);
and U9710 (N_9710,N_9500,N_9551);
xor U9711 (N_9711,N_9439,N_9406);
nor U9712 (N_9712,N_9431,N_9446);
nand U9713 (N_9713,N_9531,N_9429);
nand U9714 (N_9714,N_9484,N_9502);
nand U9715 (N_9715,N_9435,N_9549);
or U9716 (N_9716,N_9426,N_9516);
nor U9717 (N_9717,N_9576,N_9505);
nor U9718 (N_9718,N_9400,N_9583);
or U9719 (N_9719,N_9590,N_9541);
nor U9720 (N_9720,N_9410,N_9429);
nand U9721 (N_9721,N_9503,N_9441);
or U9722 (N_9722,N_9467,N_9559);
nor U9723 (N_9723,N_9494,N_9565);
nand U9724 (N_9724,N_9407,N_9503);
or U9725 (N_9725,N_9591,N_9504);
or U9726 (N_9726,N_9407,N_9560);
nand U9727 (N_9727,N_9592,N_9513);
and U9728 (N_9728,N_9507,N_9426);
and U9729 (N_9729,N_9448,N_9464);
or U9730 (N_9730,N_9505,N_9453);
nor U9731 (N_9731,N_9533,N_9524);
nor U9732 (N_9732,N_9443,N_9558);
or U9733 (N_9733,N_9564,N_9402);
and U9734 (N_9734,N_9439,N_9579);
nand U9735 (N_9735,N_9583,N_9464);
nor U9736 (N_9736,N_9463,N_9487);
or U9737 (N_9737,N_9402,N_9439);
nor U9738 (N_9738,N_9446,N_9567);
nand U9739 (N_9739,N_9404,N_9546);
or U9740 (N_9740,N_9527,N_9532);
and U9741 (N_9741,N_9464,N_9580);
and U9742 (N_9742,N_9429,N_9548);
nor U9743 (N_9743,N_9422,N_9483);
nand U9744 (N_9744,N_9462,N_9435);
and U9745 (N_9745,N_9483,N_9475);
nand U9746 (N_9746,N_9458,N_9490);
or U9747 (N_9747,N_9598,N_9510);
or U9748 (N_9748,N_9578,N_9489);
xnor U9749 (N_9749,N_9430,N_9420);
nor U9750 (N_9750,N_9598,N_9492);
and U9751 (N_9751,N_9404,N_9519);
nor U9752 (N_9752,N_9416,N_9503);
nand U9753 (N_9753,N_9565,N_9490);
nor U9754 (N_9754,N_9457,N_9515);
and U9755 (N_9755,N_9466,N_9459);
nand U9756 (N_9756,N_9562,N_9448);
nor U9757 (N_9757,N_9582,N_9426);
or U9758 (N_9758,N_9568,N_9575);
and U9759 (N_9759,N_9576,N_9483);
nand U9760 (N_9760,N_9492,N_9588);
nand U9761 (N_9761,N_9411,N_9567);
and U9762 (N_9762,N_9573,N_9507);
and U9763 (N_9763,N_9584,N_9449);
nand U9764 (N_9764,N_9443,N_9464);
or U9765 (N_9765,N_9568,N_9403);
nor U9766 (N_9766,N_9511,N_9513);
xnor U9767 (N_9767,N_9467,N_9434);
nor U9768 (N_9768,N_9533,N_9467);
xor U9769 (N_9769,N_9407,N_9411);
or U9770 (N_9770,N_9525,N_9428);
nand U9771 (N_9771,N_9560,N_9565);
nor U9772 (N_9772,N_9482,N_9497);
nor U9773 (N_9773,N_9522,N_9498);
nor U9774 (N_9774,N_9540,N_9537);
or U9775 (N_9775,N_9483,N_9457);
and U9776 (N_9776,N_9424,N_9540);
xnor U9777 (N_9777,N_9434,N_9446);
xor U9778 (N_9778,N_9422,N_9556);
and U9779 (N_9779,N_9574,N_9443);
and U9780 (N_9780,N_9434,N_9547);
or U9781 (N_9781,N_9515,N_9489);
nand U9782 (N_9782,N_9585,N_9487);
or U9783 (N_9783,N_9491,N_9434);
and U9784 (N_9784,N_9492,N_9411);
nor U9785 (N_9785,N_9513,N_9468);
nand U9786 (N_9786,N_9461,N_9563);
nor U9787 (N_9787,N_9487,N_9424);
xnor U9788 (N_9788,N_9580,N_9491);
nand U9789 (N_9789,N_9518,N_9421);
or U9790 (N_9790,N_9599,N_9400);
or U9791 (N_9791,N_9442,N_9542);
or U9792 (N_9792,N_9553,N_9452);
xnor U9793 (N_9793,N_9541,N_9499);
or U9794 (N_9794,N_9540,N_9588);
xor U9795 (N_9795,N_9403,N_9431);
xnor U9796 (N_9796,N_9468,N_9444);
nand U9797 (N_9797,N_9565,N_9457);
nand U9798 (N_9798,N_9430,N_9469);
xnor U9799 (N_9799,N_9568,N_9505);
and U9800 (N_9800,N_9685,N_9607);
or U9801 (N_9801,N_9657,N_9698);
nor U9802 (N_9802,N_9750,N_9771);
xnor U9803 (N_9803,N_9742,N_9712);
or U9804 (N_9804,N_9702,N_9673);
nand U9805 (N_9805,N_9717,N_9730);
nand U9806 (N_9806,N_9656,N_9744);
or U9807 (N_9807,N_9679,N_9608);
xor U9808 (N_9808,N_9682,N_9731);
or U9809 (N_9809,N_9670,N_9738);
and U9810 (N_9810,N_9691,N_9667);
and U9811 (N_9811,N_9622,N_9718);
nand U9812 (N_9812,N_9641,N_9797);
nor U9813 (N_9813,N_9737,N_9677);
xnor U9814 (N_9814,N_9701,N_9736);
nor U9815 (N_9815,N_9780,N_9711);
and U9816 (N_9816,N_9752,N_9774);
and U9817 (N_9817,N_9707,N_9620);
and U9818 (N_9818,N_9621,N_9669);
nand U9819 (N_9819,N_9633,N_9770);
nand U9820 (N_9820,N_9781,N_9766);
or U9821 (N_9821,N_9617,N_9626);
nand U9822 (N_9822,N_9634,N_9693);
or U9823 (N_9823,N_9603,N_9666);
or U9824 (N_9824,N_9757,N_9725);
nor U9825 (N_9825,N_9755,N_9606);
nand U9826 (N_9826,N_9709,N_9715);
nor U9827 (N_9827,N_9678,N_9688);
nor U9828 (N_9828,N_9788,N_9743);
and U9829 (N_9829,N_9655,N_9729);
nor U9830 (N_9830,N_9787,N_9630);
xor U9831 (N_9831,N_9751,N_9605);
nor U9832 (N_9832,N_9661,N_9675);
and U9833 (N_9833,N_9694,N_9676);
nand U9834 (N_9834,N_9662,N_9650);
and U9835 (N_9835,N_9628,N_9643);
and U9836 (N_9836,N_9705,N_9660);
xor U9837 (N_9837,N_9710,N_9625);
or U9838 (N_9838,N_9689,N_9719);
nand U9839 (N_9839,N_9779,N_9721);
and U9840 (N_9840,N_9767,N_9658);
or U9841 (N_9841,N_9627,N_9776);
or U9842 (N_9842,N_9614,N_9668);
and U9843 (N_9843,N_9623,N_9600);
and U9844 (N_9844,N_9611,N_9749);
xor U9845 (N_9845,N_9637,N_9758);
xor U9846 (N_9846,N_9704,N_9601);
and U9847 (N_9847,N_9610,N_9624);
nand U9848 (N_9848,N_9665,N_9681);
and U9849 (N_9849,N_9723,N_9773);
nor U9850 (N_9850,N_9746,N_9671);
and U9851 (N_9851,N_9713,N_9648);
xor U9852 (N_9852,N_9785,N_9636);
or U9853 (N_9853,N_9680,N_9708);
and U9854 (N_9854,N_9684,N_9647);
and U9855 (N_9855,N_9615,N_9799);
xor U9856 (N_9856,N_9720,N_9649);
nand U9857 (N_9857,N_9745,N_9638);
nand U9858 (N_9858,N_9795,N_9756);
xnor U9859 (N_9859,N_9672,N_9703);
xnor U9860 (N_9860,N_9659,N_9697);
and U9861 (N_9861,N_9619,N_9798);
and U9862 (N_9862,N_9635,N_9753);
xor U9863 (N_9863,N_9748,N_9663);
or U9864 (N_9864,N_9612,N_9653);
and U9865 (N_9865,N_9613,N_9645);
xor U9866 (N_9866,N_9768,N_9646);
nand U9867 (N_9867,N_9765,N_9741);
or U9868 (N_9868,N_9686,N_9792);
nor U9869 (N_9869,N_9772,N_9726);
or U9870 (N_9870,N_9674,N_9734);
xnor U9871 (N_9871,N_9696,N_9714);
and U9872 (N_9872,N_9747,N_9692);
nand U9873 (N_9873,N_9754,N_9644);
nand U9874 (N_9874,N_9790,N_9740);
xnor U9875 (N_9875,N_9796,N_9727);
nand U9876 (N_9876,N_9616,N_9735);
nand U9877 (N_9877,N_9664,N_9789);
or U9878 (N_9878,N_9739,N_9654);
xor U9879 (N_9879,N_9690,N_9777);
or U9880 (N_9880,N_9602,N_9761);
nand U9881 (N_9881,N_9760,N_9778);
or U9882 (N_9882,N_9782,N_9722);
and U9883 (N_9883,N_9683,N_9706);
xor U9884 (N_9884,N_9762,N_9716);
nand U9885 (N_9885,N_9639,N_9631);
xor U9886 (N_9886,N_9769,N_9764);
or U9887 (N_9887,N_9687,N_9786);
nor U9888 (N_9888,N_9699,N_9724);
xor U9889 (N_9889,N_9695,N_9618);
or U9890 (N_9890,N_9640,N_9759);
and U9891 (N_9891,N_9651,N_9793);
nand U9892 (N_9892,N_9763,N_9604);
or U9893 (N_9893,N_9652,N_9700);
or U9894 (N_9894,N_9728,N_9794);
nand U9895 (N_9895,N_9791,N_9733);
xnor U9896 (N_9896,N_9609,N_9784);
and U9897 (N_9897,N_9642,N_9629);
or U9898 (N_9898,N_9732,N_9775);
nor U9899 (N_9899,N_9632,N_9783);
and U9900 (N_9900,N_9661,N_9667);
xor U9901 (N_9901,N_9618,N_9772);
or U9902 (N_9902,N_9627,N_9680);
xnor U9903 (N_9903,N_9784,N_9737);
nor U9904 (N_9904,N_9625,N_9682);
nand U9905 (N_9905,N_9779,N_9742);
or U9906 (N_9906,N_9721,N_9663);
and U9907 (N_9907,N_9740,N_9686);
nor U9908 (N_9908,N_9641,N_9648);
or U9909 (N_9909,N_9718,N_9785);
xnor U9910 (N_9910,N_9765,N_9777);
and U9911 (N_9911,N_9637,N_9697);
or U9912 (N_9912,N_9755,N_9604);
xor U9913 (N_9913,N_9794,N_9784);
nor U9914 (N_9914,N_9722,N_9740);
and U9915 (N_9915,N_9716,N_9793);
and U9916 (N_9916,N_9643,N_9794);
nor U9917 (N_9917,N_9738,N_9677);
xnor U9918 (N_9918,N_9632,N_9633);
or U9919 (N_9919,N_9735,N_9628);
xor U9920 (N_9920,N_9770,N_9636);
xnor U9921 (N_9921,N_9723,N_9744);
nor U9922 (N_9922,N_9713,N_9631);
nor U9923 (N_9923,N_9630,N_9799);
nand U9924 (N_9924,N_9641,N_9656);
nor U9925 (N_9925,N_9665,N_9790);
nand U9926 (N_9926,N_9796,N_9672);
nand U9927 (N_9927,N_9630,N_9750);
xor U9928 (N_9928,N_9669,N_9604);
nand U9929 (N_9929,N_9661,N_9666);
or U9930 (N_9930,N_9635,N_9733);
or U9931 (N_9931,N_9725,N_9720);
xnor U9932 (N_9932,N_9798,N_9738);
and U9933 (N_9933,N_9605,N_9657);
or U9934 (N_9934,N_9697,N_9738);
and U9935 (N_9935,N_9641,N_9713);
or U9936 (N_9936,N_9718,N_9736);
nand U9937 (N_9937,N_9622,N_9663);
or U9938 (N_9938,N_9664,N_9682);
and U9939 (N_9939,N_9769,N_9729);
nand U9940 (N_9940,N_9694,N_9636);
or U9941 (N_9941,N_9707,N_9630);
or U9942 (N_9942,N_9688,N_9789);
nor U9943 (N_9943,N_9757,N_9708);
or U9944 (N_9944,N_9679,N_9751);
and U9945 (N_9945,N_9638,N_9760);
nand U9946 (N_9946,N_9642,N_9653);
nand U9947 (N_9947,N_9751,N_9609);
nand U9948 (N_9948,N_9640,N_9762);
nand U9949 (N_9949,N_9725,N_9706);
or U9950 (N_9950,N_9792,N_9756);
or U9951 (N_9951,N_9644,N_9649);
xor U9952 (N_9952,N_9795,N_9668);
and U9953 (N_9953,N_9673,N_9674);
or U9954 (N_9954,N_9630,N_9727);
nand U9955 (N_9955,N_9682,N_9712);
and U9956 (N_9956,N_9604,N_9713);
xor U9957 (N_9957,N_9671,N_9766);
or U9958 (N_9958,N_9740,N_9656);
nor U9959 (N_9959,N_9604,N_9688);
nor U9960 (N_9960,N_9673,N_9636);
nand U9961 (N_9961,N_9770,N_9653);
or U9962 (N_9962,N_9672,N_9755);
and U9963 (N_9963,N_9747,N_9657);
nand U9964 (N_9964,N_9713,N_9697);
nand U9965 (N_9965,N_9672,N_9630);
or U9966 (N_9966,N_9745,N_9615);
nor U9967 (N_9967,N_9623,N_9609);
and U9968 (N_9968,N_9617,N_9675);
nor U9969 (N_9969,N_9775,N_9671);
or U9970 (N_9970,N_9785,N_9717);
nand U9971 (N_9971,N_9769,N_9689);
nand U9972 (N_9972,N_9734,N_9788);
nand U9973 (N_9973,N_9664,N_9646);
nor U9974 (N_9974,N_9690,N_9786);
or U9975 (N_9975,N_9633,N_9700);
nor U9976 (N_9976,N_9716,N_9711);
nand U9977 (N_9977,N_9772,N_9754);
xor U9978 (N_9978,N_9653,N_9646);
xor U9979 (N_9979,N_9745,N_9735);
or U9980 (N_9980,N_9728,N_9634);
xnor U9981 (N_9981,N_9638,N_9787);
and U9982 (N_9982,N_9770,N_9698);
nor U9983 (N_9983,N_9792,N_9720);
nor U9984 (N_9984,N_9665,N_9743);
nor U9985 (N_9985,N_9735,N_9718);
and U9986 (N_9986,N_9786,N_9755);
xnor U9987 (N_9987,N_9692,N_9672);
and U9988 (N_9988,N_9662,N_9723);
or U9989 (N_9989,N_9704,N_9620);
xnor U9990 (N_9990,N_9699,N_9669);
or U9991 (N_9991,N_9750,N_9623);
or U9992 (N_9992,N_9712,N_9640);
and U9993 (N_9993,N_9784,N_9626);
xor U9994 (N_9994,N_9748,N_9747);
nor U9995 (N_9995,N_9780,N_9736);
xnor U9996 (N_9996,N_9778,N_9639);
nor U9997 (N_9997,N_9778,N_9789);
and U9998 (N_9998,N_9632,N_9750);
xnor U9999 (N_9999,N_9791,N_9701);
nand U10000 (N_10000,N_9924,N_9999);
and U10001 (N_10001,N_9816,N_9946);
nor U10002 (N_10002,N_9883,N_9819);
and U10003 (N_10003,N_9885,N_9833);
and U10004 (N_10004,N_9986,N_9987);
nor U10005 (N_10005,N_9855,N_9815);
and U10006 (N_10006,N_9968,N_9954);
xnor U10007 (N_10007,N_9820,N_9847);
nand U10008 (N_10008,N_9837,N_9950);
nand U10009 (N_10009,N_9982,N_9806);
nor U10010 (N_10010,N_9923,N_9817);
and U10011 (N_10011,N_9912,N_9908);
nor U10012 (N_10012,N_9869,N_9934);
nand U10013 (N_10013,N_9842,N_9905);
nand U10014 (N_10014,N_9917,N_9927);
or U10015 (N_10015,N_9832,N_9872);
xor U10016 (N_10016,N_9991,N_9861);
or U10017 (N_10017,N_9825,N_9959);
nor U10018 (N_10018,N_9926,N_9802);
nor U10019 (N_10019,N_9893,N_9848);
or U10020 (N_10020,N_9904,N_9996);
xnor U10021 (N_10021,N_9836,N_9914);
nand U10022 (N_10022,N_9894,N_9887);
nor U10023 (N_10023,N_9877,N_9918);
nor U10024 (N_10024,N_9862,N_9897);
nor U10025 (N_10025,N_9916,N_9945);
and U10026 (N_10026,N_9811,N_9866);
and U10027 (N_10027,N_9983,N_9822);
nand U10028 (N_10028,N_9834,N_9853);
nor U10029 (N_10029,N_9818,N_9981);
xnor U10030 (N_10030,N_9947,N_9903);
nor U10031 (N_10031,N_9890,N_9948);
xor U10032 (N_10032,N_9997,N_9845);
nor U10033 (N_10033,N_9857,N_9984);
xor U10034 (N_10034,N_9972,N_9846);
nand U10035 (N_10035,N_9814,N_9973);
xnor U10036 (N_10036,N_9960,N_9949);
xor U10037 (N_10037,N_9863,N_9901);
nand U10038 (N_10038,N_9868,N_9852);
and U10039 (N_10039,N_9804,N_9921);
or U10040 (N_10040,N_9849,N_9951);
or U10041 (N_10041,N_9995,N_9907);
and U10042 (N_10042,N_9958,N_9952);
nor U10043 (N_10043,N_9879,N_9882);
xnor U10044 (N_10044,N_9956,N_9993);
nor U10045 (N_10045,N_9933,N_9838);
and U10046 (N_10046,N_9876,N_9895);
nor U10047 (N_10047,N_9910,N_9967);
nand U10048 (N_10048,N_9911,N_9902);
and U10049 (N_10049,N_9940,N_9977);
and U10050 (N_10050,N_9936,N_9841);
nand U10051 (N_10051,N_9859,N_9888);
or U10052 (N_10052,N_9909,N_9827);
or U10053 (N_10053,N_9939,N_9844);
nand U10054 (N_10054,N_9942,N_9929);
and U10055 (N_10055,N_9928,N_9919);
and U10056 (N_10056,N_9899,N_9970);
nor U10057 (N_10057,N_9943,N_9864);
nand U10058 (N_10058,N_9807,N_9990);
and U10059 (N_10059,N_9920,N_9880);
and U10060 (N_10060,N_9922,N_9898);
xor U10061 (N_10061,N_9856,N_9944);
nand U10062 (N_10062,N_9961,N_9965);
nor U10063 (N_10063,N_9808,N_9858);
xor U10064 (N_10064,N_9830,N_9932);
or U10065 (N_10065,N_9874,N_9854);
nor U10066 (N_10066,N_9821,N_9812);
xnor U10067 (N_10067,N_9935,N_9925);
nand U10068 (N_10068,N_9957,N_9813);
and U10069 (N_10069,N_9875,N_9892);
nand U10070 (N_10070,N_9826,N_9955);
nor U10071 (N_10071,N_9809,N_9803);
and U10072 (N_10072,N_9913,N_9979);
nor U10073 (N_10073,N_9801,N_9966);
xor U10074 (N_10074,N_9931,N_9896);
nor U10075 (N_10075,N_9978,N_9805);
nand U10076 (N_10076,N_9938,N_9871);
nor U10077 (N_10077,N_9891,N_9998);
nor U10078 (N_10078,N_9840,N_9953);
xor U10079 (N_10079,N_9975,N_9930);
and U10080 (N_10080,N_9976,N_9870);
xnor U10081 (N_10081,N_9989,N_9937);
nand U10082 (N_10082,N_9873,N_9980);
and U10083 (N_10083,N_9831,N_9985);
or U10084 (N_10084,N_9851,N_9867);
and U10085 (N_10085,N_9941,N_9974);
and U10086 (N_10086,N_9850,N_9878);
or U10087 (N_10087,N_9889,N_9824);
and U10088 (N_10088,N_9828,N_9962);
nand U10089 (N_10089,N_9963,N_9865);
or U10090 (N_10090,N_9988,N_9915);
and U10091 (N_10091,N_9800,N_9992);
nor U10092 (N_10092,N_9964,N_9994);
or U10093 (N_10093,N_9971,N_9969);
and U10094 (N_10094,N_9839,N_9900);
or U10095 (N_10095,N_9829,N_9835);
nor U10096 (N_10096,N_9823,N_9884);
nor U10097 (N_10097,N_9881,N_9860);
nor U10098 (N_10098,N_9886,N_9810);
and U10099 (N_10099,N_9906,N_9843);
nor U10100 (N_10100,N_9926,N_9877);
and U10101 (N_10101,N_9871,N_9852);
nand U10102 (N_10102,N_9901,N_9927);
or U10103 (N_10103,N_9984,N_9947);
or U10104 (N_10104,N_9972,N_9944);
nor U10105 (N_10105,N_9988,N_9910);
nand U10106 (N_10106,N_9989,N_9837);
or U10107 (N_10107,N_9921,N_9838);
or U10108 (N_10108,N_9844,N_9971);
or U10109 (N_10109,N_9984,N_9963);
nand U10110 (N_10110,N_9917,N_9851);
and U10111 (N_10111,N_9864,N_9880);
and U10112 (N_10112,N_9967,N_9873);
or U10113 (N_10113,N_9850,N_9993);
xor U10114 (N_10114,N_9909,N_9857);
or U10115 (N_10115,N_9928,N_9909);
and U10116 (N_10116,N_9959,N_9818);
nor U10117 (N_10117,N_9809,N_9829);
nand U10118 (N_10118,N_9849,N_9831);
and U10119 (N_10119,N_9819,N_9802);
or U10120 (N_10120,N_9844,N_9860);
or U10121 (N_10121,N_9804,N_9991);
or U10122 (N_10122,N_9951,N_9924);
and U10123 (N_10123,N_9973,N_9872);
nor U10124 (N_10124,N_9867,N_9949);
or U10125 (N_10125,N_9976,N_9955);
nand U10126 (N_10126,N_9899,N_9879);
and U10127 (N_10127,N_9845,N_9867);
xor U10128 (N_10128,N_9821,N_9878);
nand U10129 (N_10129,N_9823,N_9818);
xnor U10130 (N_10130,N_9860,N_9912);
xor U10131 (N_10131,N_9862,N_9858);
nand U10132 (N_10132,N_9888,N_9897);
and U10133 (N_10133,N_9819,N_9971);
or U10134 (N_10134,N_9917,N_9913);
xnor U10135 (N_10135,N_9850,N_9989);
or U10136 (N_10136,N_9842,N_9976);
or U10137 (N_10137,N_9819,N_9892);
xor U10138 (N_10138,N_9887,N_9913);
nor U10139 (N_10139,N_9883,N_9905);
xnor U10140 (N_10140,N_9805,N_9887);
nor U10141 (N_10141,N_9808,N_9978);
and U10142 (N_10142,N_9955,N_9862);
xor U10143 (N_10143,N_9859,N_9948);
and U10144 (N_10144,N_9800,N_9844);
xnor U10145 (N_10145,N_9945,N_9851);
nor U10146 (N_10146,N_9880,N_9834);
or U10147 (N_10147,N_9891,N_9833);
nand U10148 (N_10148,N_9825,N_9830);
nor U10149 (N_10149,N_9919,N_9805);
or U10150 (N_10150,N_9928,N_9984);
xor U10151 (N_10151,N_9848,N_9965);
xor U10152 (N_10152,N_9975,N_9814);
nand U10153 (N_10153,N_9898,N_9991);
and U10154 (N_10154,N_9978,N_9919);
nor U10155 (N_10155,N_9992,N_9872);
xnor U10156 (N_10156,N_9923,N_9986);
nor U10157 (N_10157,N_9973,N_9868);
xor U10158 (N_10158,N_9933,N_9996);
nand U10159 (N_10159,N_9928,N_9904);
nor U10160 (N_10160,N_9910,N_9947);
xnor U10161 (N_10161,N_9910,N_9877);
nor U10162 (N_10162,N_9827,N_9801);
nor U10163 (N_10163,N_9923,N_9871);
nand U10164 (N_10164,N_9911,N_9968);
or U10165 (N_10165,N_9984,N_9983);
nor U10166 (N_10166,N_9836,N_9900);
or U10167 (N_10167,N_9889,N_9990);
nor U10168 (N_10168,N_9897,N_9943);
nor U10169 (N_10169,N_9895,N_9981);
xnor U10170 (N_10170,N_9849,N_9846);
nand U10171 (N_10171,N_9893,N_9891);
xor U10172 (N_10172,N_9980,N_9951);
nor U10173 (N_10173,N_9827,N_9950);
nand U10174 (N_10174,N_9957,N_9846);
nand U10175 (N_10175,N_9893,N_9975);
xnor U10176 (N_10176,N_9858,N_9932);
and U10177 (N_10177,N_9936,N_9917);
nor U10178 (N_10178,N_9931,N_9813);
or U10179 (N_10179,N_9889,N_9986);
xnor U10180 (N_10180,N_9973,N_9952);
nand U10181 (N_10181,N_9999,N_9984);
nor U10182 (N_10182,N_9855,N_9870);
nor U10183 (N_10183,N_9991,N_9893);
xor U10184 (N_10184,N_9870,N_9858);
xnor U10185 (N_10185,N_9975,N_9922);
nand U10186 (N_10186,N_9851,N_9919);
or U10187 (N_10187,N_9930,N_9833);
or U10188 (N_10188,N_9802,N_9925);
nor U10189 (N_10189,N_9989,N_9928);
or U10190 (N_10190,N_9834,N_9881);
nor U10191 (N_10191,N_9858,N_9949);
and U10192 (N_10192,N_9804,N_9835);
nor U10193 (N_10193,N_9925,N_9954);
and U10194 (N_10194,N_9890,N_9850);
or U10195 (N_10195,N_9802,N_9948);
xnor U10196 (N_10196,N_9964,N_9960);
nand U10197 (N_10197,N_9935,N_9951);
xor U10198 (N_10198,N_9934,N_9888);
nor U10199 (N_10199,N_9872,N_9962);
nor U10200 (N_10200,N_10005,N_10121);
and U10201 (N_10201,N_10001,N_10190);
and U10202 (N_10202,N_10100,N_10152);
or U10203 (N_10203,N_10108,N_10097);
xor U10204 (N_10204,N_10168,N_10133);
nor U10205 (N_10205,N_10075,N_10081);
xor U10206 (N_10206,N_10076,N_10086);
nor U10207 (N_10207,N_10025,N_10048);
and U10208 (N_10208,N_10023,N_10056);
or U10209 (N_10209,N_10116,N_10194);
and U10210 (N_10210,N_10020,N_10182);
nor U10211 (N_10211,N_10157,N_10069);
xnor U10212 (N_10212,N_10027,N_10186);
nor U10213 (N_10213,N_10191,N_10178);
nand U10214 (N_10214,N_10037,N_10145);
or U10215 (N_10215,N_10154,N_10163);
or U10216 (N_10216,N_10144,N_10196);
xor U10217 (N_10217,N_10162,N_10006);
xor U10218 (N_10218,N_10080,N_10012);
xor U10219 (N_10219,N_10046,N_10039);
or U10220 (N_10220,N_10102,N_10147);
or U10221 (N_10221,N_10013,N_10011);
or U10222 (N_10222,N_10174,N_10058);
nor U10223 (N_10223,N_10130,N_10140);
and U10224 (N_10224,N_10197,N_10078);
nor U10225 (N_10225,N_10195,N_10067);
nand U10226 (N_10226,N_10091,N_10101);
and U10227 (N_10227,N_10126,N_10095);
nand U10228 (N_10228,N_10018,N_10089);
nor U10229 (N_10229,N_10170,N_10019);
xor U10230 (N_10230,N_10028,N_10139);
and U10231 (N_10231,N_10034,N_10060);
nand U10232 (N_10232,N_10110,N_10193);
and U10233 (N_10233,N_10038,N_10159);
or U10234 (N_10234,N_10175,N_10050);
nor U10235 (N_10235,N_10141,N_10169);
or U10236 (N_10236,N_10151,N_10082);
nor U10237 (N_10237,N_10107,N_10138);
or U10238 (N_10238,N_10061,N_10087);
xnor U10239 (N_10239,N_10041,N_10047);
nand U10240 (N_10240,N_10043,N_10088);
nand U10241 (N_10241,N_10149,N_10040);
nor U10242 (N_10242,N_10137,N_10142);
nand U10243 (N_10243,N_10109,N_10068);
or U10244 (N_10244,N_10183,N_10134);
and U10245 (N_10245,N_10181,N_10003);
xor U10246 (N_10246,N_10032,N_10042);
nor U10247 (N_10247,N_10125,N_10187);
or U10248 (N_10248,N_10172,N_10055);
nor U10249 (N_10249,N_10029,N_10092);
and U10250 (N_10250,N_10173,N_10179);
nor U10251 (N_10251,N_10131,N_10167);
nand U10252 (N_10252,N_10099,N_10198);
nor U10253 (N_10253,N_10132,N_10017);
nor U10254 (N_10254,N_10084,N_10079);
or U10255 (N_10255,N_10009,N_10007);
xor U10256 (N_10256,N_10014,N_10111);
or U10257 (N_10257,N_10171,N_10010);
nand U10258 (N_10258,N_10002,N_10104);
nand U10259 (N_10259,N_10189,N_10185);
or U10260 (N_10260,N_10093,N_10030);
or U10261 (N_10261,N_10035,N_10136);
xnor U10262 (N_10262,N_10052,N_10074);
nor U10263 (N_10263,N_10192,N_10083);
nand U10264 (N_10264,N_10156,N_10016);
or U10265 (N_10265,N_10122,N_10053);
xnor U10266 (N_10266,N_10004,N_10066);
xor U10267 (N_10267,N_10085,N_10064);
nor U10268 (N_10268,N_10153,N_10062);
and U10269 (N_10269,N_10073,N_10022);
nor U10270 (N_10270,N_10127,N_10160);
nand U10271 (N_10271,N_10094,N_10033);
xnor U10272 (N_10272,N_10150,N_10148);
and U10273 (N_10273,N_10177,N_10158);
and U10274 (N_10274,N_10184,N_10051);
or U10275 (N_10275,N_10106,N_10114);
and U10276 (N_10276,N_10124,N_10072);
and U10277 (N_10277,N_10115,N_10077);
xor U10278 (N_10278,N_10065,N_10026);
or U10279 (N_10279,N_10117,N_10054);
xor U10280 (N_10280,N_10090,N_10164);
xnor U10281 (N_10281,N_10118,N_10036);
or U10282 (N_10282,N_10188,N_10063);
nor U10283 (N_10283,N_10113,N_10103);
nand U10284 (N_10284,N_10180,N_10143);
nor U10285 (N_10285,N_10199,N_10057);
or U10286 (N_10286,N_10021,N_10123);
or U10287 (N_10287,N_10112,N_10015);
nand U10288 (N_10288,N_10024,N_10161);
or U10289 (N_10289,N_10146,N_10059);
nor U10290 (N_10290,N_10008,N_10176);
nand U10291 (N_10291,N_10044,N_10000);
or U10292 (N_10292,N_10135,N_10166);
nor U10293 (N_10293,N_10128,N_10105);
or U10294 (N_10294,N_10098,N_10165);
and U10295 (N_10295,N_10119,N_10096);
xnor U10296 (N_10296,N_10070,N_10120);
or U10297 (N_10297,N_10129,N_10071);
nor U10298 (N_10298,N_10045,N_10049);
xor U10299 (N_10299,N_10031,N_10155);
or U10300 (N_10300,N_10078,N_10000);
nand U10301 (N_10301,N_10159,N_10046);
and U10302 (N_10302,N_10113,N_10017);
xor U10303 (N_10303,N_10111,N_10026);
and U10304 (N_10304,N_10194,N_10123);
nor U10305 (N_10305,N_10113,N_10063);
or U10306 (N_10306,N_10138,N_10031);
or U10307 (N_10307,N_10181,N_10019);
and U10308 (N_10308,N_10054,N_10180);
nand U10309 (N_10309,N_10195,N_10091);
and U10310 (N_10310,N_10017,N_10129);
or U10311 (N_10311,N_10083,N_10098);
nor U10312 (N_10312,N_10193,N_10145);
or U10313 (N_10313,N_10002,N_10042);
or U10314 (N_10314,N_10022,N_10131);
or U10315 (N_10315,N_10174,N_10094);
xor U10316 (N_10316,N_10090,N_10106);
or U10317 (N_10317,N_10031,N_10157);
and U10318 (N_10318,N_10135,N_10005);
or U10319 (N_10319,N_10160,N_10196);
xnor U10320 (N_10320,N_10160,N_10157);
xor U10321 (N_10321,N_10009,N_10004);
or U10322 (N_10322,N_10059,N_10120);
or U10323 (N_10323,N_10196,N_10190);
and U10324 (N_10324,N_10015,N_10152);
and U10325 (N_10325,N_10102,N_10185);
nand U10326 (N_10326,N_10078,N_10128);
nand U10327 (N_10327,N_10062,N_10061);
and U10328 (N_10328,N_10143,N_10017);
or U10329 (N_10329,N_10147,N_10148);
and U10330 (N_10330,N_10181,N_10049);
nand U10331 (N_10331,N_10126,N_10022);
or U10332 (N_10332,N_10061,N_10112);
nor U10333 (N_10333,N_10008,N_10003);
nand U10334 (N_10334,N_10058,N_10035);
and U10335 (N_10335,N_10066,N_10140);
nand U10336 (N_10336,N_10017,N_10029);
or U10337 (N_10337,N_10157,N_10176);
nand U10338 (N_10338,N_10001,N_10041);
or U10339 (N_10339,N_10121,N_10080);
or U10340 (N_10340,N_10185,N_10188);
xor U10341 (N_10341,N_10008,N_10095);
nor U10342 (N_10342,N_10114,N_10178);
nand U10343 (N_10343,N_10080,N_10148);
or U10344 (N_10344,N_10057,N_10052);
nor U10345 (N_10345,N_10162,N_10187);
nor U10346 (N_10346,N_10090,N_10109);
xnor U10347 (N_10347,N_10189,N_10079);
xnor U10348 (N_10348,N_10024,N_10039);
nand U10349 (N_10349,N_10035,N_10050);
xnor U10350 (N_10350,N_10124,N_10021);
and U10351 (N_10351,N_10089,N_10014);
and U10352 (N_10352,N_10196,N_10188);
and U10353 (N_10353,N_10009,N_10032);
and U10354 (N_10354,N_10037,N_10157);
nand U10355 (N_10355,N_10158,N_10196);
nand U10356 (N_10356,N_10080,N_10052);
or U10357 (N_10357,N_10177,N_10106);
nor U10358 (N_10358,N_10187,N_10139);
nand U10359 (N_10359,N_10127,N_10094);
and U10360 (N_10360,N_10134,N_10118);
xnor U10361 (N_10361,N_10043,N_10035);
nand U10362 (N_10362,N_10128,N_10112);
xor U10363 (N_10363,N_10053,N_10188);
and U10364 (N_10364,N_10187,N_10138);
xor U10365 (N_10365,N_10010,N_10032);
nor U10366 (N_10366,N_10063,N_10154);
xor U10367 (N_10367,N_10095,N_10124);
or U10368 (N_10368,N_10073,N_10188);
xor U10369 (N_10369,N_10008,N_10135);
xnor U10370 (N_10370,N_10182,N_10156);
and U10371 (N_10371,N_10167,N_10100);
xnor U10372 (N_10372,N_10081,N_10083);
nand U10373 (N_10373,N_10129,N_10065);
xor U10374 (N_10374,N_10123,N_10067);
or U10375 (N_10375,N_10134,N_10051);
and U10376 (N_10376,N_10175,N_10171);
nor U10377 (N_10377,N_10136,N_10054);
nand U10378 (N_10378,N_10012,N_10027);
nand U10379 (N_10379,N_10015,N_10154);
and U10380 (N_10380,N_10062,N_10070);
nor U10381 (N_10381,N_10022,N_10098);
nor U10382 (N_10382,N_10124,N_10036);
nand U10383 (N_10383,N_10110,N_10069);
nand U10384 (N_10384,N_10185,N_10130);
and U10385 (N_10385,N_10021,N_10167);
nor U10386 (N_10386,N_10097,N_10011);
xnor U10387 (N_10387,N_10050,N_10039);
and U10388 (N_10388,N_10029,N_10035);
and U10389 (N_10389,N_10131,N_10158);
or U10390 (N_10390,N_10126,N_10131);
nor U10391 (N_10391,N_10042,N_10174);
and U10392 (N_10392,N_10168,N_10056);
xnor U10393 (N_10393,N_10039,N_10000);
nor U10394 (N_10394,N_10047,N_10124);
and U10395 (N_10395,N_10069,N_10020);
or U10396 (N_10396,N_10004,N_10103);
and U10397 (N_10397,N_10132,N_10075);
or U10398 (N_10398,N_10029,N_10151);
nand U10399 (N_10399,N_10047,N_10039);
and U10400 (N_10400,N_10247,N_10264);
or U10401 (N_10401,N_10313,N_10328);
nand U10402 (N_10402,N_10315,N_10241);
xnor U10403 (N_10403,N_10251,N_10349);
or U10404 (N_10404,N_10334,N_10389);
nor U10405 (N_10405,N_10292,N_10326);
and U10406 (N_10406,N_10359,N_10351);
xor U10407 (N_10407,N_10387,N_10347);
and U10408 (N_10408,N_10312,N_10288);
nand U10409 (N_10409,N_10289,N_10262);
xnor U10410 (N_10410,N_10290,N_10371);
or U10411 (N_10411,N_10240,N_10339);
or U10412 (N_10412,N_10254,N_10203);
and U10413 (N_10413,N_10310,N_10331);
nor U10414 (N_10414,N_10305,N_10274);
nor U10415 (N_10415,N_10279,N_10329);
and U10416 (N_10416,N_10285,N_10232);
and U10417 (N_10417,N_10294,N_10260);
or U10418 (N_10418,N_10252,N_10237);
nor U10419 (N_10419,N_10327,N_10301);
nand U10420 (N_10420,N_10317,N_10300);
nor U10421 (N_10421,N_10207,N_10379);
nand U10422 (N_10422,N_10276,N_10204);
xnor U10423 (N_10423,N_10297,N_10394);
or U10424 (N_10424,N_10235,N_10293);
and U10425 (N_10425,N_10298,N_10218);
xnor U10426 (N_10426,N_10302,N_10374);
and U10427 (N_10427,N_10304,N_10299);
or U10428 (N_10428,N_10219,N_10388);
nor U10429 (N_10429,N_10200,N_10272);
and U10430 (N_10430,N_10324,N_10261);
and U10431 (N_10431,N_10287,N_10356);
nand U10432 (N_10432,N_10229,N_10248);
and U10433 (N_10433,N_10238,N_10354);
xor U10434 (N_10434,N_10314,N_10263);
xnor U10435 (N_10435,N_10378,N_10385);
nor U10436 (N_10436,N_10233,N_10363);
or U10437 (N_10437,N_10367,N_10373);
and U10438 (N_10438,N_10319,N_10375);
nand U10439 (N_10439,N_10393,N_10391);
nand U10440 (N_10440,N_10335,N_10392);
nand U10441 (N_10441,N_10355,N_10268);
nand U10442 (N_10442,N_10230,N_10205);
nor U10443 (N_10443,N_10212,N_10234);
nand U10444 (N_10444,N_10353,N_10358);
nor U10445 (N_10445,N_10361,N_10253);
or U10446 (N_10446,N_10250,N_10221);
xnor U10447 (N_10447,N_10368,N_10210);
and U10448 (N_10448,N_10365,N_10398);
and U10449 (N_10449,N_10303,N_10325);
xnor U10450 (N_10450,N_10377,N_10357);
nand U10451 (N_10451,N_10350,N_10201);
nor U10452 (N_10452,N_10364,N_10372);
and U10453 (N_10453,N_10216,N_10369);
xnor U10454 (N_10454,N_10236,N_10208);
nor U10455 (N_10455,N_10333,N_10346);
nand U10456 (N_10456,N_10281,N_10311);
nand U10457 (N_10457,N_10383,N_10270);
xor U10458 (N_10458,N_10228,N_10245);
nand U10459 (N_10459,N_10224,N_10376);
and U10460 (N_10460,N_10370,N_10257);
xor U10461 (N_10461,N_10362,N_10213);
nor U10462 (N_10462,N_10283,N_10399);
nor U10463 (N_10463,N_10226,N_10244);
and U10464 (N_10464,N_10223,N_10381);
xnor U10465 (N_10465,N_10348,N_10306);
nand U10466 (N_10466,N_10343,N_10323);
or U10467 (N_10467,N_10269,N_10266);
and U10468 (N_10468,N_10242,N_10337);
and U10469 (N_10469,N_10214,N_10278);
and U10470 (N_10470,N_10342,N_10295);
nand U10471 (N_10471,N_10209,N_10382);
and U10472 (N_10472,N_10286,N_10338);
and U10473 (N_10473,N_10215,N_10395);
nor U10474 (N_10474,N_10309,N_10296);
nand U10475 (N_10475,N_10259,N_10291);
and U10476 (N_10476,N_10202,N_10316);
nand U10477 (N_10477,N_10322,N_10220);
or U10478 (N_10478,N_10341,N_10231);
nand U10479 (N_10479,N_10336,N_10249);
nor U10480 (N_10480,N_10318,N_10256);
nand U10481 (N_10481,N_10255,N_10384);
or U10482 (N_10482,N_10330,N_10277);
and U10483 (N_10483,N_10282,N_10397);
and U10484 (N_10484,N_10321,N_10225);
and U10485 (N_10485,N_10258,N_10284);
nand U10486 (N_10486,N_10211,N_10307);
nor U10487 (N_10487,N_10345,N_10352);
nand U10488 (N_10488,N_10217,N_10239);
or U10489 (N_10489,N_10271,N_10267);
and U10490 (N_10490,N_10308,N_10366);
nor U10491 (N_10491,N_10390,N_10344);
and U10492 (N_10492,N_10332,N_10396);
nand U10493 (N_10493,N_10206,N_10340);
or U10494 (N_10494,N_10246,N_10280);
xor U10495 (N_10495,N_10320,N_10222);
xnor U10496 (N_10496,N_10265,N_10243);
nor U10497 (N_10497,N_10275,N_10380);
and U10498 (N_10498,N_10386,N_10227);
nor U10499 (N_10499,N_10360,N_10273);
and U10500 (N_10500,N_10222,N_10242);
nor U10501 (N_10501,N_10342,N_10228);
xnor U10502 (N_10502,N_10393,N_10337);
nor U10503 (N_10503,N_10368,N_10284);
nand U10504 (N_10504,N_10295,N_10213);
xnor U10505 (N_10505,N_10353,N_10370);
nand U10506 (N_10506,N_10393,N_10290);
and U10507 (N_10507,N_10211,N_10330);
nand U10508 (N_10508,N_10362,N_10296);
nor U10509 (N_10509,N_10297,N_10200);
xor U10510 (N_10510,N_10345,N_10252);
xor U10511 (N_10511,N_10270,N_10336);
or U10512 (N_10512,N_10219,N_10228);
or U10513 (N_10513,N_10375,N_10304);
or U10514 (N_10514,N_10259,N_10277);
nor U10515 (N_10515,N_10242,N_10334);
or U10516 (N_10516,N_10299,N_10360);
nor U10517 (N_10517,N_10352,N_10306);
or U10518 (N_10518,N_10384,N_10332);
xnor U10519 (N_10519,N_10384,N_10315);
nor U10520 (N_10520,N_10203,N_10365);
nand U10521 (N_10521,N_10284,N_10331);
and U10522 (N_10522,N_10212,N_10376);
or U10523 (N_10523,N_10383,N_10360);
nand U10524 (N_10524,N_10296,N_10276);
nor U10525 (N_10525,N_10244,N_10250);
and U10526 (N_10526,N_10321,N_10356);
or U10527 (N_10527,N_10208,N_10386);
and U10528 (N_10528,N_10211,N_10341);
nand U10529 (N_10529,N_10279,N_10303);
nor U10530 (N_10530,N_10295,N_10274);
or U10531 (N_10531,N_10265,N_10210);
xnor U10532 (N_10532,N_10280,N_10216);
or U10533 (N_10533,N_10206,N_10208);
nor U10534 (N_10534,N_10331,N_10202);
and U10535 (N_10535,N_10240,N_10344);
and U10536 (N_10536,N_10348,N_10288);
xnor U10537 (N_10537,N_10397,N_10268);
xnor U10538 (N_10538,N_10230,N_10382);
xor U10539 (N_10539,N_10276,N_10329);
or U10540 (N_10540,N_10387,N_10291);
or U10541 (N_10541,N_10371,N_10320);
xnor U10542 (N_10542,N_10384,N_10328);
and U10543 (N_10543,N_10278,N_10391);
nor U10544 (N_10544,N_10297,N_10301);
or U10545 (N_10545,N_10201,N_10377);
and U10546 (N_10546,N_10270,N_10330);
and U10547 (N_10547,N_10372,N_10209);
or U10548 (N_10548,N_10378,N_10369);
or U10549 (N_10549,N_10249,N_10212);
xor U10550 (N_10550,N_10253,N_10280);
and U10551 (N_10551,N_10227,N_10202);
nand U10552 (N_10552,N_10317,N_10302);
or U10553 (N_10553,N_10207,N_10201);
or U10554 (N_10554,N_10341,N_10200);
and U10555 (N_10555,N_10289,N_10321);
or U10556 (N_10556,N_10358,N_10368);
nor U10557 (N_10557,N_10308,N_10255);
nand U10558 (N_10558,N_10311,N_10347);
or U10559 (N_10559,N_10395,N_10239);
or U10560 (N_10560,N_10327,N_10312);
and U10561 (N_10561,N_10334,N_10272);
or U10562 (N_10562,N_10257,N_10226);
or U10563 (N_10563,N_10355,N_10261);
and U10564 (N_10564,N_10231,N_10263);
and U10565 (N_10565,N_10280,N_10326);
xnor U10566 (N_10566,N_10215,N_10280);
or U10567 (N_10567,N_10373,N_10205);
nand U10568 (N_10568,N_10211,N_10394);
nor U10569 (N_10569,N_10270,N_10353);
or U10570 (N_10570,N_10255,N_10238);
xnor U10571 (N_10571,N_10370,N_10284);
xor U10572 (N_10572,N_10372,N_10356);
and U10573 (N_10573,N_10307,N_10356);
xnor U10574 (N_10574,N_10330,N_10310);
or U10575 (N_10575,N_10351,N_10253);
and U10576 (N_10576,N_10391,N_10296);
or U10577 (N_10577,N_10333,N_10236);
or U10578 (N_10578,N_10271,N_10273);
nand U10579 (N_10579,N_10279,N_10342);
and U10580 (N_10580,N_10362,N_10205);
nand U10581 (N_10581,N_10299,N_10288);
nor U10582 (N_10582,N_10397,N_10331);
xor U10583 (N_10583,N_10359,N_10300);
xnor U10584 (N_10584,N_10218,N_10377);
nand U10585 (N_10585,N_10265,N_10346);
nand U10586 (N_10586,N_10334,N_10366);
nor U10587 (N_10587,N_10222,N_10201);
and U10588 (N_10588,N_10216,N_10294);
nor U10589 (N_10589,N_10322,N_10218);
nand U10590 (N_10590,N_10303,N_10302);
xor U10591 (N_10591,N_10277,N_10367);
nand U10592 (N_10592,N_10324,N_10250);
and U10593 (N_10593,N_10237,N_10251);
or U10594 (N_10594,N_10399,N_10314);
nor U10595 (N_10595,N_10256,N_10224);
or U10596 (N_10596,N_10373,N_10217);
xnor U10597 (N_10597,N_10216,N_10240);
and U10598 (N_10598,N_10226,N_10239);
or U10599 (N_10599,N_10251,N_10386);
xor U10600 (N_10600,N_10461,N_10515);
xnor U10601 (N_10601,N_10408,N_10528);
xor U10602 (N_10602,N_10451,N_10457);
xor U10603 (N_10603,N_10508,N_10525);
nand U10604 (N_10604,N_10474,N_10427);
nor U10605 (N_10605,N_10547,N_10467);
or U10606 (N_10606,N_10540,N_10439);
nand U10607 (N_10607,N_10598,N_10443);
nor U10608 (N_10608,N_10506,N_10596);
or U10609 (N_10609,N_10502,N_10458);
and U10610 (N_10610,N_10432,N_10471);
nand U10611 (N_10611,N_10588,N_10494);
xnor U10612 (N_10612,N_10568,N_10485);
or U10613 (N_10613,N_10593,N_10530);
nor U10614 (N_10614,N_10406,N_10520);
nand U10615 (N_10615,N_10483,N_10511);
nor U10616 (N_10616,N_10590,N_10534);
and U10617 (N_10617,N_10573,N_10437);
nand U10618 (N_10618,N_10463,N_10442);
or U10619 (N_10619,N_10479,N_10527);
or U10620 (N_10620,N_10415,N_10510);
or U10621 (N_10621,N_10517,N_10433);
nand U10622 (N_10622,N_10497,N_10484);
or U10623 (N_10623,N_10566,N_10401);
nor U10624 (N_10624,N_10412,N_10435);
nor U10625 (N_10625,N_10441,N_10585);
xnor U10626 (N_10626,N_10482,N_10542);
and U10627 (N_10627,N_10402,N_10560);
xnor U10628 (N_10628,N_10426,N_10545);
nor U10629 (N_10629,N_10516,N_10594);
xnor U10630 (N_10630,N_10543,N_10513);
nor U10631 (N_10631,N_10505,N_10559);
nand U10632 (N_10632,N_10551,N_10445);
and U10633 (N_10633,N_10428,N_10583);
nor U10634 (N_10634,N_10587,N_10417);
or U10635 (N_10635,N_10486,N_10538);
and U10636 (N_10636,N_10514,N_10422);
and U10637 (N_10637,N_10575,N_10521);
or U10638 (N_10638,N_10470,N_10565);
or U10639 (N_10639,N_10400,N_10546);
nand U10640 (N_10640,N_10592,N_10487);
nor U10641 (N_10641,N_10431,N_10599);
or U10642 (N_10642,N_10446,N_10450);
and U10643 (N_10643,N_10548,N_10570);
and U10644 (N_10644,N_10518,N_10492);
nand U10645 (N_10645,N_10434,N_10473);
or U10646 (N_10646,N_10569,N_10584);
nand U10647 (N_10647,N_10454,N_10581);
and U10648 (N_10648,N_10453,N_10481);
and U10649 (N_10649,N_10562,N_10448);
xor U10650 (N_10650,N_10591,N_10577);
nor U10651 (N_10651,N_10475,N_10522);
nor U10652 (N_10652,N_10444,N_10589);
nor U10653 (N_10653,N_10436,N_10491);
or U10654 (N_10654,N_10465,N_10407);
nor U10655 (N_10655,N_10567,N_10504);
nand U10656 (N_10656,N_10489,N_10424);
nand U10657 (N_10657,N_10477,N_10468);
xnor U10658 (N_10658,N_10419,N_10541);
xnor U10659 (N_10659,N_10418,N_10411);
and U10660 (N_10660,N_10531,N_10563);
nand U10661 (N_10661,N_10509,N_10440);
or U10662 (N_10662,N_10549,N_10466);
xor U10663 (N_10663,N_10574,N_10580);
xnor U10664 (N_10664,N_10552,N_10526);
or U10665 (N_10665,N_10519,N_10572);
or U10666 (N_10666,N_10423,N_10480);
or U10667 (N_10667,N_10452,N_10539);
nor U10668 (N_10668,N_10564,N_10455);
or U10669 (N_10669,N_10462,N_10533);
or U10670 (N_10670,N_10529,N_10512);
and U10671 (N_10671,N_10456,N_10558);
and U10672 (N_10672,N_10536,N_10421);
or U10673 (N_10673,N_10524,N_10576);
xor U10674 (N_10674,N_10537,N_10557);
nor U10675 (N_10675,N_10579,N_10472);
or U10676 (N_10676,N_10523,N_10405);
and U10677 (N_10677,N_10488,N_10420);
xor U10678 (N_10678,N_10501,N_10498);
or U10679 (N_10679,N_10404,N_10403);
and U10680 (N_10680,N_10447,N_10550);
nand U10681 (N_10681,N_10430,N_10459);
nor U10682 (N_10682,N_10535,N_10571);
nor U10683 (N_10683,N_10553,N_10595);
xnor U10684 (N_10684,N_10414,N_10495);
nand U10685 (N_10685,N_10469,N_10429);
xnor U10686 (N_10686,N_10582,N_10425);
xnor U10687 (N_10687,N_10496,N_10556);
nand U10688 (N_10688,N_10554,N_10410);
and U10689 (N_10689,N_10561,N_10578);
nand U10690 (N_10690,N_10507,N_10555);
xnor U10691 (N_10691,N_10503,N_10464);
nand U10692 (N_10692,N_10493,N_10597);
nor U10693 (N_10693,N_10438,N_10409);
or U10694 (N_10694,N_10490,N_10586);
xnor U10695 (N_10695,N_10413,N_10449);
nor U10696 (N_10696,N_10544,N_10416);
nor U10697 (N_10697,N_10532,N_10460);
or U10698 (N_10698,N_10499,N_10478);
nand U10699 (N_10699,N_10500,N_10476);
xnor U10700 (N_10700,N_10595,N_10560);
nand U10701 (N_10701,N_10591,N_10473);
xnor U10702 (N_10702,N_10449,N_10559);
nand U10703 (N_10703,N_10514,N_10532);
and U10704 (N_10704,N_10595,N_10429);
nand U10705 (N_10705,N_10594,N_10518);
xor U10706 (N_10706,N_10532,N_10442);
nor U10707 (N_10707,N_10493,N_10465);
nor U10708 (N_10708,N_10513,N_10402);
and U10709 (N_10709,N_10567,N_10594);
xor U10710 (N_10710,N_10566,N_10562);
or U10711 (N_10711,N_10501,N_10429);
and U10712 (N_10712,N_10482,N_10507);
nor U10713 (N_10713,N_10484,N_10576);
or U10714 (N_10714,N_10429,N_10412);
nand U10715 (N_10715,N_10436,N_10439);
nand U10716 (N_10716,N_10419,N_10496);
xnor U10717 (N_10717,N_10547,N_10462);
nand U10718 (N_10718,N_10460,N_10541);
nor U10719 (N_10719,N_10476,N_10571);
or U10720 (N_10720,N_10576,N_10497);
and U10721 (N_10721,N_10465,N_10479);
nor U10722 (N_10722,N_10515,N_10422);
nand U10723 (N_10723,N_10488,N_10554);
and U10724 (N_10724,N_10519,N_10563);
xnor U10725 (N_10725,N_10590,N_10449);
xnor U10726 (N_10726,N_10433,N_10594);
or U10727 (N_10727,N_10577,N_10414);
xnor U10728 (N_10728,N_10404,N_10406);
or U10729 (N_10729,N_10505,N_10407);
nor U10730 (N_10730,N_10437,N_10430);
nand U10731 (N_10731,N_10524,N_10536);
and U10732 (N_10732,N_10545,N_10598);
xor U10733 (N_10733,N_10516,N_10551);
and U10734 (N_10734,N_10570,N_10466);
or U10735 (N_10735,N_10453,N_10462);
or U10736 (N_10736,N_10441,N_10562);
or U10737 (N_10737,N_10439,N_10482);
or U10738 (N_10738,N_10404,N_10459);
nor U10739 (N_10739,N_10517,N_10482);
and U10740 (N_10740,N_10599,N_10421);
nand U10741 (N_10741,N_10587,N_10576);
nor U10742 (N_10742,N_10407,N_10458);
or U10743 (N_10743,N_10521,N_10410);
nor U10744 (N_10744,N_10537,N_10549);
or U10745 (N_10745,N_10429,N_10447);
or U10746 (N_10746,N_10402,N_10573);
and U10747 (N_10747,N_10423,N_10508);
or U10748 (N_10748,N_10415,N_10413);
nand U10749 (N_10749,N_10581,N_10541);
nor U10750 (N_10750,N_10403,N_10580);
xnor U10751 (N_10751,N_10540,N_10478);
and U10752 (N_10752,N_10558,N_10574);
nand U10753 (N_10753,N_10458,N_10505);
xnor U10754 (N_10754,N_10554,N_10540);
nor U10755 (N_10755,N_10535,N_10510);
nor U10756 (N_10756,N_10490,N_10527);
xor U10757 (N_10757,N_10569,N_10524);
and U10758 (N_10758,N_10512,N_10533);
nand U10759 (N_10759,N_10458,N_10541);
xnor U10760 (N_10760,N_10469,N_10478);
nor U10761 (N_10761,N_10456,N_10458);
nand U10762 (N_10762,N_10539,N_10482);
and U10763 (N_10763,N_10575,N_10565);
nor U10764 (N_10764,N_10524,N_10467);
and U10765 (N_10765,N_10466,N_10543);
and U10766 (N_10766,N_10584,N_10572);
nand U10767 (N_10767,N_10450,N_10408);
or U10768 (N_10768,N_10525,N_10496);
xor U10769 (N_10769,N_10472,N_10506);
xnor U10770 (N_10770,N_10457,N_10558);
xor U10771 (N_10771,N_10454,N_10495);
or U10772 (N_10772,N_10582,N_10455);
nor U10773 (N_10773,N_10451,N_10435);
xnor U10774 (N_10774,N_10458,N_10404);
and U10775 (N_10775,N_10526,N_10558);
or U10776 (N_10776,N_10556,N_10595);
nand U10777 (N_10777,N_10444,N_10458);
xnor U10778 (N_10778,N_10519,N_10503);
nand U10779 (N_10779,N_10521,N_10452);
and U10780 (N_10780,N_10584,N_10514);
xor U10781 (N_10781,N_10589,N_10420);
and U10782 (N_10782,N_10588,N_10514);
and U10783 (N_10783,N_10420,N_10533);
and U10784 (N_10784,N_10435,N_10545);
xnor U10785 (N_10785,N_10464,N_10445);
and U10786 (N_10786,N_10425,N_10531);
and U10787 (N_10787,N_10430,N_10476);
xor U10788 (N_10788,N_10579,N_10417);
or U10789 (N_10789,N_10534,N_10455);
nand U10790 (N_10790,N_10491,N_10417);
nand U10791 (N_10791,N_10554,N_10538);
nand U10792 (N_10792,N_10581,N_10416);
nor U10793 (N_10793,N_10553,N_10433);
or U10794 (N_10794,N_10463,N_10426);
xnor U10795 (N_10795,N_10474,N_10449);
nor U10796 (N_10796,N_10447,N_10522);
and U10797 (N_10797,N_10589,N_10487);
xnor U10798 (N_10798,N_10421,N_10519);
xor U10799 (N_10799,N_10526,N_10529);
or U10800 (N_10800,N_10718,N_10747);
or U10801 (N_10801,N_10659,N_10685);
and U10802 (N_10802,N_10712,N_10754);
xnor U10803 (N_10803,N_10603,N_10622);
nand U10804 (N_10804,N_10767,N_10757);
nor U10805 (N_10805,N_10691,N_10615);
or U10806 (N_10806,N_10710,N_10611);
nor U10807 (N_10807,N_10764,N_10794);
nand U10808 (N_10808,N_10728,N_10660);
and U10809 (N_10809,N_10662,N_10639);
nand U10810 (N_10810,N_10608,N_10657);
nor U10811 (N_10811,N_10715,N_10700);
xnor U10812 (N_10812,N_10768,N_10698);
and U10813 (N_10813,N_10630,N_10778);
nand U10814 (N_10814,N_10649,N_10644);
nand U10815 (N_10815,N_10779,N_10797);
and U10816 (N_10816,N_10762,N_10738);
nand U10817 (N_10817,N_10701,N_10618);
nor U10818 (N_10818,N_10719,N_10687);
nand U10819 (N_10819,N_10634,N_10651);
xnor U10820 (N_10820,N_10785,N_10627);
nor U10821 (N_10821,N_10777,N_10645);
xnor U10822 (N_10822,N_10646,N_10695);
nand U10823 (N_10823,N_10723,N_10722);
nand U10824 (N_10824,N_10666,N_10694);
xnor U10825 (N_10825,N_10705,N_10771);
or U10826 (N_10826,N_10652,N_10752);
or U10827 (N_10827,N_10606,N_10616);
nand U10828 (N_10828,N_10744,N_10766);
and U10829 (N_10829,N_10733,N_10671);
nor U10830 (N_10830,N_10656,N_10610);
or U10831 (N_10831,N_10650,N_10625);
nor U10832 (N_10832,N_10655,N_10780);
and U10833 (N_10833,N_10774,N_10690);
xnor U10834 (N_10834,N_10748,N_10665);
nand U10835 (N_10835,N_10612,N_10734);
and U10836 (N_10836,N_10727,N_10732);
or U10837 (N_10837,N_10654,N_10759);
xor U10838 (N_10838,N_10647,N_10729);
and U10839 (N_10839,N_10784,N_10730);
xnor U10840 (N_10840,N_10702,N_10623);
nor U10841 (N_10841,N_10772,N_10663);
nor U10842 (N_10842,N_10709,N_10721);
nor U10843 (N_10843,N_10795,N_10787);
or U10844 (N_10844,N_10624,N_10796);
nor U10845 (N_10845,N_10620,N_10628);
nor U10846 (N_10846,N_10720,N_10664);
and U10847 (N_10847,N_10783,N_10745);
or U10848 (N_10848,N_10740,N_10632);
and U10849 (N_10849,N_10776,N_10689);
or U10850 (N_10850,N_10604,N_10761);
xor U10851 (N_10851,N_10641,N_10725);
xnor U10852 (N_10852,N_10600,N_10792);
or U10853 (N_10853,N_10640,N_10708);
and U10854 (N_10854,N_10679,N_10668);
nand U10855 (N_10855,N_10683,N_10697);
xnor U10856 (N_10856,N_10706,N_10653);
nand U10857 (N_10857,N_10619,N_10642);
xnor U10858 (N_10858,N_10741,N_10799);
xor U10859 (N_10859,N_10756,N_10621);
and U10860 (N_10860,N_10688,N_10724);
xnor U10861 (N_10861,N_10613,N_10692);
or U10862 (N_10862,N_10770,N_10765);
nand U10863 (N_10863,N_10601,N_10782);
or U10864 (N_10864,N_10775,N_10677);
and U10865 (N_10865,N_10680,N_10696);
xnor U10866 (N_10866,N_10674,N_10758);
nand U10867 (N_10867,N_10763,N_10798);
xnor U10868 (N_10868,N_10617,N_10614);
and U10869 (N_10869,N_10714,N_10633);
nor U10870 (N_10870,N_10676,N_10648);
or U10871 (N_10871,N_10681,N_10751);
and U10872 (N_10872,N_10682,N_10699);
nor U10873 (N_10873,N_10661,N_10638);
nand U10874 (N_10874,N_10675,N_10791);
and U10875 (N_10875,N_10605,N_10790);
and U10876 (N_10876,N_10673,N_10789);
nor U10877 (N_10877,N_10669,N_10635);
or U10878 (N_10878,N_10755,N_10760);
nand U10879 (N_10879,N_10717,N_10667);
nand U10880 (N_10880,N_10711,N_10629);
and U10881 (N_10881,N_10786,N_10672);
and U10882 (N_10882,N_10750,N_10742);
nor U10883 (N_10883,N_10746,N_10686);
nand U10884 (N_10884,N_10753,N_10643);
nand U10885 (N_10885,N_10684,N_10735);
nand U10886 (N_10886,N_10631,N_10749);
and U10887 (N_10887,N_10703,N_10781);
nand U10888 (N_10888,N_10607,N_10693);
nand U10889 (N_10889,N_10713,N_10609);
nand U10890 (N_10890,N_10739,N_10716);
nor U10891 (N_10891,N_10731,N_10737);
and U10892 (N_10892,N_10707,N_10743);
nand U10893 (N_10893,N_10636,N_10736);
or U10894 (N_10894,N_10670,N_10726);
nor U10895 (N_10895,N_10626,N_10793);
xnor U10896 (N_10896,N_10773,N_10658);
and U10897 (N_10897,N_10637,N_10602);
xnor U10898 (N_10898,N_10704,N_10678);
xnor U10899 (N_10899,N_10769,N_10788);
or U10900 (N_10900,N_10790,N_10616);
and U10901 (N_10901,N_10637,N_10692);
xor U10902 (N_10902,N_10611,N_10746);
nand U10903 (N_10903,N_10634,N_10757);
or U10904 (N_10904,N_10630,N_10672);
nand U10905 (N_10905,N_10604,N_10717);
nand U10906 (N_10906,N_10763,N_10741);
and U10907 (N_10907,N_10750,N_10652);
nor U10908 (N_10908,N_10683,N_10611);
nor U10909 (N_10909,N_10682,N_10641);
or U10910 (N_10910,N_10687,N_10799);
and U10911 (N_10911,N_10730,N_10778);
or U10912 (N_10912,N_10678,N_10740);
nand U10913 (N_10913,N_10786,N_10788);
and U10914 (N_10914,N_10634,N_10630);
xnor U10915 (N_10915,N_10689,N_10752);
xnor U10916 (N_10916,N_10680,N_10745);
nor U10917 (N_10917,N_10790,N_10668);
and U10918 (N_10918,N_10674,N_10737);
nand U10919 (N_10919,N_10615,N_10611);
and U10920 (N_10920,N_10747,N_10731);
and U10921 (N_10921,N_10614,N_10668);
nor U10922 (N_10922,N_10770,N_10739);
xnor U10923 (N_10923,N_10673,N_10794);
and U10924 (N_10924,N_10794,N_10656);
xnor U10925 (N_10925,N_10702,N_10606);
nor U10926 (N_10926,N_10677,N_10609);
and U10927 (N_10927,N_10778,N_10608);
nor U10928 (N_10928,N_10707,N_10691);
or U10929 (N_10929,N_10693,N_10638);
and U10930 (N_10930,N_10613,N_10769);
xor U10931 (N_10931,N_10767,N_10656);
nand U10932 (N_10932,N_10687,N_10772);
nor U10933 (N_10933,N_10740,N_10630);
nand U10934 (N_10934,N_10791,N_10797);
nand U10935 (N_10935,N_10674,N_10614);
nand U10936 (N_10936,N_10794,N_10608);
xor U10937 (N_10937,N_10603,N_10646);
nor U10938 (N_10938,N_10689,N_10772);
xor U10939 (N_10939,N_10727,N_10723);
nand U10940 (N_10940,N_10689,N_10620);
or U10941 (N_10941,N_10639,N_10707);
nand U10942 (N_10942,N_10614,N_10673);
or U10943 (N_10943,N_10725,N_10777);
xnor U10944 (N_10944,N_10664,N_10685);
and U10945 (N_10945,N_10712,N_10730);
or U10946 (N_10946,N_10648,N_10647);
or U10947 (N_10947,N_10678,N_10670);
xnor U10948 (N_10948,N_10604,N_10641);
and U10949 (N_10949,N_10636,N_10776);
nand U10950 (N_10950,N_10648,N_10733);
or U10951 (N_10951,N_10676,N_10726);
nor U10952 (N_10952,N_10740,N_10749);
nand U10953 (N_10953,N_10685,N_10768);
nor U10954 (N_10954,N_10674,N_10742);
nor U10955 (N_10955,N_10755,N_10756);
and U10956 (N_10956,N_10742,N_10775);
and U10957 (N_10957,N_10681,N_10647);
or U10958 (N_10958,N_10763,N_10704);
or U10959 (N_10959,N_10642,N_10687);
nor U10960 (N_10960,N_10696,N_10692);
and U10961 (N_10961,N_10758,N_10729);
nor U10962 (N_10962,N_10616,N_10732);
xnor U10963 (N_10963,N_10684,N_10749);
or U10964 (N_10964,N_10783,N_10708);
nor U10965 (N_10965,N_10797,N_10622);
xnor U10966 (N_10966,N_10774,N_10724);
xnor U10967 (N_10967,N_10619,N_10703);
nand U10968 (N_10968,N_10737,N_10799);
or U10969 (N_10969,N_10616,N_10651);
or U10970 (N_10970,N_10662,N_10727);
and U10971 (N_10971,N_10615,N_10798);
and U10972 (N_10972,N_10655,N_10794);
xnor U10973 (N_10973,N_10789,N_10786);
nor U10974 (N_10974,N_10728,N_10653);
or U10975 (N_10975,N_10766,N_10769);
or U10976 (N_10976,N_10731,N_10742);
and U10977 (N_10977,N_10670,N_10788);
xor U10978 (N_10978,N_10660,N_10654);
xor U10979 (N_10979,N_10624,N_10799);
nand U10980 (N_10980,N_10616,N_10783);
nor U10981 (N_10981,N_10774,N_10732);
and U10982 (N_10982,N_10652,N_10609);
nand U10983 (N_10983,N_10752,N_10684);
and U10984 (N_10984,N_10799,N_10692);
nand U10985 (N_10985,N_10780,N_10744);
and U10986 (N_10986,N_10717,N_10635);
xnor U10987 (N_10987,N_10713,N_10786);
nand U10988 (N_10988,N_10798,N_10656);
or U10989 (N_10989,N_10672,N_10724);
and U10990 (N_10990,N_10695,N_10714);
nand U10991 (N_10991,N_10658,N_10791);
and U10992 (N_10992,N_10720,N_10641);
xor U10993 (N_10993,N_10709,N_10785);
and U10994 (N_10994,N_10631,N_10784);
nand U10995 (N_10995,N_10692,N_10682);
and U10996 (N_10996,N_10602,N_10688);
xor U10997 (N_10997,N_10724,N_10603);
nor U10998 (N_10998,N_10748,N_10698);
nand U10999 (N_10999,N_10746,N_10659);
nand U11000 (N_11000,N_10923,N_10845);
or U11001 (N_11001,N_10810,N_10830);
nand U11002 (N_11002,N_10939,N_10984);
xnor U11003 (N_11003,N_10801,N_10970);
or U11004 (N_11004,N_10893,N_10943);
or U11005 (N_11005,N_10915,N_10898);
or U11006 (N_11006,N_10849,N_10965);
or U11007 (N_11007,N_10877,N_10823);
nand U11008 (N_11008,N_10838,N_10944);
xor U11009 (N_11009,N_10859,N_10816);
nor U11010 (N_11010,N_10804,N_10919);
nand U11011 (N_11011,N_10864,N_10843);
nand U11012 (N_11012,N_10917,N_10950);
or U11013 (N_11013,N_10806,N_10985);
xor U11014 (N_11014,N_10883,N_10924);
nand U11015 (N_11015,N_10867,N_10896);
nor U11016 (N_11016,N_10857,N_10871);
and U11017 (N_11017,N_10821,N_10907);
xnor U11018 (N_11018,N_10987,N_10989);
nand U11019 (N_11019,N_10834,N_10892);
nand U11020 (N_11020,N_10862,N_10828);
and U11021 (N_11021,N_10929,N_10901);
and U11022 (N_11022,N_10914,N_10941);
nor U11023 (N_11023,N_10990,N_10868);
nor U11024 (N_11024,N_10889,N_10906);
or U11025 (N_11025,N_10826,N_10997);
nand U11026 (N_11026,N_10986,N_10932);
nand U11027 (N_11027,N_10820,N_10953);
or U11028 (N_11028,N_10831,N_10994);
xnor U11029 (N_11029,N_10888,N_10962);
nor U11030 (N_11030,N_10832,N_10975);
or U11031 (N_11031,N_10860,N_10957);
nand U11032 (N_11032,N_10921,N_10937);
xnor U11033 (N_11033,N_10809,N_10948);
or U11034 (N_11034,N_10951,N_10960);
and U11035 (N_11035,N_10934,N_10972);
nand U11036 (N_11036,N_10829,N_10863);
xnor U11037 (N_11037,N_10991,N_10886);
nor U11038 (N_11038,N_10813,N_10876);
or U11039 (N_11039,N_10833,N_10897);
and U11040 (N_11040,N_10865,N_10947);
or U11041 (N_11041,N_10817,N_10908);
and U11042 (N_11042,N_10979,N_10909);
nand U11043 (N_11043,N_10993,N_10861);
nand U11044 (N_11044,N_10968,N_10977);
nor U11045 (N_11045,N_10996,N_10814);
nand U11046 (N_11046,N_10920,N_10983);
and U11047 (N_11047,N_10998,N_10928);
and U11048 (N_11048,N_10959,N_10848);
nand U11049 (N_11049,N_10884,N_10899);
nor U11050 (N_11050,N_10875,N_10945);
xnor U11051 (N_11051,N_10847,N_10927);
or U11052 (N_11052,N_10811,N_10873);
and U11053 (N_11053,N_10880,N_10842);
and U11054 (N_11054,N_10827,N_10895);
nand U11055 (N_11055,N_10916,N_10851);
xnor U11056 (N_11056,N_10844,N_10995);
nand U11057 (N_11057,N_10971,N_10910);
nand U11058 (N_11058,N_10869,N_10887);
xnor U11059 (N_11059,N_10836,N_10808);
nor U11060 (N_11060,N_10913,N_10802);
nor U11061 (N_11061,N_10940,N_10964);
or U11062 (N_11062,N_10938,N_10840);
nand U11063 (N_11063,N_10803,N_10933);
nand U11064 (N_11064,N_10800,N_10812);
and U11065 (N_11065,N_10882,N_10885);
nor U11066 (N_11066,N_10963,N_10819);
nor U11067 (N_11067,N_10988,N_10822);
nor U11068 (N_11068,N_10974,N_10825);
xnor U11069 (N_11069,N_10982,N_10911);
nand U11070 (N_11070,N_10866,N_10904);
or U11071 (N_11071,N_10835,N_10903);
and U11072 (N_11072,N_10942,N_10853);
or U11073 (N_11073,N_10858,N_10855);
nand U11074 (N_11074,N_10973,N_10931);
xnor U11075 (N_11075,N_10936,N_10879);
xor U11076 (N_11076,N_10925,N_10969);
or U11077 (N_11077,N_10874,N_10992);
and U11078 (N_11078,N_10958,N_10824);
or U11079 (N_11079,N_10850,N_10905);
nand U11080 (N_11080,N_10805,N_10837);
nor U11081 (N_11081,N_10870,N_10891);
nor U11082 (N_11082,N_10976,N_10999);
or U11083 (N_11083,N_10894,N_10900);
nand U11084 (N_11084,N_10839,N_10956);
xnor U11085 (N_11085,N_10980,N_10978);
and U11086 (N_11086,N_10846,N_10815);
nor U11087 (N_11087,N_10949,N_10881);
or U11088 (N_11088,N_10918,N_10818);
nor U11089 (N_11089,N_10966,N_10872);
nand U11090 (N_11090,N_10954,N_10926);
nand U11091 (N_11091,N_10841,N_10967);
xor U11092 (N_11092,N_10878,N_10912);
nand U11093 (N_11093,N_10856,N_10961);
xor U11094 (N_11094,N_10930,N_10946);
and U11095 (N_11095,N_10922,N_10955);
xnor U11096 (N_11096,N_10807,N_10981);
or U11097 (N_11097,N_10852,N_10854);
and U11098 (N_11098,N_10935,N_10890);
and U11099 (N_11099,N_10952,N_10902);
xnor U11100 (N_11100,N_10908,N_10942);
xnor U11101 (N_11101,N_10951,N_10989);
and U11102 (N_11102,N_10946,N_10964);
nand U11103 (N_11103,N_10852,N_10828);
xor U11104 (N_11104,N_10818,N_10883);
or U11105 (N_11105,N_10898,N_10866);
nor U11106 (N_11106,N_10890,N_10922);
nor U11107 (N_11107,N_10949,N_10826);
xnor U11108 (N_11108,N_10961,N_10850);
xnor U11109 (N_11109,N_10960,N_10825);
xnor U11110 (N_11110,N_10850,N_10885);
nor U11111 (N_11111,N_10970,N_10813);
or U11112 (N_11112,N_10855,N_10831);
and U11113 (N_11113,N_10865,N_10990);
and U11114 (N_11114,N_10814,N_10997);
xor U11115 (N_11115,N_10849,N_10844);
nor U11116 (N_11116,N_10835,N_10940);
nor U11117 (N_11117,N_10850,N_10847);
or U11118 (N_11118,N_10859,N_10986);
xor U11119 (N_11119,N_10818,N_10966);
nor U11120 (N_11120,N_10899,N_10959);
nand U11121 (N_11121,N_10819,N_10823);
nor U11122 (N_11122,N_10995,N_10962);
or U11123 (N_11123,N_10819,N_10808);
nor U11124 (N_11124,N_10805,N_10813);
nor U11125 (N_11125,N_10950,N_10872);
or U11126 (N_11126,N_10841,N_10995);
nor U11127 (N_11127,N_10842,N_10962);
and U11128 (N_11128,N_10820,N_10928);
nor U11129 (N_11129,N_10865,N_10877);
or U11130 (N_11130,N_10967,N_10830);
and U11131 (N_11131,N_10904,N_10916);
and U11132 (N_11132,N_10899,N_10871);
or U11133 (N_11133,N_10926,N_10832);
or U11134 (N_11134,N_10927,N_10867);
nand U11135 (N_11135,N_10860,N_10958);
or U11136 (N_11136,N_10803,N_10993);
nor U11137 (N_11137,N_10994,N_10870);
and U11138 (N_11138,N_10941,N_10925);
xnor U11139 (N_11139,N_10922,N_10965);
or U11140 (N_11140,N_10890,N_10981);
xor U11141 (N_11141,N_10921,N_10853);
and U11142 (N_11142,N_10906,N_10959);
xor U11143 (N_11143,N_10902,N_10838);
and U11144 (N_11144,N_10861,N_10923);
nor U11145 (N_11145,N_10980,N_10808);
nand U11146 (N_11146,N_10955,N_10950);
xor U11147 (N_11147,N_10947,N_10871);
or U11148 (N_11148,N_10894,N_10932);
or U11149 (N_11149,N_10873,N_10968);
or U11150 (N_11150,N_10876,N_10810);
xor U11151 (N_11151,N_10900,N_10910);
nor U11152 (N_11152,N_10972,N_10981);
nor U11153 (N_11153,N_10803,N_10999);
nor U11154 (N_11154,N_10846,N_10833);
xnor U11155 (N_11155,N_10915,N_10848);
nor U11156 (N_11156,N_10977,N_10851);
nor U11157 (N_11157,N_10891,N_10990);
nor U11158 (N_11158,N_10979,N_10836);
and U11159 (N_11159,N_10894,N_10881);
and U11160 (N_11160,N_10965,N_10878);
or U11161 (N_11161,N_10917,N_10891);
nand U11162 (N_11162,N_10950,N_10875);
and U11163 (N_11163,N_10974,N_10908);
or U11164 (N_11164,N_10990,N_10989);
nand U11165 (N_11165,N_10846,N_10939);
xnor U11166 (N_11166,N_10911,N_10887);
nand U11167 (N_11167,N_10865,N_10938);
nor U11168 (N_11168,N_10965,N_10800);
xnor U11169 (N_11169,N_10964,N_10885);
nor U11170 (N_11170,N_10844,N_10898);
or U11171 (N_11171,N_10953,N_10836);
or U11172 (N_11172,N_10941,N_10985);
nor U11173 (N_11173,N_10930,N_10975);
or U11174 (N_11174,N_10860,N_10922);
and U11175 (N_11175,N_10945,N_10824);
or U11176 (N_11176,N_10997,N_10823);
and U11177 (N_11177,N_10955,N_10903);
nand U11178 (N_11178,N_10922,N_10928);
xnor U11179 (N_11179,N_10946,N_10967);
nor U11180 (N_11180,N_10987,N_10983);
and U11181 (N_11181,N_10943,N_10939);
nand U11182 (N_11182,N_10844,N_10838);
nand U11183 (N_11183,N_10872,N_10928);
xnor U11184 (N_11184,N_10934,N_10835);
or U11185 (N_11185,N_10873,N_10831);
or U11186 (N_11186,N_10807,N_10864);
nand U11187 (N_11187,N_10907,N_10945);
nor U11188 (N_11188,N_10810,N_10931);
or U11189 (N_11189,N_10983,N_10918);
xor U11190 (N_11190,N_10947,N_10862);
and U11191 (N_11191,N_10887,N_10805);
nand U11192 (N_11192,N_10981,N_10913);
xor U11193 (N_11193,N_10812,N_10854);
xnor U11194 (N_11194,N_10919,N_10921);
and U11195 (N_11195,N_10909,N_10954);
nor U11196 (N_11196,N_10865,N_10917);
or U11197 (N_11197,N_10991,N_10872);
xor U11198 (N_11198,N_10806,N_10842);
nor U11199 (N_11199,N_10832,N_10848);
nor U11200 (N_11200,N_11144,N_11167);
or U11201 (N_11201,N_11113,N_11044);
or U11202 (N_11202,N_11067,N_11016);
or U11203 (N_11203,N_11065,N_11026);
and U11204 (N_11204,N_11063,N_11024);
nand U11205 (N_11205,N_11136,N_11134);
nand U11206 (N_11206,N_11176,N_11150);
nor U11207 (N_11207,N_11131,N_11194);
nor U11208 (N_11208,N_11190,N_11059);
xor U11209 (N_11209,N_11186,N_11057);
and U11210 (N_11210,N_11018,N_11162);
or U11211 (N_11211,N_11062,N_11106);
nand U11212 (N_11212,N_11074,N_11165);
xor U11213 (N_11213,N_11052,N_11175);
nand U11214 (N_11214,N_11036,N_11084);
nand U11215 (N_11215,N_11172,N_11130);
and U11216 (N_11216,N_11049,N_11058);
nor U11217 (N_11217,N_11195,N_11035);
and U11218 (N_11218,N_11073,N_11086);
and U11219 (N_11219,N_11191,N_11145);
nand U11220 (N_11220,N_11091,N_11142);
xor U11221 (N_11221,N_11196,N_11140);
nand U11222 (N_11222,N_11048,N_11071);
and U11223 (N_11223,N_11043,N_11087);
nand U11224 (N_11224,N_11025,N_11115);
nand U11225 (N_11225,N_11001,N_11139);
nor U11226 (N_11226,N_11080,N_11055);
xor U11227 (N_11227,N_11119,N_11111);
or U11228 (N_11228,N_11120,N_11112);
and U11229 (N_11229,N_11011,N_11143);
xnor U11230 (N_11230,N_11008,N_11097);
nor U11231 (N_11231,N_11088,N_11183);
and U11232 (N_11232,N_11039,N_11078);
nor U11233 (N_11233,N_11041,N_11180);
nor U11234 (N_11234,N_11188,N_11015);
or U11235 (N_11235,N_11184,N_11114);
or U11236 (N_11236,N_11094,N_11138);
nand U11237 (N_11237,N_11029,N_11021);
or U11238 (N_11238,N_11161,N_11148);
nor U11239 (N_11239,N_11164,N_11066);
and U11240 (N_11240,N_11174,N_11003);
nand U11241 (N_11241,N_11040,N_11042);
xnor U11242 (N_11242,N_11095,N_11163);
and U11243 (N_11243,N_11107,N_11126);
and U11244 (N_11244,N_11198,N_11110);
and U11245 (N_11245,N_11118,N_11010);
and U11246 (N_11246,N_11081,N_11017);
xor U11247 (N_11247,N_11102,N_11159);
or U11248 (N_11248,N_11064,N_11019);
and U11249 (N_11249,N_11069,N_11076);
xnor U11250 (N_11250,N_11199,N_11009);
nand U11251 (N_11251,N_11132,N_11104);
nor U11252 (N_11252,N_11099,N_11173);
nor U11253 (N_11253,N_11053,N_11151);
nor U11254 (N_11254,N_11030,N_11149);
nor U11255 (N_11255,N_11193,N_11155);
nand U11256 (N_11256,N_11033,N_11089);
and U11257 (N_11257,N_11068,N_11135);
nor U11258 (N_11258,N_11082,N_11154);
nor U11259 (N_11259,N_11187,N_11005);
or U11260 (N_11260,N_11070,N_11027);
xnor U11261 (N_11261,N_11045,N_11038);
nor U11262 (N_11262,N_11141,N_11034);
nand U11263 (N_11263,N_11098,N_11096);
and U11264 (N_11264,N_11093,N_11122);
and U11265 (N_11265,N_11013,N_11171);
nor U11266 (N_11266,N_11023,N_11075);
nor U11267 (N_11267,N_11108,N_11169);
and U11268 (N_11268,N_11128,N_11014);
xor U11269 (N_11269,N_11158,N_11192);
nor U11270 (N_11270,N_11006,N_11072);
nand U11271 (N_11271,N_11061,N_11177);
xnor U11272 (N_11272,N_11152,N_11170);
nand U11273 (N_11273,N_11054,N_11051);
nor U11274 (N_11274,N_11123,N_11000);
nand U11275 (N_11275,N_11182,N_11116);
and U11276 (N_11276,N_11056,N_11185);
xnor U11277 (N_11277,N_11153,N_11178);
nor U11278 (N_11278,N_11168,N_11146);
and U11279 (N_11279,N_11189,N_11181);
nand U11280 (N_11280,N_11127,N_11156);
xnor U11281 (N_11281,N_11147,N_11002);
or U11282 (N_11282,N_11179,N_11032);
nand U11283 (N_11283,N_11124,N_11197);
xnor U11284 (N_11284,N_11046,N_11092);
xnor U11285 (N_11285,N_11022,N_11050);
nor U11286 (N_11286,N_11031,N_11166);
or U11287 (N_11287,N_11101,N_11100);
xor U11288 (N_11288,N_11137,N_11125);
xnor U11289 (N_11289,N_11121,N_11079);
xnor U11290 (N_11290,N_11028,N_11090);
nand U11291 (N_11291,N_11109,N_11117);
and U11292 (N_11292,N_11060,N_11129);
and U11293 (N_11293,N_11037,N_11012);
xnor U11294 (N_11294,N_11047,N_11105);
nand U11295 (N_11295,N_11103,N_11133);
or U11296 (N_11296,N_11020,N_11160);
nor U11297 (N_11297,N_11157,N_11007);
and U11298 (N_11298,N_11077,N_11004);
nor U11299 (N_11299,N_11083,N_11085);
and U11300 (N_11300,N_11019,N_11109);
and U11301 (N_11301,N_11111,N_11050);
xor U11302 (N_11302,N_11119,N_11161);
nand U11303 (N_11303,N_11075,N_11174);
xnor U11304 (N_11304,N_11093,N_11170);
xnor U11305 (N_11305,N_11176,N_11158);
nand U11306 (N_11306,N_11059,N_11005);
xnor U11307 (N_11307,N_11042,N_11033);
nand U11308 (N_11308,N_11055,N_11168);
or U11309 (N_11309,N_11159,N_11038);
and U11310 (N_11310,N_11132,N_11032);
nor U11311 (N_11311,N_11176,N_11182);
xnor U11312 (N_11312,N_11171,N_11011);
or U11313 (N_11313,N_11177,N_11016);
or U11314 (N_11314,N_11124,N_11028);
and U11315 (N_11315,N_11092,N_11107);
nand U11316 (N_11316,N_11105,N_11165);
nand U11317 (N_11317,N_11171,N_11023);
and U11318 (N_11318,N_11056,N_11054);
or U11319 (N_11319,N_11157,N_11164);
and U11320 (N_11320,N_11110,N_11179);
or U11321 (N_11321,N_11067,N_11193);
nand U11322 (N_11322,N_11068,N_11049);
or U11323 (N_11323,N_11066,N_11078);
and U11324 (N_11324,N_11138,N_11151);
or U11325 (N_11325,N_11051,N_11104);
nand U11326 (N_11326,N_11112,N_11178);
xor U11327 (N_11327,N_11125,N_11052);
nand U11328 (N_11328,N_11192,N_11105);
nor U11329 (N_11329,N_11050,N_11096);
and U11330 (N_11330,N_11109,N_11099);
xnor U11331 (N_11331,N_11119,N_11109);
and U11332 (N_11332,N_11083,N_11127);
xnor U11333 (N_11333,N_11049,N_11060);
nand U11334 (N_11334,N_11020,N_11105);
nor U11335 (N_11335,N_11048,N_11153);
and U11336 (N_11336,N_11012,N_11071);
or U11337 (N_11337,N_11012,N_11194);
nand U11338 (N_11338,N_11198,N_11022);
xor U11339 (N_11339,N_11076,N_11173);
nand U11340 (N_11340,N_11143,N_11122);
nand U11341 (N_11341,N_11028,N_11052);
nand U11342 (N_11342,N_11084,N_11059);
xor U11343 (N_11343,N_11104,N_11190);
nor U11344 (N_11344,N_11096,N_11048);
and U11345 (N_11345,N_11183,N_11058);
nor U11346 (N_11346,N_11130,N_11159);
nor U11347 (N_11347,N_11132,N_11013);
nor U11348 (N_11348,N_11061,N_11153);
or U11349 (N_11349,N_11140,N_11025);
nand U11350 (N_11350,N_11172,N_11005);
and U11351 (N_11351,N_11097,N_11041);
xnor U11352 (N_11352,N_11058,N_11167);
xnor U11353 (N_11353,N_11132,N_11063);
nand U11354 (N_11354,N_11079,N_11035);
xor U11355 (N_11355,N_11049,N_11003);
or U11356 (N_11356,N_11140,N_11172);
nor U11357 (N_11357,N_11184,N_11187);
and U11358 (N_11358,N_11128,N_11060);
and U11359 (N_11359,N_11117,N_11122);
or U11360 (N_11360,N_11181,N_11163);
and U11361 (N_11361,N_11180,N_11045);
nor U11362 (N_11362,N_11051,N_11155);
xor U11363 (N_11363,N_11113,N_11017);
or U11364 (N_11364,N_11020,N_11192);
nand U11365 (N_11365,N_11168,N_11002);
or U11366 (N_11366,N_11112,N_11051);
or U11367 (N_11367,N_11075,N_11081);
or U11368 (N_11368,N_11145,N_11184);
and U11369 (N_11369,N_11078,N_11044);
and U11370 (N_11370,N_11184,N_11026);
xnor U11371 (N_11371,N_11024,N_11089);
nand U11372 (N_11372,N_11114,N_11088);
xnor U11373 (N_11373,N_11005,N_11134);
and U11374 (N_11374,N_11136,N_11054);
nor U11375 (N_11375,N_11066,N_11012);
and U11376 (N_11376,N_11175,N_11039);
xor U11377 (N_11377,N_11016,N_11022);
nand U11378 (N_11378,N_11169,N_11089);
and U11379 (N_11379,N_11024,N_11088);
or U11380 (N_11380,N_11028,N_11168);
and U11381 (N_11381,N_11065,N_11072);
nor U11382 (N_11382,N_11106,N_11069);
nor U11383 (N_11383,N_11088,N_11180);
and U11384 (N_11384,N_11193,N_11186);
nor U11385 (N_11385,N_11100,N_11149);
or U11386 (N_11386,N_11196,N_11123);
or U11387 (N_11387,N_11035,N_11121);
nand U11388 (N_11388,N_11021,N_11166);
nand U11389 (N_11389,N_11194,N_11148);
nand U11390 (N_11390,N_11073,N_11059);
nand U11391 (N_11391,N_11040,N_11030);
nand U11392 (N_11392,N_11147,N_11104);
nor U11393 (N_11393,N_11096,N_11085);
nor U11394 (N_11394,N_11175,N_11018);
nor U11395 (N_11395,N_11076,N_11009);
and U11396 (N_11396,N_11122,N_11151);
nand U11397 (N_11397,N_11127,N_11011);
nand U11398 (N_11398,N_11058,N_11057);
and U11399 (N_11399,N_11029,N_11068);
or U11400 (N_11400,N_11246,N_11233);
xnor U11401 (N_11401,N_11274,N_11395);
or U11402 (N_11402,N_11371,N_11372);
or U11403 (N_11403,N_11273,N_11250);
nor U11404 (N_11404,N_11379,N_11399);
nor U11405 (N_11405,N_11281,N_11207);
and U11406 (N_11406,N_11334,N_11322);
and U11407 (N_11407,N_11266,N_11307);
and U11408 (N_11408,N_11324,N_11318);
or U11409 (N_11409,N_11361,N_11260);
xnor U11410 (N_11410,N_11350,N_11383);
or U11411 (N_11411,N_11227,N_11277);
or U11412 (N_11412,N_11257,N_11256);
and U11413 (N_11413,N_11289,N_11357);
and U11414 (N_11414,N_11288,N_11231);
xor U11415 (N_11415,N_11373,N_11397);
xor U11416 (N_11416,N_11249,N_11222);
or U11417 (N_11417,N_11314,N_11278);
nor U11418 (N_11418,N_11265,N_11321);
xor U11419 (N_11419,N_11346,N_11224);
xnor U11420 (N_11420,N_11347,N_11242);
and U11421 (N_11421,N_11331,N_11253);
and U11422 (N_11422,N_11287,N_11320);
nand U11423 (N_11423,N_11261,N_11319);
and U11424 (N_11424,N_11218,N_11213);
xor U11425 (N_11425,N_11294,N_11263);
nand U11426 (N_11426,N_11220,N_11272);
nor U11427 (N_11427,N_11367,N_11377);
xor U11428 (N_11428,N_11244,N_11365);
nor U11429 (N_11429,N_11340,N_11228);
and U11430 (N_11430,N_11332,N_11262);
nand U11431 (N_11431,N_11271,N_11363);
nand U11432 (N_11432,N_11300,N_11279);
xor U11433 (N_11433,N_11342,N_11270);
nand U11434 (N_11434,N_11275,N_11386);
nand U11435 (N_11435,N_11339,N_11323);
nand U11436 (N_11436,N_11338,N_11214);
or U11437 (N_11437,N_11312,N_11252);
or U11438 (N_11438,N_11248,N_11204);
xor U11439 (N_11439,N_11304,N_11235);
or U11440 (N_11440,N_11203,N_11223);
xnor U11441 (N_11441,N_11337,N_11391);
or U11442 (N_11442,N_11217,N_11243);
and U11443 (N_11443,N_11335,N_11247);
xor U11444 (N_11444,N_11313,N_11311);
and U11445 (N_11445,N_11251,N_11259);
nand U11446 (N_11446,N_11362,N_11254);
or U11447 (N_11447,N_11286,N_11310);
xor U11448 (N_11448,N_11293,N_11230);
xnor U11449 (N_11449,N_11241,N_11205);
xnor U11450 (N_11450,N_11343,N_11374);
xnor U11451 (N_11451,N_11398,N_11269);
nor U11452 (N_11452,N_11392,N_11353);
or U11453 (N_11453,N_11225,N_11388);
and U11454 (N_11454,N_11341,N_11264);
nor U11455 (N_11455,N_11369,N_11299);
and U11456 (N_11456,N_11325,N_11238);
xnor U11457 (N_11457,N_11351,N_11317);
or U11458 (N_11458,N_11258,N_11326);
or U11459 (N_11459,N_11255,N_11285);
or U11460 (N_11460,N_11236,N_11237);
xnor U11461 (N_11461,N_11229,N_11336);
xnor U11462 (N_11462,N_11328,N_11297);
nor U11463 (N_11463,N_11276,N_11316);
xnor U11464 (N_11464,N_11291,N_11354);
or U11465 (N_11465,N_11267,N_11208);
xor U11466 (N_11466,N_11352,N_11201);
nor U11467 (N_11467,N_11302,N_11368);
xnor U11468 (N_11468,N_11333,N_11348);
nand U11469 (N_11469,N_11327,N_11345);
nand U11470 (N_11470,N_11282,N_11330);
and U11471 (N_11471,N_11370,N_11382);
nor U11472 (N_11472,N_11240,N_11295);
nand U11473 (N_11473,N_11239,N_11303);
nor U11474 (N_11474,N_11280,N_11358);
nor U11475 (N_11475,N_11232,N_11290);
and U11476 (N_11476,N_11283,N_11394);
and U11477 (N_11477,N_11221,N_11298);
and U11478 (N_11478,N_11219,N_11202);
nor U11479 (N_11479,N_11385,N_11349);
xor U11480 (N_11480,N_11364,N_11245);
xnor U11481 (N_11481,N_11200,N_11390);
xor U11482 (N_11482,N_11284,N_11356);
nor U11483 (N_11483,N_11359,N_11215);
nand U11484 (N_11484,N_11216,N_11209);
nand U11485 (N_11485,N_11396,N_11212);
or U11486 (N_11486,N_11381,N_11389);
xor U11487 (N_11487,N_11308,N_11296);
nand U11488 (N_11488,N_11206,N_11306);
nand U11489 (N_11489,N_11355,N_11393);
and U11490 (N_11490,N_11226,N_11292);
or U11491 (N_11491,N_11268,N_11234);
nand U11492 (N_11492,N_11344,N_11210);
nor U11493 (N_11493,N_11387,N_11366);
nand U11494 (N_11494,N_11375,N_11360);
or U11495 (N_11495,N_11378,N_11315);
nand U11496 (N_11496,N_11309,N_11305);
and U11497 (N_11497,N_11329,N_11380);
xor U11498 (N_11498,N_11376,N_11301);
and U11499 (N_11499,N_11384,N_11211);
xnor U11500 (N_11500,N_11399,N_11313);
nand U11501 (N_11501,N_11231,N_11346);
or U11502 (N_11502,N_11316,N_11346);
nand U11503 (N_11503,N_11315,N_11275);
xor U11504 (N_11504,N_11333,N_11202);
xor U11505 (N_11505,N_11247,N_11387);
and U11506 (N_11506,N_11250,N_11213);
xnor U11507 (N_11507,N_11356,N_11216);
nand U11508 (N_11508,N_11252,N_11305);
or U11509 (N_11509,N_11218,N_11368);
nor U11510 (N_11510,N_11297,N_11261);
and U11511 (N_11511,N_11398,N_11379);
nand U11512 (N_11512,N_11372,N_11348);
nor U11513 (N_11513,N_11299,N_11329);
nor U11514 (N_11514,N_11243,N_11358);
nand U11515 (N_11515,N_11305,N_11267);
or U11516 (N_11516,N_11311,N_11252);
or U11517 (N_11517,N_11305,N_11253);
and U11518 (N_11518,N_11309,N_11204);
nand U11519 (N_11519,N_11323,N_11314);
xor U11520 (N_11520,N_11201,N_11223);
and U11521 (N_11521,N_11333,N_11203);
or U11522 (N_11522,N_11238,N_11350);
or U11523 (N_11523,N_11378,N_11397);
or U11524 (N_11524,N_11288,N_11296);
xnor U11525 (N_11525,N_11214,N_11284);
xor U11526 (N_11526,N_11259,N_11350);
xnor U11527 (N_11527,N_11390,N_11342);
or U11528 (N_11528,N_11330,N_11304);
or U11529 (N_11529,N_11227,N_11302);
or U11530 (N_11530,N_11296,N_11272);
nand U11531 (N_11531,N_11326,N_11359);
xor U11532 (N_11532,N_11244,N_11210);
nand U11533 (N_11533,N_11207,N_11338);
and U11534 (N_11534,N_11202,N_11348);
nor U11535 (N_11535,N_11368,N_11360);
and U11536 (N_11536,N_11326,N_11227);
or U11537 (N_11537,N_11277,N_11260);
and U11538 (N_11538,N_11352,N_11234);
nand U11539 (N_11539,N_11288,N_11201);
nand U11540 (N_11540,N_11389,N_11212);
nand U11541 (N_11541,N_11224,N_11394);
and U11542 (N_11542,N_11314,N_11214);
or U11543 (N_11543,N_11361,N_11342);
nor U11544 (N_11544,N_11358,N_11225);
or U11545 (N_11545,N_11294,N_11271);
nand U11546 (N_11546,N_11295,N_11306);
nand U11547 (N_11547,N_11344,N_11375);
xnor U11548 (N_11548,N_11396,N_11334);
nor U11549 (N_11549,N_11352,N_11255);
and U11550 (N_11550,N_11220,N_11244);
or U11551 (N_11551,N_11321,N_11370);
nand U11552 (N_11552,N_11324,N_11355);
or U11553 (N_11553,N_11234,N_11294);
nor U11554 (N_11554,N_11273,N_11366);
nor U11555 (N_11555,N_11349,N_11303);
nor U11556 (N_11556,N_11392,N_11337);
or U11557 (N_11557,N_11324,N_11327);
xor U11558 (N_11558,N_11365,N_11255);
xor U11559 (N_11559,N_11242,N_11269);
xor U11560 (N_11560,N_11278,N_11228);
nor U11561 (N_11561,N_11306,N_11287);
and U11562 (N_11562,N_11328,N_11292);
nand U11563 (N_11563,N_11322,N_11235);
or U11564 (N_11564,N_11381,N_11269);
xor U11565 (N_11565,N_11240,N_11378);
and U11566 (N_11566,N_11285,N_11299);
nor U11567 (N_11567,N_11296,N_11347);
or U11568 (N_11568,N_11300,N_11368);
nand U11569 (N_11569,N_11264,N_11362);
nor U11570 (N_11570,N_11319,N_11347);
or U11571 (N_11571,N_11241,N_11299);
xor U11572 (N_11572,N_11299,N_11286);
xor U11573 (N_11573,N_11344,N_11353);
or U11574 (N_11574,N_11363,N_11280);
nor U11575 (N_11575,N_11289,N_11333);
or U11576 (N_11576,N_11359,N_11396);
nor U11577 (N_11577,N_11249,N_11238);
nand U11578 (N_11578,N_11335,N_11339);
xnor U11579 (N_11579,N_11334,N_11220);
xor U11580 (N_11580,N_11233,N_11391);
and U11581 (N_11581,N_11389,N_11370);
or U11582 (N_11582,N_11206,N_11291);
and U11583 (N_11583,N_11306,N_11272);
xor U11584 (N_11584,N_11228,N_11371);
and U11585 (N_11585,N_11387,N_11265);
nor U11586 (N_11586,N_11253,N_11367);
or U11587 (N_11587,N_11296,N_11321);
nand U11588 (N_11588,N_11282,N_11212);
nand U11589 (N_11589,N_11290,N_11302);
xnor U11590 (N_11590,N_11389,N_11237);
nand U11591 (N_11591,N_11225,N_11359);
nand U11592 (N_11592,N_11314,N_11282);
nor U11593 (N_11593,N_11368,N_11260);
nand U11594 (N_11594,N_11288,N_11208);
nand U11595 (N_11595,N_11308,N_11383);
and U11596 (N_11596,N_11368,N_11315);
or U11597 (N_11597,N_11279,N_11272);
nor U11598 (N_11598,N_11376,N_11246);
nor U11599 (N_11599,N_11329,N_11395);
nor U11600 (N_11600,N_11409,N_11462);
or U11601 (N_11601,N_11598,N_11599);
nand U11602 (N_11602,N_11486,N_11415);
xor U11603 (N_11603,N_11483,N_11445);
nand U11604 (N_11604,N_11494,N_11558);
or U11605 (N_11605,N_11501,N_11427);
nor U11606 (N_11606,N_11560,N_11416);
xor U11607 (N_11607,N_11579,N_11536);
and U11608 (N_11608,N_11520,N_11547);
nor U11609 (N_11609,N_11471,N_11413);
and U11610 (N_11610,N_11472,N_11511);
and U11611 (N_11611,N_11428,N_11402);
nand U11612 (N_11612,N_11479,N_11527);
nor U11613 (N_11613,N_11485,N_11460);
or U11614 (N_11614,N_11593,N_11433);
or U11615 (N_11615,N_11574,N_11597);
or U11616 (N_11616,N_11591,N_11457);
nor U11617 (N_11617,N_11507,N_11468);
xnor U11618 (N_11618,N_11570,N_11466);
nand U11619 (N_11619,N_11498,N_11537);
xor U11620 (N_11620,N_11506,N_11522);
and U11621 (N_11621,N_11510,N_11443);
or U11622 (N_11622,N_11476,N_11513);
and U11623 (N_11623,N_11403,N_11475);
or U11624 (N_11624,N_11590,N_11592);
nor U11625 (N_11625,N_11464,N_11587);
xnor U11626 (N_11626,N_11534,N_11435);
nor U11627 (N_11627,N_11557,N_11474);
xnor U11628 (N_11628,N_11444,N_11477);
nand U11629 (N_11629,N_11407,N_11530);
or U11630 (N_11630,N_11412,N_11432);
xnor U11631 (N_11631,N_11481,N_11493);
nand U11632 (N_11632,N_11441,N_11482);
and U11633 (N_11633,N_11561,N_11496);
nor U11634 (N_11634,N_11401,N_11567);
nor U11635 (N_11635,N_11491,N_11436);
nand U11636 (N_11636,N_11449,N_11518);
nor U11637 (N_11637,N_11526,N_11509);
nand U11638 (N_11638,N_11411,N_11455);
and U11639 (N_11639,N_11495,N_11552);
or U11640 (N_11640,N_11529,N_11422);
xnor U11641 (N_11641,N_11596,N_11538);
nand U11642 (N_11642,N_11434,N_11430);
nor U11643 (N_11643,N_11431,N_11404);
nand U11644 (N_11644,N_11577,N_11488);
nor U11645 (N_11645,N_11531,N_11420);
xor U11646 (N_11646,N_11517,N_11480);
nand U11647 (N_11647,N_11400,N_11408);
nand U11648 (N_11648,N_11571,N_11446);
and U11649 (N_11649,N_11546,N_11542);
xor U11650 (N_11650,N_11572,N_11437);
nor U11651 (N_11651,N_11463,N_11539);
nand U11652 (N_11652,N_11424,N_11580);
xnor U11653 (N_11653,N_11421,N_11540);
nor U11654 (N_11654,N_11500,N_11550);
or U11655 (N_11655,N_11499,N_11418);
or U11656 (N_11656,N_11512,N_11502);
or U11657 (N_11657,N_11514,N_11442);
or U11658 (N_11658,N_11452,N_11467);
xnor U11659 (N_11659,N_11548,N_11521);
or U11660 (N_11660,N_11556,N_11516);
and U11661 (N_11661,N_11559,N_11564);
nor U11662 (N_11662,N_11575,N_11583);
nand U11663 (N_11663,N_11523,N_11489);
or U11664 (N_11664,N_11525,N_11528);
nand U11665 (N_11665,N_11419,N_11470);
nand U11666 (N_11666,N_11508,N_11519);
nand U11667 (N_11667,N_11448,N_11456);
xnor U11668 (N_11668,N_11497,N_11544);
or U11669 (N_11669,N_11532,N_11533);
nand U11670 (N_11670,N_11565,N_11562);
and U11671 (N_11671,N_11504,N_11505);
nor U11672 (N_11672,N_11405,N_11586);
or U11673 (N_11673,N_11425,N_11429);
or U11674 (N_11674,N_11503,N_11582);
nand U11675 (N_11675,N_11459,N_11535);
or U11676 (N_11676,N_11554,N_11568);
and U11677 (N_11677,N_11524,N_11541);
nor U11678 (N_11678,N_11589,N_11439);
nand U11679 (N_11679,N_11543,N_11585);
xor U11680 (N_11680,N_11569,N_11490);
nor U11681 (N_11681,N_11453,N_11545);
nand U11682 (N_11682,N_11555,N_11581);
and U11683 (N_11683,N_11473,N_11595);
and U11684 (N_11684,N_11576,N_11484);
nand U11685 (N_11685,N_11515,N_11438);
nand U11686 (N_11686,N_11414,N_11440);
or U11687 (N_11687,N_11551,N_11465);
nor U11688 (N_11688,N_11454,N_11487);
nor U11689 (N_11689,N_11423,N_11588);
and U11690 (N_11690,N_11450,N_11563);
and U11691 (N_11691,N_11451,N_11553);
xnor U11692 (N_11692,N_11417,N_11406);
and U11693 (N_11693,N_11447,N_11458);
and U11694 (N_11694,N_11469,N_11584);
nor U11695 (N_11695,N_11578,N_11478);
nand U11696 (N_11696,N_11426,N_11410);
nand U11697 (N_11697,N_11573,N_11566);
xnor U11698 (N_11698,N_11549,N_11492);
nor U11699 (N_11699,N_11461,N_11594);
nand U11700 (N_11700,N_11591,N_11481);
nand U11701 (N_11701,N_11435,N_11541);
nand U11702 (N_11702,N_11597,N_11418);
xor U11703 (N_11703,N_11522,N_11433);
xor U11704 (N_11704,N_11440,N_11509);
xor U11705 (N_11705,N_11501,N_11459);
or U11706 (N_11706,N_11419,N_11479);
or U11707 (N_11707,N_11502,N_11473);
nor U11708 (N_11708,N_11528,N_11418);
or U11709 (N_11709,N_11594,N_11555);
and U11710 (N_11710,N_11586,N_11408);
xnor U11711 (N_11711,N_11594,N_11543);
and U11712 (N_11712,N_11420,N_11407);
xor U11713 (N_11713,N_11400,N_11532);
and U11714 (N_11714,N_11452,N_11415);
nand U11715 (N_11715,N_11474,N_11565);
and U11716 (N_11716,N_11529,N_11534);
nand U11717 (N_11717,N_11575,N_11513);
or U11718 (N_11718,N_11495,N_11437);
or U11719 (N_11719,N_11575,N_11455);
and U11720 (N_11720,N_11515,N_11504);
nand U11721 (N_11721,N_11516,N_11524);
nor U11722 (N_11722,N_11484,N_11413);
nand U11723 (N_11723,N_11568,N_11518);
nand U11724 (N_11724,N_11576,N_11441);
or U11725 (N_11725,N_11491,N_11440);
nor U11726 (N_11726,N_11535,N_11409);
xnor U11727 (N_11727,N_11429,N_11434);
xor U11728 (N_11728,N_11507,N_11533);
nor U11729 (N_11729,N_11451,N_11496);
and U11730 (N_11730,N_11525,N_11428);
and U11731 (N_11731,N_11401,N_11579);
or U11732 (N_11732,N_11500,N_11461);
nand U11733 (N_11733,N_11584,N_11476);
xnor U11734 (N_11734,N_11535,N_11405);
nand U11735 (N_11735,N_11599,N_11424);
and U11736 (N_11736,N_11421,N_11409);
nor U11737 (N_11737,N_11425,N_11407);
nor U11738 (N_11738,N_11568,N_11403);
nand U11739 (N_11739,N_11413,N_11406);
nor U11740 (N_11740,N_11511,N_11412);
nor U11741 (N_11741,N_11487,N_11549);
and U11742 (N_11742,N_11435,N_11470);
or U11743 (N_11743,N_11561,N_11455);
or U11744 (N_11744,N_11478,N_11590);
nor U11745 (N_11745,N_11594,N_11435);
and U11746 (N_11746,N_11580,N_11462);
nand U11747 (N_11747,N_11585,N_11404);
and U11748 (N_11748,N_11586,N_11480);
nor U11749 (N_11749,N_11596,N_11421);
xor U11750 (N_11750,N_11451,N_11576);
xor U11751 (N_11751,N_11513,N_11483);
xor U11752 (N_11752,N_11574,N_11532);
or U11753 (N_11753,N_11518,N_11402);
and U11754 (N_11754,N_11534,N_11491);
and U11755 (N_11755,N_11537,N_11552);
or U11756 (N_11756,N_11561,N_11492);
nor U11757 (N_11757,N_11470,N_11429);
or U11758 (N_11758,N_11458,N_11547);
and U11759 (N_11759,N_11529,N_11502);
nor U11760 (N_11760,N_11479,N_11556);
and U11761 (N_11761,N_11453,N_11480);
or U11762 (N_11762,N_11522,N_11577);
nor U11763 (N_11763,N_11449,N_11493);
nand U11764 (N_11764,N_11432,N_11596);
nor U11765 (N_11765,N_11537,N_11517);
xnor U11766 (N_11766,N_11499,N_11408);
nand U11767 (N_11767,N_11497,N_11446);
and U11768 (N_11768,N_11451,N_11498);
nand U11769 (N_11769,N_11487,N_11497);
or U11770 (N_11770,N_11504,N_11457);
and U11771 (N_11771,N_11469,N_11535);
and U11772 (N_11772,N_11413,N_11462);
and U11773 (N_11773,N_11433,N_11474);
or U11774 (N_11774,N_11531,N_11577);
nand U11775 (N_11775,N_11586,N_11460);
nor U11776 (N_11776,N_11582,N_11430);
xnor U11777 (N_11777,N_11581,N_11409);
nor U11778 (N_11778,N_11565,N_11459);
or U11779 (N_11779,N_11434,N_11505);
or U11780 (N_11780,N_11463,N_11429);
nand U11781 (N_11781,N_11591,N_11461);
nand U11782 (N_11782,N_11553,N_11506);
nor U11783 (N_11783,N_11416,N_11546);
nor U11784 (N_11784,N_11460,N_11570);
nand U11785 (N_11785,N_11582,N_11424);
nand U11786 (N_11786,N_11507,N_11495);
or U11787 (N_11787,N_11557,N_11493);
nand U11788 (N_11788,N_11453,N_11500);
nand U11789 (N_11789,N_11436,N_11505);
nand U11790 (N_11790,N_11445,N_11546);
nand U11791 (N_11791,N_11450,N_11467);
nand U11792 (N_11792,N_11568,N_11422);
nor U11793 (N_11793,N_11403,N_11439);
xor U11794 (N_11794,N_11400,N_11471);
nand U11795 (N_11795,N_11423,N_11473);
or U11796 (N_11796,N_11406,N_11565);
and U11797 (N_11797,N_11534,N_11593);
and U11798 (N_11798,N_11450,N_11591);
nor U11799 (N_11799,N_11548,N_11529);
and U11800 (N_11800,N_11745,N_11679);
or U11801 (N_11801,N_11614,N_11608);
and U11802 (N_11802,N_11644,N_11600);
or U11803 (N_11803,N_11624,N_11754);
and U11804 (N_11804,N_11619,N_11674);
nor U11805 (N_11805,N_11687,N_11752);
nand U11806 (N_11806,N_11796,N_11657);
nand U11807 (N_11807,N_11723,N_11669);
and U11808 (N_11808,N_11791,N_11743);
nor U11809 (N_11809,N_11736,N_11797);
or U11810 (N_11810,N_11622,N_11615);
xor U11811 (N_11811,N_11756,N_11768);
and U11812 (N_11812,N_11747,N_11704);
nand U11813 (N_11813,N_11713,N_11604);
and U11814 (N_11814,N_11758,N_11675);
nor U11815 (N_11815,N_11610,N_11786);
nor U11816 (N_11816,N_11741,N_11770);
nor U11817 (N_11817,N_11711,N_11715);
nor U11818 (N_11818,N_11783,N_11649);
and U11819 (N_11819,N_11737,N_11774);
or U11820 (N_11820,N_11682,N_11673);
nor U11821 (N_11821,N_11751,N_11706);
xor U11822 (N_11822,N_11638,N_11647);
nor U11823 (N_11823,N_11683,N_11779);
nor U11824 (N_11824,N_11760,N_11650);
nand U11825 (N_11825,N_11661,N_11701);
or U11826 (N_11826,N_11761,N_11660);
and U11827 (N_11827,N_11666,N_11696);
or U11828 (N_11828,N_11708,N_11616);
xnor U11829 (N_11829,N_11694,N_11668);
and U11830 (N_11830,N_11705,N_11628);
xnor U11831 (N_11831,N_11606,N_11629);
nand U11832 (N_11832,N_11671,N_11625);
nand U11833 (N_11833,N_11798,N_11734);
and U11834 (N_11834,N_11688,N_11690);
nand U11835 (N_11835,N_11775,N_11709);
nand U11836 (N_11836,N_11794,N_11746);
or U11837 (N_11837,N_11722,N_11612);
nand U11838 (N_11838,N_11635,N_11654);
nand U11839 (N_11839,N_11698,N_11678);
or U11840 (N_11840,N_11670,N_11738);
and U11841 (N_11841,N_11702,N_11697);
nor U11842 (N_11842,N_11700,N_11740);
nor U11843 (N_11843,N_11727,N_11633);
xor U11844 (N_11844,N_11648,N_11640);
and U11845 (N_11845,N_11781,N_11658);
nand U11846 (N_11846,N_11699,N_11630);
nor U11847 (N_11847,N_11602,N_11714);
xnor U11848 (N_11848,N_11773,N_11776);
nor U11849 (N_11849,N_11632,N_11641);
or U11850 (N_11850,N_11686,N_11643);
xor U11851 (N_11851,N_11601,N_11636);
xor U11852 (N_11852,N_11677,N_11655);
and U11853 (N_11853,N_11787,N_11642);
or U11854 (N_11854,N_11607,N_11603);
or U11855 (N_11855,N_11665,N_11739);
xnor U11856 (N_11856,N_11672,N_11695);
nor U11857 (N_11857,N_11712,N_11605);
xor U11858 (N_11858,N_11778,N_11728);
and U11859 (N_11859,N_11692,N_11731);
xnor U11860 (N_11860,N_11680,N_11609);
and U11861 (N_11861,N_11716,N_11719);
xor U11862 (N_11862,N_11639,N_11691);
nor U11863 (N_11863,N_11784,N_11748);
nand U11864 (N_11864,N_11762,N_11676);
nand U11865 (N_11865,N_11710,N_11730);
nand U11866 (N_11866,N_11656,N_11732);
or U11867 (N_11867,N_11763,N_11617);
nor U11868 (N_11868,N_11788,N_11721);
nand U11869 (N_11869,N_11651,N_11765);
nor U11870 (N_11870,N_11689,N_11667);
nand U11871 (N_11871,N_11742,N_11664);
xnor U11872 (N_11872,N_11753,N_11693);
xnor U11873 (N_11873,N_11634,N_11718);
xor U11874 (N_11874,N_11744,N_11652);
and U11875 (N_11875,N_11749,N_11618);
or U11876 (N_11876,N_11685,N_11725);
and U11877 (N_11877,N_11626,N_11720);
and U11878 (N_11878,N_11759,N_11793);
xor U11879 (N_11879,N_11659,N_11646);
and U11880 (N_11880,N_11799,N_11611);
or U11881 (N_11881,N_11792,N_11662);
nor U11882 (N_11882,N_11750,N_11767);
xnor U11883 (N_11883,N_11627,N_11703);
nand U11884 (N_11884,N_11733,N_11790);
nand U11885 (N_11885,N_11620,N_11735);
xnor U11886 (N_11886,N_11755,N_11684);
nand U11887 (N_11887,N_11769,N_11795);
and U11888 (N_11888,N_11785,N_11764);
and U11889 (N_11889,N_11777,N_11707);
nand U11890 (N_11890,N_11757,N_11653);
or U11891 (N_11891,N_11726,N_11717);
xor U11892 (N_11892,N_11772,N_11729);
nand U11893 (N_11893,N_11645,N_11766);
nand U11894 (N_11894,N_11637,N_11771);
or U11895 (N_11895,N_11789,N_11663);
nor U11896 (N_11896,N_11724,N_11681);
and U11897 (N_11897,N_11780,N_11631);
and U11898 (N_11898,N_11613,N_11623);
nand U11899 (N_11899,N_11621,N_11782);
nand U11900 (N_11900,N_11671,N_11715);
or U11901 (N_11901,N_11716,N_11792);
xnor U11902 (N_11902,N_11724,N_11668);
xor U11903 (N_11903,N_11722,N_11791);
nand U11904 (N_11904,N_11745,N_11643);
and U11905 (N_11905,N_11622,N_11679);
and U11906 (N_11906,N_11620,N_11722);
or U11907 (N_11907,N_11776,N_11638);
and U11908 (N_11908,N_11674,N_11782);
xnor U11909 (N_11909,N_11655,N_11795);
xnor U11910 (N_11910,N_11660,N_11764);
and U11911 (N_11911,N_11611,N_11784);
nor U11912 (N_11912,N_11669,N_11749);
nor U11913 (N_11913,N_11768,N_11685);
xnor U11914 (N_11914,N_11631,N_11744);
nor U11915 (N_11915,N_11658,N_11652);
or U11916 (N_11916,N_11756,N_11623);
and U11917 (N_11917,N_11708,N_11676);
and U11918 (N_11918,N_11714,N_11724);
nand U11919 (N_11919,N_11676,N_11740);
and U11920 (N_11920,N_11774,N_11663);
nor U11921 (N_11921,N_11645,N_11794);
nor U11922 (N_11922,N_11731,N_11646);
nor U11923 (N_11923,N_11749,N_11754);
nand U11924 (N_11924,N_11648,N_11701);
nand U11925 (N_11925,N_11680,N_11613);
or U11926 (N_11926,N_11698,N_11641);
and U11927 (N_11927,N_11685,N_11646);
nor U11928 (N_11928,N_11641,N_11677);
xnor U11929 (N_11929,N_11792,N_11636);
and U11930 (N_11930,N_11774,N_11729);
nor U11931 (N_11931,N_11787,N_11608);
and U11932 (N_11932,N_11618,N_11745);
xnor U11933 (N_11933,N_11784,N_11793);
nand U11934 (N_11934,N_11785,N_11760);
nor U11935 (N_11935,N_11716,N_11763);
or U11936 (N_11936,N_11736,N_11684);
nand U11937 (N_11937,N_11787,N_11760);
or U11938 (N_11938,N_11636,N_11652);
nor U11939 (N_11939,N_11645,N_11730);
or U11940 (N_11940,N_11756,N_11698);
or U11941 (N_11941,N_11722,N_11688);
xor U11942 (N_11942,N_11655,N_11696);
and U11943 (N_11943,N_11744,N_11794);
xnor U11944 (N_11944,N_11763,N_11771);
nand U11945 (N_11945,N_11685,N_11651);
or U11946 (N_11946,N_11670,N_11613);
and U11947 (N_11947,N_11776,N_11758);
xnor U11948 (N_11948,N_11729,N_11699);
xnor U11949 (N_11949,N_11713,N_11637);
nor U11950 (N_11950,N_11710,N_11793);
nor U11951 (N_11951,N_11695,N_11701);
nand U11952 (N_11952,N_11740,N_11697);
nand U11953 (N_11953,N_11619,N_11683);
nand U11954 (N_11954,N_11600,N_11679);
and U11955 (N_11955,N_11686,N_11797);
nand U11956 (N_11956,N_11666,N_11603);
xor U11957 (N_11957,N_11703,N_11774);
or U11958 (N_11958,N_11643,N_11665);
or U11959 (N_11959,N_11722,N_11647);
and U11960 (N_11960,N_11668,N_11675);
and U11961 (N_11961,N_11792,N_11785);
or U11962 (N_11962,N_11684,N_11774);
or U11963 (N_11963,N_11671,N_11676);
and U11964 (N_11964,N_11795,N_11626);
nor U11965 (N_11965,N_11690,N_11602);
nand U11966 (N_11966,N_11771,N_11741);
or U11967 (N_11967,N_11747,N_11675);
xnor U11968 (N_11968,N_11798,N_11677);
or U11969 (N_11969,N_11609,N_11625);
or U11970 (N_11970,N_11685,N_11760);
nand U11971 (N_11971,N_11721,N_11706);
nand U11972 (N_11972,N_11639,N_11671);
and U11973 (N_11973,N_11739,N_11754);
xor U11974 (N_11974,N_11647,N_11603);
or U11975 (N_11975,N_11765,N_11666);
xnor U11976 (N_11976,N_11719,N_11674);
xnor U11977 (N_11977,N_11622,N_11791);
nor U11978 (N_11978,N_11607,N_11775);
xor U11979 (N_11979,N_11653,N_11692);
nand U11980 (N_11980,N_11657,N_11649);
nand U11981 (N_11981,N_11751,N_11741);
nand U11982 (N_11982,N_11782,N_11791);
nor U11983 (N_11983,N_11683,N_11776);
xor U11984 (N_11984,N_11666,N_11625);
nor U11985 (N_11985,N_11615,N_11663);
xnor U11986 (N_11986,N_11661,N_11615);
xnor U11987 (N_11987,N_11706,N_11679);
and U11988 (N_11988,N_11723,N_11789);
xnor U11989 (N_11989,N_11671,N_11774);
or U11990 (N_11990,N_11678,N_11676);
and U11991 (N_11991,N_11759,N_11603);
nor U11992 (N_11992,N_11737,N_11730);
nor U11993 (N_11993,N_11657,N_11788);
nand U11994 (N_11994,N_11758,N_11723);
nor U11995 (N_11995,N_11609,N_11701);
nor U11996 (N_11996,N_11669,N_11764);
xnor U11997 (N_11997,N_11721,N_11739);
nor U11998 (N_11998,N_11785,N_11663);
xnor U11999 (N_11999,N_11783,N_11704);
nor U12000 (N_12000,N_11919,N_11976);
nand U12001 (N_12001,N_11817,N_11932);
and U12002 (N_12002,N_11814,N_11887);
xor U12003 (N_12003,N_11890,N_11861);
nand U12004 (N_12004,N_11869,N_11842);
nor U12005 (N_12005,N_11974,N_11922);
xnor U12006 (N_12006,N_11859,N_11993);
xnor U12007 (N_12007,N_11882,N_11809);
and U12008 (N_12008,N_11991,N_11871);
nand U12009 (N_12009,N_11850,N_11896);
and U12010 (N_12010,N_11826,N_11881);
or U12011 (N_12011,N_11940,N_11969);
and U12012 (N_12012,N_11962,N_11885);
nor U12013 (N_12013,N_11944,N_11840);
nor U12014 (N_12014,N_11845,N_11879);
or U12015 (N_12015,N_11893,N_11989);
nand U12016 (N_12016,N_11916,N_11996);
or U12017 (N_12017,N_11992,N_11823);
xor U12018 (N_12018,N_11824,N_11910);
or U12019 (N_12019,N_11836,N_11956);
nand U12020 (N_12020,N_11902,N_11906);
xor U12021 (N_12021,N_11930,N_11883);
nand U12022 (N_12022,N_11874,N_11977);
xor U12023 (N_12023,N_11866,N_11806);
nand U12024 (N_12024,N_11920,N_11983);
or U12025 (N_12025,N_11827,N_11918);
xnor U12026 (N_12026,N_11863,N_11844);
or U12027 (N_12027,N_11815,N_11851);
or U12028 (N_12028,N_11876,N_11958);
xnor U12029 (N_12029,N_11897,N_11973);
xor U12030 (N_12030,N_11888,N_11904);
xnor U12031 (N_12031,N_11868,N_11858);
nand U12032 (N_12032,N_11835,N_11936);
nor U12033 (N_12033,N_11848,N_11975);
nand U12034 (N_12034,N_11963,N_11926);
nand U12035 (N_12035,N_11872,N_11984);
or U12036 (N_12036,N_11935,N_11933);
nor U12037 (N_12037,N_11901,N_11857);
xor U12038 (N_12038,N_11924,N_11854);
nand U12039 (N_12039,N_11966,N_11834);
nor U12040 (N_12040,N_11998,N_11913);
or U12041 (N_12041,N_11898,N_11947);
nand U12042 (N_12042,N_11931,N_11949);
or U12043 (N_12043,N_11838,N_11855);
and U12044 (N_12044,N_11945,N_11877);
xnor U12045 (N_12045,N_11929,N_11982);
or U12046 (N_12046,N_11960,N_11968);
nand U12047 (N_12047,N_11899,N_11829);
nand U12048 (N_12048,N_11997,N_11964);
and U12049 (N_12049,N_11911,N_11959);
and U12050 (N_12050,N_11865,N_11816);
nor U12051 (N_12051,N_11884,N_11828);
and U12052 (N_12052,N_11811,N_11875);
xnor U12053 (N_12053,N_11803,N_11923);
or U12054 (N_12054,N_11800,N_11946);
nand U12055 (N_12055,N_11941,N_11886);
nor U12056 (N_12056,N_11937,N_11812);
nand U12057 (N_12057,N_11927,N_11833);
xnor U12058 (N_12058,N_11917,N_11953);
or U12059 (N_12059,N_11986,N_11900);
or U12060 (N_12060,N_11810,N_11909);
or U12061 (N_12061,N_11950,N_11954);
xnor U12062 (N_12062,N_11971,N_11988);
xor U12063 (N_12063,N_11908,N_11807);
and U12064 (N_12064,N_11832,N_11939);
or U12065 (N_12065,N_11980,N_11951);
xor U12066 (N_12066,N_11860,N_11818);
or U12067 (N_12067,N_11938,N_11849);
xnor U12068 (N_12068,N_11928,N_11813);
xor U12069 (N_12069,N_11819,N_11914);
xor U12070 (N_12070,N_11805,N_11802);
xor U12071 (N_12071,N_11952,N_11990);
and U12072 (N_12072,N_11948,N_11999);
nor U12073 (N_12073,N_11943,N_11979);
nor U12074 (N_12074,N_11965,N_11873);
or U12075 (N_12075,N_11862,N_11915);
xnor U12076 (N_12076,N_11870,N_11970);
and U12077 (N_12077,N_11895,N_11894);
and U12078 (N_12078,N_11987,N_11921);
nor U12079 (N_12079,N_11942,N_11825);
and U12080 (N_12080,N_11837,N_11892);
xor U12081 (N_12081,N_11912,N_11955);
and U12082 (N_12082,N_11907,N_11903);
and U12083 (N_12083,N_11808,N_11841);
or U12084 (N_12084,N_11853,N_11831);
or U12085 (N_12085,N_11852,N_11843);
and U12086 (N_12086,N_11889,N_11847);
xor U12087 (N_12087,N_11856,N_11801);
nand U12088 (N_12088,N_11957,N_11994);
or U12089 (N_12089,N_11822,N_11978);
nor U12090 (N_12090,N_11905,N_11985);
xnor U12091 (N_12091,N_11867,N_11804);
xnor U12092 (N_12092,N_11972,N_11846);
or U12093 (N_12093,N_11880,N_11821);
and U12094 (N_12094,N_11864,N_11878);
or U12095 (N_12095,N_11981,N_11830);
nor U12096 (N_12096,N_11967,N_11820);
and U12097 (N_12097,N_11891,N_11934);
or U12098 (N_12098,N_11925,N_11961);
nor U12099 (N_12099,N_11839,N_11995);
xor U12100 (N_12100,N_11947,N_11812);
or U12101 (N_12101,N_11812,N_11896);
nand U12102 (N_12102,N_11892,N_11858);
and U12103 (N_12103,N_11988,N_11901);
nor U12104 (N_12104,N_11933,N_11928);
or U12105 (N_12105,N_11902,N_11882);
or U12106 (N_12106,N_11907,N_11967);
nor U12107 (N_12107,N_11899,N_11862);
nor U12108 (N_12108,N_11958,N_11916);
and U12109 (N_12109,N_11936,N_11997);
and U12110 (N_12110,N_11990,N_11933);
or U12111 (N_12111,N_11847,N_11815);
and U12112 (N_12112,N_11923,N_11890);
nor U12113 (N_12113,N_11907,N_11943);
or U12114 (N_12114,N_11821,N_11889);
xnor U12115 (N_12115,N_11838,N_11983);
nor U12116 (N_12116,N_11987,N_11853);
nor U12117 (N_12117,N_11880,N_11986);
and U12118 (N_12118,N_11979,N_11921);
or U12119 (N_12119,N_11871,N_11886);
xor U12120 (N_12120,N_11815,N_11864);
or U12121 (N_12121,N_11987,N_11882);
xor U12122 (N_12122,N_11945,N_11888);
nor U12123 (N_12123,N_11938,N_11851);
or U12124 (N_12124,N_11899,N_11910);
and U12125 (N_12125,N_11992,N_11863);
nor U12126 (N_12126,N_11907,N_11911);
xor U12127 (N_12127,N_11986,N_11874);
or U12128 (N_12128,N_11918,N_11983);
nor U12129 (N_12129,N_11848,N_11881);
or U12130 (N_12130,N_11885,N_11956);
nor U12131 (N_12131,N_11831,N_11817);
or U12132 (N_12132,N_11958,N_11882);
nand U12133 (N_12133,N_11827,N_11963);
and U12134 (N_12134,N_11991,N_11839);
nand U12135 (N_12135,N_11980,N_11861);
and U12136 (N_12136,N_11978,N_11999);
xor U12137 (N_12137,N_11892,N_11832);
nand U12138 (N_12138,N_11988,N_11869);
nand U12139 (N_12139,N_11924,N_11842);
nor U12140 (N_12140,N_11825,N_11995);
nor U12141 (N_12141,N_11985,N_11894);
nand U12142 (N_12142,N_11881,N_11829);
nor U12143 (N_12143,N_11997,N_11916);
xor U12144 (N_12144,N_11956,N_11939);
xnor U12145 (N_12145,N_11839,N_11974);
or U12146 (N_12146,N_11991,N_11992);
nor U12147 (N_12147,N_11855,N_11909);
or U12148 (N_12148,N_11965,N_11897);
nor U12149 (N_12149,N_11838,N_11843);
or U12150 (N_12150,N_11903,N_11977);
xnor U12151 (N_12151,N_11844,N_11952);
nor U12152 (N_12152,N_11939,N_11819);
and U12153 (N_12153,N_11852,N_11989);
nand U12154 (N_12154,N_11853,N_11819);
or U12155 (N_12155,N_11819,N_11847);
nand U12156 (N_12156,N_11956,N_11811);
and U12157 (N_12157,N_11906,N_11871);
xor U12158 (N_12158,N_11905,N_11822);
nand U12159 (N_12159,N_11806,N_11865);
nand U12160 (N_12160,N_11993,N_11832);
nand U12161 (N_12161,N_11977,N_11800);
and U12162 (N_12162,N_11804,N_11895);
xor U12163 (N_12163,N_11882,N_11984);
xor U12164 (N_12164,N_11943,N_11830);
and U12165 (N_12165,N_11853,N_11989);
xor U12166 (N_12166,N_11833,N_11828);
nand U12167 (N_12167,N_11943,N_11928);
nor U12168 (N_12168,N_11936,N_11804);
xnor U12169 (N_12169,N_11923,N_11992);
nor U12170 (N_12170,N_11928,N_11996);
nand U12171 (N_12171,N_11847,N_11904);
nand U12172 (N_12172,N_11905,N_11874);
xnor U12173 (N_12173,N_11917,N_11938);
nor U12174 (N_12174,N_11964,N_11947);
nand U12175 (N_12175,N_11840,N_11803);
xnor U12176 (N_12176,N_11953,N_11971);
and U12177 (N_12177,N_11882,N_11859);
nand U12178 (N_12178,N_11966,N_11938);
nand U12179 (N_12179,N_11850,N_11855);
nor U12180 (N_12180,N_11872,N_11956);
nor U12181 (N_12181,N_11899,N_11941);
nor U12182 (N_12182,N_11997,N_11861);
nand U12183 (N_12183,N_11865,N_11938);
and U12184 (N_12184,N_11878,N_11977);
or U12185 (N_12185,N_11960,N_11851);
or U12186 (N_12186,N_11848,N_11870);
and U12187 (N_12187,N_11800,N_11912);
nand U12188 (N_12188,N_11881,N_11992);
nor U12189 (N_12189,N_11910,N_11986);
nor U12190 (N_12190,N_11929,N_11856);
nand U12191 (N_12191,N_11922,N_11890);
nand U12192 (N_12192,N_11982,N_11881);
nor U12193 (N_12193,N_11992,N_11906);
nor U12194 (N_12194,N_11833,N_11917);
and U12195 (N_12195,N_11821,N_11979);
and U12196 (N_12196,N_11995,N_11871);
and U12197 (N_12197,N_11991,N_11862);
or U12198 (N_12198,N_11805,N_11814);
nand U12199 (N_12199,N_11983,N_11882);
nand U12200 (N_12200,N_12154,N_12145);
and U12201 (N_12201,N_12074,N_12064);
xnor U12202 (N_12202,N_12148,N_12161);
nor U12203 (N_12203,N_12030,N_12037);
nor U12204 (N_12204,N_12114,N_12071);
nor U12205 (N_12205,N_12091,N_12076);
nand U12206 (N_12206,N_12118,N_12149);
nor U12207 (N_12207,N_12178,N_12124);
xor U12208 (N_12208,N_12199,N_12164);
nor U12209 (N_12209,N_12077,N_12029);
or U12210 (N_12210,N_12107,N_12159);
nand U12211 (N_12211,N_12086,N_12033);
nor U12212 (N_12212,N_12050,N_12186);
xnor U12213 (N_12213,N_12051,N_12111);
xor U12214 (N_12214,N_12014,N_12015);
and U12215 (N_12215,N_12026,N_12194);
nor U12216 (N_12216,N_12005,N_12185);
or U12217 (N_12217,N_12122,N_12165);
and U12218 (N_12218,N_12106,N_12063);
nor U12219 (N_12219,N_12075,N_12098);
and U12220 (N_12220,N_12053,N_12127);
or U12221 (N_12221,N_12132,N_12072);
and U12222 (N_12222,N_12141,N_12073);
xnor U12223 (N_12223,N_12142,N_12174);
nand U12224 (N_12224,N_12129,N_12057);
and U12225 (N_12225,N_12179,N_12061);
nand U12226 (N_12226,N_12019,N_12109);
or U12227 (N_12227,N_12020,N_12192);
xor U12228 (N_12228,N_12018,N_12001);
xor U12229 (N_12229,N_12160,N_12130);
and U12230 (N_12230,N_12045,N_12102);
or U12231 (N_12231,N_12042,N_12139);
nor U12232 (N_12232,N_12172,N_12044);
and U12233 (N_12233,N_12092,N_12134);
nand U12234 (N_12234,N_12166,N_12152);
nand U12235 (N_12235,N_12125,N_12023);
nand U12236 (N_12236,N_12188,N_12126);
nand U12237 (N_12237,N_12116,N_12197);
nand U12238 (N_12238,N_12082,N_12183);
xor U12239 (N_12239,N_12080,N_12101);
xor U12240 (N_12240,N_12151,N_12085);
or U12241 (N_12241,N_12083,N_12024);
nor U12242 (N_12242,N_12198,N_12059);
or U12243 (N_12243,N_12120,N_12052);
xnor U12244 (N_12244,N_12117,N_12003);
and U12245 (N_12245,N_12039,N_12090);
or U12246 (N_12246,N_12121,N_12137);
nor U12247 (N_12247,N_12147,N_12135);
nor U12248 (N_12248,N_12171,N_12004);
or U12249 (N_12249,N_12055,N_12175);
nand U12250 (N_12250,N_12177,N_12079);
nand U12251 (N_12251,N_12190,N_12123);
or U12252 (N_12252,N_12038,N_12084);
or U12253 (N_12253,N_12058,N_12108);
and U12254 (N_12254,N_12105,N_12195);
or U12255 (N_12255,N_12047,N_12028);
and U12256 (N_12256,N_12062,N_12155);
nand U12257 (N_12257,N_12009,N_12022);
and U12258 (N_12258,N_12131,N_12115);
and U12259 (N_12259,N_12078,N_12007);
nand U12260 (N_12260,N_12008,N_12000);
xnor U12261 (N_12261,N_12002,N_12182);
nand U12262 (N_12262,N_12017,N_12021);
nand U12263 (N_12263,N_12043,N_12140);
nor U12264 (N_12264,N_12087,N_12070);
nor U12265 (N_12265,N_12133,N_12191);
or U12266 (N_12266,N_12184,N_12093);
xnor U12267 (N_12267,N_12136,N_12013);
nor U12268 (N_12268,N_12040,N_12112);
nor U12269 (N_12269,N_12167,N_12049);
nand U12270 (N_12270,N_12025,N_12156);
and U12271 (N_12271,N_12067,N_12187);
xor U12272 (N_12272,N_12035,N_12065);
xor U12273 (N_12273,N_12060,N_12056);
xor U12274 (N_12274,N_12034,N_12069);
or U12275 (N_12275,N_12012,N_12068);
or U12276 (N_12276,N_12146,N_12168);
and U12277 (N_12277,N_12110,N_12010);
xor U12278 (N_12278,N_12031,N_12094);
and U12279 (N_12279,N_12153,N_12176);
or U12280 (N_12280,N_12181,N_12099);
or U12281 (N_12281,N_12097,N_12150);
and U12282 (N_12282,N_12081,N_12143);
nand U12283 (N_12283,N_12144,N_12027);
and U12284 (N_12284,N_12157,N_12100);
xor U12285 (N_12285,N_12103,N_12088);
xnor U12286 (N_12286,N_12189,N_12011);
xnor U12287 (N_12287,N_12054,N_12162);
nand U12288 (N_12288,N_12006,N_12036);
xnor U12289 (N_12289,N_12170,N_12104);
and U12290 (N_12290,N_12048,N_12169);
nor U12291 (N_12291,N_12193,N_12032);
and U12292 (N_12292,N_12128,N_12180);
xnor U12293 (N_12293,N_12163,N_12113);
nand U12294 (N_12294,N_12066,N_12158);
xor U12295 (N_12295,N_12173,N_12089);
xor U12296 (N_12296,N_12119,N_12096);
nand U12297 (N_12297,N_12196,N_12095);
xnor U12298 (N_12298,N_12016,N_12046);
or U12299 (N_12299,N_12041,N_12138);
and U12300 (N_12300,N_12144,N_12113);
xor U12301 (N_12301,N_12070,N_12100);
nor U12302 (N_12302,N_12169,N_12071);
or U12303 (N_12303,N_12129,N_12084);
and U12304 (N_12304,N_12077,N_12159);
and U12305 (N_12305,N_12065,N_12010);
nand U12306 (N_12306,N_12137,N_12143);
or U12307 (N_12307,N_12070,N_12160);
and U12308 (N_12308,N_12054,N_12029);
and U12309 (N_12309,N_12167,N_12085);
nand U12310 (N_12310,N_12142,N_12075);
nor U12311 (N_12311,N_12180,N_12077);
nand U12312 (N_12312,N_12066,N_12166);
nor U12313 (N_12313,N_12131,N_12102);
or U12314 (N_12314,N_12185,N_12142);
and U12315 (N_12315,N_12049,N_12028);
nor U12316 (N_12316,N_12055,N_12027);
and U12317 (N_12317,N_12163,N_12150);
xnor U12318 (N_12318,N_12072,N_12105);
nand U12319 (N_12319,N_12185,N_12008);
and U12320 (N_12320,N_12178,N_12012);
xor U12321 (N_12321,N_12079,N_12093);
nand U12322 (N_12322,N_12193,N_12008);
nand U12323 (N_12323,N_12061,N_12178);
nor U12324 (N_12324,N_12124,N_12008);
and U12325 (N_12325,N_12120,N_12066);
or U12326 (N_12326,N_12136,N_12081);
xor U12327 (N_12327,N_12157,N_12111);
nor U12328 (N_12328,N_12130,N_12065);
nand U12329 (N_12329,N_12174,N_12121);
nor U12330 (N_12330,N_12003,N_12190);
or U12331 (N_12331,N_12140,N_12151);
nor U12332 (N_12332,N_12134,N_12084);
nor U12333 (N_12333,N_12190,N_12100);
nor U12334 (N_12334,N_12110,N_12006);
xor U12335 (N_12335,N_12000,N_12060);
and U12336 (N_12336,N_12194,N_12108);
nor U12337 (N_12337,N_12024,N_12138);
nor U12338 (N_12338,N_12044,N_12079);
or U12339 (N_12339,N_12194,N_12122);
or U12340 (N_12340,N_12166,N_12103);
xor U12341 (N_12341,N_12119,N_12188);
xor U12342 (N_12342,N_12184,N_12100);
xnor U12343 (N_12343,N_12038,N_12141);
or U12344 (N_12344,N_12194,N_12137);
or U12345 (N_12345,N_12156,N_12066);
nor U12346 (N_12346,N_12179,N_12122);
or U12347 (N_12347,N_12141,N_12194);
xnor U12348 (N_12348,N_12161,N_12065);
and U12349 (N_12349,N_12042,N_12076);
and U12350 (N_12350,N_12193,N_12024);
nand U12351 (N_12351,N_12158,N_12128);
nand U12352 (N_12352,N_12079,N_12020);
nor U12353 (N_12353,N_12065,N_12018);
xor U12354 (N_12354,N_12015,N_12028);
and U12355 (N_12355,N_12084,N_12078);
xor U12356 (N_12356,N_12054,N_12131);
nand U12357 (N_12357,N_12186,N_12097);
or U12358 (N_12358,N_12096,N_12062);
or U12359 (N_12359,N_12090,N_12197);
nor U12360 (N_12360,N_12142,N_12039);
xnor U12361 (N_12361,N_12022,N_12125);
and U12362 (N_12362,N_12128,N_12029);
nand U12363 (N_12363,N_12017,N_12096);
nor U12364 (N_12364,N_12162,N_12154);
xnor U12365 (N_12365,N_12099,N_12003);
nand U12366 (N_12366,N_12032,N_12096);
xnor U12367 (N_12367,N_12017,N_12079);
or U12368 (N_12368,N_12154,N_12053);
or U12369 (N_12369,N_12034,N_12196);
nor U12370 (N_12370,N_12124,N_12039);
xor U12371 (N_12371,N_12181,N_12131);
nand U12372 (N_12372,N_12060,N_12040);
or U12373 (N_12373,N_12108,N_12132);
or U12374 (N_12374,N_12064,N_12052);
nand U12375 (N_12375,N_12143,N_12170);
nand U12376 (N_12376,N_12001,N_12189);
or U12377 (N_12377,N_12035,N_12093);
nor U12378 (N_12378,N_12050,N_12043);
nand U12379 (N_12379,N_12175,N_12027);
or U12380 (N_12380,N_12170,N_12073);
and U12381 (N_12381,N_12108,N_12107);
or U12382 (N_12382,N_12030,N_12181);
and U12383 (N_12383,N_12096,N_12114);
nor U12384 (N_12384,N_12174,N_12010);
xnor U12385 (N_12385,N_12020,N_12130);
nor U12386 (N_12386,N_12093,N_12121);
nor U12387 (N_12387,N_12080,N_12114);
and U12388 (N_12388,N_12173,N_12165);
nor U12389 (N_12389,N_12140,N_12197);
and U12390 (N_12390,N_12138,N_12189);
and U12391 (N_12391,N_12177,N_12020);
xor U12392 (N_12392,N_12106,N_12079);
nor U12393 (N_12393,N_12152,N_12113);
and U12394 (N_12394,N_12062,N_12036);
xor U12395 (N_12395,N_12148,N_12125);
xor U12396 (N_12396,N_12196,N_12064);
xor U12397 (N_12397,N_12191,N_12142);
nand U12398 (N_12398,N_12108,N_12169);
and U12399 (N_12399,N_12001,N_12019);
nor U12400 (N_12400,N_12399,N_12324);
nand U12401 (N_12401,N_12354,N_12371);
xor U12402 (N_12402,N_12289,N_12274);
nand U12403 (N_12403,N_12308,N_12233);
nand U12404 (N_12404,N_12266,N_12322);
nor U12405 (N_12405,N_12253,N_12278);
nand U12406 (N_12406,N_12311,N_12361);
nor U12407 (N_12407,N_12220,N_12342);
nand U12408 (N_12408,N_12334,N_12338);
or U12409 (N_12409,N_12295,N_12277);
nand U12410 (N_12410,N_12370,N_12376);
xnor U12411 (N_12411,N_12333,N_12218);
and U12412 (N_12412,N_12259,N_12280);
and U12413 (N_12413,N_12283,N_12262);
nand U12414 (N_12414,N_12307,N_12201);
xor U12415 (N_12415,N_12309,N_12299);
nand U12416 (N_12416,N_12362,N_12360);
or U12417 (N_12417,N_12287,N_12230);
and U12418 (N_12418,N_12237,N_12364);
and U12419 (N_12419,N_12368,N_12288);
and U12420 (N_12420,N_12235,N_12390);
nor U12421 (N_12421,N_12365,N_12205);
xor U12422 (N_12422,N_12330,N_12264);
and U12423 (N_12423,N_12336,N_12281);
nor U12424 (N_12424,N_12378,N_12319);
nor U12425 (N_12425,N_12377,N_12258);
or U12426 (N_12426,N_12238,N_12325);
nand U12427 (N_12427,N_12306,N_12315);
nor U12428 (N_12428,N_12391,N_12380);
and U12429 (N_12429,N_12369,N_12318);
nand U12430 (N_12430,N_12292,N_12305);
nand U12431 (N_12431,N_12227,N_12393);
nor U12432 (N_12432,N_12239,N_12385);
and U12433 (N_12433,N_12351,N_12245);
or U12434 (N_12434,N_12261,N_12214);
or U12435 (N_12435,N_12303,N_12341);
and U12436 (N_12436,N_12384,N_12257);
nor U12437 (N_12437,N_12265,N_12229);
or U12438 (N_12438,N_12296,N_12359);
xor U12439 (N_12439,N_12363,N_12328);
nor U12440 (N_12440,N_12202,N_12231);
or U12441 (N_12441,N_12314,N_12252);
and U12442 (N_12442,N_12276,N_12347);
and U12443 (N_12443,N_12355,N_12343);
nand U12444 (N_12444,N_12394,N_12268);
xor U12445 (N_12445,N_12397,N_12356);
and U12446 (N_12446,N_12381,N_12249);
or U12447 (N_12447,N_12221,N_12247);
and U12448 (N_12448,N_12358,N_12386);
xnor U12449 (N_12449,N_12300,N_12367);
or U12450 (N_12450,N_12374,N_12396);
nor U12451 (N_12451,N_12241,N_12317);
nor U12452 (N_12452,N_12254,N_12327);
xor U12453 (N_12453,N_12373,N_12302);
nor U12454 (N_12454,N_12348,N_12210);
or U12455 (N_12455,N_12226,N_12248);
and U12456 (N_12456,N_12366,N_12242);
or U12457 (N_12457,N_12215,N_12345);
nand U12458 (N_12458,N_12272,N_12304);
and U12459 (N_12459,N_12375,N_12337);
nor U12460 (N_12460,N_12207,N_12383);
and U12461 (N_12461,N_12282,N_12297);
and U12462 (N_12462,N_12301,N_12326);
and U12463 (N_12463,N_12284,N_12286);
or U12464 (N_12464,N_12243,N_12224);
nor U12465 (N_12465,N_12211,N_12291);
and U12466 (N_12466,N_12349,N_12200);
nand U12467 (N_12467,N_12216,N_12331);
nand U12468 (N_12468,N_12335,N_12255);
nand U12469 (N_12469,N_12398,N_12232);
nand U12470 (N_12470,N_12234,N_12382);
nand U12471 (N_12471,N_12206,N_12388);
nor U12472 (N_12472,N_12203,N_12273);
or U12473 (N_12473,N_12323,N_12350);
nor U12474 (N_12474,N_12285,N_12387);
xnor U12475 (N_12475,N_12329,N_12204);
nor U12476 (N_12476,N_12246,N_12395);
and U12477 (N_12477,N_12339,N_12250);
xnor U12478 (N_12478,N_12213,N_12267);
nand U12479 (N_12479,N_12293,N_12312);
nor U12480 (N_12480,N_12298,N_12219);
and U12481 (N_12481,N_12310,N_12344);
nand U12482 (N_12482,N_12320,N_12294);
or U12483 (N_12483,N_12379,N_12389);
and U12484 (N_12484,N_12372,N_12271);
or U12485 (N_12485,N_12275,N_12290);
or U12486 (N_12486,N_12332,N_12240);
or U12487 (N_12487,N_12208,N_12346);
and U12488 (N_12488,N_12313,N_12316);
nand U12489 (N_12489,N_12321,N_12244);
xor U12490 (N_12490,N_12392,N_12217);
or U12491 (N_12491,N_12340,N_12357);
or U12492 (N_12492,N_12223,N_12251);
nand U12493 (N_12493,N_12270,N_12228);
and U12494 (N_12494,N_12209,N_12263);
xnor U12495 (N_12495,N_12222,N_12353);
nor U12496 (N_12496,N_12269,N_12352);
and U12497 (N_12497,N_12236,N_12212);
and U12498 (N_12498,N_12279,N_12256);
and U12499 (N_12499,N_12260,N_12225);
xnor U12500 (N_12500,N_12361,N_12302);
or U12501 (N_12501,N_12258,N_12247);
nand U12502 (N_12502,N_12223,N_12344);
nand U12503 (N_12503,N_12293,N_12314);
and U12504 (N_12504,N_12359,N_12261);
or U12505 (N_12505,N_12257,N_12382);
nand U12506 (N_12506,N_12311,N_12248);
nand U12507 (N_12507,N_12232,N_12220);
or U12508 (N_12508,N_12203,N_12320);
xnor U12509 (N_12509,N_12279,N_12378);
or U12510 (N_12510,N_12209,N_12300);
xor U12511 (N_12511,N_12236,N_12220);
nand U12512 (N_12512,N_12271,N_12341);
nor U12513 (N_12513,N_12206,N_12207);
nand U12514 (N_12514,N_12287,N_12363);
nor U12515 (N_12515,N_12302,N_12244);
nor U12516 (N_12516,N_12304,N_12380);
nand U12517 (N_12517,N_12339,N_12274);
and U12518 (N_12518,N_12342,N_12258);
and U12519 (N_12519,N_12277,N_12325);
or U12520 (N_12520,N_12249,N_12227);
and U12521 (N_12521,N_12285,N_12312);
and U12522 (N_12522,N_12213,N_12331);
or U12523 (N_12523,N_12353,N_12393);
xnor U12524 (N_12524,N_12361,N_12392);
or U12525 (N_12525,N_12339,N_12358);
nor U12526 (N_12526,N_12253,N_12293);
or U12527 (N_12527,N_12348,N_12281);
xnor U12528 (N_12528,N_12253,N_12366);
nand U12529 (N_12529,N_12381,N_12269);
xnor U12530 (N_12530,N_12347,N_12374);
or U12531 (N_12531,N_12216,N_12312);
and U12532 (N_12532,N_12234,N_12383);
and U12533 (N_12533,N_12267,N_12207);
nor U12534 (N_12534,N_12392,N_12271);
and U12535 (N_12535,N_12215,N_12270);
nand U12536 (N_12536,N_12305,N_12348);
or U12537 (N_12537,N_12225,N_12393);
and U12538 (N_12538,N_12304,N_12392);
nor U12539 (N_12539,N_12233,N_12331);
and U12540 (N_12540,N_12256,N_12337);
xnor U12541 (N_12541,N_12332,N_12244);
or U12542 (N_12542,N_12327,N_12366);
and U12543 (N_12543,N_12304,N_12393);
nand U12544 (N_12544,N_12287,N_12348);
nand U12545 (N_12545,N_12226,N_12324);
and U12546 (N_12546,N_12382,N_12239);
and U12547 (N_12547,N_12297,N_12205);
xnor U12548 (N_12548,N_12305,N_12285);
and U12549 (N_12549,N_12211,N_12276);
xnor U12550 (N_12550,N_12307,N_12360);
and U12551 (N_12551,N_12264,N_12395);
xnor U12552 (N_12552,N_12379,N_12261);
xor U12553 (N_12553,N_12278,N_12343);
nand U12554 (N_12554,N_12329,N_12237);
xnor U12555 (N_12555,N_12377,N_12313);
xnor U12556 (N_12556,N_12354,N_12284);
nand U12557 (N_12557,N_12297,N_12225);
or U12558 (N_12558,N_12386,N_12258);
xor U12559 (N_12559,N_12277,N_12235);
nor U12560 (N_12560,N_12398,N_12210);
xnor U12561 (N_12561,N_12265,N_12267);
or U12562 (N_12562,N_12349,N_12297);
xor U12563 (N_12563,N_12296,N_12246);
and U12564 (N_12564,N_12302,N_12251);
or U12565 (N_12565,N_12341,N_12267);
nand U12566 (N_12566,N_12363,N_12332);
and U12567 (N_12567,N_12230,N_12395);
and U12568 (N_12568,N_12394,N_12316);
nand U12569 (N_12569,N_12368,N_12230);
nor U12570 (N_12570,N_12316,N_12251);
nor U12571 (N_12571,N_12301,N_12384);
nor U12572 (N_12572,N_12338,N_12352);
or U12573 (N_12573,N_12369,N_12248);
nand U12574 (N_12574,N_12373,N_12320);
nor U12575 (N_12575,N_12377,N_12279);
or U12576 (N_12576,N_12391,N_12248);
or U12577 (N_12577,N_12261,N_12362);
and U12578 (N_12578,N_12233,N_12333);
xnor U12579 (N_12579,N_12309,N_12353);
nor U12580 (N_12580,N_12395,N_12306);
nand U12581 (N_12581,N_12279,N_12316);
nand U12582 (N_12582,N_12281,N_12384);
or U12583 (N_12583,N_12358,N_12311);
or U12584 (N_12584,N_12381,N_12338);
nor U12585 (N_12585,N_12363,N_12343);
xor U12586 (N_12586,N_12263,N_12308);
nand U12587 (N_12587,N_12331,N_12348);
nand U12588 (N_12588,N_12224,N_12298);
xor U12589 (N_12589,N_12319,N_12241);
nor U12590 (N_12590,N_12295,N_12333);
nor U12591 (N_12591,N_12296,N_12346);
nor U12592 (N_12592,N_12279,N_12335);
xnor U12593 (N_12593,N_12264,N_12304);
and U12594 (N_12594,N_12247,N_12269);
xnor U12595 (N_12595,N_12256,N_12250);
or U12596 (N_12596,N_12325,N_12276);
or U12597 (N_12597,N_12298,N_12370);
or U12598 (N_12598,N_12299,N_12318);
or U12599 (N_12599,N_12259,N_12226);
xor U12600 (N_12600,N_12557,N_12483);
and U12601 (N_12601,N_12508,N_12414);
nand U12602 (N_12602,N_12424,N_12467);
and U12603 (N_12603,N_12520,N_12471);
xnor U12604 (N_12604,N_12404,N_12579);
nand U12605 (N_12605,N_12554,N_12451);
nand U12606 (N_12606,N_12582,N_12443);
xnor U12607 (N_12607,N_12574,N_12409);
or U12608 (N_12608,N_12519,N_12495);
nor U12609 (N_12609,N_12400,N_12518);
and U12610 (N_12610,N_12457,N_12550);
nand U12611 (N_12611,N_12597,N_12410);
nor U12612 (N_12612,N_12419,N_12425);
or U12613 (N_12613,N_12543,N_12448);
nor U12614 (N_12614,N_12506,N_12561);
nor U12615 (N_12615,N_12526,N_12405);
xnor U12616 (N_12616,N_12403,N_12423);
or U12617 (N_12617,N_12479,N_12453);
xor U12618 (N_12618,N_12527,N_12573);
xnor U12619 (N_12619,N_12496,N_12547);
or U12620 (N_12620,N_12464,N_12489);
and U12621 (N_12621,N_12462,N_12504);
nand U12622 (N_12622,N_12456,N_12418);
nor U12623 (N_12623,N_12500,N_12583);
xnor U12624 (N_12624,N_12412,N_12524);
and U12625 (N_12625,N_12509,N_12593);
or U12626 (N_12626,N_12569,N_12580);
and U12627 (N_12627,N_12522,N_12470);
or U12628 (N_12628,N_12477,N_12570);
nand U12629 (N_12629,N_12577,N_12539);
xor U12630 (N_12630,N_12581,N_12560);
nand U12631 (N_12631,N_12502,N_12534);
nor U12632 (N_12632,N_12528,N_12490);
xnor U12633 (N_12633,N_12440,N_12562);
nor U12634 (N_12634,N_12511,N_12540);
nor U12635 (N_12635,N_12567,N_12454);
and U12636 (N_12636,N_12559,N_12594);
or U12637 (N_12637,N_12576,N_12463);
or U12638 (N_12638,N_12445,N_12564);
and U12639 (N_12639,N_12499,N_12481);
nand U12640 (N_12640,N_12523,N_12517);
nand U12641 (N_12641,N_12475,N_12406);
xor U12642 (N_12642,N_12455,N_12599);
nor U12643 (N_12643,N_12482,N_12497);
xor U12644 (N_12644,N_12461,N_12537);
or U12645 (N_12645,N_12415,N_12474);
nand U12646 (N_12646,N_12429,N_12472);
nor U12647 (N_12647,N_12563,N_12592);
or U12648 (N_12648,N_12436,N_12476);
nand U12649 (N_12649,N_12441,N_12447);
or U12650 (N_12650,N_12452,N_12469);
and U12651 (N_12651,N_12512,N_12525);
nand U12652 (N_12652,N_12551,N_12450);
nand U12653 (N_12653,N_12439,N_12434);
or U12654 (N_12654,N_12488,N_12485);
nand U12655 (N_12655,N_12468,N_12480);
and U12656 (N_12656,N_12402,N_12433);
nand U12657 (N_12657,N_12421,N_12510);
or U12658 (N_12658,N_12498,N_12531);
nor U12659 (N_12659,N_12458,N_12487);
or U12660 (N_12660,N_12493,N_12516);
nor U12661 (N_12661,N_12521,N_12478);
or U12662 (N_12662,N_12568,N_12501);
xor U12663 (N_12663,N_12558,N_12492);
xnor U12664 (N_12664,N_12432,N_12556);
xor U12665 (N_12665,N_12473,N_12588);
nand U12666 (N_12666,N_12536,N_12589);
xor U12667 (N_12667,N_12446,N_12430);
xor U12668 (N_12668,N_12428,N_12542);
nand U12669 (N_12669,N_12459,N_12532);
or U12670 (N_12670,N_12555,N_12465);
nor U12671 (N_12671,N_12438,N_12426);
and U12672 (N_12672,N_12422,N_12587);
nor U12673 (N_12673,N_12533,N_12598);
or U12674 (N_12674,N_12548,N_12553);
nand U12675 (N_12675,N_12435,N_12529);
and U12676 (N_12676,N_12444,N_12596);
nand U12677 (N_12677,N_12590,N_12575);
nor U12678 (N_12678,N_12507,N_12515);
or U12679 (N_12679,N_12431,N_12571);
nand U12680 (N_12680,N_12460,N_12514);
nor U12681 (N_12681,N_12449,N_12484);
or U12682 (N_12682,N_12535,N_12420);
and U12683 (N_12683,N_12586,N_12416);
or U12684 (N_12684,N_12584,N_12585);
nand U12685 (N_12685,N_12486,N_12552);
xnor U12686 (N_12686,N_12591,N_12541);
nor U12687 (N_12687,N_12595,N_12565);
xnor U12688 (N_12688,N_12513,N_12545);
nor U12689 (N_12689,N_12442,N_12538);
or U12690 (N_12690,N_12437,N_12491);
nor U12691 (N_12691,N_12549,N_12427);
and U12692 (N_12692,N_12503,N_12572);
xor U12693 (N_12693,N_12417,N_12411);
or U12694 (N_12694,N_12544,N_12530);
nand U12695 (N_12695,N_12413,N_12494);
nor U12696 (N_12696,N_12546,N_12466);
nor U12697 (N_12697,N_12505,N_12566);
and U12698 (N_12698,N_12407,N_12401);
nand U12699 (N_12699,N_12578,N_12408);
and U12700 (N_12700,N_12478,N_12565);
nor U12701 (N_12701,N_12460,N_12482);
and U12702 (N_12702,N_12550,N_12473);
and U12703 (N_12703,N_12413,N_12408);
xor U12704 (N_12704,N_12418,N_12446);
xor U12705 (N_12705,N_12403,N_12519);
nor U12706 (N_12706,N_12593,N_12581);
and U12707 (N_12707,N_12491,N_12405);
nor U12708 (N_12708,N_12476,N_12443);
nand U12709 (N_12709,N_12444,N_12591);
xnor U12710 (N_12710,N_12423,N_12519);
xnor U12711 (N_12711,N_12403,N_12510);
xor U12712 (N_12712,N_12403,N_12532);
nor U12713 (N_12713,N_12562,N_12490);
xnor U12714 (N_12714,N_12468,N_12465);
or U12715 (N_12715,N_12558,N_12536);
xor U12716 (N_12716,N_12435,N_12559);
and U12717 (N_12717,N_12513,N_12566);
nor U12718 (N_12718,N_12483,N_12418);
or U12719 (N_12719,N_12518,N_12556);
nand U12720 (N_12720,N_12408,N_12496);
nor U12721 (N_12721,N_12587,N_12521);
nand U12722 (N_12722,N_12434,N_12466);
and U12723 (N_12723,N_12450,N_12532);
nor U12724 (N_12724,N_12435,N_12404);
xor U12725 (N_12725,N_12487,N_12423);
and U12726 (N_12726,N_12441,N_12420);
xnor U12727 (N_12727,N_12547,N_12413);
xnor U12728 (N_12728,N_12404,N_12483);
nor U12729 (N_12729,N_12515,N_12418);
xnor U12730 (N_12730,N_12520,N_12532);
or U12731 (N_12731,N_12438,N_12597);
or U12732 (N_12732,N_12452,N_12450);
nand U12733 (N_12733,N_12452,N_12512);
and U12734 (N_12734,N_12411,N_12496);
xor U12735 (N_12735,N_12489,N_12457);
nor U12736 (N_12736,N_12494,N_12508);
and U12737 (N_12737,N_12445,N_12500);
xor U12738 (N_12738,N_12458,N_12495);
nor U12739 (N_12739,N_12542,N_12421);
or U12740 (N_12740,N_12503,N_12597);
or U12741 (N_12741,N_12438,N_12403);
nand U12742 (N_12742,N_12531,N_12530);
nand U12743 (N_12743,N_12464,N_12447);
xor U12744 (N_12744,N_12514,N_12467);
xor U12745 (N_12745,N_12544,N_12560);
nor U12746 (N_12746,N_12556,N_12427);
nor U12747 (N_12747,N_12429,N_12432);
nand U12748 (N_12748,N_12485,N_12487);
xnor U12749 (N_12749,N_12470,N_12517);
or U12750 (N_12750,N_12586,N_12423);
or U12751 (N_12751,N_12443,N_12405);
nor U12752 (N_12752,N_12530,N_12581);
xnor U12753 (N_12753,N_12582,N_12560);
xor U12754 (N_12754,N_12535,N_12530);
xor U12755 (N_12755,N_12460,N_12443);
nand U12756 (N_12756,N_12458,N_12512);
nor U12757 (N_12757,N_12416,N_12519);
and U12758 (N_12758,N_12413,N_12424);
nand U12759 (N_12759,N_12566,N_12540);
xor U12760 (N_12760,N_12432,N_12446);
xnor U12761 (N_12761,N_12592,N_12498);
and U12762 (N_12762,N_12453,N_12575);
xor U12763 (N_12763,N_12532,N_12551);
and U12764 (N_12764,N_12495,N_12589);
nand U12765 (N_12765,N_12456,N_12530);
and U12766 (N_12766,N_12540,N_12459);
nand U12767 (N_12767,N_12514,N_12435);
and U12768 (N_12768,N_12410,N_12504);
nand U12769 (N_12769,N_12548,N_12454);
or U12770 (N_12770,N_12532,N_12466);
nand U12771 (N_12771,N_12467,N_12573);
nand U12772 (N_12772,N_12535,N_12490);
nand U12773 (N_12773,N_12497,N_12540);
nor U12774 (N_12774,N_12545,N_12465);
and U12775 (N_12775,N_12596,N_12442);
nor U12776 (N_12776,N_12488,N_12440);
and U12777 (N_12777,N_12461,N_12478);
and U12778 (N_12778,N_12586,N_12593);
or U12779 (N_12779,N_12508,N_12442);
or U12780 (N_12780,N_12445,N_12483);
nor U12781 (N_12781,N_12467,N_12468);
nand U12782 (N_12782,N_12497,N_12489);
and U12783 (N_12783,N_12483,N_12536);
xor U12784 (N_12784,N_12474,N_12432);
xor U12785 (N_12785,N_12443,N_12584);
nor U12786 (N_12786,N_12442,N_12476);
or U12787 (N_12787,N_12441,N_12453);
nor U12788 (N_12788,N_12525,N_12418);
nor U12789 (N_12789,N_12568,N_12435);
nor U12790 (N_12790,N_12426,N_12479);
nand U12791 (N_12791,N_12411,N_12501);
or U12792 (N_12792,N_12551,N_12587);
nor U12793 (N_12793,N_12561,N_12518);
nand U12794 (N_12794,N_12548,N_12523);
or U12795 (N_12795,N_12518,N_12506);
nor U12796 (N_12796,N_12593,N_12549);
nand U12797 (N_12797,N_12517,N_12459);
xnor U12798 (N_12798,N_12571,N_12487);
nor U12799 (N_12799,N_12430,N_12477);
and U12800 (N_12800,N_12727,N_12613);
and U12801 (N_12801,N_12635,N_12695);
and U12802 (N_12802,N_12628,N_12605);
or U12803 (N_12803,N_12651,N_12652);
and U12804 (N_12804,N_12688,N_12729);
and U12805 (N_12805,N_12756,N_12629);
xnor U12806 (N_12806,N_12607,N_12786);
nand U12807 (N_12807,N_12743,N_12700);
xor U12808 (N_12808,N_12779,N_12775);
or U12809 (N_12809,N_12661,N_12603);
nand U12810 (N_12810,N_12722,N_12691);
nor U12811 (N_12811,N_12718,N_12634);
and U12812 (N_12812,N_12708,N_12602);
xor U12813 (N_12813,N_12793,N_12740);
xor U12814 (N_12814,N_12766,N_12707);
or U12815 (N_12815,N_12686,N_12794);
nand U12816 (N_12816,N_12697,N_12716);
and U12817 (N_12817,N_12667,N_12654);
xor U12818 (N_12818,N_12702,N_12683);
or U12819 (N_12819,N_12776,N_12730);
or U12820 (N_12820,N_12737,N_12690);
nor U12821 (N_12821,N_12642,N_12744);
and U12822 (N_12822,N_12609,N_12783);
xor U12823 (N_12823,N_12692,N_12693);
nor U12824 (N_12824,N_12770,N_12734);
nand U12825 (N_12825,N_12763,N_12610);
nand U12826 (N_12826,N_12762,N_12627);
and U12827 (N_12827,N_12694,N_12626);
nor U12828 (N_12828,N_12666,N_12752);
or U12829 (N_12829,N_12647,N_12753);
xnor U12830 (N_12830,N_12789,N_12731);
xor U12831 (N_12831,N_12780,N_12724);
and U12832 (N_12832,N_12799,N_12678);
xnor U12833 (N_12833,N_12796,N_12787);
xnor U12834 (N_12834,N_12664,N_12710);
xnor U12835 (N_12835,N_12736,N_12767);
nand U12836 (N_12836,N_12640,N_12746);
and U12837 (N_12837,N_12742,N_12791);
nand U12838 (N_12838,N_12649,N_12798);
nand U12839 (N_12839,N_12696,N_12677);
or U12840 (N_12840,N_12772,N_12738);
or U12841 (N_12841,N_12687,N_12631);
and U12842 (N_12842,N_12606,N_12726);
or U12843 (N_12843,N_12785,N_12633);
or U12844 (N_12844,N_12714,N_12689);
nor U12845 (N_12845,N_12673,N_12623);
or U12846 (N_12846,N_12725,N_12748);
nor U12847 (N_12847,N_12701,N_12675);
nor U12848 (N_12848,N_12636,N_12709);
nand U12849 (N_12849,N_12625,N_12788);
and U12850 (N_12850,N_12632,N_12717);
nor U12851 (N_12851,N_12614,N_12765);
nand U12852 (N_12852,N_12679,N_12764);
xor U12853 (N_12853,N_12622,N_12648);
and U12854 (N_12854,N_12620,N_12790);
and U12855 (N_12855,N_12618,N_12778);
and U12856 (N_12856,N_12741,N_12615);
nand U12857 (N_12857,N_12668,N_12676);
nor U12858 (N_12858,N_12604,N_12712);
or U12859 (N_12859,N_12761,N_12711);
nand U12860 (N_12860,N_12733,N_12641);
or U12861 (N_12861,N_12777,N_12728);
xor U12862 (N_12862,N_12732,N_12760);
or U12863 (N_12863,N_12784,N_12672);
xor U12864 (N_12864,N_12619,N_12656);
or U12865 (N_12865,N_12655,N_12745);
xnor U12866 (N_12866,N_12608,N_12774);
or U12867 (N_12867,N_12624,N_12768);
or U12868 (N_12868,N_12616,N_12660);
nand U12869 (N_12869,N_12755,N_12663);
xor U12870 (N_12870,N_12721,N_12751);
xnor U12871 (N_12871,N_12769,N_12637);
nor U12872 (N_12872,N_12703,N_12719);
nand U12873 (N_12873,N_12617,N_12681);
nor U12874 (N_12874,N_12758,N_12630);
xor U12875 (N_12875,N_12792,N_12644);
nand U12876 (N_12876,N_12747,N_12643);
and U12877 (N_12877,N_12680,N_12638);
or U12878 (N_12878,N_12621,N_12658);
nor U12879 (N_12879,N_12704,N_12600);
nand U12880 (N_12880,N_12662,N_12735);
nor U12881 (N_12881,N_12612,N_12781);
nand U12882 (N_12882,N_12699,N_12670);
and U12883 (N_12883,N_12650,N_12669);
nor U12884 (N_12884,N_12757,N_12771);
nand U12885 (N_12885,N_12698,N_12754);
or U12886 (N_12886,N_12797,N_12671);
nor U12887 (N_12887,N_12759,N_12706);
and U12888 (N_12888,N_12674,N_12713);
or U12889 (N_12889,N_12723,N_12682);
nor U12890 (N_12890,N_12659,N_12782);
and U12891 (N_12891,N_12715,N_12749);
xnor U12892 (N_12892,N_12639,N_12611);
nor U12893 (N_12893,N_12653,N_12795);
nor U12894 (N_12894,N_12665,N_12705);
nor U12895 (N_12895,N_12684,N_12645);
nand U12896 (N_12896,N_12739,N_12750);
nand U12897 (N_12897,N_12685,N_12657);
and U12898 (N_12898,N_12601,N_12646);
xnor U12899 (N_12899,N_12720,N_12773);
and U12900 (N_12900,N_12778,N_12760);
and U12901 (N_12901,N_12731,N_12748);
or U12902 (N_12902,N_12772,N_12743);
xor U12903 (N_12903,N_12611,N_12749);
xnor U12904 (N_12904,N_12653,N_12788);
xor U12905 (N_12905,N_12637,N_12609);
xor U12906 (N_12906,N_12624,N_12729);
nand U12907 (N_12907,N_12707,N_12602);
nand U12908 (N_12908,N_12760,N_12722);
nor U12909 (N_12909,N_12639,N_12686);
nand U12910 (N_12910,N_12774,N_12731);
xor U12911 (N_12911,N_12610,N_12734);
or U12912 (N_12912,N_12600,N_12619);
or U12913 (N_12913,N_12697,N_12609);
or U12914 (N_12914,N_12752,N_12636);
nand U12915 (N_12915,N_12674,N_12696);
nand U12916 (N_12916,N_12617,N_12690);
xnor U12917 (N_12917,N_12682,N_12687);
xor U12918 (N_12918,N_12636,N_12737);
nor U12919 (N_12919,N_12600,N_12672);
xnor U12920 (N_12920,N_12624,N_12758);
or U12921 (N_12921,N_12722,N_12725);
and U12922 (N_12922,N_12681,N_12677);
and U12923 (N_12923,N_12744,N_12735);
xor U12924 (N_12924,N_12676,N_12672);
xnor U12925 (N_12925,N_12636,N_12663);
xnor U12926 (N_12926,N_12615,N_12787);
nor U12927 (N_12927,N_12656,N_12631);
xor U12928 (N_12928,N_12650,N_12632);
xor U12929 (N_12929,N_12678,N_12613);
or U12930 (N_12930,N_12685,N_12620);
nor U12931 (N_12931,N_12635,N_12733);
xnor U12932 (N_12932,N_12675,N_12645);
or U12933 (N_12933,N_12665,N_12610);
xor U12934 (N_12934,N_12658,N_12736);
nor U12935 (N_12935,N_12615,N_12637);
or U12936 (N_12936,N_12796,N_12730);
or U12937 (N_12937,N_12771,N_12661);
nor U12938 (N_12938,N_12797,N_12686);
nor U12939 (N_12939,N_12704,N_12746);
nor U12940 (N_12940,N_12795,N_12624);
xnor U12941 (N_12941,N_12722,N_12739);
nor U12942 (N_12942,N_12648,N_12693);
xor U12943 (N_12943,N_12667,N_12617);
and U12944 (N_12944,N_12679,N_12655);
nand U12945 (N_12945,N_12789,N_12796);
nand U12946 (N_12946,N_12662,N_12642);
nand U12947 (N_12947,N_12708,N_12768);
or U12948 (N_12948,N_12641,N_12660);
xor U12949 (N_12949,N_12616,N_12790);
nor U12950 (N_12950,N_12769,N_12613);
xnor U12951 (N_12951,N_12760,N_12682);
xnor U12952 (N_12952,N_12619,N_12612);
and U12953 (N_12953,N_12633,N_12624);
xnor U12954 (N_12954,N_12772,N_12690);
nor U12955 (N_12955,N_12628,N_12643);
nand U12956 (N_12956,N_12727,N_12614);
nor U12957 (N_12957,N_12688,N_12652);
nor U12958 (N_12958,N_12654,N_12713);
nor U12959 (N_12959,N_12633,N_12681);
nand U12960 (N_12960,N_12601,N_12619);
or U12961 (N_12961,N_12643,N_12625);
or U12962 (N_12962,N_12799,N_12672);
nor U12963 (N_12963,N_12699,N_12601);
xnor U12964 (N_12964,N_12774,N_12753);
or U12965 (N_12965,N_12746,N_12625);
and U12966 (N_12966,N_12628,N_12646);
nand U12967 (N_12967,N_12787,N_12744);
nor U12968 (N_12968,N_12708,N_12728);
nor U12969 (N_12969,N_12657,N_12682);
xnor U12970 (N_12970,N_12748,N_12645);
xor U12971 (N_12971,N_12728,N_12711);
nand U12972 (N_12972,N_12646,N_12644);
xor U12973 (N_12973,N_12709,N_12722);
nand U12974 (N_12974,N_12608,N_12650);
nand U12975 (N_12975,N_12789,N_12774);
xor U12976 (N_12976,N_12694,N_12750);
nand U12977 (N_12977,N_12718,N_12639);
or U12978 (N_12978,N_12717,N_12648);
nor U12979 (N_12979,N_12675,N_12770);
xor U12980 (N_12980,N_12728,N_12733);
nand U12981 (N_12981,N_12765,N_12623);
or U12982 (N_12982,N_12615,N_12743);
nand U12983 (N_12983,N_12640,N_12685);
nor U12984 (N_12984,N_12796,N_12742);
nand U12985 (N_12985,N_12671,N_12770);
nor U12986 (N_12986,N_12665,N_12641);
nor U12987 (N_12987,N_12617,N_12640);
and U12988 (N_12988,N_12759,N_12641);
xnor U12989 (N_12989,N_12628,N_12765);
xor U12990 (N_12990,N_12724,N_12605);
and U12991 (N_12991,N_12693,N_12643);
xnor U12992 (N_12992,N_12607,N_12653);
nand U12993 (N_12993,N_12768,N_12782);
nand U12994 (N_12994,N_12698,N_12692);
nor U12995 (N_12995,N_12675,N_12630);
nor U12996 (N_12996,N_12752,N_12608);
xnor U12997 (N_12997,N_12725,N_12627);
nand U12998 (N_12998,N_12674,N_12742);
or U12999 (N_12999,N_12739,N_12719);
xor U13000 (N_13000,N_12940,N_12844);
and U13001 (N_13001,N_12986,N_12864);
nor U13002 (N_13002,N_12947,N_12835);
nand U13003 (N_13003,N_12906,N_12909);
nor U13004 (N_13004,N_12816,N_12828);
nand U13005 (N_13005,N_12978,N_12899);
and U13006 (N_13006,N_12992,N_12841);
and U13007 (N_13007,N_12920,N_12960);
nand U13008 (N_13008,N_12945,N_12866);
or U13009 (N_13009,N_12815,N_12819);
and U13010 (N_13010,N_12907,N_12865);
and U13011 (N_13011,N_12919,N_12921);
xnor U13012 (N_13012,N_12888,N_12878);
nor U13013 (N_13013,N_12814,N_12957);
or U13014 (N_13014,N_12831,N_12818);
nor U13015 (N_13015,N_12933,N_12840);
and U13016 (N_13016,N_12857,N_12853);
xnor U13017 (N_13017,N_12944,N_12953);
xor U13018 (N_13018,N_12833,N_12923);
nand U13019 (N_13019,N_12860,N_12990);
and U13020 (N_13020,N_12859,N_12809);
nand U13021 (N_13021,N_12873,N_12991);
xor U13022 (N_13022,N_12910,N_12966);
nand U13023 (N_13023,N_12823,N_12892);
nand U13024 (N_13024,N_12897,N_12961);
xnor U13025 (N_13025,N_12948,N_12874);
and U13026 (N_13026,N_12916,N_12881);
and U13027 (N_13027,N_12880,N_12882);
nand U13028 (N_13028,N_12943,N_12850);
nor U13029 (N_13029,N_12810,N_12996);
or U13030 (N_13030,N_12984,N_12847);
xnor U13031 (N_13031,N_12995,N_12958);
xor U13032 (N_13032,N_12912,N_12908);
or U13033 (N_13033,N_12855,N_12830);
or U13034 (N_13034,N_12900,N_12889);
nor U13035 (N_13035,N_12974,N_12970);
nand U13036 (N_13036,N_12851,N_12869);
or U13037 (N_13037,N_12926,N_12805);
nand U13038 (N_13038,N_12934,N_12971);
nand U13039 (N_13039,N_12885,N_12854);
or U13040 (N_13040,N_12858,N_12904);
and U13041 (N_13041,N_12849,N_12973);
and U13042 (N_13042,N_12821,N_12925);
and U13043 (N_13043,N_12965,N_12848);
nand U13044 (N_13044,N_12883,N_12988);
or U13045 (N_13045,N_12879,N_12824);
xnor U13046 (N_13046,N_12905,N_12829);
and U13047 (N_13047,N_12942,N_12817);
nor U13048 (N_13048,N_12967,N_12994);
and U13049 (N_13049,N_12915,N_12832);
or U13050 (N_13050,N_12838,N_12887);
xor U13051 (N_13051,N_12976,N_12935);
or U13052 (N_13052,N_12895,N_12964);
nor U13053 (N_13053,N_12929,N_12954);
and U13054 (N_13054,N_12890,N_12804);
nor U13055 (N_13055,N_12927,N_12914);
xnor U13056 (N_13056,N_12875,N_12977);
or U13057 (N_13057,N_12997,N_12913);
xnor U13058 (N_13058,N_12979,N_12877);
xnor U13059 (N_13059,N_12802,N_12808);
nand U13060 (N_13060,N_12839,N_12959);
and U13061 (N_13061,N_12852,N_12956);
or U13062 (N_13062,N_12918,N_12811);
nor U13063 (N_13063,N_12922,N_12803);
nand U13064 (N_13064,N_12863,N_12980);
or U13065 (N_13065,N_12872,N_12932);
nand U13066 (N_13066,N_12845,N_12972);
or U13067 (N_13067,N_12813,N_12968);
nor U13068 (N_13068,N_12820,N_12999);
nor U13069 (N_13069,N_12955,N_12938);
and U13070 (N_13070,N_12812,N_12868);
xor U13071 (N_13071,N_12951,N_12937);
xor U13072 (N_13072,N_12985,N_12806);
xor U13073 (N_13073,N_12928,N_12982);
xnor U13074 (N_13074,N_12861,N_12822);
or U13075 (N_13075,N_12876,N_12825);
nor U13076 (N_13076,N_12941,N_12901);
nand U13077 (N_13077,N_12950,N_12870);
nor U13078 (N_13078,N_12963,N_12893);
xnor U13079 (N_13079,N_12843,N_12862);
nand U13080 (N_13080,N_12989,N_12952);
and U13081 (N_13081,N_12898,N_12983);
nand U13082 (N_13082,N_12884,N_12981);
nand U13083 (N_13083,N_12834,N_12807);
nand U13084 (N_13084,N_12924,N_12800);
and U13085 (N_13085,N_12896,N_12998);
nand U13086 (N_13086,N_12826,N_12962);
nand U13087 (N_13087,N_12886,N_12891);
nor U13088 (N_13088,N_12894,N_12842);
nor U13089 (N_13089,N_12837,N_12936);
or U13090 (N_13090,N_12911,N_12969);
and U13091 (N_13091,N_12949,N_12946);
nand U13092 (N_13092,N_12856,N_12846);
nand U13093 (N_13093,N_12867,N_12827);
and U13094 (N_13094,N_12902,N_12917);
and U13095 (N_13095,N_12871,N_12931);
or U13096 (N_13096,N_12993,N_12930);
and U13097 (N_13097,N_12987,N_12939);
and U13098 (N_13098,N_12903,N_12801);
nor U13099 (N_13099,N_12836,N_12975);
nor U13100 (N_13100,N_12826,N_12972);
nand U13101 (N_13101,N_12863,N_12944);
nand U13102 (N_13102,N_12859,N_12914);
nor U13103 (N_13103,N_12951,N_12901);
or U13104 (N_13104,N_12929,N_12980);
or U13105 (N_13105,N_12995,N_12879);
xnor U13106 (N_13106,N_12918,N_12891);
nor U13107 (N_13107,N_12943,N_12958);
and U13108 (N_13108,N_12823,N_12956);
nor U13109 (N_13109,N_12978,N_12997);
xnor U13110 (N_13110,N_12983,N_12861);
or U13111 (N_13111,N_12869,N_12918);
nand U13112 (N_13112,N_12838,N_12877);
xor U13113 (N_13113,N_12852,N_12982);
nor U13114 (N_13114,N_12816,N_12834);
nor U13115 (N_13115,N_12882,N_12990);
or U13116 (N_13116,N_12914,N_12823);
xor U13117 (N_13117,N_12917,N_12836);
nand U13118 (N_13118,N_12947,N_12855);
xnor U13119 (N_13119,N_12906,N_12840);
xnor U13120 (N_13120,N_12932,N_12917);
nor U13121 (N_13121,N_12985,N_12954);
xor U13122 (N_13122,N_12915,N_12929);
xnor U13123 (N_13123,N_12809,N_12953);
xnor U13124 (N_13124,N_12892,N_12988);
xor U13125 (N_13125,N_12907,N_12922);
or U13126 (N_13126,N_12925,N_12994);
xnor U13127 (N_13127,N_12978,N_12824);
or U13128 (N_13128,N_12995,N_12903);
or U13129 (N_13129,N_12893,N_12895);
nor U13130 (N_13130,N_12986,N_12882);
nor U13131 (N_13131,N_12887,N_12977);
or U13132 (N_13132,N_12935,N_12984);
and U13133 (N_13133,N_12974,N_12953);
or U13134 (N_13134,N_12996,N_12936);
xor U13135 (N_13135,N_12993,N_12904);
nor U13136 (N_13136,N_12822,N_12942);
or U13137 (N_13137,N_12886,N_12830);
nand U13138 (N_13138,N_12878,N_12913);
nor U13139 (N_13139,N_12818,N_12808);
nand U13140 (N_13140,N_12898,N_12913);
nand U13141 (N_13141,N_12941,N_12934);
xnor U13142 (N_13142,N_12968,N_12920);
and U13143 (N_13143,N_12925,N_12923);
nor U13144 (N_13144,N_12832,N_12891);
xnor U13145 (N_13145,N_12897,N_12903);
nor U13146 (N_13146,N_12848,N_12974);
and U13147 (N_13147,N_12860,N_12975);
and U13148 (N_13148,N_12870,N_12822);
nor U13149 (N_13149,N_12981,N_12904);
and U13150 (N_13150,N_12925,N_12812);
nand U13151 (N_13151,N_12926,N_12898);
or U13152 (N_13152,N_12876,N_12873);
nand U13153 (N_13153,N_12929,N_12845);
xor U13154 (N_13154,N_12978,N_12936);
xor U13155 (N_13155,N_12844,N_12913);
or U13156 (N_13156,N_12806,N_12994);
nor U13157 (N_13157,N_12809,N_12860);
xnor U13158 (N_13158,N_12940,N_12833);
and U13159 (N_13159,N_12993,N_12983);
or U13160 (N_13160,N_12866,N_12825);
or U13161 (N_13161,N_12842,N_12995);
or U13162 (N_13162,N_12943,N_12879);
nor U13163 (N_13163,N_12987,N_12807);
xnor U13164 (N_13164,N_12838,N_12883);
or U13165 (N_13165,N_12872,N_12904);
and U13166 (N_13166,N_12841,N_12878);
nor U13167 (N_13167,N_12846,N_12821);
and U13168 (N_13168,N_12810,N_12833);
xor U13169 (N_13169,N_12828,N_12839);
xnor U13170 (N_13170,N_12950,N_12940);
nand U13171 (N_13171,N_12995,N_12869);
nand U13172 (N_13172,N_12836,N_12887);
and U13173 (N_13173,N_12844,N_12947);
and U13174 (N_13174,N_12949,N_12874);
nand U13175 (N_13175,N_12904,N_12818);
nor U13176 (N_13176,N_12832,N_12908);
nand U13177 (N_13177,N_12908,N_12837);
or U13178 (N_13178,N_12834,N_12920);
nand U13179 (N_13179,N_12951,N_12814);
nor U13180 (N_13180,N_12852,N_12936);
nor U13181 (N_13181,N_12887,N_12916);
xor U13182 (N_13182,N_12933,N_12924);
nand U13183 (N_13183,N_12831,N_12917);
and U13184 (N_13184,N_12997,N_12915);
nand U13185 (N_13185,N_12958,N_12864);
and U13186 (N_13186,N_12857,N_12815);
nor U13187 (N_13187,N_12960,N_12899);
or U13188 (N_13188,N_12912,N_12979);
nand U13189 (N_13189,N_12807,N_12950);
xor U13190 (N_13190,N_12840,N_12967);
or U13191 (N_13191,N_12845,N_12831);
nor U13192 (N_13192,N_12921,N_12939);
or U13193 (N_13193,N_12860,N_12939);
xnor U13194 (N_13194,N_12902,N_12813);
nand U13195 (N_13195,N_12803,N_12908);
or U13196 (N_13196,N_12831,N_12933);
nor U13197 (N_13197,N_12837,N_12892);
and U13198 (N_13198,N_12909,N_12934);
and U13199 (N_13199,N_12872,N_12984);
or U13200 (N_13200,N_13198,N_13038);
xnor U13201 (N_13201,N_13086,N_13121);
nor U13202 (N_13202,N_13103,N_13126);
xor U13203 (N_13203,N_13075,N_13000);
nand U13204 (N_13204,N_13181,N_13164);
xor U13205 (N_13205,N_13051,N_13183);
or U13206 (N_13206,N_13053,N_13050);
nand U13207 (N_13207,N_13008,N_13015);
nor U13208 (N_13208,N_13160,N_13009);
nand U13209 (N_13209,N_13025,N_13157);
and U13210 (N_13210,N_13057,N_13066);
or U13211 (N_13211,N_13150,N_13058);
nand U13212 (N_13212,N_13090,N_13145);
nor U13213 (N_13213,N_13135,N_13077);
and U13214 (N_13214,N_13108,N_13029);
or U13215 (N_13215,N_13113,N_13042);
nand U13216 (N_13216,N_13041,N_13191);
nand U13217 (N_13217,N_13193,N_13073);
xnor U13218 (N_13218,N_13007,N_13177);
xnor U13219 (N_13219,N_13156,N_13039);
xor U13220 (N_13220,N_13137,N_13169);
or U13221 (N_13221,N_13083,N_13030);
nand U13222 (N_13222,N_13159,N_13199);
nor U13223 (N_13223,N_13140,N_13004);
nor U13224 (N_13224,N_13054,N_13080);
nand U13225 (N_13225,N_13011,N_13104);
and U13226 (N_13226,N_13123,N_13125);
and U13227 (N_13227,N_13189,N_13153);
or U13228 (N_13228,N_13045,N_13147);
and U13229 (N_13229,N_13176,N_13163);
nand U13230 (N_13230,N_13087,N_13035);
nand U13231 (N_13231,N_13184,N_13143);
xnor U13232 (N_13232,N_13100,N_13152);
xor U13233 (N_13233,N_13052,N_13196);
xor U13234 (N_13234,N_13064,N_13119);
nand U13235 (N_13235,N_13102,N_13144);
xnor U13236 (N_13236,N_13017,N_13016);
or U13237 (N_13237,N_13168,N_13106);
xnor U13238 (N_13238,N_13118,N_13188);
and U13239 (N_13239,N_13129,N_13120);
and U13240 (N_13240,N_13138,N_13161);
nor U13241 (N_13241,N_13022,N_13142);
or U13242 (N_13242,N_13170,N_13047);
or U13243 (N_13243,N_13115,N_13018);
nor U13244 (N_13244,N_13048,N_13044);
or U13245 (N_13245,N_13026,N_13055);
and U13246 (N_13246,N_13171,N_13122);
or U13247 (N_13247,N_13010,N_13002);
nand U13248 (N_13248,N_13155,N_13056);
nor U13249 (N_13249,N_13037,N_13180);
and U13250 (N_13250,N_13076,N_13006);
nor U13251 (N_13251,N_13019,N_13148);
nor U13252 (N_13252,N_13105,N_13187);
or U13253 (N_13253,N_13166,N_13139);
xnor U13254 (N_13254,N_13067,N_13068);
xor U13255 (N_13255,N_13020,N_13043);
xnor U13256 (N_13256,N_13031,N_13013);
xnor U13257 (N_13257,N_13061,N_13179);
and U13258 (N_13258,N_13085,N_13173);
or U13259 (N_13259,N_13095,N_13185);
and U13260 (N_13260,N_13091,N_13133);
xnor U13261 (N_13261,N_13127,N_13124);
nand U13262 (N_13262,N_13063,N_13093);
xnor U13263 (N_13263,N_13178,N_13084);
and U13264 (N_13264,N_13028,N_13098);
and U13265 (N_13265,N_13071,N_13197);
nor U13266 (N_13266,N_13131,N_13001);
nor U13267 (N_13267,N_13167,N_13096);
nand U13268 (N_13268,N_13069,N_13099);
nor U13269 (N_13269,N_13149,N_13027);
nor U13270 (N_13270,N_13081,N_13154);
xnor U13271 (N_13271,N_13112,N_13109);
and U13272 (N_13272,N_13136,N_13024);
or U13273 (N_13273,N_13097,N_13021);
xor U13274 (N_13274,N_13088,N_13005);
nor U13275 (N_13275,N_13003,N_13101);
or U13276 (N_13276,N_13049,N_13141);
or U13277 (N_13277,N_13116,N_13162);
nor U13278 (N_13278,N_13092,N_13151);
nand U13279 (N_13279,N_13082,N_13114);
or U13280 (N_13280,N_13186,N_13146);
nand U13281 (N_13281,N_13062,N_13130);
or U13282 (N_13282,N_13040,N_13117);
xor U13283 (N_13283,N_13192,N_13174);
nand U13284 (N_13284,N_13194,N_13079);
xor U13285 (N_13285,N_13072,N_13111);
and U13286 (N_13286,N_13110,N_13134);
nand U13287 (N_13287,N_13128,N_13059);
nand U13288 (N_13288,N_13046,N_13195);
and U13289 (N_13289,N_13023,N_13012);
or U13290 (N_13290,N_13036,N_13172);
xnor U13291 (N_13291,N_13032,N_13034);
nand U13292 (N_13292,N_13182,N_13089);
nand U13293 (N_13293,N_13065,N_13074);
and U13294 (N_13294,N_13175,N_13033);
or U13295 (N_13295,N_13014,N_13107);
nor U13296 (N_13296,N_13165,N_13070);
or U13297 (N_13297,N_13060,N_13078);
nor U13298 (N_13298,N_13158,N_13094);
xnor U13299 (N_13299,N_13132,N_13190);
nor U13300 (N_13300,N_13195,N_13187);
or U13301 (N_13301,N_13056,N_13084);
and U13302 (N_13302,N_13155,N_13093);
or U13303 (N_13303,N_13167,N_13124);
or U13304 (N_13304,N_13057,N_13026);
and U13305 (N_13305,N_13076,N_13115);
xnor U13306 (N_13306,N_13086,N_13131);
nand U13307 (N_13307,N_13097,N_13119);
xor U13308 (N_13308,N_13141,N_13159);
and U13309 (N_13309,N_13132,N_13034);
and U13310 (N_13310,N_13101,N_13030);
nor U13311 (N_13311,N_13089,N_13132);
or U13312 (N_13312,N_13055,N_13148);
nand U13313 (N_13313,N_13154,N_13044);
or U13314 (N_13314,N_13176,N_13154);
nor U13315 (N_13315,N_13024,N_13142);
nor U13316 (N_13316,N_13042,N_13116);
and U13317 (N_13317,N_13040,N_13043);
and U13318 (N_13318,N_13008,N_13059);
nand U13319 (N_13319,N_13137,N_13040);
nand U13320 (N_13320,N_13108,N_13190);
nand U13321 (N_13321,N_13136,N_13087);
nand U13322 (N_13322,N_13057,N_13110);
nand U13323 (N_13323,N_13035,N_13027);
and U13324 (N_13324,N_13197,N_13085);
or U13325 (N_13325,N_13141,N_13132);
xnor U13326 (N_13326,N_13069,N_13165);
nand U13327 (N_13327,N_13021,N_13162);
nand U13328 (N_13328,N_13077,N_13185);
and U13329 (N_13329,N_13105,N_13052);
and U13330 (N_13330,N_13058,N_13194);
nor U13331 (N_13331,N_13065,N_13068);
nor U13332 (N_13332,N_13006,N_13111);
and U13333 (N_13333,N_13165,N_13101);
xnor U13334 (N_13334,N_13149,N_13148);
nor U13335 (N_13335,N_13068,N_13175);
or U13336 (N_13336,N_13060,N_13033);
and U13337 (N_13337,N_13189,N_13198);
and U13338 (N_13338,N_13185,N_13045);
nand U13339 (N_13339,N_13125,N_13162);
and U13340 (N_13340,N_13182,N_13137);
nor U13341 (N_13341,N_13147,N_13063);
and U13342 (N_13342,N_13154,N_13042);
nor U13343 (N_13343,N_13132,N_13072);
or U13344 (N_13344,N_13082,N_13067);
nand U13345 (N_13345,N_13087,N_13197);
nand U13346 (N_13346,N_13117,N_13069);
xnor U13347 (N_13347,N_13025,N_13164);
and U13348 (N_13348,N_13058,N_13193);
nand U13349 (N_13349,N_13073,N_13056);
nor U13350 (N_13350,N_13138,N_13172);
or U13351 (N_13351,N_13011,N_13102);
or U13352 (N_13352,N_13087,N_13133);
nand U13353 (N_13353,N_13099,N_13022);
nor U13354 (N_13354,N_13171,N_13008);
nor U13355 (N_13355,N_13108,N_13137);
xnor U13356 (N_13356,N_13010,N_13110);
or U13357 (N_13357,N_13009,N_13198);
nand U13358 (N_13358,N_13043,N_13113);
xnor U13359 (N_13359,N_13106,N_13199);
xor U13360 (N_13360,N_13183,N_13040);
or U13361 (N_13361,N_13010,N_13150);
nand U13362 (N_13362,N_13071,N_13142);
nand U13363 (N_13363,N_13029,N_13123);
nand U13364 (N_13364,N_13106,N_13135);
nand U13365 (N_13365,N_13160,N_13084);
or U13366 (N_13366,N_13062,N_13170);
or U13367 (N_13367,N_13103,N_13114);
nor U13368 (N_13368,N_13142,N_13177);
nor U13369 (N_13369,N_13008,N_13161);
xnor U13370 (N_13370,N_13015,N_13192);
and U13371 (N_13371,N_13194,N_13054);
nor U13372 (N_13372,N_13125,N_13128);
nor U13373 (N_13373,N_13191,N_13179);
nor U13374 (N_13374,N_13031,N_13068);
nor U13375 (N_13375,N_13199,N_13198);
and U13376 (N_13376,N_13085,N_13195);
nand U13377 (N_13377,N_13091,N_13173);
or U13378 (N_13378,N_13193,N_13031);
nand U13379 (N_13379,N_13038,N_13124);
nor U13380 (N_13380,N_13110,N_13072);
nand U13381 (N_13381,N_13087,N_13147);
nor U13382 (N_13382,N_13126,N_13002);
xor U13383 (N_13383,N_13182,N_13107);
or U13384 (N_13384,N_13163,N_13154);
or U13385 (N_13385,N_13048,N_13191);
and U13386 (N_13386,N_13139,N_13113);
or U13387 (N_13387,N_13088,N_13078);
nor U13388 (N_13388,N_13033,N_13193);
nand U13389 (N_13389,N_13169,N_13052);
xnor U13390 (N_13390,N_13168,N_13059);
or U13391 (N_13391,N_13104,N_13180);
or U13392 (N_13392,N_13140,N_13099);
nor U13393 (N_13393,N_13043,N_13188);
nor U13394 (N_13394,N_13059,N_13049);
or U13395 (N_13395,N_13018,N_13000);
or U13396 (N_13396,N_13054,N_13069);
or U13397 (N_13397,N_13190,N_13128);
and U13398 (N_13398,N_13193,N_13034);
or U13399 (N_13399,N_13164,N_13050);
nor U13400 (N_13400,N_13356,N_13292);
nor U13401 (N_13401,N_13209,N_13334);
nor U13402 (N_13402,N_13287,N_13311);
nand U13403 (N_13403,N_13343,N_13310);
and U13404 (N_13404,N_13251,N_13390);
xnor U13405 (N_13405,N_13276,N_13346);
and U13406 (N_13406,N_13312,N_13229);
nor U13407 (N_13407,N_13262,N_13329);
or U13408 (N_13408,N_13246,N_13241);
xnor U13409 (N_13409,N_13375,N_13270);
nor U13410 (N_13410,N_13374,N_13323);
xor U13411 (N_13411,N_13217,N_13285);
or U13412 (N_13412,N_13349,N_13252);
nand U13413 (N_13413,N_13378,N_13392);
nand U13414 (N_13414,N_13273,N_13244);
and U13415 (N_13415,N_13250,N_13382);
and U13416 (N_13416,N_13353,N_13279);
and U13417 (N_13417,N_13361,N_13377);
and U13418 (N_13418,N_13372,N_13274);
nor U13419 (N_13419,N_13219,N_13260);
nand U13420 (N_13420,N_13326,N_13317);
and U13421 (N_13421,N_13302,N_13315);
or U13422 (N_13422,N_13322,N_13298);
nor U13423 (N_13423,N_13271,N_13380);
xor U13424 (N_13424,N_13210,N_13218);
or U13425 (N_13425,N_13389,N_13247);
nor U13426 (N_13426,N_13257,N_13320);
and U13427 (N_13427,N_13367,N_13242);
xnor U13428 (N_13428,N_13245,N_13370);
or U13429 (N_13429,N_13300,N_13280);
nor U13430 (N_13430,N_13297,N_13254);
xnor U13431 (N_13431,N_13284,N_13200);
nand U13432 (N_13432,N_13253,N_13202);
or U13433 (N_13433,N_13266,N_13396);
nand U13434 (N_13434,N_13363,N_13395);
nand U13435 (N_13435,N_13385,N_13272);
nand U13436 (N_13436,N_13319,N_13358);
or U13437 (N_13437,N_13327,N_13314);
or U13438 (N_13438,N_13340,N_13359);
xnor U13439 (N_13439,N_13376,N_13208);
xor U13440 (N_13440,N_13211,N_13325);
or U13441 (N_13441,N_13296,N_13240);
and U13442 (N_13442,N_13345,N_13335);
xor U13443 (N_13443,N_13336,N_13386);
and U13444 (N_13444,N_13225,N_13399);
nand U13445 (N_13445,N_13291,N_13239);
or U13446 (N_13446,N_13351,N_13206);
nand U13447 (N_13447,N_13234,N_13201);
nor U13448 (N_13448,N_13379,N_13255);
xor U13449 (N_13449,N_13277,N_13350);
nor U13450 (N_13450,N_13313,N_13224);
xnor U13451 (N_13451,N_13235,N_13393);
nand U13452 (N_13452,N_13331,N_13293);
xnor U13453 (N_13453,N_13364,N_13337);
xnor U13454 (N_13454,N_13223,N_13330);
nand U13455 (N_13455,N_13268,N_13258);
and U13456 (N_13456,N_13221,N_13230);
xnor U13457 (N_13457,N_13263,N_13283);
nor U13458 (N_13458,N_13352,N_13204);
xor U13459 (N_13459,N_13299,N_13397);
and U13460 (N_13460,N_13339,N_13308);
or U13461 (N_13461,N_13354,N_13233);
nand U13462 (N_13462,N_13215,N_13324);
xnor U13463 (N_13463,N_13342,N_13387);
nand U13464 (N_13464,N_13394,N_13341);
nand U13465 (N_13465,N_13303,N_13214);
and U13466 (N_13466,N_13290,N_13309);
or U13467 (N_13467,N_13355,N_13316);
nand U13468 (N_13468,N_13371,N_13226);
nand U13469 (N_13469,N_13321,N_13231);
nand U13470 (N_13470,N_13338,N_13212);
nand U13471 (N_13471,N_13348,N_13304);
xor U13472 (N_13472,N_13373,N_13332);
xnor U13473 (N_13473,N_13237,N_13318);
xor U13474 (N_13474,N_13301,N_13227);
and U13475 (N_13475,N_13391,N_13357);
xor U13476 (N_13476,N_13360,N_13295);
nand U13477 (N_13477,N_13243,N_13222);
or U13478 (N_13478,N_13269,N_13366);
or U13479 (N_13479,N_13281,N_13388);
xor U13480 (N_13480,N_13220,N_13278);
nand U13481 (N_13481,N_13282,N_13267);
nand U13482 (N_13482,N_13236,N_13232);
xor U13483 (N_13483,N_13368,N_13207);
nand U13484 (N_13484,N_13203,N_13256);
xor U13485 (N_13485,N_13306,N_13286);
nor U13486 (N_13486,N_13383,N_13384);
nor U13487 (N_13487,N_13216,N_13307);
xor U13488 (N_13488,N_13249,N_13213);
and U13489 (N_13489,N_13261,N_13344);
xor U13490 (N_13490,N_13369,N_13238);
xor U13491 (N_13491,N_13288,N_13381);
and U13492 (N_13492,N_13264,N_13259);
nor U13493 (N_13493,N_13328,N_13248);
and U13494 (N_13494,N_13228,N_13333);
or U13495 (N_13495,N_13398,N_13362);
or U13496 (N_13496,N_13347,N_13205);
xnor U13497 (N_13497,N_13294,N_13265);
and U13498 (N_13498,N_13365,N_13275);
nor U13499 (N_13499,N_13289,N_13305);
nor U13500 (N_13500,N_13332,N_13277);
nor U13501 (N_13501,N_13222,N_13368);
or U13502 (N_13502,N_13222,N_13256);
nand U13503 (N_13503,N_13305,N_13273);
and U13504 (N_13504,N_13345,N_13300);
and U13505 (N_13505,N_13239,N_13320);
nor U13506 (N_13506,N_13376,N_13369);
and U13507 (N_13507,N_13209,N_13305);
xor U13508 (N_13508,N_13251,N_13276);
nand U13509 (N_13509,N_13222,N_13274);
nor U13510 (N_13510,N_13318,N_13343);
or U13511 (N_13511,N_13205,N_13303);
nand U13512 (N_13512,N_13285,N_13366);
or U13513 (N_13513,N_13395,N_13329);
and U13514 (N_13514,N_13230,N_13345);
nor U13515 (N_13515,N_13283,N_13394);
xnor U13516 (N_13516,N_13317,N_13365);
nor U13517 (N_13517,N_13348,N_13391);
nor U13518 (N_13518,N_13204,N_13228);
nor U13519 (N_13519,N_13346,N_13350);
and U13520 (N_13520,N_13317,N_13233);
xor U13521 (N_13521,N_13338,N_13364);
and U13522 (N_13522,N_13360,N_13339);
nand U13523 (N_13523,N_13264,N_13288);
and U13524 (N_13524,N_13375,N_13250);
xor U13525 (N_13525,N_13357,N_13203);
nand U13526 (N_13526,N_13269,N_13281);
or U13527 (N_13527,N_13332,N_13243);
nor U13528 (N_13528,N_13272,N_13234);
and U13529 (N_13529,N_13324,N_13227);
nor U13530 (N_13530,N_13270,N_13399);
and U13531 (N_13531,N_13305,N_13384);
or U13532 (N_13532,N_13235,N_13356);
and U13533 (N_13533,N_13247,N_13386);
xnor U13534 (N_13534,N_13277,N_13247);
xnor U13535 (N_13535,N_13238,N_13328);
nor U13536 (N_13536,N_13342,N_13204);
and U13537 (N_13537,N_13257,N_13287);
xnor U13538 (N_13538,N_13393,N_13298);
xnor U13539 (N_13539,N_13284,N_13216);
or U13540 (N_13540,N_13386,N_13215);
or U13541 (N_13541,N_13280,N_13308);
nand U13542 (N_13542,N_13372,N_13245);
or U13543 (N_13543,N_13329,N_13217);
nor U13544 (N_13544,N_13200,N_13274);
xnor U13545 (N_13545,N_13263,N_13244);
nor U13546 (N_13546,N_13375,N_13388);
nor U13547 (N_13547,N_13364,N_13240);
nand U13548 (N_13548,N_13245,N_13378);
xor U13549 (N_13549,N_13228,N_13292);
nor U13550 (N_13550,N_13238,N_13271);
nand U13551 (N_13551,N_13396,N_13211);
and U13552 (N_13552,N_13294,N_13395);
nor U13553 (N_13553,N_13306,N_13329);
nor U13554 (N_13554,N_13245,N_13299);
nor U13555 (N_13555,N_13323,N_13392);
or U13556 (N_13556,N_13317,N_13347);
nand U13557 (N_13557,N_13362,N_13291);
and U13558 (N_13558,N_13244,N_13296);
or U13559 (N_13559,N_13288,N_13367);
or U13560 (N_13560,N_13209,N_13294);
nand U13561 (N_13561,N_13264,N_13394);
nand U13562 (N_13562,N_13344,N_13269);
or U13563 (N_13563,N_13389,N_13280);
and U13564 (N_13564,N_13205,N_13265);
nand U13565 (N_13565,N_13319,N_13398);
and U13566 (N_13566,N_13365,N_13345);
nand U13567 (N_13567,N_13360,N_13302);
nand U13568 (N_13568,N_13308,N_13382);
xor U13569 (N_13569,N_13207,N_13382);
or U13570 (N_13570,N_13318,N_13377);
and U13571 (N_13571,N_13337,N_13334);
nor U13572 (N_13572,N_13386,N_13314);
nor U13573 (N_13573,N_13258,N_13395);
and U13574 (N_13574,N_13341,N_13270);
or U13575 (N_13575,N_13315,N_13388);
nor U13576 (N_13576,N_13393,N_13224);
xnor U13577 (N_13577,N_13228,N_13399);
xor U13578 (N_13578,N_13254,N_13312);
nand U13579 (N_13579,N_13282,N_13279);
xor U13580 (N_13580,N_13284,N_13322);
nor U13581 (N_13581,N_13337,N_13239);
xnor U13582 (N_13582,N_13281,N_13380);
or U13583 (N_13583,N_13313,N_13255);
or U13584 (N_13584,N_13253,N_13239);
nand U13585 (N_13585,N_13259,N_13354);
or U13586 (N_13586,N_13222,N_13321);
nor U13587 (N_13587,N_13307,N_13367);
nor U13588 (N_13588,N_13396,N_13321);
or U13589 (N_13589,N_13353,N_13209);
or U13590 (N_13590,N_13399,N_13345);
and U13591 (N_13591,N_13350,N_13204);
nand U13592 (N_13592,N_13395,N_13225);
nor U13593 (N_13593,N_13298,N_13253);
nor U13594 (N_13594,N_13233,N_13373);
xor U13595 (N_13595,N_13251,N_13317);
and U13596 (N_13596,N_13367,N_13247);
nor U13597 (N_13597,N_13288,N_13246);
and U13598 (N_13598,N_13318,N_13261);
nor U13599 (N_13599,N_13387,N_13240);
and U13600 (N_13600,N_13595,N_13487);
nor U13601 (N_13601,N_13550,N_13587);
or U13602 (N_13602,N_13574,N_13483);
or U13603 (N_13603,N_13422,N_13521);
nand U13604 (N_13604,N_13592,N_13533);
xor U13605 (N_13605,N_13453,N_13529);
xor U13606 (N_13606,N_13412,N_13423);
or U13607 (N_13607,N_13551,N_13534);
xnor U13608 (N_13608,N_13447,N_13597);
nand U13609 (N_13609,N_13593,N_13434);
or U13610 (N_13610,N_13584,N_13465);
nor U13611 (N_13611,N_13490,N_13576);
nor U13612 (N_13612,N_13589,N_13572);
xnor U13613 (N_13613,N_13579,N_13508);
and U13614 (N_13614,N_13520,N_13558);
xor U13615 (N_13615,N_13421,N_13485);
nor U13616 (N_13616,N_13457,N_13401);
nand U13617 (N_13617,N_13569,N_13435);
and U13618 (N_13618,N_13492,N_13438);
or U13619 (N_13619,N_13556,N_13578);
nor U13620 (N_13620,N_13429,N_13524);
nand U13621 (N_13621,N_13583,N_13460);
nand U13622 (N_13622,N_13507,N_13498);
or U13623 (N_13623,N_13479,N_13446);
or U13624 (N_13624,N_13542,N_13528);
nor U13625 (N_13625,N_13462,N_13505);
nor U13626 (N_13626,N_13437,N_13568);
nand U13627 (N_13627,N_13486,N_13552);
nand U13628 (N_13628,N_13445,N_13458);
and U13629 (N_13629,N_13439,N_13580);
or U13630 (N_13630,N_13459,N_13428);
nor U13631 (N_13631,N_13554,N_13530);
nand U13632 (N_13632,N_13469,N_13413);
or U13633 (N_13633,N_13594,N_13563);
nor U13634 (N_13634,N_13436,N_13567);
nor U13635 (N_13635,N_13561,N_13588);
xor U13636 (N_13636,N_13535,N_13596);
and U13637 (N_13637,N_13514,N_13400);
nor U13638 (N_13638,N_13450,N_13405);
nor U13639 (N_13639,N_13546,N_13482);
xor U13640 (N_13640,N_13471,N_13553);
xnor U13641 (N_13641,N_13454,N_13577);
or U13642 (N_13642,N_13491,N_13461);
and U13643 (N_13643,N_13484,N_13590);
or U13644 (N_13644,N_13493,N_13506);
or U13645 (N_13645,N_13463,N_13502);
or U13646 (N_13646,N_13557,N_13455);
and U13647 (N_13647,N_13476,N_13545);
nor U13648 (N_13648,N_13473,N_13424);
xor U13649 (N_13649,N_13411,N_13420);
nor U13650 (N_13650,N_13573,N_13407);
nand U13651 (N_13651,N_13494,N_13430);
or U13652 (N_13652,N_13559,N_13562);
nor U13653 (N_13653,N_13467,N_13544);
nor U13654 (N_13654,N_13495,N_13539);
nand U13655 (N_13655,N_13477,N_13409);
and U13656 (N_13656,N_13517,N_13503);
or U13657 (N_13657,N_13523,N_13488);
nor U13658 (N_13658,N_13541,N_13540);
and U13659 (N_13659,N_13598,N_13575);
nor U13660 (N_13660,N_13526,N_13451);
nor U13661 (N_13661,N_13418,N_13481);
and U13662 (N_13662,N_13527,N_13555);
or U13663 (N_13663,N_13504,N_13415);
nand U13664 (N_13664,N_13472,N_13496);
and U13665 (N_13665,N_13432,N_13549);
nor U13666 (N_13666,N_13591,N_13410);
and U13667 (N_13667,N_13509,N_13499);
nand U13668 (N_13668,N_13442,N_13443);
nand U13669 (N_13669,N_13403,N_13532);
and U13670 (N_13670,N_13543,N_13433);
and U13671 (N_13671,N_13525,N_13513);
xnor U13672 (N_13672,N_13474,N_13475);
nand U13673 (N_13673,N_13489,N_13468);
nand U13674 (N_13674,N_13441,N_13571);
xnor U13675 (N_13675,N_13464,N_13512);
or U13676 (N_13676,N_13516,N_13497);
xnor U13677 (N_13677,N_13466,N_13444);
nor U13678 (N_13678,N_13564,N_13478);
and U13679 (N_13679,N_13406,N_13519);
nor U13680 (N_13680,N_13537,N_13538);
and U13681 (N_13681,N_13585,N_13511);
nor U13682 (N_13682,N_13548,N_13566);
nor U13683 (N_13683,N_13522,N_13531);
or U13684 (N_13684,N_13586,N_13480);
or U13685 (N_13685,N_13427,N_13515);
or U13686 (N_13686,N_13440,N_13581);
or U13687 (N_13687,N_13518,N_13547);
xnor U13688 (N_13688,N_13565,N_13570);
nand U13689 (N_13689,N_13448,N_13470);
xnor U13690 (N_13690,N_13452,N_13449);
nor U13691 (N_13691,N_13456,N_13500);
or U13692 (N_13692,N_13599,N_13501);
nor U13693 (N_13693,N_13416,N_13426);
or U13694 (N_13694,N_13536,N_13404);
or U13695 (N_13695,N_13417,N_13431);
nand U13696 (N_13696,N_13414,N_13560);
and U13697 (N_13697,N_13419,N_13408);
and U13698 (N_13698,N_13425,N_13402);
or U13699 (N_13699,N_13582,N_13510);
nor U13700 (N_13700,N_13506,N_13448);
and U13701 (N_13701,N_13542,N_13436);
xor U13702 (N_13702,N_13586,N_13483);
and U13703 (N_13703,N_13499,N_13517);
or U13704 (N_13704,N_13541,N_13504);
nand U13705 (N_13705,N_13507,N_13502);
xor U13706 (N_13706,N_13416,N_13540);
xnor U13707 (N_13707,N_13496,N_13501);
xor U13708 (N_13708,N_13571,N_13584);
nand U13709 (N_13709,N_13437,N_13590);
nor U13710 (N_13710,N_13496,N_13434);
xnor U13711 (N_13711,N_13501,N_13444);
and U13712 (N_13712,N_13582,N_13406);
and U13713 (N_13713,N_13430,N_13534);
nor U13714 (N_13714,N_13572,N_13524);
or U13715 (N_13715,N_13403,N_13481);
nand U13716 (N_13716,N_13443,N_13492);
nor U13717 (N_13717,N_13494,N_13523);
xnor U13718 (N_13718,N_13470,N_13435);
or U13719 (N_13719,N_13439,N_13512);
nand U13720 (N_13720,N_13521,N_13447);
or U13721 (N_13721,N_13491,N_13515);
and U13722 (N_13722,N_13536,N_13521);
xnor U13723 (N_13723,N_13591,N_13565);
nor U13724 (N_13724,N_13410,N_13455);
xor U13725 (N_13725,N_13525,N_13406);
nand U13726 (N_13726,N_13506,N_13417);
nor U13727 (N_13727,N_13516,N_13494);
and U13728 (N_13728,N_13573,N_13493);
nor U13729 (N_13729,N_13547,N_13510);
xor U13730 (N_13730,N_13488,N_13589);
nand U13731 (N_13731,N_13460,N_13553);
and U13732 (N_13732,N_13546,N_13569);
nor U13733 (N_13733,N_13464,N_13503);
nor U13734 (N_13734,N_13570,N_13415);
or U13735 (N_13735,N_13433,N_13406);
nand U13736 (N_13736,N_13454,N_13403);
nor U13737 (N_13737,N_13536,N_13570);
xor U13738 (N_13738,N_13539,N_13594);
nor U13739 (N_13739,N_13441,N_13536);
or U13740 (N_13740,N_13573,N_13487);
nand U13741 (N_13741,N_13536,N_13461);
nor U13742 (N_13742,N_13447,N_13446);
xnor U13743 (N_13743,N_13550,N_13558);
nand U13744 (N_13744,N_13568,N_13542);
and U13745 (N_13745,N_13590,N_13467);
or U13746 (N_13746,N_13491,N_13459);
xor U13747 (N_13747,N_13597,N_13533);
nor U13748 (N_13748,N_13432,N_13597);
nand U13749 (N_13749,N_13555,N_13440);
nand U13750 (N_13750,N_13461,N_13571);
or U13751 (N_13751,N_13474,N_13573);
or U13752 (N_13752,N_13518,N_13510);
or U13753 (N_13753,N_13474,N_13400);
nor U13754 (N_13754,N_13428,N_13483);
or U13755 (N_13755,N_13452,N_13466);
xnor U13756 (N_13756,N_13554,N_13518);
or U13757 (N_13757,N_13501,N_13512);
and U13758 (N_13758,N_13522,N_13452);
and U13759 (N_13759,N_13535,N_13593);
nor U13760 (N_13760,N_13436,N_13494);
nor U13761 (N_13761,N_13441,N_13567);
nor U13762 (N_13762,N_13433,N_13594);
and U13763 (N_13763,N_13403,N_13530);
and U13764 (N_13764,N_13434,N_13512);
and U13765 (N_13765,N_13521,N_13423);
and U13766 (N_13766,N_13582,N_13483);
nor U13767 (N_13767,N_13544,N_13434);
nand U13768 (N_13768,N_13537,N_13440);
or U13769 (N_13769,N_13468,N_13437);
xnor U13770 (N_13770,N_13579,N_13401);
xor U13771 (N_13771,N_13593,N_13559);
or U13772 (N_13772,N_13561,N_13487);
xor U13773 (N_13773,N_13418,N_13566);
nand U13774 (N_13774,N_13478,N_13579);
or U13775 (N_13775,N_13522,N_13567);
nor U13776 (N_13776,N_13498,N_13440);
nand U13777 (N_13777,N_13548,N_13428);
nand U13778 (N_13778,N_13492,N_13519);
nand U13779 (N_13779,N_13488,N_13401);
and U13780 (N_13780,N_13510,N_13415);
nand U13781 (N_13781,N_13585,N_13410);
nand U13782 (N_13782,N_13471,N_13547);
and U13783 (N_13783,N_13422,N_13498);
and U13784 (N_13784,N_13510,N_13460);
xor U13785 (N_13785,N_13584,N_13500);
or U13786 (N_13786,N_13594,N_13477);
xnor U13787 (N_13787,N_13472,N_13485);
nor U13788 (N_13788,N_13544,N_13493);
or U13789 (N_13789,N_13502,N_13491);
or U13790 (N_13790,N_13563,N_13417);
nand U13791 (N_13791,N_13470,N_13517);
nand U13792 (N_13792,N_13460,N_13478);
nand U13793 (N_13793,N_13419,N_13485);
or U13794 (N_13794,N_13544,N_13473);
xnor U13795 (N_13795,N_13555,N_13401);
nand U13796 (N_13796,N_13435,N_13469);
xnor U13797 (N_13797,N_13520,N_13446);
nor U13798 (N_13798,N_13418,N_13509);
and U13799 (N_13799,N_13418,N_13561);
xor U13800 (N_13800,N_13730,N_13753);
or U13801 (N_13801,N_13602,N_13729);
xnor U13802 (N_13802,N_13605,N_13751);
xor U13803 (N_13803,N_13625,N_13694);
and U13804 (N_13804,N_13709,N_13693);
nor U13805 (N_13805,N_13757,N_13610);
and U13806 (N_13806,N_13712,N_13669);
nand U13807 (N_13807,N_13628,N_13608);
xnor U13808 (N_13808,N_13711,N_13769);
xor U13809 (N_13809,N_13792,N_13738);
and U13810 (N_13810,N_13692,N_13786);
and U13811 (N_13811,N_13779,N_13773);
xor U13812 (N_13812,N_13687,N_13766);
or U13813 (N_13813,N_13667,N_13741);
or U13814 (N_13814,N_13781,N_13698);
nor U13815 (N_13815,N_13679,N_13629);
xor U13816 (N_13816,N_13641,N_13722);
xnor U13817 (N_13817,N_13622,N_13645);
xor U13818 (N_13818,N_13618,N_13714);
or U13819 (N_13819,N_13737,N_13656);
or U13820 (N_13820,N_13775,N_13765);
or U13821 (N_13821,N_13735,N_13674);
nand U13822 (N_13822,N_13724,N_13665);
and U13823 (N_13823,N_13604,N_13678);
nand U13824 (N_13824,N_13710,N_13655);
or U13825 (N_13825,N_13696,N_13739);
or U13826 (N_13826,N_13788,N_13721);
nand U13827 (N_13827,N_13783,N_13728);
and U13828 (N_13828,N_13770,N_13630);
and U13829 (N_13829,N_13725,N_13755);
and U13830 (N_13830,N_13791,N_13695);
nor U13831 (N_13831,N_13648,N_13774);
nor U13832 (N_13832,N_13671,N_13651);
and U13833 (N_13833,N_13603,N_13633);
and U13834 (N_13834,N_13746,N_13708);
or U13835 (N_13835,N_13606,N_13790);
nand U13836 (N_13836,N_13632,N_13657);
xnor U13837 (N_13837,N_13650,N_13713);
nand U13838 (N_13838,N_13756,N_13764);
and U13839 (N_13839,N_13750,N_13745);
xor U13840 (N_13840,N_13776,N_13705);
nor U13841 (N_13841,N_13703,N_13787);
nand U13842 (N_13842,N_13662,N_13672);
nand U13843 (N_13843,N_13706,N_13720);
nand U13844 (N_13844,N_13624,N_13626);
or U13845 (N_13845,N_13701,N_13620);
nand U13846 (N_13846,N_13771,N_13680);
and U13847 (N_13847,N_13675,N_13638);
nor U13848 (N_13848,N_13799,N_13600);
xor U13849 (N_13849,N_13707,N_13736);
and U13850 (N_13850,N_13748,N_13639);
xor U13851 (N_13851,N_13688,N_13697);
nor U13852 (N_13852,N_13691,N_13634);
and U13853 (N_13853,N_13683,N_13686);
or U13854 (N_13854,N_13752,N_13777);
and U13855 (N_13855,N_13663,N_13636);
or U13856 (N_13856,N_13785,N_13658);
and U13857 (N_13857,N_13740,N_13732);
or U13858 (N_13858,N_13616,N_13623);
and U13859 (N_13859,N_13798,N_13702);
nor U13860 (N_13860,N_13758,N_13609);
or U13861 (N_13861,N_13716,N_13761);
nand U13862 (N_13862,N_13733,N_13673);
nand U13863 (N_13863,N_13796,N_13653);
xor U13864 (N_13864,N_13778,N_13666);
and U13865 (N_13865,N_13619,N_13780);
nand U13866 (N_13866,N_13699,N_13644);
nor U13867 (N_13867,N_13642,N_13749);
or U13868 (N_13868,N_13744,N_13727);
and U13869 (N_13869,N_13760,N_13768);
nand U13870 (N_13870,N_13647,N_13654);
nor U13871 (N_13871,N_13685,N_13613);
or U13872 (N_13872,N_13617,N_13668);
xnor U13873 (N_13873,N_13637,N_13734);
or U13874 (N_13874,N_13700,N_13601);
and U13875 (N_13875,N_13607,N_13631);
xor U13876 (N_13876,N_13782,N_13797);
nand U13877 (N_13877,N_13754,N_13661);
or U13878 (N_13878,N_13793,N_13772);
nor U13879 (N_13879,N_13611,N_13742);
and U13880 (N_13880,N_13704,N_13640);
and U13881 (N_13881,N_13762,N_13684);
and U13882 (N_13882,N_13689,N_13643);
and U13883 (N_13883,N_13718,N_13767);
and U13884 (N_13884,N_13795,N_13726);
and U13885 (N_13885,N_13723,N_13763);
and U13886 (N_13886,N_13743,N_13670);
nand U13887 (N_13887,N_13652,N_13681);
or U13888 (N_13888,N_13717,N_13646);
and U13889 (N_13889,N_13664,N_13676);
nor U13890 (N_13890,N_13690,N_13615);
xnor U13891 (N_13891,N_13627,N_13660);
and U13892 (N_13892,N_13794,N_13659);
xnor U13893 (N_13893,N_13731,N_13789);
nand U13894 (N_13894,N_13715,N_13677);
nand U13895 (N_13895,N_13635,N_13614);
or U13896 (N_13896,N_13747,N_13649);
xor U13897 (N_13897,N_13612,N_13784);
nor U13898 (N_13898,N_13759,N_13682);
nand U13899 (N_13899,N_13719,N_13621);
nand U13900 (N_13900,N_13682,N_13706);
and U13901 (N_13901,N_13799,N_13722);
nor U13902 (N_13902,N_13601,N_13687);
nand U13903 (N_13903,N_13767,N_13634);
and U13904 (N_13904,N_13768,N_13641);
nand U13905 (N_13905,N_13733,N_13601);
nand U13906 (N_13906,N_13615,N_13696);
nor U13907 (N_13907,N_13665,N_13686);
xor U13908 (N_13908,N_13717,N_13643);
xnor U13909 (N_13909,N_13602,N_13751);
xor U13910 (N_13910,N_13691,N_13785);
nand U13911 (N_13911,N_13603,N_13684);
nand U13912 (N_13912,N_13792,N_13618);
nand U13913 (N_13913,N_13680,N_13636);
and U13914 (N_13914,N_13623,N_13641);
nor U13915 (N_13915,N_13672,N_13765);
nor U13916 (N_13916,N_13724,N_13622);
nor U13917 (N_13917,N_13765,N_13642);
nor U13918 (N_13918,N_13671,N_13654);
or U13919 (N_13919,N_13797,N_13657);
nor U13920 (N_13920,N_13790,N_13755);
nand U13921 (N_13921,N_13690,N_13774);
or U13922 (N_13922,N_13601,N_13654);
nand U13923 (N_13923,N_13601,N_13641);
or U13924 (N_13924,N_13641,N_13628);
xnor U13925 (N_13925,N_13662,N_13724);
or U13926 (N_13926,N_13785,N_13600);
and U13927 (N_13927,N_13758,N_13642);
and U13928 (N_13928,N_13708,N_13684);
or U13929 (N_13929,N_13663,N_13717);
or U13930 (N_13930,N_13607,N_13664);
and U13931 (N_13931,N_13702,N_13711);
nor U13932 (N_13932,N_13659,N_13706);
nor U13933 (N_13933,N_13679,N_13673);
or U13934 (N_13934,N_13750,N_13659);
and U13935 (N_13935,N_13699,N_13617);
and U13936 (N_13936,N_13799,N_13673);
nand U13937 (N_13937,N_13628,N_13621);
and U13938 (N_13938,N_13719,N_13765);
or U13939 (N_13939,N_13763,N_13659);
nor U13940 (N_13940,N_13799,N_13643);
and U13941 (N_13941,N_13782,N_13769);
nand U13942 (N_13942,N_13790,N_13777);
xnor U13943 (N_13943,N_13791,N_13607);
or U13944 (N_13944,N_13785,N_13638);
nand U13945 (N_13945,N_13763,N_13666);
xor U13946 (N_13946,N_13734,N_13665);
nand U13947 (N_13947,N_13798,N_13604);
xor U13948 (N_13948,N_13644,N_13716);
or U13949 (N_13949,N_13628,N_13684);
nor U13950 (N_13950,N_13755,N_13636);
nor U13951 (N_13951,N_13766,N_13792);
xnor U13952 (N_13952,N_13797,N_13647);
xor U13953 (N_13953,N_13741,N_13695);
xnor U13954 (N_13954,N_13647,N_13782);
or U13955 (N_13955,N_13638,N_13724);
nor U13956 (N_13956,N_13709,N_13675);
or U13957 (N_13957,N_13780,N_13672);
xnor U13958 (N_13958,N_13755,N_13680);
nor U13959 (N_13959,N_13756,N_13632);
and U13960 (N_13960,N_13723,N_13682);
nor U13961 (N_13961,N_13697,N_13652);
and U13962 (N_13962,N_13778,N_13775);
and U13963 (N_13963,N_13619,N_13664);
or U13964 (N_13964,N_13749,N_13785);
nand U13965 (N_13965,N_13644,N_13622);
nand U13966 (N_13966,N_13699,N_13730);
nor U13967 (N_13967,N_13753,N_13698);
nand U13968 (N_13968,N_13633,N_13775);
nor U13969 (N_13969,N_13789,N_13619);
nand U13970 (N_13970,N_13788,N_13799);
xor U13971 (N_13971,N_13799,N_13647);
nand U13972 (N_13972,N_13683,N_13707);
nor U13973 (N_13973,N_13677,N_13639);
or U13974 (N_13974,N_13750,N_13680);
and U13975 (N_13975,N_13669,N_13737);
and U13976 (N_13976,N_13786,N_13701);
or U13977 (N_13977,N_13669,N_13647);
and U13978 (N_13978,N_13629,N_13612);
nor U13979 (N_13979,N_13774,N_13607);
or U13980 (N_13980,N_13773,N_13694);
nand U13981 (N_13981,N_13633,N_13792);
or U13982 (N_13982,N_13736,N_13670);
and U13983 (N_13983,N_13666,N_13768);
and U13984 (N_13984,N_13738,N_13640);
or U13985 (N_13985,N_13656,N_13763);
or U13986 (N_13986,N_13787,N_13609);
nor U13987 (N_13987,N_13664,N_13691);
and U13988 (N_13988,N_13673,N_13691);
nor U13989 (N_13989,N_13721,N_13646);
xor U13990 (N_13990,N_13708,N_13782);
and U13991 (N_13991,N_13708,N_13730);
nand U13992 (N_13992,N_13615,N_13682);
and U13993 (N_13993,N_13799,N_13781);
nor U13994 (N_13994,N_13654,N_13609);
and U13995 (N_13995,N_13610,N_13775);
or U13996 (N_13996,N_13723,N_13653);
and U13997 (N_13997,N_13614,N_13629);
xor U13998 (N_13998,N_13789,N_13660);
or U13999 (N_13999,N_13767,N_13736);
or U14000 (N_14000,N_13939,N_13937);
or U14001 (N_14001,N_13954,N_13976);
xnor U14002 (N_14002,N_13858,N_13817);
nor U14003 (N_14003,N_13904,N_13820);
xor U14004 (N_14004,N_13964,N_13902);
and U14005 (N_14005,N_13984,N_13883);
xnor U14006 (N_14006,N_13982,N_13808);
and U14007 (N_14007,N_13860,N_13812);
xor U14008 (N_14008,N_13863,N_13877);
xor U14009 (N_14009,N_13862,N_13871);
and U14010 (N_14010,N_13920,N_13923);
xor U14011 (N_14011,N_13943,N_13850);
nor U14012 (N_14012,N_13844,N_13922);
nand U14013 (N_14013,N_13842,N_13809);
xor U14014 (N_14014,N_13806,N_13906);
or U14015 (N_14015,N_13991,N_13992);
nand U14016 (N_14016,N_13834,N_13886);
nor U14017 (N_14017,N_13872,N_13859);
nor U14018 (N_14018,N_13855,N_13905);
nand U14019 (N_14019,N_13876,N_13965);
or U14020 (N_14020,N_13831,N_13949);
nand U14021 (N_14021,N_13885,N_13951);
nor U14022 (N_14022,N_13967,N_13810);
or U14023 (N_14023,N_13802,N_13899);
nor U14024 (N_14024,N_13945,N_13924);
or U14025 (N_14025,N_13938,N_13837);
nand U14026 (N_14026,N_13933,N_13889);
nand U14027 (N_14027,N_13957,N_13926);
and U14028 (N_14028,N_13870,N_13856);
and U14029 (N_14029,N_13900,N_13921);
and U14030 (N_14030,N_13830,N_13960);
and U14031 (N_14031,N_13878,N_13804);
or U14032 (N_14032,N_13910,N_13998);
nor U14033 (N_14033,N_13931,N_13890);
nand U14034 (N_14034,N_13917,N_13981);
or U14035 (N_14035,N_13866,N_13935);
and U14036 (N_14036,N_13881,N_13819);
nor U14037 (N_14037,N_13973,N_13942);
nand U14038 (N_14038,N_13854,N_13907);
or U14039 (N_14039,N_13880,N_13891);
and U14040 (N_14040,N_13977,N_13823);
xnor U14041 (N_14041,N_13853,N_13800);
nand U14042 (N_14042,N_13829,N_13840);
nand U14043 (N_14043,N_13944,N_13827);
xor U14044 (N_14044,N_13887,N_13836);
xnor U14045 (N_14045,N_13959,N_13995);
nor U14046 (N_14046,N_13929,N_13974);
nand U14047 (N_14047,N_13822,N_13879);
nand U14048 (N_14048,N_13824,N_13861);
nand U14049 (N_14049,N_13961,N_13828);
nand U14050 (N_14050,N_13989,N_13898);
nand U14051 (N_14051,N_13952,N_13940);
xnor U14052 (N_14052,N_13803,N_13867);
xnor U14053 (N_14053,N_13845,N_13912);
or U14054 (N_14054,N_13970,N_13852);
xnor U14055 (N_14055,N_13956,N_13999);
nor U14056 (N_14056,N_13972,N_13930);
and U14057 (N_14057,N_13997,N_13915);
nand U14058 (N_14058,N_13848,N_13932);
and U14059 (N_14059,N_13847,N_13919);
nand U14060 (N_14060,N_13978,N_13941);
nand U14061 (N_14061,N_13821,N_13838);
or U14062 (N_14062,N_13893,N_13996);
or U14063 (N_14063,N_13963,N_13816);
or U14064 (N_14064,N_13841,N_13969);
nand U14065 (N_14065,N_13839,N_13927);
or U14066 (N_14066,N_13826,N_13925);
nor U14067 (N_14067,N_13990,N_13903);
nor U14068 (N_14068,N_13892,N_13993);
xnor U14069 (N_14069,N_13868,N_13869);
xor U14070 (N_14070,N_13936,N_13918);
and U14071 (N_14071,N_13911,N_13947);
nor U14072 (N_14072,N_13987,N_13864);
and U14073 (N_14073,N_13966,N_13994);
xnor U14074 (N_14074,N_13874,N_13843);
xnor U14075 (N_14075,N_13875,N_13986);
nor U14076 (N_14076,N_13897,N_13888);
nand U14077 (N_14077,N_13825,N_13980);
nor U14078 (N_14078,N_13873,N_13814);
or U14079 (N_14079,N_13913,N_13983);
nand U14080 (N_14080,N_13958,N_13832);
nor U14081 (N_14081,N_13948,N_13807);
nor U14082 (N_14082,N_13908,N_13857);
xor U14083 (N_14083,N_13985,N_13813);
nor U14084 (N_14084,N_13988,N_13894);
and U14085 (N_14085,N_13901,N_13895);
and U14086 (N_14086,N_13928,N_13818);
or U14087 (N_14087,N_13851,N_13979);
and U14088 (N_14088,N_13909,N_13946);
or U14089 (N_14089,N_13815,N_13811);
or U14090 (N_14090,N_13805,N_13971);
and U14091 (N_14091,N_13950,N_13882);
nand U14092 (N_14092,N_13849,N_13955);
nand U14093 (N_14093,N_13914,N_13833);
xnor U14094 (N_14094,N_13865,N_13975);
nor U14095 (N_14095,N_13884,N_13962);
or U14096 (N_14096,N_13801,N_13896);
nand U14097 (N_14097,N_13934,N_13916);
xnor U14098 (N_14098,N_13835,N_13968);
nand U14099 (N_14099,N_13846,N_13953);
nor U14100 (N_14100,N_13925,N_13818);
or U14101 (N_14101,N_13997,N_13923);
and U14102 (N_14102,N_13813,N_13965);
xor U14103 (N_14103,N_13868,N_13974);
and U14104 (N_14104,N_13825,N_13851);
nor U14105 (N_14105,N_13968,N_13941);
xnor U14106 (N_14106,N_13832,N_13862);
or U14107 (N_14107,N_13826,N_13940);
xor U14108 (N_14108,N_13990,N_13962);
xnor U14109 (N_14109,N_13851,N_13820);
nand U14110 (N_14110,N_13913,N_13961);
xnor U14111 (N_14111,N_13949,N_13868);
and U14112 (N_14112,N_13940,N_13931);
nor U14113 (N_14113,N_13840,N_13915);
xnor U14114 (N_14114,N_13923,N_13836);
xnor U14115 (N_14115,N_13855,N_13983);
nor U14116 (N_14116,N_13911,N_13812);
xnor U14117 (N_14117,N_13825,N_13946);
nor U14118 (N_14118,N_13907,N_13936);
or U14119 (N_14119,N_13811,N_13988);
and U14120 (N_14120,N_13837,N_13915);
and U14121 (N_14121,N_13901,N_13992);
or U14122 (N_14122,N_13893,N_13912);
nand U14123 (N_14123,N_13893,N_13879);
or U14124 (N_14124,N_13913,N_13984);
xor U14125 (N_14125,N_13899,N_13955);
nor U14126 (N_14126,N_13813,N_13927);
xor U14127 (N_14127,N_13821,N_13937);
xor U14128 (N_14128,N_13941,N_13870);
and U14129 (N_14129,N_13811,N_13987);
nor U14130 (N_14130,N_13873,N_13863);
nor U14131 (N_14131,N_13826,N_13968);
xor U14132 (N_14132,N_13904,N_13968);
nor U14133 (N_14133,N_13881,N_13855);
xor U14134 (N_14134,N_13832,N_13818);
and U14135 (N_14135,N_13956,N_13801);
or U14136 (N_14136,N_13952,N_13836);
nand U14137 (N_14137,N_13868,N_13981);
or U14138 (N_14138,N_13991,N_13843);
and U14139 (N_14139,N_13852,N_13992);
and U14140 (N_14140,N_13904,N_13967);
or U14141 (N_14141,N_13825,N_13970);
nor U14142 (N_14142,N_13841,N_13819);
and U14143 (N_14143,N_13932,N_13817);
nor U14144 (N_14144,N_13861,N_13911);
and U14145 (N_14145,N_13893,N_13801);
nor U14146 (N_14146,N_13924,N_13961);
xor U14147 (N_14147,N_13987,N_13945);
and U14148 (N_14148,N_13972,N_13906);
and U14149 (N_14149,N_13984,N_13863);
nand U14150 (N_14150,N_13906,N_13807);
nor U14151 (N_14151,N_13994,N_13990);
nand U14152 (N_14152,N_13910,N_13846);
and U14153 (N_14153,N_13894,N_13903);
nand U14154 (N_14154,N_13896,N_13910);
and U14155 (N_14155,N_13817,N_13895);
and U14156 (N_14156,N_13857,N_13979);
or U14157 (N_14157,N_13852,N_13869);
nand U14158 (N_14158,N_13825,N_13948);
nand U14159 (N_14159,N_13904,N_13911);
nor U14160 (N_14160,N_13880,N_13803);
and U14161 (N_14161,N_13998,N_13851);
and U14162 (N_14162,N_13920,N_13891);
nor U14163 (N_14163,N_13988,N_13996);
or U14164 (N_14164,N_13846,N_13907);
or U14165 (N_14165,N_13966,N_13828);
nand U14166 (N_14166,N_13820,N_13863);
and U14167 (N_14167,N_13995,N_13856);
nand U14168 (N_14168,N_13979,N_13944);
nor U14169 (N_14169,N_13813,N_13884);
and U14170 (N_14170,N_13977,N_13989);
xnor U14171 (N_14171,N_13917,N_13824);
xor U14172 (N_14172,N_13996,N_13810);
or U14173 (N_14173,N_13992,N_13853);
and U14174 (N_14174,N_13983,N_13886);
and U14175 (N_14175,N_13984,N_13875);
nor U14176 (N_14176,N_13941,N_13908);
nand U14177 (N_14177,N_13983,N_13874);
or U14178 (N_14178,N_13883,N_13804);
and U14179 (N_14179,N_13925,N_13845);
xor U14180 (N_14180,N_13850,N_13827);
and U14181 (N_14181,N_13938,N_13967);
or U14182 (N_14182,N_13929,N_13931);
nor U14183 (N_14183,N_13880,N_13941);
xor U14184 (N_14184,N_13954,N_13877);
or U14185 (N_14185,N_13870,N_13831);
xor U14186 (N_14186,N_13965,N_13845);
nand U14187 (N_14187,N_13885,N_13852);
or U14188 (N_14188,N_13947,N_13854);
xnor U14189 (N_14189,N_13904,N_13960);
xnor U14190 (N_14190,N_13866,N_13819);
or U14191 (N_14191,N_13993,N_13861);
xor U14192 (N_14192,N_13867,N_13842);
and U14193 (N_14193,N_13814,N_13832);
or U14194 (N_14194,N_13892,N_13862);
xnor U14195 (N_14195,N_13834,N_13997);
or U14196 (N_14196,N_13871,N_13986);
nand U14197 (N_14197,N_13889,N_13967);
nor U14198 (N_14198,N_13825,N_13840);
xor U14199 (N_14199,N_13973,N_13992);
nor U14200 (N_14200,N_14029,N_14009);
and U14201 (N_14201,N_14081,N_14174);
nor U14202 (N_14202,N_14013,N_14151);
nand U14203 (N_14203,N_14005,N_14026);
xnor U14204 (N_14204,N_14150,N_14032);
nand U14205 (N_14205,N_14078,N_14075);
or U14206 (N_14206,N_14071,N_14191);
xor U14207 (N_14207,N_14036,N_14055);
and U14208 (N_14208,N_14196,N_14061);
nor U14209 (N_14209,N_14126,N_14108);
and U14210 (N_14210,N_14084,N_14141);
or U14211 (N_14211,N_14004,N_14098);
or U14212 (N_14212,N_14116,N_14198);
xnor U14213 (N_14213,N_14040,N_14161);
and U14214 (N_14214,N_14158,N_14076);
nor U14215 (N_14215,N_14073,N_14169);
nor U14216 (N_14216,N_14090,N_14106);
and U14217 (N_14217,N_14007,N_14016);
or U14218 (N_14218,N_14143,N_14117);
nor U14219 (N_14219,N_14109,N_14102);
nand U14220 (N_14220,N_14012,N_14093);
or U14221 (N_14221,N_14164,N_14124);
xor U14222 (N_14222,N_14092,N_14027);
nor U14223 (N_14223,N_14064,N_14039);
xnor U14224 (N_14224,N_14068,N_14183);
and U14225 (N_14225,N_14030,N_14003);
and U14226 (N_14226,N_14031,N_14054);
and U14227 (N_14227,N_14085,N_14052);
nand U14228 (N_14228,N_14129,N_14080);
and U14229 (N_14229,N_14063,N_14144);
nor U14230 (N_14230,N_14065,N_14053);
or U14231 (N_14231,N_14096,N_14127);
nand U14232 (N_14232,N_14135,N_14179);
xnor U14233 (N_14233,N_14149,N_14067);
nand U14234 (N_14234,N_14033,N_14171);
and U14235 (N_14235,N_14056,N_14074);
and U14236 (N_14236,N_14022,N_14095);
nor U14237 (N_14237,N_14042,N_14172);
xnor U14238 (N_14238,N_14132,N_14062);
nand U14239 (N_14239,N_14111,N_14048);
nor U14240 (N_14240,N_14166,N_14023);
or U14241 (N_14241,N_14104,N_14131);
nand U14242 (N_14242,N_14180,N_14087);
and U14243 (N_14243,N_14066,N_14058);
nand U14244 (N_14244,N_14008,N_14120);
xor U14245 (N_14245,N_14178,N_14086);
nor U14246 (N_14246,N_14177,N_14189);
nand U14247 (N_14247,N_14100,N_14142);
or U14248 (N_14248,N_14049,N_14047);
or U14249 (N_14249,N_14186,N_14155);
xor U14250 (N_14250,N_14157,N_14193);
or U14251 (N_14251,N_14101,N_14014);
and U14252 (N_14252,N_14082,N_14148);
and U14253 (N_14253,N_14021,N_14188);
and U14254 (N_14254,N_14103,N_14165);
nand U14255 (N_14255,N_14197,N_14044);
or U14256 (N_14256,N_14043,N_14037);
and U14257 (N_14257,N_14114,N_14045);
nand U14258 (N_14258,N_14019,N_14105);
xor U14259 (N_14259,N_14028,N_14110);
nand U14260 (N_14260,N_14182,N_14025);
xor U14261 (N_14261,N_14118,N_14140);
and U14262 (N_14262,N_14162,N_14145);
xor U14263 (N_14263,N_14057,N_14112);
xor U14264 (N_14264,N_14097,N_14059);
xnor U14265 (N_14265,N_14195,N_14041);
nor U14266 (N_14266,N_14168,N_14185);
xor U14267 (N_14267,N_14156,N_14194);
nand U14268 (N_14268,N_14175,N_14160);
nand U14269 (N_14269,N_14035,N_14079);
nor U14270 (N_14270,N_14123,N_14113);
or U14271 (N_14271,N_14181,N_14015);
nor U14272 (N_14272,N_14011,N_14192);
and U14273 (N_14273,N_14147,N_14138);
xor U14274 (N_14274,N_14122,N_14077);
nor U14275 (N_14275,N_14034,N_14153);
nand U14276 (N_14276,N_14154,N_14069);
and U14277 (N_14277,N_14046,N_14094);
nor U14278 (N_14278,N_14006,N_14163);
xor U14279 (N_14279,N_14173,N_14167);
nand U14280 (N_14280,N_14002,N_14146);
xnor U14281 (N_14281,N_14017,N_14091);
xnor U14282 (N_14282,N_14024,N_14038);
or U14283 (N_14283,N_14128,N_14099);
or U14284 (N_14284,N_14115,N_14152);
or U14285 (N_14285,N_14139,N_14051);
or U14286 (N_14286,N_14133,N_14121);
nand U14287 (N_14287,N_14050,N_14083);
nand U14288 (N_14288,N_14072,N_14010);
nand U14289 (N_14289,N_14018,N_14136);
and U14290 (N_14290,N_14001,N_14089);
or U14291 (N_14291,N_14134,N_14187);
nor U14292 (N_14292,N_14088,N_14170);
xor U14293 (N_14293,N_14119,N_14199);
nand U14294 (N_14294,N_14107,N_14159);
nor U14295 (N_14295,N_14060,N_14020);
and U14296 (N_14296,N_14176,N_14130);
xor U14297 (N_14297,N_14184,N_14125);
or U14298 (N_14298,N_14190,N_14137);
or U14299 (N_14299,N_14000,N_14070);
and U14300 (N_14300,N_14006,N_14160);
or U14301 (N_14301,N_14081,N_14132);
xnor U14302 (N_14302,N_14169,N_14185);
and U14303 (N_14303,N_14112,N_14048);
xor U14304 (N_14304,N_14010,N_14033);
nor U14305 (N_14305,N_14015,N_14151);
and U14306 (N_14306,N_14056,N_14032);
and U14307 (N_14307,N_14085,N_14076);
nand U14308 (N_14308,N_14174,N_14091);
or U14309 (N_14309,N_14154,N_14047);
nor U14310 (N_14310,N_14098,N_14196);
and U14311 (N_14311,N_14084,N_14094);
nor U14312 (N_14312,N_14181,N_14174);
and U14313 (N_14313,N_14068,N_14158);
nor U14314 (N_14314,N_14178,N_14023);
nand U14315 (N_14315,N_14145,N_14090);
nor U14316 (N_14316,N_14114,N_14096);
nand U14317 (N_14317,N_14138,N_14196);
nor U14318 (N_14318,N_14157,N_14135);
xnor U14319 (N_14319,N_14146,N_14159);
nand U14320 (N_14320,N_14189,N_14092);
nand U14321 (N_14321,N_14152,N_14167);
or U14322 (N_14322,N_14064,N_14180);
nand U14323 (N_14323,N_14180,N_14175);
nand U14324 (N_14324,N_14108,N_14093);
and U14325 (N_14325,N_14178,N_14183);
xnor U14326 (N_14326,N_14196,N_14099);
xnor U14327 (N_14327,N_14101,N_14175);
and U14328 (N_14328,N_14090,N_14030);
xor U14329 (N_14329,N_14107,N_14050);
or U14330 (N_14330,N_14042,N_14170);
nor U14331 (N_14331,N_14144,N_14163);
nor U14332 (N_14332,N_14132,N_14106);
nor U14333 (N_14333,N_14124,N_14096);
nor U14334 (N_14334,N_14067,N_14141);
xnor U14335 (N_14335,N_14040,N_14197);
xor U14336 (N_14336,N_14108,N_14161);
xor U14337 (N_14337,N_14092,N_14080);
nand U14338 (N_14338,N_14086,N_14142);
nor U14339 (N_14339,N_14188,N_14163);
xor U14340 (N_14340,N_14150,N_14068);
or U14341 (N_14341,N_14110,N_14179);
nand U14342 (N_14342,N_14142,N_14155);
nor U14343 (N_14343,N_14120,N_14064);
or U14344 (N_14344,N_14103,N_14027);
nand U14345 (N_14345,N_14169,N_14188);
xor U14346 (N_14346,N_14199,N_14056);
or U14347 (N_14347,N_14004,N_14019);
and U14348 (N_14348,N_14020,N_14000);
xnor U14349 (N_14349,N_14077,N_14182);
and U14350 (N_14350,N_14131,N_14025);
and U14351 (N_14351,N_14096,N_14053);
xor U14352 (N_14352,N_14027,N_14156);
or U14353 (N_14353,N_14095,N_14059);
nand U14354 (N_14354,N_14039,N_14079);
xor U14355 (N_14355,N_14031,N_14187);
nor U14356 (N_14356,N_14105,N_14170);
nor U14357 (N_14357,N_14124,N_14008);
or U14358 (N_14358,N_14002,N_14173);
nand U14359 (N_14359,N_14099,N_14101);
nor U14360 (N_14360,N_14051,N_14178);
and U14361 (N_14361,N_14186,N_14141);
nor U14362 (N_14362,N_14152,N_14009);
or U14363 (N_14363,N_14015,N_14058);
xor U14364 (N_14364,N_14140,N_14182);
nand U14365 (N_14365,N_14045,N_14135);
nand U14366 (N_14366,N_14199,N_14035);
nor U14367 (N_14367,N_14172,N_14090);
xnor U14368 (N_14368,N_14024,N_14081);
or U14369 (N_14369,N_14131,N_14127);
xor U14370 (N_14370,N_14025,N_14066);
nand U14371 (N_14371,N_14196,N_14126);
nor U14372 (N_14372,N_14048,N_14005);
xor U14373 (N_14373,N_14101,N_14053);
nand U14374 (N_14374,N_14090,N_14083);
xor U14375 (N_14375,N_14128,N_14091);
nor U14376 (N_14376,N_14091,N_14185);
or U14377 (N_14377,N_14169,N_14013);
and U14378 (N_14378,N_14004,N_14074);
nand U14379 (N_14379,N_14135,N_14122);
or U14380 (N_14380,N_14166,N_14163);
nor U14381 (N_14381,N_14134,N_14041);
and U14382 (N_14382,N_14092,N_14030);
nand U14383 (N_14383,N_14189,N_14014);
and U14384 (N_14384,N_14169,N_14135);
nor U14385 (N_14385,N_14174,N_14194);
xor U14386 (N_14386,N_14170,N_14035);
and U14387 (N_14387,N_14190,N_14115);
xor U14388 (N_14388,N_14184,N_14095);
xor U14389 (N_14389,N_14193,N_14091);
nand U14390 (N_14390,N_14073,N_14090);
xnor U14391 (N_14391,N_14016,N_14061);
nand U14392 (N_14392,N_14112,N_14097);
xor U14393 (N_14393,N_14041,N_14109);
nor U14394 (N_14394,N_14010,N_14180);
or U14395 (N_14395,N_14156,N_14051);
nand U14396 (N_14396,N_14190,N_14077);
xnor U14397 (N_14397,N_14139,N_14022);
or U14398 (N_14398,N_14118,N_14072);
xor U14399 (N_14399,N_14021,N_14103);
or U14400 (N_14400,N_14333,N_14327);
or U14401 (N_14401,N_14245,N_14366);
nand U14402 (N_14402,N_14260,N_14362);
or U14403 (N_14403,N_14310,N_14301);
xor U14404 (N_14404,N_14321,N_14356);
or U14405 (N_14405,N_14300,N_14303);
and U14406 (N_14406,N_14374,N_14244);
nand U14407 (N_14407,N_14346,N_14288);
nor U14408 (N_14408,N_14391,N_14361);
nor U14409 (N_14409,N_14360,N_14250);
nor U14410 (N_14410,N_14287,N_14231);
and U14411 (N_14411,N_14225,N_14229);
xor U14412 (N_14412,N_14305,N_14282);
nand U14413 (N_14413,N_14240,N_14338);
xnor U14414 (N_14414,N_14398,N_14258);
nor U14415 (N_14415,N_14370,N_14389);
and U14416 (N_14416,N_14241,N_14378);
nor U14417 (N_14417,N_14239,N_14252);
nand U14418 (N_14418,N_14270,N_14236);
nand U14419 (N_14419,N_14213,N_14281);
nor U14420 (N_14420,N_14312,N_14266);
nor U14421 (N_14421,N_14347,N_14379);
or U14422 (N_14422,N_14284,N_14218);
nand U14423 (N_14423,N_14232,N_14326);
or U14424 (N_14424,N_14279,N_14291);
or U14425 (N_14425,N_14337,N_14259);
nand U14426 (N_14426,N_14324,N_14355);
or U14427 (N_14427,N_14304,N_14350);
nand U14428 (N_14428,N_14354,N_14399);
nor U14429 (N_14429,N_14221,N_14204);
or U14430 (N_14430,N_14383,N_14323);
or U14431 (N_14431,N_14271,N_14382);
and U14432 (N_14432,N_14249,N_14254);
xor U14433 (N_14433,N_14268,N_14214);
nand U14434 (N_14434,N_14344,N_14205);
xnor U14435 (N_14435,N_14216,N_14209);
nor U14436 (N_14436,N_14319,N_14377);
and U14437 (N_14437,N_14234,N_14299);
or U14438 (N_14438,N_14395,N_14207);
xnor U14439 (N_14439,N_14340,N_14336);
nor U14440 (N_14440,N_14325,N_14329);
or U14441 (N_14441,N_14373,N_14265);
and U14442 (N_14442,N_14330,N_14348);
xnor U14443 (N_14443,N_14210,N_14385);
or U14444 (N_14444,N_14211,N_14261);
xnor U14445 (N_14445,N_14369,N_14292);
nand U14446 (N_14446,N_14308,N_14313);
xnor U14447 (N_14447,N_14212,N_14215);
and U14448 (N_14448,N_14226,N_14248);
or U14449 (N_14449,N_14334,N_14298);
nor U14450 (N_14450,N_14311,N_14328);
and U14451 (N_14451,N_14372,N_14388);
nor U14452 (N_14452,N_14237,N_14256);
and U14453 (N_14453,N_14290,N_14243);
nor U14454 (N_14454,N_14387,N_14316);
nand U14455 (N_14455,N_14339,N_14341);
xnor U14456 (N_14456,N_14267,N_14320);
xor U14457 (N_14457,N_14233,N_14371);
nand U14458 (N_14458,N_14269,N_14368);
or U14459 (N_14459,N_14263,N_14314);
nor U14460 (N_14460,N_14295,N_14206);
xnor U14461 (N_14461,N_14381,N_14358);
nor U14462 (N_14462,N_14276,N_14217);
nor U14463 (N_14463,N_14247,N_14353);
xor U14464 (N_14464,N_14201,N_14365);
nand U14465 (N_14465,N_14309,N_14224);
or U14466 (N_14466,N_14296,N_14246);
nand U14467 (N_14467,N_14332,N_14202);
xnor U14468 (N_14468,N_14235,N_14200);
and U14469 (N_14469,N_14222,N_14384);
nand U14470 (N_14470,N_14335,N_14331);
and U14471 (N_14471,N_14390,N_14280);
and U14472 (N_14472,N_14357,N_14396);
xnor U14473 (N_14473,N_14285,N_14203);
and U14474 (N_14474,N_14275,N_14345);
and U14475 (N_14475,N_14317,N_14272);
nand U14476 (N_14476,N_14297,N_14318);
or U14477 (N_14477,N_14251,N_14283);
nor U14478 (N_14478,N_14278,N_14262);
xnor U14479 (N_14479,N_14349,N_14315);
and U14480 (N_14480,N_14273,N_14359);
or U14481 (N_14481,N_14255,N_14257);
xor U14482 (N_14482,N_14277,N_14230);
nor U14483 (N_14483,N_14264,N_14363);
xnor U14484 (N_14484,N_14228,N_14219);
and U14485 (N_14485,N_14238,N_14227);
xnor U14486 (N_14486,N_14343,N_14394);
or U14487 (N_14487,N_14375,N_14286);
nand U14488 (N_14488,N_14386,N_14289);
or U14489 (N_14489,N_14364,N_14274);
or U14490 (N_14490,N_14376,N_14223);
or U14491 (N_14491,N_14302,N_14293);
and U14492 (N_14492,N_14307,N_14294);
nand U14493 (N_14493,N_14352,N_14380);
and U14494 (N_14494,N_14253,N_14306);
or U14495 (N_14495,N_14342,N_14393);
nand U14496 (N_14496,N_14351,N_14397);
and U14497 (N_14497,N_14242,N_14392);
and U14498 (N_14498,N_14367,N_14220);
nand U14499 (N_14499,N_14322,N_14208);
xnor U14500 (N_14500,N_14374,N_14271);
nand U14501 (N_14501,N_14309,N_14282);
and U14502 (N_14502,N_14399,N_14321);
and U14503 (N_14503,N_14256,N_14383);
nand U14504 (N_14504,N_14368,N_14358);
nor U14505 (N_14505,N_14202,N_14302);
and U14506 (N_14506,N_14231,N_14300);
nor U14507 (N_14507,N_14239,N_14397);
nor U14508 (N_14508,N_14241,N_14213);
or U14509 (N_14509,N_14349,N_14244);
xor U14510 (N_14510,N_14316,N_14284);
nand U14511 (N_14511,N_14329,N_14287);
or U14512 (N_14512,N_14204,N_14345);
and U14513 (N_14513,N_14310,N_14387);
nor U14514 (N_14514,N_14213,N_14246);
xnor U14515 (N_14515,N_14373,N_14306);
xor U14516 (N_14516,N_14326,N_14371);
and U14517 (N_14517,N_14331,N_14342);
nand U14518 (N_14518,N_14204,N_14263);
nor U14519 (N_14519,N_14230,N_14336);
nand U14520 (N_14520,N_14301,N_14252);
xnor U14521 (N_14521,N_14313,N_14225);
xnor U14522 (N_14522,N_14291,N_14275);
nand U14523 (N_14523,N_14333,N_14229);
or U14524 (N_14524,N_14304,N_14289);
xor U14525 (N_14525,N_14289,N_14264);
or U14526 (N_14526,N_14348,N_14380);
and U14527 (N_14527,N_14342,N_14349);
xnor U14528 (N_14528,N_14361,N_14376);
nand U14529 (N_14529,N_14318,N_14381);
or U14530 (N_14530,N_14315,N_14384);
and U14531 (N_14531,N_14394,N_14350);
and U14532 (N_14532,N_14243,N_14359);
or U14533 (N_14533,N_14329,N_14379);
or U14534 (N_14534,N_14262,N_14225);
nand U14535 (N_14535,N_14223,N_14208);
nor U14536 (N_14536,N_14214,N_14270);
and U14537 (N_14537,N_14370,N_14247);
nand U14538 (N_14538,N_14279,N_14312);
nand U14539 (N_14539,N_14384,N_14373);
xor U14540 (N_14540,N_14249,N_14352);
nor U14541 (N_14541,N_14295,N_14237);
nor U14542 (N_14542,N_14312,N_14383);
or U14543 (N_14543,N_14228,N_14362);
nor U14544 (N_14544,N_14238,N_14205);
nand U14545 (N_14545,N_14213,N_14296);
nand U14546 (N_14546,N_14204,N_14331);
xnor U14547 (N_14547,N_14315,N_14280);
xnor U14548 (N_14548,N_14279,N_14394);
nand U14549 (N_14549,N_14241,N_14246);
nor U14550 (N_14550,N_14232,N_14210);
nor U14551 (N_14551,N_14269,N_14348);
nand U14552 (N_14552,N_14361,N_14314);
xor U14553 (N_14553,N_14236,N_14323);
xor U14554 (N_14554,N_14370,N_14240);
nand U14555 (N_14555,N_14274,N_14222);
or U14556 (N_14556,N_14225,N_14288);
and U14557 (N_14557,N_14374,N_14249);
or U14558 (N_14558,N_14317,N_14273);
nor U14559 (N_14559,N_14231,N_14322);
nor U14560 (N_14560,N_14203,N_14321);
and U14561 (N_14561,N_14246,N_14351);
nand U14562 (N_14562,N_14269,N_14385);
nor U14563 (N_14563,N_14294,N_14365);
nor U14564 (N_14564,N_14297,N_14240);
nand U14565 (N_14565,N_14379,N_14235);
and U14566 (N_14566,N_14203,N_14210);
and U14567 (N_14567,N_14358,N_14232);
xor U14568 (N_14568,N_14320,N_14251);
and U14569 (N_14569,N_14358,N_14394);
and U14570 (N_14570,N_14328,N_14248);
or U14571 (N_14571,N_14307,N_14245);
nor U14572 (N_14572,N_14209,N_14384);
and U14573 (N_14573,N_14302,N_14209);
nor U14574 (N_14574,N_14378,N_14242);
nor U14575 (N_14575,N_14324,N_14314);
nand U14576 (N_14576,N_14227,N_14307);
or U14577 (N_14577,N_14210,N_14380);
xor U14578 (N_14578,N_14370,N_14282);
or U14579 (N_14579,N_14249,N_14353);
or U14580 (N_14580,N_14364,N_14201);
xnor U14581 (N_14581,N_14218,N_14301);
or U14582 (N_14582,N_14283,N_14286);
or U14583 (N_14583,N_14398,N_14360);
and U14584 (N_14584,N_14278,N_14387);
nor U14585 (N_14585,N_14389,N_14378);
nand U14586 (N_14586,N_14216,N_14293);
nor U14587 (N_14587,N_14264,N_14387);
xnor U14588 (N_14588,N_14236,N_14366);
and U14589 (N_14589,N_14237,N_14223);
xor U14590 (N_14590,N_14337,N_14237);
xnor U14591 (N_14591,N_14208,N_14283);
nand U14592 (N_14592,N_14216,N_14336);
nor U14593 (N_14593,N_14279,N_14313);
or U14594 (N_14594,N_14225,N_14232);
nor U14595 (N_14595,N_14201,N_14284);
xor U14596 (N_14596,N_14367,N_14323);
and U14597 (N_14597,N_14393,N_14335);
xnor U14598 (N_14598,N_14348,N_14297);
and U14599 (N_14599,N_14241,N_14272);
and U14600 (N_14600,N_14520,N_14403);
or U14601 (N_14601,N_14479,N_14430);
or U14602 (N_14602,N_14507,N_14443);
nor U14603 (N_14603,N_14435,N_14491);
xnor U14604 (N_14604,N_14453,N_14501);
or U14605 (N_14605,N_14413,N_14431);
nand U14606 (N_14606,N_14547,N_14532);
or U14607 (N_14607,N_14508,N_14405);
and U14608 (N_14608,N_14425,N_14452);
nor U14609 (N_14609,N_14416,N_14462);
nor U14610 (N_14610,N_14559,N_14589);
or U14611 (N_14611,N_14423,N_14498);
nand U14612 (N_14612,N_14410,N_14455);
and U14613 (N_14613,N_14463,N_14546);
nor U14614 (N_14614,N_14527,N_14414);
and U14615 (N_14615,N_14480,N_14581);
and U14616 (N_14616,N_14468,N_14402);
xnor U14617 (N_14617,N_14499,N_14444);
nor U14618 (N_14618,N_14524,N_14580);
or U14619 (N_14619,N_14458,N_14556);
nand U14620 (N_14620,N_14436,N_14495);
xnor U14621 (N_14621,N_14449,N_14528);
nor U14622 (N_14622,N_14597,N_14534);
nor U14623 (N_14623,N_14418,N_14427);
nand U14624 (N_14624,N_14522,N_14471);
or U14625 (N_14625,N_14584,N_14486);
or U14626 (N_14626,N_14497,N_14407);
xor U14627 (N_14627,N_14561,N_14516);
xnor U14628 (N_14628,N_14485,N_14482);
xnor U14629 (N_14629,N_14529,N_14511);
and U14630 (N_14630,N_14473,N_14493);
xnor U14631 (N_14631,N_14563,N_14446);
xnor U14632 (N_14632,N_14437,N_14543);
nand U14633 (N_14633,N_14533,N_14577);
nor U14634 (N_14634,N_14417,N_14429);
or U14635 (N_14635,N_14445,N_14475);
nor U14636 (N_14636,N_14474,N_14494);
xor U14637 (N_14637,N_14510,N_14596);
nor U14638 (N_14638,N_14585,N_14448);
and U14639 (N_14639,N_14515,N_14464);
nand U14640 (N_14640,N_14588,N_14558);
or U14641 (N_14641,N_14582,N_14538);
and U14642 (N_14642,N_14566,N_14504);
and U14643 (N_14643,N_14487,N_14496);
or U14644 (N_14644,N_14573,N_14512);
and U14645 (N_14645,N_14579,N_14544);
xnor U14646 (N_14646,N_14426,N_14564);
nand U14647 (N_14647,N_14459,N_14574);
xnor U14648 (N_14648,N_14535,N_14412);
or U14649 (N_14649,N_14433,N_14409);
nor U14650 (N_14650,N_14441,N_14466);
nor U14651 (N_14651,N_14434,N_14583);
and U14652 (N_14652,N_14551,N_14470);
nand U14653 (N_14653,N_14484,N_14541);
xor U14654 (N_14654,N_14456,N_14531);
xor U14655 (N_14655,N_14525,N_14571);
or U14656 (N_14656,N_14472,N_14552);
and U14657 (N_14657,N_14505,N_14521);
and U14658 (N_14658,N_14545,N_14404);
and U14659 (N_14659,N_14595,N_14415);
nor U14660 (N_14660,N_14424,N_14461);
nand U14661 (N_14661,N_14549,N_14526);
nor U14662 (N_14662,N_14506,N_14518);
nor U14663 (N_14663,N_14509,N_14578);
nor U14664 (N_14664,N_14565,N_14478);
and U14665 (N_14665,N_14451,N_14587);
and U14666 (N_14666,N_14489,N_14592);
nor U14667 (N_14667,N_14557,N_14530);
and U14668 (N_14668,N_14465,N_14502);
nand U14669 (N_14669,N_14568,N_14590);
and U14670 (N_14670,N_14420,N_14490);
xnor U14671 (N_14671,N_14567,N_14569);
or U14672 (N_14672,N_14481,N_14598);
or U14673 (N_14673,N_14492,N_14439);
nor U14674 (N_14674,N_14553,N_14519);
and U14675 (N_14675,N_14457,N_14503);
xnor U14676 (N_14676,N_14406,N_14476);
nand U14677 (N_14677,N_14554,N_14517);
xor U14678 (N_14678,N_14539,N_14440);
or U14679 (N_14679,N_14523,N_14488);
xor U14680 (N_14680,N_14454,N_14483);
nor U14681 (N_14681,N_14548,N_14555);
xnor U14682 (N_14682,N_14593,N_14562);
xor U14683 (N_14683,N_14411,N_14477);
and U14684 (N_14684,N_14460,N_14428);
nor U14685 (N_14685,N_14432,N_14438);
and U14686 (N_14686,N_14576,N_14442);
and U14687 (N_14687,N_14421,N_14542);
xor U14688 (N_14688,N_14599,N_14560);
or U14689 (N_14689,N_14400,N_14419);
nor U14690 (N_14690,N_14572,N_14450);
nor U14691 (N_14691,N_14514,N_14570);
nand U14692 (N_14692,N_14540,N_14422);
or U14693 (N_14693,N_14550,N_14401);
xor U14694 (N_14694,N_14586,N_14447);
and U14695 (N_14695,N_14469,N_14537);
xor U14696 (N_14696,N_14594,N_14536);
xor U14697 (N_14697,N_14408,N_14575);
nand U14698 (N_14698,N_14591,N_14500);
or U14699 (N_14699,N_14513,N_14467);
and U14700 (N_14700,N_14412,N_14463);
nor U14701 (N_14701,N_14521,N_14450);
nor U14702 (N_14702,N_14524,N_14507);
and U14703 (N_14703,N_14429,N_14468);
nor U14704 (N_14704,N_14529,N_14567);
xor U14705 (N_14705,N_14510,N_14599);
xnor U14706 (N_14706,N_14520,N_14428);
nor U14707 (N_14707,N_14500,N_14454);
xor U14708 (N_14708,N_14531,N_14505);
xor U14709 (N_14709,N_14540,N_14586);
nand U14710 (N_14710,N_14575,N_14440);
nor U14711 (N_14711,N_14419,N_14580);
nor U14712 (N_14712,N_14558,N_14483);
or U14713 (N_14713,N_14558,N_14541);
xor U14714 (N_14714,N_14416,N_14473);
nor U14715 (N_14715,N_14407,N_14545);
or U14716 (N_14716,N_14463,N_14482);
or U14717 (N_14717,N_14518,N_14530);
xnor U14718 (N_14718,N_14599,N_14413);
nor U14719 (N_14719,N_14467,N_14468);
and U14720 (N_14720,N_14400,N_14401);
and U14721 (N_14721,N_14575,N_14475);
nor U14722 (N_14722,N_14518,N_14445);
nand U14723 (N_14723,N_14405,N_14529);
nor U14724 (N_14724,N_14467,N_14486);
nand U14725 (N_14725,N_14550,N_14500);
nand U14726 (N_14726,N_14471,N_14555);
nor U14727 (N_14727,N_14533,N_14554);
nand U14728 (N_14728,N_14513,N_14524);
nand U14729 (N_14729,N_14570,N_14551);
nor U14730 (N_14730,N_14486,N_14594);
nor U14731 (N_14731,N_14476,N_14486);
and U14732 (N_14732,N_14535,N_14461);
and U14733 (N_14733,N_14466,N_14495);
nor U14734 (N_14734,N_14415,N_14585);
and U14735 (N_14735,N_14406,N_14552);
nand U14736 (N_14736,N_14483,N_14523);
and U14737 (N_14737,N_14553,N_14541);
nand U14738 (N_14738,N_14545,N_14416);
nand U14739 (N_14739,N_14463,N_14573);
or U14740 (N_14740,N_14517,N_14473);
nor U14741 (N_14741,N_14426,N_14402);
and U14742 (N_14742,N_14440,N_14463);
or U14743 (N_14743,N_14470,N_14429);
nor U14744 (N_14744,N_14557,N_14495);
xnor U14745 (N_14745,N_14414,N_14488);
and U14746 (N_14746,N_14466,N_14434);
xor U14747 (N_14747,N_14597,N_14554);
xor U14748 (N_14748,N_14497,N_14413);
nor U14749 (N_14749,N_14524,N_14585);
nand U14750 (N_14750,N_14547,N_14582);
nand U14751 (N_14751,N_14540,N_14481);
xor U14752 (N_14752,N_14505,N_14510);
nand U14753 (N_14753,N_14545,N_14569);
or U14754 (N_14754,N_14560,N_14474);
nor U14755 (N_14755,N_14427,N_14439);
or U14756 (N_14756,N_14525,N_14469);
and U14757 (N_14757,N_14459,N_14561);
and U14758 (N_14758,N_14493,N_14563);
and U14759 (N_14759,N_14477,N_14526);
nand U14760 (N_14760,N_14579,N_14596);
xor U14761 (N_14761,N_14582,N_14463);
xor U14762 (N_14762,N_14565,N_14571);
nor U14763 (N_14763,N_14563,N_14480);
nor U14764 (N_14764,N_14561,N_14478);
nor U14765 (N_14765,N_14541,N_14490);
nand U14766 (N_14766,N_14574,N_14434);
xor U14767 (N_14767,N_14583,N_14495);
or U14768 (N_14768,N_14555,N_14411);
xor U14769 (N_14769,N_14519,N_14476);
xor U14770 (N_14770,N_14539,N_14516);
xor U14771 (N_14771,N_14442,N_14586);
nor U14772 (N_14772,N_14442,N_14484);
or U14773 (N_14773,N_14422,N_14463);
nor U14774 (N_14774,N_14451,N_14419);
and U14775 (N_14775,N_14418,N_14489);
nand U14776 (N_14776,N_14528,N_14470);
nor U14777 (N_14777,N_14498,N_14512);
or U14778 (N_14778,N_14570,N_14476);
nand U14779 (N_14779,N_14585,N_14431);
nor U14780 (N_14780,N_14458,N_14505);
xnor U14781 (N_14781,N_14401,N_14559);
and U14782 (N_14782,N_14594,N_14403);
xnor U14783 (N_14783,N_14409,N_14596);
or U14784 (N_14784,N_14565,N_14556);
nand U14785 (N_14785,N_14424,N_14422);
nor U14786 (N_14786,N_14508,N_14495);
nor U14787 (N_14787,N_14596,N_14555);
xor U14788 (N_14788,N_14456,N_14586);
or U14789 (N_14789,N_14516,N_14599);
nand U14790 (N_14790,N_14564,N_14441);
and U14791 (N_14791,N_14401,N_14520);
or U14792 (N_14792,N_14525,N_14411);
nor U14793 (N_14793,N_14577,N_14499);
xor U14794 (N_14794,N_14451,N_14555);
xnor U14795 (N_14795,N_14428,N_14445);
and U14796 (N_14796,N_14516,N_14484);
or U14797 (N_14797,N_14420,N_14532);
nor U14798 (N_14798,N_14435,N_14473);
xnor U14799 (N_14799,N_14508,N_14574);
nand U14800 (N_14800,N_14717,N_14655);
nor U14801 (N_14801,N_14721,N_14778);
or U14802 (N_14802,N_14705,N_14627);
nor U14803 (N_14803,N_14748,N_14790);
nor U14804 (N_14804,N_14641,N_14690);
nor U14805 (N_14805,N_14751,N_14729);
xnor U14806 (N_14806,N_14685,N_14648);
or U14807 (N_14807,N_14747,N_14724);
nand U14808 (N_14808,N_14638,N_14665);
or U14809 (N_14809,N_14640,N_14735);
xnor U14810 (N_14810,N_14743,N_14669);
or U14811 (N_14811,N_14770,N_14662);
and U14812 (N_14812,N_14712,N_14782);
or U14813 (N_14813,N_14642,N_14795);
or U14814 (N_14814,N_14773,N_14613);
nor U14815 (N_14815,N_14736,N_14737);
nand U14816 (N_14816,N_14785,N_14787);
nor U14817 (N_14817,N_14769,N_14749);
or U14818 (N_14818,N_14664,N_14723);
nor U14819 (N_14819,N_14606,N_14626);
nor U14820 (N_14820,N_14744,N_14754);
and U14821 (N_14821,N_14714,N_14651);
or U14822 (N_14822,N_14756,N_14783);
nand U14823 (N_14823,N_14686,N_14630);
or U14824 (N_14824,N_14682,N_14605);
nand U14825 (N_14825,N_14760,N_14789);
and U14826 (N_14826,N_14659,N_14732);
xnor U14827 (N_14827,N_14713,N_14708);
xnor U14828 (N_14828,N_14687,N_14740);
nor U14829 (N_14829,N_14727,N_14710);
xnor U14830 (N_14830,N_14791,N_14611);
nor U14831 (N_14831,N_14702,N_14632);
xnor U14832 (N_14832,N_14679,N_14601);
and U14833 (N_14833,N_14750,N_14767);
or U14834 (N_14834,N_14772,N_14633);
nor U14835 (N_14835,N_14635,N_14761);
or U14836 (N_14836,N_14624,N_14643);
nand U14837 (N_14837,N_14618,N_14762);
xor U14838 (N_14838,N_14670,N_14718);
xor U14839 (N_14839,N_14608,N_14777);
nor U14840 (N_14840,N_14614,N_14768);
and U14841 (N_14841,N_14706,N_14607);
xor U14842 (N_14842,N_14674,N_14646);
xor U14843 (N_14843,N_14726,N_14771);
nor U14844 (N_14844,N_14745,N_14738);
and U14845 (N_14845,N_14684,N_14683);
nor U14846 (N_14846,N_14629,N_14623);
and U14847 (N_14847,N_14673,N_14720);
nand U14848 (N_14848,N_14779,N_14715);
and U14849 (N_14849,N_14661,N_14700);
xnor U14850 (N_14850,N_14620,N_14628);
xnor U14851 (N_14851,N_14647,N_14796);
or U14852 (N_14852,N_14739,N_14728);
xor U14853 (N_14853,N_14780,N_14704);
nand U14854 (N_14854,N_14616,N_14652);
nor U14855 (N_14855,N_14758,N_14681);
xnor U14856 (N_14856,N_14658,N_14609);
nand U14857 (N_14857,N_14730,N_14699);
or U14858 (N_14858,N_14716,N_14656);
or U14859 (N_14859,N_14703,N_14698);
nor U14860 (N_14860,N_14733,N_14695);
and U14861 (N_14861,N_14766,N_14786);
and U14862 (N_14862,N_14731,N_14741);
or U14863 (N_14863,N_14711,N_14657);
or U14864 (N_14864,N_14784,N_14603);
nand U14865 (N_14865,N_14645,N_14781);
and U14866 (N_14866,N_14719,N_14615);
xor U14867 (N_14867,N_14763,N_14755);
and U14868 (N_14868,N_14637,N_14600);
nor U14869 (N_14869,N_14691,N_14649);
xnor U14870 (N_14870,N_14676,N_14610);
xnor U14871 (N_14871,N_14666,N_14622);
xnor U14872 (N_14872,N_14742,N_14631);
nand U14873 (N_14873,N_14604,N_14672);
nand U14874 (N_14874,N_14764,N_14668);
nand U14875 (N_14875,N_14722,N_14654);
xor U14876 (N_14876,N_14619,N_14653);
or U14877 (N_14877,N_14612,N_14697);
nand U14878 (N_14878,N_14678,N_14693);
nor U14879 (N_14879,N_14650,N_14759);
nor U14880 (N_14880,N_14765,N_14663);
nor U14881 (N_14881,N_14671,N_14644);
nand U14882 (N_14882,N_14776,N_14798);
nand U14883 (N_14883,N_14675,N_14677);
nor U14884 (N_14884,N_14794,N_14701);
nand U14885 (N_14885,N_14757,N_14752);
nand U14886 (N_14886,N_14753,N_14634);
or U14887 (N_14887,N_14696,N_14680);
xnor U14888 (N_14888,N_14694,N_14775);
nor U14889 (N_14889,N_14797,N_14660);
nor U14890 (N_14890,N_14689,N_14602);
and U14891 (N_14891,N_14621,N_14636);
xor U14892 (N_14892,N_14725,N_14707);
or U14893 (N_14893,N_14793,N_14799);
or U14894 (N_14894,N_14734,N_14639);
and U14895 (N_14895,N_14692,N_14774);
nor U14896 (N_14896,N_14792,N_14788);
nand U14897 (N_14897,N_14617,N_14625);
nand U14898 (N_14898,N_14667,N_14746);
nor U14899 (N_14899,N_14688,N_14709);
and U14900 (N_14900,N_14632,N_14668);
xor U14901 (N_14901,N_14608,N_14779);
nor U14902 (N_14902,N_14666,N_14781);
and U14903 (N_14903,N_14714,N_14725);
and U14904 (N_14904,N_14787,N_14751);
and U14905 (N_14905,N_14785,N_14649);
nor U14906 (N_14906,N_14704,N_14748);
and U14907 (N_14907,N_14784,N_14753);
nand U14908 (N_14908,N_14771,N_14695);
nand U14909 (N_14909,N_14663,N_14751);
or U14910 (N_14910,N_14793,N_14608);
nor U14911 (N_14911,N_14719,N_14756);
xnor U14912 (N_14912,N_14660,N_14774);
and U14913 (N_14913,N_14616,N_14608);
nand U14914 (N_14914,N_14782,N_14711);
or U14915 (N_14915,N_14771,N_14640);
nand U14916 (N_14916,N_14736,N_14631);
nand U14917 (N_14917,N_14675,N_14722);
xor U14918 (N_14918,N_14799,N_14704);
and U14919 (N_14919,N_14668,N_14657);
xnor U14920 (N_14920,N_14670,N_14707);
and U14921 (N_14921,N_14785,N_14742);
and U14922 (N_14922,N_14623,N_14613);
or U14923 (N_14923,N_14614,N_14758);
or U14924 (N_14924,N_14705,N_14634);
xnor U14925 (N_14925,N_14716,N_14605);
nand U14926 (N_14926,N_14618,N_14629);
xor U14927 (N_14927,N_14797,N_14622);
and U14928 (N_14928,N_14670,N_14783);
and U14929 (N_14929,N_14757,N_14607);
or U14930 (N_14930,N_14662,N_14693);
and U14931 (N_14931,N_14710,N_14775);
and U14932 (N_14932,N_14700,N_14733);
nand U14933 (N_14933,N_14729,N_14694);
nand U14934 (N_14934,N_14670,N_14630);
nand U14935 (N_14935,N_14752,N_14754);
nand U14936 (N_14936,N_14623,N_14724);
nor U14937 (N_14937,N_14656,N_14643);
nor U14938 (N_14938,N_14749,N_14787);
nor U14939 (N_14939,N_14690,N_14717);
or U14940 (N_14940,N_14702,N_14641);
nor U14941 (N_14941,N_14782,N_14654);
and U14942 (N_14942,N_14629,N_14677);
nor U14943 (N_14943,N_14721,N_14772);
nand U14944 (N_14944,N_14784,N_14797);
nand U14945 (N_14945,N_14664,N_14732);
xnor U14946 (N_14946,N_14666,N_14629);
or U14947 (N_14947,N_14719,N_14792);
nand U14948 (N_14948,N_14695,N_14601);
xor U14949 (N_14949,N_14707,N_14700);
and U14950 (N_14950,N_14722,N_14681);
nand U14951 (N_14951,N_14653,N_14746);
nand U14952 (N_14952,N_14646,N_14724);
or U14953 (N_14953,N_14634,N_14671);
or U14954 (N_14954,N_14657,N_14771);
or U14955 (N_14955,N_14790,N_14747);
nor U14956 (N_14956,N_14764,N_14770);
nand U14957 (N_14957,N_14781,N_14692);
nor U14958 (N_14958,N_14622,N_14741);
or U14959 (N_14959,N_14783,N_14782);
or U14960 (N_14960,N_14696,N_14760);
nand U14961 (N_14961,N_14601,N_14775);
or U14962 (N_14962,N_14765,N_14687);
or U14963 (N_14963,N_14764,N_14632);
and U14964 (N_14964,N_14794,N_14746);
or U14965 (N_14965,N_14732,N_14654);
or U14966 (N_14966,N_14758,N_14637);
or U14967 (N_14967,N_14680,N_14612);
or U14968 (N_14968,N_14657,N_14715);
nor U14969 (N_14969,N_14770,N_14760);
or U14970 (N_14970,N_14756,N_14793);
xnor U14971 (N_14971,N_14704,N_14626);
nand U14972 (N_14972,N_14633,N_14653);
and U14973 (N_14973,N_14709,N_14713);
or U14974 (N_14974,N_14654,N_14610);
nand U14975 (N_14975,N_14638,N_14762);
and U14976 (N_14976,N_14604,N_14632);
nand U14977 (N_14977,N_14661,N_14744);
nand U14978 (N_14978,N_14765,N_14680);
nand U14979 (N_14979,N_14712,N_14664);
xor U14980 (N_14980,N_14748,N_14682);
and U14981 (N_14981,N_14738,N_14686);
and U14982 (N_14982,N_14770,N_14762);
or U14983 (N_14983,N_14647,N_14710);
nor U14984 (N_14984,N_14769,N_14695);
nand U14985 (N_14985,N_14682,N_14793);
and U14986 (N_14986,N_14605,N_14612);
and U14987 (N_14987,N_14649,N_14725);
nor U14988 (N_14988,N_14713,N_14703);
or U14989 (N_14989,N_14745,N_14783);
xnor U14990 (N_14990,N_14683,N_14776);
nor U14991 (N_14991,N_14721,N_14765);
nor U14992 (N_14992,N_14697,N_14747);
and U14993 (N_14993,N_14661,N_14710);
or U14994 (N_14994,N_14739,N_14637);
or U14995 (N_14995,N_14612,N_14677);
nor U14996 (N_14996,N_14769,N_14626);
or U14997 (N_14997,N_14698,N_14612);
nor U14998 (N_14998,N_14654,N_14688);
xor U14999 (N_14999,N_14737,N_14607);
nand U15000 (N_15000,N_14928,N_14860);
nor U15001 (N_15001,N_14936,N_14995);
or U15002 (N_15002,N_14805,N_14957);
or U15003 (N_15003,N_14898,N_14837);
nor U15004 (N_15004,N_14842,N_14962);
nor U15005 (N_15005,N_14945,N_14810);
or U15006 (N_15006,N_14985,N_14987);
xor U15007 (N_15007,N_14951,N_14980);
xnor U15008 (N_15008,N_14887,N_14940);
or U15009 (N_15009,N_14979,N_14981);
and U15010 (N_15010,N_14930,N_14884);
or U15011 (N_15011,N_14872,N_14809);
nand U15012 (N_15012,N_14913,N_14974);
nand U15013 (N_15013,N_14840,N_14891);
xor U15014 (N_15014,N_14841,N_14829);
nand U15015 (N_15015,N_14915,N_14944);
xor U15016 (N_15016,N_14852,N_14911);
and U15017 (N_15017,N_14893,N_14935);
and U15018 (N_15018,N_14836,N_14997);
nand U15019 (N_15019,N_14952,N_14938);
and U15020 (N_15020,N_14978,N_14819);
nor U15021 (N_15021,N_14948,N_14916);
and U15022 (N_15022,N_14831,N_14811);
xnor U15023 (N_15023,N_14814,N_14932);
and U15024 (N_15024,N_14823,N_14953);
nand U15025 (N_15025,N_14975,N_14888);
and U15026 (N_15026,N_14881,N_14950);
xnor U15027 (N_15027,N_14863,N_14870);
nand U15028 (N_15028,N_14942,N_14896);
xnor U15029 (N_15029,N_14868,N_14966);
nand U15030 (N_15030,N_14990,N_14969);
xnor U15031 (N_15031,N_14924,N_14808);
or U15032 (N_15032,N_14968,N_14854);
xor U15033 (N_15033,N_14834,N_14965);
nand U15034 (N_15034,N_14897,N_14835);
and U15035 (N_15035,N_14925,N_14851);
nor U15036 (N_15036,N_14933,N_14844);
nand U15037 (N_15037,N_14977,N_14964);
and U15038 (N_15038,N_14867,N_14906);
nand U15039 (N_15039,N_14830,N_14857);
nand U15040 (N_15040,N_14845,N_14826);
nand U15041 (N_15041,N_14972,N_14878);
nand U15042 (N_15042,N_14873,N_14838);
nor U15043 (N_15043,N_14992,N_14832);
nand U15044 (N_15044,N_14880,N_14994);
and U15045 (N_15045,N_14989,N_14879);
or U15046 (N_15046,N_14939,N_14864);
nand U15047 (N_15047,N_14943,N_14803);
xor U15048 (N_15048,N_14902,N_14920);
or U15049 (N_15049,N_14883,N_14865);
nand U15050 (N_15050,N_14806,N_14914);
and U15051 (N_15051,N_14846,N_14859);
xnor U15052 (N_15052,N_14890,N_14947);
or U15053 (N_15053,N_14991,N_14801);
xor U15054 (N_15054,N_14812,N_14949);
nor U15055 (N_15055,N_14905,N_14946);
or U15056 (N_15056,N_14959,N_14847);
nand U15057 (N_15057,N_14804,N_14999);
and U15058 (N_15058,N_14998,N_14869);
nor U15059 (N_15059,N_14875,N_14967);
nor U15060 (N_15060,N_14912,N_14954);
or U15061 (N_15061,N_14922,N_14923);
and U15062 (N_15062,N_14816,N_14856);
nand U15063 (N_15063,N_14926,N_14843);
nand U15064 (N_15064,N_14988,N_14800);
or U15065 (N_15065,N_14861,N_14821);
or U15066 (N_15066,N_14970,N_14825);
or U15067 (N_15067,N_14982,N_14827);
xnor U15068 (N_15068,N_14886,N_14918);
nor U15069 (N_15069,N_14910,N_14958);
xor U15070 (N_15070,N_14931,N_14822);
and U15071 (N_15071,N_14895,N_14839);
or U15072 (N_15072,N_14955,N_14815);
xnor U15073 (N_15073,N_14862,N_14904);
nand U15074 (N_15074,N_14901,N_14900);
xor U15075 (N_15075,N_14802,N_14871);
xor U15076 (N_15076,N_14971,N_14828);
xor U15077 (N_15077,N_14853,N_14889);
nor U15078 (N_15078,N_14921,N_14961);
nor U15079 (N_15079,N_14986,N_14820);
nand U15080 (N_15080,N_14892,N_14973);
and U15081 (N_15081,N_14807,N_14907);
nor U15082 (N_15082,N_14996,N_14929);
nor U15083 (N_15083,N_14937,N_14833);
or U15084 (N_15084,N_14882,N_14984);
nor U15085 (N_15085,N_14850,N_14855);
nand U15086 (N_15086,N_14848,N_14899);
nor U15087 (N_15087,N_14963,N_14919);
or U15088 (N_15088,N_14858,N_14877);
and U15089 (N_15089,N_14817,N_14909);
xnor U15090 (N_15090,N_14976,N_14941);
and U15091 (N_15091,N_14876,N_14866);
or U15092 (N_15092,N_14894,N_14956);
xnor U15093 (N_15093,N_14874,N_14934);
or U15094 (N_15094,N_14818,N_14908);
or U15095 (N_15095,N_14849,N_14903);
and U15096 (N_15096,N_14917,N_14993);
or U15097 (N_15097,N_14813,N_14960);
and U15098 (N_15098,N_14885,N_14927);
nand U15099 (N_15099,N_14824,N_14983);
or U15100 (N_15100,N_14990,N_14911);
and U15101 (N_15101,N_14888,N_14812);
or U15102 (N_15102,N_14950,N_14949);
xnor U15103 (N_15103,N_14930,N_14888);
and U15104 (N_15104,N_14814,N_14915);
nor U15105 (N_15105,N_14982,N_14952);
and U15106 (N_15106,N_14866,N_14845);
nand U15107 (N_15107,N_14975,N_14863);
or U15108 (N_15108,N_14983,N_14855);
nor U15109 (N_15109,N_14898,N_14900);
and U15110 (N_15110,N_14947,N_14817);
nand U15111 (N_15111,N_14866,N_14981);
xor U15112 (N_15112,N_14974,N_14971);
xnor U15113 (N_15113,N_14904,N_14978);
xor U15114 (N_15114,N_14820,N_14942);
nor U15115 (N_15115,N_14975,N_14898);
nand U15116 (N_15116,N_14817,N_14837);
xnor U15117 (N_15117,N_14962,N_14824);
nor U15118 (N_15118,N_14896,N_14876);
or U15119 (N_15119,N_14988,N_14954);
and U15120 (N_15120,N_14995,N_14982);
xor U15121 (N_15121,N_14937,N_14994);
and U15122 (N_15122,N_14834,N_14977);
xnor U15123 (N_15123,N_14931,N_14814);
nand U15124 (N_15124,N_14965,N_14995);
and U15125 (N_15125,N_14978,N_14881);
and U15126 (N_15126,N_14902,N_14897);
nor U15127 (N_15127,N_14870,N_14953);
and U15128 (N_15128,N_14809,N_14940);
and U15129 (N_15129,N_14853,N_14814);
nor U15130 (N_15130,N_14807,N_14881);
nand U15131 (N_15131,N_14845,N_14855);
xnor U15132 (N_15132,N_14952,N_14805);
and U15133 (N_15133,N_14972,N_14851);
xor U15134 (N_15134,N_14827,N_14916);
xnor U15135 (N_15135,N_14807,N_14827);
nor U15136 (N_15136,N_14955,N_14862);
or U15137 (N_15137,N_14970,N_14992);
nand U15138 (N_15138,N_14869,N_14941);
and U15139 (N_15139,N_14907,N_14967);
nor U15140 (N_15140,N_14909,N_14927);
nand U15141 (N_15141,N_14881,N_14932);
nor U15142 (N_15142,N_14945,N_14826);
nor U15143 (N_15143,N_14988,N_14942);
nor U15144 (N_15144,N_14903,N_14951);
and U15145 (N_15145,N_14903,N_14873);
and U15146 (N_15146,N_14929,N_14849);
nor U15147 (N_15147,N_14949,N_14928);
nor U15148 (N_15148,N_14911,N_14910);
and U15149 (N_15149,N_14815,N_14997);
nor U15150 (N_15150,N_14937,N_14949);
and U15151 (N_15151,N_14818,N_14938);
xnor U15152 (N_15152,N_14812,N_14802);
nor U15153 (N_15153,N_14958,N_14966);
and U15154 (N_15154,N_14968,N_14988);
nand U15155 (N_15155,N_14973,N_14817);
and U15156 (N_15156,N_14867,N_14944);
xnor U15157 (N_15157,N_14962,N_14974);
xor U15158 (N_15158,N_14807,N_14893);
xnor U15159 (N_15159,N_14830,N_14896);
nor U15160 (N_15160,N_14856,N_14963);
nor U15161 (N_15161,N_14959,N_14951);
and U15162 (N_15162,N_14933,N_14918);
xor U15163 (N_15163,N_14872,N_14930);
xnor U15164 (N_15164,N_14883,N_14902);
xnor U15165 (N_15165,N_14809,N_14973);
or U15166 (N_15166,N_14836,N_14923);
xnor U15167 (N_15167,N_14984,N_14946);
xor U15168 (N_15168,N_14992,N_14922);
nor U15169 (N_15169,N_14904,N_14842);
xor U15170 (N_15170,N_14879,N_14819);
xnor U15171 (N_15171,N_14933,N_14956);
nand U15172 (N_15172,N_14922,N_14905);
xor U15173 (N_15173,N_14824,N_14815);
and U15174 (N_15174,N_14868,N_14934);
and U15175 (N_15175,N_14947,N_14859);
nand U15176 (N_15176,N_14967,N_14896);
or U15177 (N_15177,N_14927,N_14853);
or U15178 (N_15178,N_14953,N_14974);
nor U15179 (N_15179,N_14956,N_14839);
xnor U15180 (N_15180,N_14966,N_14827);
nor U15181 (N_15181,N_14878,N_14970);
and U15182 (N_15182,N_14898,N_14891);
nand U15183 (N_15183,N_14960,N_14993);
nor U15184 (N_15184,N_14974,N_14878);
nand U15185 (N_15185,N_14804,N_14822);
and U15186 (N_15186,N_14878,N_14865);
nand U15187 (N_15187,N_14875,N_14835);
or U15188 (N_15188,N_14835,N_14815);
nor U15189 (N_15189,N_14859,N_14825);
nor U15190 (N_15190,N_14820,N_14953);
nor U15191 (N_15191,N_14800,N_14872);
nor U15192 (N_15192,N_14873,N_14946);
and U15193 (N_15193,N_14824,N_14819);
xor U15194 (N_15194,N_14900,N_14814);
nand U15195 (N_15195,N_14983,N_14827);
nor U15196 (N_15196,N_14853,N_14949);
or U15197 (N_15197,N_14971,N_14949);
xor U15198 (N_15198,N_14894,N_14957);
nor U15199 (N_15199,N_14999,N_14844);
nor U15200 (N_15200,N_15036,N_15122);
xnor U15201 (N_15201,N_15170,N_15181);
nor U15202 (N_15202,N_15195,N_15004);
xnor U15203 (N_15203,N_15185,N_15065);
nand U15204 (N_15204,N_15120,N_15045);
xor U15205 (N_15205,N_15127,N_15021);
nor U15206 (N_15206,N_15081,N_15174);
or U15207 (N_15207,N_15161,N_15037);
nor U15208 (N_15208,N_15156,N_15098);
nor U15209 (N_15209,N_15190,N_15018);
nor U15210 (N_15210,N_15051,N_15013);
nor U15211 (N_15211,N_15192,N_15175);
nor U15212 (N_15212,N_15109,N_15147);
nor U15213 (N_15213,N_15140,N_15153);
or U15214 (N_15214,N_15135,N_15113);
xnor U15215 (N_15215,N_15087,N_15064);
or U15216 (N_15216,N_15006,N_15168);
or U15217 (N_15217,N_15080,N_15139);
and U15218 (N_15218,N_15030,N_15083);
nor U15219 (N_15219,N_15182,N_15000);
and U15220 (N_15220,N_15119,N_15075);
xor U15221 (N_15221,N_15049,N_15062);
xnor U15222 (N_15222,N_15059,N_15040);
or U15223 (N_15223,N_15033,N_15148);
xor U15224 (N_15224,N_15189,N_15115);
xnor U15225 (N_15225,N_15060,N_15101);
nand U15226 (N_15226,N_15166,N_15043);
or U15227 (N_15227,N_15145,N_15138);
and U15228 (N_15228,N_15025,N_15047);
xor U15229 (N_15229,N_15003,N_15094);
or U15230 (N_15230,N_15146,N_15011);
or U15231 (N_15231,N_15034,N_15014);
xnor U15232 (N_15232,N_15050,N_15088);
xor U15233 (N_15233,N_15130,N_15017);
or U15234 (N_15234,N_15117,N_15184);
xnor U15235 (N_15235,N_15169,N_15155);
nand U15236 (N_15236,N_15152,N_15046);
nor U15237 (N_15237,N_15171,N_15091);
and U15238 (N_15238,N_15134,N_15068);
or U15239 (N_15239,N_15188,N_15137);
and U15240 (N_15240,N_15044,N_15024);
and U15241 (N_15241,N_15150,N_15095);
nand U15242 (N_15242,N_15199,N_15183);
and U15243 (N_15243,N_15114,N_15077);
or U15244 (N_15244,N_15015,N_15103);
nor U15245 (N_15245,N_15142,N_15067);
xnor U15246 (N_15246,N_15154,N_15052);
and U15247 (N_15247,N_15159,N_15141);
or U15248 (N_15248,N_15026,N_15076);
nor U15249 (N_15249,N_15010,N_15071);
nor U15250 (N_15250,N_15023,N_15032);
xor U15251 (N_15251,N_15100,N_15099);
nor U15252 (N_15252,N_15187,N_15131);
xnor U15253 (N_15253,N_15019,N_15151);
or U15254 (N_15254,N_15186,N_15085);
nand U15255 (N_15255,N_15078,N_15001);
or U15256 (N_15256,N_15097,N_15086);
and U15257 (N_15257,N_15163,N_15180);
nand U15258 (N_15258,N_15123,N_15106);
nor U15259 (N_15259,N_15111,N_15008);
and U15260 (N_15260,N_15162,N_15167);
nor U15261 (N_15261,N_15110,N_15193);
xor U15262 (N_15262,N_15038,N_15028);
nand U15263 (N_15263,N_15079,N_15031);
and U15264 (N_15264,N_15063,N_15020);
or U15265 (N_15265,N_15012,N_15125);
and U15266 (N_15266,N_15118,N_15089);
nor U15267 (N_15267,N_15176,N_15108);
or U15268 (N_15268,N_15056,N_15173);
nor U15269 (N_15269,N_15121,N_15194);
and U15270 (N_15270,N_15196,N_15053);
nand U15271 (N_15271,N_15061,N_15058);
nand U15272 (N_15272,N_15082,N_15116);
or U15273 (N_15273,N_15074,N_15164);
nor U15274 (N_15274,N_15112,N_15042);
nor U15275 (N_15275,N_15102,N_15096);
or U15276 (N_15276,N_15129,N_15090);
xor U15277 (N_15277,N_15179,N_15092);
nand U15278 (N_15278,N_15143,N_15126);
or U15279 (N_15279,N_15128,N_15066);
nor U15280 (N_15280,N_15165,N_15104);
nand U15281 (N_15281,N_15048,N_15070);
or U15282 (N_15282,N_15191,N_15197);
or U15283 (N_15283,N_15039,N_15007);
nand U15284 (N_15284,N_15035,N_15132);
nor U15285 (N_15285,N_15022,N_15009);
nor U15286 (N_15286,N_15124,N_15172);
or U15287 (N_15287,N_15069,N_15054);
or U15288 (N_15288,N_15041,N_15027);
or U15289 (N_15289,N_15133,N_15149);
and U15290 (N_15290,N_15005,N_15055);
or U15291 (N_15291,N_15016,N_15198);
xor U15292 (N_15292,N_15157,N_15002);
xnor U15293 (N_15293,N_15073,N_15057);
nand U15294 (N_15294,N_15093,N_15160);
nand U15295 (N_15295,N_15144,N_15158);
and U15296 (N_15296,N_15107,N_15084);
and U15297 (N_15297,N_15072,N_15177);
or U15298 (N_15298,N_15105,N_15029);
xor U15299 (N_15299,N_15178,N_15136);
nand U15300 (N_15300,N_15068,N_15196);
xnor U15301 (N_15301,N_15110,N_15047);
and U15302 (N_15302,N_15017,N_15081);
and U15303 (N_15303,N_15030,N_15198);
nor U15304 (N_15304,N_15053,N_15118);
or U15305 (N_15305,N_15100,N_15090);
nand U15306 (N_15306,N_15019,N_15175);
nor U15307 (N_15307,N_15055,N_15183);
nor U15308 (N_15308,N_15187,N_15038);
and U15309 (N_15309,N_15151,N_15140);
and U15310 (N_15310,N_15148,N_15069);
nand U15311 (N_15311,N_15187,N_15119);
nor U15312 (N_15312,N_15052,N_15044);
xor U15313 (N_15313,N_15094,N_15061);
xor U15314 (N_15314,N_15175,N_15021);
nand U15315 (N_15315,N_15084,N_15006);
or U15316 (N_15316,N_15143,N_15048);
nor U15317 (N_15317,N_15131,N_15080);
nor U15318 (N_15318,N_15145,N_15062);
xnor U15319 (N_15319,N_15058,N_15132);
xor U15320 (N_15320,N_15036,N_15194);
nand U15321 (N_15321,N_15035,N_15164);
or U15322 (N_15322,N_15067,N_15088);
and U15323 (N_15323,N_15198,N_15058);
and U15324 (N_15324,N_15084,N_15131);
xor U15325 (N_15325,N_15062,N_15039);
xor U15326 (N_15326,N_15180,N_15165);
nor U15327 (N_15327,N_15058,N_15123);
nand U15328 (N_15328,N_15076,N_15087);
nor U15329 (N_15329,N_15054,N_15007);
and U15330 (N_15330,N_15011,N_15013);
or U15331 (N_15331,N_15107,N_15177);
nor U15332 (N_15332,N_15055,N_15010);
xor U15333 (N_15333,N_15168,N_15175);
xor U15334 (N_15334,N_15173,N_15002);
nor U15335 (N_15335,N_15020,N_15158);
or U15336 (N_15336,N_15152,N_15088);
and U15337 (N_15337,N_15133,N_15040);
or U15338 (N_15338,N_15167,N_15188);
xnor U15339 (N_15339,N_15111,N_15102);
nand U15340 (N_15340,N_15176,N_15052);
and U15341 (N_15341,N_15188,N_15104);
or U15342 (N_15342,N_15196,N_15058);
nand U15343 (N_15343,N_15101,N_15002);
xnor U15344 (N_15344,N_15027,N_15147);
nor U15345 (N_15345,N_15143,N_15115);
xor U15346 (N_15346,N_15074,N_15108);
nand U15347 (N_15347,N_15134,N_15000);
nand U15348 (N_15348,N_15125,N_15151);
xor U15349 (N_15349,N_15162,N_15070);
nand U15350 (N_15350,N_15155,N_15069);
xor U15351 (N_15351,N_15076,N_15027);
nand U15352 (N_15352,N_15099,N_15110);
or U15353 (N_15353,N_15150,N_15080);
xor U15354 (N_15354,N_15002,N_15145);
nand U15355 (N_15355,N_15183,N_15173);
and U15356 (N_15356,N_15030,N_15173);
and U15357 (N_15357,N_15007,N_15182);
and U15358 (N_15358,N_15081,N_15178);
nand U15359 (N_15359,N_15090,N_15134);
xor U15360 (N_15360,N_15066,N_15176);
xnor U15361 (N_15361,N_15074,N_15174);
or U15362 (N_15362,N_15100,N_15167);
nand U15363 (N_15363,N_15189,N_15084);
or U15364 (N_15364,N_15079,N_15075);
and U15365 (N_15365,N_15049,N_15024);
nor U15366 (N_15366,N_15170,N_15082);
or U15367 (N_15367,N_15178,N_15000);
nand U15368 (N_15368,N_15009,N_15123);
or U15369 (N_15369,N_15020,N_15155);
xor U15370 (N_15370,N_15178,N_15100);
nand U15371 (N_15371,N_15146,N_15098);
or U15372 (N_15372,N_15092,N_15172);
and U15373 (N_15373,N_15026,N_15162);
xor U15374 (N_15374,N_15181,N_15088);
and U15375 (N_15375,N_15064,N_15124);
xor U15376 (N_15376,N_15029,N_15000);
or U15377 (N_15377,N_15037,N_15120);
nor U15378 (N_15378,N_15116,N_15181);
or U15379 (N_15379,N_15182,N_15145);
and U15380 (N_15380,N_15096,N_15120);
nor U15381 (N_15381,N_15074,N_15166);
nand U15382 (N_15382,N_15066,N_15040);
xnor U15383 (N_15383,N_15137,N_15092);
or U15384 (N_15384,N_15174,N_15177);
nor U15385 (N_15385,N_15017,N_15062);
nor U15386 (N_15386,N_15107,N_15118);
xnor U15387 (N_15387,N_15152,N_15155);
xnor U15388 (N_15388,N_15177,N_15101);
nor U15389 (N_15389,N_15038,N_15043);
xor U15390 (N_15390,N_15198,N_15108);
nor U15391 (N_15391,N_15121,N_15016);
and U15392 (N_15392,N_15148,N_15158);
or U15393 (N_15393,N_15085,N_15136);
or U15394 (N_15394,N_15013,N_15017);
xnor U15395 (N_15395,N_15002,N_15043);
nor U15396 (N_15396,N_15136,N_15061);
nand U15397 (N_15397,N_15073,N_15155);
or U15398 (N_15398,N_15168,N_15065);
nand U15399 (N_15399,N_15128,N_15051);
and U15400 (N_15400,N_15382,N_15218);
nand U15401 (N_15401,N_15214,N_15395);
xor U15402 (N_15402,N_15365,N_15247);
nor U15403 (N_15403,N_15370,N_15213);
nor U15404 (N_15404,N_15226,N_15210);
xor U15405 (N_15405,N_15308,N_15332);
and U15406 (N_15406,N_15239,N_15291);
nand U15407 (N_15407,N_15333,N_15259);
or U15408 (N_15408,N_15327,N_15256);
nor U15409 (N_15409,N_15389,N_15258);
and U15410 (N_15410,N_15349,N_15233);
nor U15411 (N_15411,N_15205,N_15310);
nand U15412 (N_15412,N_15377,N_15300);
nand U15413 (N_15413,N_15385,N_15374);
nor U15414 (N_15414,N_15270,N_15284);
and U15415 (N_15415,N_15208,N_15371);
xnor U15416 (N_15416,N_15297,N_15224);
nor U15417 (N_15417,N_15222,N_15219);
and U15418 (N_15418,N_15250,N_15343);
nor U15419 (N_15419,N_15306,N_15257);
and U15420 (N_15420,N_15325,N_15293);
or U15421 (N_15421,N_15207,N_15227);
nand U15422 (N_15422,N_15265,N_15268);
xnor U15423 (N_15423,N_15369,N_15215);
xnor U15424 (N_15424,N_15311,N_15290);
and U15425 (N_15425,N_15328,N_15393);
and U15426 (N_15426,N_15249,N_15229);
nand U15427 (N_15427,N_15361,N_15288);
xnor U15428 (N_15428,N_15301,N_15271);
nor U15429 (N_15429,N_15335,N_15359);
nor U15430 (N_15430,N_15201,N_15292);
or U15431 (N_15431,N_15299,N_15321);
nand U15432 (N_15432,N_15309,N_15355);
nand U15433 (N_15433,N_15275,N_15254);
xor U15434 (N_15434,N_15375,N_15357);
and U15435 (N_15435,N_15347,N_15220);
nor U15436 (N_15436,N_15320,N_15302);
or U15437 (N_15437,N_15336,N_15312);
nor U15438 (N_15438,N_15317,N_15245);
or U15439 (N_15439,N_15203,N_15381);
and U15440 (N_15440,N_15294,N_15286);
xor U15441 (N_15441,N_15234,N_15253);
xor U15442 (N_15442,N_15238,N_15240);
and U15443 (N_15443,N_15366,N_15358);
xor U15444 (N_15444,N_15237,N_15241);
nor U15445 (N_15445,N_15346,N_15352);
or U15446 (N_15446,N_15266,N_15331);
nor U15447 (N_15447,N_15396,N_15243);
and U15448 (N_15448,N_15379,N_15260);
nand U15449 (N_15449,N_15350,N_15264);
xnor U15450 (N_15450,N_15384,N_15282);
nand U15451 (N_15451,N_15206,N_15211);
nor U15452 (N_15452,N_15236,N_15277);
nor U15453 (N_15453,N_15383,N_15334);
xor U15454 (N_15454,N_15399,N_15209);
and U15455 (N_15455,N_15318,N_15315);
nor U15456 (N_15456,N_15373,N_15267);
nand U15457 (N_15457,N_15340,N_15280);
nor U15458 (N_15458,N_15263,N_15202);
or U15459 (N_15459,N_15360,N_15281);
xor U15460 (N_15460,N_15269,N_15363);
xor U15461 (N_15461,N_15394,N_15329);
or U15462 (N_15462,N_15216,N_15390);
nand U15463 (N_15463,N_15348,N_15303);
nor U15464 (N_15464,N_15295,N_15376);
or U15465 (N_15465,N_15304,N_15338);
or U15466 (N_15466,N_15232,N_15353);
or U15467 (N_15467,N_15242,N_15344);
xnor U15468 (N_15468,N_15262,N_15319);
nand U15469 (N_15469,N_15223,N_15200);
nand U15470 (N_15470,N_15378,N_15313);
nor U15471 (N_15471,N_15285,N_15341);
xnor U15472 (N_15472,N_15272,N_15387);
nor U15473 (N_15473,N_15398,N_15204);
and U15474 (N_15474,N_15316,N_15337);
nand U15475 (N_15475,N_15342,N_15289);
nor U15476 (N_15476,N_15252,N_15279);
xnor U15477 (N_15477,N_15305,N_15217);
nor U15478 (N_15478,N_15339,N_15367);
or U15479 (N_15479,N_15261,N_15274);
and U15480 (N_15480,N_15212,N_15397);
nor U15481 (N_15481,N_15296,N_15278);
xor U15482 (N_15482,N_15244,N_15364);
or U15483 (N_15483,N_15283,N_15246);
nor U15484 (N_15484,N_15356,N_15225);
or U15485 (N_15485,N_15248,N_15380);
xor U15486 (N_15486,N_15228,N_15354);
and U15487 (N_15487,N_15323,N_15231);
nand U15488 (N_15488,N_15330,N_15345);
and U15489 (N_15489,N_15298,N_15287);
xor U15490 (N_15490,N_15388,N_15221);
xor U15491 (N_15491,N_15276,N_15372);
nand U15492 (N_15492,N_15314,N_15251);
and U15493 (N_15493,N_15235,N_15273);
xor U15494 (N_15494,N_15351,N_15391);
and U15495 (N_15495,N_15322,N_15326);
and U15496 (N_15496,N_15362,N_15307);
nand U15497 (N_15497,N_15230,N_15392);
nor U15498 (N_15498,N_15324,N_15368);
nor U15499 (N_15499,N_15386,N_15255);
nand U15500 (N_15500,N_15364,N_15207);
nand U15501 (N_15501,N_15350,N_15250);
and U15502 (N_15502,N_15386,N_15238);
xor U15503 (N_15503,N_15323,N_15288);
nand U15504 (N_15504,N_15351,N_15209);
or U15505 (N_15505,N_15335,N_15394);
xnor U15506 (N_15506,N_15224,N_15294);
nand U15507 (N_15507,N_15223,N_15315);
or U15508 (N_15508,N_15223,N_15320);
xnor U15509 (N_15509,N_15230,N_15249);
and U15510 (N_15510,N_15241,N_15272);
nand U15511 (N_15511,N_15380,N_15203);
nand U15512 (N_15512,N_15246,N_15378);
and U15513 (N_15513,N_15365,N_15356);
nand U15514 (N_15514,N_15218,N_15360);
or U15515 (N_15515,N_15235,N_15315);
nand U15516 (N_15516,N_15293,N_15291);
and U15517 (N_15517,N_15352,N_15324);
xor U15518 (N_15518,N_15278,N_15253);
xor U15519 (N_15519,N_15313,N_15329);
xnor U15520 (N_15520,N_15228,N_15318);
nor U15521 (N_15521,N_15249,N_15290);
and U15522 (N_15522,N_15222,N_15354);
or U15523 (N_15523,N_15200,N_15367);
or U15524 (N_15524,N_15389,N_15321);
or U15525 (N_15525,N_15331,N_15312);
or U15526 (N_15526,N_15351,N_15231);
nand U15527 (N_15527,N_15276,N_15317);
and U15528 (N_15528,N_15322,N_15371);
and U15529 (N_15529,N_15328,N_15223);
xnor U15530 (N_15530,N_15391,N_15396);
and U15531 (N_15531,N_15257,N_15399);
xnor U15532 (N_15532,N_15393,N_15292);
xor U15533 (N_15533,N_15370,N_15312);
nor U15534 (N_15534,N_15259,N_15388);
and U15535 (N_15535,N_15383,N_15235);
nor U15536 (N_15536,N_15295,N_15361);
and U15537 (N_15537,N_15204,N_15332);
or U15538 (N_15538,N_15321,N_15329);
nor U15539 (N_15539,N_15233,N_15281);
and U15540 (N_15540,N_15246,N_15306);
xnor U15541 (N_15541,N_15282,N_15209);
and U15542 (N_15542,N_15362,N_15380);
and U15543 (N_15543,N_15226,N_15339);
nand U15544 (N_15544,N_15204,N_15394);
and U15545 (N_15545,N_15363,N_15380);
and U15546 (N_15546,N_15371,N_15280);
nand U15547 (N_15547,N_15242,N_15374);
and U15548 (N_15548,N_15295,N_15348);
or U15549 (N_15549,N_15201,N_15290);
and U15550 (N_15550,N_15312,N_15265);
nor U15551 (N_15551,N_15343,N_15355);
nand U15552 (N_15552,N_15322,N_15231);
or U15553 (N_15553,N_15317,N_15320);
or U15554 (N_15554,N_15273,N_15346);
xnor U15555 (N_15555,N_15381,N_15287);
nor U15556 (N_15556,N_15352,N_15283);
nand U15557 (N_15557,N_15346,N_15319);
xor U15558 (N_15558,N_15332,N_15342);
nor U15559 (N_15559,N_15237,N_15379);
nor U15560 (N_15560,N_15315,N_15203);
nor U15561 (N_15561,N_15298,N_15338);
and U15562 (N_15562,N_15253,N_15345);
and U15563 (N_15563,N_15264,N_15337);
and U15564 (N_15564,N_15285,N_15380);
or U15565 (N_15565,N_15390,N_15316);
nand U15566 (N_15566,N_15239,N_15388);
xor U15567 (N_15567,N_15263,N_15376);
and U15568 (N_15568,N_15346,N_15367);
nor U15569 (N_15569,N_15279,N_15239);
xnor U15570 (N_15570,N_15329,N_15257);
and U15571 (N_15571,N_15275,N_15207);
nor U15572 (N_15572,N_15232,N_15253);
xnor U15573 (N_15573,N_15285,N_15391);
nand U15574 (N_15574,N_15308,N_15274);
or U15575 (N_15575,N_15216,N_15370);
or U15576 (N_15576,N_15368,N_15395);
nor U15577 (N_15577,N_15278,N_15211);
and U15578 (N_15578,N_15325,N_15320);
nand U15579 (N_15579,N_15279,N_15202);
or U15580 (N_15580,N_15216,N_15221);
and U15581 (N_15581,N_15305,N_15392);
nor U15582 (N_15582,N_15377,N_15237);
nand U15583 (N_15583,N_15329,N_15264);
xor U15584 (N_15584,N_15224,N_15292);
nand U15585 (N_15585,N_15319,N_15344);
nand U15586 (N_15586,N_15337,N_15334);
nand U15587 (N_15587,N_15300,N_15283);
or U15588 (N_15588,N_15293,N_15258);
nor U15589 (N_15589,N_15380,N_15209);
and U15590 (N_15590,N_15294,N_15299);
nor U15591 (N_15591,N_15388,N_15286);
and U15592 (N_15592,N_15229,N_15318);
and U15593 (N_15593,N_15316,N_15366);
xnor U15594 (N_15594,N_15232,N_15331);
nor U15595 (N_15595,N_15273,N_15311);
or U15596 (N_15596,N_15251,N_15275);
xor U15597 (N_15597,N_15277,N_15279);
or U15598 (N_15598,N_15235,N_15308);
xor U15599 (N_15599,N_15353,N_15387);
and U15600 (N_15600,N_15566,N_15595);
nand U15601 (N_15601,N_15466,N_15436);
or U15602 (N_15602,N_15464,N_15522);
and U15603 (N_15603,N_15480,N_15468);
nand U15604 (N_15604,N_15452,N_15430);
and U15605 (N_15605,N_15451,N_15579);
nand U15606 (N_15606,N_15502,N_15409);
xnor U15607 (N_15607,N_15527,N_15467);
nand U15608 (N_15608,N_15557,N_15532);
nor U15609 (N_15609,N_15514,N_15441);
xnor U15610 (N_15610,N_15418,N_15541);
xor U15611 (N_15611,N_15587,N_15599);
or U15612 (N_15612,N_15513,N_15564);
or U15613 (N_15613,N_15412,N_15421);
xor U15614 (N_15614,N_15463,N_15448);
nor U15615 (N_15615,N_15563,N_15507);
or U15616 (N_15616,N_15497,N_15420);
nor U15617 (N_15617,N_15492,N_15465);
nand U15618 (N_15618,N_15509,N_15444);
nand U15619 (N_15619,N_15403,N_15489);
nor U15620 (N_15620,N_15469,N_15455);
and U15621 (N_15621,N_15598,N_15560);
or U15622 (N_15622,N_15400,N_15594);
nand U15623 (N_15623,N_15581,N_15439);
xor U15624 (N_15624,N_15591,N_15588);
nor U15625 (N_15625,N_15445,N_15506);
or U15626 (N_15626,N_15434,N_15553);
nor U15627 (N_15627,N_15470,N_15578);
or U15628 (N_15628,N_15475,N_15411);
nand U15629 (N_15629,N_15437,N_15562);
or U15630 (N_15630,N_15414,N_15481);
nand U15631 (N_15631,N_15567,N_15556);
nand U15632 (N_15632,N_15534,N_15461);
nor U15633 (N_15633,N_15558,N_15431);
nor U15634 (N_15634,N_15424,N_15416);
and U15635 (N_15635,N_15586,N_15597);
nand U15636 (N_15636,N_15404,N_15550);
and U15637 (N_15637,N_15576,N_15410);
and U15638 (N_15638,N_15406,N_15443);
nand U15639 (N_15639,N_15524,N_15542);
nand U15640 (N_15640,N_15505,N_15545);
nand U15641 (N_15641,N_15495,N_15584);
xnor U15642 (N_15642,N_15433,N_15554);
nand U15643 (N_15643,N_15575,N_15548);
or U15644 (N_15644,N_15508,N_15582);
or U15645 (N_15645,N_15478,N_15498);
nor U15646 (N_15646,N_15453,N_15511);
xor U15647 (N_15647,N_15539,N_15474);
or U15648 (N_15648,N_15486,N_15457);
or U15649 (N_15649,N_15459,N_15547);
or U15650 (N_15650,N_15408,N_15561);
xnor U15651 (N_15651,N_15460,N_15458);
nor U15652 (N_15652,N_15425,N_15555);
nor U15653 (N_15653,N_15573,N_15426);
and U15654 (N_15654,N_15523,N_15485);
or U15655 (N_15655,N_15520,N_15405);
and U15656 (N_15656,N_15442,N_15535);
nand U15657 (N_15657,N_15501,N_15515);
nor U15658 (N_15658,N_15574,N_15544);
nand U15659 (N_15659,N_15490,N_15543);
and U15660 (N_15660,N_15538,N_15590);
and U15661 (N_15661,N_15552,N_15536);
and U15662 (N_15662,N_15519,N_15585);
xor U15663 (N_15663,N_15589,N_15484);
and U15664 (N_15664,N_15549,N_15477);
nor U15665 (N_15665,N_15537,N_15592);
nand U15666 (N_15666,N_15521,N_15551);
nor U15667 (N_15667,N_15517,N_15510);
xor U15668 (N_15668,N_15568,N_15415);
and U15669 (N_15669,N_15540,N_15572);
nor U15670 (N_15670,N_15454,N_15569);
nor U15671 (N_15671,N_15446,N_15427);
nand U15672 (N_15672,N_15559,N_15518);
or U15673 (N_15673,N_15456,N_15422);
nor U15674 (N_15674,N_15479,N_15440);
and U15675 (N_15675,N_15473,N_15583);
xor U15676 (N_15676,N_15565,N_15462);
nor U15677 (N_15677,N_15493,N_15423);
nor U15678 (N_15678,N_15571,N_15516);
nor U15679 (N_15679,N_15533,N_15530);
or U15680 (N_15680,N_15546,N_15402);
nor U15681 (N_15681,N_15472,N_15526);
and U15682 (N_15682,N_15471,N_15417);
nand U15683 (N_15683,N_15496,N_15435);
xnor U15684 (N_15684,N_15512,N_15500);
nand U15685 (N_15685,N_15593,N_15531);
xnor U15686 (N_15686,N_15504,N_15428);
nor U15687 (N_15687,N_15482,N_15487);
and U15688 (N_15688,N_15570,N_15432);
or U15689 (N_15689,N_15528,N_15449);
xor U15690 (N_15690,N_15413,N_15580);
xnor U15691 (N_15691,N_15503,N_15499);
or U15692 (N_15692,N_15529,N_15483);
nor U15693 (N_15693,N_15577,N_15488);
xnor U15694 (N_15694,N_15407,N_15429);
xor U15695 (N_15695,N_15596,N_15450);
and U15696 (N_15696,N_15401,N_15438);
xor U15697 (N_15697,N_15476,N_15491);
nor U15698 (N_15698,N_15419,N_15494);
nand U15699 (N_15699,N_15525,N_15447);
nand U15700 (N_15700,N_15556,N_15417);
or U15701 (N_15701,N_15419,N_15471);
nor U15702 (N_15702,N_15568,N_15556);
and U15703 (N_15703,N_15461,N_15500);
and U15704 (N_15704,N_15443,N_15541);
nand U15705 (N_15705,N_15468,N_15404);
or U15706 (N_15706,N_15402,N_15529);
or U15707 (N_15707,N_15419,N_15423);
and U15708 (N_15708,N_15544,N_15412);
nand U15709 (N_15709,N_15462,N_15489);
nor U15710 (N_15710,N_15481,N_15522);
or U15711 (N_15711,N_15502,N_15526);
or U15712 (N_15712,N_15591,N_15466);
nand U15713 (N_15713,N_15482,N_15597);
nand U15714 (N_15714,N_15418,N_15589);
and U15715 (N_15715,N_15508,N_15424);
xor U15716 (N_15716,N_15443,N_15536);
nor U15717 (N_15717,N_15486,N_15596);
nand U15718 (N_15718,N_15539,N_15553);
and U15719 (N_15719,N_15446,N_15555);
nand U15720 (N_15720,N_15470,N_15442);
xnor U15721 (N_15721,N_15448,N_15549);
nand U15722 (N_15722,N_15502,N_15588);
nor U15723 (N_15723,N_15489,N_15573);
and U15724 (N_15724,N_15537,N_15586);
xnor U15725 (N_15725,N_15479,N_15441);
nor U15726 (N_15726,N_15517,N_15469);
and U15727 (N_15727,N_15562,N_15547);
nand U15728 (N_15728,N_15454,N_15410);
nand U15729 (N_15729,N_15481,N_15562);
or U15730 (N_15730,N_15579,N_15456);
nor U15731 (N_15731,N_15426,N_15513);
xnor U15732 (N_15732,N_15520,N_15599);
nor U15733 (N_15733,N_15510,N_15434);
nor U15734 (N_15734,N_15492,N_15444);
xor U15735 (N_15735,N_15598,N_15534);
nand U15736 (N_15736,N_15464,N_15485);
and U15737 (N_15737,N_15476,N_15464);
or U15738 (N_15738,N_15552,N_15532);
and U15739 (N_15739,N_15451,N_15599);
or U15740 (N_15740,N_15568,N_15489);
xor U15741 (N_15741,N_15407,N_15561);
nor U15742 (N_15742,N_15548,N_15556);
and U15743 (N_15743,N_15418,N_15594);
and U15744 (N_15744,N_15585,N_15402);
xor U15745 (N_15745,N_15515,N_15514);
xor U15746 (N_15746,N_15480,N_15479);
or U15747 (N_15747,N_15459,N_15555);
xnor U15748 (N_15748,N_15450,N_15505);
nand U15749 (N_15749,N_15532,N_15588);
nand U15750 (N_15750,N_15569,N_15480);
or U15751 (N_15751,N_15414,N_15455);
xor U15752 (N_15752,N_15427,N_15425);
nor U15753 (N_15753,N_15446,N_15537);
nor U15754 (N_15754,N_15475,N_15448);
and U15755 (N_15755,N_15490,N_15418);
nand U15756 (N_15756,N_15536,N_15480);
xnor U15757 (N_15757,N_15460,N_15450);
and U15758 (N_15758,N_15569,N_15464);
or U15759 (N_15759,N_15419,N_15444);
nand U15760 (N_15760,N_15550,N_15493);
nor U15761 (N_15761,N_15512,N_15451);
or U15762 (N_15762,N_15578,N_15496);
or U15763 (N_15763,N_15438,N_15477);
xor U15764 (N_15764,N_15594,N_15499);
nand U15765 (N_15765,N_15502,N_15444);
or U15766 (N_15766,N_15489,N_15493);
xnor U15767 (N_15767,N_15552,N_15534);
xor U15768 (N_15768,N_15466,N_15444);
nand U15769 (N_15769,N_15432,N_15486);
and U15770 (N_15770,N_15593,N_15415);
or U15771 (N_15771,N_15483,N_15521);
and U15772 (N_15772,N_15406,N_15446);
and U15773 (N_15773,N_15460,N_15597);
nor U15774 (N_15774,N_15586,N_15484);
or U15775 (N_15775,N_15458,N_15401);
nand U15776 (N_15776,N_15409,N_15437);
nand U15777 (N_15777,N_15528,N_15469);
nor U15778 (N_15778,N_15547,N_15538);
and U15779 (N_15779,N_15554,N_15574);
xor U15780 (N_15780,N_15522,N_15473);
nand U15781 (N_15781,N_15558,N_15446);
xnor U15782 (N_15782,N_15508,N_15443);
nand U15783 (N_15783,N_15594,N_15565);
xnor U15784 (N_15784,N_15579,N_15470);
nor U15785 (N_15785,N_15433,N_15488);
or U15786 (N_15786,N_15460,N_15492);
nor U15787 (N_15787,N_15543,N_15452);
or U15788 (N_15788,N_15533,N_15440);
xnor U15789 (N_15789,N_15553,N_15444);
xnor U15790 (N_15790,N_15446,N_15461);
xor U15791 (N_15791,N_15590,N_15427);
nor U15792 (N_15792,N_15475,N_15577);
xor U15793 (N_15793,N_15469,N_15438);
nand U15794 (N_15794,N_15413,N_15524);
and U15795 (N_15795,N_15468,N_15401);
nand U15796 (N_15796,N_15491,N_15420);
xor U15797 (N_15797,N_15552,N_15507);
or U15798 (N_15798,N_15569,N_15559);
and U15799 (N_15799,N_15520,N_15449);
xnor U15800 (N_15800,N_15755,N_15621);
nand U15801 (N_15801,N_15679,N_15725);
nand U15802 (N_15802,N_15650,N_15683);
nand U15803 (N_15803,N_15688,N_15671);
and U15804 (N_15804,N_15618,N_15646);
and U15805 (N_15805,N_15750,N_15705);
xor U15806 (N_15806,N_15625,N_15785);
xor U15807 (N_15807,N_15732,N_15788);
nor U15808 (N_15808,N_15699,N_15713);
and U15809 (N_15809,N_15685,N_15702);
xor U15810 (N_15810,N_15665,N_15652);
and U15811 (N_15811,N_15739,N_15793);
nand U15812 (N_15812,N_15669,N_15765);
or U15813 (N_15813,N_15745,N_15603);
nand U15814 (N_15814,N_15609,N_15734);
or U15815 (N_15815,N_15778,N_15626);
xor U15816 (N_15816,N_15619,N_15795);
and U15817 (N_15817,N_15747,N_15620);
and U15818 (N_15818,N_15744,N_15756);
and U15819 (N_15819,N_15730,N_15703);
nor U15820 (N_15820,N_15704,N_15658);
and U15821 (N_15821,N_15753,N_15754);
and U15822 (N_15822,N_15727,N_15799);
nand U15823 (N_15823,N_15656,N_15726);
nor U15824 (N_15824,N_15711,N_15742);
nor U15825 (N_15825,N_15694,N_15772);
nor U15826 (N_15826,N_15654,N_15653);
and U15827 (N_15827,N_15718,N_15636);
xnor U15828 (N_15828,N_15686,N_15708);
or U15829 (N_15829,N_15712,N_15696);
and U15830 (N_15830,N_15600,N_15616);
nand U15831 (N_15831,N_15783,N_15647);
xnor U15832 (N_15832,N_15627,N_15645);
and U15833 (N_15833,N_15638,N_15667);
xnor U15834 (N_15834,N_15786,N_15698);
xor U15835 (N_15835,N_15700,N_15673);
xor U15836 (N_15836,N_15615,N_15623);
nor U15837 (N_15837,N_15635,N_15630);
nand U15838 (N_15838,N_15674,N_15752);
nand U15839 (N_15839,N_15723,N_15748);
or U15840 (N_15840,N_15749,N_15682);
nand U15841 (N_15841,N_15709,N_15779);
and U15842 (N_15842,N_15695,N_15759);
xor U15843 (N_15843,N_15776,N_15605);
nor U15844 (N_15844,N_15681,N_15606);
xor U15845 (N_15845,N_15782,N_15791);
xor U15846 (N_15846,N_15763,N_15648);
xnor U15847 (N_15847,N_15758,N_15641);
and U15848 (N_15848,N_15787,N_15670);
nand U15849 (N_15849,N_15773,N_15660);
nor U15850 (N_15850,N_15719,N_15736);
nand U15851 (N_15851,N_15684,N_15720);
nand U15852 (N_15852,N_15613,N_15659);
nand U15853 (N_15853,N_15722,N_15666);
and U15854 (N_15854,N_15633,N_15716);
xor U15855 (N_15855,N_15678,N_15737);
nor U15856 (N_15856,N_15717,N_15611);
nor U15857 (N_15857,N_15769,N_15746);
or U15858 (N_15858,N_15691,N_15687);
or U15859 (N_15859,N_15639,N_15707);
or U15860 (N_15860,N_15770,N_15697);
xnor U15861 (N_15861,N_15774,N_15760);
nor U15862 (N_15862,N_15612,N_15604);
xnor U15863 (N_15863,N_15608,N_15735);
nor U15864 (N_15864,N_15740,N_15796);
or U15865 (N_15865,N_15643,N_15661);
nand U15866 (N_15866,N_15655,N_15797);
nand U15867 (N_15867,N_15794,N_15689);
or U15868 (N_15868,N_15798,N_15714);
xnor U15869 (N_15869,N_15629,N_15729);
or U15870 (N_15870,N_15614,N_15784);
nand U15871 (N_15871,N_15610,N_15789);
or U15872 (N_15872,N_15657,N_15677);
xor U15873 (N_15873,N_15624,N_15668);
xor U15874 (N_15874,N_15780,N_15662);
and U15875 (N_15875,N_15706,N_15651);
xnor U15876 (N_15876,N_15731,N_15634);
and U15877 (N_15877,N_15733,N_15607);
or U15878 (N_15878,N_15775,N_15728);
nand U15879 (N_15879,N_15767,N_15622);
nand U15880 (N_15880,N_15762,N_15632);
and U15881 (N_15881,N_15766,N_15601);
xor U15882 (N_15882,N_15771,N_15676);
nor U15883 (N_15883,N_15764,N_15768);
or U15884 (N_15884,N_15738,N_15637);
and U15885 (N_15885,N_15617,N_15790);
or U15886 (N_15886,N_15690,N_15631);
nor U15887 (N_15887,N_15692,N_15693);
nand U15888 (N_15888,N_15675,N_15781);
or U15889 (N_15889,N_15672,N_15701);
or U15890 (N_15890,N_15710,N_15777);
xor U15891 (N_15891,N_15721,N_15761);
and U15892 (N_15892,N_15664,N_15792);
nand U15893 (N_15893,N_15724,N_15743);
and U15894 (N_15894,N_15663,N_15602);
or U15895 (N_15895,N_15640,N_15757);
nor U15896 (N_15896,N_15680,N_15644);
and U15897 (N_15897,N_15741,N_15649);
nor U15898 (N_15898,N_15715,N_15642);
xor U15899 (N_15899,N_15751,N_15628);
xor U15900 (N_15900,N_15614,N_15693);
xnor U15901 (N_15901,N_15624,N_15694);
or U15902 (N_15902,N_15691,N_15695);
nand U15903 (N_15903,N_15777,N_15795);
or U15904 (N_15904,N_15676,N_15697);
or U15905 (N_15905,N_15693,N_15687);
and U15906 (N_15906,N_15754,N_15701);
and U15907 (N_15907,N_15674,N_15609);
or U15908 (N_15908,N_15749,N_15602);
nor U15909 (N_15909,N_15684,N_15702);
xor U15910 (N_15910,N_15697,N_15692);
or U15911 (N_15911,N_15703,N_15765);
or U15912 (N_15912,N_15737,N_15734);
xnor U15913 (N_15913,N_15682,N_15641);
nand U15914 (N_15914,N_15649,N_15719);
nor U15915 (N_15915,N_15693,N_15751);
nor U15916 (N_15916,N_15724,N_15638);
and U15917 (N_15917,N_15766,N_15704);
nand U15918 (N_15918,N_15620,N_15654);
and U15919 (N_15919,N_15701,N_15715);
and U15920 (N_15920,N_15771,N_15795);
nand U15921 (N_15921,N_15795,N_15701);
nor U15922 (N_15922,N_15705,N_15636);
and U15923 (N_15923,N_15698,N_15610);
nor U15924 (N_15924,N_15695,N_15688);
nand U15925 (N_15925,N_15663,N_15780);
nor U15926 (N_15926,N_15751,N_15603);
or U15927 (N_15927,N_15799,N_15751);
nand U15928 (N_15928,N_15779,N_15627);
nand U15929 (N_15929,N_15607,N_15799);
or U15930 (N_15930,N_15661,N_15766);
xor U15931 (N_15931,N_15607,N_15749);
nor U15932 (N_15932,N_15644,N_15768);
and U15933 (N_15933,N_15773,N_15704);
or U15934 (N_15934,N_15616,N_15745);
and U15935 (N_15935,N_15672,N_15622);
and U15936 (N_15936,N_15709,N_15743);
or U15937 (N_15937,N_15716,N_15737);
xnor U15938 (N_15938,N_15686,N_15681);
and U15939 (N_15939,N_15696,N_15793);
nand U15940 (N_15940,N_15740,N_15685);
nand U15941 (N_15941,N_15674,N_15681);
xor U15942 (N_15942,N_15770,N_15667);
and U15943 (N_15943,N_15715,N_15712);
nand U15944 (N_15944,N_15607,N_15727);
nor U15945 (N_15945,N_15609,N_15738);
xnor U15946 (N_15946,N_15693,N_15766);
xnor U15947 (N_15947,N_15671,N_15757);
xnor U15948 (N_15948,N_15760,N_15746);
nor U15949 (N_15949,N_15613,N_15603);
nor U15950 (N_15950,N_15659,N_15742);
or U15951 (N_15951,N_15650,N_15777);
and U15952 (N_15952,N_15669,N_15741);
xor U15953 (N_15953,N_15761,N_15772);
and U15954 (N_15954,N_15643,N_15625);
nor U15955 (N_15955,N_15757,N_15754);
nor U15956 (N_15956,N_15627,N_15625);
nor U15957 (N_15957,N_15743,N_15623);
xor U15958 (N_15958,N_15772,N_15643);
nor U15959 (N_15959,N_15654,N_15797);
and U15960 (N_15960,N_15787,N_15713);
xnor U15961 (N_15961,N_15627,N_15686);
or U15962 (N_15962,N_15650,N_15651);
nor U15963 (N_15963,N_15720,N_15649);
nand U15964 (N_15964,N_15792,N_15670);
xor U15965 (N_15965,N_15665,N_15749);
nand U15966 (N_15966,N_15695,N_15773);
or U15967 (N_15967,N_15703,N_15678);
and U15968 (N_15968,N_15763,N_15750);
nor U15969 (N_15969,N_15679,N_15782);
or U15970 (N_15970,N_15688,N_15768);
xnor U15971 (N_15971,N_15687,N_15773);
nand U15972 (N_15972,N_15649,N_15736);
or U15973 (N_15973,N_15703,N_15609);
xor U15974 (N_15974,N_15603,N_15633);
nand U15975 (N_15975,N_15743,N_15637);
or U15976 (N_15976,N_15648,N_15719);
xnor U15977 (N_15977,N_15712,N_15738);
nor U15978 (N_15978,N_15739,N_15697);
xnor U15979 (N_15979,N_15681,N_15740);
or U15980 (N_15980,N_15682,N_15754);
and U15981 (N_15981,N_15753,N_15692);
nor U15982 (N_15982,N_15741,N_15799);
nand U15983 (N_15983,N_15639,N_15676);
xnor U15984 (N_15984,N_15784,N_15600);
and U15985 (N_15985,N_15791,N_15645);
nand U15986 (N_15986,N_15645,N_15772);
or U15987 (N_15987,N_15781,N_15797);
nand U15988 (N_15988,N_15704,N_15670);
xnor U15989 (N_15989,N_15671,N_15792);
nor U15990 (N_15990,N_15634,N_15784);
nor U15991 (N_15991,N_15765,N_15619);
nor U15992 (N_15992,N_15768,N_15663);
nor U15993 (N_15993,N_15742,N_15777);
or U15994 (N_15994,N_15782,N_15659);
xnor U15995 (N_15995,N_15687,N_15793);
nand U15996 (N_15996,N_15604,N_15735);
xnor U15997 (N_15997,N_15711,N_15778);
and U15998 (N_15998,N_15600,N_15749);
or U15999 (N_15999,N_15682,N_15707);
nor U16000 (N_16000,N_15970,N_15967);
xnor U16001 (N_16001,N_15871,N_15832);
or U16002 (N_16002,N_15981,N_15813);
or U16003 (N_16003,N_15994,N_15891);
or U16004 (N_16004,N_15931,N_15973);
nand U16005 (N_16005,N_15854,N_15989);
xnor U16006 (N_16006,N_15917,N_15905);
or U16007 (N_16007,N_15982,N_15828);
or U16008 (N_16008,N_15975,N_15887);
and U16009 (N_16009,N_15878,N_15962);
or U16010 (N_16010,N_15993,N_15952);
and U16011 (N_16011,N_15807,N_15923);
nor U16012 (N_16012,N_15851,N_15977);
xnor U16013 (N_16013,N_15960,N_15873);
nor U16014 (N_16014,N_15961,N_15944);
nand U16015 (N_16015,N_15872,N_15950);
and U16016 (N_16016,N_15838,N_15978);
nand U16017 (N_16017,N_15829,N_15914);
or U16018 (N_16018,N_15818,N_15949);
xnor U16019 (N_16019,N_15830,N_15897);
nand U16020 (N_16020,N_15968,N_15825);
xnor U16021 (N_16021,N_15995,N_15913);
or U16022 (N_16022,N_15869,N_15925);
or U16023 (N_16023,N_15937,N_15881);
and U16024 (N_16024,N_15951,N_15898);
nor U16025 (N_16025,N_15964,N_15958);
xnor U16026 (N_16026,N_15842,N_15804);
nand U16027 (N_16027,N_15976,N_15948);
nor U16028 (N_16028,N_15808,N_15922);
nand U16029 (N_16029,N_15884,N_15864);
nor U16030 (N_16030,N_15929,N_15957);
nor U16031 (N_16031,N_15852,N_15894);
xor U16032 (N_16032,N_15936,N_15947);
or U16033 (N_16033,N_15844,N_15827);
nand U16034 (N_16034,N_15833,N_15940);
xor U16035 (N_16035,N_15927,N_15810);
nor U16036 (N_16036,N_15990,N_15971);
xor U16037 (N_16037,N_15910,N_15900);
and U16038 (N_16038,N_15826,N_15892);
nor U16039 (N_16039,N_15814,N_15903);
and U16040 (N_16040,N_15904,N_15984);
nand U16041 (N_16041,N_15901,N_15885);
nor U16042 (N_16042,N_15959,N_15979);
or U16043 (N_16043,N_15845,N_15856);
or U16044 (N_16044,N_15867,N_15911);
nand U16045 (N_16045,N_15837,N_15916);
nor U16046 (N_16046,N_15966,N_15935);
or U16047 (N_16047,N_15835,N_15843);
xor U16048 (N_16048,N_15877,N_15907);
nor U16049 (N_16049,N_15806,N_15924);
or U16050 (N_16050,N_15805,N_15819);
xor U16051 (N_16051,N_15899,N_15853);
nor U16052 (N_16052,N_15841,N_15938);
nand U16053 (N_16053,N_15939,N_15850);
nand U16054 (N_16054,N_15840,N_15886);
nand U16055 (N_16055,N_15946,N_15824);
nand U16056 (N_16056,N_15987,N_15956);
nor U16057 (N_16057,N_15908,N_15986);
nand U16058 (N_16058,N_15875,N_15889);
or U16059 (N_16059,N_15811,N_15921);
nand U16060 (N_16060,N_15919,N_15926);
nand U16061 (N_16061,N_15953,N_15920);
nand U16062 (N_16062,N_15800,N_15876);
or U16063 (N_16063,N_15870,N_15801);
xor U16064 (N_16064,N_15803,N_15915);
nand U16065 (N_16065,N_15863,N_15836);
and U16066 (N_16066,N_15912,N_15890);
nand U16067 (N_16067,N_15882,N_15932);
nand U16068 (N_16068,N_15963,N_15941);
xnor U16069 (N_16069,N_15879,N_15985);
nand U16070 (N_16070,N_15972,N_15906);
nand U16071 (N_16071,N_15933,N_15997);
and U16072 (N_16072,N_15895,N_15943);
or U16073 (N_16073,N_15822,N_15866);
and U16074 (N_16074,N_15857,N_15848);
nor U16075 (N_16075,N_15809,N_15902);
nand U16076 (N_16076,N_15934,N_15865);
xnor U16077 (N_16077,N_15928,N_15991);
nand U16078 (N_16078,N_15945,N_15909);
or U16079 (N_16079,N_15817,N_15942);
and U16080 (N_16080,N_15918,N_15820);
nor U16081 (N_16081,N_15874,N_15930);
and U16082 (N_16082,N_15896,N_15847);
xnor U16083 (N_16083,N_15996,N_15861);
nand U16084 (N_16084,N_15834,N_15868);
xnor U16085 (N_16085,N_15839,N_15954);
nor U16086 (N_16086,N_15823,N_15880);
nor U16087 (N_16087,N_15816,N_15955);
nand U16088 (N_16088,N_15821,N_15999);
and U16089 (N_16089,N_15980,N_15858);
xnor U16090 (N_16090,N_15893,N_15862);
and U16091 (N_16091,N_15831,N_15965);
or U16092 (N_16092,N_15983,N_15815);
xnor U16093 (N_16093,N_15888,N_15855);
nor U16094 (N_16094,N_15974,N_15860);
nor U16095 (N_16095,N_15992,N_15883);
nor U16096 (N_16096,N_15802,N_15969);
nor U16097 (N_16097,N_15988,N_15998);
nand U16098 (N_16098,N_15859,N_15846);
nor U16099 (N_16099,N_15812,N_15849);
nand U16100 (N_16100,N_15869,N_15804);
nand U16101 (N_16101,N_15998,N_15862);
nor U16102 (N_16102,N_15944,N_15976);
nand U16103 (N_16103,N_15987,N_15992);
nor U16104 (N_16104,N_15908,N_15872);
nor U16105 (N_16105,N_15860,N_15867);
and U16106 (N_16106,N_15985,N_15961);
or U16107 (N_16107,N_15915,N_15892);
nand U16108 (N_16108,N_15880,N_15833);
xnor U16109 (N_16109,N_15814,N_15851);
or U16110 (N_16110,N_15916,N_15988);
nor U16111 (N_16111,N_15877,N_15855);
nand U16112 (N_16112,N_15996,N_15944);
and U16113 (N_16113,N_15936,N_15920);
and U16114 (N_16114,N_15946,N_15844);
and U16115 (N_16115,N_15906,N_15883);
and U16116 (N_16116,N_15978,N_15904);
xor U16117 (N_16117,N_15898,N_15858);
nor U16118 (N_16118,N_15954,N_15967);
xnor U16119 (N_16119,N_15945,N_15938);
and U16120 (N_16120,N_15976,N_15809);
nor U16121 (N_16121,N_15970,N_15862);
and U16122 (N_16122,N_15942,N_15961);
and U16123 (N_16123,N_15947,N_15887);
or U16124 (N_16124,N_15813,N_15937);
nand U16125 (N_16125,N_15883,N_15864);
and U16126 (N_16126,N_15871,N_15980);
nand U16127 (N_16127,N_15995,N_15958);
and U16128 (N_16128,N_15867,N_15842);
xnor U16129 (N_16129,N_15899,N_15975);
nor U16130 (N_16130,N_15818,N_15866);
and U16131 (N_16131,N_15843,N_15868);
and U16132 (N_16132,N_15866,N_15960);
xor U16133 (N_16133,N_15850,N_15888);
or U16134 (N_16134,N_15880,N_15964);
nor U16135 (N_16135,N_15819,N_15835);
or U16136 (N_16136,N_15984,N_15858);
or U16137 (N_16137,N_15848,N_15849);
nand U16138 (N_16138,N_15878,N_15936);
nand U16139 (N_16139,N_15901,N_15881);
and U16140 (N_16140,N_15867,N_15932);
nor U16141 (N_16141,N_15857,N_15900);
xor U16142 (N_16142,N_15831,N_15850);
and U16143 (N_16143,N_15805,N_15851);
xor U16144 (N_16144,N_15983,N_15892);
or U16145 (N_16145,N_15938,N_15803);
nor U16146 (N_16146,N_15836,N_15987);
or U16147 (N_16147,N_15972,N_15800);
nor U16148 (N_16148,N_15818,N_15941);
xor U16149 (N_16149,N_15929,N_15869);
nand U16150 (N_16150,N_15839,N_15868);
or U16151 (N_16151,N_15817,N_15883);
nor U16152 (N_16152,N_15917,N_15934);
xor U16153 (N_16153,N_15935,N_15934);
and U16154 (N_16154,N_15957,N_15945);
nand U16155 (N_16155,N_15970,N_15997);
or U16156 (N_16156,N_15940,N_15831);
xor U16157 (N_16157,N_15990,N_15833);
or U16158 (N_16158,N_15812,N_15965);
nand U16159 (N_16159,N_15858,N_15989);
nor U16160 (N_16160,N_15877,N_15808);
nand U16161 (N_16161,N_15814,N_15825);
and U16162 (N_16162,N_15893,N_15987);
nand U16163 (N_16163,N_15917,N_15948);
xor U16164 (N_16164,N_15904,N_15824);
and U16165 (N_16165,N_15992,N_15900);
xor U16166 (N_16166,N_15834,N_15805);
nor U16167 (N_16167,N_15919,N_15873);
or U16168 (N_16168,N_15873,N_15988);
or U16169 (N_16169,N_15814,N_15844);
or U16170 (N_16170,N_15975,N_15869);
or U16171 (N_16171,N_15855,N_15924);
or U16172 (N_16172,N_15903,N_15950);
nor U16173 (N_16173,N_15985,N_15941);
nor U16174 (N_16174,N_15989,N_15935);
nor U16175 (N_16175,N_15929,N_15966);
or U16176 (N_16176,N_15843,N_15881);
or U16177 (N_16177,N_15808,N_15890);
or U16178 (N_16178,N_15949,N_15910);
nor U16179 (N_16179,N_15851,N_15862);
and U16180 (N_16180,N_15842,N_15955);
or U16181 (N_16181,N_15916,N_15801);
nand U16182 (N_16182,N_15855,N_15911);
and U16183 (N_16183,N_15946,N_15982);
and U16184 (N_16184,N_15820,N_15888);
nor U16185 (N_16185,N_15883,N_15988);
nor U16186 (N_16186,N_15808,N_15829);
nand U16187 (N_16187,N_15851,N_15914);
nand U16188 (N_16188,N_15848,N_15889);
and U16189 (N_16189,N_15868,N_15840);
nand U16190 (N_16190,N_15943,N_15963);
and U16191 (N_16191,N_15912,N_15921);
and U16192 (N_16192,N_15823,N_15958);
nand U16193 (N_16193,N_15803,N_15808);
nor U16194 (N_16194,N_15968,N_15902);
xnor U16195 (N_16195,N_15905,N_15881);
and U16196 (N_16196,N_15871,N_15842);
or U16197 (N_16197,N_15933,N_15889);
nor U16198 (N_16198,N_15992,N_15914);
and U16199 (N_16199,N_15863,N_15876);
nor U16200 (N_16200,N_16175,N_16044);
or U16201 (N_16201,N_16180,N_16065);
and U16202 (N_16202,N_16128,N_16076);
nor U16203 (N_16203,N_16183,N_16169);
xor U16204 (N_16204,N_16164,N_16138);
xor U16205 (N_16205,N_16143,N_16016);
nand U16206 (N_16206,N_16093,N_16073);
and U16207 (N_16207,N_16012,N_16104);
and U16208 (N_16208,N_16032,N_16191);
and U16209 (N_16209,N_16075,N_16102);
and U16210 (N_16210,N_16148,N_16139);
xor U16211 (N_16211,N_16179,N_16052);
nor U16212 (N_16212,N_16094,N_16070);
and U16213 (N_16213,N_16092,N_16035);
nand U16214 (N_16214,N_16011,N_16066);
xor U16215 (N_16215,N_16170,N_16187);
xor U16216 (N_16216,N_16064,N_16025);
or U16217 (N_16217,N_16114,N_16178);
xor U16218 (N_16218,N_16033,N_16173);
xnor U16219 (N_16219,N_16054,N_16015);
and U16220 (N_16220,N_16026,N_16137);
nand U16221 (N_16221,N_16000,N_16156);
xor U16222 (N_16222,N_16067,N_16113);
or U16223 (N_16223,N_16023,N_16136);
or U16224 (N_16224,N_16184,N_16106);
or U16225 (N_16225,N_16043,N_16101);
or U16226 (N_16226,N_16182,N_16154);
or U16227 (N_16227,N_16071,N_16135);
nor U16228 (N_16228,N_16057,N_16091);
nand U16229 (N_16229,N_16022,N_16116);
nand U16230 (N_16230,N_16125,N_16149);
and U16231 (N_16231,N_16047,N_16181);
xor U16232 (N_16232,N_16050,N_16155);
nor U16233 (N_16233,N_16079,N_16074);
and U16234 (N_16234,N_16053,N_16009);
xor U16235 (N_16235,N_16157,N_16172);
nand U16236 (N_16236,N_16083,N_16163);
xnor U16237 (N_16237,N_16002,N_16100);
xor U16238 (N_16238,N_16099,N_16122);
and U16239 (N_16239,N_16115,N_16048);
or U16240 (N_16240,N_16124,N_16121);
and U16241 (N_16241,N_16123,N_16039);
xor U16242 (N_16242,N_16008,N_16117);
and U16243 (N_16243,N_16186,N_16086);
or U16244 (N_16244,N_16001,N_16013);
nor U16245 (N_16245,N_16177,N_16142);
nand U16246 (N_16246,N_16072,N_16061);
xor U16247 (N_16247,N_16078,N_16188);
nor U16248 (N_16248,N_16108,N_16165);
xnor U16249 (N_16249,N_16036,N_16063);
nor U16250 (N_16250,N_16021,N_16162);
and U16251 (N_16251,N_16112,N_16040);
nand U16252 (N_16252,N_16062,N_16046);
or U16253 (N_16253,N_16151,N_16107);
nand U16254 (N_16254,N_16185,N_16174);
and U16255 (N_16255,N_16084,N_16118);
or U16256 (N_16256,N_16027,N_16031);
nor U16257 (N_16257,N_16127,N_16134);
xnor U16258 (N_16258,N_16131,N_16176);
nor U16259 (N_16259,N_16029,N_16006);
nor U16260 (N_16260,N_16194,N_16005);
and U16261 (N_16261,N_16049,N_16171);
or U16262 (N_16262,N_16017,N_16147);
and U16263 (N_16263,N_16037,N_16056);
nand U16264 (N_16264,N_16069,N_16024);
nor U16265 (N_16265,N_16130,N_16095);
or U16266 (N_16266,N_16119,N_16019);
xnor U16267 (N_16267,N_16028,N_16018);
nand U16268 (N_16268,N_16198,N_16080);
nand U16269 (N_16269,N_16193,N_16197);
and U16270 (N_16270,N_16158,N_16051);
nand U16271 (N_16271,N_16068,N_16153);
xnor U16272 (N_16272,N_16089,N_16189);
or U16273 (N_16273,N_16110,N_16190);
and U16274 (N_16274,N_16098,N_16034);
nor U16275 (N_16275,N_16133,N_16003);
or U16276 (N_16276,N_16140,N_16146);
nand U16277 (N_16277,N_16060,N_16103);
nor U16278 (N_16278,N_16097,N_16141);
xor U16279 (N_16279,N_16042,N_16120);
xor U16280 (N_16280,N_16010,N_16087);
nor U16281 (N_16281,N_16196,N_16109);
and U16282 (N_16282,N_16159,N_16090);
nor U16283 (N_16283,N_16105,N_16161);
nor U16284 (N_16284,N_16077,N_16055);
or U16285 (N_16285,N_16088,N_16038);
nor U16286 (N_16286,N_16058,N_16132);
or U16287 (N_16287,N_16007,N_16192);
or U16288 (N_16288,N_16195,N_16004);
or U16289 (N_16289,N_16045,N_16082);
or U16290 (N_16290,N_16014,N_16041);
nand U16291 (N_16291,N_16126,N_16085);
or U16292 (N_16292,N_16167,N_16145);
nor U16293 (N_16293,N_16096,N_16111);
xnor U16294 (N_16294,N_16166,N_16059);
xnor U16295 (N_16295,N_16129,N_16020);
nand U16296 (N_16296,N_16150,N_16030);
nand U16297 (N_16297,N_16144,N_16160);
and U16298 (N_16298,N_16199,N_16152);
xor U16299 (N_16299,N_16168,N_16081);
and U16300 (N_16300,N_16193,N_16071);
nand U16301 (N_16301,N_16091,N_16112);
nand U16302 (N_16302,N_16065,N_16052);
nor U16303 (N_16303,N_16160,N_16161);
nor U16304 (N_16304,N_16173,N_16020);
nor U16305 (N_16305,N_16099,N_16199);
or U16306 (N_16306,N_16199,N_16048);
nor U16307 (N_16307,N_16067,N_16028);
and U16308 (N_16308,N_16127,N_16095);
xor U16309 (N_16309,N_16172,N_16186);
or U16310 (N_16310,N_16132,N_16188);
or U16311 (N_16311,N_16194,N_16017);
nor U16312 (N_16312,N_16158,N_16159);
and U16313 (N_16313,N_16151,N_16042);
and U16314 (N_16314,N_16183,N_16167);
or U16315 (N_16315,N_16017,N_16108);
or U16316 (N_16316,N_16125,N_16008);
nor U16317 (N_16317,N_16154,N_16108);
xor U16318 (N_16318,N_16144,N_16107);
or U16319 (N_16319,N_16080,N_16076);
or U16320 (N_16320,N_16194,N_16004);
or U16321 (N_16321,N_16060,N_16181);
xnor U16322 (N_16322,N_16068,N_16033);
xnor U16323 (N_16323,N_16045,N_16068);
nand U16324 (N_16324,N_16179,N_16061);
xor U16325 (N_16325,N_16013,N_16042);
nand U16326 (N_16326,N_16089,N_16142);
or U16327 (N_16327,N_16198,N_16019);
and U16328 (N_16328,N_16052,N_16049);
nand U16329 (N_16329,N_16051,N_16029);
and U16330 (N_16330,N_16034,N_16170);
or U16331 (N_16331,N_16054,N_16043);
xor U16332 (N_16332,N_16005,N_16199);
nand U16333 (N_16333,N_16037,N_16011);
nor U16334 (N_16334,N_16159,N_16038);
nor U16335 (N_16335,N_16191,N_16017);
or U16336 (N_16336,N_16151,N_16193);
nor U16337 (N_16337,N_16115,N_16127);
nand U16338 (N_16338,N_16110,N_16123);
and U16339 (N_16339,N_16089,N_16038);
xor U16340 (N_16340,N_16153,N_16196);
nor U16341 (N_16341,N_16135,N_16016);
or U16342 (N_16342,N_16160,N_16072);
nor U16343 (N_16343,N_16097,N_16154);
and U16344 (N_16344,N_16053,N_16046);
nor U16345 (N_16345,N_16164,N_16019);
xor U16346 (N_16346,N_16111,N_16050);
nor U16347 (N_16347,N_16036,N_16061);
xnor U16348 (N_16348,N_16094,N_16001);
or U16349 (N_16349,N_16148,N_16100);
and U16350 (N_16350,N_16197,N_16175);
nor U16351 (N_16351,N_16013,N_16090);
nor U16352 (N_16352,N_16082,N_16056);
nor U16353 (N_16353,N_16005,N_16163);
or U16354 (N_16354,N_16177,N_16147);
nor U16355 (N_16355,N_16168,N_16133);
nand U16356 (N_16356,N_16047,N_16085);
and U16357 (N_16357,N_16099,N_16143);
or U16358 (N_16358,N_16121,N_16152);
xor U16359 (N_16359,N_16013,N_16040);
xor U16360 (N_16360,N_16060,N_16121);
xnor U16361 (N_16361,N_16095,N_16100);
nand U16362 (N_16362,N_16182,N_16132);
or U16363 (N_16363,N_16193,N_16184);
nand U16364 (N_16364,N_16149,N_16054);
nand U16365 (N_16365,N_16177,N_16148);
nor U16366 (N_16366,N_16142,N_16123);
nand U16367 (N_16367,N_16144,N_16141);
xnor U16368 (N_16368,N_16037,N_16069);
xnor U16369 (N_16369,N_16034,N_16100);
nor U16370 (N_16370,N_16163,N_16075);
and U16371 (N_16371,N_16068,N_16187);
xor U16372 (N_16372,N_16072,N_16028);
and U16373 (N_16373,N_16158,N_16194);
xnor U16374 (N_16374,N_16175,N_16055);
or U16375 (N_16375,N_16192,N_16085);
xor U16376 (N_16376,N_16004,N_16028);
or U16377 (N_16377,N_16071,N_16138);
or U16378 (N_16378,N_16008,N_16082);
or U16379 (N_16379,N_16066,N_16019);
or U16380 (N_16380,N_16015,N_16031);
and U16381 (N_16381,N_16183,N_16080);
or U16382 (N_16382,N_16021,N_16020);
nand U16383 (N_16383,N_16193,N_16107);
and U16384 (N_16384,N_16088,N_16194);
and U16385 (N_16385,N_16107,N_16059);
nand U16386 (N_16386,N_16108,N_16069);
or U16387 (N_16387,N_16136,N_16017);
nand U16388 (N_16388,N_16089,N_16004);
nand U16389 (N_16389,N_16049,N_16096);
or U16390 (N_16390,N_16109,N_16067);
xnor U16391 (N_16391,N_16025,N_16063);
and U16392 (N_16392,N_16038,N_16195);
and U16393 (N_16393,N_16135,N_16040);
nor U16394 (N_16394,N_16130,N_16046);
or U16395 (N_16395,N_16118,N_16119);
nand U16396 (N_16396,N_16016,N_16183);
and U16397 (N_16397,N_16166,N_16110);
nor U16398 (N_16398,N_16124,N_16118);
or U16399 (N_16399,N_16081,N_16051);
nor U16400 (N_16400,N_16229,N_16348);
xor U16401 (N_16401,N_16356,N_16231);
nor U16402 (N_16402,N_16233,N_16268);
nor U16403 (N_16403,N_16363,N_16324);
nor U16404 (N_16404,N_16200,N_16395);
nor U16405 (N_16405,N_16206,N_16353);
xor U16406 (N_16406,N_16327,N_16323);
xor U16407 (N_16407,N_16252,N_16388);
nand U16408 (N_16408,N_16357,N_16301);
or U16409 (N_16409,N_16285,N_16373);
nor U16410 (N_16410,N_16251,N_16276);
nand U16411 (N_16411,N_16279,N_16397);
and U16412 (N_16412,N_16288,N_16396);
or U16413 (N_16413,N_16321,N_16326);
and U16414 (N_16414,N_16345,N_16267);
and U16415 (N_16415,N_16394,N_16307);
xor U16416 (N_16416,N_16383,N_16304);
nor U16417 (N_16417,N_16214,N_16314);
and U16418 (N_16418,N_16296,N_16305);
or U16419 (N_16419,N_16386,N_16256);
and U16420 (N_16420,N_16244,N_16259);
nor U16421 (N_16421,N_16202,N_16336);
xor U16422 (N_16422,N_16366,N_16333);
and U16423 (N_16423,N_16207,N_16220);
xnor U16424 (N_16424,N_16315,N_16219);
and U16425 (N_16425,N_16349,N_16230);
nor U16426 (N_16426,N_16216,N_16380);
nor U16427 (N_16427,N_16215,N_16280);
nor U16428 (N_16428,N_16350,N_16303);
or U16429 (N_16429,N_16302,N_16300);
or U16430 (N_16430,N_16275,N_16289);
nor U16431 (N_16431,N_16254,N_16360);
and U16432 (N_16432,N_16311,N_16375);
nand U16433 (N_16433,N_16266,N_16271);
xor U16434 (N_16434,N_16330,N_16298);
nor U16435 (N_16435,N_16261,N_16218);
nor U16436 (N_16436,N_16378,N_16212);
nand U16437 (N_16437,N_16258,N_16299);
nor U16438 (N_16438,N_16263,N_16234);
nand U16439 (N_16439,N_16293,N_16253);
nand U16440 (N_16440,N_16269,N_16379);
and U16441 (N_16441,N_16203,N_16309);
or U16442 (N_16442,N_16284,N_16328);
xnor U16443 (N_16443,N_16354,N_16381);
nor U16444 (N_16444,N_16246,N_16255);
or U16445 (N_16445,N_16260,N_16358);
xor U16446 (N_16446,N_16390,N_16376);
xnor U16447 (N_16447,N_16264,N_16338);
nand U16448 (N_16448,N_16274,N_16277);
or U16449 (N_16449,N_16295,N_16362);
or U16450 (N_16450,N_16243,N_16281);
and U16451 (N_16451,N_16290,N_16239);
nand U16452 (N_16452,N_16213,N_16292);
nand U16453 (N_16453,N_16398,N_16310);
and U16454 (N_16454,N_16232,N_16211);
xnor U16455 (N_16455,N_16225,N_16364);
xnor U16456 (N_16456,N_16312,N_16210);
nand U16457 (N_16457,N_16222,N_16365);
nor U16458 (N_16458,N_16369,N_16359);
nor U16459 (N_16459,N_16287,N_16331);
nand U16460 (N_16460,N_16238,N_16343);
nand U16461 (N_16461,N_16208,N_16313);
nor U16462 (N_16462,N_16329,N_16242);
xor U16463 (N_16463,N_16217,N_16372);
or U16464 (N_16464,N_16344,N_16387);
or U16465 (N_16465,N_16399,N_16248);
nand U16466 (N_16466,N_16283,N_16265);
nor U16467 (N_16467,N_16389,N_16235);
and U16468 (N_16468,N_16319,N_16316);
nand U16469 (N_16469,N_16392,N_16382);
nand U16470 (N_16470,N_16374,N_16250);
xor U16471 (N_16471,N_16337,N_16209);
nand U16472 (N_16472,N_16384,N_16332);
xor U16473 (N_16473,N_16236,N_16370);
xor U16474 (N_16474,N_16221,N_16393);
or U16475 (N_16475,N_16355,N_16291);
xor U16476 (N_16476,N_16371,N_16308);
nor U16477 (N_16477,N_16341,N_16247);
xnor U16478 (N_16478,N_16272,N_16385);
nor U16479 (N_16479,N_16270,N_16205);
nor U16480 (N_16480,N_16294,N_16347);
nand U16481 (N_16481,N_16377,N_16237);
nor U16482 (N_16482,N_16361,N_16335);
nand U16483 (N_16483,N_16262,N_16367);
and U16484 (N_16484,N_16322,N_16273);
nor U16485 (N_16485,N_16339,N_16278);
or U16486 (N_16486,N_16224,N_16340);
xnor U16487 (N_16487,N_16342,N_16257);
xnor U16488 (N_16488,N_16201,N_16282);
and U16489 (N_16489,N_16286,N_16334);
nand U16490 (N_16490,N_16223,N_16351);
nand U16491 (N_16491,N_16306,N_16346);
nand U16492 (N_16492,N_16318,N_16245);
xor U16493 (N_16493,N_16226,N_16352);
or U16494 (N_16494,N_16241,N_16204);
and U16495 (N_16495,N_16320,N_16391);
and U16496 (N_16496,N_16297,N_16240);
nor U16497 (N_16497,N_16317,N_16227);
and U16498 (N_16498,N_16325,N_16368);
xor U16499 (N_16499,N_16228,N_16249);
nor U16500 (N_16500,N_16379,N_16357);
xnor U16501 (N_16501,N_16338,N_16269);
xnor U16502 (N_16502,N_16227,N_16313);
or U16503 (N_16503,N_16339,N_16377);
nor U16504 (N_16504,N_16255,N_16312);
nand U16505 (N_16505,N_16244,N_16206);
xnor U16506 (N_16506,N_16330,N_16221);
and U16507 (N_16507,N_16229,N_16394);
xor U16508 (N_16508,N_16370,N_16287);
xnor U16509 (N_16509,N_16203,N_16315);
nor U16510 (N_16510,N_16354,N_16281);
or U16511 (N_16511,N_16240,N_16339);
nand U16512 (N_16512,N_16267,N_16287);
and U16513 (N_16513,N_16363,N_16248);
and U16514 (N_16514,N_16391,N_16246);
nor U16515 (N_16515,N_16242,N_16382);
or U16516 (N_16516,N_16281,N_16218);
nor U16517 (N_16517,N_16220,N_16293);
xor U16518 (N_16518,N_16255,N_16279);
nand U16519 (N_16519,N_16230,N_16279);
xor U16520 (N_16520,N_16260,N_16223);
and U16521 (N_16521,N_16329,N_16385);
or U16522 (N_16522,N_16345,N_16382);
nor U16523 (N_16523,N_16228,N_16312);
nor U16524 (N_16524,N_16363,N_16314);
or U16525 (N_16525,N_16328,N_16301);
nand U16526 (N_16526,N_16314,N_16343);
or U16527 (N_16527,N_16289,N_16283);
nand U16528 (N_16528,N_16298,N_16321);
or U16529 (N_16529,N_16319,N_16363);
xor U16530 (N_16530,N_16375,N_16255);
or U16531 (N_16531,N_16361,N_16255);
or U16532 (N_16532,N_16346,N_16215);
and U16533 (N_16533,N_16372,N_16227);
and U16534 (N_16534,N_16385,N_16285);
or U16535 (N_16535,N_16347,N_16261);
xnor U16536 (N_16536,N_16333,N_16290);
or U16537 (N_16537,N_16352,N_16375);
xnor U16538 (N_16538,N_16202,N_16344);
nor U16539 (N_16539,N_16301,N_16260);
xnor U16540 (N_16540,N_16256,N_16329);
or U16541 (N_16541,N_16326,N_16399);
nand U16542 (N_16542,N_16213,N_16309);
nor U16543 (N_16543,N_16293,N_16379);
nor U16544 (N_16544,N_16306,N_16328);
xor U16545 (N_16545,N_16330,N_16228);
xnor U16546 (N_16546,N_16309,N_16305);
or U16547 (N_16547,N_16285,N_16272);
nand U16548 (N_16548,N_16220,N_16231);
nand U16549 (N_16549,N_16329,N_16276);
nand U16550 (N_16550,N_16300,N_16235);
nand U16551 (N_16551,N_16322,N_16355);
nor U16552 (N_16552,N_16260,N_16321);
or U16553 (N_16553,N_16207,N_16244);
xor U16554 (N_16554,N_16297,N_16238);
and U16555 (N_16555,N_16383,N_16227);
or U16556 (N_16556,N_16261,N_16206);
and U16557 (N_16557,N_16248,N_16210);
xnor U16558 (N_16558,N_16294,N_16348);
nor U16559 (N_16559,N_16258,N_16202);
xor U16560 (N_16560,N_16204,N_16287);
and U16561 (N_16561,N_16332,N_16316);
or U16562 (N_16562,N_16386,N_16346);
and U16563 (N_16563,N_16302,N_16249);
or U16564 (N_16564,N_16380,N_16266);
xnor U16565 (N_16565,N_16216,N_16267);
and U16566 (N_16566,N_16243,N_16313);
and U16567 (N_16567,N_16365,N_16304);
and U16568 (N_16568,N_16354,N_16224);
nor U16569 (N_16569,N_16206,N_16228);
and U16570 (N_16570,N_16289,N_16201);
or U16571 (N_16571,N_16234,N_16366);
and U16572 (N_16572,N_16334,N_16387);
nor U16573 (N_16573,N_16266,N_16298);
nand U16574 (N_16574,N_16363,N_16354);
nand U16575 (N_16575,N_16279,N_16388);
and U16576 (N_16576,N_16294,N_16288);
nand U16577 (N_16577,N_16218,N_16305);
or U16578 (N_16578,N_16378,N_16328);
or U16579 (N_16579,N_16389,N_16203);
xor U16580 (N_16580,N_16248,N_16344);
nor U16581 (N_16581,N_16356,N_16293);
nor U16582 (N_16582,N_16331,N_16244);
xnor U16583 (N_16583,N_16238,N_16200);
and U16584 (N_16584,N_16292,N_16330);
or U16585 (N_16585,N_16372,N_16329);
and U16586 (N_16586,N_16370,N_16309);
nor U16587 (N_16587,N_16399,N_16330);
nand U16588 (N_16588,N_16278,N_16243);
xor U16589 (N_16589,N_16232,N_16270);
xor U16590 (N_16590,N_16244,N_16322);
or U16591 (N_16591,N_16311,N_16248);
nand U16592 (N_16592,N_16252,N_16381);
nand U16593 (N_16593,N_16378,N_16391);
or U16594 (N_16594,N_16213,N_16283);
xnor U16595 (N_16595,N_16303,N_16209);
or U16596 (N_16596,N_16257,N_16362);
or U16597 (N_16597,N_16219,N_16217);
or U16598 (N_16598,N_16204,N_16253);
and U16599 (N_16599,N_16312,N_16248);
xnor U16600 (N_16600,N_16405,N_16452);
xor U16601 (N_16601,N_16522,N_16467);
or U16602 (N_16602,N_16581,N_16562);
xnor U16603 (N_16603,N_16520,N_16457);
nand U16604 (N_16604,N_16535,N_16404);
nor U16605 (N_16605,N_16545,N_16560);
nor U16606 (N_16606,N_16556,N_16519);
nand U16607 (N_16607,N_16466,N_16420);
or U16608 (N_16608,N_16547,N_16568);
and U16609 (N_16609,N_16448,N_16505);
xnor U16610 (N_16610,N_16591,N_16550);
and U16611 (N_16611,N_16496,N_16412);
xnor U16612 (N_16612,N_16436,N_16504);
nor U16613 (N_16613,N_16426,N_16423);
or U16614 (N_16614,N_16461,N_16416);
nand U16615 (N_16615,N_16417,N_16469);
or U16616 (N_16616,N_16512,N_16418);
xor U16617 (N_16617,N_16538,N_16422);
or U16618 (N_16618,N_16566,N_16493);
nand U16619 (N_16619,N_16518,N_16557);
and U16620 (N_16620,N_16433,N_16454);
xor U16621 (N_16621,N_16577,N_16587);
xor U16622 (N_16622,N_16553,N_16530);
nor U16623 (N_16623,N_16597,N_16567);
or U16624 (N_16624,N_16424,N_16470);
nor U16625 (N_16625,N_16491,N_16528);
nor U16626 (N_16626,N_16419,N_16584);
xor U16627 (N_16627,N_16532,N_16589);
nor U16628 (N_16628,N_16576,N_16438);
and U16629 (N_16629,N_16571,N_16552);
nand U16630 (N_16630,N_16445,N_16435);
and U16631 (N_16631,N_16427,N_16558);
nand U16632 (N_16632,N_16511,N_16430);
nor U16633 (N_16633,N_16506,N_16563);
nor U16634 (N_16634,N_16437,N_16569);
xnor U16635 (N_16635,N_16462,N_16514);
nand U16636 (N_16636,N_16573,N_16513);
xnor U16637 (N_16637,N_16549,N_16486);
xor U16638 (N_16638,N_16559,N_16451);
nand U16639 (N_16639,N_16555,N_16421);
or U16640 (N_16640,N_16444,N_16543);
xnor U16641 (N_16641,N_16510,N_16551);
nand U16642 (N_16642,N_16459,N_16482);
and U16643 (N_16643,N_16585,N_16400);
and U16644 (N_16644,N_16494,N_16484);
nand U16645 (N_16645,N_16490,N_16471);
and U16646 (N_16646,N_16453,N_16432);
or U16647 (N_16647,N_16402,N_16447);
xnor U16648 (N_16648,N_16594,N_16565);
nand U16649 (N_16649,N_16578,N_16546);
xnor U16650 (N_16650,N_16595,N_16431);
xnor U16651 (N_16651,N_16596,N_16521);
nand U16652 (N_16652,N_16598,N_16499);
xnor U16653 (N_16653,N_16586,N_16542);
nand U16654 (N_16654,N_16411,N_16570);
xnor U16655 (N_16655,N_16472,N_16475);
nand U16656 (N_16656,N_16561,N_16536);
and U16657 (N_16657,N_16502,N_16582);
xnor U16658 (N_16658,N_16401,N_16523);
and U16659 (N_16659,N_16503,N_16409);
xor U16660 (N_16660,N_16410,N_16537);
xnor U16661 (N_16661,N_16554,N_16548);
and U16662 (N_16662,N_16516,N_16439);
nor U16663 (N_16663,N_16440,N_16458);
and U16664 (N_16664,N_16413,N_16478);
xnor U16665 (N_16665,N_16474,N_16500);
nor U16666 (N_16666,N_16464,N_16534);
and U16667 (N_16667,N_16477,N_16524);
nor U16668 (N_16668,N_16443,N_16429);
and U16669 (N_16669,N_16495,N_16509);
xnor U16670 (N_16670,N_16599,N_16476);
nand U16671 (N_16671,N_16468,N_16480);
or U16672 (N_16672,N_16592,N_16407);
and U16673 (N_16673,N_16408,N_16580);
or U16674 (N_16674,N_16415,N_16485);
xnor U16675 (N_16675,N_16434,N_16406);
and U16676 (N_16676,N_16526,N_16446);
nand U16677 (N_16677,N_16465,N_16481);
xor U16678 (N_16678,N_16489,N_16539);
nand U16679 (N_16679,N_16492,N_16583);
and U16680 (N_16680,N_16479,N_16593);
xnor U16681 (N_16681,N_16574,N_16442);
nor U16682 (N_16682,N_16428,N_16487);
xor U16683 (N_16683,N_16527,N_16507);
xor U16684 (N_16684,N_16541,N_16540);
xnor U16685 (N_16685,N_16441,N_16414);
xor U16686 (N_16686,N_16517,N_16403);
xnor U16687 (N_16687,N_16588,N_16590);
xnor U16688 (N_16688,N_16460,N_16473);
xor U16689 (N_16689,N_16544,N_16501);
nor U16690 (N_16690,N_16533,N_16497);
xor U16691 (N_16691,N_16498,N_16575);
or U16692 (N_16692,N_16525,N_16455);
nand U16693 (N_16693,N_16572,N_16564);
nor U16694 (N_16694,N_16508,N_16450);
nand U16695 (N_16695,N_16425,N_16488);
nor U16696 (N_16696,N_16579,N_16456);
nor U16697 (N_16697,N_16529,N_16515);
and U16698 (N_16698,N_16463,N_16531);
and U16699 (N_16699,N_16449,N_16483);
nor U16700 (N_16700,N_16554,N_16445);
or U16701 (N_16701,N_16515,N_16490);
xnor U16702 (N_16702,N_16484,N_16512);
nor U16703 (N_16703,N_16451,N_16558);
or U16704 (N_16704,N_16499,N_16595);
or U16705 (N_16705,N_16408,N_16412);
xnor U16706 (N_16706,N_16469,N_16484);
nor U16707 (N_16707,N_16590,N_16595);
nor U16708 (N_16708,N_16568,N_16401);
nand U16709 (N_16709,N_16564,N_16448);
nor U16710 (N_16710,N_16421,N_16551);
or U16711 (N_16711,N_16594,N_16441);
nand U16712 (N_16712,N_16458,N_16491);
and U16713 (N_16713,N_16459,N_16594);
nand U16714 (N_16714,N_16561,N_16568);
and U16715 (N_16715,N_16530,N_16575);
nor U16716 (N_16716,N_16475,N_16588);
nand U16717 (N_16717,N_16455,N_16421);
or U16718 (N_16718,N_16449,N_16460);
or U16719 (N_16719,N_16518,N_16595);
or U16720 (N_16720,N_16427,N_16406);
nor U16721 (N_16721,N_16531,N_16527);
or U16722 (N_16722,N_16448,N_16569);
xnor U16723 (N_16723,N_16424,N_16456);
nor U16724 (N_16724,N_16504,N_16587);
and U16725 (N_16725,N_16562,N_16542);
xnor U16726 (N_16726,N_16443,N_16596);
and U16727 (N_16727,N_16568,N_16541);
or U16728 (N_16728,N_16482,N_16450);
nand U16729 (N_16729,N_16533,N_16428);
xor U16730 (N_16730,N_16593,N_16429);
or U16731 (N_16731,N_16513,N_16412);
nor U16732 (N_16732,N_16445,N_16493);
or U16733 (N_16733,N_16515,N_16545);
nand U16734 (N_16734,N_16592,N_16581);
xor U16735 (N_16735,N_16517,N_16417);
or U16736 (N_16736,N_16485,N_16458);
or U16737 (N_16737,N_16515,N_16462);
nor U16738 (N_16738,N_16459,N_16548);
xor U16739 (N_16739,N_16599,N_16438);
and U16740 (N_16740,N_16546,N_16455);
or U16741 (N_16741,N_16429,N_16584);
and U16742 (N_16742,N_16469,N_16588);
nand U16743 (N_16743,N_16427,N_16567);
xor U16744 (N_16744,N_16588,N_16439);
nor U16745 (N_16745,N_16474,N_16590);
xor U16746 (N_16746,N_16495,N_16405);
or U16747 (N_16747,N_16593,N_16468);
nor U16748 (N_16748,N_16421,N_16552);
and U16749 (N_16749,N_16583,N_16459);
nor U16750 (N_16750,N_16435,N_16425);
and U16751 (N_16751,N_16480,N_16587);
nand U16752 (N_16752,N_16509,N_16583);
or U16753 (N_16753,N_16500,N_16565);
nor U16754 (N_16754,N_16415,N_16403);
nand U16755 (N_16755,N_16545,N_16565);
nand U16756 (N_16756,N_16438,N_16505);
and U16757 (N_16757,N_16578,N_16565);
or U16758 (N_16758,N_16513,N_16514);
nand U16759 (N_16759,N_16458,N_16564);
nor U16760 (N_16760,N_16455,N_16559);
or U16761 (N_16761,N_16574,N_16571);
xor U16762 (N_16762,N_16507,N_16441);
or U16763 (N_16763,N_16492,N_16438);
and U16764 (N_16764,N_16412,N_16464);
nand U16765 (N_16765,N_16423,N_16540);
nor U16766 (N_16766,N_16530,N_16582);
nand U16767 (N_16767,N_16508,N_16431);
or U16768 (N_16768,N_16573,N_16461);
nor U16769 (N_16769,N_16598,N_16490);
or U16770 (N_16770,N_16545,N_16569);
and U16771 (N_16771,N_16480,N_16534);
nand U16772 (N_16772,N_16426,N_16538);
nor U16773 (N_16773,N_16586,N_16446);
nor U16774 (N_16774,N_16489,N_16594);
or U16775 (N_16775,N_16409,N_16523);
nor U16776 (N_16776,N_16575,N_16468);
or U16777 (N_16777,N_16427,N_16481);
xor U16778 (N_16778,N_16401,N_16452);
nand U16779 (N_16779,N_16535,N_16568);
or U16780 (N_16780,N_16572,N_16467);
or U16781 (N_16781,N_16505,N_16479);
and U16782 (N_16782,N_16420,N_16535);
and U16783 (N_16783,N_16574,N_16436);
or U16784 (N_16784,N_16544,N_16448);
xnor U16785 (N_16785,N_16449,N_16497);
and U16786 (N_16786,N_16476,N_16583);
xnor U16787 (N_16787,N_16431,N_16451);
or U16788 (N_16788,N_16469,N_16404);
and U16789 (N_16789,N_16569,N_16519);
or U16790 (N_16790,N_16491,N_16429);
nor U16791 (N_16791,N_16595,N_16514);
nor U16792 (N_16792,N_16527,N_16523);
and U16793 (N_16793,N_16576,N_16479);
and U16794 (N_16794,N_16435,N_16530);
and U16795 (N_16795,N_16580,N_16558);
nand U16796 (N_16796,N_16535,N_16491);
nand U16797 (N_16797,N_16415,N_16452);
nand U16798 (N_16798,N_16582,N_16537);
xor U16799 (N_16799,N_16544,N_16413);
and U16800 (N_16800,N_16708,N_16733);
nor U16801 (N_16801,N_16687,N_16744);
xor U16802 (N_16802,N_16635,N_16686);
xor U16803 (N_16803,N_16767,N_16717);
xor U16804 (N_16804,N_16722,N_16702);
nor U16805 (N_16805,N_16757,N_16704);
or U16806 (N_16806,N_16720,N_16657);
xor U16807 (N_16807,N_16667,N_16798);
xnor U16808 (N_16808,N_16713,N_16771);
nand U16809 (N_16809,N_16616,N_16602);
and U16810 (N_16810,N_16731,N_16628);
and U16811 (N_16811,N_16673,N_16745);
and U16812 (N_16812,N_16754,N_16759);
and U16813 (N_16813,N_16659,N_16793);
nand U16814 (N_16814,N_16703,N_16625);
xnor U16815 (N_16815,N_16640,N_16753);
or U16816 (N_16816,N_16768,N_16651);
nor U16817 (N_16817,N_16648,N_16697);
and U16818 (N_16818,N_16791,N_16779);
xnor U16819 (N_16819,N_16658,N_16799);
nor U16820 (N_16820,N_16626,N_16780);
nand U16821 (N_16821,N_16634,N_16642);
xor U16822 (N_16822,N_16775,N_16674);
xor U16823 (N_16823,N_16706,N_16665);
xor U16824 (N_16824,N_16772,N_16756);
and U16825 (N_16825,N_16668,N_16617);
nand U16826 (N_16826,N_16664,N_16699);
xnor U16827 (N_16827,N_16661,N_16607);
nand U16828 (N_16828,N_16789,N_16794);
nor U16829 (N_16829,N_16654,N_16729);
or U16830 (N_16830,N_16777,N_16620);
and U16831 (N_16831,N_16709,N_16695);
xnor U16832 (N_16832,N_16646,N_16601);
xor U16833 (N_16833,N_16726,N_16685);
xnor U16834 (N_16834,N_16688,N_16751);
and U16835 (N_16835,N_16638,N_16630);
xor U16836 (N_16836,N_16752,N_16636);
and U16837 (N_16837,N_16747,N_16740);
and U16838 (N_16838,N_16797,N_16623);
xor U16839 (N_16839,N_16749,N_16608);
nand U16840 (N_16840,N_16762,N_16641);
and U16841 (N_16841,N_16715,N_16725);
or U16842 (N_16842,N_16766,N_16770);
or U16843 (N_16843,N_16711,N_16652);
or U16844 (N_16844,N_16790,N_16684);
nor U16845 (N_16845,N_16691,N_16796);
nand U16846 (N_16846,N_16619,N_16627);
xnor U16847 (N_16847,N_16765,N_16693);
nand U16848 (N_16848,N_16716,N_16610);
nor U16849 (N_16849,N_16776,N_16644);
and U16850 (N_16850,N_16622,N_16750);
xor U16851 (N_16851,N_16730,N_16707);
or U16852 (N_16852,N_16727,N_16660);
and U16853 (N_16853,N_16633,N_16643);
xnor U16854 (N_16854,N_16795,N_16738);
or U16855 (N_16855,N_16662,N_16792);
nand U16856 (N_16856,N_16786,N_16624);
nand U16857 (N_16857,N_16788,N_16632);
or U16858 (N_16858,N_16676,N_16618);
and U16859 (N_16859,N_16782,N_16672);
nor U16860 (N_16860,N_16677,N_16760);
or U16861 (N_16861,N_16600,N_16721);
nor U16862 (N_16862,N_16647,N_16783);
nand U16863 (N_16863,N_16714,N_16696);
nor U16864 (N_16864,N_16764,N_16778);
xnor U16865 (N_16865,N_16774,N_16604);
and U16866 (N_16866,N_16653,N_16737);
nor U16867 (N_16867,N_16690,N_16736);
nor U16868 (N_16868,N_16781,N_16773);
and U16869 (N_16869,N_16631,N_16732);
and U16870 (N_16870,N_16718,N_16629);
or U16871 (N_16871,N_16621,N_16615);
xor U16872 (N_16872,N_16694,N_16769);
or U16873 (N_16873,N_16785,N_16758);
and U16874 (N_16874,N_16606,N_16612);
nand U16875 (N_16875,N_16755,N_16650);
and U16876 (N_16876,N_16719,N_16671);
and U16877 (N_16877,N_16700,N_16698);
nor U16878 (N_16878,N_16739,N_16603);
or U16879 (N_16879,N_16675,N_16689);
nand U16880 (N_16880,N_16746,N_16614);
and U16881 (N_16881,N_16763,N_16639);
nor U16882 (N_16882,N_16743,N_16681);
nor U16883 (N_16883,N_16613,N_16741);
and U16884 (N_16884,N_16712,N_16680);
and U16885 (N_16885,N_16655,N_16666);
nand U16886 (N_16886,N_16742,N_16649);
or U16887 (N_16887,N_16605,N_16682);
nand U16888 (N_16888,N_16663,N_16701);
xor U16889 (N_16889,N_16679,N_16710);
nor U16890 (N_16890,N_16670,N_16748);
or U16891 (N_16891,N_16637,N_16611);
nand U16892 (N_16892,N_16683,N_16787);
xor U16893 (N_16893,N_16645,N_16728);
nor U16894 (N_16894,N_16656,N_16724);
nor U16895 (N_16895,N_16678,N_16692);
or U16896 (N_16896,N_16735,N_16761);
and U16897 (N_16897,N_16784,N_16723);
xnor U16898 (N_16898,N_16609,N_16734);
nand U16899 (N_16899,N_16705,N_16669);
and U16900 (N_16900,N_16604,N_16615);
or U16901 (N_16901,N_16605,N_16769);
nor U16902 (N_16902,N_16729,N_16785);
or U16903 (N_16903,N_16726,N_16687);
xnor U16904 (N_16904,N_16745,N_16765);
nor U16905 (N_16905,N_16735,N_16634);
xor U16906 (N_16906,N_16611,N_16747);
xnor U16907 (N_16907,N_16646,N_16686);
nand U16908 (N_16908,N_16671,N_16667);
nor U16909 (N_16909,N_16614,N_16668);
nor U16910 (N_16910,N_16756,N_16660);
and U16911 (N_16911,N_16675,N_16600);
nand U16912 (N_16912,N_16770,N_16720);
or U16913 (N_16913,N_16786,N_16709);
nand U16914 (N_16914,N_16620,N_16644);
xor U16915 (N_16915,N_16733,N_16795);
xor U16916 (N_16916,N_16782,N_16787);
nor U16917 (N_16917,N_16782,N_16660);
nand U16918 (N_16918,N_16634,N_16682);
xor U16919 (N_16919,N_16682,N_16703);
nor U16920 (N_16920,N_16738,N_16780);
nand U16921 (N_16921,N_16755,N_16605);
or U16922 (N_16922,N_16786,N_16761);
or U16923 (N_16923,N_16641,N_16792);
nand U16924 (N_16924,N_16689,N_16709);
nand U16925 (N_16925,N_16718,N_16757);
nand U16926 (N_16926,N_16646,N_16684);
and U16927 (N_16927,N_16643,N_16612);
xor U16928 (N_16928,N_16600,N_16782);
nand U16929 (N_16929,N_16710,N_16732);
nor U16930 (N_16930,N_16615,N_16639);
nor U16931 (N_16931,N_16617,N_16662);
nor U16932 (N_16932,N_16685,N_16774);
and U16933 (N_16933,N_16751,N_16760);
nor U16934 (N_16934,N_16650,N_16630);
xnor U16935 (N_16935,N_16652,N_16700);
nand U16936 (N_16936,N_16708,N_16617);
and U16937 (N_16937,N_16638,N_16770);
nor U16938 (N_16938,N_16793,N_16785);
xor U16939 (N_16939,N_16747,N_16738);
nor U16940 (N_16940,N_16639,N_16745);
nand U16941 (N_16941,N_16793,N_16675);
nand U16942 (N_16942,N_16777,N_16692);
nand U16943 (N_16943,N_16617,N_16769);
nand U16944 (N_16944,N_16605,N_16618);
xnor U16945 (N_16945,N_16636,N_16624);
nor U16946 (N_16946,N_16765,N_16714);
nor U16947 (N_16947,N_16725,N_16773);
xor U16948 (N_16948,N_16740,N_16688);
xor U16949 (N_16949,N_16752,N_16720);
and U16950 (N_16950,N_16770,N_16655);
nand U16951 (N_16951,N_16789,N_16786);
nand U16952 (N_16952,N_16753,N_16614);
xnor U16953 (N_16953,N_16646,N_16657);
nand U16954 (N_16954,N_16720,N_16795);
or U16955 (N_16955,N_16715,N_16677);
xnor U16956 (N_16956,N_16766,N_16612);
nor U16957 (N_16957,N_16793,N_16614);
or U16958 (N_16958,N_16743,N_16768);
xnor U16959 (N_16959,N_16634,N_16664);
nand U16960 (N_16960,N_16779,N_16624);
nor U16961 (N_16961,N_16605,N_16712);
xnor U16962 (N_16962,N_16766,N_16760);
xnor U16963 (N_16963,N_16779,N_16781);
nand U16964 (N_16964,N_16638,N_16739);
nor U16965 (N_16965,N_16621,N_16780);
nor U16966 (N_16966,N_16782,N_16769);
xor U16967 (N_16967,N_16666,N_16708);
xor U16968 (N_16968,N_16641,N_16799);
or U16969 (N_16969,N_16667,N_16730);
nand U16970 (N_16970,N_16780,N_16684);
nand U16971 (N_16971,N_16610,N_16774);
xnor U16972 (N_16972,N_16631,N_16660);
or U16973 (N_16973,N_16756,N_16780);
xor U16974 (N_16974,N_16621,N_16619);
or U16975 (N_16975,N_16678,N_16682);
or U16976 (N_16976,N_16632,N_16764);
and U16977 (N_16977,N_16744,N_16608);
or U16978 (N_16978,N_16609,N_16788);
nor U16979 (N_16979,N_16795,N_16793);
and U16980 (N_16980,N_16620,N_16794);
nand U16981 (N_16981,N_16754,N_16657);
nor U16982 (N_16982,N_16751,N_16719);
xnor U16983 (N_16983,N_16698,N_16706);
nand U16984 (N_16984,N_16639,N_16691);
or U16985 (N_16985,N_16798,N_16790);
or U16986 (N_16986,N_16744,N_16695);
nor U16987 (N_16987,N_16791,N_16759);
or U16988 (N_16988,N_16773,N_16728);
or U16989 (N_16989,N_16648,N_16728);
or U16990 (N_16990,N_16625,N_16626);
xor U16991 (N_16991,N_16697,N_16617);
nor U16992 (N_16992,N_16757,N_16742);
or U16993 (N_16993,N_16761,N_16696);
nor U16994 (N_16994,N_16777,N_16682);
and U16995 (N_16995,N_16682,N_16662);
xnor U16996 (N_16996,N_16600,N_16655);
or U16997 (N_16997,N_16790,N_16611);
and U16998 (N_16998,N_16638,N_16718);
nor U16999 (N_16999,N_16612,N_16656);
xor U17000 (N_17000,N_16913,N_16882);
nand U17001 (N_17001,N_16829,N_16834);
xor U17002 (N_17002,N_16861,N_16864);
or U17003 (N_17003,N_16967,N_16963);
xor U17004 (N_17004,N_16927,N_16958);
or U17005 (N_17005,N_16803,N_16941);
nor U17006 (N_17006,N_16823,N_16966);
and U17007 (N_17007,N_16810,N_16935);
and U17008 (N_17008,N_16843,N_16868);
nor U17009 (N_17009,N_16859,N_16902);
and U17010 (N_17010,N_16897,N_16894);
nand U17011 (N_17011,N_16965,N_16855);
or U17012 (N_17012,N_16874,N_16920);
and U17013 (N_17013,N_16987,N_16943);
nor U17014 (N_17014,N_16817,N_16905);
and U17015 (N_17015,N_16995,N_16860);
xnor U17016 (N_17016,N_16901,N_16884);
nor U17017 (N_17017,N_16820,N_16858);
nand U17018 (N_17018,N_16994,N_16997);
xnor U17019 (N_17019,N_16947,N_16915);
nor U17020 (N_17020,N_16828,N_16937);
nand U17021 (N_17021,N_16989,N_16980);
and U17022 (N_17022,N_16856,N_16988);
nor U17023 (N_17023,N_16805,N_16951);
xor U17024 (N_17024,N_16887,N_16847);
xor U17025 (N_17025,N_16972,N_16993);
or U17026 (N_17026,N_16949,N_16996);
nor U17027 (N_17027,N_16835,N_16819);
nand U17028 (N_17028,N_16931,N_16890);
nand U17029 (N_17029,N_16886,N_16853);
nand U17030 (N_17030,N_16991,N_16973);
nand U17031 (N_17031,N_16986,N_16892);
or U17032 (N_17032,N_16909,N_16811);
and U17033 (N_17033,N_16812,N_16815);
nand U17034 (N_17034,N_16827,N_16969);
xor U17035 (N_17035,N_16844,N_16932);
or U17036 (N_17036,N_16830,N_16831);
or U17037 (N_17037,N_16875,N_16974);
nor U17038 (N_17038,N_16903,N_16910);
xnor U17039 (N_17039,N_16837,N_16857);
or U17040 (N_17040,N_16872,N_16977);
nand U17041 (N_17041,N_16880,N_16826);
nor U17042 (N_17042,N_16940,N_16804);
nor U17043 (N_17043,N_16992,N_16933);
nor U17044 (N_17044,N_16985,N_16982);
nor U17045 (N_17045,N_16816,N_16800);
or U17046 (N_17046,N_16961,N_16948);
nor U17047 (N_17047,N_16938,N_16968);
nor U17048 (N_17048,N_16833,N_16945);
or U17049 (N_17049,N_16984,N_16832);
nor U17050 (N_17050,N_16893,N_16962);
or U17051 (N_17051,N_16873,N_16824);
nand U17052 (N_17052,N_16900,N_16929);
nand U17053 (N_17053,N_16908,N_16990);
and U17054 (N_17054,N_16904,N_16952);
and U17055 (N_17055,N_16802,N_16923);
nor U17056 (N_17056,N_16975,N_16926);
and U17057 (N_17057,N_16906,N_16960);
xor U17058 (N_17058,N_16801,N_16976);
nor U17059 (N_17059,N_16881,N_16867);
nand U17060 (N_17060,N_16849,N_16955);
nor U17061 (N_17061,N_16877,N_16959);
or U17062 (N_17062,N_16865,N_16862);
xor U17063 (N_17063,N_16928,N_16939);
nand U17064 (N_17064,N_16848,N_16934);
nand U17065 (N_17065,N_16916,N_16979);
nand U17066 (N_17066,N_16813,N_16845);
and U17067 (N_17067,N_16889,N_16954);
nor U17068 (N_17068,N_16956,N_16871);
nor U17069 (N_17069,N_16891,N_16842);
nand U17070 (N_17070,N_16846,N_16888);
nand U17071 (N_17071,N_16869,N_16885);
nand U17072 (N_17072,N_16922,N_16838);
xor U17073 (N_17073,N_16912,N_16911);
nor U17074 (N_17074,N_16807,N_16852);
or U17075 (N_17075,N_16850,N_16925);
and U17076 (N_17076,N_16953,N_16821);
or U17077 (N_17077,N_16942,N_16814);
and U17078 (N_17078,N_16879,N_16919);
or U17079 (N_17079,N_16840,N_16918);
nor U17080 (N_17080,N_16978,N_16899);
nor U17081 (N_17081,N_16863,N_16883);
xor U17082 (N_17082,N_16998,N_16983);
and U17083 (N_17083,N_16896,N_16876);
xnor U17084 (N_17084,N_16878,N_16981);
or U17085 (N_17085,N_16870,N_16944);
nand U17086 (N_17086,N_16914,N_16921);
or U17087 (N_17087,N_16971,N_16808);
or U17088 (N_17088,N_16950,N_16907);
nor U17089 (N_17089,N_16836,N_16825);
nand U17090 (N_17090,N_16999,N_16917);
nor U17091 (N_17091,N_16806,N_16809);
xnor U17092 (N_17092,N_16957,N_16851);
nand U17093 (N_17093,N_16924,N_16866);
nor U17094 (N_17094,N_16970,N_16818);
or U17095 (N_17095,N_16930,N_16854);
or U17096 (N_17096,N_16936,N_16898);
and U17097 (N_17097,N_16895,N_16822);
nor U17098 (N_17098,N_16841,N_16946);
nand U17099 (N_17099,N_16839,N_16964);
or U17100 (N_17100,N_16807,N_16942);
nor U17101 (N_17101,N_16927,N_16947);
nor U17102 (N_17102,N_16927,N_16946);
and U17103 (N_17103,N_16865,N_16917);
xnor U17104 (N_17104,N_16833,N_16995);
nor U17105 (N_17105,N_16857,N_16800);
nand U17106 (N_17106,N_16855,N_16912);
and U17107 (N_17107,N_16847,N_16939);
xor U17108 (N_17108,N_16898,N_16877);
nor U17109 (N_17109,N_16816,N_16838);
xnor U17110 (N_17110,N_16955,N_16848);
nor U17111 (N_17111,N_16916,N_16993);
nand U17112 (N_17112,N_16842,N_16984);
or U17113 (N_17113,N_16906,N_16871);
or U17114 (N_17114,N_16821,N_16942);
and U17115 (N_17115,N_16917,N_16871);
and U17116 (N_17116,N_16855,N_16992);
nor U17117 (N_17117,N_16899,N_16989);
or U17118 (N_17118,N_16902,N_16932);
xnor U17119 (N_17119,N_16942,N_16911);
nor U17120 (N_17120,N_16858,N_16983);
xor U17121 (N_17121,N_16962,N_16859);
and U17122 (N_17122,N_16835,N_16881);
nand U17123 (N_17123,N_16972,N_16896);
xnor U17124 (N_17124,N_16908,N_16922);
and U17125 (N_17125,N_16944,N_16943);
xnor U17126 (N_17126,N_16990,N_16933);
xor U17127 (N_17127,N_16940,N_16851);
xor U17128 (N_17128,N_16808,N_16859);
or U17129 (N_17129,N_16935,N_16861);
nor U17130 (N_17130,N_16840,N_16845);
nand U17131 (N_17131,N_16877,N_16909);
or U17132 (N_17132,N_16919,N_16813);
nand U17133 (N_17133,N_16891,N_16910);
nand U17134 (N_17134,N_16998,N_16808);
and U17135 (N_17135,N_16861,N_16806);
or U17136 (N_17136,N_16995,N_16930);
and U17137 (N_17137,N_16929,N_16899);
and U17138 (N_17138,N_16879,N_16862);
nand U17139 (N_17139,N_16937,N_16986);
xnor U17140 (N_17140,N_16815,N_16836);
and U17141 (N_17141,N_16983,N_16862);
and U17142 (N_17142,N_16874,N_16903);
or U17143 (N_17143,N_16939,N_16982);
and U17144 (N_17144,N_16925,N_16912);
nor U17145 (N_17145,N_16928,N_16999);
nand U17146 (N_17146,N_16949,N_16807);
and U17147 (N_17147,N_16807,N_16872);
or U17148 (N_17148,N_16844,N_16945);
xor U17149 (N_17149,N_16991,N_16863);
xnor U17150 (N_17150,N_16867,N_16966);
nor U17151 (N_17151,N_16998,N_16942);
xnor U17152 (N_17152,N_16991,N_16994);
nand U17153 (N_17153,N_16987,N_16920);
or U17154 (N_17154,N_16921,N_16911);
and U17155 (N_17155,N_16973,N_16903);
or U17156 (N_17156,N_16910,N_16911);
nor U17157 (N_17157,N_16829,N_16896);
or U17158 (N_17158,N_16809,N_16978);
or U17159 (N_17159,N_16872,N_16958);
xnor U17160 (N_17160,N_16831,N_16821);
xnor U17161 (N_17161,N_16862,N_16803);
or U17162 (N_17162,N_16946,N_16993);
nand U17163 (N_17163,N_16855,N_16850);
and U17164 (N_17164,N_16918,N_16845);
nor U17165 (N_17165,N_16879,N_16831);
nor U17166 (N_17166,N_16854,N_16993);
xnor U17167 (N_17167,N_16943,N_16925);
and U17168 (N_17168,N_16920,N_16995);
nor U17169 (N_17169,N_16919,N_16874);
xnor U17170 (N_17170,N_16816,N_16927);
nand U17171 (N_17171,N_16832,N_16853);
nand U17172 (N_17172,N_16835,N_16861);
xnor U17173 (N_17173,N_16911,N_16812);
or U17174 (N_17174,N_16825,N_16860);
xor U17175 (N_17175,N_16836,N_16813);
nand U17176 (N_17176,N_16885,N_16803);
and U17177 (N_17177,N_16931,N_16915);
or U17178 (N_17178,N_16919,N_16922);
or U17179 (N_17179,N_16919,N_16818);
xnor U17180 (N_17180,N_16831,N_16809);
nand U17181 (N_17181,N_16806,N_16919);
nand U17182 (N_17182,N_16806,N_16952);
xor U17183 (N_17183,N_16973,N_16823);
nor U17184 (N_17184,N_16861,N_16933);
or U17185 (N_17185,N_16822,N_16836);
nand U17186 (N_17186,N_16850,N_16984);
nor U17187 (N_17187,N_16973,N_16817);
nor U17188 (N_17188,N_16912,N_16981);
nand U17189 (N_17189,N_16996,N_16842);
xnor U17190 (N_17190,N_16878,N_16967);
nand U17191 (N_17191,N_16918,N_16960);
and U17192 (N_17192,N_16832,N_16908);
and U17193 (N_17193,N_16878,N_16950);
xnor U17194 (N_17194,N_16923,N_16820);
and U17195 (N_17195,N_16838,N_16899);
nand U17196 (N_17196,N_16901,N_16918);
or U17197 (N_17197,N_16965,N_16838);
or U17198 (N_17198,N_16845,N_16902);
and U17199 (N_17199,N_16894,N_16905);
and U17200 (N_17200,N_17095,N_17061);
or U17201 (N_17201,N_17060,N_17087);
or U17202 (N_17202,N_17049,N_17114);
xnor U17203 (N_17203,N_17057,N_17038);
and U17204 (N_17204,N_17159,N_17099);
and U17205 (N_17205,N_17163,N_17093);
or U17206 (N_17206,N_17071,N_17083);
nor U17207 (N_17207,N_17145,N_17023);
and U17208 (N_17208,N_17006,N_17096);
xor U17209 (N_17209,N_17183,N_17188);
or U17210 (N_17210,N_17115,N_17190);
or U17211 (N_17211,N_17170,N_17085);
or U17212 (N_17212,N_17008,N_17155);
nor U17213 (N_17213,N_17044,N_17091);
nand U17214 (N_17214,N_17147,N_17072);
and U17215 (N_17215,N_17162,N_17020);
nand U17216 (N_17216,N_17100,N_17131);
nand U17217 (N_17217,N_17033,N_17056);
nor U17218 (N_17218,N_17164,N_17053);
nand U17219 (N_17219,N_17019,N_17129);
and U17220 (N_17220,N_17180,N_17015);
and U17221 (N_17221,N_17154,N_17104);
and U17222 (N_17222,N_17030,N_17192);
nand U17223 (N_17223,N_17031,N_17181);
xor U17224 (N_17224,N_17141,N_17175);
or U17225 (N_17225,N_17042,N_17032);
nor U17226 (N_17226,N_17134,N_17011);
xor U17227 (N_17227,N_17149,N_17138);
and U17228 (N_17228,N_17121,N_17101);
and U17229 (N_17229,N_17078,N_17116);
xor U17230 (N_17230,N_17133,N_17172);
and U17231 (N_17231,N_17127,N_17080);
and U17232 (N_17232,N_17001,N_17022);
nand U17233 (N_17233,N_17045,N_17197);
nor U17234 (N_17234,N_17108,N_17055);
and U17235 (N_17235,N_17195,N_17140);
xnor U17236 (N_17236,N_17067,N_17184);
and U17237 (N_17237,N_17081,N_17107);
nor U17238 (N_17238,N_17089,N_17168);
or U17239 (N_17239,N_17028,N_17113);
nor U17240 (N_17240,N_17103,N_17090);
or U17241 (N_17241,N_17068,N_17178);
nand U17242 (N_17242,N_17097,N_17132);
xor U17243 (N_17243,N_17075,N_17017);
or U17244 (N_17244,N_17148,N_17004);
xor U17245 (N_17245,N_17156,N_17171);
xor U17246 (N_17246,N_17174,N_17191);
nand U17247 (N_17247,N_17034,N_17036);
or U17248 (N_17248,N_17076,N_17064);
nand U17249 (N_17249,N_17094,N_17082);
nand U17250 (N_17250,N_17182,N_17194);
and U17251 (N_17251,N_17157,N_17029);
nor U17252 (N_17252,N_17074,N_17063);
nor U17253 (N_17253,N_17088,N_17092);
nor U17254 (N_17254,N_17048,N_17144);
xnor U17255 (N_17255,N_17073,N_17166);
nor U17256 (N_17256,N_17198,N_17024);
xor U17257 (N_17257,N_17069,N_17013);
or U17258 (N_17258,N_17047,N_17137);
nor U17259 (N_17259,N_17169,N_17125);
and U17260 (N_17260,N_17193,N_17143);
or U17261 (N_17261,N_17050,N_17158);
or U17262 (N_17262,N_17120,N_17039);
xor U17263 (N_17263,N_17070,N_17035);
xnor U17264 (N_17264,N_17040,N_17065);
nand U17265 (N_17265,N_17110,N_17041);
nor U17266 (N_17266,N_17186,N_17046);
nor U17267 (N_17267,N_17014,N_17153);
nand U17268 (N_17268,N_17160,N_17106);
nor U17269 (N_17269,N_17142,N_17151);
and U17270 (N_17270,N_17025,N_17021);
nand U17271 (N_17271,N_17002,N_17119);
and U17272 (N_17272,N_17005,N_17043);
or U17273 (N_17273,N_17112,N_17084);
or U17274 (N_17274,N_17062,N_17136);
xnor U17275 (N_17275,N_17139,N_17196);
nand U17276 (N_17276,N_17051,N_17102);
nor U17277 (N_17277,N_17007,N_17161);
or U17278 (N_17278,N_17098,N_17122);
nor U17279 (N_17279,N_17054,N_17118);
nand U17280 (N_17280,N_17079,N_17128);
and U17281 (N_17281,N_17165,N_17123);
nor U17282 (N_17282,N_17086,N_17126);
or U17283 (N_17283,N_17009,N_17018);
nor U17284 (N_17284,N_17010,N_17150);
xor U17285 (N_17285,N_17105,N_17146);
and U17286 (N_17286,N_17058,N_17124);
or U17287 (N_17287,N_17037,N_17135);
and U17288 (N_17288,N_17130,N_17026);
and U17289 (N_17289,N_17003,N_17199);
or U17290 (N_17290,N_17152,N_17000);
or U17291 (N_17291,N_17185,N_17189);
or U17292 (N_17292,N_17066,N_17027);
xor U17293 (N_17293,N_17179,N_17012);
nor U17294 (N_17294,N_17117,N_17176);
nand U17295 (N_17295,N_17059,N_17109);
and U17296 (N_17296,N_17173,N_17177);
and U17297 (N_17297,N_17077,N_17052);
and U17298 (N_17298,N_17167,N_17016);
nand U17299 (N_17299,N_17111,N_17187);
xor U17300 (N_17300,N_17038,N_17102);
xor U17301 (N_17301,N_17120,N_17102);
nor U17302 (N_17302,N_17141,N_17066);
xnor U17303 (N_17303,N_17099,N_17199);
nand U17304 (N_17304,N_17135,N_17174);
xnor U17305 (N_17305,N_17162,N_17165);
or U17306 (N_17306,N_17136,N_17107);
and U17307 (N_17307,N_17133,N_17084);
or U17308 (N_17308,N_17114,N_17153);
nand U17309 (N_17309,N_17098,N_17192);
or U17310 (N_17310,N_17152,N_17116);
nor U17311 (N_17311,N_17005,N_17100);
nor U17312 (N_17312,N_17023,N_17029);
nand U17313 (N_17313,N_17058,N_17011);
nand U17314 (N_17314,N_17072,N_17049);
nor U17315 (N_17315,N_17022,N_17149);
xnor U17316 (N_17316,N_17153,N_17085);
and U17317 (N_17317,N_17069,N_17074);
or U17318 (N_17318,N_17184,N_17055);
nor U17319 (N_17319,N_17015,N_17035);
or U17320 (N_17320,N_17079,N_17084);
or U17321 (N_17321,N_17017,N_17183);
and U17322 (N_17322,N_17080,N_17179);
and U17323 (N_17323,N_17061,N_17041);
nand U17324 (N_17324,N_17129,N_17071);
or U17325 (N_17325,N_17177,N_17143);
and U17326 (N_17326,N_17077,N_17122);
nor U17327 (N_17327,N_17120,N_17041);
nor U17328 (N_17328,N_17174,N_17183);
xnor U17329 (N_17329,N_17078,N_17130);
nor U17330 (N_17330,N_17157,N_17100);
nand U17331 (N_17331,N_17190,N_17182);
xnor U17332 (N_17332,N_17043,N_17054);
xnor U17333 (N_17333,N_17118,N_17094);
and U17334 (N_17334,N_17166,N_17147);
xor U17335 (N_17335,N_17159,N_17158);
or U17336 (N_17336,N_17022,N_17165);
xor U17337 (N_17337,N_17115,N_17138);
xnor U17338 (N_17338,N_17079,N_17179);
or U17339 (N_17339,N_17013,N_17131);
xor U17340 (N_17340,N_17010,N_17157);
nand U17341 (N_17341,N_17191,N_17081);
xor U17342 (N_17342,N_17147,N_17168);
nand U17343 (N_17343,N_17043,N_17171);
or U17344 (N_17344,N_17036,N_17180);
nand U17345 (N_17345,N_17054,N_17088);
xnor U17346 (N_17346,N_17103,N_17076);
nor U17347 (N_17347,N_17149,N_17122);
nor U17348 (N_17348,N_17045,N_17134);
nand U17349 (N_17349,N_17036,N_17147);
xnor U17350 (N_17350,N_17165,N_17119);
or U17351 (N_17351,N_17031,N_17194);
xnor U17352 (N_17352,N_17128,N_17103);
or U17353 (N_17353,N_17003,N_17091);
nor U17354 (N_17354,N_17116,N_17107);
or U17355 (N_17355,N_17024,N_17177);
and U17356 (N_17356,N_17063,N_17183);
nor U17357 (N_17357,N_17169,N_17180);
and U17358 (N_17358,N_17144,N_17176);
xor U17359 (N_17359,N_17093,N_17144);
xor U17360 (N_17360,N_17018,N_17127);
and U17361 (N_17361,N_17084,N_17150);
or U17362 (N_17362,N_17081,N_17094);
and U17363 (N_17363,N_17055,N_17142);
and U17364 (N_17364,N_17135,N_17001);
nand U17365 (N_17365,N_17168,N_17150);
or U17366 (N_17366,N_17056,N_17082);
or U17367 (N_17367,N_17186,N_17198);
nor U17368 (N_17368,N_17012,N_17145);
nand U17369 (N_17369,N_17195,N_17069);
and U17370 (N_17370,N_17001,N_17167);
xor U17371 (N_17371,N_17147,N_17055);
xnor U17372 (N_17372,N_17069,N_17172);
or U17373 (N_17373,N_17195,N_17144);
xnor U17374 (N_17374,N_17150,N_17077);
and U17375 (N_17375,N_17117,N_17063);
nor U17376 (N_17376,N_17184,N_17051);
and U17377 (N_17377,N_17116,N_17002);
nor U17378 (N_17378,N_17166,N_17070);
nor U17379 (N_17379,N_17029,N_17004);
nor U17380 (N_17380,N_17157,N_17084);
xor U17381 (N_17381,N_17076,N_17119);
xnor U17382 (N_17382,N_17195,N_17028);
nand U17383 (N_17383,N_17040,N_17019);
nand U17384 (N_17384,N_17081,N_17154);
and U17385 (N_17385,N_17159,N_17163);
nand U17386 (N_17386,N_17091,N_17185);
or U17387 (N_17387,N_17183,N_17038);
nor U17388 (N_17388,N_17174,N_17111);
nand U17389 (N_17389,N_17183,N_17156);
xnor U17390 (N_17390,N_17087,N_17081);
or U17391 (N_17391,N_17137,N_17011);
nand U17392 (N_17392,N_17154,N_17018);
or U17393 (N_17393,N_17181,N_17135);
or U17394 (N_17394,N_17005,N_17196);
and U17395 (N_17395,N_17031,N_17177);
nor U17396 (N_17396,N_17001,N_17035);
or U17397 (N_17397,N_17176,N_17130);
xnor U17398 (N_17398,N_17037,N_17166);
or U17399 (N_17399,N_17126,N_17010);
and U17400 (N_17400,N_17254,N_17297);
or U17401 (N_17401,N_17304,N_17229);
and U17402 (N_17402,N_17377,N_17356);
nand U17403 (N_17403,N_17281,N_17385);
or U17404 (N_17404,N_17342,N_17364);
nand U17405 (N_17405,N_17379,N_17228);
xor U17406 (N_17406,N_17201,N_17273);
xor U17407 (N_17407,N_17352,N_17382);
nand U17408 (N_17408,N_17348,N_17373);
nor U17409 (N_17409,N_17223,N_17208);
nand U17410 (N_17410,N_17398,N_17294);
or U17411 (N_17411,N_17328,N_17245);
xor U17412 (N_17412,N_17368,N_17248);
or U17413 (N_17413,N_17291,N_17286);
or U17414 (N_17414,N_17320,N_17347);
and U17415 (N_17415,N_17299,N_17218);
nand U17416 (N_17416,N_17302,N_17202);
nor U17417 (N_17417,N_17258,N_17307);
and U17418 (N_17418,N_17311,N_17203);
and U17419 (N_17419,N_17261,N_17361);
or U17420 (N_17420,N_17345,N_17386);
nor U17421 (N_17421,N_17390,N_17334);
and U17422 (N_17422,N_17381,N_17240);
xor U17423 (N_17423,N_17253,N_17214);
or U17424 (N_17424,N_17354,N_17296);
and U17425 (N_17425,N_17272,N_17392);
and U17426 (N_17426,N_17389,N_17359);
nand U17427 (N_17427,N_17251,N_17293);
or U17428 (N_17428,N_17282,N_17301);
xor U17429 (N_17429,N_17244,N_17225);
nor U17430 (N_17430,N_17204,N_17220);
or U17431 (N_17431,N_17306,N_17232);
nand U17432 (N_17432,N_17351,N_17310);
xnor U17433 (N_17433,N_17265,N_17399);
xor U17434 (N_17434,N_17367,N_17316);
nand U17435 (N_17435,N_17274,N_17243);
xnor U17436 (N_17436,N_17239,N_17262);
nor U17437 (N_17437,N_17215,N_17329);
or U17438 (N_17438,N_17231,N_17234);
and U17439 (N_17439,N_17312,N_17211);
nand U17440 (N_17440,N_17380,N_17308);
and U17441 (N_17441,N_17255,N_17270);
and U17442 (N_17442,N_17300,N_17370);
and U17443 (N_17443,N_17263,N_17357);
and U17444 (N_17444,N_17363,N_17339);
or U17445 (N_17445,N_17349,N_17384);
and U17446 (N_17446,N_17396,N_17327);
xor U17447 (N_17447,N_17287,N_17383);
and U17448 (N_17448,N_17219,N_17366);
xnor U17449 (N_17449,N_17242,N_17246);
and U17450 (N_17450,N_17205,N_17346);
or U17451 (N_17451,N_17280,N_17252);
nand U17452 (N_17452,N_17317,N_17212);
xor U17453 (N_17453,N_17341,N_17315);
nor U17454 (N_17454,N_17227,N_17319);
or U17455 (N_17455,N_17372,N_17290);
nand U17456 (N_17456,N_17314,N_17309);
or U17457 (N_17457,N_17295,N_17344);
and U17458 (N_17458,N_17230,N_17237);
nor U17459 (N_17459,N_17369,N_17335);
or U17460 (N_17460,N_17285,N_17371);
xnor U17461 (N_17461,N_17292,N_17200);
nor U17462 (N_17462,N_17325,N_17397);
and U17463 (N_17463,N_17353,N_17387);
or U17464 (N_17464,N_17217,N_17360);
or U17465 (N_17465,N_17283,N_17330);
nand U17466 (N_17466,N_17362,N_17276);
nor U17467 (N_17467,N_17350,N_17206);
nand U17468 (N_17468,N_17391,N_17303);
and U17469 (N_17469,N_17222,N_17264);
xor U17470 (N_17470,N_17375,N_17257);
or U17471 (N_17471,N_17298,N_17388);
and U17472 (N_17472,N_17331,N_17332);
nand U17473 (N_17473,N_17241,N_17247);
xnor U17474 (N_17474,N_17250,N_17365);
nor U17475 (N_17475,N_17233,N_17322);
or U17476 (N_17476,N_17324,N_17338);
nor U17477 (N_17477,N_17224,N_17321);
xnor U17478 (N_17478,N_17323,N_17213);
and U17479 (N_17479,N_17221,N_17216);
or U17480 (N_17480,N_17336,N_17340);
or U17481 (N_17481,N_17378,N_17266);
or U17482 (N_17482,N_17355,N_17337);
or U17483 (N_17483,N_17209,N_17260);
nor U17484 (N_17484,N_17267,N_17288);
or U17485 (N_17485,N_17275,N_17374);
or U17486 (N_17486,N_17279,N_17393);
and U17487 (N_17487,N_17238,N_17259);
and U17488 (N_17488,N_17277,N_17249);
xnor U17489 (N_17489,N_17333,N_17395);
nor U17490 (N_17490,N_17318,N_17271);
or U17491 (N_17491,N_17326,N_17278);
xor U17492 (N_17492,N_17207,N_17394);
nand U17493 (N_17493,N_17289,N_17236);
and U17494 (N_17494,N_17226,N_17358);
xnor U17495 (N_17495,N_17376,N_17343);
and U17496 (N_17496,N_17268,N_17269);
nor U17497 (N_17497,N_17256,N_17210);
nand U17498 (N_17498,N_17313,N_17305);
nor U17499 (N_17499,N_17284,N_17235);
and U17500 (N_17500,N_17300,N_17266);
nor U17501 (N_17501,N_17314,N_17365);
and U17502 (N_17502,N_17213,N_17283);
nand U17503 (N_17503,N_17275,N_17387);
xnor U17504 (N_17504,N_17394,N_17288);
xor U17505 (N_17505,N_17225,N_17216);
xor U17506 (N_17506,N_17299,N_17209);
nor U17507 (N_17507,N_17273,N_17319);
and U17508 (N_17508,N_17222,N_17230);
xnor U17509 (N_17509,N_17391,N_17234);
nor U17510 (N_17510,N_17332,N_17317);
nor U17511 (N_17511,N_17398,N_17274);
nor U17512 (N_17512,N_17385,N_17302);
nor U17513 (N_17513,N_17215,N_17229);
nor U17514 (N_17514,N_17370,N_17251);
nand U17515 (N_17515,N_17266,N_17386);
xor U17516 (N_17516,N_17380,N_17367);
nand U17517 (N_17517,N_17281,N_17246);
or U17518 (N_17518,N_17229,N_17383);
or U17519 (N_17519,N_17348,N_17293);
nand U17520 (N_17520,N_17317,N_17263);
nor U17521 (N_17521,N_17360,N_17246);
nand U17522 (N_17522,N_17260,N_17311);
nand U17523 (N_17523,N_17232,N_17260);
or U17524 (N_17524,N_17235,N_17344);
and U17525 (N_17525,N_17306,N_17202);
or U17526 (N_17526,N_17296,N_17235);
nor U17527 (N_17527,N_17240,N_17228);
nand U17528 (N_17528,N_17353,N_17256);
and U17529 (N_17529,N_17307,N_17212);
nor U17530 (N_17530,N_17369,N_17366);
or U17531 (N_17531,N_17258,N_17354);
xor U17532 (N_17532,N_17368,N_17319);
xor U17533 (N_17533,N_17324,N_17391);
nor U17534 (N_17534,N_17255,N_17226);
nand U17535 (N_17535,N_17212,N_17235);
nor U17536 (N_17536,N_17218,N_17327);
nor U17537 (N_17537,N_17391,N_17237);
nor U17538 (N_17538,N_17282,N_17290);
xnor U17539 (N_17539,N_17318,N_17397);
or U17540 (N_17540,N_17290,N_17376);
or U17541 (N_17541,N_17356,N_17333);
nor U17542 (N_17542,N_17285,N_17211);
xnor U17543 (N_17543,N_17270,N_17364);
or U17544 (N_17544,N_17367,N_17217);
nand U17545 (N_17545,N_17212,N_17357);
and U17546 (N_17546,N_17303,N_17379);
xor U17547 (N_17547,N_17203,N_17294);
nand U17548 (N_17548,N_17246,N_17268);
nand U17549 (N_17549,N_17234,N_17210);
xnor U17550 (N_17550,N_17354,N_17373);
and U17551 (N_17551,N_17257,N_17210);
xor U17552 (N_17552,N_17391,N_17366);
and U17553 (N_17553,N_17379,N_17336);
nor U17554 (N_17554,N_17270,N_17361);
xor U17555 (N_17555,N_17247,N_17316);
nand U17556 (N_17556,N_17388,N_17224);
or U17557 (N_17557,N_17312,N_17304);
xor U17558 (N_17558,N_17364,N_17244);
nor U17559 (N_17559,N_17207,N_17282);
xnor U17560 (N_17560,N_17282,N_17305);
nand U17561 (N_17561,N_17375,N_17320);
xnor U17562 (N_17562,N_17305,N_17286);
or U17563 (N_17563,N_17239,N_17381);
nand U17564 (N_17564,N_17325,N_17250);
nand U17565 (N_17565,N_17237,N_17334);
nand U17566 (N_17566,N_17316,N_17243);
nand U17567 (N_17567,N_17382,N_17346);
or U17568 (N_17568,N_17322,N_17251);
xnor U17569 (N_17569,N_17200,N_17368);
and U17570 (N_17570,N_17295,N_17359);
and U17571 (N_17571,N_17207,N_17244);
or U17572 (N_17572,N_17257,N_17307);
nor U17573 (N_17573,N_17385,N_17322);
or U17574 (N_17574,N_17230,N_17207);
xnor U17575 (N_17575,N_17263,N_17383);
nor U17576 (N_17576,N_17242,N_17257);
nand U17577 (N_17577,N_17330,N_17319);
nor U17578 (N_17578,N_17266,N_17363);
and U17579 (N_17579,N_17372,N_17260);
or U17580 (N_17580,N_17227,N_17235);
and U17581 (N_17581,N_17311,N_17392);
xnor U17582 (N_17582,N_17266,N_17332);
xnor U17583 (N_17583,N_17392,N_17377);
nand U17584 (N_17584,N_17351,N_17242);
nor U17585 (N_17585,N_17370,N_17335);
nor U17586 (N_17586,N_17220,N_17214);
or U17587 (N_17587,N_17377,N_17358);
xor U17588 (N_17588,N_17348,N_17388);
xor U17589 (N_17589,N_17267,N_17255);
nor U17590 (N_17590,N_17287,N_17307);
nand U17591 (N_17591,N_17201,N_17368);
or U17592 (N_17592,N_17201,N_17219);
xnor U17593 (N_17593,N_17208,N_17284);
xnor U17594 (N_17594,N_17383,N_17322);
nor U17595 (N_17595,N_17227,N_17307);
and U17596 (N_17596,N_17233,N_17296);
and U17597 (N_17597,N_17228,N_17285);
nor U17598 (N_17598,N_17234,N_17372);
nand U17599 (N_17599,N_17388,N_17331);
nor U17600 (N_17600,N_17491,N_17507);
or U17601 (N_17601,N_17458,N_17505);
xor U17602 (N_17602,N_17504,N_17476);
and U17603 (N_17603,N_17435,N_17574);
xor U17604 (N_17604,N_17542,N_17596);
and U17605 (N_17605,N_17463,N_17443);
or U17606 (N_17606,N_17418,N_17599);
or U17607 (N_17607,N_17469,N_17433);
or U17608 (N_17608,N_17481,N_17534);
or U17609 (N_17609,N_17556,N_17401);
or U17610 (N_17610,N_17506,N_17410);
xnor U17611 (N_17611,N_17594,N_17529);
and U17612 (N_17612,N_17412,N_17595);
or U17613 (N_17613,N_17495,N_17598);
or U17614 (N_17614,N_17503,N_17572);
nand U17615 (N_17615,N_17456,N_17497);
nor U17616 (N_17616,N_17436,N_17462);
xor U17617 (N_17617,N_17553,N_17409);
xor U17618 (N_17618,N_17400,N_17512);
or U17619 (N_17619,N_17474,N_17588);
and U17620 (N_17620,N_17597,N_17516);
and U17621 (N_17621,N_17550,N_17475);
or U17622 (N_17622,N_17533,N_17459);
and U17623 (N_17623,N_17508,N_17416);
and U17624 (N_17624,N_17407,N_17521);
nand U17625 (N_17625,N_17515,N_17483);
nand U17626 (N_17626,N_17546,N_17403);
or U17627 (N_17627,N_17423,N_17540);
or U17628 (N_17628,N_17580,N_17451);
or U17629 (N_17629,N_17582,N_17581);
and U17630 (N_17630,N_17501,N_17405);
nand U17631 (N_17631,N_17496,N_17535);
nor U17632 (N_17632,N_17419,N_17492);
and U17633 (N_17633,N_17532,N_17593);
or U17634 (N_17634,N_17537,N_17525);
nor U17635 (N_17635,N_17570,N_17452);
or U17636 (N_17636,N_17518,N_17558);
or U17637 (N_17637,N_17590,N_17488);
or U17638 (N_17638,N_17404,N_17592);
or U17639 (N_17639,N_17408,N_17520);
or U17640 (N_17640,N_17519,N_17438);
or U17641 (N_17641,N_17539,N_17531);
xor U17642 (N_17642,N_17464,N_17559);
and U17643 (N_17643,N_17552,N_17490);
xor U17644 (N_17644,N_17579,N_17447);
xnor U17645 (N_17645,N_17484,N_17541);
and U17646 (N_17646,N_17437,N_17494);
or U17647 (N_17647,N_17528,N_17426);
xor U17648 (N_17648,N_17575,N_17493);
or U17649 (N_17649,N_17479,N_17568);
and U17650 (N_17650,N_17414,N_17444);
and U17651 (N_17651,N_17563,N_17536);
nor U17652 (N_17652,N_17467,N_17465);
and U17653 (N_17653,N_17545,N_17578);
and U17654 (N_17654,N_17470,N_17487);
nand U17655 (N_17655,N_17522,N_17560);
or U17656 (N_17656,N_17468,N_17513);
nand U17657 (N_17657,N_17448,N_17565);
xor U17658 (N_17658,N_17544,N_17530);
nor U17659 (N_17659,N_17573,N_17586);
nor U17660 (N_17660,N_17510,N_17526);
xnor U17661 (N_17661,N_17538,N_17432);
or U17662 (N_17662,N_17431,N_17486);
or U17663 (N_17663,N_17472,N_17454);
and U17664 (N_17664,N_17461,N_17449);
or U17665 (N_17665,N_17427,N_17523);
or U17666 (N_17666,N_17569,N_17477);
nor U17667 (N_17667,N_17554,N_17499);
nor U17668 (N_17668,N_17425,N_17441);
nand U17669 (N_17669,N_17548,N_17584);
and U17670 (N_17670,N_17567,N_17406);
nor U17671 (N_17671,N_17457,N_17413);
and U17672 (N_17672,N_17561,N_17524);
xor U17673 (N_17673,N_17428,N_17402);
nor U17674 (N_17674,N_17411,N_17439);
xnor U17675 (N_17675,N_17446,N_17466);
nand U17676 (N_17676,N_17473,N_17589);
and U17677 (N_17677,N_17571,N_17450);
nor U17678 (N_17678,N_17514,N_17562);
or U17679 (N_17679,N_17442,N_17547);
or U17680 (N_17680,N_17424,N_17583);
nor U17681 (N_17681,N_17555,N_17471);
nor U17682 (N_17682,N_17440,N_17564);
xnor U17683 (N_17683,N_17453,N_17551);
and U17684 (N_17684,N_17422,N_17577);
and U17685 (N_17685,N_17417,N_17576);
and U17686 (N_17686,N_17543,N_17485);
xor U17687 (N_17687,N_17527,N_17415);
nor U17688 (N_17688,N_17585,N_17480);
nor U17689 (N_17689,N_17498,N_17429);
or U17690 (N_17690,N_17502,N_17500);
and U17691 (N_17691,N_17455,N_17566);
xnor U17692 (N_17692,N_17421,N_17434);
nor U17693 (N_17693,N_17549,N_17557);
nor U17694 (N_17694,N_17509,N_17478);
nor U17695 (N_17695,N_17587,N_17511);
nor U17696 (N_17696,N_17482,N_17460);
or U17697 (N_17697,N_17591,N_17517);
or U17698 (N_17698,N_17420,N_17445);
or U17699 (N_17699,N_17430,N_17489);
and U17700 (N_17700,N_17479,N_17545);
xor U17701 (N_17701,N_17553,N_17506);
or U17702 (N_17702,N_17418,N_17554);
and U17703 (N_17703,N_17531,N_17586);
or U17704 (N_17704,N_17411,N_17579);
nand U17705 (N_17705,N_17534,N_17515);
nor U17706 (N_17706,N_17440,N_17437);
and U17707 (N_17707,N_17443,N_17489);
xor U17708 (N_17708,N_17570,N_17519);
xnor U17709 (N_17709,N_17556,N_17484);
or U17710 (N_17710,N_17498,N_17537);
nor U17711 (N_17711,N_17496,N_17443);
xor U17712 (N_17712,N_17529,N_17491);
or U17713 (N_17713,N_17598,N_17503);
nor U17714 (N_17714,N_17549,N_17432);
nand U17715 (N_17715,N_17580,N_17574);
or U17716 (N_17716,N_17495,N_17568);
nor U17717 (N_17717,N_17539,N_17579);
nand U17718 (N_17718,N_17558,N_17476);
nand U17719 (N_17719,N_17507,N_17560);
and U17720 (N_17720,N_17576,N_17477);
nand U17721 (N_17721,N_17429,N_17591);
nand U17722 (N_17722,N_17595,N_17592);
xnor U17723 (N_17723,N_17493,N_17450);
xor U17724 (N_17724,N_17531,N_17460);
nor U17725 (N_17725,N_17548,N_17420);
and U17726 (N_17726,N_17416,N_17527);
xnor U17727 (N_17727,N_17542,N_17518);
nand U17728 (N_17728,N_17519,N_17425);
nor U17729 (N_17729,N_17578,N_17512);
xor U17730 (N_17730,N_17598,N_17467);
xnor U17731 (N_17731,N_17471,N_17532);
nor U17732 (N_17732,N_17502,N_17417);
nand U17733 (N_17733,N_17498,N_17478);
nor U17734 (N_17734,N_17565,N_17520);
nand U17735 (N_17735,N_17405,N_17473);
nand U17736 (N_17736,N_17445,N_17408);
xor U17737 (N_17737,N_17511,N_17466);
nand U17738 (N_17738,N_17525,N_17583);
and U17739 (N_17739,N_17510,N_17408);
nor U17740 (N_17740,N_17423,N_17456);
nor U17741 (N_17741,N_17402,N_17484);
xor U17742 (N_17742,N_17451,N_17582);
nand U17743 (N_17743,N_17467,N_17575);
and U17744 (N_17744,N_17512,N_17533);
and U17745 (N_17745,N_17516,N_17509);
nor U17746 (N_17746,N_17562,N_17487);
and U17747 (N_17747,N_17530,N_17532);
and U17748 (N_17748,N_17538,N_17492);
nand U17749 (N_17749,N_17548,N_17529);
xor U17750 (N_17750,N_17588,N_17468);
xor U17751 (N_17751,N_17581,N_17415);
xor U17752 (N_17752,N_17498,N_17475);
and U17753 (N_17753,N_17501,N_17531);
or U17754 (N_17754,N_17562,N_17473);
nand U17755 (N_17755,N_17501,N_17585);
and U17756 (N_17756,N_17414,N_17498);
and U17757 (N_17757,N_17499,N_17454);
nor U17758 (N_17758,N_17562,N_17504);
or U17759 (N_17759,N_17424,N_17539);
or U17760 (N_17760,N_17505,N_17592);
xor U17761 (N_17761,N_17522,N_17448);
xnor U17762 (N_17762,N_17560,N_17480);
xnor U17763 (N_17763,N_17567,N_17582);
nor U17764 (N_17764,N_17510,N_17598);
nand U17765 (N_17765,N_17457,N_17445);
xor U17766 (N_17766,N_17501,N_17572);
nand U17767 (N_17767,N_17421,N_17562);
and U17768 (N_17768,N_17565,N_17500);
or U17769 (N_17769,N_17533,N_17442);
nor U17770 (N_17770,N_17409,N_17415);
and U17771 (N_17771,N_17448,N_17575);
xnor U17772 (N_17772,N_17558,N_17507);
xor U17773 (N_17773,N_17441,N_17401);
xor U17774 (N_17774,N_17434,N_17430);
nor U17775 (N_17775,N_17473,N_17438);
nor U17776 (N_17776,N_17416,N_17511);
xnor U17777 (N_17777,N_17440,N_17490);
nor U17778 (N_17778,N_17448,N_17524);
xor U17779 (N_17779,N_17541,N_17495);
and U17780 (N_17780,N_17441,N_17475);
nand U17781 (N_17781,N_17445,N_17527);
and U17782 (N_17782,N_17555,N_17430);
nor U17783 (N_17783,N_17449,N_17448);
xnor U17784 (N_17784,N_17459,N_17433);
xnor U17785 (N_17785,N_17484,N_17406);
xnor U17786 (N_17786,N_17437,N_17589);
or U17787 (N_17787,N_17415,N_17556);
nand U17788 (N_17788,N_17512,N_17513);
nor U17789 (N_17789,N_17503,N_17511);
nor U17790 (N_17790,N_17440,N_17581);
or U17791 (N_17791,N_17429,N_17496);
or U17792 (N_17792,N_17414,N_17458);
xnor U17793 (N_17793,N_17598,N_17589);
or U17794 (N_17794,N_17483,N_17531);
nand U17795 (N_17795,N_17417,N_17572);
xnor U17796 (N_17796,N_17478,N_17555);
nor U17797 (N_17797,N_17565,N_17599);
and U17798 (N_17798,N_17550,N_17507);
nor U17799 (N_17799,N_17594,N_17560);
xnor U17800 (N_17800,N_17725,N_17648);
nand U17801 (N_17801,N_17647,N_17697);
nand U17802 (N_17802,N_17709,N_17679);
and U17803 (N_17803,N_17727,N_17636);
nor U17804 (N_17804,N_17701,N_17649);
nand U17805 (N_17805,N_17635,N_17688);
xnor U17806 (N_17806,N_17626,N_17617);
or U17807 (N_17807,N_17750,N_17706);
or U17808 (N_17808,N_17668,N_17759);
or U17809 (N_17809,N_17621,N_17673);
or U17810 (N_17810,N_17777,N_17631);
and U17811 (N_17811,N_17717,N_17629);
nor U17812 (N_17812,N_17784,N_17646);
and U17813 (N_17813,N_17684,N_17654);
and U17814 (N_17814,N_17793,N_17796);
nor U17815 (N_17815,N_17756,N_17786);
xnor U17816 (N_17816,N_17734,N_17704);
and U17817 (N_17817,N_17669,N_17686);
xnor U17818 (N_17818,N_17656,N_17715);
or U17819 (N_17819,N_17644,N_17719);
and U17820 (N_17820,N_17702,N_17741);
nand U17821 (N_17821,N_17724,N_17768);
nor U17822 (N_17822,N_17752,N_17735);
nor U17823 (N_17823,N_17770,N_17781);
xnor U17824 (N_17824,N_17634,N_17795);
and U17825 (N_17825,N_17604,N_17671);
and U17826 (N_17826,N_17609,N_17678);
nor U17827 (N_17827,N_17682,N_17699);
nor U17828 (N_17828,N_17675,N_17651);
nand U17829 (N_17829,N_17757,N_17645);
xor U17830 (N_17830,N_17751,N_17600);
nand U17831 (N_17831,N_17794,N_17625);
xor U17832 (N_17832,N_17790,N_17791);
nor U17833 (N_17833,N_17722,N_17742);
and U17834 (N_17834,N_17611,N_17639);
nand U17835 (N_17835,N_17762,N_17713);
nor U17836 (N_17836,N_17758,N_17774);
and U17837 (N_17837,N_17681,N_17707);
or U17838 (N_17838,N_17653,N_17664);
or U17839 (N_17839,N_17642,N_17710);
nor U17840 (N_17840,N_17665,N_17663);
xor U17841 (N_17841,N_17680,N_17705);
or U17842 (N_17842,N_17737,N_17780);
xnor U17843 (N_17843,N_17789,N_17782);
or U17844 (N_17844,N_17732,N_17615);
xnor U17845 (N_17845,N_17743,N_17728);
and U17846 (N_17846,N_17687,N_17637);
or U17847 (N_17847,N_17661,N_17603);
and U17848 (N_17848,N_17667,N_17783);
or U17849 (N_17849,N_17754,N_17712);
nor U17850 (N_17850,N_17753,N_17624);
nor U17851 (N_17851,N_17767,N_17623);
and U17852 (N_17852,N_17630,N_17622);
nor U17853 (N_17853,N_17788,N_17776);
xnor U17854 (N_17854,N_17726,N_17723);
or U17855 (N_17855,N_17677,N_17674);
or U17856 (N_17856,N_17766,N_17708);
xor U17857 (N_17857,N_17763,N_17655);
xor U17858 (N_17858,N_17659,N_17749);
or U17859 (N_17859,N_17694,N_17605);
nand U17860 (N_17860,N_17628,N_17672);
nor U17861 (N_17861,N_17778,N_17711);
and U17862 (N_17862,N_17755,N_17606);
nand U17863 (N_17863,N_17658,N_17736);
or U17864 (N_17864,N_17792,N_17641);
and U17865 (N_17865,N_17703,N_17612);
nor U17866 (N_17866,N_17761,N_17733);
nor U17867 (N_17867,N_17714,N_17695);
nand U17868 (N_17868,N_17633,N_17608);
nand U17869 (N_17869,N_17607,N_17798);
xnor U17870 (N_17870,N_17640,N_17632);
and U17871 (N_17871,N_17721,N_17650);
nand U17872 (N_17872,N_17772,N_17657);
and U17873 (N_17873,N_17773,N_17619);
nor U17874 (N_17874,N_17739,N_17685);
or U17875 (N_17875,N_17620,N_17720);
or U17876 (N_17876,N_17618,N_17785);
nand U17877 (N_17877,N_17696,N_17693);
nor U17878 (N_17878,N_17601,N_17775);
xnor U17879 (N_17879,N_17689,N_17799);
or U17880 (N_17880,N_17716,N_17691);
or U17881 (N_17881,N_17692,N_17731);
or U17882 (N_17882,N_17676,N_17771);
nor U17883 (N_17883,N_17797,N_17616);
xor U17884 (N_17884,N_17760,N_17660);
nand U17885 (N_17885,N_17602,N_17718);
or U17886 (N_17886,N_17745,N_17683);
nor U17887 (N_17887,N_17764,N_17613);
nor U17888 (N_17888,N_17666,N_17698);
xor U17889 (N_17889,N_17747,N_17730);
nand U17890 (N_17890,N_17740,N_17638);
and U17891 (N_17891,N_17738,N_17690);
and U17892 (N_17892,N_17700,N_17610);
nand U17893 (N_17893,N_17662,N_17670);
xnor U17894 (N_17894,N_17652,N_17779);
nor U17895 (N_17895,N_17746,N_17729);
nor U17896 (N_17896,N_17744,N_17643);
xor U17897 (N_17897,N_17627,N_17748);
xnor U17898 (N_17898,N_17769,N_17614);
or U17899 (N_17899,N_17787,N_17765);
and U17900 (N_17900,N_17720,N_17765);
nor U17901 (N_17901,N_17710,N_17773);
xor U17902 (N_17902,N_17772,N_17669);
nor U17903 (N_17903,N_17681,N_17688);
nand U17904 (N_17904,N_17644,N_17624);
nand U17905 (N_17905,N_17788,N_17721);
nand U17906 (N_17906,N_17784,N_17749);
xnor U17907 (N_17907,N_17765,N_17795);
xnor U17908 (N_17908,N_17670,N_17764);
nand U17909 (N_17909,N_17769,N_17668);
and U17910 (N_17910,N_17719,N_17729);
or U17911 (N_17911,N_17739,N_17635);
and U17912 (N_17912,N_17661,N_17681);
xor U17913 (N_17913,N_17662,N_17700);
nor U17914 (N_17914,N_17733,N_17726);
and U17915 (N_17915,N_17793,N_17699);
nand U17916 (N_17916,N_17659,N_17612);
or U17917 (N_17917,N_17639,N_17647);
xnor U17918 (N_17918,N_17616,N_17741);
and U17919 (N_17919,N_17603,N_17674);
and U17920 (N_17920,N_17739,N_17772);
nor U17921 (N_17921,N_17749,N_17798);
and U17922 (N_17922,N_17662,N_17787);
nor U17923 (N_17923,N_17616,N_17707);
or U17924 (N_17924,N_17664,N_17668);
and U17925 (N_17925,N_17759,N_17777);
or U17926 (N_17926,N_17721,N_17656);
nand U17927 (N_17927,N_17692,N_17604);
or U17928 (N_17928,N_17784,N_17619);
or U17929 (N_17929,N_17648,N_17695);
xnor U17930 (N_17930,N_17665,N_17714);
nor U17931 (N_17931,N_17678,N_17684);
nand U17932 (N_17932,N_17665,N_17609);
nand U17933 (N_17933,N_17635,N_17624);
nor U17934 (N_17934,N_17746,N_17685);
nand U17935 (N_17935,N_17654,N_17758);
xor U17936 (N_17936,N_17760,N_17651);
and U17937 (N_17937,N_17715,N_17601);
and U17938 (N_17938,N_17676,N_17729);
xnor U17939 (N_17939,N_17631,N_17701);
nand U17940 (N_17940,N_17609,N_17656);
nor U17941 (N_17941,N_17601,N_17646);
nand U17942 (N_17942,N_17770,N_17658);
and U17943 (N_17943,N_17780,N_17759);
and U17944 (N_17944,N_17665,N_17657);
xnor U17945 (N_17945,N_17689,N_17610);
and U17946 (N_17946,N_17697,N_17666);
and U17947 (N_17947,N_17633,N_17604);
nor U17948 (N_17948,N_17783,N_17636);
xor U17949 (N_17949,N_17610,N_17785);
nor U17950 (N_17950,N_17716,N_17601);
xnor U17951 (N_17951,N_17612,N_17733);
and U17952 (N_17952,N_17636,N_17632);
xnor U17953 (N_17953,N_17658,N_17799);
or U17954 (N_17954,N_17731,N_17728);
xor U17955 (N_17955,N_17705,N_17729);
or U17956 (N_17956,N_17729,N_17762);
nand U17957 (N_17957,N_17769,N_17645);
or U17958 (N_17958,N_17735,N_17723);
nand U17959 (N_17959,N_17629,N_17707);
and U17960 (N_17960,N_17623,N_17666);
xnor U17961 (N_17961,N_17783,N_17677);
nand U17962 (N_17962,N_17781,N_17661);
or U17963 (N_17963,N_17769,N_17758);
xnor U17964 (N_17964,N_17681,N_17687);
and U17965 (N_17965,N_17680,N_17685);
nand U17966 (N_17966,N_17762,N_17707);
xnor U17967 (N_17967,N_17738,N_17656);
and U17968 (N_17968,N_17659,N_17671);
nor U17969 (N_17969,N_17717,N_17680);
and U17970 (N_17970,N_17670,N_17767);
and U17971 (N_17971,N_17712,N_17671);
xnor U17972 (N_17972,N_17714,N_17774);
xnor U17973 (N_17973,N_17778,N_17603);
or U17974 (N_17974,N_17749,N_17631);
or U17975 (N_17975,N_17790,N_17680);
or U17976 (N_17976,N_17612,N_17623);
nor U17977 (N_17977,N_17741,N_17626);
xor U17978 (N_17978,N_17616,N_17605);
or U17979 (N_17979,N_17711,N_17793);
xnor U17980 (N_17980,N_17683,N_17680);
or U17981 (N_17981,N_17781,N_17678);
and U17982 (N_17982,N_17753,N_17745);
and U17983 (N_17983,N_17687,N_17759);
and U17984 (N_17984,N_17789,N_17719);
and U17985 (N_17985,N_17679,N_17772);
xnor U17986 (N_17986,N_17714,N_17789);
nor U17987 (N_17987,N_17651,N_17736);
nand U17988 (N_17988,N_17691,N_17710);
nor U17989 (N_17989,N_17763,N_17642);
nor U17990 (N_17990,N_17741,N_17645);
nand U17991 (N_17991,N_17784,N_17641);
nor U17992 (N_17992,N_17660,N_17606);
and U17993 (N_17993,N_17750,N_17658);
xnor U17994 (N_17994,N_17622,N_17600);
or U17995 (N_17995,N_17620,N_17797);
nand U17996 (N_17996,N_17619,N_17662);
and U17997 (N_17997,N_17653,N_17642);
and U17998 (N_17998,N_17760,N_17677);
or U17999 (N_17999,N_17638,N_17762);
nor U18000 (N_18000,N_17826,N_17965);
nor U18001 (N_18001,N_17929,N_17926);
nor U18002 (N_18002,N_17988,N_17879);
or U18003 (N_18003,N_17905,N_17847);
and U18004 (N_18004,N_17995,N_17954);
nor U18005 (N_18005,N_17890,N_17928);
or U18006 (N_18006,N_17915,N_17886);
or U18007 (N_18007,N_17942,N_17855);
nor U18008 (N_18008,N_17863,N_17891);
or U18009 (N_18009,N_17958,N_17922);
nand U18010 (N_18010,N_17974,N_17964);
nand U18011 (N_18011,N_17851,N_17979);
or U18012 (N_18012,N_17978,N_17893);
and U18013 (N_18013,N_17875,N_17892);
nor U18014 (N_18014,N_17802,N_17931);
or U18015 (N_18015,N_17808,N_17940);
or U18016 (N_18016,N_17852,N_17814);
and U18017 (N_18017,N_17921,N_17920);
and U18018 (N_18018,N_17866,N_17956);
and U18019 (N_18019,N_17946,N_17980);
or U18020 (N_18020,N_17914,N_17927);
nand U18021 (N_18021,N_17837,N_17945);
nor U18022 (N_18022,N_17960,N_17824);
nand U18023 (N_18023,N_17831,N_17815);
nor U18024 (N_18024,N_17903,N_17962);
and U18025 (N_18025,N_17898,N_17884);
nand U18026 (N_18026,N_17934,N_17801);
or U18027 (N_18027,N_17846,N_17818);
nand U18028 (N_18028,N_17849,N_17806);
nor U18029 (N_18029,N_17901,N_17805);
nor U18030 (N_18030,N_17895,N_17829);
xor U18031 (N_18031,N_17944,N_17984);
nand U18032 (N_18032,N_17843,N_17850);
and U18033 (N_18033,N_17904,N_17845);
nor U18034 (N_18034,N_17870,N_17957);
or U18035 (N_18035,N_17813,N_17830);
or U18036 (N_18036,N_17894,N_17867);
and U18037 (N_18037,N_17912,N_17918);
and U18038 (N_18038,N_17857,N_17888);
xor U18039 (N_18039,N_17865,N_17937);
nor U18040 (N_18040,N_17932,N_17985);
or U18041 (N_18041,N_17935,N_17878);
or U18042 (N_18042,N_17933,N_17963);
or U18043 (N_18043,N_17812,N_17938);
nand U18044 (N_18044,N_17976,N_17874);
or U18045 (N_18045,N_17916,N_17924);
xor U18046 (N_18046,N_17816,N_17968);
nand U18047 (N_18047,N_17919,N_17835);
or U18048 (N_18048,N_17950,N_17839);
xnor U18049 (N_18049,N_17883,N_17871);
nand U18050 (N_18050,N_17907,N_17911);
nor U18051 (N_18051,N_17993,N_17949);
xnor U18052 (N_18052,N_17820,N_17811);
nor U18053 (N_18053,N_17882,N_17951);
nand U18054 (N_18054,N_17889,N_17943);
or U18055 (N_18055,N_17864,N_17840);
nor U18056 (N_18056,N_17969,N_17860);
or U18057 (N_18057,N_17971,N_17827);
or U18058 (N_18058,N_17982,N_17999);
xor U18059 (N_18059,N_17981,N_17841);
and U18060 (N_18060,N_17947,N_17910);
nand U18061 (N_18061,N_17909,N_17885);
and U18062 (N_18062,N_17997,N_17939);
nor U18063 (N_18063,N_17856,N_17868);
nor U18064 (N_18064,N_17804,N_17819);
nand U18065 (N_18065,N_17897,N_17832);
nand U18066 (N_18066,N_17822,N_17880);
nor U18067 (N_18067,N_17930,N_17809);
or U18068 (N_18068,N_17821,N_17994);
nand U18069 (N_18069,N_17967,N_17817);
nand U18070 (N_18070,N_17998,N_17836);
nor U18071 (N_18071,N_17800,N_17952);
nand U18072 (N_18072,N_17970,N_17803);
nand U18073 (N_18073,N_17906,N_17872);
nor U18074 (N_18074,N_17858,N_17877);
nand U18075 (N_18075,N_17810,N_17989);
or U18076 (N_18076,N_17854,N_17842);
nor U18077 (N_18077,N_17896,N_17869);
or U18078 (N_18078,N_17996,N_17936);
or U18079 (N_18079,N_17948,N_17983);
or U18080 (N_18080,N_17991,N_17955);
nor U18081 (N_18081,N_17834,N_17838);
xnor U18082 (N_18082,N_17961,N_17992);
or U18083 (N_18083,N_17925,N_17913);
xnor U18084 (N_18084,N_17923,N_17844);
nor U18085 (N_18085,N_17859,N_17902);
or U18086 (N_18086,N_17807,N_17861);
nand U18087 (N_18087,N_17873,N_17917);
nor U18088 (N_18088,N_17941,N_17848);
nand U18089 (N_18089,N_17887,N_17975);
and U18090 (N_18090,N_17853,N_17959);
xor U18091 (N_18091,N_17828,N_17972);
nor U18092 (N_18092,N_17881,N_17987);
nand U18093 (N_18093,N_17862,N_17973);
or U18094 (N_18094,N_17977,N_17823);
xnor U18095 (N_18095,N_17833,N_17966);
or U18096 (N_18096,N_17986,N_17908);
and U18097 (N_18097,N_17900,N_17990);
xnor U18098 (N_18098,N_17876,N_17899);
and U18099 (N_18099,N_17953,N_17825);
or U18100 (N_18100,N_17919,N_17851);
nand U18101 (N_18101,N_17996,N_17879);
xnor U18102 (N_18102,N_17810,N_17832);
nand U18103 (N_18103,N_17999,N_17903);
nor U18104 (N_18104,N_17978,N_17983);
nor U18105 (N_18105,N_17957,N_17864);
or U18106 (N_18106,N_17876,N_17930);
and U18107 (N_18107,N_17996,N_17883);
nor U18108 (N_18108,N_17938,N_17845);
or U18109 (N_18109,N_17821,N_17939);
xnor U18110 (N_18110,N_17967,N_17897);
and U18111 (N_18111,N_17983,N_17995);
and U18112 (N_18112,N_17865,N_17927);
xor U18113 (N_18113,N_17898,N_17926);
nor U18114 (N_18114,N_17821,N_17930);
xor U18115 (N_18115,N_17958,N_17819);
xor U18116 (N_18116,N_17804,N_17861);
and U18117 (N_18117,N_17845,N_17808);
and U18118 (N_18118,N_17945,N_17824);
or U18119 (N_18119,N_17875,N_17807);
or U18120 (N_18120,N_17956,N_17995);
xor U18121 (N_18121,N_17851,N_17837);
nand U18122 (N_18122,N_17976,N_17846);
and U18123 (N_18123,N_17841,N_17894);
xor U18124 (N_18124,N_17908,N_17822);
and U18125 (N_18125,N_17815,N_17935);
and U18126 (N_18126,N_17844,N_17861);
nor U18127 (N_18127,N_17837,N_17975);
and U18128 (N_18128,N_17885,N_17959);
nand U18129 (N_18129,N_17847,N_17939);
nand U18130 (N_18130,N_17837,N_17855);
or U18131 (N_18131,N_17885,N_17953);
and U18132 (N_18132,N_17863,N_17874);
nor U18133 (N_18133,N_17881,N_17944);
or U18134 (N_18134,N_17800,N_17898);
nand U18135 (N_18135,N_17923,N_17943);
nor U18136 (N_18136,N_17835,N_17885);
or U18137 (N_18137,N_17917,N_17912);
or U18138 (N_18138,N_17928,N_17836);
or U18139 (N_18139,N_17883,N_17874);
nand U18140 (N_18140,N_17987,N_17976);
nand U18141 (N_18141,N_17810,N_17843);
or U18142 (N_18142,N_17849,N_17963);
or U18143 (N_18143,N_17816,N_17942);
nor U18144 (N_18144,N_17917,N_17879);
nor U18145 (N_18145,N_17916,N_17958);
or U18146 (N_18146,N_17989,N_17871);
xnor U18147 (N_18147,N_17897,N_17819);
nand U18148 (N_18148,N_17941,N_17937);
and U18149 (N_18149,N_17923,N_17916);
nor U18150 (N_18150,N_17934,N_17982);
and U18151 (N_18151,N_17870,N_17811);
xnor U18152 (N_18152,N_17857,N_17813);
xnor U18153 (N_18153,N_17874,N_17993);
nor U18154 (N_18154,N_17892,N_17956);
nor U18155 (N_18155,N_17876,N_17856);
nand U18156 (N_18156,N_17877,N_17934);
xnor U18157 (N_18157,N_17877,N_17901);
and U18158 (N_18158,N_17948,N_17970);
xor U18159 (N_18159,N_17845,N_17827);
nor U18160 (N_18160,N_17920,N_17915);
nor U18161 (N_18161,N_17987,N_17913);
xor U18162 (N_18162,N_17843,N_17934);
nand U18163 (N_18163,N_17891,N_17883);
or U18164 (N_18164,N_17871,N_17907);
and U18165 (N_18165,N_17823,N_17900);
nor U18166 (N_18166,N_17858,N_17991);
or U18167 (N_18167,N_17879,N_17949);
xnor U18168 (N_18168,N_17923,N_17881);
or U18169 (N_18169,N_17880,N_17965);
and U18170 (N_18170,N_17988,N_17888);
xor U18171 (N_18171,N_17964,N_17954);
nand U18172 (N_18172,N_17857,N_17820);
nor U18173 (N_18173,N_17815,N_17890);
or U18174 (N_18174,N_17889,N_17838);
and U18175 (N_18175,N_17981,N_17994);
xnor U18176 (N_18176,N_17825,N_17918);
or U18177 (N_18177,N_17963,N_17944);
and U18178 (N_18178,N_17937,N_17852);
and U18179 (N_18179,N_17820,N_17982);
xor U18180 (N_18180,N_17891,N_17871);
xnor U18181 (N_18181,N_17973,N_17813);
and U18182 (N_18182,N_17996,N_17824);
and U18183 (N_18183,N_17827,N_17840);
nand U18184 (N_18184,N_17834,N_17916);
or U18185 (N_18185,N_17871,N_17912);
nor U18186 (N_18186,N_17979,N_17975);
nor U18187 (N_18187,N_17828,N_17965);
xnor U18188 (N_18188,N_17980,N_17807);
or U18189 (N_18189,N_17991,N_17873);
nor U18190 (N_18190,N_17918,N_17863);
nor U18191 (N_18191,N_17868,N_17876);
xnor U18192 (N_18192,N_17907,N_17899);
and U18193 (N_18193,N_17976,N_17834);
and U18194 (N_18194,N_17873,N_17901);
nor U18195 (N_18195,N_17962,N_17937);
nand U18196 (N_18196,N_17864,N_17960);
xnor U18197 (N_18197,N_17938,N_17816);
nor U18198 (N_18198,N_17848,N_17959);
xnor U18199 (N_18199,N_17934,N_17829);
nor U18200 (N_18200,N_18121,N_18180);
or U18201 (N_18201,N_18046,N_18199);
nor U18202 (N_18202,N_18054,N_18113);
nand U18203 (N_18203,N_18143,N_18138);
or U18204 (N_18204,N_18150,N_18170);
nand U18205 (N_18205,N_18073,N_18078);
or U18206 (N_18206,N_18061,N_18177);
or U18207 (N_18207,N_18185,N_18037);
nand U18208 (N_18208,N_18144,N_18011);
xor U18209 (N_18209,N_18187,N_18049);
nor U18210 (N_18210,N_18053,N_18154);
nand U18211 (N_18211,N_18125,N_18094);
nand U18212 (N_18212,N_18083,N_18039);
xnor U18213 (N_18213,N_18171,N_18044);
nand U18214 (N_18214,N_18142,N_18184);
or U18215 (N_18215,N_18065,N_18024);
nor U18216 (N_18216,N_18147,N_18060);
nor U18217 (N_18217,N_18106,N_18156);
nand U18218 (N_18218,N_18016,N_18148);
nor U18219 (N_18219,N_18071,N_18139);
nor U18220 (N_18220,N_18015,N_18020);
nor U18221 (N_18221,N_18038,N_18152);
or U18222 (N_18222,N_18000,N_18032);
xnor U18223 (N_18223,N_18127,N_18157);
and U18224 (N_18224,N_18174,N_18081);
nand U18225 (N_18225,N_18048,N_18105);
nor U18226 (N_18226,N_18183,N_18059);
xor U18227 (N_18227,N_18196,N_18045);
nand U18228 (N_18228,N_18191,N_18128);
nor U18229 (N_18229,N_18124,N_18074);
nor U18230 (N_18230,N_18192,N_18175);
xnor U18231 (N_18231,N_18066,N_18120);
nand U18232 (N_18232,N_18093,N_18135);
or U18233 (N_18233,N_18022,N_18086);
or U18234 (N_18234,N_18136,N_18188);
xnor U18235 (N_18235,N_18146,N_18034);
xor U18236 (N_18236,N_18162,N_18092);
xnor U18237 (N_18237,N_18089,N_18197);
nor U18238 (N_18238,N_18107,N_18153);
or U18239 (N_18239,N_18067,N_18030);
or U18240 (N_18240,N_18003,N_18178);
nand U18241 (N_18241,N_18176,N_18036);
nand U18242 (N_18242,N_18064,N_18195);
nand U18243 (N_18243,N_18099,N_18096);
nor U18244 (N_18244,N_18117,N_18166);
nor U18245 (N_18245,N_18070,N_18161);
nand U18246 (N_18246,N_18155,N_18141);
nand U18247 (N_18247,N_18123,N_18190);
nand U18248 (N_18248,N_18186,N_18042);
nand U18249 (N_18249,N_18068,N_18160);
nand U18250 (N_18250,N_18017,N_18173);
xor U18251 (N_18251,N_18090,N_18026);
nand U18252 (N_18252,N_18108,N_18167);
and U18253 (N_18253,N_18057,N_18035);
nand U18254 (N_18254,N_18149,N_18122);
or U18255 (N_18255,N_18047,N_18084);
nor U18256 (N_18256,N_18012,N_18041);
nand U18257 (N_18257,N_18133,N_18088);
and U18258 (N_18258,N_18006,N_18114);
and U18259 (N_18259,N_18019,N_18013);
or U18260 (N_18260,N_18025,N_18145);
and U18261 (N_18261,N_18062,N_18029);
xor U18262 (N_18262,N_18040,N_18151);
nor U18263 (N_18263,N_18069,N_18023);
or U18264 (N_18264,N_18132,N_18172);
and U18265 (N_18265,N_18158,N_18103);
nand U18266 (N_18266,N_18119,N_18168);
or U18267 (N_18267,N_18014,N_18164);
and U18268 (N_18268,N_18010,N_18193);
xnor U18269 (N_18269,N_18002,N_18181);
xor U18270 (N_18270,N_18095,N_18087);
or U18271 (N_18271,N_18137,N_18104);
and U18272 (N_18272,N_18076,N_18009);
or U18273 (N_18273,N_18194,N_18134);
or U18274 (N_18274,N_18075,N_18031);
nor U18275 (N_18275,N_18163,N_18052);
or U18276 (N_18276,N_18116,N_18189);
xnor U18277 (N_18277,N_18159,N_18100);
nor U18278 (N_18278,N_18050,N_18109);
or U18279 (N_18279,N_18058,N_18021);
nor U18280 (N_18280,N_18043,N_18169);
nor U18281 (N_18281,N_18007,N_18102);
xnor U18282 (N_18282,N_18063,N_18129);
or U18283 (N_18283,N_18005,N_18079);
and U18284 (N_18284,N_18182,N_18118);
nand U18285 (N_18285,N_18198,N_18110);
xor U18286 (N_18286,N_18165,N_18056);
nand U18287 (N_18287,N_18018,N_18001);
or U18288 (N_18288,N_18055,N_18051);
or U18289 (N_18289,N_18080,N_18115);
and U18290 (N_18290,N_18085,N_18004);
xnor U18291 (N_18291,N_18098,N_18140);
xnor U18292 (N_18292,N_18179,N_18033);
and U18293 (N_18293,N_18077,N_18111);
or U18294 (N_18294,N_18008,N_18027);
nand U18295 (N_18295,N_18091,N_18097);
and U18296 (N_18296,N_18028,N_18082);
and U18297 (N_18297,N_18072,N_18126);
nor U18298 (N_18298,N_18131,N_18112);
nor U18299 (N_18299,N_18101,N_18130);
or U18300 (N_18300,N_18006,N_18143);
nand U18301 (N_18301,N_18198,N_18084);
or U18302 (N_18302,N_18053,N_18178);
and U18303 (N_18303,N_18101,N_18120);
and U18304 (N_18304,N_18109,N_18139);
nor U18305 (N_18305,N_18130,N_18014);
or U18306 (N_18306,N_18057,N_18186);
or U18307 (N_18307,N_18006,N_18059);
nor U18308 (N_18308,N_18110,N_18167);
nor U18309 (N_18309,N_18141,N_18110);
nor U18310 (N_18310,N_18008,N_18068);
or U18311 (N_18311,N_18080,N_18097);
nor U18312 (N_18312,N_18179,N_18196);
nand U18313 (N_18313,N_18165,N_18075);
and U18314 (N_18314,N_18144,N_18116);
xnor U18315 (N_18315,N_18090,N_18180);
nor U18316 (N_18316,N_18079,N_18119);
nor U18317 (N_18317,N_18141,N_18093);
xnor U18318 (N_18318,N_18100,N_18146);
and U18319 (N_18319,N_18117,N_18103);
xor U18320 (N_18320,N_18161,N_18025);
nor U18321 (N_18321,N_18016,N_18146);
xor U18322 (N_18322,N_18155,N_18048);
or U18323 (N_18323,N_18111,N_18057);
and U18324 (N_18324,N_18036,N_18178);
nand U18325 (N_18325,N_18129,N_18195);
nand U18326 (N_18326,N_18117,N_18116);
or U18327 (N_18327,N_18084,N_18117);
xor U18328 (N_18328,N_18048,N_18140);
or U18329 (N_18329,N_18114,N_18035);
nor U18330 (N_18330,N_18090,N_18133);
nand U18331 (N_18331,N_18006,N_18173);
nand U18332 (N_18332,N_18091,N_18149);
nand U18333 (N_18333,N_18052,N_18040);
or U18334 (N_18334,N_18100,N_18130);
nand U18335 (N_18335,N_18045,N_18064);
nor U18336 (N_18336,N_18116,N_18197);
and U18337 (N_18337,N_18151,N_18149);
nor U18338 (N_18338,N_18137,N_18112);
and U18339 (N_18339,N_18102,N_18095);
nor U18340 (N_18340,N_18182,N_18007);
xor U18341 (N_18341,N_18062,N_18183);
or U18342 (N_18342,N_18042,N_18154);
or U18343 (N_18343,N_18146,N_18029);
nor U18344 (N_18344,N_18102,N_18055);
and U18345 (N_18345,N_18053,N_18166);
and U18346 (N_18346,N_18150,N_18182);
nand U18347 (N_18347,N_18175,N_18165);
nor U18348 (N_18348,N_18102,N_18123);
and U18349 (N_18349,N_18121,N_18003);
nand U18350 (N_18350,N_18110,N_18003);
nand U18351 (N_18351,N_18022,N_18018);
xor U18352 (N_18352,N_18157,N_18014);
and U18353 (N_18353,N_18177,N_18005);
nand U18354 (N_18354,N_18096,N_18165);
or U18355 (N_18355,N_18105,N_18103);
nand U18356 (N_18356,N_18060,N_18188);
or U18357 (N_18357,N_18065,N_18108);
xor U18358 (N_18358,N_18110,N_18079);
or U18359 (N_18359,N_18144,N_18048);
xor U18360 (N_18360,N_18048,N_18015);
nand U18361 (N_18361,N_18128,N_18175);
nand U18362 (N_18362,N_18050,N_18070);
and U18363 (N_18363,N_18030,N_18192);
or U18364 (N_18364,N_18040,N_18036);
nand U18365 (N_18365,N_18191,N_18017);
xor U18366 (N_18366,N_18055,N_18174);
xor U18367 (N_18367,N_18165,N_18101);
nor U18368 (N_18368,N_18014,N_18180);
xor U18369 (N_18369,N_18199,N_18110);
nor U18370 (N_18370,N_18000,N_18164);
nor U18371 (N_18371,N_18104,N_18085);
xor U18372 (N_18372,N_18041,N_18110);
xor U18373 (N_18373,N_18163,N_18134);
nand U18374 (N_18374,N_18091,N_18041);
xnor U18375 (N_18375,N_18114,N_18088);
or U18376 (N_18376,N_18016,N_18187);
xor U18377 (N_18377,N_18025,N_18123);
nor U18378 (N_18378,N_18101,N_18071);
nand U18379 (N_18379,N_18147,N_18131);
and U18380 (N_18380,N_18172,N_18112);
and U18381 (N_18381,N_18132,N_18037);
xor U18382 (N_18382,N_18013,N_18072);
nand U18383 (N_18383,N_18128,N_18171);
and U18384 (N_18384,N_18133,N_18060);
and U18385 (N_18385,N_18025,N_18112);
xnor U18386 (N_18386,N_18006,N_18145);
nand U18387 (N_18387,N_18087,N_18034);
and U18388 (N_18388,N_18077,N_18184);
nor U18389 (N_18389,N_18141,N_18047);
nor U18390 (N_18390,N_18174,N_18118);
nor U18391 (N_18391,N_18004,N_18093);
or U18392 (N_18392,N_18135,N_18177);
and U18393 (N_18393,N_18116,N_18187);
and U18394 (N_18394,N_18005,N_18029);
xor U18395 (N_18395,N_18151,N_18153);
nor U18396 (N_18396,N_18048,N_18119);
nor U18397 (N_18397,N_18198,N_18057);
and U18398 (N_18398,N_18128,N_18199);
xnor U18399 (N_18399,N_18023,N_18054);
nor U18400 (N_18400,N_18226,N_18309);
xnor U18401 (N_18401,N_18207,N_18215);
or U18402 (N_18402,N_18393,N_18369);
xor U18403 (N_18403,N_18315,N_18323);
and U18404 (N_18404,N_18240,N_18244);
nand U18405 (N_18405,N_18253,N_18383);
xor U18406 (N_18406,N_18341,N_18306);
nor U18407 (N_18407,N_18227,N_18360);
or U18408 (N_18408,N_18345,N_18373);
nor U18409 (N_18409,N_18353,N_18209);
nor U18410 (N_18410,N_18334,N_18238);
xor U18411 (N_18411,N_18230,N_18324);
xor U18412 (N_18412,N_18302,N_18242);
nand U18413 (N_18413,N_18214,N_18250);
nand U18414 (N_18414,N_18319,N_18362);
and U18415 (N_18415,N_18274,N_18263);
or U18416 (N_18416,N_18267,N_18304);
and U18417 (N_18417,N_18228,N_18285);
and U18418 (N_18418,N_18296,N_18355);
or U18419 (N_18419,N_18299,N_18288);
nand U18420 (N_18420,N_18337,N_18248);
or U18421 (N_18421,N_18282,N_18204);
nor U18422 (N_18422,N_18245,N_18232);
nand U18423 (N_18423,N_18303,N_18284);
nand U18424 (N_18424,N_18213,N_18301);
xor U18425 (N_18425,N_18394,N_18384);
or U18426 (N_18426,N_18330,N_18203);
nand U18427 (N_18427,N_18235,N_18387);
nor U18428 (N_18428,N_18381,N_18390);
nand U18429 (N_18429,N_18208,N_18254);
xnor U18430 (N_18430,N_18222,N_18261);
xor U18431 (N_18431,N_18257,N_18367);
or U18432 (N_18432,N_18329,N_18347);
and U18433 (N_18433,N_18379,N_18243);
xor U18434 (N_18434,N_18365,N_18311);
nand U18435 (N_18435,N_18325,N_18398);
and U18436 (N_18436,N_18358,N_18357);
nand U18437 (N_18437,N_18395,N_18295);
nand U18438 (N_18438,N_18221,N_18291);
xnor U18439 (N_18439,N_18316,N_18371);
or U18440 (N_18440,N_18307,N_18259);
nand U18441 (N_18441,N_18231,N_18270);
xnor U18442 (N_18442,N_18246,N_18287);
nand U18443 (N_18443,N_18312,N_18266);
and U18444 (N_18444,N_18351,N_18342);
or U18445 (N_18445,N_18352,N_18374);
nor U18446 (N_18446,N_18262,N_18382);
and U18447 (N_18447,N_18300,N_18280);
nand U18448 (N_18448,N_18366,N_18335);
or U18449 (N_18449,N_18210,N_18224);
xnor U18450 (N_18450,N_18255,N_18361);
or U18451 (N_18451,N_18348,N_18219);
nor U18452 (N_18452,N_18294,N_18350);
nor U18453 (N_18453,N_18217,N_18239);
or U18454 (N_18454,N_18375,N_18308);
nor U18455 (N_18455,N_18223,N_18326);
nand U18456 (N_18456,N_18377,N_18289);
xor U18457 (N_18457,N_18317,N_18310);
nand U18458 (N_18458,N_18290,N_18336);
xor U18459 (N_18459,N_18380,N_18252);
or U18460 (N_18460,N_18305,N_18272);
or U18461 (N_18461,N_18322,N_18225);
xnor U18462 (N_18462,N_18389,N_18376);
and U18463 (N_18463,N_18281,N_18229);
xnor U18464 (N_18464,N_18397,N_18396);
or U18465 (N_18465,N_18268,N_18320);
nand U18466 (N_18466,N_18216,N_18349);
and U18467 (N_18467,N_18314,N_18364);
xnor U18468 (N_18468,N_18333,N_18321);
xnor U18469 (N_18469,N_18318,N_18385);
and U18470 (N_18470,N_18265,N_18368);
nor U18471 (N_18471,N_18200,N_18269);
xnor U18472 (N_18472,N_18338,N_18332);
nand U18473 (N_18473,N_18339,N_18344);
and U18474 (N_18474,N_18392,N_18346);
or U18475 (N_18475,N_18372,N_18391);
nor U18476 (N_18476,N_18343,N_18328);
nor U18477 (N_18477,N_18279,N_18297);
nand U18478 (N_18478,N_18206,N_18256);
and U18479 (N_18479,N_18264,N_18247);
or U18480 (N_18480,N_18340,N_18388);
nand U18481 (N_18481,N_18399,N_18273);
nand U18482 (N_18482,N_18276,N_18220);
nor U18483 (N_18483,N_18370,N_18260);
nor U18484 (N_18484,N_18354,N_18298);
or U18485 (N_18485,N_18212,N_18234);
and U18486 (N_18486,N_18277,N_18237);
xor U18487 (N_18487,N_18271,N_18211);
xor U18488 (N_18488,N_18202,N_18286);
nor U18489 (N_18489,N_18275,N_18218);
nand U18490 (N_18490,N_18278,N_18249);
and U18491 (N_18491,N_18236,N_18331);
or U18492 (N_18492,N_18356,N_18251);
xor U18493 (N_18493,N_18292,N_18293);
nor U18494 (N_18494,N_18378,N_18363);
nor U18495 (N_18495,N_18327,N_18386);
nand U18496 (N_18496,N_18201,N_18205);
or U18497 (N_18497,N_18313,N_18233);
or U18498 (N_18498,N_18283,N_18241);
or U18499 (N_18499,N_18258,N_18359);
or U18500 (N_18500,N_18301,N_18328);
xor U18501 (N_18501,N_18229,N_18291);
nor U18502 (N_18502,N_18375,N_18208);
xor U18503 (N_18503,N_18291,N_18367);
nand U18504 (N_18504,N_18287,N_18347);
nand U18505 (N_18505,N_18381,N_18269);
nor U18506 (N_18506,N_18272,N_18323);
nor U18507 (N_18507,N_18205,N_18259);
xor U18508 (N_18508,N_18333,N_18235);
nor U18509 (N_18509,N_18322,N_18361);
nand U18510 (N_18510,N_18324,N_18284);
xnor U18511 (N_18511,N_18220,N_18395);
nand U18512 (N_18512,N_18218,N_18206);
nand U18513 (N_18513,N_18330,N_18334);
and U18514 (N_18514,N_18356,N_18242);
xnor U18515 (N_18515,N_18261,N_18263);
and U18516 (N_18516,N_18373,N_18297);
or U18517 (N_18517,N_18326,N_18217);
nor U18518 (N_18518,N_18227,N_18348);
nand U18519 (N_18519,N_18225,N_18375);
and U18520 (N_18520,N_18294,N_18308);
and U18521 (N_18521,N_18298,N_18229);
nor U18522 (N_18522,N_18257,N_18215);
xor U18523 (N_18523,N_18239,N_18213);
and U18524 (N_18524,N_18365,N_18209);
nand U18525 (N_18525,N_18328,N_18325);
and U18526 (N_18526,N_18328,N_18292);
xor U18527 (N_18527,N_18239,N_18256);
xor U18528 (N_18528,N_18268,N_18292);
or U18529 (N_18529,N_18246,N_18230);
nor U18530 (N_18530,N_18279,N_18223);
nand U18531 (N_18531,N_18228,N_18302);
nand U18532 (N_18532,N_18217,N_18240);
nand U18533 (N_18533,N_18261,N_18355);
xnor U18534 (N_18534,N_18289,N_18317);
nand U18535 (N_18535,N_18330,N_18228);
nor U18536 (N_18536,N_18205,N_18287);
nor U18537 (N_18537,N_18344,N_18232);
xor U18538 (N_18538,N_18306,N_18349);
nor U18539 (N_18539,N_18382,N_18278);
xnor U18540 (N_18540,N_18343,N_18224);
or U18541 (N_18541,N_18297,N_18383);
and U18542 (N_18542,N_18368,N_18314);
nand U18543 (N_18543,N_18358,N_18245);
nor U18544 (N_18544,N_18261,N_18349);
or U18545 (N_18545,N_18236,N_18260);
nor U18546 (N_18546,N_18366,N_18200);
xnor U18547 (N_18547,N_18398,N_18246);
xnor U18548 (N_18548,N_18303,N_18322);
nor U18549 (N_18549,N_18279,N_18298);
nor U18550 (N_18550,N_18314,N_18339);
or U18551 (N_18551,N_18226,N_18201);
and U18552 (N_18552,N_18273,N_18253);
and U18553 (N_18553,N_18285,N_18295);
and U18554 (N_18554,N_18319,N_18276);
xnor U18555 (N_18555,N_18367,N_18258);
and U18556 (N_18556,N_18236,N_18295);
or U18557 (N_18557,N_18226,N_18321);
xor U18558 (N_18558,N_18394,N_18260);
or U18559 (N_18559,N_18240,N_18267);
or U18560 (N_18560,N_18363,N_18235);
and U18561 (N_18561,N_18321,N_18292);
xor U18562 (N_18562,N_18322,N_18273);
and U18563 (N_18563,N_18202,N_18360);
xor U18564 (N_18564,N_18336,N_18396);
nand U18565 (N_18565,N_18348,N_18294);
and U18566 (N_18566,N_18286,N_18219);
xor U18567 (N_18567,N_18237,N_18347);
and U18568 (N_18568,N_18399,N_18258);
or U18569 (N_18569,N_18202,N_18317);
nor U18570 (N_18570,N_18253,N_18261);
nand U18571 (N_18571,N_18210,N_18320);
xor U18572 (N_18572,N_18249,N_18358);
and U18573 (N_18573,N_18205,N_18340);
xor U18574 (N_18574,N_18252,N_18368);
xnor U18575 (N_18575,N_18263,N_18273);
or U18576 (N_18576,N_18238,N_18208);
or U18577 (N_18577,N_18256,N_18310);
xor U18578 (N_18578,N_18279,N_18219);
xor U18579 (N_18579,N_18381,N_18397);
or U18580 (N_18580,N_18297,N_18340);
xnor U18581 (N_18581,N_18297,N_18328);
and U18582 (N_18582,N_18297,N_18352);
and U18583 (N_18583,N_18311,N_18307);
nand U18584 (N_18584,N_18279,N_18295);
nor U18585 (N_18585,N_18297,N_18371);
and U18586 (N_18586,N_18274,N_18333);
nor U18587 (N_18587,N_18288,N_18241);
or U18588 (N_18588,N_18393,N_18340);
nor U18589 (N_18589,N_18241,N_18270);
xor U18590 (N_18590,N_18227,N_18314);
or U18591 (N_18591,N_18219,N_18255);
nand U18592 (N_18592,N_18279,N_18258);
nand U18593 (N_18593,N_18326,N_18210);
nand U18594 (N_18594,N_18206,N_18327);
nand U18595 (N_18595,N_18314,N_18210);
nor U18596 (N_18596,N_18283,N_18225);
nor U18597 (N_18597,N_18312,N_18279);
nor U18598 (N_18598,N_18309,N_18316);
or U18599 (N_18599,N_18278,N_18276);
or U18600 (N_18600,N_18545,N_18521);
or U18601 (N_18601,N_18411,N_18450);
or U18602 (N_18602,N_18441,N_18554);
nand U18603 (N_18603,N_18562,N_18525);
nor U18604 (N_18604,N_18446,N_18409);
and U18605 (N_18605,N_18419,N_18460);
nor U18606 (N_18606,N_18566,N_18591);
and U18607 (N_18607,N_18474,N_18570);
xor U18608 (N_18608,N_18414,N_18582);
nand U18609 (N_18609,N_18470,N_18538);
nor U18610 (N_18610,N_18451,N_18468);
or U18611 (N_18611,N_18431,N_18506);
or U18612 (N_18612,N_18495,N_18483);
nor U18613 (N_18613,N_18498,N_18432);
nand U18614 (N_18614,N_18514,N_18406);
nor U18615 (N_18615,N_18449,N_18471);
nor U18616 (N_18616,N_18539,N_18421);
and U18617 (N_18617,N_18412,N_18430);
or U18618 (N_18618,N_18489,N_18465);
or U18619 (N_18619,N_18475,N_18546);
nor U18620 (N_18620,N_18517,N_18523);
nand U18621 (N_18621,N_18462,N_18416);
or U18622 (N_18622,N_18590,N_18408);
nand U18623 (N_18623,N_18487,N_18556);
nor U18624 (N_18624,N_18583,N_18469);
nor U18625 (N_18625,N_18433,N_18456);
nor U18626 (N_18626,N_18494,N_18404);
xor U18627 (N_18627,N_18434,N_18544);
or U18628 (N_18628,N_18422,N_18575);
nand U18629 (N_18629,N_18476,N_18400);
or U18630 (N_18630,N_18407,N_18572);
nand U18631 (N_18631,N_18531,N_18542);
xor U18632 (N_18632,N_18423,N_18427);
nand U18633 (N_18633,N_18459,N_18505);
xor U18634 (N_18634,N_18574,N_18563);
xor U18635 (N_18635,N_18442,N_18481);
or U18636 (N_18636,N_18508,N_18581);
or U18637 (N_18637,N_18402,N_18437);
or U18638 (N_18638,N_18403,N_18594);
nor U18639 (N_18639,N_18596,N_18597);
or U18640 (N_18640,N_18503,N_18405);
xnor U18641 (N_18641,N_18435,N_18458);
nor U18642 (N_18642,N_18533,N_18488);
or U18643 (N_18643,N_18477,N_18499);
nor U18644 (N_18644,N_18492,N_18558);
xnor U18645 (N_18645,N_18578,N_18467);
or U18646 (N_18646,N_18576,N_18510);
nand U18647 (N_18647,N_18453,N_18420);
xnor U18648 (N_18648,N_18568,N_18580);
or U18649 (N_18649,N_18532,N_18444);
and U18650 (N_18650,N_18513,N_18585);
xor U18651 (N_18651,N_18452,N_18579);
and U18652 (N_18652,N_18577,N_18536);
and U18653 (N_18653,N_18482,N_18463);
or U18654 (N_18654,N_18418,N_18550);
nor U18655 (N_18655,N_18543,N_18526);
and U18656 (N_18656,N_18501,N_18518);
nor U18657 (N_18657,N_18569,N_18565);
xnor U18658 (N_18658,N_18428,N_18493);
xnor U18659 (N_18659,N_18448,N_18593);
nor U18660 (N_18660,N_18541,N_18595);
nand U18661 (N_18661,N_18571,N_18537);
and U18662 (N_18662,N_18424,N_18520);
nor U18663 (N_18663,N_18425,N_18485);
nand U18664 (N_18664,N_18511,N_18436);
xor U18665 (N_18665,N_18560,N_18496);
nor U18666 (N_18666,N_18417,N_18557);
xor U18667 (N_18667,N_18478,N_18454);
or U18668 (N_18668,N_18559,N_18561);
or U18669 (N_18669,N_18586,N_18551);
nor U18670 (N_18670,N_18464,N_18549);
nand U18671 (N_18671,N_18516,N_18429);
nand U18672 (N_18672,N_18527,N_18415);
nor U18673 (N_18673,N_18472,N_18587);
xnor U18674 (N_18674,N_18445,N_18484);
nor U18675 (N_18675,N_18455,N_18598);
nand U18676 (N_18676,N_18447,N_18401);
and U18677 (N_18677,N_18473,N_18443);
or U18678 (N_18678,N_18410,N_18491);
xnor U18679 (N_18679,N_18479,N_18555);
nor U18680 (N_18680,N_18530,N_18519);
and U18681 (N_18681,N_18457,N_18515);
or U18682 (N_18682,N_18573,N_18413);
xnor U18683 (N_18683,N_18548,N_18461);
nand U18684 (N_18684,N_18438,N_18507);
or U18685 (N_18685,N_18528,N_18584);
nor U18686 (N_18686,N_18552,N_18504);
nor U18687 (N_18687,N_18439,N_18440);
xnor U18688 (N_18688,N_18466,N_18540);
and U18689 (N_18689,N_18480,N_18502);
nor U18690 (N_18690,N_18534,N_18564);
and U18691 (N_18691,N_18588,N_18490);
xnor U18692 (N_18692,N_18529,N_18500);
or U18693 (N_18693,N_18599,N_18567);
and U18694 (N_18694,N_18524,N_18547);
and U18695 (N_18695,N_18589,N_18512);
or U18696 (N_18696,N_18535,N_18553);
xor U18697 (N_18697,N_18497,N_18426);
and U18698 (N_18698,N_18522,N_18509);
and U18699 (N_18699,N_18592,N_18486);
xor U18700 (N_18700,N_18540,N_18404);
xnor U18701 (N_18701,N_18573,N_18480);
nor U18702 (N_18702,N_18453,N_18459);
xnor U18703 (N_18703,N_18479,N_18557);
and U18704 (N_18704,N_18409,N_18528);
and U18705 (N_18705,N_18478,N_18579);
nor U18706 (N_18706,N_18449,N_18549);
nor U18707 (N_18707,N_18507,N_18497);
nand U18708 (N_18708,N_18455,N_18587);
nand U18709 (N_18709,N_18513,N_18459);
nand U18710 (N_18710,N_18549,N_18505);
or U18711 (N_18711,N_18429,N_18411);
or U18712 (N_18712,N_18447,N_18559);
and U18713 (N_18713,N_18450,N_18505);
xnor U18714 (N_18714,N_18405,N_18492);
and U18715 (N_18715,N_18517,N_18568);
nor U18716 (N_18716,N_18472,N_18546);
xnor U18717 (N_18717,N_18578,N_18584);
nand U18718 (N_18718,N_18571,N_18458);
nand U18719 (N_18719,N_18435,N_18403);
and U18720 (N_18720,N_18541,N_18567);
xnor U18721 (N_18721,N_18531,N_18478);
and U18722 (N_18722,N_18506,N_18461);
and U18723 (N_18723,N_18436,N_18415);
and U18724 (N_18724,N_18574,N_18552);
nor U18725 (N_18725,N_18549,N_18467);
nor U18726 (N_18726,N_18562,N_18534);
and U18727 (N_18727,N_18430,N_18438);
xor U18728 (N_18728,N_18509,N_18460);
nand U18729 (N_18729,N_18478,N_18561);
or U18730 (N_18730,N_18405,N_18417);
xor U18731 (N_18731,N_18542,N_18446);
nor U18732 (N_18732,N_18477,N_18425);
nor U18733 (N_18733,N_18597,N_18580);
or U18734 (N_18734,N_18567,N_18577);
or U18735 (N_18735,N_18472,N_18452);
xor U18736 (N_18736,N_18572,N_18593);
or U18737 (N_18737,N_18442,N_18528);
nand U18738 (N_18738,N_18476,N_18463);
or U18739 (N_18739,N_18550,N_18537);
nor U18740 (N_18740,N_18421,N_18419);
xor U18741 (N_18741,N_18536,N_18553);
nand U18742 (N_18742,N_18480,N_18415);
nor U18743 (N_18743,N_18492,N_18583);
xnor U18744 (N_18744,N_18596,N_18576);
or U18745 (N_18745,N_18454,N_18419);
nor U18746 (N_18746,N_18419,N_18414);
and U18747 (N_18747,N_18597,N_18583);
nand U18748 (N_18748,N_18528,N_18570);
and U18749 (N_18749,N_18583,N_18479);
or U18750 (N_18750,N_18475,N_18428);
nand U18751 (N_18751,N_18509,N_18498);
nand U18752 (N_18752,N_18438,N_18569);
nand U18753 (N_18753,N_18467,N_18561);
nor U18754 (N_18754,N_18480,N_18529);
nand U18755 (N_18755,N_18440,N_18510);
nor U18756 (N_18756,N_18475,N_18478);
nor U18757 (N_18757,N_18567,N_18560);
or U18758 (N_18758,N_18444,N_18591);
nand U18759 (N_18759,N_18475,N_18430);
xnor U18760 (N_18760,N_18519,N_18432);
nor U18761 (N_18761,N_18411,N_18561);
nand U18762 (N_18762,N_18591,N_18572);
xnor U18763 (N_18763,N_18524,N_18585);
nand U18764 (N_18764,N_18525,N_18421);
nand U18765 (N_18765,N_18446,N_18439);
xnor U18766 (N_18766,N_18597,N_18442);
or U18767 (N_18767,N_18433,N_18425);
xnor U18768 (N_18768,N_18402,N_18513);
and U18769 (N_18769,N_18588,N_18536);
nor U18770 (N_18770,N_18509,N_18504);
or U18771 (N_18771,N_18573,N_18546);
nor U18772 (N_18772,N_18564,N_18405);
nand U18773 (N_18773,N_18498,N_18585);
nor U18774 (N_18774,N_18596,N_18534);
nand U18775 (N_18775,N_18414,N_18482);
and U18776 (N_18776,N_18419,N_18552);
and U18777 (N_18777,N_18458,N_18441);
nand U18778 (N_18778,N_18545,N_18518);
nand U18779 (N_18779,N_18561,N_18534);
xnor U18780 (N_18780,N_18493,N_18438);
xnor U18781 (N_18781,N_18528,N_18486);
nand U18782 (N_18782,N_18533,N_18557);
and U18783 (N_18783,N_18557,N_18532);
or U18784 (N_18784,N_18477,N_18412);
nand U18785 (N_18785,N_18476,N_18565);
nor U18786 (N_18786,N_18586,N_18448);
xnor U18787 (N_18787,N_18494,N_18570);
and U18788 (N_18788,N_18435,N_18454);
and U18789 (N_18789,N_18592,N_18532);
nor U18790 (N_18790,N_18503,N_18567);
nor U18791 (N_18791,N_18570,N_18577);
and U18792 (N_18792,N_18586,N_18491);
or U18793 (N_18793,N_18443,N_18584);
xnor U18794 (N_18794,N_18583,N_18503);
xor U18795 (N_18795,N_18500,N_18598);
or U18796 (N_18796,N_18429,N_18408);
xor U18797 (N_18797,N_18538,N_18565);
nor U18798 (N_18798,N_18590,N_18541);
nand U18799 (N_18799,N_18594,N_18574);
or U18800 (N_18800,N_18661,N_18763);
and U18801 (N_18801,N_18774,N_18624);
nand U18802 (N_18802,N_18625,N_18606);
nor U18803 (N_18803,N_18717,N_18758);
nor U18804 (N_18804,N_18618,N_18724);
and U18805 (N_18805,N_18674,N_18739);
nor U18806 (N_18806,N_18619,N_18630);
and U18807 (N_18807,N_18643,N_18760);
and U18808 (N_18808,N_18692,N_18667);
xnor U18809 (N_18809,N_18783,N_18778);
and U18810 (N_18810,N_18775,N_18652);
xnor U18811 (N_18811,N_18700,N_18642);
and U18812 (N_18812,N_18715,N_18638);
nor U18813 (N_18813,N_18666,N_18679);
and U18814 (N_18814,N_18678,N_18664);
xnor U18815 (N_18815,N_18725,N_18626);
nand U18816 (N_18816,N_18653,N_18749);
xor U18817 (N_18817,N_18672,N_18733);
or U18818 (N_18818,N_18776,N_18744);
and U18819 (N_18819,N_18721,N_18622);
nand U18820 (N_18820,N_18699,N_18732);
nand U18821 (N_18821,N_18704,N_18691);
nor U18822 (N_18822,N_18791,N_18735);
and U18823 (N_18823,N_18787,N_18604);
nand U18824 (N_18824,N_18779,N_18714);
and U18825 (N_18825,N_18764,N_18756);
nor U18826 (N_18826,N_18670,N_18723);
xnor U18827 (N_18827,N_18683,N_18798);
nand U18828 (N_18828,N_18752,N_18689);
nor U18829 (N_18829,N_18617,N_18680);
nor U18830 (N_18830,N_18633,N_18623);
nor U18831 (N_18831,N_18757,N_18637);
or U18832 (N_18832,N_18602,N_18611);
nand U18833 (N_18833,N_18712,N_18770);
and U18834 (N_18834,N_18707,N_18709);
xnor U18835 (N_18835,N_18729,N_18645);
xor U18836 (N_18836,N_18655,N_18613);
and U18837 (N_18837,N_18656,N_18659);
and U18838 (N_18838,N_18657,N_18675);
nor U18839 (N_18839,N_18647,N_18658);
and U18840 (N_18840,N_18650,N_18706);
nand U18841 (N_18841,N_18765,N_18614);
or U18842 (N_18842,N_18740,N_18671);
nand U18843 (N_18843,N_18681,N_18730);
nand U18844 (N_18844,N_18665,N_18693);
or U18845 (N_18845,N_18748,N_18685);
nand U18846 (N_18846,N_18621,N_18651);
nor U18847 (N_18847,N_18690,N_18603);
nand U18848 (N_18848,N_18608,N_18792);
nand U18849 (N_18849,N_18629,N_18640);
nand U18850 (N_18850,N_18612,N_18795);
nor U18851 (N_18851,N_18677,N_18694);
or U18852 (N_18852,N_18610,N_18703);
xnor U18853 (N_18853,N_18627,N_18639);
nor U18854 (N_18854,N_18719,N_18766);
or U18855 (N_18855,N_18772,N_18669);
and U18856 (N_18856,N_18620,N_18785);
nor U18857 (N_18857,N_18796,N_18701);
xnor U18858 (N_18858,N_18648,N_18695);
nand U18859 (N_18859,N_18663,N_18747);
or U18860 (N_18860,N_18682,N_18716);
nand U18861 (N_18861,N_18790,N_18781);
nor U18862 (N_18862,N_18754,N_18722);
and U18863 (N_18863,N_18718,N_18607);
xor U18864 (N_18864,N_18726,N_18759);
xor U18865 (N_18865,N_18710,N_18762);
and U18866 (N_18866,N_18777,N_18780);
nor U18867 (N_18867,N_18646,N_18686);
nand U18868 (N_18868,N_18676,N_18734);
nor U18869 (N_18869,N_18746,N_18649);
xnor U18870 (N_18870,N_18673,N_18768);
xnor U18871 (N_18871,N_18727,N_18767);
nand U18872 (N_18872,N_18794,N_18684);
and U18873 (N_18873,N_18713,N_18687);
nand U18874 (N_18874,N_18741,N_18697);
nand U18875 (N_18875,N_18668,N_18662);
xor U18876 (N_18876,N_18745,N_18631);
xnor U18877 (N_18877,N_18743,N_18696);
and U18878 (N_18878,N_18742,N_18786);
xnor U18879 (N_18879,N_18751,N_18635);
nand U18880 (N_18880,N_18615,N_18605);
xnor U18881 (N_18881,N_18788,N_18688);
nor U18882 (N_18882,N_18769,N_18797);
and U18883 (N_18883,N_18782,N_18736);
and U18884 (N_18884,N_18600,N_18711);
or U18885 (N_18885,N_18789,N_18632);
nor U18886 (N_18886,N_18616,N_18771);
and U18887 (N_18887,N_18702,N_18644);
nor U18888 (N_18888,N_18601,N_18750);
xnor U18889 (N_18889,N_18753,N_18737);
nor U18890 (N_18890,N_18784,N_18720);
nor U18891 (N_18891,N_18728,N_18698);
or U18892 (N_18892,N_18773,N_18793);
xnor U18893 (N_18893,N_18761,N_18654);
nor U18894 (N_18894,N_18609,N_18799);
or U18895 (N_18895,N_18636,N_18660);
or U18896 (N_18896,N_18628,N_18708);
and U18897 (N_18897,N_18755,N_18634);
nor U18898 (N_18898,N_18738,N_18731);
nand U18899 (N_18899,N_18705,N_18641);
or U18900 (N_18900,N_18758,N_18750);
and U18901 (N_18901,N_18621,N_18755);
or U18902 (N_18902,N_18734,N_18711);
and U18903 (N_18903,N_18690,N_18668);
or U18904 (N_18904,N_18600,N_18617);
nand U18905 (N_18905,N_18708,N_18677);
or U18906 (N_18906,N_18712,N_18649);
or U18907 (N_18907,N_18668,N_18632);
nor U18908 (N_18908,N_18709,N_18740);
or U18909 (N_18909,N_18636,N_18659);
nor U18910 (N_18910,N_18667,N_18677);
nor U18911 (N_18911,N_18632,N_18759);
or U18912 (N_18912,N_18745,N_18756);
nor U18913 (N_18913,N_18649,N_18617);
nor U18914 (N_18914,N_18611,N_18640);
nor U18915 (N_18915,N_18714,N_18798);
nor U18916 (N_18916,N_18664,N_18617);
and U18917 (N_18917,N_18777,N_18639);
nor U18918 (N_18918,N_18743,N_18729);
nor U18919 (N_18919,N_18668,N_18752);
and U18920 (N_18920,N_18657,N_18620);
xor U18921 (N_18921,N_18605,N_18788);
or U18922 (N_18922,N_18791,N_18721);
xor U18923 (N_18923,N_18755,N_18655);
and U18924 (N_18924,N_18781,N_18718);
and U18925 (N_18925,N_18737,N_18651);
nor U18926 (N_18926,N_18731,N_18765);
xnor U18927 (N_18927,N_18621,N_18703);
or U18928 (N_18928,N_18780,N_18741);
nor U18929 (N_18929,N_18669,N_18719);
or U18930 (N_18930,N_18720,N_18741);
and U18931 (N_18931,N_18613,N_18617);
xor U18932 (N_18932,N_18658,N_18703);
nand U18933 (N_18933,N_18730,N_18634);
nor U18934 (N_18934,N_18607,N_18724);
xnor U18935 (N_18935,N_18733,N_18780);
and U18936 (N_18936,N_18763,N_18724);
or U18937 (N_18937,N_18690,N_18645);
and U18938 (N_18938,N_18660,N_18662);
xnor U18939 (N_18939,N_18723,N_18634);
xnor U18940 (N_18940,N_18783,N_18676);
or U18941 (N_18941,N_18715,N_18689);
and U18942 (N_18942,N_18682,N_18715);
xor U18943 (N_18943,N_18757,N_18799);
nand U18944 (N_18944,N_18763,N_18677);
xor U18945 (N_18945,N_18618,N_18677);
nor U18946 (N_18946,N_18642,N_18694);
nand U18947 (N_18947,N_18655,N_18785);
or U18948 (N_18948,N_18772,N_18725);
nand U18949 (N_18949,N_18763,N_18744);
nand U18950 (N_18950,N_18728,N_18681);
xor U18951 (N_18951,N_18617,N_18697);
or U18952 (N_18952,N_18732,N_18789);
and U18953 (N_18953,N_18714,N_18673);
nor U18954 (N_18954,N_18624,N_18719);
or U18955 (N_18955,N_18703,N_18740);
or U18956 (N_18956,N_18705,N_18693);
nor U18957 (N_18957,N_18733,N_18639);
or U18958 (N_18958,N_18693,N_18646);
nand U18959 (N_18959,N_18701,N_18626);
nor U18960 (N_18960,N_18746,N_18795);
or U18961 (N_18961,N_18732,N_18744);
xor U18962 (N_18962,N_18652,N_18735);
and U18963 (N_18963,N_18733,N_18616);
nor U18964 (N_18964,N_18633,N_18618);
nor U18965 (N_18965,N_18763,N_18786);
xor U18966 (N_18966,N_18795,N_18796);
and U18967 (N_18967,N_18634,N_18725);
xor U18968 (N_18968,N_18621,N_18788);
and U18969 (N_18969,N_18784,N_18771);
nand U18970 (N_18970,N_18663,N_18745);
nor U18971 (N_18971,N_18775,N_18692);
or U18972 (N_18972,N_18626,N_18718);
nor U18973 (N_18973,N_18683,N_18715);
nand U18974 (N_18974,N_18734,N_18759);
nand U18975 (N_18975,N_18793,N_18756);
nand U18976 (N_18976,N_18772,N_18709);
and U18977 (N_18977,N_18736,N_18613);
nand U18978 (N_18978,N_18603,N_18777);
xor U18979 (N_18979,N_18766,N_18605);
nand U18980 (N_18980,N_18768,N_18699);
and U18981 (N_18981,N_18754,N_18760);
xnor U18982 (N_18982,N_18699,N_18795);
xor U18983 (N_18983,N_18625,N_18609);
and U18984 (N_18984,N_18742,N_18795);
nand U18985 (N_18985,N_18684,N_18753);
xnor U18986 (N_18986,N_18627,N_18617);
or U18987 (N_18987,N_18714,N_18748);
xnor U18988 (N_18988,N_18742,N_18639);
nand U18989 (N_18989,N_18739,N_18606);
and U18990 (N_18990,N_18647,N_18793);
or U18991 (N_18991,N_18717,N_18640);
nor U18992 (N_18992,N_18735,N_18678);
nand U18993 (N_18993,N_18709,N_18608);
nand U18994 (N_18994,N_18749,N_18693);
nand U18995 (N_18995,N_18769,N_18753);
nor U18996 (N_18996,N_18659,N_18722);
or U18997 (N_18997,N_18759,N_18750);
xor U18998 (N_18998,N_18649,N_18771);
xnor U18999 (N_18999,N_18711,N_18645);
nand U19000 (N_19000,N_18822,N_18886);
xnor U19001 (N_19001,N_18838,N_18939);
xor U19002 (N_19002,N_18846,N_18821);
or U19003 (N_19003,N_18842,N_18930);
nand U19004 (N_19004,N_18830,N_18924);
or U19005 (N_19005,N_18909,N_18845);
nor U19006 (N_19006,N_18938,N_18804);
or U19007 (N_19007,N_18933,N_18835);
nand U19008 (N_19008,N_18942,N_18992);
and U19009 (N_19009,N_18919,N_18853);
nor U19010 (N_19010,N_18917,N_18827);
nand U19011 (N_19011,N_18994,N_18892);
or U19012 (N_19012,N_18864,N_18894);
or U19013 (N_19013,N_18929,N_18801);
nor U19014 (N_19014,N_18854,N_18876);
nand U19015 (N_19015,N_18998,N_18884);
or U19016 (N_19016,N_18972,N_18875);
and U19017 (N_19017,N_18979,N_18848);
xor U19018 (N_19018,N_18840,N_18809);
nor U19019 (N_19019,N_18949,N_18996);
xnor U19020 (N_19020,N_18953,N_18865);
xnor U19021 (N_19021,N_18993,N_18916);
nand U19022 (N_19022,N_18817,N_18813);
nand U19023 (N_19023,N_18831,N_18874);
or U19024 (N_19024,N_18815,N_18877);
xor U19025 (N_19025,N_18971,N_18983);
or U19026 (N_19026,N_18989,N_18987);
xor U19027 (N_19027,N_18948,N_18891);
and U19028 (N_19028,N_18986,N_18873);
nor U19029 (N_19029,N_18946,N_18910);
nand U19030 (N_19030,N_18926,N_18920);
xnor U19031 (N_19031,N_18834,N_18960);
nor U19032 (N_19032,N_18837,N_18867);
nor U19033 (N_19033,N_18925,N_18912);
nor U19034 (N_19034,N_18961,N_18857);
and U19035 (N_19035,N_18868,N_18870);
xnor U19036 (N_19036,N_18962,N_18914);
nand U19037 (N_19037,N_18955,N_18880);
nor U19038 (N_19038,N_18847,N_18802);
xnor U19039 (N_19039,N_18881,N_18940);
or U19040 (N_19040,N_18849,N_18969);
and U19041 (N_19041,N_18997,N_18851);
nand U19042 (N_19042,N_18990,N_18820);
and U19043 (N_19043,N_18826,N_18980);
nand U19044 (N_19044,N_18843,N_18952);
or U19045 (N_19045,N_18887,N_18812);
or U19046 (N_19046,N_18800,N_18988);
xnor U19047 (N_19047,N_18860,N_18901);
nor U19048 (N_19048,N_18811,N_18839);
and U19049 (N_19049,N_18890,N_18808);
nand U19050 (N_19050,N_18819,N_18810);
and U19051 (N_19051,N_18844,N_18906);
and U19052 (N_19052,N_18937,N_18967);
nand U19053 (N_19053,N_18828,N_18872);
or U19054 (N_19054,N_18833,N_18985);
xnor U19055 (N_19055,N_18941,N_18871);
nor U19056 (N_19056,N_18858,N_18862);
or U19057 (N_19057,N_18861,N_18902);
or U19058 (N_19058,N_18883,N_18899);
or U19059 (N_19059,N_18896,N_18970);
nand U19060 (N_19060,N_18977,N_18856);
xnor U19061 (N_19061,N_18878,N_18911);
xnor U19062 (N_19062,N_18931,N_18841);
and U19063 (N_19063,N_18824,N_18895);
nor U19064 (N_19064,N_18978,N_18951);
and U19065 (N_19065,N_18968,N_18921);
xnor U19066 (N_19066,N_18943,N_18958);
xor U19067 (N_19067,N_18947,N_18855);
and U19068 (N_19068,N_18832,N_18866);
nor U19069 (N_19069,N_18957,N_18806);
xnor U19070 (N_19070,N_18918,N_18915);
xor U19071 (N_19071,N_18974,N_18869);
xor U19072 (N_19072,N_18818,N_18807);
xnor U19073 (N_19073,N_18932,N_18905);
and U19074 (N_19074,N_18963,N_18803);
nor U19075 (N_19075,N_18852,N_18825);
nand U19076 (N_19076,N_18836,N_18882);
nand U19077 (N_19077,N_18956,N_18814);
nor U19078 (N_19078,N_18888,N_18816);
or U19079 (N_19079,N_18823,N_18975);
nor U19080 (N_19080,N_18950,N_18965);
and U19081 (N_19081,N_18805,N_18954);
and U19082 (N_19082,N_18934,N_18973);
and U19083 (N_19083,N_18959,N_18928);
nand U19084 (N_19084,N_18984,N_18964);
nand U19085 (N_19085,N_18927,N_18976);
nand U19086 (N_19086,N_18863,N_18999);
or U19087 (N_19087,N_18885,N_18859);
nor U19088 (N_19088,N_18893,N_18907);
nand U19089 (N_19089,N_18908,N_18922);
nor U19090 (N_19090,N_18936,N_18904);
and U19091 (N_19091,N_18898,N_18829);
xnor U19092 (N_19092,N_18982,N_18897);
xor U19093 (N_19093,N_18900,N_18850);
or U19094 (N_19094,N_18995,N_18903);
xnor U19095 (N_19095,N_18945,N_18889);
or U19096 (N_19096,N_18944,N_18879);
and U19097 (N_19097,N_18991,N_18923);
and U19098 (N_19098,N_18935,N_18981);
or U19099 (N_19099,N_18913,N_18966);
or U19100 (N_19100,N_18821,N_18875);
xnor U19101 (N_19101,N_18854,N_18906);
nor U19102 (N_19102,N_18963,N_18922);
nor U19103 (N_19103,N_18833,N_18981);
nand U19104 (N_19104,N_18933,N_18876);
xor U19105 (N_19105,N_18972,N_18952);
or U19106 (N_19106,N_18995,N_18913);
and U19107 (N_19107,N_18952,N_18962);
nand U19108 (N_19108,N_18822,N_18989);
and U19109 (N_19109,N_18922,N_18890);
nand U19110 (N_19110,N_18953,N_18946);
and U19111 (N_19111,N_18822,N_18922);
or U19112 (N_19112,N_18985,N_18853);
and U19113 (N_19113,N_18957,N_18858);
nor U19114 (N_19114,N_18884,N_18995);
and U19115 (N_19115,N_18839,N_18807);
nor U19116 (N_19116,N_18949,N_18979);
and U19117 (N_19117,N_18984,N_18910);
or U19118 (N_19118,N_18953,N_18888);
nor U19119 (N_19119,N_18928,N_18918);
and U19120 (N_19120,N_18924,N_18901);
nor U19121 (N_19121,N_18827,N_18918);
nand U19122 (N_19122,N_18852,N_18828);
or U19123 (N_19123,N_18883,N_18859);
nor U19124 (N_19124,N_18956,N_18985);
nand U19125 (N_19125,N_18868,N_18826);
xor U19126 (N_19126,N_18992,N_18848);
nor U19127 (N_19127,N_18931,N_18880);
or U19128 (N_19128,N_18910,N_18860);
xnor U19129 (N_19129,N_18922,N_18966);
or U19130 (N_19130,N_18935,N_18878);
xor U19131 (N_19131,N_18824,N_18844);
xor U19132 (N_19132,N_18883,N_18984);
and U19133 (N_19133,N_18800,N_18804);
xnor U19134 (N_19134,N_18977,N_18914);
xnor U19135 (N_19135,N_18804,N_18933);
xor U19136 (N_19136,N_18967,N_18816);
nor U19137 (N_19137,N_18871,N_18919);
or U19138 (N_19138,N_18943,N_18952);
nand U19139 (N_19139,N_18862,N_18816);
and U19140 (N_19140,N_18945,N_18897);
nor U19141 (N_19141,N_18918,N_18980);
nand U19142 (N_19142,N_18959,N_18871);
or U19143 (N_19143,N_18885,N_18838);
and U19144 (N_19144,N_18906,N_18886);
xnor U19145 (N_19145,N_18821,N_18804);
nor U19146 (N_19146,N_18882,N_18805);
nand U19147 (N_19147,N_18931,N_18825);
and U19148 (N_19148,N_18901,N_18963);
nor U19149 (N_19149,N_18847,N_18899);
nor U19150 (N_19150,N_18967,N_18980);
or U19151 (N_19151,N_18998,N_18990);
nand U19152 (N_19152,N_18854,N_18979);
or U19153 (N_19153,N_18886,N_18956);
nor U19154 (N_19154,N_18835,N_18908);
nand U19155 (N_19155,N_18962,N_18996);
or U19156 (N_19156,N_18946,N_18836);
or U19157 (N_19157,N_18936,N_18951);
nor U19158 (N_19158,N_18903,N_18937);
or U19159 (N_19159,N_18802,N_18973);
or U19160 (N_19160,N_18871,N_18888);
nand U19161 (N_19161,N_18828,N_18875);
nor U19162 (N_19162,N_18901,N_18914);
xor U19163 (N_19163,N_18954,N_18947);
nand U19164 (N_19164,N_18937,N_18929);
and U19165 (N_19165,N_18997,N_18993);
nand U19166 (N_19166,N_18910,N_18838);
and U19167 (N_19167,N_18912,N_18927);
xor U19168 (N_19168,N_18890,N_18948);
nand U19169 (N_19169,N_18871,N_18978);
and U19170 (N_19170,N_18831,N_18884);
and U19171 (N_19171,N_18924,N_18880);
xor U19172 (N_19172,N_18963,N_18913);
or U19173 (N_19173,N_18826,N_18917);
xor U19174 (N_19174,N_18870,N_18954);
or U19175 (N_19175,N_18830,N_18863);
or U19176 (N_19176,N_18955,N_18972);
or U19177 (N_19177,N_18851,N_18815);
nand U19178 (N_19178,N_18888,N_18975);
xnor U19179 (N_19179,N_18826,N_18878);
and U19180 (N_19180,N_18901,N_18909);
xnor U19181 (N_19181,N_18905,N_18884);
xor U19182 (N_19182,N_18945,N_18900);
xor U19183 (N_19183,N_18935,N_18828);
or U19184 (N_19184,N_18900,N_18943);
nor U19185 (N_19185,N_18827,N_18982);
and U19186 (N_19186,N_18830,N_18818);
and U19187 (N_19187,N_18815,N_18856);
or U19188 (N_19188,N_18945,N_18986);
xnor U19189 (N_19189,N_18992,N_18987);
nor U19190 (N_19190,N_18817,N_18966);
xnor U19191 (N_19191,N_18958,N_18901);
xnor U19192 (N_19192,N_18803,N_18859);
xor U19193 (N_19193,N_18914,N_18858);
nand U19194 (N_19194,N_18947,N_18918);
xnor U19195 (N_19195,N_18900,N_18982);
or U19196 (N_19196,N_18934,N_18979);
nand U19197 (N_19197,N_18959,N_18880);
nand U19198 (N_19198,N_18900,N_18942);
nand U19199 (N_19199,N_18926,N_18829);
nand U19200 (N_19200,N_19128,N_19010);
nand U19201 (N_19201,N_19021,N_19170);
nor U19202 (N_19202,N_19012,N_19095);
and U19203 (N_19203,N_19055,N_19193);
xor U19204 (N_19204,N_19109,N_19098);
nor U19205 (N_19205,N_19062,N_19103);
xnor U19206 (N_19206,N_19172,N_19023);
and U19207 (N_19207,N_19184,N_19153);
nand U19208 (N_19208,N_19087,N_19118);
nor U19209 (N_19209,N_19187,N_19086);
or U19210 (N_19210,N_19112,N_19052);
nor U19211 (N_19211,N_19132,N_19093);
and U19212 (N_19212,N_19158,N_19114);
or U19213 (N_19213,N_19143,N_19129);
nand U19214 (N_19214,N_19006,N_19159);
nand U19215 (N_19215,N_19022,N_19008);
or U19216 (N_19216,N_19091,N_19066);
or U19217 (N_19217,N_19189,N_19175);
or U19218 (N_19218,N_19041,N_19191);
nand U19219 (N_19219,N_19038,N_19043);
nor U19220 (N_19220,N_19176,N_19009);
xor U19221 (N_19221,N_19037,N_19157);
nand U19222 (N_19222,N_19099,N_19156);
xor U19223 (N_19223,N_19131,N_19192);
nand U19224 (N_19224,N_19130,N_19011);
nand U19225 (N_19225,N_19155,N_19137);
xor U19226 (N_19226,N_19180,N_19127);
nand U19227 (N_19227,N_19135,N_19019);
nand U19228 (N_19228,N_19122,N_19162);
or U19229 (N_19229,N_19015,N_19173);
or U19230 (N_19230,N_19164,N_19097);
and U19231 (N_19231,N_19003,N_19120);
nor U19232 (N_19232,N_19057,N_19072);
or U19233 (N_19233,N_19074,N_19005);
nor U19234 (N_19234,N_19088,N_19029);
nor U19235 (N_19235,N_19194,N_19160);
nor U19236 (N_19236,N_19061,N_19040);
xnor U19237 (N_19237,N_19167,N_19145);
nand U19238 (N_19238,N_19059,N_19136);
nand U19239 (N_19239,N_19096,N_19007);
nand U19240 (N_19240,N_19016,N_19105);
and U19241 (N_19241,N_19020,N_19169);
nor U19242 (N_19242,N_19035,N_19177);
or U19243 (N_19243,N_19102,N_19094);
nand U19244 (N_19244,N_19108,N_19048);
nor U19245 (N_19245,N_19090,N_19163);
xnor U19246 (N_19246,N_19196,N_19183);
and U19247 (N_19247,N_19116,N_19150);
xor U19248 (N_19248,N_19190,N_19085);
nand U19249 (N_19249,N_19078,N_19113);
xor U19250 (N_19250,N_19199,N_19034);
or U19251 (N_19251,N_19028,N_19161);
or U19252 (N_19252,N_19068,N_19147);
or U19253 (N_19253,N_19146,N_19031);
nand U19254 (N_19254,N_19138,N_19179);
nand U19255 (N_19255,N_19053,N_19125);
nor U19256 (N_19256,N_19018,N_19151);
or U19257 (N_19257,N_19171,N_19198);
and U19258 (N_19258,N_19082,N_19002);
nor U19259 (N_19259,N_19026,N_19104);
nand U19260 (N_19260,N_19111,N_19077);
xor U19261 (N_19261,N_19185,N_19107);
or U19262 (N_19262,N_19106,N_19092);
and U19263 (N_19263,N_19030,N_19154);
nor U19264 (N_19264,N_19166,N_19124);
xnor U19265 (N_19265,N_19110,N_19168);
nand U19266 (N_19266,N_19083,N_19134);
or U19267 (N_19267,N_19042,N_19064);
xor U19268 (N_19268,N_19050,N_19032);
nand U19269 (N_19269,N_19119,N_19075);
nor U19270 (N_19270,N_19186,N_19081);
and U19271 (N_19271,N_19047,N_19045);
nor U19272 (N_19272,N_19080,N_19181);
and U19273 (N_19273,N_19148,N_19056);
or U19274 (N_19274,N_19060,N_19025);
nor U19275 (N_19275,N_19063,N_19142);
xor U19276 (N_19276,N_19065,N_19079);
xor U19277 (N_19277,N_19000,N_19049);
or U19278 (N_19278,N_19004,N_19076);
xor U19279 (N_19279,N_19140,N_19036);
nor U19280 (N_19280,N_19117,N_19144);
nor U19281 (N_19281,N_19149,N_19044);
or U19282 (N_19282,N_19195,N_19188);
nor U19283 (N_19283,N_19197,N_19070);
nand U19284 (N_19284,N_19014,N_19141);
or U19285 (N_19285,N_19121,N_19027);
and U19286 (N_19286,N_19046,N_19174);
or U19287 (N_19287,N_19017,N_19033);
or U19288 (N_19288,N_19100,N_19139);
xor U19289 (N_19289,N_19133,N_19039);
nand U19290 (N_19290,N_19182,N_19024);
xnor U19291 (N_19291,N_19101,N_19178);
and U19292 (N_19292,N_19058,N_19054);
nand U19293 (N_19293,N_19084,N_19067);
xnor U19294 (N_19294,N_19152,N_19165);
and U19295 (N_19295,N_19126,N_19051);
nor U19296 (N_19296,N_19071,N_19123);
and U19297 (N_19297,N_19013,N_19089);
xnor U19298 (N_19298,N_19001,N_19069);
nand U19299 (N_19299,N_19115,N_19073);
or U19300 (N_19300,N_19049,N_19078);
nor U19301 (N_19301,N_19066,N_19138);
nand U19302 (N_19302,N_19088,N_19021);
nor U19303 (N_19303,N_19153,N_19138);
or U19304 (N_19304,N_19006,N_19047);
or U19305 (N_19305,N_19004,N_19001);
nand U19306 (N_19306,N_19122,N_19012);
and U19307 (N_19307,N_19089,N_19134);
and U19308 (N_19308,N_19120,N_19004);
and U19309 (N_19309,N_19015,N_19141);
xor U19310 (N_19310,N_19149,N_19075);
nand U19311 (N_19311,N_19150,N_19076);
or U19312 (N_19312,N_19141,N_19074);
and U19313 (N_19313,N_19133,N_19104);
xor U19314 (N_19314,N_19017,N_19148);
and U19315 (N_19315,N_19152,N_19168);
and U19316 (N_19316,N_19124,N_19061);
and U19317 (N_19317,N_19006,N_19090);
or U19318 (N_19318,N_19064,N_19023);
nor U19319 (N_19319,N_19090,N_19013);
or U19320 (N_19320,N_19066,N_19163);
nor U19321 (N_19321,N_19098,N_19074);
or U19322 (N_19322,N_19133,N_19125);
and U19323 (N_19323,N_19140,N_19155);
nor U19324 (N_19324,N_19097,N_19196);
or U19325 (N_19325,N_19022,N_19090);
nand U19326 (N_19326,N_19155,N_19003);
nor U19327 (N_19327,N_19058,N_19108);
and U19328 (N_19328,N_19172,N_19179);
or U19329 (N_19329,N_19137,N_19104);
xor U19330 (N_19330,N_19054,N_19047);
or U19331 (N_19331,N_19197,N_19163);
xor U19332 (N_19332,N_19161,N_19059);
and U19333 (N_19333,N_19069,N_19152);
nand U19334 (N_19334,N_19083,N_19161);
xnor U19335 (N_19335,N_19041,N_19198);
nand U19336 (N_19336,N_19108,N_19172);
xnor U19337 (N_19337,N_19105,N_19195);
nand U19338 (N_19338,N_19024,N_19084);
xnor U19339 (N_19339,N_19138,N_19096);
nor U19340 (N_19340,N_19025,N_19134);
xor U19341 (N_19341,N_19065,N_19177);
nor U19342 (N_19342,N_19175,N_19050);
or U19343 (N_19343,N_19072,N_19149);
nand U19344 (N_19344,N_19156,N_19163);
nor U19345 (N_19345,N_19036,N_19034);
or U19346 (N_19346,N_19077,N_19130);
or U19347 (N_19347,N_19064,N_19053);
nand U19348 (N_19348,N_19056,N_19187);
nand U19349 (N_19349,N_19188,N_19006);
or U19350 (N_19350,N_19004,N_19089);
xnor U19351 (N_19351,N_19180,N_19177);
nor U19352 (N_19352,N_19056,N_19150);
or U19353 (N_19353,N_19085,N_19142);
or U19354 (N_19354,N_19142,N_19198);
nor U19355 (N_19355,N_19089,N_19033);
nand U19356 (N_19356,N_19094,N_19158);
or U19357 (N_19357,N_19152,N_19117);
and U19358 (N_19358,N_19093,N_19094);
nand U19359 (N_19359,N_19133,N_19170);
and U19360 (N_19360,N_19027,N_19082);
or U19361 (N_19361,N_19043,N_19031);
and U19362 (N_19362,N_19077,N_19087);
and U19363 (N_19363,N_19002,N_19083);
nor U19364 (N_19364,N_19125,N_19144);
or U19365 (N_19365,N_19167,N_19035);
or U19366 (N_19366,N_19037,N_19140);
nor U19367 (N_19367,N_19077,N_19058);
xor U19368 (N_19368,N_19011,N_19119);
xnor U19369 (N_19369,N_19088,N_19026);
nand U19370 (N_19370,N_19038,N_19152);
nor U19371 (N_19371,N_19056,N_19110);
nand U19372 (N_19372,N_19186,N_19120);
and U19373 (N_19373,N_19049,N_19134);
nand U19374 (N_19374,N_19009,N_19061);
nor U19375 (N_19375,N_19189,N_19065);
and U19376 (N_19376,N_19174,N_19102);
xnor U19377 (N_19377,N_19022,N_19137);
xnor U19378 (N_19378,N_19144,N_19080);
xnor U19379 (N_19379,N_19077,N_19107);
xnor U19380 (N_19380,N_19010,N_19171);
nor U19381 (N_19381,N_19035,N_19078);
and U19382 (N_19382,N_19004,N_19059);
nor U19383 (N_19383,N_19193,N_19063);
and U19384 (N_19384,N_19020,N_19129);
nand U19385 (N_19385,N_19001,N_19025);
xnor U19386 (N_19386,N_19126,N_19109);
xnor U19387 (N_19387,N_19027,N_19146);
nand U19388 (N_19388,N_19042,N_19182);
or U19389 (N_19389,N_19110,N_19066);
nor U19390 (N_19390,N_19118,N_19145);
and U19391 (N_19391,N_19157,N_19185);
nor U19392 (N_19392,N_19045,N_19050);
or U19393 (N_19393,N_19029,N_19092);
xor U19394 (N_19394,N_19034,N_19085);
and U19395 (N_19395,N_19006,N_19087);
or U19396 (N_19396,N_19035,N_19147);
or U19397 (N_19397,N_19191,N_19025);
xnor U19398 (N_19398,N_19162,N_19031);
xnor U19399 (N_19399,N_19094,N_19031);
nor U19400 (N_19400,N_19371,N_19306);
nor U19401 (N_19401,N_19236,N_19329);
nand U19402 (N_19402,N_19388,N_19394);
and U19403 (N_19403,N_19339,N_19311);
nand U19404 (N_19404,N_19301,N_19319);
nand U19405 (N_19405,N_19354,N_19205);
xor U19406 (N_19406,N_19234,N_19286);
xor U19407 (N_19407,N_19359,N_19328);
xnor U19408 (N_19408,N_19245,N_19362);
nand U19409 (N_19409,N_19357,N_19368);
xnor U19410 (N_19410,N_19338,N_19295);
and U19411 (N_19411,N_19299,N_19211);
or U19412 (N_19412,N_19298,N_19314);
xor U19413 (N_19413,N_19335,N_19214);
nand U19414 (N_19414,N_19209,N_19223);
or U19415 (N_19415,N_19316,N_19349);
nand U19416 (N_19416,N_19248,N_19230);
nor U19417 (N_19417,N_19274,N_19386);
nor U19418 (N_19418,N_19256,N_19264);
and U19419 (N_19419,N_19337,N_19383);
nor U19420 (N_19420,N_19332,N_19333);
nor U19421 (N_19421,N_19285,N_19372);
nor U19422 (N_19422,N_19389,N_19290);
nand U19423 (N_19423,N_19215,N_19302);
xnor U19424 (N_19424,N_19224,N_19217);
nor U19425 (N_19425,N_19346,N_19387);
and U19426 (N_19426,N_19255,N_19397);
xnor U19427 (N_19427,N_19208,N_19304);
and U19428 (N_19428,N_19206,N_19212);
nor U19429 (N_19429,N_19326,N_19262);
nand U19430 (N_19430,N_19296,N_19327);
nand U19431 (N_19431,N_19219,N_19272);
nor U19432 (N_19432,N_19345,N_19266);
nand U19433 (N_19433,N_19292,N_19373);
nand U19434 (N_19434,N_19287,N_19228);
nand U19435 (N_19435,N_19231,N_19277);
nand U19436 (N_19436,N_19369,N_19251);
nand U19437 (N_19437,N_19376,N_19378);
nand U19438 (N_19438,N_19269,N_19293);
nor U19439 (N_19439,N_19375,N_19233);
nand U19440 (N_19440,N_19237,N_19379);
xnor U19441 (N_19441,N_19343,N_19320);
xnor U19442 (N_19442,N_19324,N_19267);
nor U19443 (N_19443,N_19330,N_19384);
nor U19444 (N_19444,N_19307,N_19281);
or U19445 (N_19445,N_19351,N_19280);
nand U19446 (N_19446,N_19263,N_19395);
or U19447 (N_19447,N_19225,N_19352);
or U19448 (N_19448,N_19200,N_19348);
nor U19449 (N_19449,N_19322,N_19385);
xor U19450 (N_19450,N_19270,N_19350);
and U19451 (N_19451,N_19291,N_19318);
or U19452 (N_19452,N_19391,N_19241);
xor U19453 (N_19453,N_19271,N_19294);
nor U19454 (N_19454,N_19252,N_19315);
or U19455 (N_19455,N_19258,N_19377);
nand U19456 (N_19456,N_19275,N_19398);
and U19457 (N_19457,N_19365,N_19268);
xnor U19458 (N_19458,N_19232,N_19355);
xor U19459 (N_19459,N_19222,N_19207);
xnor U19460 (N_19460,N_19229,N_19247);
or U19461 (N_19461,N_19312,N_19273);
and U19462 (N_19462,N_19308,N_19278);
and U19463 (N_19463,N_19334,N_19238);
xor U19464 (N_19464,N_19390,N_19218);
nand U19465 (N_19465,N_19243,N_19261);
xor U19466 (N_19466,N_19344,N_19340);
or U19467 (N_19467,N_19249,N_19204);
xor U19468 (N_19468,N_19265,N_19380);
or U19469 (N_19469,N_19347,N_19367);
nand U19470 (N_19470,N_19393,N_19254);
and U19471 (N_19471,N_19313,N_19288);
nand U19472 (N_19472,N_19227,N_19250);
or U19473 (N_19473,N_19360,N_19399);
or U19474 (N_19474,N_19221,N_19374);
and U19475 (N_19475,N_19216,N_19244);
nor U19476 (N_19476,N_19364,N_19257);
nand U19477 (N_19477,N_19382,N_19203);
and U19478 (N_19478,N_19310,N_19303);
or U19479 (N_19479,N_19240,N_19392);
nand U19480 (N_19480,N_19279,N_19226);
or U19481 (N_19481,N_19321,N_19297);
nand U19482 (N_19482,N_19220,N_19305);
nor U19483 (N_19483,N_19396,N_19342);
nor U19484 (N_19484,N_19300,N_19370);
nor U19485 (N_19485,N_19260,N_19358);
nand U19486 (N_19486,N_19284,N_19202);
nor U19487 (N_19487,N_19289,N_19246);
xnor U19488 (N_19488,N_19235,N_19213);
nand U19489 (N_19489,N_19282,N_19210);
nor U19490 (N_19490,N_19253,N_19201);
nor U19491 (N_19491,N_19361,N_19363);
or U19492 (N_19492,N_19323,N_19331);
xnor U19493 (N_19493,N_19309,N_19276);
or U19494 (N_19494,N_19381,N_19325);
or U19495 (N_19495,N_19317,N_19366);
nor U19496 (N_19496,N_19242,N_19283);
or U19497 (N_19497,N_19259,N_19239);
nand U19498 (N_19498,N_19353,N_19356);
nor U19499 (N_19499,N_19341,N_19336);
xnor U19500 (N_19500,N_19259,N_19361);
and U19501 (N_19501,N_19364,N_19323);
nor U19502 (N_19502,N_19253,N_19268);
and U19503 (N_19503,N_19226,N_19356);
nand U19504 (N_19504,N_19313,N_19291);
nand U19505 (N_19505,N_19261,N_19277);
xor U19506 (N_19506,N_19210,N_19243);
xor U19507 (N_19507,N_19359,N_19234);
or U19508 (N_19508,N_19257,N_19390);
xor U19509 (N_19509,N_19246,N_19296);
nand U19510 (N_19510,N_19360,N_19342);
and U19511 (N_19511,N_19311,N_19285);
and U19512 (N_19512,N_19325,N_19326);
nand U19513 (N_19513,N_19219,N_19368);
or U19514 (N_19514,N_19378,N_19341);
nand U19515 (N_19515,N_19258,N_19348);
nor U19516 (N_19516,N_19290,N_19223);
nand U19517 (N_19517,N_19266,N_19349);
and U19518 (N_19518,N_19351,N_19369);
xnor U19519 (N_19519,N_19365,N_19232);
or U19520 (N_19520,N_19277,N_19221);
and U19521 (N_19521,N_19374,N_19282);
nor U19522 (N_19522,N_19336,N_19330);
and U19523 (N_19523,N_19260,N_19306);
nand U19524 (N_19524,N_19333,N_19308);
and U19525 (N_19525,N_19344,N_19375);
or U19526 (N_19526,N_19239,N_19233);
and U19527 (N_19527,N_19264,N_19248);
or U19528 (N_19528,N_19278,N_19271);
nand U19529 (N_19529,N_19359,N_19308);
nor U19530 (N_19530,N_19249,N_19382);
and U19531 (N_19531,N_19298,N_19277);
and U19532 (N_19532,N_19267,N_19209);
and U19533 (N_19533,N_19319,N_19220);
nand U19534 (N_19534,N_19337,N_19330);
nor U19535 (N_19535,N_19244,N_19274);
or U19536 (N_19536,N_19323,N_19259);
nor U19537 (N_19537,N_19385,N_19365);
nor U19538 (N_19538,N_19237,N_19332);
nand U19539 (N_19539,N_19294,N_19355);
or U19540 (N_19540,N_19310,N_19316);
nor U19541 (N_19541,N_19393,N_19326);
or U19542 (N_19542,N_19250,N_19273);
nor U19543 (N_19543,N_19254,N_19387);
xor U19544 (N_19544,N_19294,N_19221);
or U19545 (N_19545,N_19273,N_19223);
xnor U19546 (N_19546,N_19371,N_19277);
and U19547 (N_19547,N_19378,N_19269);
xor U19548 (N_19548,N_19226,N_19233);
or U19549 (N_19549,N_19339,N_19371);
and U19550 (N_19550,N_19345,N_19391);
nor U19551 (N_19551,N_19273,N_19325);
xnor U19552 (N_19552,N_19357,N_19274);
nor U19553 (N_19553,N_19276,N_19326);
and U19554 (N_19554,N_19244,N_19202);
and U19555 (N_19555,N_19248,N_19357);
or U19556 (N_19556,N_19304,N_19291);
and U19557 (N_19557,N_19364,N_19366);
or U19558 (N_19558,N_19375,N_19299);
nor U19559 (N_19559,N_19244,N_19386);
xnor U19560 (N_19560,N_19345,N_19245);
xnor U19561 (N_19561,N_19388,N_19398);
xor U19562 (N_19562,N_19259,N_19317);
nor U19563 (N_19563,N_19283,N_19245);
or U19564 (N_19564,N_19390,N_19369);
and U19565 (N_19565,N_19296,N_19201);
and U19566 (N_19566,N_19353,N_19329);
xor U19567 (N_19567,N_19237,N_19206);
xnor U19568 (N_19568,N_19325,N_19231);
and U19569 (N_19569,N_19258,N_19252);
and U19570 (N_19570,N_19341,N_19316);
xor U19571 (N_19571,N_19283,N_19359);
and U19572 (N_19572,N_19221,N_19309);
and U19573 (N_19573,N_19220,N_19217);
or U19574 (N_19574,N_19232,N_19364);
and U19575 (N_19575,N_19263,N_19232);
or U19576 (N_19576,N_19379,N_19331);
xor U19577 (N_19577,N_19295,N_19307);
nand U19578 (N_19578,N_19391,N_19268);
or U19579 (N_19579,N_19294,N_19370);
or U19580 (N_19580,N_19369,N_19360);
nor U19581 (N_19581,N_19387,N_19242);
and U19582 (N_19582,N_19362,N_19249);
nand U19583 (N_19583,N_19361,N_19282);
nor U19584 (N_19584,N_19309,N_19361);
and U19585 (N_19585,N_19373,N_19243);
nand U19586 (N_19586,N_19296,N_19289);
xor U19587 (N_19587,N_19264,N_19314);
and U19588 (N_19588,N_19273,N_19210);
nor U19589 (N_19589,N_19242,N_19316);
nor U19590 (N_19590,N_19253,N_19261);
nand U19591 (N_19591,N_19259,N_19284);
nand U19592 (N_19592,N_19266,N_19245);
nor U19593 (N_19593,N_19318,N_19287);
or U19594 (N_19594,N_19219,N_19335);
or U19595 (N_19595,N_19289,N_19388);
nand U19596 (N_19596,N_19378,N_19301);
nor U19597 (N_19597,N_19241,N_19342);
nor U19598 (N_19598,N_19365,N_19294);
or U19599 (N_19599,N_19207,N_19277);
or U19600 (N_19600,N_19499,N_19475);
nand U19601 (N_19601,N_19407,N_19543);
nor U19602 (N_19602,N_19590,N_19422);
and U19603 (N_19603,N_19466,N_19402);
nor U19604 (N_19604,N_19593,N_19498);
xnor U19605 (N_19605,N_19572,N_19566);
or U19606 (N_19606,N_19589,N_19536);
and U19607 (N_19607,N_19519,N_19439);
or U19608 (N_19608,N_19477,N_19530);
nand U19609 (N_19609,N_19487,N_19413);
and U19610 (N_19610,N_19552,N_19493);
nor U19611 (N_19611,N_19534,N_19599);
nand U19612 (N_19612,N_19521,N_19411);
and U19613 (N_19613,N_19503,N_19541);
xnor U19614 (N_19614,N_19406,N_19482);
and U19615 (N_19615,N_19443,N_19551);
nand U19616 (N_19616,N_19502,N_19400);
or U19617 (N_19617,N_19433,N_19462);
or U19618 (N_19618,N_19456,N_19403);
nand U19619 (N_19619,N_19457,N_19579);
xnor U19620 (N_19620,N_19404,N_19538);
nor U19621 (N_19621,N_19588,N_19467);
nand U19622 (N_19622,N_19416,N_19461);
or U19623 (N_19623,N_19414,N_19597);
xor U19624 (N_19624,N_19516,N_19561);
or U19625 (N_19625,N_19472,N_19442);
nor U19626 (N_19626,N_19495,N_19594);
and U19627 (N_19627,N_19524,N_19426);
nand U19628 (N_19628,N_19424,N_19483);
nor U19629 (N_19629,N_19558,N_19592);
nor U19630 (N_19630,N_19522,N_19546);
nand U19631 (N_19631,N_19533,N_19408);
nor U19632 (N_19632,N_19469,N_19515);
and U19633 (N_19633,N_19528,N_19435);
nor U19634 (N_19634,N_19582,N_19506);
xor U19635 (N_19635,N_19480,N_19527);
and U19636 (N_19636,N_19450,N_19556);
and U19637 (N_19637,N_19434,N_19553);
xor U19638 (N_19638,N_19577,N_19501);
xor U19639 (N_19639,N_19517,N_19571);
or U19640 (N_19640,N_19465,N_19481);
or U19641 (N_19641,N_19446,N_19464);
nor U19642 (N_19642,N_19419,N_19580);
or U19643 (N_19643,N_19401,N_19478);
nor U19644 (N_19644,N_19468,N_19532);
nor U19645 (N_19645,N_19567,N_19454);
and U19646 (N_19646,N_19578,N_19479);
nand U19647 (N_19647,N_19526,N_19451);
nor U19648 (N_19648,N_19427,N_19489);
nor U19649 (N_19649,N_19470,N_19586);
xor U19650 (N_19650,N_19412,N_19520);
or U19651 (N_19651,N_19473,N_19565);
xnor U19652 (N_19652,N_19448,N_19542);
nand U19653 (N_19653,N_19555,N_19485);
and U19654 (N_19654,N_19486,N_19511);
nor U19655 (N_19655,N_19494,N_19595);
and U19656 (N_19656,N_19507,N_19425);
and U19657 (N_19657,N_19510,N_19539);
and U19658 (N_19658,N_19497,N_19490);
nor U19659 (N_19659,N_19428,N_19509);
xor U19660 (N_19660,N_19548,N_19460);
or U19661 (N_19661,N_19458,N_19569);
xnor U19662 (N_19662,N_19437,N_19444);
nor U19663 (N_19663,N_19423,N_19484);
xor U19664 (N_19664,N_19417,N_19544);
nor U19665 (N_19665,N_19488,N_19508);
or U19666 (N_19666,N_19449,N_19540);
nand U19667 (N_19667,N_19547,N_19550);
or U19668 (N_19668,N_19575,N_19574);
and U19669 (N_19669,N_19459,N_19410);
nand U19670 (N_19670,N_19584,N_19554);
xnor U19671 (N_19671,N_19440,N_19549);
and U19672 (N_19672,N_19409,N_19491);
xnor U19673 (N_19673,N_19523,N_19441);
nand U19674 (N_19674,N_19476,N_19518);
or U19675 (N_19675,N_19525,N_19474);
nor U19676 (N_19676,N_19537,N_19447);
and U19677 (N_19677,N_19418,N_19581);
nor U19678 (N_19678,N_19405,N_19557);
nor U19679 (N_19679,N_19452,N_19585);
nor U19680 (N_19680,N_19564,N_19562);
xor U19681 (N_19681,N_19492,N_19570);
xor U19682 (N_19682,N_19587,N_19471);
nor U19683 (N_19683,N_19563,N_19568);
nand U19684 (N_19684,N_19415,N_19430);
nor U19685 (N_19685,N_19512,N_19591);
or U19686 (N_19686,N_19531,N_19529);
xnor U19687 (N_19687,N_19500,N_19598);
nor U19688 (N_19688,N_19513,N_19504);
and U19689 (N_19689,N_19438,N_19496);
or U19690 (N_19690,N_19429,N_19445);
or U19691 (N_19691,N_19559,N_19431);
and U19692 (N_19692,N_19455,N_19463);
or U19693 (N_19693,N_19583,N_19420);
nand U19694 (N_19694,N_19432,N_19505);
xnor U19695 (N_19695,N_19514,N_19545);
and U19696 (N_19696,N_19573,N_19453);
nand U19697 (N_19697,N_19596,N_19421);
xor U19698 (N_19698,N_19560,N_19576);
and U19699 (N_19699,N_19436,N_19535);
nor U19700 (N_19700,N_19562,N_19535);
nand U19701 (N_19701,N_19458,N_19553);
nand U19702 (N_19702,N_19400,N_19434);
or U19703 (N_19703,N_19572,N_19587);
or U19704 (N_19704,N_19540,N_19451);
xor U19705 (N_19705,N_19530,N_19550);
or U19706 (N_19706,N_19503,N_19573);
nor U19707 (N_19707,N_19562,N_19538);
nand U19708 (N_19708,N_19534,N_19504);
nor U19709 (N_19709,N_19547,N_19560);
or U19710 (N_19710,N_19522,N_19538);
nor U19711 (N_19711,N_19448,N_19526);
and U19712 (N_19712,N_19453,N_19595);
nor U19713 (N_19713,N_19413,N_19524);
nand U19714 (N_19714,N_19437,N_19532);
xnor U19715 (N_19715,N_19402,N_19516);
and U19716 (N_19716,N_19409,N_19418);
nand U19717 (N_19717,N_19497,N_19441);
xnor U19718 (N_19718,N_19566,N_19551);
or U19719 (N_19719,N_19550,N_19592);
or U19720 (N_19720,N_19546,N_19583);
nor U19721 (N_19721,N_19465,N_19408);
nand U19722 (N_19722,N_19472,N_19406);
nand U19723 (N_19723,N_19465,N_19447);
nor U19724 (N_19724,N_19439,N_19422);
nor U19725 (N_19725,N_19514,N_19473);
nor U19726 (N_19726,N_19591,N_19515);
nor U19727 (N_19727,N_19458,N_19452);
nand U19728 (N_19728,N_19417,N_19460);
or U19729 (N_19729,N_19448,N_19544);
nand U19730 (N_19730,N_19461,N_19441);
nand U19731 (N_19731,N_19556,N_19535);
nor U19732 (N_19732,N_19509,N_19598);
or U19733 (N_19733,N_19554,N_19561);
nand U19734 (N_19734,N_19566,N_19565);
nor U19735 (N_19735,N_19448,N_19484);
nor U19736 (N_19736,N_19454,N_19422);
or U19737 (N_19737,N_19524,N_19494);
nor U19738 (N_19738,N_19503,N_19557);
nand U19739 (N_19739,N_19500,N_19502);
and U19740 (N_19740,N_19567,N_19515);
nand U19741 (N_19741,N_19538,N_19561);
nor U19742 (N_19742,N_19463,N_19537);
nor U19743 (N_19743,N_19530,N_19446);
and U19744 (N_19744,N_19573,N_19431);
xor U19745 (N_19745,N_19496,N_19455);
and U19746 (N_19746,N_19542,N_19569);
nand U19747 (N_19747,N_19463,N_19559);
nand U19748 (N_19748,N_19550,N_19532);
and U19749 (N_19749,N_19555,N_19494);
nor U19750 (N_19750,N_19564,N_19486);
nor U19751 (N_19751,N_19407,N_19453);
nor U19752 (N_19752,N_19474,N_19451);
nand U19753 (N_19753,N_19595,N_19560);
or U19754 (N_19754,N_19529,N_19405);
xor U19755 (N_19755,N_19482,N_19452);
nand U19756 (N_19756,N_19438,N_19536);
nand U19757 (N_19757,N_19509,N_19533);
or U19758 (N_19758,N_19446,N_19562);
or U19759 (N_19759,N_19493,N_19417);
and U19760 (N_19760,N_19492,N_19591);
xnor U19761 (N_19761,N_19595,N_19552);
and U19762 (N_19762,N_19408,N_19515);
nand U19763 (N_19763,N_19437,N_19555);
and U19764 (N_19764,N_19417,N_19530);
nor U19765 (N_19765,N_19500,N_19450);
and U19766 (N_19766,N_19510,N_19472);
xor U19767 (N_19767,N_19424,N_19481);
nor U19768 (N_19768,N_19534,N_19408);
xnor U19769 (N_19769,N_19528,N_19448);
nor U19770 (N_19770,N_19400,N_19472);
nor U19771 (N_19771,N_19511,N_19422);
nor U19772 (N_19772,N_19529,N_19450);
nor U19773 (N_19773,N_19557,N_19515);
or U19774 (N_19774,N_19552,N_19456);
nand U19775 (N_19775,N_19550,N_19477);
nor U19776 (N_19776,N_19571,N_19516);
nand U19777 (N_19777,N_19499,N_19493);
nor U19778 (N_19778,N_19492,N_19456);
nor U19779 (N_19779,N_19451,N_19488);
xnor U19780 (N_19780,N_19471,N_19547);
and U19781 (N_19781,N_19575,N_19485);
xnor U19782 (N_19782,N_19410,N_19409);
xor U19783 (N_19783,N_19509,N_19530);
xnor U19784 (N_19784,N_19489,N_19514);
or U19785 (N_19785,N_19566,N_19550);
nand U19786 (N_19786,N_19476,N_19419);
and U19787 (N_19787,N_19466,N_19578);
xor U19788 (N_19788,N_19486,N_19463);
xnor U19789 (N_19789,N_19599,N_19581);
and U19790 (N_19790,N_19407,N_19521);
or U19791 (N_19791,N_19594,N_19591);
and U19792 (N_19792,N_19574,N_19591);
nor U19793 (N_19793,N_19480,N_19445);
xor U19794 (N_19794,N_19495,N_19496);
and U19795 (N_19795,N_19459,N_19496);
nor U19796 (N_19796,N_19559,N_19450);
nand U19797 (N_19797,N_19431,N_19486);
and U19798 (N_19798,N_19480,N_19458);
nand U19799 (N_19799,N_19427,N_19578);
xnor U19800 (N_19800,N_19610,N_19718);
nor U19801 (N_19801,N_19665,N_19742);
and U19802 (N_19802,N_19619,N_19673);
nand U19803 (N_19803,N_19615,N_19706);
xor U19804 (N_19804,N_19613,N_19627);
nor U19805 (N_19805,N_19605,N_19785);
and U19806 (N_19806,N_19780,N_19713);
or U19807 (N_19807,N_19683,N_19633);
and U19808 (N_19808,N_19716,N_19795);
xnor U19809 (N_19809,N_19638,N_19798);
xnor U19810 (N_19810,N_19679,N_19714);
nand U19811 (N_19811,N_19735,N_19702);
or U19812 (N_19812,N_19736,N_19697);
xnor U19813 (N_19813,N_19695,N_19779);
nand U19814 (N_19814,N_19681,N_19641);
xor U19815 (N_19815,N_19637,N_19773);
and U19816 (N_19816,N_19783,N_19643);
and U19817 (N_19817,N_19687,N_19626);
xnor U19818 (N_19818,N_19606,N_19634);
xor U19819 (N_19819,N_19651,N_19745);
or U19820 (N_19820,N_19793,N_19676);
nand U19821 (N_19821,N_19692,N_19758);
or U19822 (N_19822,N_19636,N_19760);
xor U19823 (N_19823,N_19655,N_19693);
nand U19824 (N_19824,N_19658,N_19631);
and U19825 (N_19825,N_19787,N_19649);
nand U19826 (N_19826,N_19734,N_19796);
nand U19827 (N_19827,N_19704,N_19729);
and U19828 (N_19828,N_19746,N_19756);
nor U19829 (N_19829,N_19703,N_19624);
nor U19830 (N_19830,N_19674,N_19726);
or U19831 (N_19831,N_19720,N_19685);
nor U19832 (N_19832,N_19646,N_19677);
nor U19833 (N_19833,N_19752,N_19622);
and U19834 (N_19834,N_19715,N_19740);
xor U19835 (N_19835,N_19712,N_19663);
and U19836 (N_19836,N_19753,N_19645);
xnor U19837 (N_19837,N_19733,N_19770);
xnor U19838 (N_19838,N_19721,N_19701);
or U19839 (N_19839,N_19680,N_19709);
nor U19840 (N_19840,N_19732,N_19600);
nor U19841 (N_19841,N_19608,N_19755);
nor U19842 (N_19842,N_19784,N_19777);
nor U19843 (N_19843,N_19710,N_19660);
and U19844 (N_19844,N_19616,N_19604);
nand U19845 (N_19845,N_19614,N_19696);
or U19846 (N_19846,N_19799,N_19654);
xnor U19847 (N_19847,N_19698,N_19738);
and U19848 (N_19848,N_19666,N_19632);
and U19849 (N_19849,N_19625,N_19764);
nor U19850 (N_19850,N_19700,N_19659);
nor U19851 (N_19851,N_19618,N_19761);
xnor U19852 (N_19852,N_19757,N_19776);
or U19853 (N_19853,N_19630,N_19617);
nor U19854 (N_19854,N_19717,N_19763);
nand U19855 (N_19855,N_19754,N_19648);
nor U19856 (N_19856,N_19688,N_19668);
nor U19857 (N_19857,N_19778,N_19724);
nand U19858 (N_19858,N_19731,N_19647);
nor U19859 (N_19859,N_19794,N_19728);
xnor U19860 (N_19860,N_19767,N_19684);
nor U19861 (N_19861,N_19682,N_19743);
nand U19862 (N_19862,N_19708,N_19744);
or U19863 (N_19863,N_19772,N_19750);
or U19864 (N_19864,N_19781,N_19797);
or U19865 (N_19865,N_19749,N_19629);
and U19866 (N_19866,N_19690,N_19694);
nor U19867 (N_19867,N_19628,N_19769);
xnor U19868 (N_19868,N_19789,N_19672);
xnor U19869 (N_19869,N_19727,N_19691);
and U19870 (N_19870,N_19730,N_19669);
nand U19871 (N_19871,N_19768,N_19705);
and U19872 (N_19872,N_19656,N_19601);
nand U19873 (N_19873,N_19671,N_19748);
xnor U19874 (N_19874,N_19675,N_19782);
xor U19875 (N_19875,N_19774,N_19602);
and U19876 (N_19876,N_19739,N_19612);
and U19877 (N_19877,N_19786,N_19689);
and U19878 (N_19878,N_19640,N_19707);
xor U19879 (N_19879,N_19667,N_19652);
xor U19880 (N_19880,N_19722,N_19771);
xor U19881 (N_19881,N_19661,N_19642);
nor U19882 (N_19882,N_19644,N_19788);
and U19883 (N_19883,N_19611,N_19623);
or U19884 (N_19884,N_19686,N_19603);
and U19885 (N_19885,N_19741,N_19699);
and U19886 (N_19886,N_19635,N_19621);
nand U19887 (N_19887,N_19751,N_19670);
and U19888 (N_19888,N_19653,N_19723);
nor U19889 (N_19889,N_19792,N_19678);
nor U19890 (N_19890,N_19747,N_19775);
xnor U19891 (N_19891,N_19664,N_19607);
or U19892 (N_19892,N_19759,N_19609);
xor U19893 (N_19893,N_19662,N_19711);
xnor U19894 (N_19894,N_19762,N_19765);
nand U19895 (N_19895,N_19620,N_19639);
or U19896 (N_19896,N_19737,N_19791);
nand U19897 (N_19897,N_19766,N_19725);
or U19898 (N_19898,N_19719,N_19650);
xnor U19899 (N_19899,N_19790,N_19657);
and U19900 (N_19900,N_19734,N_19772);
nand U19901 (N_19901,N_19688,N_19653);
nand U19902 (N_19902,N_19697,N_19677);
nand U19903 (N_19903,N_19702,N_19773);
xor U19904 (N_19904,N_19639,N_19714);
nor U19905 (N_19905,N_19626,N_19709);
nand U19906 (N_19906,N_19671,N_19781);
nor U19907 (N_19907,N_19799,N_19764);
nor U19908 (N_19908,N_19626,N_19618);
nand U19909 (N_19909,N_19701,N_19623);
xnor U19910 (N_19910,N_19708,N_19686);
nand U19911 (N_19911,N_19669,N_19614);
nor U19912 (N_19912,N_19634,N_19747);
xnor U19913 (N_19913,N_19651,N_19609);
xor U19914 (N_19914,N_19753,N_19788);
and U19915 (N_19915,N_19751,N_19649);
nor U19916 (N_19916,N_19706,N_19744);
and U19917 (N_19917,N_19610,N_19749);
and U19918 (N_19918,N_19649,N_19718);
nor U19919 (N_19919,N_19660,N_19777);
nor U19920 (N_19920,N_19684,N_19679);
nor U19921 (N_19921,N_19657,N_19632);
or U19922 (N_19922,N_19675,N_19790);
nand U19923 (N_19923,N_19715,N_19699);
nor U19924 (N_19924,N_19697,N_19699);
or U19925 (N_19925,N_19756,N_19691);
nand U19926 (N_19926,N_19709,N_19657);
xnor U19927 (N_19927,N_19676,N_19742);
or U19928 (N_19928,N_19606,N_19747);
and U19929 (N_19929,N_19792,N_19762);
nand U19930 (N_19930,N_19710,N_19618);
xor U19931 (N_19931,N_19662,N_19685);
nand U19932 (N_19932,N_19627,N_19672);
nor U19933 (N_19933,N_19742,N_19764);
xnor U19934 (N_19934,N_19783,N_19722);
nand U19935 (N_19935,N_19744,N_19643);
and U19936 (N_19936,N_19718,N_19730);
nor U19937 (N_19937,N_19721,N_19709);
xor U19938 (N_19938,N_19727,N_19639);
nor U19939 (N_19939,N_19738,N_19661);
and U19940 (N_19940,N_19642,N_19613);
nor U19941 (N_19941,N_19772,N_19616);
nor U19942 (N_19942,N_19619,N_19646);
nand U19943 (N_19943,N_19787,N_19738);
or U19944 (N_19944,N_19709,N_19649);
or U19945 (N_19945,N_19630,N_19631);
nand U19946 (N_19946,N_19640,N_19651);
xnor U19947 (N_19947,N_19773,N_19618);
or U19948 (N_19948,N_19729,N_19718);
xnor U19949 (N_19949,N_19679,N_19618);
and U19950 (N_19950,N_19712,N_19612);
or U19951 (N_19951,N_19715,N_19687);
xor U19952 (N_19952,N_19785,N_19771);
nor U19953 (N_19953,N_19665,N_19694);
and U19954 (N_19954,N_19725,N_19741);
xor U19955 (N_19955,N_19674,N_19725);
nand U19956 (N_19956,N_19751,N_19730);
xor U19957 (N_19957,N_19714,N_19629);
nor U19958 (N_19958,N_19785,N_19630);
nor U19959 (N_19959,N_19741,N_19614);
nand U19960 (N_19960,N_19615,N_19713);
nor U19961 (N_19961,N_19638,N_19768);
nand U19962 (N_19962,N_19668,N_19626);
or U19963 (N_19963,N_19612,N_19741);
xor U19964 (N_19964,N_19658,N_19610);
or U19965 (N_19965,N_19633,N_19722);
or U19966 (N_19966,N_19699,N_19683);
xor U19967 (N_19967,N_19763,N_19637);
and U19968 (N_19968,N_19742,N_19744);
or U19969 (N_19969,N_19630,N_19685);
and U19970 (N_19970,N_19736,N_19773);
or U19971 (N_19971,N_19653,N_19608);
nand U19972 (N_19972,N_19709,N_19616);
or U19973 (N_19973,N_19629,N_19671);
and U19974 (N_19974,N_19658,N_19616);
nor U19975 (N_19975,N_19638,N_19767);
xnor U19976 (N_19976,N_19780,N_19730);
or U19977 (N_19977,N_19605,N_19674);
nand U19978 (N_19978,N_19617,N_19751);
or U19979 (N_19979,N_19707,N_19718);
and U19980 (N_19980,N_19724,N_19777);
nor U19981 (N_19981,N_19759,N_19792);
or U19982 (N_19982,N_19614,N_19781);
or U19983 (N_19983,N_19650,N_19619);
nor U19984 (N_19984,N_19734,N_19714);
nand U19985 (N_19985,N_19784,N_19774);
xnor U19986 (N_19986,N_19723,N_19695);
nor U19987 (N_19987,N_19735,N_19707);
and U19988 (N_19988,N_19609,N_19639);
nor U19989 (N_19989,N_19658,N_19751);
and U19990 (N_19990,N_19620,N_19692);
nor U19991 (N_19991,N_19720,N_19712);
and U19992 (N_19992,N_19628,N_19609);
or U19993 (N_19993,N_19765,N_19689);
xnor U19994 (N_19994,N_19784,N_19792);
and U19995 (N_19995,N_19741,N_19759);
xnor U19996 (N_19996,N_19623,N_19662);
nand U19997 (N_19997,N_19756,N_19671);
xnor U19998 (N_19998,N_19678,N_19697);
and U19999 (N_19999,N_19642,N_19715);
nand UO_0 (O_0,N_19959,N_19910);
or UO_1 (O_1,N_19819,N_19982);
xnor UO_2 (O_2,N_19924,N_19941);
xor UO_3 (O_3,N_19877,N_19881);
nor UO_4 (O_4,N_19976,N_19993);
or UO_5 (O_5,N_19804,N_19902);
and UO_6 (O_6,N_19822,N_19886);
nor UO_7 (O_7,N_19890,N_19865);
nor UO_8 (O_8,N_19896,N_19970);
and UO_9 (O_9,N_19894,N_19884);
nand UO_10 (O_10,N_19810,N_19916);
and UO_11 (O_11,N_19934,N_19879);
xnor UO_12 (O_12,N_19957,N_19885);
xor UO_13 (O_13,N_19901,N_19805);
and UO_14 (O_14,N_19987,N_19992);
and UO_15 (O_15,N_19814,N_19847);
nor UO_16 (O_16,N_19917,N_19815);
and UO_17 (O_17,N_19843,N_19835);
xnor UO_18 (O_18,N_19802,N_19882);
nand UO_19 (O_19,N_19907,N_19842);
nor UO_20 (O_20,N_19958,N_19828);
nor UO_21 (O_21,N_19988,N_19928);
or UO_22 (O_22,N_19960,N_19892);
xor UO_23 (O_23,N_19997,N_19969);
nand UO_24 (O_24,N_19812,N_19820);
nand UO_25 (O_25,N_19813,N_19834);
or UO_26 (O_26,N_19953,N_19854);
xor UO_27 (O_27,N_19871,N_19999);
nor UO_28 (O_28,N_19998,N_19921);
nor UO_29 (O_29,N_19913,N_19850);
nor UO_30 (O_30,N_19839,N_19965);
xnor UO_31 (O_31,N_19833,N_19837);
nand UO_32 (O_32,N_19887,N_19899);
nand UO_33 (O_33,N_19829,N_19977);
or UO_34 (O_34,N_19922,N_19836);
nand UO_35 (O_35,N_19940,N_19844);
nor UO_36 (O_36,N_19849,N_19831);
nand UO_37 (O_37,N_19889,N_19860);
nor UO_38 (O_38,N_19906,N_19967);
nor UO_39 (O_39,N_19990,N_19898);
nand UO_40 (O_40,N_19868,N_19840);
nor UO_41 (O_41,N_19827,N_19862);
and UO_42 (O_42,N_19873,N_19980);
and UO_43 (O_43,N_19874,N_19955);
and UO_44 (O_44,N_19878,N_19948);
xnor UO_45 (O_45,N_19925,N_19848);
or UO_46 (O_46,N_19989,N_19944);
nand UO_47 (O_47,N_19893,N_19912);
nor UO_48 (O_48,N_19986,N_19864);
nor UO_49 (O_49,N_19908,N_19818);
and UO_50 (O_50,N_19876,N_19947);
and UO_51 (O_51,N_19938,N_19920);
or UO_52 (O_52,N_19852,N_19954);
xor UO_53 (O_53,N_19996,N_19811);
and UO_54 (O_54,N_19949,N_19933);
and UO_55 (O_55,N_19929,N_19891);
or UO_56 (O_56,N_19951,N_19909);
or UO_57 (O_57,N_19883,N_19966);
xnor UO_58 (O_58,N_19816,N_19861);
xor UO_59 (O_59,N_19950,N_19935);
nand UO_60 (O_60,N_19964,N_19923);
or UO_61 (O_61,N_19900,N_19832);
or UO_62 (O_62,N_19809,N_19939);
xor UO_63 (O_63,N_19825,N_19895);
and UO_64 (O_64,N_19888,N_19973);
nor UO_65 (O_65,N_19845,N_19838);
and UO_66 (O_66,N_19978,N_19905);
or UO_67 (O_67,N_19851,N_19943);
and UO_68 (O_68,N_19870,N_19956);
and UO_69 (O_69,N_19826,N_19994);
and UO_70 (O_70,N_19869,N_19821);
and UO_71 (O_71,N_19936,N_19962);
xnor UO_72 (O_72,N_19981,N_19857);
xor UO_73 (O_73,N_19972,N_19853);
xor UO_74 (O_74,N_19866,N_19856);
nand UO_75 (O_75,N_19937,N_19927);
xnor UO_76 (O_76,N_19995,N_19946);
and UO_77 (O_77,N_19983,N_19904);
and UO_78 (O_78,N_19846,N_19915);
nor UO_79 (O_79,N_19823,N_19824);
or UO_80 (O_80,N_19918,N_19926);
xor UO_81 (O_81,N_19961,N_19919);
nor UO_82 (O_82,N_19808,N_19963);
nor UO_83 (O_83,N_19872,N_19903);
and UO_84 (O_84,N_19855,N_19875);
nand UO_85 (O_85,N_19968,N_19952);
nor UO_86 (O_86,N_19800,N_19830);
xnor UO_87 (O_87,N_19897,N_19841);
nand UO_88 (O_88,N_19858,N_19975);
or UO_89 (O_89,N_19942,N_19974);
xor UO_90 (O_90,N_19971,N_19801);
nor UO_91 (O_91,N_19803,N_19931);
and UO_92 (O_92,N_19979,N_19985);
nand UO_93 (O_93,N_19859,N_19807);
and UO_94 (O_94,N_19930,N_19806);
or UO_95 (O_95,N_19911,N_19945);
nor UO_96 (O_96,N_19932,N_19991);
xor UO_97 (O_97,N_19867,N_19914);
or UO_98 (O_98,N_19880,N_19817);
or UO_99 (O_99,N_19863,N_19984);
nor UO_100 (O_100,N_19959,N_19985);
and UO_101 (O_101,N_19932,N_19930);
nor UO_102 (O_102,N_19954,N_19931);
and UO_103 (O_103,N_19941,N_19954);
nor UO_104 (O_104,N_19882,N_19900);
and UO_105 (O_105,N_19831,N_19850);
and UO_106 (O_106,N_19845,N_19813);
nand UO_107 (O_107,N_19869,N_19924);
or UO_108 (O_108,N_19888,N_19941);
nand UO_109 (O_109,N_19944,N_19815);
xor UO_110 (O_110,N_19969,N_19883);
or UO_111 (O_111,N_19875,N_19892);
or UO_112 (O_112,N_19923,N_19902);
nand UO_113 (O_113,N_19938,N_19946);
xnor UO_114 (O_114,N_19814,N_19976);
and UO_115 (O_115,N_19873,N_19811);
xor UO_116 (O_116,N_19958,N_19951);
and UO_117 (O_117,N_19829,N_19803);
nand UO_118 (O_118,N_19864,N_19817);
or UO_119 (O_119,N_19904,N_19925);
nor UO_120 (O_120,N_19823,N_19813);
nand UO_121 (O_121,N_19978,N_19998);
nand UO_122 (O_122,N_19811,N_19905);
xor UO_123 (O_123,N_19951,N_19992);
and UO_124 (O_124,N_19947,N_19852);
or UO_125 (O_125,N_19819,N_19925);
or UO_126 (O_126,N_19814,N_19956);
nor UO_127 (O_127,N_19917,N_19970);
nor UO_128 (O_128,N_19927,N_19930);
or UO_129 (O_129,N_19894,N_19898);
nor UO_130 (O_130,N_19938,N_19871);
and UO_131 (O_131,N_19981,N_19993);
nand UO_132 (O_132,N_19940,N_19863);
and UO_133 (O_133,N_19845,N_19920);
nand UO_134 (O_134,N_19904,N_19953);
xnor UO_135 (O_135,N_19853,N_19945);
nor UO_136 (O_136,N_19808,N_19814);
and UO_137 (O_137,N_19842,N_19968);
xnor UO_138 (O_138,N_19917,N_19848);
nor UO_139 (O_139,N_19837,N_19962);
xor UO_140 (O_140,N_19875,N_19983);
xor UO_141 (O_141,N_19891,N_19890);
or UO_142 (O_142,N_19860,N_19880);
or UO_143 (O_143,N_19834,N_19936);
and UO_144 (O_144,N_19845,N_19997);
and UO_145 (O_145,N_19987,N_19944);
nor UO_146 (O_146,N_19815,N_19933);
or UO_147 (O_147,N_19945,N_19880);
nand UO_148 (O_148,N_19933,N_19841);
xor UO_149 (O_149,N_19886,N_19845);
nand UO_150 (O_150,N_19961,N_19808);
nand UO_151 (O_151,N_19944,N_19900);
xor UO_152 (O_152,N_19938,N_19847);
xnor UO_153 (O_153,N_19846,N_19857);
nand UO_154 (O_154,N_19953,N_19861);
or UO_155 (O_155,N_19991,N_19870);
or UO_156 (O_156,N_19861,N_19997);
xor UO_157 (O_157,N_19887,N_19877);
xor UO_158 (O_158,N_19838,N_19976);
xnor UO_159 (O_159,N_19816,N_19981);
nand UO_160 (O_160,N_19964,N_19938);
xnor UO_161 (O_161,N_19870,N_19884);
or UO_162 (O_162,N_19822,N_19899);
and UO_163 (O_163,N_19924,N_19948);
nor UO_164 (O_164,N_19857,N_19858);
nor UO_165 (O_165,N_19873,N_19943);
xor UO_166 (O_166,N_19877,N_19979);
and UO_167 (O_167,N_19897,N_19857);
or UO_168 (O_168,N_19861,N_19945);
and UO_169 (O_169,N_19884,N_19982);
and UO_170 (O_170,N_19856,N_19839);
nor UO_171 (O_171,N_19866,N_19810);
nand UO_172 (O_172,N_19859,N_19856);
nand UO_173 (O_173,N_19827,N_19958);
or UO_174 (O_174,N_19822,N_19880);
or UO_175 (O_175,N_19942,N_19820);
nand UO_176 (O_176,N_19908,N_19999);
or UO_177 (O_177,N_19995,N_19930);
nor UO_178 (O_178,N_19874,N_19817);
xnor UO_179 (O_179,N_19940,N_19827);
nand UO_180 (O_180,N_19869,N_19953);
nor UO_181 (O_181,N_19816,N_19847);
nand UO_182 (O_182,N_19955,N_19979);
xor UO_183 (O_183,N_19864,N_19992);
nand UO_184 (O_184,N_19840,N_19881);
nor UO_185 (O_185,N_19869,N_19941);
or UO_186 (O_186,N_19895,N_19914);
or UO_187 (O_187,N_19897,N_19868);
nor UO_188 (O_188,N_19884,N_19873);
nand UO_189 (O_189,N_19949,N_19825);
nor UO_190 (O_190,N_19902,N_19838);
xor UO_191 (O_191,N_19888,N_19966);
xor UO_192 (O_192,N_19929,N_19987);
nor UO_193 (O_193,N_19936,N_19838);
or UO_194 (O_194,N_19866,N_19822);
nor UO_195 (O_195,N_19866,N_19970);
nor UO_196 (O_196,N_19856,N_19901);
nand UO_197 (O_197,N_19894,N_19947);
nor UO_198 (O_198,N_19800,N_19960);
nand UO_199 (O_199,N_19891,N_19803);
or UO_200 (O_200,N_19863,N_19989);
and UO_201 (O_201,N_19917,N_19905);
or UO_202 (O_202,N_19808,N_19994);
or UO_203 (O_203,N_19844,N_19930);
and UO_204 (O_204,N_19935,N_19932);
nor UO_205 (O_205,N_19883,N_19939);
xnor UO_206 (O_206,N_19851,N_19899);
and UO_207 (O_207,N_19803,N_19971);
xor UO_208 (O_208,N_19957,N_19939);
or UO_209 (O_209,N_19820,N_19876);
nor UO_210 (O_210,N_19935,N_19993);
nand UO_211 (O_211,N_19952,N_19853);
xor UO_212 (O_212,N_19910,N_19832);
xnor UO_213 (O_213,N_19909,N_19851);
and UO_214 (O_214,N_19873,N_19838);
nor UO_215 (O_215,N_19966,N_19822);
nor UO_216 (O_216,N_19972,N_19969);
nor UO_217 (O_217,N_19850,N_19855);
nand UO_218 (O_218,N_19827,N_19913);
nor UO_219 (O_219,N_19831,N_19835);
or UO_220 (O_220,N_19903,N_19832);
and UO_221 (O_221,N_19921,N_19800);
xnor UO_222 (O_222,N_19812,N_19956);
and UO_223 (O_223,N_19973,N_19970);
nand UO_224 (O_224,N_19811,N_19872);
or UO_225 (O_225,N_19997,N_19873);
and UO_226 (O_226,N_19950,N_19874);
nand UO_227 (O_227,N_19947,N_19813);
or UO_228 (O_228,N_19819,N_19831);
nor UO_229 (O_229,N_19942,N_19956);
and UO_230 (O_230,N_19878,N_19876);
nand UO_231 (O_231,N_19853,N_19873);
nand UO_232 (O_232,N_19996,N_19858);
nand UO_233 (O_233,N_19946,N_19808);
nor UO_234 (O_234,N_19819,N_19991);
xor UO_235 (O_235,N_19954,N_19994);
nor UO_236 (O_236,N_19974,N_19997);
nor UO_237 (O_237,N_19812,N_19938);
nor UO_238 (O_238,N_19916,N_19862);
xor UO_239 (O_239,N_19824,N_19921);
and UO_240 (O_240,N_19890,N_19971);
nand UO_241 (O_241,N_19933,N_19965);
or UO_242 (O_242,N_19864,N_19932);
nand UO_243 (O_243,N_19951,N_19896);
xnor UO_244 (O_244,N_19941,N_19881);
xnor UO_245 (O_245,N_19954,N_19807);
and UO_246 (O_246,N_19867,N_19902);
nand UO_247 (O_247,N_19818,N_19864);
or UO_248 (O_248,N_19989,N_19928);
nand UO_249 (O_249,N_19849,N_19937);
nand UO_250 (O_250,N_19973,N_19911);
nor UO_251 (O_251,N_19866,N_19809);
and UO_252 (O_252,N_19901,N_19926);
or UO_253 (O_253,N_19982,N_19898);
nand UO_254 (O_254,N_19932,N_19834);
xnor UO_255 (O_255,N_19936,N_19873);
or UO_256 (O_256,N_19897,N_19984);
nor UO_257 (O_257,N_19850,N_19912);
nand UO_258 (O_258,N_19807,N_19936);
nor UO_259 (O_259,N_19979,N_19833);
nand UO_260 (O_260,N_19952,N_19886);
nand UO_261 (O_261,N_19990,N_19926);
xor UO_262 (O_262,N_19962,N_19904);
nand UO_263 (O_263,N_19843,N_19915);
xnor UO_264 (O_264,N_19919,N_19917);
or UO_265 (O_265,N_19910,N_19901);
xnor UO_266 (O_266,N_19828,N_19809);
or UO_267 (O_267,N_19851,N_19813);
xnor UO_268 (O_268,N_19873,N_19960);
xor UO_269 (O_269,N_19854,N_19929);
xnor UO_270 (O_270,N_19800,N_19875);
nand UO_271 (O_271,N_19952,N_19807);
xor UO_272 (O_272,N_19993,N_19876);
nor UO_273 (O_273,N_19885,N_19852);
and UO_274 (O_274,N_19906,N_19869);
nor UO_275 (O_275,N_19942,N_19927);
nor UO_276 (O_276,N_19899,N_19815);
nand UO_277 (O_277,N_19804,N_19811);
or UO_278 (O_278,N_19831,N_19946);
xnor UO_279 (O_279,N_19918,N_19884);
and UO_280 (O_280,N_19817,N_19845);
nand UO_281 (O_281,N_19849,N_19855);
nor UO_282 (O_282,N_19887,N_19915);
nand UO_283 (O_283,N_19958,N_19950);
and UO_284 (O_284,N_19836,N_19907);
or UO_285 (O_285,N_19804,N_19833);
nand UO_286 (O_286,N_19811,N_19901);
nand UO_287 (O_287,N_19895,N_19844);
nand UO_288 (O_288,N_19841,N_19921);
nand UO_289 (O_289,N_19898,N_19822);
nor UO_290 (O_290,N_19929,N_19983);
xor UO_291 (O_291,N_19946,N_19817);
nor UO_292 (O_292,N_19923,N_19860);
nor UO_293 (O_293,N_19949,N_19954);
nor UO_294 (O_294,N_19866,N_19944);
xor UO_295 (O_295,N_19824,N_19857);
xor UO_296 (O_296,N_19821,N_19937);
or UO_297 (O_297,N_19923,N_19891);
and UO_298 (O_298,N_19927,N_19894);
nor UO_299 (O_299,N_19988,N_19929);
or UO_300 (O_300,N_19813,N_19992);
nor UO_301 (O_301,N_19807,N_19938);
nor UO_302 (O_302,N_19823,N_19952);
and UO_303 (O_303,N_19808,N_19886);
and UO_304 (O_304,N_19862,N_19895);
or UO_305 (O_305,N_19948,N_19839);
nand UO_306 (O_306,N_19855,N_19906);
nand UO_307 (O_307,N_19858,N_19803);
nand UO_308 (O_308,N_19807,N_19841);
xnor UO_309 (O_309,N_19806,N_19952);
nor UO_310 (O_310,N_19896,N_19883);
or UO_311 (O_311,N_19954,N_19871);
nor UO_312 (O_312,N_19994,N_19854);
and UO_313 (O_313,N_19870,N_19920);
and UO_314 (O_314,N_19942,N_19802);
nor UO_315 (O_315,N_19985,N_19890);
nand UO_316 (O_316,N_19811,N_19862);
or UO_317 (O_317,N_19821,N_19944);
xor UO_318 (O_318,N_19993,N_19803);
and UO_319 (O_319,N_19966,N_19943);
xor UO_320 (O_320,N_19990,N_19961);
and UO_321 (O_321,N_19835,N_19936);
xor UO_322 (O_322,N_19902,N_19899);
nor UO_323 (O_323,N_19993,N_19853);
nand UO_324 (O_324,N_19815,N_19988);
nor UO_325 (O_325,N_19872,N_19877);
nor UO_326 (O_326,N_19966,N_19857);
xor UO_327 (O_327,N_19837,N_19854);
xnor UO_328 (O_328,N_19997,N_19884);
xnor UO_329 (O_329,N_19862,N_19934);
xor UO_330 (O_330,N_19959,N_19895);
or UO_331 (O_331,N_19847,N_19920);
or UO_332 (O_332,N_19866,N_19994);
nand UO_333 (O_333,N_19953,N_19838);
nand UO_334 (O_334,N_19909,N_19956);
xor UO_335 (O_335,N_19984,N_19829);
nor UO_336 (O_336,N_19802,N_19832);
xnor UO_337 (O_337,N_19921,N_19975);
nand UO_338 (O_338,N_19852,N_19848);
and UO_339 (O_339,N_19944,N_19957);
nand UO_340 (O_340,N_19800,N_19976);
xor UO_341 (O_341,N_19993,N_19869);
nor UO_342 (O_342,N_19942,N_19830);
xor UO_343 (O_343,N_19813,N_19913);
or UO_344 (O_344,N_19826,N_19882);
nor UO_345 (O_345,N_19991,N_19864);
nand UO_346 (O_346,N_19976,N_19884);
or UO_347 (O_347,N_19831,N_19893);
and UO_348 (O_348,N_19860,N_19850);
xnor UO_349 (O_349,N_19974,N_19876);
and UO_350 (O_350,N_19883,N_19886);
nor UO_351 (O_351,N_19802,N_19992);
nand UO_352 (O_352,N_19939,N_19802);
xor UO_353 (O_353,N_19950,N_19903);
nor UO_354 (O_354,N_19801,N_19848);
nor UO_355 (O_355,N_19921,N_19918);
nor UO_356 (O_356,N_19911,N_19924);
nor UO_357 (O_357,N_19854,N_19894);
nand UO_358 (O_358,N_19947,N_19990);
and UO_359 (O_359,N_19803,N_19894);
xor UO_360 (O_360,N_19969,N_19819);
xnor UO_361 (O_361,N_19936,N_19923);
nor UO_362 (O_362,N_19885,N_19937);
xnor UO_363 (O_363,N_19917,N_19819);
nor UO_364 (O_364,N_19893,N_19947);
nand UO_365 (O_365,N_19810,N_19890);
or UO_366 (O_366,N_19942,N_19822);
nor UO_367 (O_367,N_19847,N_19979);
xnor UO_368 (O_368,N_19999,N_19918);
nand UO_369 (O_369,N_19984,N_19940);
xnor UO_370 (O_370,N_19808,N_19839);
nor UO_371 (O_371,N_19824,N_19938);
and UO_372 (O_372,N_19894,N_19957);
or UO_373 (O_373,N_19907,N_19824);
nor UO_374 (O_374,N_19922,N_19911);
nand UO_375 (O_375,N_19897,N_19961);
xor UO_376 (O_376,N_19961,N_19906);
and UO_377 (O_377,N_19949,N_19814);
or UO_378 (O_378,N_19814,N_19936);
nor UO_379 (O_379,N_19806,N_19860);
xor UO_380 (O_380,N_19823,N_19940);
nor UO_381 (O_381,N_19826,N_19801);
and UO_382 (O_382,N_19992,N_19869);
or UO_383 (O_383,N_19981,N_19875);
nor UO_384 (O_384,N_19927,N_19898);
nand UO_385 (O_385,N_19918,N_19851);
nor UO_386 (O_386,N_19836,N_19829);
nand UO_387 (O_387,N_19864,N_19843);
nor UO_388 (O_388,N_19896,N_19879);
and UO_389 (O_389,N_19946,N_19842);
or UO_390 (O_390,N_19955,N_19910);
xor UO_391 (O_391,N_19801,N_19915);
xor UO_392 (O_392,N_19990,N_19885);
xnor UO_393 (O_393,N_19828,N_19887);
xnor UO_394 (O_394,N_19996,N_19849);
nor UO_395 (O_395,N_19919,N_19996);
or UO_396 (O_396,N_19950,N_19805);
xor UO_397 (O_397,N_19836,N_19981);
and UO_398 (O_398,N_19826,N_19855);
or UO_399 (O_399,N_19924,N_19843);
nor UO_400 (O_400,N_19981,N_19847);
and UO_401 (O_401,N_19817,N_19899);
xnor UO_402 (O_402,N_19801,N_19830);
nor UO_403 (O_403,N_19907,N_19967);
and UO_404 (O_404,N_19854,N_19961);
nand UO_405 (O_405,N_19925,N_19975);
nand UO_406 (O_406,N_19813,N_19943);
nand UO_407 (O_407,N_19867,N_19849);
and UO_408 (O_408,N_19880,N_19907);
xnor UO_409 (O_409,N_19973,N_19912);
xnor UO_410 (O_410,N_19821,N_19963);
xor UO_411 (O_411,N_19954,N_19802);
nand UO_412 (O_412,N_19975,N_19869);
nand UO_413 (O_413,N_19804,N_19800);
and UO_414 (O_414,N_19854,N_19958);
nor UO_415 (O_415,N_19828,N_19929);
nand UO_416 (O_416,N_19857,N_19960);
xnor UO_417 (O_417,N_19912,N_19946);
and UO_418 (O_418,N_19904,N_19872);
nand UO_419 (O_419,N_19993,N_19957);
nor UO_420 (O_420,N_19815,N_19903);
nor UO_421 (O_421,N_19888,N_19873);
nor UO_422 (O_422,N_19837,N_19929);
xnor UO_423 (O_423,N_19860,N_19924);
nor UO_424 (O_424,N_19901,N_19826);
xnor UO_425 (O_425,N_19860,N_19996);
and UO_426 (O_426,N_19929,N_19964);
nor UO_427 (O_427,N_19956,N_19889);
xnor UO_428 (O_428,N_19931,N_19917);
and UO_429 (O_429,N_19830,N_19859);
and UO_430 (O_430,N_19855,N_19959);
and UO_431 (O_431,N_19920,N_19994);
nor UO_432 (O_432,N_19889,N_19969);
xnor UO_433 (O_433,N_19977,N_19872);
or UO_434 (O_434,N_19958,N_19896);
nand UO_435 (O_435,N_19832,N_19951);
or UO_436 (O_436,N_19803,N_19836);
or UO_437 (O_437,N_19921,N_19830);
or UO_438 (O_438,N_19948,N_19824);
nand UO_439 (O_439,N_19976,N_19977);
nor UO_440 (O_440,N_19919,N_19938);
nor UO_441 (O_441,N_19818,N_19835);
and UO_442 (O_442,N_19809,N_19813);
nor UO_443 (O_443,N_19992,N_19820);
nor UO_444 (O_444,N_19955,N_19863);
xnor UO_445 (O_445,N_19874,N_19839);
or UO_446 (O_446,N_19920,N_19929);
nand UO_447 (O_447,N_19897,N_19982);
and UO_448 (O_448,N_19871,N_19881);
nand UO_449 (O_449,N_19909,N_19816);
xnor UO_450 (O_450,N_19827,N_19938);
nand UO_451 (O_451,N_19988,N_19836);
xor UO_452 (O_452,N_19834,N_19987);
xor UO_453 (O_453,N_19903,N_19908);
or UO_454 (O_454,N_19909,N_19813);
nor UO_455 (O_455,N_19828,N_19827);
nand UO_456 (O_456,N_19848,N_19884);
nor UO_457 (O_457,N_19903,N_19996);
nand UO_458 (O_458,N_19906,N_19960);
nor UO_459 (O_459,N_19979,N_19876);
and UO_460 (O_460,N_19935,N_19961);
or UO_461 (O_461,N_19815,N_19926);
xnor UO_462 (O_462,N_19841,N_19931);
nor UO_463 (O_463,N_19875,N_19988);
xnor UO_464 (O_464,N_19823,N_19801);
nand UO_465 (O_465,N_19892,N_19817);
and UO_466 (O_466,N_19998,N_19888);
and UO_467 (O_467,N_19894,N_19920);
nand UO_468 (O_468,N_19894,N_19870);
and UO_469 (O_469,N_19915,N_19807);
nor UO_470 (O_470,N_19816,N_19836);
and UO_471 (O_471,N_19800,N_19932);
nand UO_472 (O_472,N_19992,N_19833);
and UO_473 (O_473,N_19995,N_19889);
nor UO_474 (O_474,N_19983,N_19917);
or UO_475 (O_475,N_19819,N_19810);
nor UO_476 (O_476,N_19989,N_19886);
xnor UO_477 (O_477,N_19845,N_19913);
or UO_478 (O_478,N_19953,N_19911);
or UO_479 (O_479,N_19949,N_19974);
and UO_480 (O_480,N_19991,N_19916);
nor UO_481 (O_481,N_19908,N_19892);
nor UO_482 (O_482,N_19815,N_19983);
and UO_483 (O_483,N_19868,N_19822);
nor UO_484 (O_484,N_19957,N_19824);
and UO_485 (O_485,N_19805,N_19823);
nand UO_486 (O_486,N_19914,N_19836);
and UO_487 (O_487,N_19913,N_19950);
xor UO_488 (O_488,N_19894,N_19950);
xnor UO_489 (O_489,N_19900,N_19903);
xor UO_490 (O_490,N_19812,N_19863);
or UO_491 (O_491,N_19855,N_19820);
nor UO_492 (O_492,N_19889,N_19976);
nand UO_493 (O_493,N_19849,N_19941);
nand UO_494 (O_494,N_19970,N_19847);
or UO_495 (O_495,N_19806,N_19980);
nor UO_496 (O_496,N_19978,N_19928);
nor UO_497 (O_497,N_19848,N_19937);
or UO_498 (O_498,N_19869,N_19947);
or UO_499 (O_499,N_19913,N_19877);
nand UO_500 (O_500,N_19923,N_19801);
and UO_501 (O_501,N_19824,N_19873);
nor UO_502 (O_502,N_19887,N_19843);
or UO_503 (O_503,N_19854,N_19987);
nand UO_504 (O_504,N_19803,N_19920);
nand UO_505 (O_505,N_19809,N_19816);
and UO_506 (O_506,N_19843,N_19992);
and UO_507 (O_507,N_19895,N_19804);
nor UO_508 (O_508,N_19992,N_19944);
or UO_509 (O_509,N_19850,N_19996);
or UO_510 (O_510,N_19891,N_19902);
nor UO_511 (O_511,N_19937,N_19893);
xnor UO_512 (O_512,N_19902,N_19999);
nor UO_513 (O_513,N_19835,N_19808);
nand UO_514 (O_514,N_19948,N_19900);
and UO_515 (O_515,N_19960,N_19881);
nand UO_516 (O_516,N_19927,N_19994);
xor UO_517 (O_517,N_19850,N_19908);
xor UO_518 (O_518,N_19917,N_19865);
or UO_519 (O_519,N_19935,N_19805);
nor UO_520 (O_520,N_19828,N_19905);
nand UO_521 (O_521,N_19801,N_19862);
and UO_522 (O_522,N_19960,N_19974);
xnor UO_523 (O_523,N_19997,N_19972);
nor UO_524 (O_524,N_19915,N_19837);
nor UO_525 (O_525,N_19880,N_19804);
nor UO_526 (O_526,N_19822,N_19968);
or UO_527 (O_527,N_19890,N_19820);
nand UO_528 (O_528,N_19942,N_19930);
or UO_529 (O_529,N_19899,N_19985);
or UO_530 (O_530,N_19903,N_19917);
nor UO_531 (O_531,N_19889,N_19821);
nand UO_532 (O_532,N_19879,N_19959);
or UO_533 (O_533,N_19835,N_19849);
and UO_534 (O_534,N_19986,N_19985);
nor UO_535 (O_535,N_19957,N_19847);
and UO_536 (O_536,N_19823,N_19838);
or UO_537 (O_537,N_19848,N_19820);
nand UO_538 (O_538,N_19951,N_19827);
xor UO_539 (O_539,N_19819,N_19921);
nand UO_540 (O_540,N_19979,N_19898);
xor UO_541 (O_541,N_19986,N_19866);
or UO_542 (O_542,N_19931,N_19977);
xnor UO_543 (O_543,N_19926,N_19974);
or UO_544 (O_544,N_19915,N_19826);
nand UO_545 (O_545,N_19889,N_19943);
nor UO_546 (O_546,N_19990,N_19959);
or UO_547 (O_547,N_19872,N_19821);
nor UO_548 (O_548,N_19904,N_19830);
nand UO_549 (O_549,N_19837,N_19937);
nand UO_550 (O_550,N_19896,N_19874);
and UO_551 (O_551,N_19844,N_19842);
xor UO_552 (O_552,N_19826,N_19911);
and UO_553 (O_553,N_19942,N_19893);
nand UO_554 (O_554,N_19990,N_19911);
nor UO_555 (O_555,N_19812,N_19869);
or UO_556 (O_556,N_19922,N_19897);
nand UO_557 (O_557,N_19936,N_19876);
xnor UO_558 (O_558,N_19841,N_19817);
nand UO_559 (O_559,N_19819,N_19930);
or UO_560 (O_560,N_19926,N_19871);
nor UO_561 (O_561,N_19816,N_19996);
nor UO_562 (O_562,N_19834,N_19900);
xnor UO_563 (O_563,N_19968,N_19901);
xor UO_564 (O_564,N_19815,N_19950);
and UO_565 (O_565,N_19954,N_19848);
and UO_566 (O_566,N_19833,N_19927);
nor UO_567 (O_567,N_19940,N_19842);
nor UO_568 (O_568,N_19980,N_19916);
or UO_569 (O_569,N_19828,N_19837);
nand UO_570 (O_570,N_19840,N_19810);
or UO_571 (O_571,N_19953,N_19927);
xnor UO_572 (O_572,N_19861,N_19905);
nand UO_573 (O_573,N_19861,N_19913);
nand UO_574 (O_574,N_19818,N_19853);
and UO_575 (O_575,N_19978,N_19847);
and UO_576 (O_576,N_19837,N_19979);
or UO_577 (O_577,N_19962,N_19980);
or UO_578 (O_578,N_19901,N_19862);
and UO_579 (O_579,N_19861,N_19932);
and UO_580 (O_580,N_19935,N_19945);
xor UO_581 (O_581,N_19995,N_19819);
nor UO_582 (O_582,N_19826,N_19962);
nor UO_583 (O_583,N_19914,N_19972);
or UO_584 (O_584,N_19881,N_19819);
or UO_585 (O_585,N_19830,N_19819);
nand UO_586 (O_586,N_19869,N_19868);
or UO_587 (O_587,N_19940,N_19838);
nand UO_588 (O_588,N_19848,N_19845);
and UO_589 (O_589,N_19852,N_19818);
nand UO_590 (O_590,N_19837,N_19874);
xor UO_591 (O_591,N_19803,N_19876);
or UO_592 (O_592,N_19864,N_19911);
xor UO_593 (O_593,N_19813,N_19862);
nand UO_594 (O_594,N_19863,N_19861);
and UO_595 (O_595,N_19969,N_19851);
nor UO_596 (O_596,N_19914,N_19911);
nand UO_597 (O_597,N_19840,N_19851);
nor UO_598 (O_598,N_19971,N_19848);
xor UO_599 (O_599,N_19907,N_19990);
nor UO_600 (O_600,N_19808,N_19998);
nor UO_601 (O_601,N_19850,N_19942);
xnor UO_602 (O_602,N_19873,N_19933);
xnor UO_603 (O_603,N_19809,N_19977);
xor UO_604 (O_604,N_19889,N_19910);
nor UO_605 (O_605,N_19810,N_19822);
and UO_606 (O_606,N_19945,N_19838);
nand UO_607 (O_607,N_19846,N_19822);
xor UO_608 (O_608,N_19832,N_19908);
nand UO_609 (O_609,N_19844,N_19877);
and UO_610 (O_610,N_19940,N_19891);
nand UO_611 (O_611,N_19851,N_19841);
nand UO_612 (O_612,N_19807,N_19978);
nor UO_613 (O_613,N_19916,N_19859);
nor UO_614 (O_614,N_19804,N_19959);
xor UO_615 (O_615,N_19826,N_19902);
xor UO_616 (O_616,N_19865,N_19921);
nand UO_617 (O_617,N_19883,N_19952);
or UO_618 (O_618,N_19944,N_19947);
nand UO_619 (O_619,N_19846,N_19881);
nand UO_620 (O_620,N_19918,N_19902);
nand UO_621 (O_621,N_19870,N_19971);
or UO_622 (O_622,N_19969,N_19875);
xnor UO_623 (O_623,N_19808,N_19995);
nor UO_624 (O_624,N_19959,N_19861);
nor UO_625 (O_625,N_19911,N_19895);
nor UO_626 (O_626,N_19928,N_19901);
xor UO_627 (O_627,N_19960,N_19891);
nor UO_628 (O_628,N_19861,N_19960);
nor UO_629 (O_629,N_19991,N_19994);
xnor UO_630 (O_630,N_19816,N_19913);
or UO_631 (O_631,N_19989,N_19986);
and UO_632 (O_632,N_19980,N_19863);
nand UO_633 (O_633,N_19810,N_19902);
nor UO_634 (O_634,N_19852,N_19803);
and UO_635 (O_635,N_19872,N_19863);
xnor UO_636 (O_636,N_19977,N_19911);
or UO_637 (O_637,N_19909,N_19819);
nand UO_638 (O_638,N_19953,N_19954);
nand UO_639 (O_639,N_19988,N_19938);
and UO_640 (O_640,N_19825,N_19938);
nor UO_641 (O_641,N_19863,N_19848);
nand UO_642 (O_642,N_19883,N_19910);
nand UO_643 (O_643,N_19931,N_19851);
nand UO_644 (O_644,N_19801,N_19879);
nor UO_645 (O_645,N_19904,N_19929);
nand UO_646 (O_646,N_19834,N_19877);
nor UO_647 (O_647,N_19902,N_19905);
or UO_648 (O_648,N_19986,N_19888);
xor UO_649 (O_649,N_19856,N_19804);
nor UO_650 (O_650,N_19820,N_19996);
nand UO_651 (O_651,N_19960,N_19997);
nand UO_652 (O_652,N_19907,N_19886);
nand UO_653 (O_653,N_19817,N_19853);
xnor UO_654 (O_654,N_19847,N_19869);
nor UO_655 (O_655,N_19907,N_19912);
nand UO_656 (O_656,N_19834,N_19837);
or UO_657 (O_657,N_19924,N_19872);
and UO_658 (O_658,N_19863,N_19917);
and UO_659 (O_659,N_19865,N_19978);
xor UO_660 (O_660,N_19908,N_19843);
or UO_661 (O_661,N_19897,N_19883);
xor UO_662 (O_662,N_19852,N_19862);
xor UO_663 (O_663,N_19834,N_19884);
or UO_664 (O_664,N_19875,N_19900);
nor UO_665 (O_665,N_19922,N_19890);
xor UO_666 (O_666,N_19941,N_19978);
nand UO_667 (O_667,N_19981,N_19961);
and UO_668 (O_668,N_19858,N_19952);
xnor UO_669 (O_669,N_19963,N_19949);
and UO_670 (O_670,N_19818,N_19931);
xnor UO_671 (O_671,N_19978,N_19858);
nor UO_672 (O_672,N_19978,N_19866);
nor UO_673 (O_673,N_19857,N_19997);
nor UO_674 (O_674,N_19906,N_19972);
and UO_675 (O_675,N_19869,N_19944);
nand UO_676 (O_676,N_19882,N_19869);
xor UO_677 (O_677,N_19843,N_19961);
and UO_678 (O_678,N_19865,N_19892);
or UO_679 (O_679,N_19947,N_19879);
and UO_680 (O_680,N_19997,N_19894);
and UO_681 (O_681,N_19895,N_19983);
nand UO_682 (O_682,N_19808,N_19951);
nand UO_683 (O_683,N_19832,N_19932);
nor UO_684 (O_684,N_19902,N_19952);
nand UO_685 (O_685,N_19842,N_19831);
xnor UO_686 (O_686,N_19801,N_19970);
xor UO_687 (O_687,N_19859,N_19938);
nand UO_688 (O_688,N_19913,N_19954);
nor UO_689 (O_689,N_19975,N_19982);
xor UO_690 (O_690,N_19853,N_19868);
nand UO_691 (O_691,N_19838,N_19911);
or UO_692 (O_692,N_19910,N_19951);
nand UO_693 (O_693,N_19827,N_19876);
or UO_694 (O_694,N_19945,N_19944);
xnor UO_695 (O_695,N_19999,N_19801);
xor UO_696 (O_696,N_19867,N_19812);
nand UO_697 (O_697,N_19864,N_19889);
xnor UO_698 (O_698,N_19973,N_19959);
and UO_699 (O_699,N_19962,N_19959);
nand UO_700 (O_700,N_19865,N_19884);
and UO_701 (O_701,N_19883,N_19859);
xor UO_702 (O_702,N_19875,N_19822);
nor UO_703 (O_703,N_19839,N_19807);
and UO_704 (O_704,N_19970,N_19958);
nand UO_705 (O_705,N_19957,N_19830);
and UO_706 (O_706,N_19931,N_19830);
nor UO_707 (O_707,N_19977,N_19854);
nor UO_708 (O_708,N_19972,N_19854);
nand UO_709 (O_709,N_19891,N_19885);
or UO_710 (O_710,N_19968,N_19924);
nor UO_711 (O_711,N_19969,N_19849);
and UO_712 (O_712,N_19850,N_19980);
nor UO_713 (O_713,N_19958,N_19856);
xnor UO_714 (O_714,N_19911,N_19818);
nand UO_715 (O_715,N_19934,N_19850);
and UO_716 (O_716,N_19904,N_19862);
or UO_717 (O_717,N_19875,N_19923);
xnor UO_718 (O_718,N_19882,N_19953);
nand UO_719 (O_719,N_19874,N_19947);
nand UO_720 (O_720,N_19899,N_19885);
or UO_721 (O_721,N_19828,N_19814);
nand UO_722 (O_722,N_19933,N_19853);
nor UO_723 (O_723,N_19970,N_19915);
nor UO_724 (O_724,N_19956,N_19906);
or UO_725 (O_725,N_19916,N_19874);
or UO_726 (O_726,N_19939,N_19994);
xnor UO_727 (O_727,N_19854,N_19868);
or UO_728 (O_728,N_19990,N_19840);
nand UO_729 (O_729,N_19866,N_19963);
xnor UO_730 (O_730,N_19983,N_19837);
nand UO_731 (O_731,N_19986,N_19967);
nand UO_732 (O_732,N_19935,N_19989);
nor UO_733 (O_733,N_19987,N_19942);
xor UO_734 (O_734,N_19802,N_19856);
nand UO_735 (O_735,N_19840,N_19928);
or UO_736 (O_736,N_19844,N_19831);
and UO_737 (O_737,N_19897,N_19871);
nor UO_738 (O_738,N_19966,N_19875);
nor UO_739 (O_739,N_19962,N_19811);
and UO_740 (O_740,N_19865,N_19906);
xor UO_741 (O_741,N_19845,N_19842);
xor UO_742 (O_742,N_19931,N_19808);
nor UO_743 (O_743,N_19959,N_19858);
or UO_744 (O_744,N_19909,N_19894);
and UO_745 (O_745,N_19868,N_19947);
nor UO_746 (O_746,N_19899,N_19994);
nor UO_747 (O_747,N_19848,N_19901);
nand UO_748 (O_748,N_19931,N_19813);
or UO_749 (O_749,N_19860,N_19934);
or UO_750 (O_750,N_19867,N_19853);
nor UO_751 (O_751,N_19912,N_19975);
nand UO_752 (O_752,N_19907,N_19997);
or UO_753 (O_753,N_19913,N_19880);
nand UO_754 (O_754,N_19853,N_19890);
nor UO_755 (O_755,N_19866,N_19996);
xor UO_756 (O_756,N_19825,N_19933);
xor UO_757 (O_757,N_19869,N_19881);
nor UO_758 (O_758,N_19922,N_19889);
and UO_759 (O_759,N_19808,N_19867);
or UO_760 (O_760,N_19940,N_19919);
and UO_761 (O_761,N_19911,N_19940);
xnor UO_762 (O_762,N_19956,N_19946);
and UO_763 (O_763,N_19975,N_19857);
or UO_764 (O_764,N_19941,N_19815);
or UO_765 (O_765,N_19885,N_19963);
nand UO_766 (O_766,N_19864,N_19846);
nand UO_767 (O_767,N_19857,N_19911);
nor UO_768 (O_768,N_19835,N_19905);
and UO_769 (O_769,N_19911,N_19904);
nor UO_770 (O_770,N_19940,N_19812);
nand UO_771 (O_771,N_19806,N_19872);
xor UO_772 (O_772,N_19822,N_19818);
nand UO_773 (O_773,N_19939,N_19858);
nand UO_774 (O_774,N_19916,N_19889);
or UO_775 (O_775,N_19978,N_19892);
xnor UO_776 (O_776,N_19812,N_19881);
and UO_777 (O_777,N_19894,N_19805);
or UO_778 (O_778,N_19805,N_19997);
and UO_779 (O_779,N_19904,N_19952);
xor UO_780 (O_780,N_19863,N_19821);
xnor UO_781 (O_781,N_19873,N_19948);
nand UO_782 (O_782,N_19998,N_19974);
nand UO_783 (O_783,N_19861,N_19873);
nand UO_784 (O_784,N_19965,N_19806);
and UO_785 (O_785,N_19848,N_19822);
and UO_786 (O_786,N_19872,N_19804);
or UO_787 (O_787,N_19912,N_19888);
nand UO_788 (O_788,N_19848,N_19859);
or UO_789 (O_789,N_19934,N_19984);
and UO_790 (O_790,N_19832,N_19920);
nand UO_791 (O_791,N_19902,N_19903);
xor UO_792 (O_792,N_19869,N_19843);
xor UO_793 (O_793,N_19866,N_19993);
xor UO_794 (O_794,N_19983,N_19892);
nand UO_795 (O_795,N_19825,N_19976);
and UO_796 (O_796,N_19823,N_19848);
or UO_797 (O_797,N_19814,N_19840);
nor UO_798 (O_798,N_19847,N_19975);
nor UO_799 (O_799,N_19802,N_19861);
xor UO_800 (O_800,N_19947,N_19882);
or UO_801 (O_801,N_19915,N_19835);
nand UO_802 (O_802,N_19820,N_19808);
and UO_803 (O_803,N_19866,N_19928);
nor UO_804 (O_804,N_19841,N_19896);
nand UO_805 (O_805,N_19815,N_19820);
and UO_806 (O_806,N_19817,N_19831);
or UO_807 (O_807,N_19902,N_19879);
xor UO_808 (O_808,N_19885,N_19813);
nand UO_809 (O_809,N_19851,N_19952);
nand UO_810 (O_810,N_19869,N_19859);
nor UO_811 (O_811,N_19902,N_19860);
and UO_812 (O_812,N_19953,N_19964);
nor UO_813 (O_813,N_19998,N_19943);
nor UO_814 (O_814,N_19933,N_19916);
nor UO_815 (O_815,N_19969,N_19894);
xor UO_816 (O_816,N_19984,N_19899);
xor UO_817 (O_817,N_19891,N_19889);
or UO_818 (O_818,N_19966,N_19823);
or UO_819 (O_819,N_19957,N_19862);
nand UO_820 (O_820,N_19897,N_19907);
nor UO_821 (O_821,N_19900,N_19925);
nand UO_822 (O_822,N_19886,N_19941);
and UO_823 (O_823,N_19863,N_19971);
nor UO_824 (O_824,N_19947,N_19927);
xor UO_825 (O_825,N_19913,N_19951);
and UO_826 (O_826,N_19984,N_19968);
xnor UO_827 (O_827,N_19966,N_19889);
xor UO_828 (O_828,N_19861,N_19804);
or UO_829 (O_829,N_19818,N_19817);
nand UO_830 (O_830,N_19860,N_19997);
nor UO_831 (O_831,N_19800,N_19999);
or UO_832 (O_832,N_19967,N_19872);
nand UO_833 (O_833,N_19873,N_19903);
nor UO_834 (O_834,N_19822,N_19975);
xnor UO_835 (O_835,N_19923,N_19982);
or UO_836 (O_836,N_19805,N_19858);
nor UO_837 (O_837,N_19965,N_19803);
or UO_838 (O_838,N_19938,N_19841);
and UO_839 (O_839,N_19935,N_19857);
or UO_840 (O_840,N_19851,N_19983);
xnor UO_841 (O_841,N_19987,N_19909);
and UO_842 (O_842,N_19815,N_19989);
nor UO_843 (O_843,N_19880,N_19980);
and UO_844 (O_844,N_19911,N_19883);
nor UO_845 (O_845,N_19844,N_19814);
nand UO_846 (O_846,N_19882,N_19977);
nand UO_847 (O_847,N_19874,N_19965);
or UO_848 (O_848,N_19856,N_19822);
nor UO_849 (O_849,N_19922,N_19983);
xnor UO_850 (O_850,N_19986,N_19996);
nor UO_851 (O_851,N_19940,N_19996);
and UO_852 (O_852,N_19945,N_19909);
xor UO_853 (O_853,N_19989,N_19866);
and UO_854 (O_854,N_19819,N_19892);
and UO_855 (O_855,N_19947,N_19979);
xor UO_856 (O_856,N_19981,N_19899);
nand UO_857 (O_857,N_19903,N_19817);
nor UO_858 (O_858,N_19921,N_19812);
or UO_859 (O_859,N_19868,N_19824);
xnor UO_860 (O_860,N_19886,N_19958);
nor UO_861 (O_861,N_19869,N_19972);
and UO_862 (O_862,N_19882,N_19962);
or UO_863 (O_863,N_19910,N_19939);
or UO_864 (O_864,N_19829,N_19878);
or UO_865 (O_865,N_19876,N_19950);
nor UO_866 (O_866,N_19908,N_19933);
or UO_867 (O_867,N_19903,N_19982);
or UO_868 (O_868,N_19924,N_19877);
nor UO_869 (O_869,N_19817,N_19916);
nand UO_870 (O_870,N_19820,N_19964);
and UO_871 (O_871,N_19802,N_19948);
and UO_872 (O_872,N_19806,N_19949);
or UO_873 (O_873,N_19998,N_19996);
nor UO_874 (O_874,N_19918,N_19907);
or UO_875 (O_875,N_19896,N_19911);
xor UO_876 (O_876,N_19965,N_19951);
xnor UO_877 (O_877,N_19830,N_19827);
nor UO_878 (O_878,N_19822,N_19943);
xor UO_879 (O_879,N_19838,N_19811);
xor UO_880 (O_880,N_19865,N_19929);
nand UO_881 (O_881,N_19994,N_19982);
and UO_882 (O_882,N_19892,N_19885);
xnor UO_883 (O_883,N_19812,N_19843);
or UO_884 (O_884,N_19914,N_19825);
nor UO_885 (O_885,N_19835,N_19926);
or UO_886 (O_886,N_19827,N_19826);
nand UO_887 (O_887,N_19981,N_19881);
and UO_888 (O_888,N_19838,N_19855);
xor UO_889 (O_889,N_19992,N_19876);
nor UO_890 (O_890,N_19942,N_19821);
or UO_891 (O_891,N_19870,N_19809);
nand UO_892 (O_892,N_19979,N_19820);
nor UO_893 (O_893,N_19882,N_19859);
and UO_894 (O_894,N_19907,N_19917);
or UO_895 (O_895,N_19942,N_19812);
and UO_896 (O_896,N_19822,N_19806);
and UO_897 (O_897,N_19915,N_19957);
nor UO_898 (O_898,N_19826,N_19924);
xor UO_899 (O_899,N_19929,N_19813);
and UO_900 (O_900,N_19864,N_19972);
xnor UO_901 (O_901,N_19837,N_19839);
or UO_902 (O_902,N_19909,N_19868);
and UO_903 (O_903,N_19938,N_19869);
and UO_904 (O_904,N_19894,N_19823);
xor UO_905 (O_905,N_19995,N_19816);
and UO_906 (O_906,N_19821,N_19935);
nor UO_907 (O_907,N_19957,N_19873);
and UO_908 (O_908,N_19986,N_19875);
nand UO_909 (O_909,N_19838,N_19931);
xor UO_910 (O_910,N_19853,N_19935);
xor UO_911 (O_911,N_19852,N_19997);
or UO_912 (O_912,N_19843,N_19940);
nand UO_913 (O_913,N_19916,N_19926);
nand UO_914 (O_914,N_19992,N_19974);
nor UO_915 (O_915,N_19881,N_19912);
or UO_916 (O_916,N_19814,N_19963);
nand UO_917 (O_917,N_19878,N_19888);
or UO_918 (O_918,N_19943,N_19963);
nor UO_919 (O_919,N_19804,N_19957);
nor UO_920 (O_920,N_19941,N_19892);
and UO_921 (O_921,N_19882,N_19868);
and UO_922 (O_922,N_19876,N_19823);
xor UO_923 (O_923,N_19990,N_19858);
or UO_924 (O_924,N_19886,N_19914);
nand UO_925 (O_925,N_19923,N_19848);
nand UO_926 (O_926,N_19844,N_19988);
and UO_927 (O_927,N_19908,N_19813);
nand UO_928 (O_928,N_19982,N_19930);
and UO_929 (O_929,N_19994,N_19859);
nor UO_930 (O_930,N_19922,N_19932);
and UO_931 (O_931,N_19833,N_19999);
xnor UO_932 (O_932,N_19956,N_19925);
and UO_933 (O_933,N_19831,N_19926);
and UO_934 (O_934,N_19989,N_19831);
or UO_935 (O_935,N_19949,N_19817);
nand UO_936 (O_936,N_19978,N_19940);
or UO_937 (O_937,N_19886,N_19973);
and UO_938 (O_938,N_19836,N_19820);
nand UO_939 (O_939,N_19907,N_19931);
or UO_940 (O_940,N_19953,N_19921);
xnor UO_941 (O_941,N_19947,N_19800);
nand UO_942 (O_942,N_19945,N_19932);
and UO_943 (O_943,N_19939,N_19820);
xor UO_944 (O_944,N_19861,N_19969);
and UO_945 (O_945,N_19958,N_19992);
nand UO_946 (O_946,N_19931,N_19964);
and UO_947 (O_947,N_19957,N_19985);
xnor UO_948 (O_948,N_19974,N_19845);
xor UO_949 (O_949,N_19825,N_19812);
nor UO_950 (O_950,N_19826,N_19876);
xnor UO_951 (O_951,N_19852,N_19964);
nor UO_952 (O_952,N_19999,N_19809);
nand UO_953 (O_953,N_19955,N_19900);
xnor UO_954 (O_954,N_19854,N_19827);
xnor UO_955 (O_955,N_19996,N_19810);
nand UO_956 (O_956,N_19918,N_19820);
xnor UO_957 (O_957,N_19934,N_19920);
and UO_958 (O_958,N_19977,N_19837);
and UO_959 (O_959,N_19868,N_19915);
nor UO_960 (O_960,N_19984,N_19978);
nor UO_961 (O_961,N_19955,N_19883);
nand UO_962 (O_962,N_19995,N_19944);
and UO_963 (O_963,N_19854,N_19957);
nor UO_964 (O_964,N_19820,N_19875);
xor UO_965 (O_965,N_19990,N_19996);
nand UO_966 (O_966,N_19985,N_19808);
and UO_967 (O_967,N_19857,N_19844);
or UO_968 (O_968,N_19991,N_19838);
nand UO_969 (O_969,N_19880,N_19867);
nand UO_970 (O_970,N_19927,N_19962);
nor UO_971 (O_971,N_19852,N_19872);
nand UO_972 (O_972,N_19911,N_19963);
or UO_973 (O_973,N_19978,N_19840);
nor UO_974 (O_974,N_19981,N_19992);
xor UO_975 (O_975,N_19907,N_19866);
and UO_976 (O_976,N_19859,N_19971);
xor UO_977 (O_977,N_19909,N_19828);
or UO_978 (O_978,N_19999,N_19932);
nand UO_979 (O_979,N_19971,N_19862);
and UO_980 (O_980,N_19862,N_19919);
and UO_981 (O_981,N_19835,N_19854);
or UO_982 (O_982,N_19977,N_19832);
nand UO_983 (O_983,N_19916,N_19827);
or UO_984 (O_984,N_19970,N_19820);
and UO_985 (O_985,N_19815,N_19874);
and UO_986 (O_986,N_19847,N_19940);
or UO_987 (O_987,N_19829,N_19805);
xor UO_988 (O_988,N_19896,N_19960);
xnor UO_989 (O_989,N_19815,N_19974);
xor UO_990 (O_990,N_19989,N_19870);
xnor UO_991 (O_991,N_19814,N_19939);
nand UO_992 (O_992,N_19879,N_19849);
and UO_993 (O_993,N_19920,N_19999);
xnor UO_994 (O_994,N_19996,N_19808);
or UO_995 (O_995,N_19923,N_19876);
xnor UO_996 (O_996,N_19944,N_19836);
xor UO_997 (O_997,N_19880,N_19868);
or UO_998 (O_998,N_19829,N_19899);
xnor UO_999 (O_999,N_19885,N_19809);
nand UO_1000 (O_1000,N_19826,N_19842);
xnor UO_1001 (O_1001,N_19829,N_19873);
xnor UO_1002 (O_1002,N_19963,N_19980);
and UO_1003 (O_1003,N_19938,N_19872);
nand UO_1004 (O_1004,N_19935,N_19947);
nand UO_1005 (O_1005,N_19913,N_19835);
nor UO_1006 (O_1006,N_19895,N_19945);
or UO_1007 (O_1007,N_19895,N_19931);
and UO_1008 (O_1008,N_19837,N_19955);
nand UO_1009 (O_1009,N_19916,N_19922);
and UO_1010 (O_1010,N_19878,N_19835);
nor UO_1011 (O_1011,N_19876,N_19937);
xnor UO_1012 (O_1012,N_19893,N_19909);
xor UO_1013 (O_1013,N_19906,N_19925);
or UO_1014 (O_1014,N_19929,N_19878);
and UO_1015 (O_1015,N_19816,N_19834);
and UO_1016 (O_1016,N_19911,N_19991);
nand UO_1017 (O_1017,N_19855,N_19843);
nand UO_1018 (O_1018,N_19815,N_19936);
nor UO_1019 (O_1019,N_19828,N_19877);
nor UO_1020 (O_1020,N_19949,N_19977);
nor UO_1021 (O_1021,N_19898,N_19968);
and UO_1022 (O_1022,N_19887,N_19835);
xnor UO_1023 (O_1023,N_19903,N_19985);
nor UO_1024 (O_1024,N_19944,N_19860);
nand UO_1025 (O_1025,N_19845,N_19956);
nor UO_1026 (O_1026,N_19972,N_19824);
nor UO_1027 (O_1027,N_19912,N_19904);
nor UO_1028 (O_1028,N_19944,N_19894);
xor UO_1029 (O_1029,N_19947,N_19921);
nand UO_1030 (O_1030,N_19870,N_19847);
or UO_1031 (O_1031,N_19959,N_19829);
xor UO_1032 (O_1032,N_19935,N_19875);
and UO_1033 (O_1033,N_19872,N_19951);
nor UO_1034 (O_1034,N_19862,N_19993);
and UO_1035 (O_1035,N_19901,N_19842);
nor UO_1036 (O_1036,N_19984,N_19913);
nand UO_1037 (O_1037,N_19962,N_19835);
nand UO_1038 (O_1038,N_19859,N_19981);
nor UO_1039 (O_1039,N_19822,N_19870);
and UO_1040 (O_1040,N_19855,N_19973);
and UO_1041 (O_1041,N_19976,N_19820);
nand UO_1042 (O_1042,N_19839,N_19905);
or UO_1043 (O_1043,N_19987,N_19986);
nand UO_1044 (O_1044,N_19963,N_19835);
and UO_1045 (O_1045,N_19954,N_19958);
xnor UO_1046 (O_1046,N_19923,N_19944);
xor UO_1047 (O_1047,N_19829,N_19824);
nor UO_1048 (O_1048,N_19976,N_19861);
nand UO_1049 (O_1049,N_19904,N_19937);
nor UO_1050 (O_1050,N_19875,N_19941);
xor UO_1051 (O_1051,N_19850,N_19802);
xnor UO_1052 (O_1052,N_19850,N_19844);
xor UO_1053 (O_1053,N_19945,N_19875);
or UO_1054 (O_1054,N_19904,N_19986);
or UO_1055 (O_1055,N_19943,N_19980);
nand UO_1056 (O_1056,N_19819,N_19967);
nand UO_1057 (O_1057,N_19885,N_19859);
nand UO_1058 (O_1058,N_19966,N_19880);
xor UO_1059 (O_1059,N_19810,N_19804);
and UO_1060 (O_1060,N_19965,N_19848);
or UO_1061 (O_1061,N_19843,N_19878);
and UO_1062 (O_1062,N_19955,N_19936);
xor UO_1063 (O_1063,N_19942,N_19857);
nand UO_1064 (O_1064,N_19989,N_19857);
nand UO_1065 (O_1065,N_19964,N_19877);
or UO_1066 (O_1066,N_19819,N_19941);
or UO_1067 (O_1067,N_19832,N_19876);
nor UO_1068 (O_1068,N_19876,N_19946);
or UO_1069 (O_1069,N_19951,N_19915);
and UO_1070 (O_1070,N_19847,N_19965);
or UO_1071 (O_1071,N_19962,N_19863);
nor UO_1072 (O_1072,N_19828,N_19811);
nand UO_1073 (O_1073,N_19841,N_19850);
nand UO_1074 (O_1074,N_19954,N_19910);
nand UO_1075 (O_1075,N_19869,N_19905);
nand UO_1076 (O_1076,N_19898,N_19951);
nand UO_1077 (O_1077,N_19804,N_19825);
nor UO_1078 (O_1078,N_19847,N_19849);
xnor UO_1079 (O_1079,N_19865,N_19968);
xnor UO_1080 (O_1080,N_19936,N_19965);
and UO_1081 (O_1081,N_19973,N_19922);
nand UO_1082 (O_1082,N_19885,N_19842);
nand UO_1083 (O_1083,N_19935,N_19991);
nand UO_1084 (O_1084,N_19811,N_19845);
nand UO_1085 (O_1085,N_19931,N_19843);
nor UO_1086 (O_1086,N_19865,N_19828);
nand UO_1087 (O_1087,N_19908,N_19937);
nor UO_1088 (O_1088,N_19893,N_19931);
xnor UO_1089 (O_1089,N_19828,N_19893);
nor UO_1090 (O_1090,N_19923,N_19969);
and UO_1091 (O_1091,N_19933,N_19923);
xnor UO_1092 (O_1092,N_19886,N_19975);
and UO_1093 (O_1093,N_19966,N_19942);
nand UO_1094 (O_1094,N_19932,N_19885);
nor UO_1095 (O_1095,N_19871,N_19942);
nor UO_1096 (O_1096,N_19814,N_19911);
nand UO_1097 (O_1097,N_19822,N_19948);
xnor UO_1098 (O_1098,N_19882,N_19956);
nor UO_1099 (O_1099,N_19968,N_19869);
or UO_1100 (O_1100,N_19881,N_19935);
and UO_1101 (O_1101,N_19902,N_19994);
or UO_1102 (O_1102,N_19972,N_19803);
or UO_1103 (O_1103,N_19990,N_19970);
or UO_1104 (O_1104,N_19983,N_19950);
nor UO_1105 (O_1105,N_19963,N_19950);
or UO_1106 (O_1106,N_19821,N_19885);
or UO_1107 (O_1107,N_19867,N_19912);
nor UO_1108 (O_1108,N_19836,N_19852);
xnor UO_1109 (O_1109,N_19854,N_19916);
or UO_1110 (O_1110,N_19835,N_19994);
nand UO_1111 (O_1111,N_19814,N_19983);
nand UO_1112 (O_1112,N_19821,N_19835);
nor UO_1113 (O_1113,N_19886,N_19966);
xor UO_1114 (O_1114,N_19830,N_19953);
nand UO_1115 (O_1115,N_19848,N_19907);
xor UO_1116 (O_1116,N_19998,N_19953);
nor UO_1117 (O_1117,N_19806,N_19905);
xnor UO_1118 (O_1118,N_19901,N_19931);
xor UO_1119 (O_1119,N_19865,N_19949);
or UO_1120 (O_1120,N_19965,N_19827);
nor UO_1121 (O_1121,N_19951,N_19815);
and UO_1122 (O_1122,N_19935,N_19900);
nor UO_1123 (O_1123,N_19803,N_19867);
xor UO_1124 (O_1124,N_19994,N_19965);
and UO_1125 (O_1125,N_19802,N_19824);
nand UO_1126 (O_1126,N_19983,N_19946);
and UO_1127 (O_1127,N_19857,N_19874);
xnor UO_1128 (O_1128,N_19935,N_19915);
and UO_1129 (O_1129,N_19823,N_19948);
or UO_1130 (O_1130,N_19814,N_19950);
xor UO_1131 (O_1131,N_19998,N_19882);
nand UO_1132 (O_1132,N_19978,N_19863);
nand UO_1133 (O_1133,N_19972,N_19976);
nand UO_1134 (O_1134,N_19951,N_19949);
xor UO_1135 (O_1135,N_19860,N_19900);
xnor UO_1136 (O_1136,N_19802,N_19825);
xnor UO_1137 (O_1137,N_19978,N_19875);
xnor UO_1138 (O_1138,N_19849,N_19872);
and UO_1139 (O_1139,N_19931,N_19889);
xor UO_1140 (O_1140,N_19838,N_19874);
xnor UO_1141 (O_1141,N_19887,N_19852);
nand UO_1142 (O_1142,N_19909,N_19869);
or UO_1143 (O_1143,N_19875,N_19883);
xor UO_1144 (O_1144,N_19830,N_19935);
nor UO_1145 (O_1145,N_19972,N_19827);
or UO_1146 (O_1146,N_19928,N_19861);
nand UO_1147 (O_1147,N_19968,N_19903);
xor UO_1148 (O_1148,N_19916,N_19880);
or UO_1149 (O_1149,N_19959,N_19898);
and UO_1150 (O_1150,N_19828,N_19882);
nor UO_1151 (O_1151,N_19998,N_19897);
xor UO_1152 (O_1152,N_19874,N_19848);
or UO_1153 (O_1153,N_19815,N_19985);
and UO_1154 (O_1154,N_19893,N_19953);
and UO_1155 (O_1155,N_19885,N_19921);
nand UO_1156 (O_1156,N_19866,N_19921);
or UO_1157 (O_1157,N_19861,N_19985);
nor UO_1158 (O_1158,N_19895,N_19817);
and UO_1159 (O_1159,N_19840,N_19993);
and UO_1160 (O_1160,N_19817,N_19809);
and UO_1161 (O_1161,N_19830,N_19922);
nand UO_1162 (O_1162,N_19963,N_19974);
or UO_1163 (O_1163,N_19911,N_19842);
xnor UO_1164 (O_1164,N_19827,N_19861);
nand UO_1165 (O_1165,N_19830,N_19952);
xnor UO_1166 (O_1166,N_19962,N_19822);
and UO_1167 (O_1167,N_19967,N_19805);
xnor UO_1168 (O_1168,N_19940,N_19805);
nand UO_1169 (O_1169,N_19839,N_19997);
xor UO_1170 (O_1170,N_19993,N_19953);
xnor UO_1171 (O_1171,N_19815,N_19878);
nand UO_1172 (O_1172,N_19916,N_19867);
and UO_1173 (O_1173,N_19835,N_19932);
xor UO_1174 (O_1174,N_19805,N_19910);
or UO_1175 (O_1175,N_19868,N_19962);
nor UO_1176 (O_1176,N_19901,N_19972);
xor UO_1177 (O_1177,N_19929,N_19850);
or UO_1178 (O_1178,N_19837,N_19945);
or UO_1179 (O_1179,N_19977,N_19831);
nand UO_1180 (O_1180,N_19827,N_19963);
or UO_1181 (O_1181,N_19985,N_19873);
nand UO_1182 (O_1182,N_19806,N_19903);
nor UO_1183 (O_1183,N_19890,N_19958);
nor UO_1184 (O_1184,N_19953,N_19875);
nand UO_1185 (O_1185,N_19843,N_19936);
xnor UO_1186 (O_1186,N_19984,N_19816);
and UO_1187 (O_1187,N_19906,N_19873);
and UO_1188 (O_1188,N_19906,N_19991);
nor UO_1189 (O_1189,N_19823,N_19995);
and UO_1190 (O_1190,N_19823,N_19917);
and UO_1191 (O_1191,N_19937,N_19891);
nand UO_1192 (O_1192,N_19978,N_19823);
or UO_1193 (O_1193,N_19981,N_19959);
and UO_1194 (O_1194,N_19804,N_19878);
xor UO_1195 (O_1195,N_19829,N_19879);
nand UO_1196 (O_1196,N_19986,N_19912);
xnor UO_1197 (O_1197,N_19812,N_19932);
xnor UO_1198 (O_1198,N_19940,N_19972);
and UO_1199 (O_1199,N_19803,N_19914);
and UO_1200 (O_1200,N_19960,N_19953);
and UO_1201 (O_1201,N_19876,N_19999);
nor UO_1202 (O_1202,N_19854,N_19996);
or UO_1203 (O_1203,N_19956,N_19878);
and UO_1204 (O_1204,N_19996,N_19822);
xor UO_1205 (O_1205,N_19816,N_19969);
xor UO_1206 (O_1206,N_19869,N_19860);
xnor UO_1207 (O_1207,N_19912,N_19923);
nor UO_1208 (O_1208,N_19990,N_19857);
and UO_1209 (O_1209,N_19801,N_19832);
nor UO_1210 (O_1210,N_19875,N_19931);
nor UO_1211 (O_1211,N_19841,N_19983);
nor UO_1212 (O_1212,N_19990,N_19972);
and UO_1213 (O_1213,N_19808,N_19822);
nor UO_1214 (O_1214,N_19990,N_19997);
or UO_1215 (O_1215,N_19884,N_19854);
or UO_1216 (O_1216,N_19937,N_19944);
xor UO_1217 (O_1217,N_19931,N_19867);
nor UO_1218 (O_1218,N_19852,N_19855);
xor UO_1219 (O_1219,N_19990,N_19813);
xnor UO_1220 (O_1220,N_19866,N_19870);
xnor UO_1221 (O_1221,N_19985,N_19870);
and UO_1222 (O_1222,N_19855,N_19904);
and UO_1223 (O_1223,N_19960,N_19838);
and UO_1224 (O_1224,N_19945,N_19936);
nand UO_1225 (O_1225,N_19817,N_19807);
and UO_1226 (O_1226,N_19955,N_19844);
or UO_1227 (O_1227,N_19900,N_19964);
and UO_1228 (O_1228,N_19899,N_19997);
and UO_1229 (O_1229,N_19844,N_19941);
nand UO_1230 (O_1230,N_19804,N_19946);
nand UO_1231 (O_1231,N_19935,N_19813);
and UO_1232 (O_1232,N_19843,N_19960);
nand UO_1233 (O_1233,N_19977,N_19875);
nor UO_1234 (O_1234,N_19879,N_19819);
and UO_1235 (O_1235,N_19826,N_19919);
nor UO_1236 (O_1236,N_19871,N_19841);
and UO_1237 (O_1237,N_19913,N_19919);
and UO_1238 (O_1238,N_19865,N_19904);
nand UO_1239 (O_1239,N_19801,N_19919);
nor UO_1240 (O_1240,N_19887,N_19949);
and UO_1241 (O_1241,N_19851,N_19825);
and UO_1242 (O_1242,N_19931,N_19926);
or UO_1243 (O_1243,N_19873,N_19912);
nand UO_1244 (O_1244,N_19879,N_19965);
xnor UO_1245 (O_1245,N_19852,N_19924);
nand UO_1246 (O_1246,N_19977,N_19861);
and UO_1247 (O_1247,N_19924,N_19815);
nand UO_1248 (O_1248,N_19904,N_19993);
nand UO_1249 (O_1249,N_19844,N_19965);
nor UO_1250 (O_1250,N_19946,N_19935);
nor UO_1251 (O_1251,N_19974,N_19908);
xor UO_1252 (O_1252,N_19847,N_19959);
and UO_1253 (O_1253,N_19806,N_19911);
or UO_1254 (O_1254,N_19832,N_19905);
or UO_1255 (O_1255,N_19927,N_19890);
nand UO_1256 (O_1256,N_19976,N_19856);
or UO_1257 (O_1257,N_19806,N_19871);
nand UO_1258 (O_1258,N_19942,N_19973);
xor UO_1259 (O_1259,N_19867,N_19929);
or UO_1260 (O_1260,N_19853,N_19851);
or UO_1261 (O_1261,N_19819,N_19993);
or UO_1262 (O_1262,N_19972,N_19935);
or UO_1263 (O_1263,N_19987,N_19934);
nor UO_1264 (O_1264,N_19803,N_19885);
xnor UO_1265 (O_1265,N_19957,N_19807);
nand UO_1266 (O_1266,N_19843,N_19805);
nor UO_1267 (O_1267,N_19834,N_19970);
xor UO_1268 (O_1268,N_19936,N_19991);
xor UO_1269 (O_1269,N_19975,N_19972);
or UO_1270 (O_1270,N_19893,N_19811);
xnor UO_1271 (O_1271,N_19983,N_19848);
nand UO_1272 (O_1272,N_19852,N_19957);
xor UO_1273 (O_1273,N_19811,N_19936);
nor UO_1274 (O_1274,N_19863,N_19877);
nor UO_1275 (O_1275,N_19960,N_19977);
and UO_1276 (O_1276,N_19889,N_19963);
xor UO_1277 (O_1277,N_19981,N_19915);
or UO_1278 (O_1278,N_19863,N_19931);
nor UO_1279 (O_1279,N_19944,N_19926);
nand UO_1280 (O_1280,N_19916,N_19997);
or UO_1281 (O_1281,N_19832,N_19826);
and UO_1282 (O_1282,N_19873,N_19883);
xor UO_1283 (O_1283,N_19981,N_19918);
nand UO_1284 (O_1284,N_19893,N_19922);
nor UO_1285 (O_1285,N_19891,N_19907);
nor UO_1286 (O_1286,N_19996,N_19964);
xnor UO_1287 (O_1287,N_19813,N_19974);
nor UO_1288 (O_1288,N_19915,N_19947);
or UO_1289 (O_1289,N_19817,N_19802);
nor UO_1290 (O_1290,N_19935,N_19981);
nand UO_1291 (O_1291,N_19950,N_19858);
nor UO_1292 (O_1292,N_19855,N_19955);
and UO_1293 (O_1293,N_19965,N_19976);
or UO_1294 (O_1294,N_19890,N_19899);
and UO_1295 (O_1295,N_19922,N_19851);
nor UO_1296 (O_1296,N_19820,N_19929);
or UO_1297 (O_1297,N_19909,N_19938);
nor UO_1298 (O_1298,N_19924,N_19859);
and UO_1299 (O_1299,N_19863,N_19858);
or UO_1300 (O_1300,N_19877,N_19990);
xor UO_1301 (O_1301,N_19967,N_19913);
nor UO_1302 (O_1302,N_19954,N_19833);
or UO_1303 (O_1303,N_19821,N_19916);
nor UO_1304 (O_1304,N_19836,N_19847);
nor UO_1305 (O_1305,N_19809,N_19860);
nor UO_1306 (O_1306,N_19863,N_19944);
and UO_1307 (O_1307,N_19962,N_19849);
nand UO_1308 (O_1308,N_19955,N_19911);
nand UO_1309 (O_1309,N_19825,N_19868);
nor UO_1310 (O_1310,N_19958,N_19838);
nor UO_1311 (O_1311,N_19800,N_19823);
nor UO_1312 (O_1312,N_19831,N_19851);
or UO_1313 (O_1313,N_19949,N_19925);
nor UO_1314 (O_1314,N_19866,N_19865);
xor UO_1315 (O_1315,N_19900,N_19873);
xnor UO_1316 (O_1316,N_19859,N_19906);
and UO_1317 (O_1317,N_19972,N_19968);
and UO_1318 (O_1318,N_19939,N_19996);
and UO_1319 (O_1319,N_19836,N_19970);
or UO_1320 (O_1320,N_19902,N_19926);
nand UO_1321 (O_1321,N_19947,N_19857);
and UO_1322 (O_1322,N_19833,N_19828);
or UO_1323 (O_1323,N_19880,N_19991);
nand UO_1324 (O_1324,N_19894,N_19907);
nand UO_1325 (O_1325,N_19806,N_19962);
xnor UO_1326 (O_1326,N_19867,N_19895);
nand UO_1327 (O_1327,N_19954,N_19812);
nand UO_1328 (O_1328,N_19927,N_19920);
or UO_1329 (O_1329,N_19815,N_19841);
nand UO_1330 (O_1330,N_19869,N_19822);
nor UO_1331 (O_1331,N_19991,N_19900);
and UO_1332 (O_1332,N_19906,N_19883);
nand UO_1333 (O_1333,N_19917,N_19918);
nand UO_1334 (O_1334,N_19810,N_19909);
xor UO_1335 (O_1335,N_19960,N_19889);
xnor UO_1336 (O_1336,N_19957,N_19895);
and UO_1337 (O_1337,N_19961,N_19964);
or UO_1338 (O_1338,N_19819,N_19940);
nor UO_1339 (O_1339,N_19951,N_19914);
and UO_1340 (O_1340,N_19992,N_19904);
nor UO_1341 (O_1341,N_19936,N_19891);
nand UO_1342 (O_1342,N_19849,N_19992);
nand UO_1343 (O_1343,N_19933,N_19924);
xor UO_1344 (O_1344,N_19966,N_19982);
nand UO_1345 (O_1345,N_19840,N_19807);
or UO_1346 (O_1346,N_19902,N_19841);
xnor UO_1347 (O_1347,N_19874,N_19830);
nand UO_1348 (O_1348,N_19847,N_19990);
xnor UO_1349 (O_1349,N_19999,N_19928);
nand UO_1350 (O_1350,N_19877,N_19820);
xor UO_1351 (O_1351,N_19970,N_19981);
and UO_1352 (O_1352,N_19805,N_19838);
or UO_1353 (O_1353,N_19954,N_19977);
or UO_1354 (O_1354,N_19928,N_19938);
nand UO_1355 (O_1355,N_19802,N_19920);
and UO_1356 (O_1356,N_19878,N_19949);
nor UO_1357 (O_1357,N_19952,N_19936);
and UO_1358 (O_1358,N_19927,N_19859);
and UO_1359 (O_1359,N_19898,N_19992);
xor UO_1360 (O_1360,N_19842,N_19944);
or UO_1361 (O_1361,N_19934,N_19954);
nand UO_1362 (O_1362,N_19837,N_19867);
or UO_1363 (O_1363,N_19813,N_19897);
nand UO_1364 (O_1364,N_19902,N_19939);
xnor UO_1365 (O_1365,N_19994,N_19942);
nor UO_1366 (O_1366,N_19997,N_19802);
xor UO_1367 (O_1367,N_19876,N_19967);
nor UO_1368 (O_1368,N_19956,N_19831);
nor UO_1369 (O_1369,N_19854,N_19822);
and UO_1370 (O_1370,N_19863,N_19916);
xor UO_1371 (O_1371,N_19866,N_19913);
or UO_1372 (O_1372,N_19991,N_19929);
and UO_1373 (O_1373,N_19927,N_19905);
or UO_1374 (O_1374,N_19979,N_19975);
nor UO_1375 (O_1375,N_19888,N_19808);
or UO_1376 (O_1376,N_19922,N_19887);
nand UO_1377 (O_1377,N_19888,N_19926);
nand UO_1378 (O_1378,N_19991,N_19845);
nand UO_1379 (O_1379,N_19900,N_19908);
nor UO_1380 (O_1380,N_19875,N_19869);
and UO_1381 (O_1381,N_19946,N_19835);
nand UO_1382 (O_1382,N_19893,N_19925);
nor UO_1383 (O_1383,N_19906,N_19989);
xnor UO_1384 (O_1384,N_19893,N_19964);
nand UO_1385 (O_1385,N_19975,N_19854);
or UO_1386 (O_1386,N_19949,N_19988);
nor UO_1387 (O_1387,N_19923,N_19868);
and UO_1388 (O_1388,N_19845,N_19933);
xor UO_1389 (O_1389,N_19928,N_19850);
nand UO_1390 (O_1390,N_19890,N_19867);
nand UO_1391 (O_1391,N_19986,N_19846);
nor UO_1392 (O_1392,N_19915,N_19805);
nor UO_1393 (O_1393,N_19823,N_19810);
or UO_1394 (O_1394,N_19965,N_19982);
nand UO_1395 (O_1395,N_19925,N_19828);
and UO_1396 (O_1396,N_19993,N_19802);
nand UO_1397 (O_1397,N_19983,N_19840);
or UO_1398 (O_1398,N_19808,N_19874);
or UO_1399 (O_1399,N_19841,N_19906);
nand UO_1400 (O_1400,N_19928,N_19879);
or UO_1401 (O_1401,N_19953,N_19999);
nand UO_1402 (O_1402,N_19910,N_19990);
nand UO_1403 (O_1403,N_19946,N_19903);
or UO_1404 (O_1404,N_19859,N_19901);
nor UO_1405 (O_1405,N_19965,N_19901);
and UO_1406 (O_1406,N_19958,N_19929);
nor UO_1407 (O_1407,N_19810,N_19879);
and UO_1408 (O_1408,N_19871,N_19959);
xor UO_1409 (O_1409,N_19803,N_19857);
nor UO_1410 (O_1410,N_19916,N_19938);
xor UO_1411 (O_1411,N_19957,N_19983);
or UO_1412 (O_1412,N_19890,N_19843);
and UO_1413 (O_1413,N_19856,N_19940);
nor UO_1414 (O_1414,N_19997,N_19874);
xnor UO_1415 (O_1415,N_19841,N_19993);
or UO_1416 (O_1416,N_19925,N_19983);
or UO_1417 (O_1417,N_19826,N_19982);
nand UO_1418 (O_1418,N_19813,N_19805);
and UO_1419 (O_1419,N_19905,N_19858);
and UO_1420 (O_1420,N_19900,N_19870);
or UO_1421 (O_1421,N_19974,N_19829);
nor UO_1422 (O_1422,N_19986,N_19842);
and UO_1423 (O_1423,N_19865,N_19971);
and UO_1424 (O_1424,N_19835,N_19801);
and UO_1425 (O_1425,N_19990,N_19859);
nor UO_1426 (O_1426,N_19968,N_19886);
and UO_1427 (O_1427,N_19986,N_19998);
or UO_1428 (O_1428,N_19885,N_19972);
nor UO_1429 (O_1429,N_19804,N_19828);
or UO_1430 (O_1430,N_19811,N_19823);
and UO_1431 (O_1431,N_19833,N_19921);
nand UO_1432 (O_1432,N_19830,N_19861);
xor UO_1433 (O_1433,N_19818,N_19891);
and UO_1434 (O_1434,N_19856,N_19945);
nand UO_1435 (O_1435,N_19866,N_19915);
or UO_1436 (O_1436,N_19815,N_19822);
nor UO_1437 (O_1437,N_19883,N_19942);
and UO_1438 (O_1438,N_19929,N_19999);
or UO_1439 (O_1439,N_19986,N_19804);
or UO_1440 (O_1440,N_19892,N_19944);
or UO_1441 (O_1441,N_19851,N_19944);
or UO_1442 (O_1442,N_19838,N_19842);
or UO_1443 (O_1443,N_19902,N_19970);
or UO_1444 (O_1444,N_19813,N_19800);
nor UO_1445 (O_1445,N_19997,N_19898);
nor UO_1446 (O_1446,N_19941,N_19876);
nor UO_1447 (O_1447,N_19990,N_19814);
xor UO_1448 (O_1448,N_19900,N_19851);
xnor UO_1449 (O_1449,N_19907,N_19913);
nand UO_1450 (O_1450,N_19812,N_19830);
xor UO_1451 (O_1451,N_19878,N_19933);
or UO_1452 (O_1452,N_19822,N_19926);
and UO_1453 (O_1453,N_19950,N_19945);
nor UO_1454 (O_1454,N_19853,N_19806);
and UO_1455 (O_1455,N_19826,N_19927);
nor UO_1456 (O_1456,N_19881,N_19864);
and UO_1457 (O_1457,N_19918,N_19952);
xnor UO_1458 (O_1458,N_19950,N_19822);
xor UO_1459 (O_1459,N_19967,N_19858);
xnor UO_1460 (O_1460,N_19816,N_19800);
and UO_1461 (O_1461,N_19984,N_19970);
and UO_1462 (O_1462,N_19871,N_19878);
or UO_1463 (O_1463,N_19870,N_19863);
nand UO_1464 (O_1464,N_19973,N_19838);
xnor UO_1465 (O_1465,N_19974,N_19901);
xor UO_1466 (O_1466,N_19813,N_19985);
and UO_1467 (O_1467,N_19812,N_19969);
nand UO_1468 (O_1468,N_19830,N_19919);
xor UO_1469 (O_1469,N_19884,N_19899);
nand UO_1470 (O_1470,N_19944,N_19981);
nand UO_1471 (O_1471,N_19936,N_19868);
and UO_1472 (O_1472,N_19870,N_19980);
and UO_1473 (O_1473,N_19912,N_19927);
or UO_1474 (O_1474,N_19954,N_19948);
nor UO_1475 (O_1475,N_19979,N_19861);
xor UO_1476 (O_1476,N_19821,N_19890);
nor UO_1477 (O_1477,N_19920,N_19889);
nor UO_1478 (O_1478,N_19892,N_19808);
or UO_1479 (O_1479,N_19987,N_19805);
nand UO_1480 (O_1480,N_19993,N_19805);
or UO_1481 (O_1481,N_19965,N_19986);
nor UO_1482 (O_1482,N_19993,N_19958);
and UO_1483 (O_1483,N_19846,N_19893);
xor UO_1484 (O_1484,N_19844,N_19881);
or UO_1485 (O_1485,N_19858,N_19916);
nand UO_1486 (O_1486,N_19964,N_19973);
nor UO_1487 (O_1487,N_19811,N_19906);
or UO_1488 (O_1488,N_19874,N_19954);
or UO_1489 (O_1489,N_19957,N_19914);
xnor UO_1490 (O_1490,N_19961,N_19802);
xnor UO_1491 (O_1491,N_19936,N_19881);
or UO_1492 (O_1492,N_19997,N_19814);
nand UO_1493 (O_1493,N_19871,N_19973);
nor UO_1494 (O_1494,N_19830,N_19898);
nor UO_1495 (O_1495,N_19832,N_19853);
xor UO_1496 (O_1496,N_19884,N_19908);
and UO_1497 (O_1497,N_19825,N_19883);
and UO_1498 (O_1498,N_19908,N_19985);
xor UO_1499 (O_1499,N_19932,N_19938);
and UO_1500 (O_1500,N_19850,N_19848);
nand UO_1501 (O_1501,N_19979,N_19856);
or UO_1502 (O_1502,N_19836,N_19994);
and UO_1503 (O_1503,N_19833,N_19849);
xnor UO_1504 (O_1504,N_19850,N_19865);
xor UO_1505 (O_1505,N_19905,N_19932);
or UO_1506 (O_1506,N_19844,N_19973);
or UO_1507 (O_1507,N_19924,N_19833);
nor UO_1508 (O_1508,N_19931,N_19911);
nand UO_1509 (O_1509,N_19941,N_19884);
nand UO_1510 (O_1510,N_19946,N_19884);
or UO_1511 (O_1511,N_19828,N_19997);
and UO_1512 (O_1512,N_19987,N_19831);
nand UO_1513 (O_1513,N_19977,N_19953);
or UO_1514 (O_1514,N_19977,N_19899);
or UO_1515 (O_1515,N_19845,N_19855);
xor UO_1516 (O_1516,N_19950,N_19956);
xor UO_1517 (O_1517,N_19919,N_19811);
nand UO_1518 (O_1518,N_19948,N_19945);
and UO_1519 (O_1519,N_19855,N_19886);
nor UO_1520 (O_1520,N_19931,N_19974);
nor UO_1521 (O_1521,N_19975,N_19820);
nor UO_1522 (O_1522,N_19810,N_19891);
or UO_1523 (O_1523,N_19988,N_19977);
nor UO_1524 (O_1524,N_19970,N_19911);
nor UO_1525 (O_1525,N_19960,N_19867);
nand UO_1526 (O_1526,N_19974,N_19804);
and UO_1527 (O_1527,N_19899,N_19904);
xnor UO_1528 (O_1528,N_19806,N_19924);
nand UO_1529 (O_1529,N_19952,N_19977);
or UO_1530 (O_1530,N_19901,N_19994);
nor UO_1531 (O_1531,N_19870,N_19804);
or UO_1532 (O_1532,N_19865,N_19999);
nand UO_1533 (O_1533,N_19837,N_19897);
and UO_1534 (O_1534,N_19815,N_19952);
and UO_1535 (O_1535,N_19973,N_19818);
and UO_1536 (O_1536,N_19861,N_19879);
or UO_1537 (O_1537,N_19961,N_19926);
nor UO_1538 (O_1538,N_19934,N_19981);
and UO_1539 (O_1539,N_19860,N_19827);
and UO_1540 (O_1540,N_19835,N_19964);
xor UO_1541 (O_1541,N_19894,N_19936);
nor UO_1542 (O_1542,N_19822,N_19986);
nor UO_1543 (O_1543,N_19983,N_19971);
xnor UO_1544 (O_1544,N_19823,N_19925);
nor UO_1545 (O_1545,N_19946,N_19950);
and UO_1546 (O_1546,N_19829,N_19833);
nand UO_1547 (O_1547,N_19889,N_19854);
or UO_1548 (O_1548,N_19881,N_19930);
xor UO_1549 (O_1549,N_19900,N_19896);
nor UO_1550 (O_1550,N_19949,N_19889);
or UO_1551 (O_1551,N_19957,N_19909);
nor UO_1552 (O_1552,N_19896,N_19807);
nand UO_1553 (O_1553,N_19942,N_19841);
or UO_1554 (O_1554,N_19951,N_19933);
and UO_1555 (O_1555,N_19856,N_19977);
and UO_1556 (O_1556,N_19802,N_19870);
nor UO_1557 (O_1557,N_19858,N_19836);
nand UO_1558 (O_1558,N_19859,N_19890);
or UO_1559 (O_1559,N_19877,N_19941);
nor UO_1560 (O_1560,N_19839,N_19866);
or UO_1561 (O_1561,N_19868,N_19928);
nor UO_1562 (O_1562,N_19803,N_19968);
nand UO_1563 (O_1563,N_19831,N_19958);
nand UO_1564 (O_1564,N_19918,N_19832);
xnor UO_1565 (O_1565,N_19865,N_19809);
and UO_1566 (O_1566,N_19815,N_19860);
and UO_1567 (O_1567,N_19873,N_19915);
nor UO_1568 (O_1568,N_19902,N_19874);
or UO_1569 (O_1569,N_19818,N_19982);
and UO_1570 (O_1570,N_19954,N_19805);
xor UO_1571 (O_1571,N_19847,N_19853);
and UO_1572 (O_1572,N_19834,N_19910);
and UO_1573 (O_1573,N_19973,N_19840);
nand UO_1574 (O_1574,N_19891,N_19988);
and UO_1575 (O_1575,N_19970,N_19994);
and UO_1576 (O_1576,N_19859,N_19819);
nor UO_1577 (O_1577,N_19835,N_19909);
and UO_1578 (O_1578,N_19881,N_19959);
and UO_1579 (O_1579,N_19816,N_19943);
or UO_1580 (O_1580,N_19844,N_19956);
or UO_1581 (O_1581,N_19936,N_19871);
nand UO_1582 (O_1582,N_19971,N_19820);
xnor UO_1583 (O_1583,N_19902,N_19829);
nor UO_1584 (O_1584,N_19811,N_19888);
nand UO_1585 (O_1585,N_19867,N_19816);
or UO_1586 (O_1586,N_19878,N_19906);
nand UO_1587 (O_1587,N_19899,N_19909);
xnor UO_1588 (O_1588,N_19985,N_19865);
and UO_1589 (O_1589,N_19855,N_19967);
and UO_1590 (O_1590,N_19801,N_19920);
xnor UO_1591 (O_1591,N_19914,N_19887);
and UO_1592 (O_1592,N_19812,N_19821);
xor UO_1593 (O_1593,N_19846,N_19934);
nand UO_1594 (O_1594,N_19843,N_19874);
or UO_1595 (O_1595,N_19871,N_19839);
and UO_1596 (O_1596,N_19801,N_19973);
and UO_1597 (O_1597,N_19915,N_19829);
xor UO_1598 (O_1598,N_19915,N_19966);
or UO_1599 (O_1599,N_19808,N_19826);
or UO_1600 (O_1600,N_19891,N_19845);
or UO_1601 (O_1601,N_19901,N_19911);
nand UO_1602 (O_1602,N_19957,N_19926);
xor UO_1603 (O_1603,N_19874,N_19899);
nand UO_1604 (O_1604,N_19967,N_19915);
or UO_1605 (O_1605,N_19903,N_19912);
nor UO_1606 (O_1606,N_19847,N_19999);
and UO_1607 (O_1607,N_19935,N_19916);
xnor UO_1608 (O_1608,N_19953,N_19902);
or UO_1609 (O_1609,N_19823,N_19921);
nand UO_1610 (O_1610,N_19828,N_19985);
nand UO_1611 (O_1611,N_19909,N_19824);
or UO_1612 (O_1612,N_19861,N_19845);
nor UO_1613 (O_1613,N_19977,N_19939);
xor UO_1614 (O_1614,N_19816,N_19926);
or UO_1615 (O_1615,N_19966,N_19945);
nand UO_1616 (O_1616,N_19992,N_19868);
xnor UO_1617 (O_1617,N_19931,N_19959);
nor UO_1618 (O_1618,N_19960,N_19899);
nand UO_1619 (O_1619,N_19838,N_19970);
or UO_1620 (O_1620,N_19810,N_19967);
nand UO_1621 (O_1621,N_19807,N_19838);
nand UO_1622 (O_1622,N_19960,N_19914);
xor UO_1623 (O_1623,N_19918,N_19986);
and UO_1624 (O_1624,N_19971,N_19840);
nor UO_1625 (O_1625,N_19819,N_19990);
and UO_1626 (O_1626,N_19842,N_19937);
nand UO_1627 (O_1627,N_19887,N_19907);
nor UO_1628 (O_1628,N_19820,N_19851);
and UO_1629 (O_1629,N_19977,N_19965);
or UO_1630 (O_1630,N_19920,N_19800);
or UO_1631 (O_1631,N_19917,N_19838);
and UO_1632 (O_1632,N_19867,N_19889);
xnor UO_1633 (O_1633,N_19889,N_19826);
and UO_1634 (O_1634,N_19918,N_19965);
xnor UO_1635 (O_1635,N_19871,N_19932);
xor UO_1636 (O_1636,N_19800,N_19930);
nand UO_1637 (O_1637,N_19940,N_19864);
nor UO_1638 (O_1638,N_19833,N_19931);
and UO_1639 (O_1639,N_19968,N_19871);
or UO_1640 (O_1640,N_19875,N_19812);
nand UO_1641 (O_1641,N_19893,N_19808);
nand UO_1642 (O_1642,N_19849,N_19944);
or UO_1643 (O_1643,N_19958,N_19937);
or UO_1644 (O_1644,N_19996,N_19959);
and UO_1645 (O_1645,N_19818,N_19871);
nand UO_1646 (O_1646,N_19908,N_19959);
nand UO_1647 (O_1647,N_19893,N_19957);
xor UO_1648 (O_1648,N_19917,N_19859);
nor UO_1649 (O_1649,N_19832,N_19986);
nand UO_1650 (O_1650,N_19914,N_19820);
and UO_1651 (O_1651,N_19917,N_19888);
and UO_1652 (O_1652,N_19925,N_19847);
and UO_1653 (O_1653,N_19874,N_19842);
or UO_1654 (O_1654,N_19998,N_19817);
or UO_1655 (O_1655,N_19986,N_19844);
nand UO_1656 (O_1656,N_19895,N_19883);
and UO_1657 (O_1657,N_19919,N_19849);
xor UO_1658 (O_1658,N_19824,N_19903);
nand UO_1659 (O_1659,N_19890,N_19938);
xor UO_1660 (O_1660,N_19841,N_19861);
and UO_1661 (O_1661,N_19905,N_19936);
nand UO_1662 (O_1662,N_19909,N_19878);
xnor UO_1663 (O_1663,N_19889,N_19870);
and UO_1664 (O_1664,N_19870,N_19922);
nor UO_1665 (O_1665,N_19807,N_19959);
and UO_1666 (O_1666,N_19812,N_19944);
and UO_1667 (O_1667,N_19993,N_19821);
xnor UO_1668 (O_1668,N_19916,N_19904);
nor UO_1669 (O_1669,N_19817,N_19945);
or UO_1670 (O_1670,N_19936,N_19922);
nor UO_1671 (O_1671,N_19845,N_19925);
and UO_1672 (O_1672,N_19815,N_19946);
and UO_1673 (O_1673,N_19832,N_19983);
and UO_1674 (O_1674,N_19843,N_19934);
nor UO_1675 (O_1675,N_19825,N_19911);
or UO_1676 (O_1676,N_19808,N_19997);
or UO_1677 (O_1677,N_19815,N_19991);
and UO_1678 (O_1678,N_19994,N_19801);
xnor UO_1679 (O_1679,N_19856,N_19999);
nor UO_1680 (O_1680,N_19871,N_19853);
and UO_1681 (O_1681,N_19800,N_19811);
xor UO_1682 (O_1682,N_19890,N_19906);
and UO_1683 (O_1683,N_19961,N_19894);
xnor UO_1684 (O_1684,N_19944,N_19985);
nor UO_1685 (O_1685,N_19820,N_19891);
or UO_1686 (O_1686,N_19978,N_19907);
nor UO_1687 (O_1687,N_19909,N_19946);
nand UO_1688 (O_1688,N_19819,N_19874);
or UO_1689 (O_1689,N_19821,N_19945);
and UO_1690 (O_1690,N_19950,N_19811);
xor UO_1691 (O_1691,N_19940,N_19829);
xnor UO_1692 (O_1692,N_19966,N_19920);
and UO_1693 (O_1693,N_19940,N_19813);
nor UO_1694 (O_1694,N_19921,N_19896);
or UO_1695 (O_1695,N_19849,N_19891);
or UO_1696 (O_1696,N_19889,N_19984);
nand UO_1697 (O_1697,N_19861,N_19946);
nand UO_1698 (O_1698,N_19966,N_19819);
nand UO_1699 (O_1699,N_19847,N_19828);
xor UO_1700 (O_1700,N_19973,N_19915);
nand UO_1701 (O_1701,N_19996,N_19918);
nor UO_1702 (O_1702,N_19893,N_19834);
xnor UO_1703 (O_1703,N_19829,N_19908);
nor UO_1704 (O_1704,N_19981,N_19939);
and UO_1705 (O_1705,N_19882,N_19983);
and UO_1706 (O_1706,N_19884,N_19823);
and UO_1707 (O_1707,N_19990,N_19976);
xor UO_1708 (O_1708,N_19890,N_19910);
and UO_1709 (O_1709,N_19974,N_19827);
xor UO_1710 (O_1710,N_19982,N_19937);
and UO_1711 (O_1711,N_19920,N_19974);
nor UO_1712 (O_1712,N_19976,N_19841);
and UO_1713 (O_1713,N_19996,N_19890);
nand UO_1714 (O_1714,N_19930,N_19997);
and UO_1715 (O_1715,N_19944,N_19867);
or UO_1716 (O_1716,N_19951,N_19927);
xnor UO_1717 (O_1717,N_19821,N_19856);
nand UO_1718 (O_1718,N_19951,N_19969);
nor UO_1719 (O_1719,N_19877,N_19912);
or UO_1720 (O_1720,N_19821,N_19913);
and UO_1721 (O_1721,N_19962,N_19805);
nand UO_1722 (O_1722,N_19935,N_19983);
and UO_1723 (O_1723,N_19967,N_19838);
nand UO_1724 (O_1724,N_19843,N_19819);
nor UO_1725 (O_1725,N_19961,N_19980);
nor UO_1726 (O_1726,N_19977,N_19883);
xor UO_1727 (O_1727,N_19950,N_19868);
xnor UO_1728 (O_1728,N_19926,N_19962);
nand UO_1729 (O_1729,N_19955,N_19918);
nand UO_1730 (O_1730,N_19932,N_19886);
xor UO_1731 (O_1731,N_19956,N_19949);
nand UO_1732 (O_1732,N_19975,N_19826);
nor UO_1733 (O_1733,N_19902,N_19909);
nand UO_1734 (O_1734,N_19992,N_19950);
nor UO_1735 (O_1735,N_19824,N_19987);
nand UO_1736 (O_1736,N_19847,N_19971);
and UO_1737 (O_1737,N_19960,N_19847);
and UO_1738 (O_1738,N_19932,N_19841);
nor UO_1739 (O_1739,N_19921,N_19886);
nor UO_1740 (O_1740,N_19957,N_19990);
and UO_1741 (O_1741,N_19811,N_19825);
nand UO_1742 (O_1742,N_19921,N_19860);
nor UO_1743 (O_1743,N_19887,N_19927);
nand UO_1744 (O_1744,N_19829,N_19893);
nand UO_1745 (O_1745,N_19989,N_19994);
and UO_1746 (O_1746,N_19981,N_19999);
nand UO_1747 (O_1747,N_19891,N_19814);
xnor UO_1748 (O_1748,N_19868,N_19953);
xnor UO_1749 (O_1749,N_19986,N_19891);
xor UO_1750 (O_1750,N_19935,N_19817);
or UO_1751 (O_1751,N_19935,N_19831);
and UO_1752 (O_1752,N_19840,N_19834);
and UO_1753 (O_1753,N_19935,N_19910);
xnor UO_1754 (O_1754,N_19965,N_19970);
xor UO_1755 (O_1755,N_19841,N_19927);
and UO_1756 (O_1756,N_19913,N_19867);
or UO_1757 (O_1757,N_19978,N_19885);
or UO_1758 (O_1758,N_19850,N_19961);
or UO_1759 (O_1759,N_19829,N_19807);
and UO_1760 (O_1760,N_19847,N_19987);
nand UO_1761 (O_1761,N_19980,N_19941);
nor UO_1762 (O_1762,N_19853,N_19959);
nor UO_1763 (O_1763,N_19943,N_19940);
or UO_1764 (O_1764,N_19941,N_19962);
xor UO_1765 (O_1765,N_19820,N_19927);
xor UO_1766 (O_1766,N_19829,N_19918);
nor UO_1767 (O_1767,N_19905,N_19994);
and UO_1768 (O_1768,N_19880,N_19812);
xor UO_1769 (O_1769,N_19891,N_19873);
nor UO_1770 (O_1770,N_19831,N_19910);
xor UO_1771 (O_1771,N_19946,N_19928);
and UO_1772 (O_1772,N_19824,N_19919);
and UO_1773 (O_1773,N_19863,N_19804);
and UO_1774 (O_1774,N_19995,N_19958);
or UO_1775 (O_1775,N_19985,N_19869);
nand UO_1776 (O_1776,N_19828,N_19956);
nand UO_1777 (O_1777,N_19946,N_19940);
xor UO_1778 (O_1778,N_19945,N_19863);
or UO_1779 (O_1779,N_19984,N_19880);
and UO_1780 (O_1780,N_19885,N_19836);
xnor UO_1781 (O_1781,N_19907,N_19996);
and UO_1782 (O_1782,N_19968,N_19824);
or UO_1783 (O_1783,N_19981,N_19921);
or UO_1784 (O_1784,N_19809,N_19875);
nand UO_1785 (O_1785,N_19910,N_19981);
nand UO_1786 (O_1786,N_19828,N_19823);
or UO_1787 (O_1787,N_19913,N_19830);
nand UO_1788 (O_1788,N_19946,N_19837);
and UO_1789 (O_1789,N_19927,N_19861);
xnor UO_1790 (O_1790,N_19972,N_19865);
xnor UO_1791 (O_1791,N_19862,N_19912);
or UO_1792 (O_1792,N_19904,N_19982);
and UO_1793 (O_1793,N_19880,N_19936);
nor UO_1794 (O_1794,N_19804,N_19888);
xor UO_1795 (O_1795,N_19886,N_19959);
and UO_1796 (O_1796,N_19864,N_19878);
xor UO_1797 (O_1797,N_19828,N_19982);
nand UO_1798 (O_1798,N_19906,N_19918);
nand UO_1799 (O_1799,N_19970,N_19983);
or UO_1800 (O_1800,N_19985,N_19809);
nor UO_1801 (O_1801,N_19895,N_19998);
or UO_1802 (O_1802,N_19890,N_19991);
xnor UO_1803 (O_1803,N_19805,N_19988);
and UO_1804 (O_1804,N_19897,N_19911);
and UO_1805 (O_1805,N_19993,N_19936);
or UO_1806 (O_1806,N_19806,N_19939);
or UO_1807 (O_1807,N_19872,N_19992);
nand UO_1808 (O_1808,N_19948,N_19919);
and UO_1809 (O_1809,N_19926,N_19971);
and UO_1810 (O_1810,N_19913,N_19948);
xor UO_1811 (O_1811,N_19851,N_19979);
or UO_1812 (O_1812,N_19847,N_19848);
nor UO_1813 (O_1813,N_19978,N_19808);
nand UO_1814 (O_1814,N_19989,N_19950);
nand UO_1815 (O_1815,N_19864,N_19950);
or UO_1816 (O_1816,N_19920,N_19993);
nand UO_1817 (O_1817,N_19812,N_19971);
xnor UO_1818 (O_1818,N_19938,N_19966);
nand UO_1819 (O_1819,N_19973,N_19826);
xnor UO_1820 (O_1820,N_19968,N_19829);
nor UO_1821 (O_1821,N_19938,N_19877);
nand UO_1822 (O_1822,N_19967,N_19973);
or UO_1823 (O_1823,N_19862,N_19974);
nand UO_1824 (O_1824,N_19862,N_19845);
and UO_1825 (O_1825,N_19916,N_19899);
or UO_1826 (O_1826,N_19818,N_19896);
nand UO_1827 (O_1827,N_19922,N_19927);
or UO_1828 (O_1828,N_19949,N_19832);
nor UO_1829 (O_1829,N_19868,N_19814);
or UO_1830 (O_1830,N_19871,N_19960);
xor UO_1831 (O_1831,N_19880,N_19948);
and UO_1832 (O_1832,N_19945,N_19953);
nor UO_1833 (O_1833,N_19899,N_19908);
nor UO_1834 (O_1834,N_19883,N_19819);
xnor UO_1835 (O_1835,N_19874,N_19821);
xnor UO_1836 (O_1836,N_19829,N_19848);
or UO_1837 (O_1837,N_19840,N_19805);
or UO_1838 (O_1838,N_19925,N_19805);
nor UO_1839 (O_1839,N_19939,N_19990);
nand UO_1840 (O_1840,N_19882,N_19861);
nor UO_1841 (O_1841,N_19862,N_19892);
xnor UO_1842 (O_1842,N_19980,N_19856);
or UO_1843 (O_1843,N_19962,N_19860);
or UO_1844 (O_1844,N_19877,N_19893);
and UO_1845 (O_1845,N_19963,N_19855);
or UO_1846 (O_1846,N_19860,N_19847);
xor UO_1847 (O_1847,N_19889,N_19849);
nand UO_1848 (O_1848,N_19933,N_19920);
and UO_1849 (O_1849,N_19969,N_19949);
and UO_1850 (O_1850,N_19805,N_19883);
xnor UO_1851 (O_1851,N_19839,N_19918);
nor UO_1852 (O_1852,N_19906,N_19940);
nor UO_1853 (O_1853,N_19865,N_19997);
xnor UO_1854 (O_1854,N_19957,N_19837);
and UO_1855 (O_1855,N_19900,N_19996);
nand UO_1856 (O_1856,N_19937,N_19894);
or UO_1857 (O_1857,N_19822,N_19995);
nand UO_1858 (O_1858,N_19933,N_19801);
and UO_1859 (O_1859,N_19903,N_19959);
nand UO_1860 (O_1860,N_19978,N_19936);
nor UO_1861 (O_1861,N_19863,N_19827);
xnor UO_1862 (O_1862,N_19839,N_19820);
xor UO_1863 (O_1863,N_19904,N_19807);
and UO_1864 (O_1864,N_19835,N_19865);
or UO_1865 (O_1865,N_19876,N_19928);
nor UO_1866 (O_1866,N_19937,N_19971);
nor UO_1867 (O_1867,N_19946,N_19960);
and UO_1868 (O_1868,N_19853,N_19999);
or UO_1869 (O_1869,N_19944,N_19970);
nand UO_1870 (O_1870,N_19868,N_19918);
and UO_1871 (O_1871,N_19889,N_19919);
or UO_1872 (O_1872,N_19871,N_19912);
and UO_1873 (O_1873,N_19981,N_19987);
xnor UO_1874 (O_1874,N_19895,N_19928);
and UO_1875 (O_1875,N_19961,N_19969);
xor UO_1876 (O_1876,N_19904,N_19868);
nand UO_1877 (O_1877,N_19845,N_19979);
nand UO_1878 (O_1878,N_19917,N_19989);
or UO_1879 (O_1879,N_19977,N_19910);
or UO_1880 (O_1880,N_19902,N_19819);
nand UO_1881 (O_1881,N_19807,N_19903);
nand UO_1882 (O_1882,N_19970,N_19825);
xnor UO_1883 (O_1883,N_19818,N_19970);
or UO_1884 (O_1884,N_19998,N_19871);
xor UO_1885 (O_1885,N_19907,N_19854);
xor UO_1886 (O_1886,N_19815,N_19947);
nand UO_1887 (O_1887,N_19994,N_19924);
and UO_1888 (O_1888,N_19884,N_19827);
nand UO_1889 (O_1889,N_19859,N_19811);
nand UO_1890 (O_1890,N_19917,N_19998);
nand UO_1891 (O_1891,N_19818,N_19917);
xor UO_1892 (O_1892,N_19994,N_19967);
xor UO_1893 (O_1893,N_19960,N_19801);
or UO_1894 (O_1894,N_19877,N_19812);
nor UO_1895 (O_1895,N_19924,N_19980);
and UO_1896 (O_1896,N_19894,N_19996);
or UO_1897 (O_1897,N_19967,N_19890);
xor UO_1898 (O_1898,N_19814,N_19845);
or UO_1899 (O_1899,N_19916,N_19994);
nor UO_1900 (O_1900,N_19820,N_19895);
xnor UO_1901 (O_1901,N_19830,N_19862);
or UO_1902 (O_1902,N_19893,N_19904);
or UO_1903 (O_1903,N_19872,N_19855);
and UO_1904 (O_1904,N_19818,N_19934);
nand UO_1905 (O_1905,N_19925,N_19803);
and UO_1906 (O_1906,N_19909,N_19969);
xnor UO_1907 (O_1907,N_19823,N_19877);
xor UO_1908 (O_1908,N_19940,N_19865);
nand UO_1909 (O_1909,N_19902,N_19854);
xor UO_1910 (O_1910,N_19892,N_19900);
xor UO_1911 (O_1911,N_19883,N_19842);
nand UO_1912 (O_1912,N_19980,N_19817);
xor UO_1913 (O_1913,N_19851,N_19887);
nand UO_1914 (O_1914,N_19847,N_19878);
nand UO_1915 (O_1915,N_19831,N_19943);
nand UO_1916 (O_1916,N_19864,N_19989);
nand UO_1917 (O_1917,N_19986,N_19851);
xor UO_1918 (O_1918,N_19879,N_19914);
or UO_1919 (O_1919,N_19968,N_19958);
nor UO_1920 (O_1920,N_19940,N_19834);
nor UO_1921 (O_1921,N_19963,N_19947);
nor UO_1922 (O_1922,N_19990,N_19882);
nand UO_1923 (O_1923,N_19850,N_19946);
and UO_1924 (O_1924,N_19967,N_19916);
xnor UO_1925 (O_1925,N_19863,N_19893);
nand UO_1926 (O_1926,N_19813,N_19942);
xnor UO_1927 (O_1927,N_19822,N_19862);
nor UO_1928 (O_1928,N_19811,N_19983);
nand UO_1929 (O_1929,N_19848,N_19870);
nand UO_1930 (O_1930,N_19858,N_19862);
and UO_1931 (O_1931,N_19812,N_19972);
xor UO_1932 (O_1932,N_19958,N_19925);
and UO_1933 (O_1933,N_19847,N_19968);
xor UO_1934 (O_1934,N_19830,N_19856);
or UO_1935 (O_1935,N_19997,N_19970);
and UO_1936 (O_1936,N_19951,N_19901);
nand UO_1937 (O_1937,N_19872,N_19914);
nand UO_1938 (O_1938,N_19810,N_19968);
or UO_1939 (O_1939,N_19991,N_19946);
nor UO_1940 (O_1940,N_19867,N_19971);
and UO_1941 (O_1941,N_19969,N_19856);
nand UO_1942 (O_1942,N_19897,N_19904);
or UO_1943 (O_1943,N_19936,N_19833);
or UO_1944 (O_1944,N_19996,N_19948);
nor UO_1945 (O_1945,N_19938,N_19861);
xnor UO_1946 (O_1946,N_19850,N_19993);
and UO_1947 (O_1947,N_19999,N_19882);
and UO_1948 (O_1948,N_19911,N_19824);
nor UO_1949 (O_1949,N_19805,N_19807);
and UO_1950 (O_1950,N_19800,N_19864);
xor UO_1951 (O_1951,N_19957,N_19980);
and UO_1952 (O_1952,N_19851,N_19935);
nor UO_1953 (O_1953,N_19952,N_19827);
or UO_1954 (O_1954,N_19816,N_19860);
nand UO_1955 (O_1955,N_19849,N_19998);
nor UO_1956 (O_1956,N_19837,N_19819);
nand UO_1957 (O_1957,N_19907,N_19922);
and UO_1958 (O_1958,N_19924,N_19900);
nand UO_1959 (O_1959,N_19947,N_19958);
and UO_1960 (O_1960,N_19904,N_19806);
nor UO_1961 (O_1961,N_19810,N_19936);
and UO_1962 (O_1962,N_19998,N_19966);
and UO_1963 (O_1963,N_19932,N_19853);
and UO_1964 (O_1964,N_19875,N_19996);
xnor UO_1965 (O_1965,N_19959,N_19980);
or UO_1966 (O_1966,N_19812,N_19862);
nor UO_1967 (O_1967,N_19939,N_19928);
and UO_1968 (O_1968,N_19882,N_19845);
nor UO_1969 (O_1969,N_19946,N_19824);
nor UO_1970 (O_1970,N_19890,N_19841);
or UO_1971 (O_1971,N_19935,N_19982);
xor UO_1972 (O_1972,N_19814,N_19861);
xnor UO_1973 (O_1973,N_19868,N_19832);
nor UO_1974 (O_1974,N_19971,N_19959);
nor UO_1975 (O_1975,N_19941,N_19916);
nor UO_1976 (O_1976,N_19876,N_19868);
nor UO_1977 (O_1977,N_19967,N_19888);
nand UO_1978 (O_1978,N_19967,N_19952);
nand UO_1979 (O_1979,N_19821,N_19841);
and UO_1980 (O_1980,N_19875,N_19837);
nor UO_1981 (O_1981,N_19925,N_19935);
and UO_1982 (O_1982,N_19990,N_19989);
nor UO_1983 (O_1983,N_19802,N_19869);
and UO_1984 (O_1984,N_19914,N_19885);
xnor UO_1985 (O_1985,N_19957,N_19861);
and UO_1986 (O_1986,N_19809,N_19852);
nand UO_1987 (O_1987,N_19949,N_19835);
nor UO_1988 (O_1988,N_19998,N_19912);
nand UO_1989 (O_1989,N_19956,N_19869);
xor UO_1990 (O_1990,N_19969,N_19930);
nor UO_1991 (O_1991,N_19891,N_19808);
nand UO_1992 (O_1992,N_19816,N_19881);
and UO_1993 (O_1993,N_19820,N_19861);
nor UO_1994 (O_1994,N_19869,N_19955);
nor UO_1995 (O_1995,N_19908,N_19940);
nor UO_1996 (O_1996,N_19841,N_19845);
nor UO_1997 (O_1997,N_19852,N_19882);
nor UO_1998 (O_1998,N_19880,N_19930);
or UO_1999 (O_1999,N_19837,N_19801);
or UO_2000 (O_2000,N_19884,N_19948);
or UO_2001 (O_2001,N_19955,N_19922);
nand UO_2002 (O_2002,N_19849,N_19861);
nand UO_2003 (O_2003,N_19803,N_19927);
xnor UO_2004 (O_2004,N_19994,N_19944);
nor UO_2005 (O_2005,N_19828,N_19841);
nor UO_2006 (O_2006,N_19876,N_19828);
xor UO_2007 (O_2007,N_19965,N_19812);
xnor UO_2008 (O_2008,N_19837,N_19890);
or UO_2009 (O_2009,N_19855,N_19851);
xnor UO_2010 (O_2010,N_19819,N_19825);
and UO_2011 (O_2011,N_19832,N_19942);
or UO_2012 (O_2012,N_19880,N_19848);
nand UO_2013 (O_2013,N_19849,N_19940);
nor UO_2014 (O_2014,N_19904,N_19951);
and UO_2015 (O_2015,N_19823,N_19889);
or UO_2016 (O_2016,N_19809,N_19982);
nand UO_2017 (O_2017,N_19851,N_19861);
xor UO_2018 (O_2018,N_19850,N_19906);
nand UO_2019 (O_2019,N_19871,N_19820);
xnor UO_2020 (O_2020,N_19811,N_19924);
nand UO_2021 (O_2021,N_19986,N_19894);
and UO_2022 (O_2022,N_19814,N_19889);
nor UO_2023 (O_2023,N_19895,N_19870);
xor UO_2024 (O_2024,N_19891,N_19979);
nor UO_2025 (O_2025,N_19921,N_19895);
and UO_2026 (O_2026,N_19872,N_19801);
or UO_2027 (O_2027,N_19872,N_19874);
or UO_2028 (O_2028,N_19910,N_19852);
xnor UO_2029 (O_2029,N_19976,N_19898);
xnor UO_2030 (O_2030,N_19938,N_19860);
or UO_2031 (O_2031,N_19838,N_19952);
and UO_2032 (O_2032,N_19993,N_19965);
and UO_2033 (O_2033,N_19949,N_19911);
nand UO_2034 (O_2034,N_19830,N_19988);
nand UO_2035 (O_2035,N_19963,N_19844);
nand UO_2036 (O_2036,N_19846,N_19842);
xnor UO_2037 (O_2037,N_19896,N_19831);
and UO_2038 (O_2038,N_19962,N_19884);
nor UO_2039 (O_2039,N_19857,N_19819);
or UO_2040 (O_2040,N_19881,N_19896);
nand UO_2041 (O_2041,N_19909,N_19821);
or UO_2042 (O_2042,N_19859,N_19801);
xnor UO_2043 (O_2043,N_19975,N_19803);
nor UO_2044 (O_2044,N_19932,N_19924);
nand UO_2045 (O_2045,N_19806,N_19841);
nor UO_2046 (O_2046,N_19998,N_19823);
nand UO_2047 (O_2047,N_19957,N_19988);
nor UO_2048 (O_2048,N_19879,N_19837);
nand UO_2049 (O_2049,N_19976,N_19857);
nor UO_2050 (O_2050,N_19952,N_19847);
nand UO_2051 (O_2051,N_19857,N_19878);
or UO_2052 (O_2052,N_19921,N_19908);
nor UO_2053 (O_2053,N_19993,N_19807);
or UO_2054 (O_2054,N_19832,N_19888);
xnor UO_2055 (O_2055,N_19844,N_19912);
or UO_2056 (O_2056,N_19810,N_19868);
xnor UO_2057 (O_2057,N_19891,N_19921);
xor UO_2058 (O_2058,N_19920,N_19952);
or UO_2059 (O_2059,N_19935,N_19931);
and UO_2060 (O_2060,N_19994,N_19907);
and UO_2061 (O_2061,N_19940,N_19872);
nand UO_2062 (O_2062,N_19915,N_19955);
xnor UO_2063 (O_2063,N_19837,N_19814);
or UO_2064 (O_2064,N_19923,N_19845);
or UO_2065 (O_2065,N_19983,N_19902);
or UO_2066 (O_2066,N_19858,N_19845);
nand UO_2067 (O_2067,N_19823,N_19967);
or UO_2068 (O_2068,N_19906,N_19888);
nand UO_2069 (O_2069,N_19996,N_19944);
xnor UO_2070 (O_2070,N_19825,N_19967);
nand UO_2071 (O_2071,N_19895,N_19955);
nand UO_2072 (O_2072,N_19980,N_19802);
or UO_2073 (O_2073,N_19874,N_19901);
nor UO_2074 (O_2074,N_19935,N_19977);
and UO_2075 (O_2075,N_19908,N_19849);
or UO_2076 (O_2076,N_19834,N_19988);
nand UO_2077 (O_2077,N_19922,N_19818);
nor UO_2078 (O_2078,N_19953,N_19984);
xnor UO_2079 (O_2079,N_19940,N_19858);
or UO_2080 (O_2080,N_19928,N_19970);
nand UO_2081 (O_2081,N_19802,N_19837);
or UO_2082 (O_2082,N_19935,N_19923);
nand UO_2083 (O_2083,N_19877,N_19852);
nand UO_2084 (O_2084,N_19995,N_19826);
nor UO_2085 (O_2085,N_19843,N_19871);
nor UO_2086 (O_2086,N_19877,N_19920);
or UO_2087 (O_2087,N_19840,N_19856);
xor UO_2088 (O_2088,N_19878,N_19877);
and UO_2089 (O_2089,N_19979,N_19869);
or UO_2090 (O_2090,N_19863,N_19853);
or UO_2091 (O_2091,N_19915,N_19903);
nand UO_2092 (O_2092,N_19873,N_19988);
xor UO_2093 (O_2093,N_19851,N_19994);
or UO_2094 (O_2094,N_19895,N_19948);
nor UO_2095 (O_2095,N_19866,N_19910);
and UO_2096 (O_2096,N_19999,N_19822);
or UO_2097 (O_2097,N_19885,N_19867);
nand UO_2098 (O_2098,N_19847,N_19901);
or UO_2099 (O_2099,N_19943,N_19982);
nor UO_2100 (O_2100,N_19998,N_19886);
nor UO_2101 (O_2101,N_19849,N_19957);
nand UO_2102 (O_2102,N_19824,N_19812);
nand UO_2103 (O_2103,N_19844,N_19862);
and UO_2104 (O_2104,N_19808,N_19986);
and UO_2105 (O_2105,N_19928,N_19922);
or UO_2106 (O_2106,N_19935,N_19934);
nor UO_2107 (O_2107,N_19867,N_19833);
and UO_2108 (O_2108,N_19800,N_19819);
or UO_2109 (O_2109,N_19831,N_19864);
nor UO_2110 (O_2110,N_19854,N_19904);
nand UO_2111 (O_2111,N_19866,N_19972);
xnor UO_2112 (O_2112,N_19904,N_19873);
or UO_2113 (O_2113,N_19901,N_19921);
nand UO_2114 (O_2114,N_19837,N_19838);
nand UO_2115 (O_2115,N_19996,N_19960);
and UO_2116 (O_2116,N_19863,N_19834);
and UO_2117 (O_2117,N_19819,N_19889);
nor UO_2118 (O_2118,N_19933,N_19936);
and UO_2119 (O_2119,N_19903,N_19943);
nor UO_2120 (O_2120,N_19859,N_19834);
nor UO_2121 (O_2121,N_19957,N_19960);
xor UO_2122 (O_2122,N_19812,N_19973);
nand UO_2123 (O_2123,N_19981,N_19969);
nand UO_2124 (O_2124,N_19911,N_19984);
nor UO_2125 (O_2125,N_19826,N_19908);
xor UO_2126 (O_2126,N_19823,N_19954);
nor UO_2127 (O_2127,N_19862,N_19931);
or UO_2128 (O_2128,N_19929,N_19907);
xnor UO_2129 (O_2129,N_19910,N_19823);
nor UO_2130 (O_2130,N_19888,N_19846);
xnor UO_2131 (O_2131,N_19811,N_19898);
nand UO_2132 (O_2132,N_19944,N_19909);
and UO_2133 (O_2133,N_19841,N_19829);
nor UO_2134 (O_2134,N_19873,N_19939);
and UO_2135 (O_2135,N_19917,N_19960);
nor UO_2136 (O_2136,N_19937,N_19934);
xnor UO_2137 (O_2137,N_19982,N_19845);
nand UO_2138 (O_2138,N_19987,N_19913);
xor UO_2139 (O_2139,N_19986,N_19970);
or UO_2140 (O_2140,N_19810,N_19844);
nor UO_2141 (O_2141,N_19814,N_19867);
and UO_2142 (O_2142,N_19802,N_19840);
and UO_2143 (O_2143,N_19800,N_19889);
or UO_2144 (O_2144,N_19942,N_19924);
xor UO_2145 (O_2145,N_19804,N_19864);
nand UO_2146 (O_2146,N_19868,N_19926);
xor UO_2147 (O_2147,N_19920,N_19997);
nor UO_2148 (O_2148,N_19952,N_19922);
nand UO_2149 (O_2149,N_19936,N_19930);
or UO_2150 (O_2150,N_19920,N_19965);
and UO_2151 (O_2151,N_19964,N_19857);
or UO_2152 (O_2152,N_19812,N_19835);
or UO_2153 (O_2153,N_19995,N_19818);
or UO_2154 (O_2154,N_19826,N_19966);
and UO_2155 (O_2155,N_19908,N_19804);
nor UO_2156 (O_2156,N_19870,N_19861);
nand UO_2157 (O_2157,N_19996,N_19935);
nand UO_2158 (O_2158,N_19970,N_19974);
or UO_2159 (O_2159,N_19947,N_19817);
xnor UO_2160 (O_2160,N_19925,N_19894);
or UO_2161 (O_2161,N_19800,N_19987);
nor UO_2162 (O_2162,N_19869,N_19861);
nand UO_2163 (O_2163,N_19843,N_19955);
and UO_2164 (O_2164,N_19813,N_19894);
nor UO_2165 (O_2165,N_19898,N_19858);
or UO_2166 (O_2166,N_19801,N_19852);
or UO_2167 (O_2167,N_19966,N_19994);
or UO_2168 (O_2168,N_19979,N_19977);
nor UO_2169 (O_2169,N_19887,N_19908);
nand UO_2170 (O_2170,N_19899,N_19966);
or UO_2171 (O_2171,N_19931,N_19902);
nand UO_2172 (O_2172,N_19825,N_19838);
xor UO_2173 (O_2173,N_19998,N_19994);
and UO_2174 (O_2174,N_19999,N_19820);
xnor UO_2175 (O_2175,N_19943,N_19925);
or UO_2176 (O_2176,N_19887,N_19975);
nand UO_2177 (O_2177,N_19876,N_19930);
and UO_2178 (O_2178,N_19897,N_19852);
or UO_2179 (O_2179,N_19859,N_19939);
and UO_2180 (O_2180,N_19964,N_19914);
nand UO_2181 (O_2181,N_19918,N_19807);
and UO_2182 (O_2182,N_19910,N_19819);
xor UO_2183 (O_2183,N_19911,N_19899);
xor UO_2184 (O_2184,N_19861,N_19920);
xor UO_2185 (O_2185,N_19969,N_19884);
or UO_2186 (O_2186,N_19834,N_19948);
xnor UO_2187 (O_2187,N_19941,N_19952);
xnor UO_2188 (O_2188,N_19841,N_19963);
or UO_2189 (O_2189,N_19820,N_19872);
nand UO_2190 (O_2190,N_19874,N_19908);
nand UO_2191 (O_2191,N_19917,N_19943);
nor UO_2192 (O_2192,N_19804,N_19913);
xnor UO_2193 (O_2193,N_19972,N_19941);
nand UO_2194 (O_2194,N_19840,N_19950);
or UO_2195 (O_2195,N_19838,N_19924);
xnor UO_2196 (O_2196,N_19932,N_19897);
xor UO_2197 (O_2197,N_19946,N_19996);
and UO_2198 (O_2198,N_19828,N_19924);
or UO_2199 (O_2199,N_19807,N_19867);
nor UO_2200 (O_2200,N_19980,N_19932);
or UO_2201 (O_2201,N_19864,N_19907);
and UO_2202 (O_2202,N_19921,N_19832);
nor UO_2203 (O_2203,N_19829,N_19927);
nor UO_2204 (O_2204,N_19942,N_19856);
nand UO_2205 (O_2205,N_19963,N_19998);
or UO_2206 (O_2206,N_19836,N_19870);
nand UO_2207 (O_2207,N_19946,N_19947);
and UO_2208 (O_2208,N_19883,N_19860);
nor UO_2209 (O_2209,N_19813,N_19895);
and UO_2210 (O_2210,N_19879,N_19873);
nand UO_2211 (O_2211,N_19978,N_19935);
xnor UO_2212 (O_2212,N_19986,N_19988);
xnor UO_2213 (O_2213,N_19954,N_19804);
or UO_2214 (O_2214,N_19861,N_19993);
nor UO_2215 (O_2215,N_19864,N_19926);
and UO_2216 (O_2216,N_19954,N_19854);
and UO_2217 (O_2217,N_19887,N_19942);
nor UO_2218 (O_2218,N_19925,N_19814);
xnor UO_2219 (O_2219,N_19904,N_19871);
xnor UO_2220 (O_2220,N_19988,N_19900);
nor UO_2221 (O_2221,N_19819,N_19973);
nand UO_2222 (O_2222,N_19830,N_19970);
xor UO_2223 (O_2223,N_19873,N_19847);
and UO_2224 (O_2224,N_19894,N_19929);
xnor UO_2225 (O_2225,N_19936,N_19805);
xnor UO_2226 (O_2226,N_19816,N_19817);
nor UO_2227 (O_2227,N_19928,N_19992);
nand UO_2228 (O_2228,N_19910,N_19811);
or UO_2229 (O_2229,N_19928,N_19918);
and UO_2230 (O_2230,N_19857,N_19813);
nand UO_2231 (O_2231,N_19922,N_19900);
nand UO_2232 (O_2232,N_19877,N_19829);
and UO_2233 (O_2233,N_19999,N_19880);
nor UO_2234 (O_2234,N_19899,N_19819);
or UO_2235 (O_2235,N_19859,N_19928);
xnor UO_2236 (O_2236,N_19865,N_19807);
xor UO_2237 (O_2237,N_19838,N_19909);
or UO_2238 (O_2238,N_19957,N_19882);
or UO_2239 (O_2239,N_19975,N_19960);
nor UO_2240 (O_2240,N_19841,N_19804);
or UO_2241 (O_2241,N_19891,N_19851);
xor UO_2242 (O_2242,N_19922,N_19888);
and UO_2243 (O_2243,N_19998,N_19920);
nand UO_2244 (O_2244,N_19900,N_19867);
and UO_2245 (O_2245,N_19800,N_19969);
and UO_2246 (O_2246,N_19905,N_19833);
nor UO_2247 (O_2247,N_19885,N_19812);
or UO_2248 (O_2248,N_19832,N_19981);
and UO_2249 (O_2249,N_19811,N_19959);
or UO_2250 (O_2250,N_19915,N_19946);
and UO_2251 (O_2251,N_19986,N_19903);
xnor UO_2252 (O_2252,N_19999,N_19855);
nand UO_2253 (O_2253,N_19819,N_19994);
and UO_2254 (O_2254,N_19901,N_19940);
nand UO_2255 (O_2255,N_19970,N_19939);
or UO_2256 (O_2256,N_19891,N_19918);
xor UO_2257 (O_2257,N_19946,N_19873);
xor UO_2258 (O_2258,N_19851,N_19863);
xor UO_2259 (O_2259,N_19945,N_19844);
nand UO_2260 (O_2260,N_19929,N_19900);
nand UO_2261 (O_2261,N_19967,N_19948);
xnor UO_2262 (O_2262,N_19925,N_19898);
nor UO_2263 (O_2263,N_19811,N_19993);
nor UO_2264 (O_2264,N_19974,N_19925);
nand UO_2265 (O_2265,N_19920,N_19940);
nor UO_2266 (O_2266,N_19941,N_19919);
nor UO_2267 (O_2267,N_19936,N_19851);
xnor UO_2268 (O_2268,N_19815,N_19845);
nand UO_2269 (O_2269,N_19855,N_19951);
xnor UO_2270 (O_2270,N_19809,N_19837);
and UO_2271 (O_2271,N_19980,N_19956);
and UO_2272 (O_2272,N_19997,N_19977);
nor UO_2273 (O_2273,N_19963,N_19875);
nand UO_2274 (O_2274,N_19954,N_19906);
or UO_2275 (O_2275,N_19978,N_19869);
and UO_2276 (O_2276,N_19866,N_19948);
nor UO_2277 (O_2277,N_19837,N_19831);
nand UO_2278 (O_2278,N_19995,N_19998);
xor UO_2279 (O_2279,N_19807,N_19891);
xor UO_2280 (O_2280,N_19937,N_19943);
nand UO_2281 (O_2281,N_19921,N_19911);
xnor UO_2282 (O_2282,N_19828,N_19853);
xor UO_2283 (O_2283,N_19918,N_19935);
nand UO_2284 (O_2284,N_19831,N_19959);
nor UO_2285 (O_2285,N_19998,N_19852);
nand UO_2286 (O_2286,N_19936,N_19895);
or UO_2287 (O_2287,N_19907,N_19840);
and UO_2288 (O_2288,N_19806,N_19820);
nand UO_2289 (O_2289,N_19900,N_19863);
nand UO_2290 (O_2290,N_19846,N_19865);
nor UO_2291 (O_2291,N_19878,N_19986);
and UO_2292 (O_2292,N_19987,N_19896);
nand UO_2293 (O_2293,N_19805,N_19966);
or UO_2294 (O_2294,N_19805,N_19944);
and UO_2295 (O_2295,N_19972,N_19986);
xor UO_2296 (O_2296,N_19984,N_19857);
nor UO_2297 (O_2297,N_19845,N_19993);
xor UO_2298 (O_2298,N_19967,N_19954);
xnor UO_2299 (O_2299,N_19879,N_19971);
nor UO_2300 (O_2300,N_19876,N_19854);
or UO_2301 (O_2301,N_19978,N_19946);
xor UO_2302 (O_2302,N_19940,N_19877);
nor UO_2303 (O_2303,N_19831,N_19962);
xor UO_2304 (O_2304,N_19926,N_19817);
and UO_2305 (O_2305,N_19886,N_19940);
nor UO_2306 (O_2306,N_19800,N_19988);
or UO_2307 (O_2307,N_19933,N_19945);
nand UO_2308 (O_2308,N_19957,N_19978);
nand UO_2309 (O_2309,N_19948,N_19818);
xor UO_2310 (O_2310,N_19968,N_19885);
and UO_2311 (O_2311,N_19835,N_19886);
nor UO_2312 (O_2312,N_19982,N_19874);
nor UO_2313 (O_2313,N_19987,N_19888);
xnor UO_2314 (O_2314,N_19926,N_19982);
xnor UO_2315 (O_2315,N_19883,N_19885);
or UO_2316 (O_2316,N_19928,N_19956);
xor UO_2317 (O_2317,N_19864,N_19967);
and UO_2318 (O_2318,N_19905,N_19973);
nand UO_2319 (O_2319,N_19914,N_19811);
nand UO_2320 (O_2320,N_19927,N_19909);
nand UO_2321 (O_2321,N_19855,N_19819);
nor UO_2322 (O_2322,N_19834,N_19857);
nor UO_2323 (O_2323,N_19872,N_19813);
or UO_2324 (O_2324,N_19995,N_19987);
and UO_2325 (O_2325,N_19923,N_19904);
and UO_2326 (O_2326,N_19844,N_19985);
xnor UO_2327 (O_2327,N_19967,N_19889);
and UO_2328 (O_2328,N_19867,N_19961);
and UO_2329 (O_2329,N_19995,N_19931);
nor UO_2330 (O_2330,N_19990,N_19928);
and UO_2331 (O_2331,N_19953,N_19922);
nor UO_2332 (O_2332,N_19960,N_19908);
or UO_2333 (O_2333,N_19945,N_19804);
nor UO_2334 (O_2334,N_19914,N_19949);
nor UO_2335 (O_2335,N_19891,N_19882);
nor UO_2336 (O_2336,N_19960,N_19944);
xnor UO_2337 (O_2337,N_19918,N_19912);
nor UO_2338 (O_2338,N_19913,N_19977);
or UO_2339 (O_2339,N_19803,N_19806);
xnor UO_2340 (O_2340,N_19805,N_19941);
nand UO_2341 (O_2341,N_19815,N_19972);
or UO_2342 (O_2342,N_19934,N_19810);
xor UO_2343 (O_2343,N_19866,N_19919);
or UO_2344 (O_2344,N_19886,N_19891);
and UO_2345 (O_2345,N_19962,N_19915);
and UO_2346 (O_2346,N_19914,N_19853);
or UO_2347 (O_2347,N_19932,N_19866);
nand UO_2348 (O_2348,N_19963,N_19933);
nand UO_2349 (O_2349,N_19882,N_19889);
nor UO_2350 (O_2350,N_19820,N_19829);
xnor UO_2351 (O_2351,N_19845,N_19908);
nand UO_2352 (O_2352,N_19931,N_19836);
xor UO_2353 (O_2353,N_19954,N_19925);
nand UO_2354 (O_2354,N_19862,N_19870);
and UO_2355 (O_2355,N_19854,N_19820);
and UO_2356 (O_2356,N_19826,N_19823);
nor UO_2357 (O_2357,N_19936,N_19960);
nor UO_2358 (O_2358,N_19899,N_19967);
nor UO_2359 (O_2359,N_19939,N_19854);
and UO_2360 (O_2360,N_19814,N_19904);
nand UO_2361 (O_2361,N_19990,N_19869);
or UO_2362 (O_2362,N_19963,N_19874);
nor UO_2363 (O_2363,N_19886,N_19812);
or UO_2364 (O_2364,N_19939,N_19834);
and UO_2365 (O_2365,N_19942,N_19925);
xor UO_2366 (O_2366,N_19897,N_19981);
nand UO_2367 (O_2367,N_19881,N_19843);
nor UO_2368 (O_2368,N_19893,N_19858);
nor UO_2369 (O_2369,N_19903,N_19977);
nor UO_2370 (O_2370,N_19994,N_19880);
xnor UO_2371 (O_2371,N_19895,N_19874);
or UO_2372 (O_2372,N_19917,N_19967);
nand UO_2373 (O_2373,N_19898,N_19903);
and UO_2374 (O_2374,N_19927,N_19963);
xnor UO_2375 (O_2375,N_19896,N_19931);
nor UO_2376 (O_2376,N_19841,N_19968);
nand UO_2377 (O_2377,N_19832,N_19859);
nand UO_2378 (O_2378,N_19806,N_19897);
or UO_2379 (O_2379,N_19834,N_19905);
xor UO_2380 (O_2380,N_19920,N_19881);
or UO_2381 (O_2381,N_19896,N_19978);
or UO_2382 (O_2382,N_19895,N_19915);
nor UO_2383 (O_2383,N_19923,N_19937);
xnor UO_2384 (O_2384,N_19987,N_19851);
nand UO_2385 (O_2385,N_19812,N_19962);
nor UO_2386 (O_2386,N_19994,N_19883);
and UO_2387 (O_2387,N_19851,N_19882);
xor UO_2388 (O_2388,N_19986,N_19942);
xnor UO_2389 (O_2389,N_19924,N_19847);
or UO_2390 (O_2390,N_19848,N_19810);
nor UO_2391 (O_2391,N_19896,N_19823);
or UO_2392 (O_2392,N_19801,N_19814);
or UO_2393 (O_2393,N_19894,N_19865);
xor UO_2394 (O_2394,N_19929,N_19841);
nor UO_2395 (O_2395,N_19829,N_19993);
nor UO_2396 (O_2396,N_19999,N_19975);
xor UO_2397 (O_2397,N_19897,N_19823);
or UO_2398 (O_2398,N_19975,N_19878);
or UO_2399 (O_2399,N_19809,N_19988);
nand UO_2400 (O_2400,N_19917,N_19927);
xnor UO_2401 (O_2401,N_19809,N_19915);
or UO_2402 (O_2402,N_19985,N_19879);
or UO_2403 (O_2403,N_19806,N_19817);
and UO_2404 (O_2404,N_19973,N_19996);
xnor UO_2405 (O_2405,N_19826,N_19847);
or UO_2406 (O_2406,N_19847,N_19811);
nor UO_2407 (O_2407,N_19906,N_19838);
and UO_2408 (O_2408,N_19821,N_19955);
nor UO_2409 (O_2409,N_19870,N_19892);
nand UO_2410 (O_2410,N_19967,N_19908);
and UO_2411 (O_2411,N_19855,N_19897);
nor UO_2412 (O_2412,N_19863,N_19906);
and UO_2413 (O_2413,N_19818,N_19836);
xor UO_2414 (O_2414,N_19888,N_19961);
or UO_2415 (O_2415,N_19951,N_19983);
or UO_2416 (O_2416,N_19862,N_19890);
or UO_2417 (O_2417,N_19995,N_19911);
or UO_2418 (O_2418,N_19989,N_19931);
or UO_2419 (O_2419,N_19808,N_19890);
xnor UO_2420 (O_2420,N_19885,N_19934);
or UO_2421 (O_2421,N_19831,N_19973);
nor UO_2422 (O_2422,N_19806,N_19929);
nor UO_2423 (O_2423,N_19994,N_19868);
nand UO_2424 (O_2424,N_19925,N_19884);
and UO_2425 (O_2425,N_19940,N_19866);
xnor UO_2426 (O_2426,N_19801,N_19817);
nor UO_2427 (O_2427,N_19826,N_19865);
nand UO_2428 (O_2428,N_19978,N_19889);
or UO_2429 (O_2429,N_19806,N_19914);
xor UO_2430 (O_2430,N_19890,N_19914);
nor UO_2431 (O_2431,N_19839,N_19867);
and UO_2432 (O_2432,N_19815,N_19854);
nand UO_2433 (O_2433,N_19886,N_19814);
and UO_2434 (O_2434,N_19938,N_19898);
or UO_2435 (O_2435,N_19804,N_19899);
and UO_2436 (O_2436,N_19858,N_19970);
and UO_2437 (O_2437,N_19823,N_19905);
or UO_2438 (O_2438,N_19853,N_19989);
xor UO_2439 (O_2439,N_19869,N_19915);
nor UO_2440 (O_2440,N_19937,N_19858);
and UO_2441 (O_2441,N_19892,N_19859);
xnor UO_2442 (O_2442,N_19835,N_19967);
xnor UO_2443 (O_2443,N_19892,N_19926);
nand UO_2444 (O_2444,N_19965,N_19952);
nand UO_2445 (O_2445,N_19810,N_19938);
nand UO_2446 (O_2446,N_19899,N_19963);
and UO_2447 (O_2447,N_19929,N_19846);
and UO_2448 (O_2448,N_19815,N_19978);
and UO_2449 (O_2449,N_19805,N_19916);
nor UO_2450 (O_2450,N_19987,N_19950);
nand UO_2451 (O_2451,N_19877,N_19897);
and UO_2452 (O_2452,N_19902,N_19908);
and UO_2453 (O_2453,N_19925,N_19882);
nor UO_2454 (O_2454,N_19825,N_19832);
nand UO_2455 (O_2455,N_19877,N_19864);
or UO_2456 (O_2456,N_19922,N_19920);
nor UO_2457 (O_2457,N_19873,N_19893);
or UO_2458 (O_2458,N_19900,N_19898);
nor UO_2459 (O_2459,N_19828,N_19821);
nor UO_2460 (O_2460,N_19970,N_19985);
nand UO_2461 (O_2461,N_19871,N_19977);
xnor UO_2462 (O_2462,N_19923,N_19877);
or UO_2463 (O_2463,N_19916,N_19982);
and UO_2464 (O_2464,N_19985,N_19920);
or UO_2465 (O_2465,N_19870,N_19828);
or UO_2466 (O_2466,N_19821,N_19855);
and UO_2467 (O_2467,N_19974,N_19896);
and UO_2468 (O_2468,N_19861,N_19817);
and UO_2469 (O_2469,N_19870,N_19869);
xnor UO_2470 (O_2470,N_19977,N_19808);
and UO_2471 (O_2471,N_19920,N_19876);
or UO_2472 (O_2472,N_19936,N_19837);
and UO_2473 (O_2473,N_19926,N_19981);
xnor UO_2474 (O_2474,N_19846,N_19994);
and UO_2475 (O_2475,N_19835,N_19947);
xor UO_2476 (O_2476,N_19860,N_19864);
xor UO_2477 (O_2477,N_19881,N_19932);
xnor UO_2478 (O_2478,N_19977,N_19845);
nand UO_2479 (O_2479,N_19837,N_19859);
and UO_2480 (O_2480,N_19809,N_19892);
nor UO_2481 (O_2481,N_19807,N_19825);
xor UO_2482 (O_2482,N_19997,N_19905);
or UO_2483 (O_2483,N_19905,N_19953);
and UO_2484 (O_2484,N_19928,N_19911);
nand UO_2485 (O_2485,N_19853,N_19947);
or UO_2486 (O_2486,N_19872,N_19899);
and UO_2487 (O_2487,N_19928,N_19899);
or UO_2488 (O_2488,N_19883,N_19923);
xnor UO_2489 (O_2489,N_19947,N_19983);
nor UO_2490 (O_2490,N_19858,N_19901);
xnor UO_2491 (O_2491,N_19985,N_19968);
or UO_2492 (O_2492,N_19969,N_19867);
xor UO_2493 (O_2493,N_19841,N_19984);
nand UO_2494 (O_2494,N_19878,N_19957);
and UO_2495 (O_2495,N_19996,N_19950);
and UO_2496 (O_2496,N_19839,N_19968);
and UO_2497 (O_2497,N_19887,N_19964);
nor UO_2498 (O_2498,N_19876,N_19842);
xor UO_2499 (O_2499,N_19976,N_19880);
endmodule