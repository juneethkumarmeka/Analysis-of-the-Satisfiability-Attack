module basic_500_3000_500_5_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_371,In_444);
xor U1 (N_1,In_75,In_415);
nand U2 (N_2,In_443,In_489);
nor U3 (N_3,In_67,In_327);
or U4 (N_4,In_181,In_49);
nand U5 (N_5,In_141,In_457);
nor U6 (N_6,In_143,In_122);
or U7 (N_7,In_78,In_442);
or U8 (N_8,In_179,In_365);
nor U9 (N_9,In_171,In_2);
or U10 (N_10,In_211,In_379);
or U11 (N_11,In_302,In_445);
nand U12 (N_12,In_128,In_50);
xor U13 (N_13,In_285,In_293);
nand U14 (N_14,In_0,In_334);
nand U15 (N_15,In_27,In_235);
nand U16 (N_16,In_324,In_167);
nand U17 (N_17,In_116,In_155);
nor U18 (N_18,In_372,In_418);
or U19 (N_19,In_483,In_45);
nor U20 (N_20,In_97,In_219);
and U21 (N_21,In_168,In_383);
or U22 (N_22,In_195,In_103);
nor U23 (N_23,In_190,In_300);
nor U24 (N_24,In_189,In_298);
xnor U25 (N_25,In_255,In_478);
or U26 (N_26,In_311,In_290);
nor U27 (N_27,In_209,In_173);
or U28 (N_28,In_362,In_391);
or U29 (N_29,In_140,In_249);
nand U30 (N_30,In_339,In_191);
or U31 (N_31,In_412,In_257);
nor U32 (N_32,In_46,In_403);
and U33 (N_33,In_107,In_109);
nand U34 (N_34,In_20,In_366);
nor U35 (N_35,In_259,In_69);
and U36 (N_36,In_175,In_202);
nand U37 (N_37,In_388,In_204);
xnor U38 (N_38,In_14,In_454);
and U39 (N_39,In_91,In_121);
nor U40 (N_40,In_41,In_342);
nand U41 (N_41,In_270,In_26);
nor U42 (N_42,In_263,In_356);
or U43 (N_43,In_315,In_410);
nor U44 (N_44,In_15,In_110);
and U45 (N_45,In_199,In_353);
and U46 (N_46,In_495,In_449);
or U47 (N_47,In_258,In_9);
nor U48 (N_48,In_446,In_299);
nor U49 (N_49,In_100,In_177);
or U50 (N_50,In_486,In_36);
nor U51 (N_51,In_289,In_321);
and U52 (N_52,In_44,In_10);
or U53 (N_53,In_294,In_174);
or U54 (N_54,In_22,In_104);
nand U55 (N_55,In_431,In_276);
nand U56 (N_56,In_316,In_292);
or U57 (N_57,In_3,In_248);
or U58 (N_58,In_402,In_164);
nand U59 (N_59,In_262,In_134);
nand U60 (N_60,In_212,In_384);
and U61 (N_61,In_268,In_435);
nor U62 (N_62,In_367,In_360);
and U63 (N_63,In_480,In_198);
or U64 (N_64,In_222,In_196);
and U65 (N_65,In_393,In_35);
nor U66 (N_66,In_266,In_398);
or U67 (N_67,In_18,In_423);
nand U68 (N_68,In_139,In_4);
and U69 (N_69,In_210,In_7);
and U70 (N_70,In_172,In_207);
nand U71 (N_71,In_129,In_80);
and U72 (N_72,In_326,In_317);
and U73 (N_73,In_216,In_83);
nor U74 (N_74,In_162,In_484);
or U75 (N_75,In_193,In_377);
or U76 (N_76,In_272,In_427);
xor U77 (N_77,In_253,In_331);
nor U78 (N_78,In_381,In_126);
xor U79 (N_79,In_346,In_21);
xor U80 (N_80,In_429,In_250);
nor U81 (N_81,In_369,In_71);
xnor U82 (N_82,In_341,In_386);
nor U83 (N_83,In_245,In_413);
nor U84 (N_84,In_70,In_147);
or U85 (N_85,In_284,In_434);
nand U86 (N_86,In_430,In_425);
or U87 (N_87,In_424,In_62);
nor U88 (N_88,In_467,In_240);
and U89 (N_89,In_53,In_90);
or U90 (N_90,In_187,In_12);
or U91 (N_91,In_477,In_405);
or U92 (N_92,In_120,In_251);
or U93 (N_93,In_400,In_458);
nand U94 (N_94,In_448,In_254);
nor U95 (N_95,In_479,In_114);
nor U96 (N_96,In_395,In_460);
or U97 (N_97,In_355,In_416);
and U98 (N_98,In_345,In_124);
xor U99 (N_99,In_323,In_73);
or U100 (N_100,In_309,In_34);
xor U101 (N_101,In_82,In_176);
and U102 (N_102,In_488,In_374);
or U103 (N_103,In_312,In_225);
xor U104 (N_104,In_496,In_319);
and U105 (N_105,In_81,In_420);
nor U106 (N_106,In_280,In_498);
or U107 (N_107,In_275,In_428);
and U108 (N_108,In_343,In_227);
or U109 (N_109,In_117,In_389);
and U110 (N_110,In_464,In_159);
and U111 (N_111,In_320,In_264);
xor U112 (N_112,In_279,In_241);
and U113 (N_113,In_54,In_11);
nand U114 (N_114,In_146,In_336);
nor U115 (N_115,In_37,In_399);
and U116 (N_116,In_165,In_170);
or U117 (N_117,In_340,In_93);
nand U118 (N_118,In_118,In_19);
nand U119 (N_119,In_281,In_491);
and U120 (N_120,In_358,In_89);
and U121 (N_121,In_132,In_499);
xor U122 (N_122,In_58,In_376);
and U123 (N_123,In_1,In_150);
nand U124 (N_124,In_297,In_414);
nor U125 (N_125,In_238,In_468);
and U126 (N_126,In_63,In_99);
nand U127 (N_127,In_350,In_322);
xor U128 (N_128,In_392,In_214);
nor U129 (N_129,In_13,In_137);
or U130 (N_130,In_375,In_476);
nor U131 (N_131,In_145,In_39);
nor U132 (N_132,In_74,In_66);
nand U133 (N_133,In_8,In_182);
nor U134 (N_134,In_380,In_396);
nor U135 (N_135,In_96,In_94);
nand U136 (N_136,In_201,In_314);
and U137 (N_137,In_456,In_230);
nand U138 (N_138,In_490,In_261);
nand U139 (N_139,In_455,In_28);
nand U140 (N_140,In_287,In_283);
xor U141 (N_141,In_106,In_493);
and U142 (N_142,In_87,In_382);
and U143 (N_143,In_135,In_92);
or U144 (N_144,In_277,In_5);
or U145 (N_145,In_197,In_136);
nor U146 (N_146,In_131,In_218);
nand U147 (N_147,In_370,In_295);
and U148 (N_148,In_180,In_308);
nor U149 (N_149,In_84,In_439);
nor U150 (N_150,In_252,In_291);
nand U151 (N_151,In_43,In_56);
or U152 (N_152,In_304,In_329);
nand U153 (N_153,In_385,In_463);
xnor U154 (N_154,In_364,In_95);
or U155 (N_155,In_473,In_60);
nand U156 (N_156,In_57,In_144);
nor U157 (N_157,In_194,In_347);
nor U158 (N_158,In_466,In_465);
xor U159 (N_159,In_492,In_77);
xor U160 (N_160,In_166,In_359);
xor U161 (N_161,In_217,In_475);
nor U162 (N_162,In_462,In_127);
nor U163 (N_163,In_55,In_33);
xor U164 (N_164,In_282,In_25);
nor U165 (N_165,In_390,In_228);
nand U166 (N_166,In_169,In_40);
or U167 (N_167,In_42,In_244);
nor U168 (N_168,In_351,In_313);
nand U169 (N_169,In_192,In_178);
xnor U170 (N_170,In_226,In_481);
or U171 (N_171,In_85,In_406);
nor U172 (N_172,In_206,In_474);
or U173 (N_173,In_436,In_23);
and U174 (N_174,In_265,In_76);
and U175 (N_175,In_108,In_378);
xnor U176 (N_176,In_337,In_223);
nor U177 (N_177,In_330,In_31);
or U178 (N_178,In_494,In_422);
xor U179 (N_179,In_105,In_305);
nor U180 (N_180,In_186,In_274);
or U181 (N_181,In_432,In_200);
or U182 (N_182,In_215,In_352);
nand U183 (N_183,In_273,In_232);
nand U184 (N_184,In_451,In_79);
nor U185 (N_185,In_459,In_111);
xnor U186 (N_186,In_243,In_158);
nand U187 (N_187,In_318,In_394);
and U188 (N_188,In_123,In_47);
or U189 (N_189,In_183,In_59);
xor U190 (N_190,In_286,In_17);
and U191 (N_191,In_152,In_401);
or U192 (N_192,In_437,In_301);
xnor U193 (N_193,In_98,In_224);
and U194 (N_194,In_188,In_373);
nand U195 (N_195,In_154,In_310);
nand U196 (N_196,In_469,In_112);
or U197 (N_197,In_363,In_450);
nand U198 (N_198,In_213,In_357);
nor U199 (N_199,In_115,In_497);
xnor U200 (N_200,In_16,In_328);
and U201 (N_201,In_156,In_397);
nor U202 (N_202,In_61,In_231);
nand U203 (N_203,In_441,In_344);
or U204 (N_204,In_269,In_472);
nor U205 (N_205,In_153,In_86);
and U206 (N_206,In_221,In_485);
and U207 (N_207,In_239,In_220);
nor U208 (N_208,In_24,In_338);
nor U209 (N_209,In_471,In_65);
nand U210 (N_210,In_303,In_361);
and U211 (N_211,In_205,In_426);
nor U212 (N_212,In_229,In_242);
nor U213 (N_213,In_411,In_149);
or U214 (N_214,In_48,In_163);
xor U215 (N_215,In_267,In_185);
xnor U216 (N_216,In_151,In_433);
nor U217 (N_217,In_125,In_452);
nand U218 (N_218,In_349,In_307);
xor U219 (N_219,In_236,In_119);
or U220 (N_220,In_421,In_161);
nor U221 (N_221,In_288,In_404);
nor U222 (N_222,In_52,In_447);
and U223 (N_223,In_296,In_237);
or U224 (N_224,In_233,In_325);
nor U225 (N_225,In_246,In_453);
nor U226 (N_226,In_260,In_271);
and U227 (N_227,In_256,In_438);
xnor U228 (N_228,In_419,In_38);
nand U229 (N_229,In_407,In_461);
xor U230 (N_230,In_470,In_333);
nor U231 (N_231,In_409,In_368);
and U232 (N_232,In_30,In_101);
nand U233 (N_233,In_102,In_482);
nand U234 (N_234,In_487,In_417);
nor U235 (N_235,In_68,In_32);
and U236 (N_236,In_203,In_64);
nand U237 (N_237,In_113,In_138);
or U238 (N_238,In_234,In_408);
nand U239 (N_239,In_29,In_208);
and U240 (N_240,In_133,In_157);
nand U241 (N_241,In_306,In_354);
nor U242 (N_242,In_335,In_130);
or U243 (N_243,In_51,In_88);
and U244 (N_244,In_6,In_440);
nor U245 (N_245,In_148,In_184);
nand U246 (N_246,In_142,In_72);
and U247 (N_247,In_332,In_278);
nand U248 (N_248,In_247,In_160);
or U249 (N_249,In_387,In_348);
nor U250 (N_250,In_233,In_84);
nand U251 (N_251,In_37,In_126);
and U252 (N_252,In_14,In_298);
and U253 (N_253,In_17,In_198);
nand U254 (N_254,In_327,In_142);
and U255 (N_255,In_234,In_3);
and U256 (N_256,In_415,In_358);
and U257 (N_257,In_126,In_385);
or U258 (N_258,In_327,In_394);
and U259 (N_259,In_148,In_211);
and U260 (N_260,In_5,In_359);
nand U261 (N_261,In_54,In_362);
and U262 (N_262,In_26,In_373);
nor U263 (N_263,In_28,In_40);
and U264 (N_264,In_14,In_438);
nand U265 (N_265,In_256,In_272);
nand U266 (N_266,In_492,In_398);
nor U267 (N_267,In_218,In_300);
nor U268 (N_268,In_415,In_475);
or U269 (N_269,In_23,In_211);
nand U270 (N_270,In_346,In_395);
nor U271 (N_271,In_219,In_234);
or U272 (N_272,In_321,In_185);
and U273 (N_273,In_160,In_159);
nor U274 (N_274,In_361,In_448);
xor U275 (N_275,In_162,In_442);
nand U276 (N_276,In_348,In_98);
nor U277 (N_277,In_481,In_229);
nand U278 (N_278,In_387,In_475);
nor U279 (N_279,In_448,In_42);
nand U280 (N_280,In_490,In_430);
or U281 (N_281,In_409,In_267);
and U282 (N_282,In_51,In_250);
or U283 (N_283,In_237,In_408);
nand U284 (N_284,In_53,In_403);
and U285 (N_285,In_390,In_284);
xor U286 (N_286,In_284,In_396);
nor U287 (N_287,In_39,In_437);
and U288 (N_288,In_3,In_39);
and U289 (N_289,In_431,In_468);
xor U290 (N_290,In_201,In_380);
nand U291 (N_291,In_5,In_252);
nor U292 (N_292,In_118,In_232);
and U293 (N_293,In_290,In_281);
or U294 (N_294,In_265,In_472);
or U295 (N_295,In_99,In_444);
and U296 (N_296,In_324,In_180);
nor U297 (N_297,In_188,In_289);
nand U298 (N_298,In_153,In_128);
nor U299 (N_299,In_16,In_187);
and U300 (N_300,In_203,In_460);
nand U301 (N_301,In_307,In_431);
or U302 (N_302,In_44,In_319);
and U303 (N_303,In_319,In_140);
nor U304 (N_304,In_266,In_180);
or U305 (N_305,In_121,In_60);
and U306 (N_306,In_106,In_479);
or U307 (N_307,In_450,In_81);
and U308 (N_308,In_321,In_100);
nor U309 (N_309,In_114,In_71);
or U310 (N_310,In_307,In_176);
nand U311 (N_311,In_333,In_358);
and U312 (N_312,In_276,In_167);
nor U313 (N_313,In_139,In_205);
and U314 (N_314,In_442,In_375);
or U315 (N_315,In_296,In_193);
nor U316 (N_316,In_412,In_83);
and U317 (N_317,In_138,In_216);
or U318 (N_318,In_451,In_327);
and U319 (N_319,In_269,In_325);
nor U320 (N_320,In_361,In_487);
nand U321 (N_321,In_146,In_319);
and U322 (N_322,In_77,In_145);
nor U323 (N_323,In_40,In_161);
nand U324 (N_324,In_347,In_340);
and U325 (N_325,In_473,In_115);
nand U326 (N_326,In_320,In_411);
and U327 (N_327,In_385,In_245);
and U328 (N_328,In_31,In_297);
and U329 (N_329,In_68,In_389);
and U330 (N_330,In_477,In_45);
nor U331 (N_331,In_260,In_84);
and U332 (N_332,In_63,In_117);
and U333 (N_333,In_251,In_241);
or U334 (N_334,In_66,In_63);
nand U335 (N_335,In_430,In_486);
and U336 (N_336,In_36,In_207);
nor U337 (N_337,In_397,In_349);
nor U338 (N_338,In_60,In_96);
or U339 (N_339,In_449,In_127);
or U340 (N_340,In_132,In_294);
or U341 (N_341,In_186,In_439);
nand U342 (N_342,In_123,In_417);
nand U343 (N_343,In_198,In_342);
and U344 (N_344,In_153,In_415);
or U345 (N_345,In_368,In_192);
nand U346 (N_346,In_278,In_161);
nand U347 (N_347,In_193,In_152);
nor U348 (N_348,In_385,In_272);
xnor U349 (N_349,In_12,In_278);
and U350 (N_350,In_79,In_391);
nand U351 (N_351,In_266,In_33);
and U352 (N_352,In_197,In_89);
or U353 (N_353,In_244,In_335);
and U354 (N_354,In_388,In_277);
nand U355 (N_355,In_128,In_249);
nor U356 (N_356,In_423,In_489);
and U357 (N_357,In_458,In_210);
xnor U358 (N_358,In_124,In_255);
nor U359 (N_359,In_318,In_438);
or U360 (N_360,In_266,In_162);
nor U361 (N_361,In_23,In_477);
nor U362 (N_362,In_174,In_4);
xnor U363 (N_363,In_318,In_6);
nor U364 (N_364,In_37,In_341);
and U365 (N_365,In_47,In_361);
or U366 (N_366,In_120,In_83);
nor U367 (N_367,In_431,In_15);
nand U368 (N_368,In_57,In_110);
and U369 (N_369,In_30,In_0);
or U370 (N_370,In_263,In_169);
or U371 (N_371,In_215,In_212);
or U372 (N_372,In_133,In_307);
or U373 (N_373,In_79,In_436);
and U374 (N_374,In_470,In_75);
nor U375 (N_375,In_190,In_81);
nand U376 (N_376,In_19,In_261);
and U377 (N_377,In_382,In_200);
and U378 (N_378,In_290,In_177);
or U379 (N_379,In_193,In_311);
nor U380 (N_380,In_147,In_349);
nor U381 (N_381,In_122,In_337);
nand U382 (N_382,In_314,In_419);
and U383 (N_383,In_206,In_413);
or U384 (N_384,In_227,In_410);
nor U385 (N_385,In_93,In_322);
nor U386 (N_386,In_343,In_204);
nand U387 (N_387,In_4,In_49);
nand U388 (N_388,In_18,In_222);
nor U389 (N_389,In_391,In_352);
xnor U390 (N_390,In_356,In_56);
xor U391 (N_391,In_184,In_137);
nor U392 (N_392,In_203,In_72);
nor U393 (N_393,In_203,In_449);
or U394 (N_394,In_494,In_290);
or U395 (N_395,In_184,In_178);
nor U396 (N_396,In_368,In_335);
nor U397 (N_397,In_37,In_225);
or U398 (N_398,In_477,In_119);
and U399 (N_399,In_22,In_267);
nor U400 (N_400,In_283,In_143);
and U401 (N_401,In_288,In_85);
and U402 (N_402,In_301,In_167);
nand U403 (N_403,In_65,In_152);
nor U404 (N_404,In_410,In_430);
or U405 (N_405,In_108,In_73);
nor U406 (N_406,In_315,In_419);
xor U407 (N_407,In_288,In_42);
nor U408 (N_408,In_182,In_232);
nand U409 (N_409,In_143,In_386);
nor U410 (N_410,In_211,In_163);
nand U411 (N_411,In_33,In_202);
or U412 (N_412,In_316,In_407);
or U413 (N_413,In_448,In_14);
nand U414 (N_414,In_212,In_177);
or U415 (N_415,In_467,In_58);
nand U416 (N_416,In_422,In_490);
nor U417 (N_417,In_382,In_287);
nand U418 (N_418,In_488,In_447);
and U419 (N_419,In_28,In_422);
or U420 (N_420,In_445,In_256);
nor U421 (N_421,In_213,In_151);
nor U422 (N_422,In_38,In_316);
and U423 (N_423,In_467,In_328);
nand U424 (N_424,In_34,In_200);
nor U425 (N_425,In_145,In_487);
nand U426 (N_426,In_265,In_133);
nor U427 (N_427,In_274,In_209);
xor U428 (N_428,In_467,In_211);
and U429 (N_429,In_44,In_111);
nor U430 (N_430,In_405,In_97);
nand U431 (N_431,In_197,In_427);
and U432 (N_432,In_336,In_172);
nor U433 (N_433,In_169,In_326);
nor U434 (N_434,In_386,In_355);
xor U435 (N_435,In_323,In_479);
nand U436 (N_436,In_283,In_359);
nor U437 (N_437,In_404,In_446);
and U438 (N_438,In_474,In_194);
nor U439 (N_439,In_83,In_6);
nor U440 (N_440,In_15,In_132);
xnor U441 (N_441,In_342,In_385);
nor U442 (N_442,In_205,In_147);
nand U443 (N_443,In_201,In_317);
xor U444 (N_444,In_60,In_351);
and U445 (N_445,In_94,In_174);
nand U446 (N_446,In_187,In_45);
nor U447 (N_447,In_475,In_141);
and U448 (N_448,In_19,In_102);
xor U449 (N_449,In_31,In_110);
nand U450 (N_450,In_51,In_265);
xnor U451 (N_451,In_218,In_159);
and U452 (N_452,In_107,In_81);
nor U453 (N_453,In_391,In_413);
nor U454 (N_454,In_472,In_145);
nand U455 (N_455,In_192,In_54);
nor U456 (N_456,In_227,In_442);
nor U457 (N_457,In_68,In_292);
nor U458 (N_458,In_109,In_104);
xnor U459 (N_459,In_452,In_451);
xnor U460 (N_460,In_298,In_467);
xor U461 (N_461,In_420,In_170);
and U462 (N_462,In_169,In_457);
and U463 (N_463,In_327,In_273);
nor U464 (N_464,In_110,In_392);
nand U465 (N_465,In_64,In_117);
nor U466 (N_466,In_393,In_379);
nor U467 (N_467,In_365,In_397);
and U468 (N_468,In_317,In_173);
nand U469 (N_469,In_165,In_180);
or U470 (N_470,In_377,In_330);
xnor U471 (N_471,In_401,In_55);
nor U472 (N_472,In_112,In_10);
or U473 (N_473,In_67,In_77);
and U474 (N_474,In_433,In_383);
nand U475 (N_475,In_496,In_397);
and U476 (N_476,In_269,In_331);
and U477 (N_477,In_40,In_348);
nor U478 (N_478,In_197,In_291);
or U479 (N_479,In_385,In_352);
or U480 (N_480,In_352,In_443);
and U481 (N_481,In_213,In_219);
nor U482 (N_482,In_394,In_317);
and U483 (N_483,In_298,In_242);
or U484 (N_484,In_146,In_304);
nand U485 (N_485,In_145,In_277);
nor U486 (N_486,In_2,In_304);
or U487 (N_487,In_52,In_446);
nand U488 (N_488,In_7,In_391);
xor U489 (N_489,In_319,In_313);
nor U490 (N_490,In_21,In_299);
or U491 (N_491,In_447,In_268);
nand U492 (N_492,In_164,In_110);
and U493 (N_493,In_374,In_478);
nor U494 (N_494,In_197,In_180);
nand U495 (N_495,In_250,In_237);
nor U496 (N_496,In_476,In_193);
nor U497 (N_497,In_448,In_366);
xnor U498 (N_498,In_324,In_313);
nor U499 (N_499,In_326,In_372);
nor U500 (N_500,In_70,In_77);
and U501 (N_501,In_247,In_11);
nor U502 (N_502,In_100,In_0);
nor U503 (N_503,In_481,In_70);
nand U504 (N_504,In_199,In_183);
nand U505 (N_505,In_235,In_217);
nor U506 (N_506,In_322,In_407);
nor U507 (N_507,In_308,In_242);
nor U508 (N_508,In_81,In_309);
or U509 (N_509,In_9,In_210);
nor U510 (N_510,In_222,In_280);
xor U511 (N_511,In_41,In_357);
nand U512 (N_512,In_467,In_249);
nand U513 (N_513,In_301,In_85);
nor U514 (N_514,In_100,In_370);
nand U515 (N_515,In_210,In_149);
or U516 (N_516,In_191,In_225);
xor U517 (N_517,In_145,In_408);
and U518 (N_518,In_374,In_114);
or U519 (N_519,In_129,In_338);
and U520 (N_520,In_33,In_8);
or U521 (N_521,In_47,In_2);
xnor U522 (N_522,In_168,In_19);
nand U523 (N_523,In_65,In_48);
nand U524 (N_524,In_253,In_27);
and U525 (N_525,In_43,In_428);
nand U526 (N_526,In_433,In_53);
nor U527 (N_527,In_162,In_249);
and U528 (N_528,In_89,In_374);
and U529 (N_529,In_311,In_7);
and U530 (N_530,In_178,In_85);
or U531 (N_531,In_330,In_368);
nor U532 (N_532,In_249,In_375);
or U533 (N_533,In_394,In_344);
nand U534 (N_534,In_330,In_39);
and U535 (N_535,In_409,In_412);
nor U536 (N_536,In_385,In_0);
nand U537 (N_537,In_212,In_257);
and U538 (N_538,In_318,In_16);
and U539 (N_539,In_398,In_63);
xnor U540 (N_540,In_382,In_288);
and U541 (N_541,In_206,In_4);
and U542 (N_542,In_425,In_0);
or U543 (N_543,In_155,In_358);
and U544 (N_544,In_377,In_368);
or U545 (N_545,In_30,In_440);
and U546 (N_546,In_395,In_135);
nor U547 (N_547,In_267,In_477);
nand U548 (N_548,In_461,In_454);
or U549 (N_549,In_351,In_192);
nand U550 (N_550,In_407,In_75);
or U551 (N_551,In_190,In_388);
and U552 (N_552,In_387,In_333);
or U553 (N_553,In_428,In_354);
xor U554 (N_554,In_392,In_191);
nand U555 (N_555,In_319,In_393);
nand U556 (N_556,In_273,In_138);
or U557 (N_557,In_12,In_335);
nand U558 (N_558,In_376,In_275);
and U559 (N_559,In_90,In_350);
nor U560 (N_560,In_314,In_324);
nor U561 (N_561,In_130,In_11);
nor U562 (N_562,In_438,In_288);
nor U563 (N_563,In_372,In_79);
xnor U564 (N_564,In_161,In_44);
and U565 (N_565,In_139,In_109);
or U566 (N_566,In_320,In_126);
xor U567 (N_567,In_329,In_493);
nor U568 (N_568,In_377,In_301);
nor U569 (N_569,In_352,In_6);
nor U570 (N_570,In_129,In_3);
xor U571 (N_571,In_164,In_423);
and U572 (N_572,In_437,In_168);
or U573 (N_573,In_489,In_163);
or U574 (N_574,In_57,In_192);
and U575 (N_575,In_384,In_165);
nand U576 (N_576,In_186,In_50);
or U577 (N_577,In_262,In_212);
and U578 (N_578,In_201,In_29);
nand U579 (N_579,In_48,In_485);
nor U580 (N_580,In_421,In_93);
nand U581 (N_581,In_442,In_444);
nor U582 (N_582,In_198,In_220);
nor U583 (N_583,In_209,In_347);
nand U584 (N_584,In_172,In_268);
xor U585 (N_585,In_348,In_148);
and U586 (N_586,In_422,In_65);
nand U587 (N_587,In_478,In_378);
nor U588 (N_588,In_294,In_251);
xnor U589 (N_589,In_176,In_414);
or U590 (N_590,In_27,In_359);
nor U591 (N_591,In_374,In_69);
nor U592 (N_592,In_419,In_468);
xnor U593 (N_593,In_33,In_315);
nor U594 (N_594,In_43,In_264);
nand U595 (N_595,In_282,In_261);
nand U596 (N_596,In_428,In_333);
nor U597 (N_597,In_292,In_161);
nand U598 (N_598,In_330,In_424);
and U599 (N_599,In_16,In_236);
or U600 (N_600,N_270,N_182);
or U601 (N_601,N_387,N_346);
nor U602 (N_602,N_52,N_121);
and U603 (N_603,N_226,N_595);
or U604 (N_604,N_18,N_166);
or U605 (N_605,N_526,N_296);
nand U606 (N_606,N_297,N_581);
and U607 (N_607,N_88,N_122);
and U608 (N_608,N_223,N_328);
or U609 (N_609,N_415,N_219);
nor U610 (N_610,N_522,N_485);
nor U611 (N_611,N_108,N_50);
and U612 (N_612,N_364,N_592);
nor U613 (N_613,N_220,N_32);
xnor U614 (N_614,N_36,N_584);
nand U615 (N_615,N_375,N_285);
and U616 (N_616,N_318,N_56);
or U617 (N_617,N_254,N_347);
and U618 (N_618,N_411,N_282);
or U619 (N_619,N_523,N_110);
or U620 (N_620,N_235,N_437);
and U621 (N_621,N_569,N_567);
xor U622 (N_622,N_113,N_206);
xor U623 (N_623,N_257,N_350);
nor U624 (N_624,N_243,N_76);
nand U625 (N_625,N_172,N_461);
xnor U626 (N_626,N_449,N_87);
xor U627 (N_627,N_16,N_348);
and U628 (N_628,N_86,N_214);
or U629 (N_629,N_309,N_42);
nor U630 (N_630,N_126,N_490);
or U631 (N_631,N_136,N_140);
or U632 (N_632,N_343,N_527);
or U633 (N_633,N_428,N_365);
or U634 (N_634,N_273,N_450);
and U635 (N_635,N_574,N_420);
and U636 (N_636,N_455,N_436);
or U637 (N_637,N_176,N_425);
nor U638 (N_638,N_286,N_211);
nand U639 (N_639,N_9,N_483);
or U640 (N_640,N_535,N_475);
nor U641 (N_641,N_540,N_85);
nor U642 (N_642,N_506,N_217);
or U643 (N_643,N_300,N_359);
nand U644 (N_644,N_61,N_43);
and U645 (N_645,N_105,N_575);
nor U646 (N_646,N_491,N_432);
and U647 (N_647,N_128,N_355);
or U648 (N_648,N_508,N_67);
xnor U649 (N_649,N_204,N_497);
or U650 (N_650,N_591,N_13);
nand U651 (N_651,N_403,N_64);
or U652 (N_652,N_54,N_45);
nand U653 (N_653,N_144,N_384);
nor U654 (N_654,N_555,N_493);
and U655 (N_655,N_440,N_307);
or U656 (N_656,N_345,N_230);
nand U657 (N_657,N_580,N_317);
and U658 (N_658,N_380,N_287);
xor U659 (N_659,N_196,N_304);
or U660 (N_660,N_542,N_53);
xnor U661 (N_661,N_504,N_404);
and U662 (N_662,N_103,N_325);
nand U663 (N_663,N_114,N_92);
nor U664 (N_664,N_118,N_258);
nor U665 (N_665,N_549,N_78);
xor U666 (N_666,N_167,N_84);
or U667 (N_667,N_502,N_530);
and U668 (N_668,N_181,N_568);
nand U669 (N_669,N_561,N_119);
xnor U670 (N_670,N_252,N_495);
nand U671 (N_671,N_259,N_330);
nor U672 (N_672,N_338,N_533);
and U673 (N_673,N_227,N_202);
and U674 (N_674,N_138,N_12);
or U675 (N_675,N_298,N_102);
and U676 (N_676,N_131,N_283);
or U677 (N_677,N_543,N_168);
nor U678 (N_678,N_71,N_448);
xor U679 (N_679,N_412,N_583);
or U680 (N_680,N_556,N_409);
or U681 (N_681,N_547,N_154);
nand U682 (N_682,N_165,N_472);
and U683 (N_683,N_344,N_210);
or U684 (N_684,N_231,N_130);
and U685 (N_685,N_517,N_190);
or U686 (N_686,N_189,N_185);
nand U687 (N_687,N_510,N_70);
nand U688 (N_688,N_200,N_498);
nor U689 (N_689,N_319,N_478);
xnor U690 (N_690,N_303,N_145);
and U691 (N_691,N_80,N_596);
nor U692 (N_692,N_435,N_418);
nor U693 (N_693,N_22,N_25);
and U694 (N_694,N_201,N_10);
nor U695 (N_695,N_51,N_101);
nand U696 (N_696,N_323,N_492);
and U697 (N_697,N_470,N_577);
and U698 (N_698,N_321,N_315);
and U699 (N_699,N_163,N_6);
and U700 (N_700,N_38,N_207);
nand U701 (N_701,N_479,N_46);
nand U702 (N_702,N_310,N_228);
xor U703 (N_703,N_594,N_55);
nor U704 (N_704,N_139,N_597);
xnor U705 (N_705,N_7,N_520);
and U706 (N_706,N_388,N_566);
or U707 (N_707,N_209,N_271);
xor U708 (N_708,N_75,N_39);
and U709 (N_709,N_353,N_93);
nor U710 (N_710,N_289,N_153);
nand U711 (N_711,N_586,N_494);
xor U712 (N_712,N_35,N_374);
or U713 (N_713,N_593,N_143);
nand U714 (N_714,N_77,N_473);
or U715 (N_715,N_134,N_312);
and U716 (N_716,N_534,N_573);
xor U717 (N_717,N_147,N_135);
or U718 (N_718,N_554,N_314);
nor U719 (N_719,N_326,N_571);
nand U720 (N_720,N_394,N_419);
or U721 (N_721,N_268,N_550);
nor U722 (N_722,N_170,N_358);
nand U723 (N_723,N_553,N_74);
or U724 (N_724,N_557,N_213);
nand U725 (N_725,N_302,N_8);
nand U726 (N_726,N_249,N_447);
nand U727 (N_727,N_261,N_565);
nor U728 (N_728,N_162,N_322);
or U729 (N_729,N_247,N_188);
xnor U730 (N_730,N_15,N_57);
nor U731 (N_731,N_332,N_149);
or U732 (N_732,N_212,N_292);
nor U733 (N_733,N_260,N_352);
nor U734 (N_734,N_240,N_552);
nor U735 (N_735,N_205,N_469);
nand U736 (N_736,N_416,N_14);
and U737 (N_737,N_465,N_487);
or U738 (N_738,N_59,N_241);
nor U739 (N_739,N_117,N_486);
or U740 (N_740,N_429,N_41);
or U741 (N_741,N_445,N_203);
nor U742 (N_742,N_104,N_439);
and U743 (N_743,N_360,N_524);
nor U744 (N_744,N_293,N_127);
and U745 (N_745,N_578,N_393);
xnor U746 (N_746,N_367,N_512);
xnor U747 (N_747,N_266,N_458);
nand U748 (N_748,N_408,N_146);
and U749 (N_749,N_528,N_137);
nand U750 (N_750,N_539,N_161);
and U751 (N_751,N_19,N_320);
or U752 (N_752,N_109,N_208);
or U753 (N_753,N_399,N_224);
xnor U754 (N_754,N_288,N_3);
and U755 (N_755,N_99,N_541);
xnor U756 (N_756,N_65,N_180);
or U757 (N_757,N_467,N_96);
or U758 (N_758,N_284,N_372);
nor U759 (N_759,N_521,N_152);
or U760 (N_760,N_516,N_563);
nand U761 (N_761,N_545,N_171);
nand U762 (N_762,N_299,N_68);
nand U763 (N_763,N_587,N_503);
nor U764 (N_764,N_385,N_337);
nor U765 (N_765,N_335,N_383);
and U766 (N_766,N_395,N_468);
nor U767 (N_767,N_390,N_576);
and U768 (N_768,N_525,N_115);
nor U769 (N_769,N_216,N_471);
or U770 (N_770,N_301,N_81);
and U771 (N_771,N_476,N_444);
nor U772 (N_772,N_111,N_351);
and U773 (N_773,N_294,N_397);
nor U774 (N_774,N_482,N_234);
and U775 (N_775,N_150,N_278);
xnor U776 (N_776,N_178,N_169);
and U777 (N_777,N_373,N_441);
nor U778 (N_778,N_489,N_499);
nand U779 (N_779,N_187,N_463);
and U780 (N_780,N_237,N_66);
nor U781 (N_781,N_164,N_116);
nor U782 (N_782,N_221,N_267);
and U783 (N_783,N_398,N_590);
and U784 (N_784,N_244,N_157);
nand U785 (N_785,N_598,N_481);
and U786 (N_786,N_342,N_434);
nand U787 (N_787,N_277,N_329);
and U788 (N_788,N_69,N_446);
and U789 (N_789,N_97,N_290);
or U790 (N_790,N_120,N_269);
xnor U791 (N_791,N_48,N_107);
nand U792 (N_792,N_464,N_431);
nand U793 (N_793,N_148,N_391);
or U794 (N_794,N_60,N_133);
nor U795 (N_795,N_215,N_132);
nand U796 (N_796,N_23,N_378);
and U797 (N_797,N_197,N_73);
and U798 (N_798,N_379,N_381);
nand U799 (N_799,N_406,N_225);
and U800 (N_800,N_401,N_537);
nand U801 (N_801,N_564,N_459);
or U802 (N_802,N_79,N_232);
nand U803 (N_803,N_155,N_536);
and U804 (N_804,N_513,N_529);
nand U805 (N_805,N_392,N_366);
or U806 (N_806,N_179,N_194);
xnor U807 (N_807,N_173,N_106);
nor U808 (N_808,N_100,N_239);
and U809 (N_809,N_251,N_123);
or U810 (N_810,N_21,N_313);
nand U811 (N_811,N_183,N_558);
and U812 (N_812,N_514,N_82);
and U813 (N_813,N_443,N_363);
and U814 (N_814,N_47,N_361);
nor U815 (N_815,N_0,N_334);
or U816 (N_816,N_280,N_191);
nor U817 (N_817,N_245,N_177);
nand U818 (N_818,N_20,N_386);
nor U819 (N_819,N_570,N_442);
nand U820 (N_820,N_272,N_40);
nand U821 (N_821,N_400,N_238);
and U822 (N_822,N_34,N_263);
nor U823 (N_823,N_256,N_305);
or U824 (N_824,N_11,N_474);
xor U825 (N_825,N_233,N_496);
nand U826 (N_826,N_63,N_341);
or U827 (N_827,N_327,N_422);
or U828 (N_828,N_264,N_27);
nand U829 (N_829,N_585,N_572);
nand U830 (N_830,N_370,N_453);
nor U831 (N_831,N_414,N_349);
and U832 (N_832,N_324,N_37);
nor U833 (N_833,N_262,N_62);
and U834 (N_834,N_253,N_2);
or U835 (N_835,N_396,N_454);
or U836 (N_836,N_462,N_427);
or U837 (N_837,N_89,N_31);
nand U838 (N_838,N_369,N_426);
or U839 (N_839,N_466,N_274);
or U840 (N_840,N_579,N_507);
nor U841 (N_841,N_582,N_589);
nor U842 (N_842,N_281,N_222);
nand U843 (N_843,N_246,N_389);
nand U844 (N_844,N_265,N_94);
nand U845 (N_845,N_308,N_410);
nand U846 (N_846,N_546,N_402);
and U847 (N_847,N_509,N_186);
nand U848 (N_848,N_28,N_518);
or U849 (N_849,N_279,N_548);
and U850 (N_850,N_44,N_58);
nor U851 (N_851,N_480,N_377);
and U852 (N_852,N_457,N_538);
and U853 (N_853,N_24,N_112);
or U854 (N_854,N_515,N_248);
nor U855 (N_855,N_433,N_339);
and U856 (N_856,N_421,N_588);
or U857 (N_857,N_438,N_505);
or U858 (N_858,N_255,N_1);
xnor U859 (N_859,N_26,N_423);
and U860 (N_860,N_417,N_405);
xor U861 (N_861,N_159,N_291);
nand U862 (N_862,N_174,N_141);
and U863 (N_863,N_532,N_275);
nand U864 (N_864,N_488,N_371);
or U865 (N_865,N_562,N_17);
and U866 (N_866,N_151,N_460);
nor U867 (N_867,N_184,N_356);
nor U868 (N_868,N_336,N_306);
nor U869 (N_869,N_551,N_362);
nor U870 (N_870,N_218,N_451);
nand U871 (N_871,N_229,N_236);
xor U872 (N_872,N_158,N_368);
and U873 (N_873,N_599,N_95);
and U874 (N_874,N_83,N_90);
nor U875 (N_875,N_125,N_129);
or U876 (N_876,N_160,N_519);
nand U877 (N_877,N_316,N_452);
or U878 (N_878,N_193,N_276);
or U879 (N_879,N_413,N_5);
and U880 (N_880,N_30,N_376);
xor U881 (N_881,N_242,N_199);
and U882 (N_882,N_198,N_124);
nand U883 (N_883,N_195,N_511);
and U884 (N_884,N_142,N_250);
nand U885 (N_885,N_72,N_382);
and U886 (N_886,N_333,N_29);
xor U887 (N_887,N_331,N_484);
nand U888 (N_888,N_311,N_430);
nand U889 (N_889,N_49,N_424);
or U890 (N_890,N_544,N_98);
nor U891 (N_891,N_500,N_407);
nor U892 (N_892,N_560,N_91);
and U893 (N_893,N_354,N_175);
or U894 (N_894,N_33,N_477);
and U895 (N_895,N_456,N_156);
xor U896 (N_896,N_531,N_501);
or U897 (N_897,N_340,N_357);
and U898 (N_898,N_295,N_192);
nand U899 (N_899,N_559,N_4);
and U900 (N_900,N_358,N_396);
nor U901 (N_901,N_556,N_15);
nor U902 (N_902,N_482,N_104);
nand U903 (N_903,N_582,N_147);
nor U904 (N_904,N_212,N_534);
nor U905 (N_905,N_414,N_282);
or U906 (N_906,N_289,N_57);
or U907 (N_907,N_129,N_58);
or U908 (N_908,N_143,N_246);
or U909 (N_909,N_39,N_77);
or U910 (N_910,N_24,N_271);
and U911 (N_911,N_330,N_409);
or U912 (N_912,N_590,N_418);
or U913 (N_913,N_270,N_199);
and U914 (N_914,N_556,N_542);
nor U915 (N_915,N_565,N_276);
xnor U916 (N_916,N_208,N_402);
nand U917 (N_917,N_403,N_485);
nor U918 (N_918,N_158,N_192);
or U919 (N_919,N_10,N_394);
and U920 (N_920,N_170,N_256);
xor U921 (N_921,N_66,N_478);
nand U922 (N_922,N_354,N_99);
nor U923 (N_923,N_591,N_549);
and U924 (N_924,N_117,N_387);
nand U925 (N_925,N_109,N_73);
xor U926 (N_926,N_271,N_503);
and U927 (N_927,N_50,N_153);
or U928 (N_928,N_410,N_205);
nor U929 (N_929,N_1,N_361);
and U930 (N_930,N_78,N_199);
or U931 (N_931,N_233,N_38);
or U932 (N_932,N_286,N_359);
nand U933 (N_933,N_458,N_211);
nand U934 (N_934,N_216,N_240);
nor U935 (N_935,N_13,N_588);
nor U936 (N_936,N_113,N_55);
nor U937 (N_937,N_445,N_256);
nand U938 (N_938,N_471,N_537);
and U939 (N_939,N_135,N_63);
nor U940 (N_940,N_342,N_520);
or U941 (N_941,N_304,N_419);
nor U942 (N_942,N_269,N_211);
nand U943 (N_943,N_161,N_529);
nand U944 (N_944,N_31,N_549);
or U945 (N_945,N_564,N_107);
nand U946 (N_946,N_382,N_5);
nand U947 (N_947,N_33,N_442);
and U948 (N_948,N_79,N_479);
nor U949 (N_949,N_445,N_310);
xor U950 (N_950,N_438,N_160);
and U951 (N_951,N_412,N_149);
or U952 (N_952,N_418,N_72);
xor U953 (N_953,N_278,N_231);
and U954 (N_954,N_591,N_583);
or U955 (N_955,N_518,N_296);
nand U956 (N_956,N_557,N_499);
xnor U957 (N_957,N_341,N_292);
xor U958 (N_958,N_567,N_259);
nand U959 (N_959,N_18,N_66);
nand U960 (N_960,N_88,N_426);
and U961 (N_961,N_38,N_409);
xnor U962 (N_962,N_302,N_63);
nand U963 (N_963,N_381,N_320);
nor U964 (N_964,N_339,N_553);
or U965 (N_965,N_199,N_107);
nor U966 (N_966,N_570,N_435);
xnor U967 (N_967,N_547,N_576);
and U968 (N_968,N_557,N_359);
or U969 (N_969,N_168,N_503);
and U970 (N_970,N_365,N_203);
nand U971 (N_971,N_578,N_42);
nand U972 (N_972,N_262,N_160);
nor U973 (N_973,N_257,N_560);
nor U974 (N_974,N_159,N_449);
nand U975 (N_975,N_37,N_467);
nand U976 (N_976,N_563,N_9);
xnor U977 (N_977,N_214,N_242);
or U978 (N_978,N_384,N_1);
or U979 (N_979,N_131,N_369);
or U980 (N_980,N_504,N_39);
and U981 (N_981,N_148,N_399);
or U982 (N_982,N_151,N_402);
nand U983 (N_983,N_196,N_330);
and U984 (N_984,N_555,N_100);
or U985 (N_985,N_36,N_247);
or U986 (N_986,N_504,N_390);
and U987 (N_987,N_438,N_332);
and U988 (N_988,N_38,N_179);
and U989 (N_989,N_255,N_51);
or U990 (N_990,N_456,N_28);
nor U991 (N_991,N_132,N_288);
and U992 (N_992,N_68,N_354);
xor U993 (N_993,N_82,N_384);
and U994 (N_994,N_75,N_167);
nand U995 (N_995,N_345,N_431);
nor U996 (N_996,N_216,N_496);
or U997 (N_997,N_154,N_163);
nor U998 (N_998,N_509,N_169);
nor U999 (N_999,N_243,N_355);
and U1000 (N_1000,N_333,N_148);
nor U1001 (N_1001,N_332,N_132);
or U1002 (N_1002,N_91,N_102);
xnor U1003 (N_1003,N_596,N_271);
nor U1004 (N_1004,N_149,N_506);
and U1005 (N_1005,N_344,N_258);
or U1006 (N_1006,N_539,N_48);
or U1007 (N_1007,N_596,N_390);
nor U1008 (N_1008,N_525,N_246);
nand U1009 (N_1009,N_227,N_34);
or U1010 (N_1010,N_14,N_57);
and U1011 (N_1011,N_354,N_385);
xnor U1012 (N_1012,N_484,N_135);
nor U1013 (N_1013,N_526,N_450);
and U1014 (N_1014,N_278,N_539);
nor U1015 (N_1015,N_499,N_494);
xor U1016 (N_1016,N_69,N_170);
nor U1017 (N_1017,N_530,N_226);
nor U1018 (N_1018,N_598,N_502);
or U1019 (N_1019,N_357,N_502);
nor U1020 (N_1020,N_58,N_229);
or U1021 (N_1021,N_266,N_448);
or U1022 (N_1022,N_363,N_126);
nand U1023 (N_1023,N_5,N_217);
nor U1024 (N_1024,N_491,N_481);
and U1025 (N_1025,N_98,N_213);
or U1026 (N_1026,N_311,N_307);
xor U1027 (N_1027,N_393,N_91);
or U1028 (N_1028,N_279,N_571);
nor U1029 (N_1029,N_50,N_141);
nor U1030 (N_1030,N_557,N_147);
or U1031 (N_1031,N_185,N_598);
nand U1032 (N_1032,N_87,N_510);
or U1033 (N_1033,N_103,N_524);
nand U1034 (N_1034,N_352,N_358);
nand U1035 (N_1035,N_441,N_239);
and U1036 (N_1036,N_586,N_248);
nand U1037 (N_1037,N_413,N_255);
and U1038 (N_1038,N_225,N_453);
or U1039 (N_1039,N_90,N_220);
or U1040 (N_1040,N_568,N_318);
nand U1041 (N_1041,N_275,N_254);
and U1042 (N_1042,N_518,N_178);
nand U1043 (N_1043,N_344,N_524);
nand U1044 (N_1044,N_496,N_14);
nand U1045 (N_1045,N_472,N_18);
nor U1046 (N_1046,N_459,N_316);
nand U1047 (N_1047,N_141,N_495);
xnor U1048 (N_1048,N_352,N_528);
xor U1049 (N_1049,N_293,N_510);
xor U1050 (N_1050,N_157,N_265);
nor U1051 (N_1051,N_311,N_472);
or U1052 (N_1052,N_156,N_543);
nand U1053 (N_1053,N_168,N_458);
or U1054 (N_1054,N_316,N_327);
or U1055 (N_1055,N_96,N_219);
nor U1056 (N_1056,N_476,N_84);
nand U1057 (N_1057,N_333,N_313);
nor U1058 (N_1058,N_337,N_11);
nor U1059 (N_1059,N_153,N_328);
nand U1060 (N_1060,N_9,N_83);
nor U1061 (N_1061,N_67,N_422);
xor U1062 (N_1062,N_42,N_452);
or U1063 (N_1063,N_226,N_313);
nand U1064 (N_1064,N_507,N_416);
or U1065 (N_1065,N_442,N_384);
or U1066 (N_1066,N_46,N_439);
nor U1067 (N_1067,N_106,N_442);
xor U1068 (N_1068,N_516,N_583);
nand U1069 (N_1069,N_449,N_588);
nor U1070 (N_1070,N_380,N_228);
nor U1071 (N_1071,N_242,N_101);
and U1072 (N_1072,N_306,N_89);
and U1073 (N_1073,N_205,N_184);
and U1074 (N_1074,N_299,N_318);
or U1075 (N_1075,N_534,N_111);
or U1076 (N_1076,N_93,N_340);
or U1077 (N_1077,N_117,N_458);
and U1078 (N_1078,N_299,N_257);
nand U1079 (N_1079,N_563,N_76);
nor U1080 (N_1080,N_406,N_558);
and U1081 (N_1081,N_32,N_74);
nand U1082 (N_1082,N_302,N_401);
or U1083 (N_1083,N_470,N_60);
and U1084 (N_1084,N_325,N_497);
nor U1085 (N_1085,N_53,N_346);
and U1086 (N_1086,N_67,N_576);
or U1087 (N_1087,N_465,N_130);
xor U1088 (N_1088,N_425,N_593);
and U1089 (N_1089,N_247,N_479);
nand U1090 (N_1090,N_534,N_166);
or U1091 (N_1091,N_76,N_522);
xor U1092 (N_1092,N_374,N_12);
or U1093 (N_1093,N_550,N_182);
nand U1094 (N_1094,N_581,N_477);
nor U1095 (N_1095,N_384,N_202);
nor U1096 (N_1096,N_113,N_303);
nor U1097 (N_1097,N_290,N_525);
or U1098 (N_1098,N_165,N_230);
nor U1099 (N_1099,N_476,N_433);
and U1100 (N_1100,N_203,N_60);
and U1101 (N_1101,N_217,N_355);
xor U1102 (N_1102,N_587,N_542);
and U1103 (N_1103,N_456,N_143);
nand U1104 (N_1104,N_164,N_227);
or U1105 (N_1105,N_275,N_181);
nor U1106 (N_1106,N_348,N_208);
and U1107 (N_1107,N_69,N_485);
or U1108 (N_1108,N_92,N_324);
xnor U1109 (N_1109,N_80,N_452);
nor U1110 (N_1110,N_291,N_399);
or U1111 (N_1111,N_374,N_328);
and U1112 (N_1112,N_519,N_282);
or U1113 (N_1113,N_181,N_288);
xor U1114 (N_1114,N_582,N_59);
and U1115 (N_1115,N_24,N_117);
and U1116 (N_1116,N_335,N_217);
nor U1117 (N_1117,N_315,N_384);
and U1118 (N_1118,N_295,N_124);
or U1119 (N_1119,N_90,N_282);
nand U1120 (N_1120,N_201,N_488);
or U1121 (N_1121,N_581,N_159);
nor U1122 (N_1122,N_563,N_40);
nor U1123 (N_1123,N_558,N_154);
or U1124 (N_1124,N_547,N_533);
or U1125 (N_1125,N_371,N_483);
and U1126 (N_1126,N_480,N_444);
xnor U1127 (N_1127,N_554,N_539);
and U1128 (N_1128,N_185,N_14);
xor U1129 (N_1129,N_148,N_92);
nor U1130 (N_1130,N_375,N_57);
nand U1131 (N_1131,N_77,N_156);
nand U1132 (N_1132,N_204,N_596);
nand U1133 (N_1133,N_173,N_194);
nor U1134 (N_1134,N_30,N_309);
or U1135 (N_1135,N_598,N_179);
xnor U1136 (N_1136,N_372,N_22);
nor U1137 (N_1137,N_321,N_522);
or U1138 (N_1138,N_361,N_109);
and U1139 (N_1139,N_92,N_452);
nand U1140 (N_1140,N_484,N_247);
and U1141 (N_1141,N_136,N_59);
nor U1142 (N_1142,N_75,N_527);
and U1143 (N_1143,N_563,N_141);
and U1144 (N_1144,N_307,N_399);
and U1145 (N_1145,N_487,N_99);
nor U1146 (N_1146,N_27,N_212);
nand U1147 (N_1147,N_252,N_331);
nand U1148 (N_1148,N_314,N_49);
nor U1149 (N_1149,N_105,N_52);
nor U1150 (N_1150,N_313,N_227);
or U1151 (N_1151,N_119,N_438);
and U1152 (N_1152,N_567,N_320);
nand U1153 (N_1153,N_340,N_1);
or U1154 (N_1154,N_76,N_281);
and U1155 (N_1155,N_197,N_88);
nand U1156 (N_1156,N_105,N_396);
or U1157 (N_1157,N_595,N_193);
nand U1158 (N_1158,N_355,N_586);
nand U1159 (N_1159,N_304,N_577);
and U1160 (N_1160,N_320,N_574);
or U1161 (N_1161,N_79,N_118);
and U1162 (N_1162,N_79,N_50);
or U1163 (N_1163,N_515,N_514);
nor U1164 (N_1164,N_568,N_522);
nand U1165 (N_1165,N_409,N_58);
or U1166 (N_1166,N_442,N_193);
nand U1167 (N_1167,N_268,N_364);
nand U1168 (N_1168,N_492,N_168);
xnor U1169 (N_1169,N_548,N_294);
nor U1170 (N_1170,N_379,N_541);
nand U1171 (N_1171,N_250,N_144);
or U1172 (N_1172,N_358,N_87);
nand U1173 (N_1173,N_278,N_155);
and U1174 (N_1174,N_170,N_407);
and U1175 (N_1175,N_483,N_132);
or U1176 (N_1176,N_479,N_40);
nand U1177 (N_1177,N_346,N_229);
or U1178 (N_1178,N_463,N_170);
nand U1179 (N_1179,N_322,N_170);
nor U1180 (N_1180,N_232,N_59);
or U1181 (N_1181,N_221,N_478);
and U1182 (N_1182,N_68,N_330);
and U1183 (N_1183,N_455,N_570);
nor U1184 (N_1184,N_326,N_183);
xor U1185 (N_1185,N_227,N_104);
and U1186 (N_1186,N_439,N_463);
or U1187 (N_1187,N_204,N_80);
nand U1188 (N_1188,N_134,N_441);
nand U1189 (N_1189,N_355,N_390);
and U1190 (N_1190,N_226,N_431);
xor U1191 (N_1191,N_141,N_151);
or U1192 (N_1192,N_415,N_533);
and U1193 (N_1193,N_474,N_43);
or U1194 (N_1194,N_154,N_241);
nor U1195 (N_1195,N_523,N_81);
or U1196 (N_1196,N_324,N_0);
or U1197 (N_1197,N_457,N_85);
nand U1198 (N_1198,N_302,N_213);
and U1199 (N_1199,N_305,N_60);
or U1200 (N_1200,N_1194,N_1052);
nor U1201 (N_1201,N_1141,N_815);
nand U1202 (N_1202,N_1042,N_869);
nand U1203 (N_1203,N_765,N_690);
nand U1204 (N_1204,N_941,N_798);
and U1205 (N_1205,N_1094,N_943);
nand U1206 (N_1206,N_1104,N_861);
or U1207 (N_1207,N_1162,N_944);
nor U1208 (N_1208,N_923,N_809);
nand U1209 (N_1209,N_1036,N_703);
xor U1210 (N_1210,N_977,N_1101);
nor U1211 (N_1211,N_1181,N_752);
nor U1212 (N_1212,N_1176,N_1033);
nor U1213 (N_1213,N_931,N_785);
and U1214 (N_1214,N_937,N_699);
and U1215 (N_1215,N_805,N_773);
or U1216 (N_1216,N_762,N_1166);
nor U1217 (N_1217,N_613,N_863);
nand U1218 (N_1218,N_1048,N_1108);
nand U1219 (N_1219,N_1085,N_634);
and U1220 (N_1220,N_600,N_656);
nand U1221 (N_1221,N_767,N_741);
xnor U1222 (N_1222,N_950,N_1148);
and U1223 (N_1223,N_654,N_802);
nor U1224 (N_1224,N_640,N_832);
and U1225 (N_1225,N_947,N_826);
xnor U1226 (N_1226,N_1103,N_786);
nor U1227 (N_1227,N_845,N_751);
or U1228 (N_1228,N_632,N_687);
nand U1229 (N_1229,N_1045,N_1002);
nor U1230 (N_1230,N_669,N_747);
or U1231 (N_1231,N_966,N_898);
nor U1232 (N_1232,N_917,N_840);
nor U1233 (N_1233,N_1161,N_666);
or U1234 (N_1234,N_987,N_1113);
and U1235 (N_1235,N_776,N_738);
or U1236 (N_1236,N_736,N_1060);
nand U1237 (N_1237,N_761,N_1071);
xnor U1238 (N_1238,N_719,N_1032);
xnor U1239 (N_1239,N_828,N_1139);
nor U1240 (N_1240,N_760,N_695);
nor U1241 (N_1241,N_994,N_718);
or U1242 (N_1242,N_1000,N_1023);
or U1243 (N_1243,N_755,N_928);
or U1244 (N_1244,N_920,N_880);
nand U1245 (N_1245,N_862,N_866);
or U1246 (N_1246,N_721,N_1169);
xor U1247 (N_1247,N_1018,N_812);
xor U1248 (N_1248,N_919,N_1190);
or U1249 (N_1249,N_650,N_1009);
nand U1250 (N_1250,N_681,N_713);
and U1251 (N_1251,N_1159,N_1037);
nor U1252 (N_1252,N_636,N_745);
and U1253 (N_1253,N_924,N_670);
or U1254 (N_1254,N_817,N_1152);
and U1255 (N_1255,N_649,N_953);
nand U1256 (N_1256,N_1074,N_971);
and U1257 (N_1257,N_1046,N_1021);
nor U1258 (N_1258,N_975,N_1167);
nand U1259 (N_1259,N_1006,N_852);
nor U1260 (N_1260,N_693,N_1112);
xor U1261 (N_1261,N_878,N_968);
and U1262 (N_1262,N_609,N_897);
or U1263 (N_1263,N_874,N_691);
and U1264 (N_1264,N_668,N_888);
nand U1265 (N_1265,N_1040,N_1007);
nor U1266 (N_1266,N_715,N_934);
nor U1267 (N_1267,N_659,N_955);
nor U1268 (N_1268,N_611,N_633);
nand U1269 (N_1269,N_1043,N_729);
or U1270 (N_1270,N_638,N_932);
nor U1271 (N_1271,N_1090,N_885);
or U1272 (N_1272,N_743,N_1053);
or U1273 (N_1273,N_744,N_637);
nor U1274 (N_1274,N_856,N_855);
xor U1275 (N_1275,N_635,N_696);
or U1276 (N_1276,N_607,N_688);
nor U1277 (N_1277,N_1063,N_835);
xnor U1278 (N_1278,N_782,N_922);
nand U1279 (N_1279,N_972,N_1135);
nor U1280 (N_1280,N_877,N_1182);
nor U1281 (N_1281,N_959,N_1069);
nand U1282 (N_1282,N_653,N_896);
xor U1283 (N_1283,N_1030,N_1127);
nand U1284 (N_1284,N_842,N_882);
nor U1285 (N_1285,N_851,N_1082);
nor U1286 (N_1286,N_1058,N_889);
and U1287 (N_1287,N_999,N_1184);
nor U1288 (N_1288,N_868,N_992);
or U1289 (N_1289,N_870,N_1196);
nor U1290 (N_1290,N_720,N_887);
nor U1291 (N_1291,N_914,N_1140);
and U1292 (N_1292,N_908,N_929);
or U1293 (N_1293,N_819,N_854);
and U1294 (N_1294,N_1128,N_705);
and U1295 (N_1295,N_630,N_1143);
nand U1296 (N_1296,N_871,N_772);
or U1297 (N_1297,N_1137,N_1056);
or U1298 (N_1298,N_652,N_1034);
xor U1299 (N_1299,N_1197,N_686);
and U1300 (N_1300,N_1189,N_876);
and U1301 (N_1301,N_1163,N_1003);
xor U1302 (N_1302,N_683,N_831);
or U1303 (N_1303,N_682,N_619);
or U1304 (N_1304,N_958,N_872);
nor U1305 (N_1305,N_764,N_701);
and U1306 (N_1306,N_671,N_811);
nand U1307 (N_1307,N_757,N_1049);
nand U1308 (N_1308,N_1022,N_787);
or U1309 (N_1309,N_1026,N_796);
or U1310 (N_1310,N_1099,N_1079);
nand U1311 (N_1311,N_1100,N_753);
nand U1312 (N_1312,N_672,N_1156);
nor U1313 (N_1313,N_1177,N_935);
and U1314 (N_1314,N_961,N_865);
nand U1315 (N_1315,N_980,N_1096);
xor U1316 (N_1316,N_1076,N_900);
and U1317 (N_1317,N_1129,N_833);
or U1318 (N_1318,N_601,N_879);
nor U1319 (N_1319,N_1155,N_1198);
nand U1320 (N_1320,N_899,N_912);
and U1321 (N_1321,N_771,N_620);
nor U1322 (N_1322,N_881,N_1111);
or U1323 (N_1323,N_604,N_822);
or U1324 (N_1324,N_742,N_1067);
and U1325 (N_1325,N_1149,N_960);
and U1326 (N_1326,N_847,N_892);
nand U1327 (N_1327,N_1070,N_1133);
or U1328 (N_1328,N_841,N_1154);
nor U1329 (N_1329,N_915,N_970);
and U1330 (N_1330,N_665,N_722);
nand U1331 (N_1331,N_952,N_731);
nand U1332 (N_1332,N_1017,N_926);
and U1333 (N_1333,N_1125,N_991);
nand U1334 (N_1334,N_1012,N_702);
xor U1335 (N_1335,N_1029,N_698);
nand U1336 (N_1336,N_711,N_990);
or U1337 (N_1337,N_774,N_618);
and U1338 (N_1338,N_1024,N_939);
nor U1339 (N_1339,N_694,N_820);
nor U1340 (N_1340,N_1150,N_1057);
nand U1341 (N_1341,N_766,N_1118);
or U1342 (N_1342,N_989,N_967);
nor U1343 (N_1343,N_1164,N_1047);
or U1344 (N_1344,N_647,N_1008);
or U1345 (N_1345,N_1130,N_602);
nand U1346 (N_1346,N_1146,N_986);
and U1347 (N_1347,N_1039,N_838);
nor U1348 (N_1348,N_737,N_976);
or U1349 (N_1349,N_1110,N_685);
nor U1350 (N_1350,N_853,N_843);
nor U1351 (N_1351,N_846,N_1171);
nor U1352 (N_1352,N_645,N_735);
or U1353 (N_1353,N_995,N_1142);
xor U1354 (N_1354,N_603,N_756);
or U1355 (N_1355,N_1170,N_824);
nor U1356 (N_1356,N_697,N_1001);
xor U1357 (N_1357,N_749,N_918);
nand U1358 (N_1358,N_978,N_617);
xor U1359 (N_1359,N_951,N_710);
and U1360 (N_1360,N_606,N_740);
nor U1361 (N_1361,N_655,N_1134);
nor U1362 (N_1362,N_837,N_848);
and U1363 (N_1363,N_883,N_827);
nand U1364 (N_1364,N_792,N_732);
and U1365 (N_1365,N_621,N_657);
or U1366 (N_1366,N_1019,N_615);
xnor U1367 (N_1367,N_954,N_823);
nand U1368 (N_1368,N_708,N_763);
nor U1369 (N_1369,N_804,N_769);
nor U1370 (N_1370,N_1165,N_723);
xor U1371 (N_1371,N_906,N_921);
and U1372 (N_1372,N_631,N_974);
xor U1373 (N_1373,N_1072,N_608);
nand U1374 (N_1374,N_1124,N_689);
or U1375 (N_1375,N_795,N_1175);
nor U1376 (N_1376,N_909,N_849);
xnor U1377 (N_1377,N_628,N_662);
and U1378 (N_1378,N_1028,N_675);
and U1379 (N_1379,N_1116,N_783);
nor U1380 (N_1380,N_1095,N_1011);
nand U1381 (N_1381,N_777,N_907);
nor U1382 (N_1382,N_1087,N_1084);
nand U1383 (N_1383,N_1187,N_780);
nor U1384 (N_1384,N_902,N_816);
or U1385 (N_1385,N_680,N_988);
or U1386 (N_1386,N_1015,N_1105);
and U1387 (N_1387,N_768,N_1035);
nand U1388 (N_1388,N_624,N_981);
or U1389 (N_1389,N_1120,N_754);
or U1390 (N_1390,N_790,N_1080);
or U1391 (N_1391,N_1098,N_1050);
nor U1392 (N_1392,N_810,N_948);
nand U1393 (N_1393,N_1173,N_748);
or U1394 (N_1394,N_1126,N_873);
or U1395 (N_1395,N_884,N_1183);
or U1396 (N_1396,N_1083,N_1066);
and U1397 (N_1397,N_904,N_933);
nand U1398 (N_1398,N_1172,N_1157);
or U1399 (N_1399,N_679,N_836);
nand U1400 (N_1400,N_1147,N_979);
nand U1401 (N_1401,N_734,N_1121);
and U1402 (N_1402,N_676,N_1062);
or U1403 (N_1403,N_1119,N_724);
xnor U1404 (N_1404,N_684,N_1174);
nor U1405 (N_1405,N_886,N_1123);
nand U1406 (N_1406,N_1109,N_1115);
nand U1407 (N_1407,N_1075,N_901);
nand U1408 (N_1408,N_692,N_623);
or U1409 (N_1409,N_674,N_864);
and U1410 (N_1410,N_1151,N_818);
or U1411 (N_1411,N_629,N_890);
or U1412 (N_1412,N_1092,N_813);
and U1413 (N_1413,N_1014,N_646);
or U1414 (N_1414,N_739,N_969);
and U1415 (N_1415,N_949,N_717);
and U1416 (N_1416,N_984,N_895);
or U1417 (N_1417,N_660,N_806);
nand U1418 (N_1418,N_982,N_1077);
and U1419 (N_1419,N_1068,N_998);
nand U1420 (N_1420,N_1088,N_1020);
or U1421 (N_1421,N_1144,N_728);
nor U1422 (N_1422,N_1195,N_985);
and U1423 (N_1423,N_643,N_891);
nand U1424 (N_1424,N_1114,N_605);
nor U1425 (N_1425,N_661,N_1192);
or U1426 (N_1426,N_1131,N_791);
nor U1427 (N_1427,N_1055,N_614);
nor U1428 (N_1428,N_867,N_610);
nand U1429 (N_1429,N_1086,N_858);
or U1430 (N_1430,N_778,N_1027);
and U1431 (N_1431,N_1059,N_1185);
nand U1432 (N_1432,N_1044,N_1179);
xnor U1433 (N_1433,N_910,N_775);
and U1434 (N_1434,N_973,N_834);
nand U1435 (N_1435,N_639,N_803);
nand U1436 (N_1436,N_797,N_799);
nand U1437 (N_1437,N_641,N_648);
nand U1438 (N_1438,N_770,N_658);
nor U1439 (N_1439,N_1031,N_746);
nor U1440 (N_1440,N_1132,N_1016);
and U1441 (N_1441,N_700,N_1186);
nor U1442 (N_1442,N_627,N_814);
and U1443 (N_1443,N_1188,N_789);
and U1444 (N_1444,N_801,N_1122);
nand U1445 (N_1445,N_850,N_794);
nand U1446 (N_1446,N_626,N_616);
nand U1447 (N_1447,N_667,N_829);
nor U1448 (N_1448,N_821,N_726);
or U1449 (N_1449,N_625,N_859);
nand U1450 (N_1450,N_1199,N_1078);
nand U1451 (N_1451,N_1073,N_733);
nor U1452 (N_1452,N_1145,N_730);
xnor U1453 (N_1453,N_905,N_844);
nor U1454 (N_1454,N_857,N_825);
or U1455 (N_1455,N_938,N_1102);
nor U1456 (N_1456,N_1097,N_1081);
xor U1457 (N_1457,N_1004,N_1013);
xnor U1458 (N_1458,N_916,N_663);
and U1459 (N_1459,N_642,N_893);
or U1460 (N_1460,N_716,N_750);
or U1461 (N_1461,N_983,N_839);
xor U1462 (N_1462,N_1191,N_788);
nand U1463 (N_1463,N_1158,N_942);
xor U1464 (N_1464,N_793,N_1089);
xor U1465 (N_1465,N_1093,N_677);
nor U1466 (N_1466,N_1054,N_1005);
nand U1467 (N_1467,N_1168,N_964);
nand U1468 (N_1468,N_622,N_808);
or U1469 (N_1469,N_913,N_612);
or U1470 (N_1470,N_1117,N_712);
and U1471 (N_1471,N_894,N_781);
and U1472 (N_1472,N_927,N_903);
nand U1473 (N_1473,N_678,N_930);
nand U1474 (N_1474,N_1025,N_940);
or U1475 (N_1475,N_725,N_1038);
nor U1476 (N_1476,N_875,N_956);
and U1477 (N_1477,N_779,N_830);
nor U1478 (N_1478,N_1106,N_1010);
nor U1479 (N_1479,N_759,N_673);
xor U1480 (N_1480,N_704,N_1193);
nand U1481 (N_1481,N_925,N_644);
and U1482 (N_1482,N_800,N_997);
and U1483 (N_1483,N_993,N_1153);
nand U1484 (N_1484,N_1138,N_996);
nor U1485 (N_1485,N_807,N_664);
nor U1486 (N_1486,N_1180,N_1136);
nand U1487 (N_1487,N_1065,N_1091);
or U1488 (N_1488,N_758,N_957);
and U1489 (N_1489,N_1178,N_965);
nand U1490 (N_1490,N_714,N_651);
nor U1491 (N_1491,N_784,N_709);
or U1492 (N_1492,N_727,N_963);
xnor U1493 (N_1493,N_706,N_946);
and U1494 (N_1494,N_1051,N_1064);
nand U1495 (N_1495,N_945,N_707);
or U1496 (N_1496,N_936,N_1160);
nand U1497 (N_1497,N_1041,N_860);
nor U1498 (N_1498,N_962,N_911);
nand U1499 (N_1499,N_1107,N_1061);
nor U1500 (N_1500,N_881,N_1163);
xor U1501 (N_1501,N_1127,N_992);
and U1502 (N_1502,N_693,N_988);
nand U1503 (N_1503,N_778,N_732);
and U1504 (N_1504,N_1013,N_633);
nor U1505 (N_1505,N_1003,N_973);
and U1506 (N_1506,N_656,N_844);
and U1507 (N_1507,N_955,N_1187);
nand U1508 (N_1508,N_829,N_661);
and U1509 (N_1509,N_755,N_789);
or U1510 (N_1510,N_731,N_719);
and U1511 (N_1511,N_718,N_1149);
or U1512 (N_1512,N_606,N_755);
or U1513 (N_1513,N_840,N_736);
xor U1514 (N_1514,N_838,N_1160);
nand U1515 (N_1515,N_884,N_1155);
nor U1516 (N_1516,N_937,N_1003);
and U1517 (N_1517,N_1149,N_1008);
xnor U1518 (N_1518,N_1150,N_908);
nor U1519 (N_1519,N_644,N_1029);
or U1520 (N_1520,N_1100,N_1168);
xor U1521 (N_1521,N_838,N_804);
nor U1522 (N_1522,N_670,N_1083);
nor U1523 (N_1523,N_781,N_853);
or U1524 (N_1524,N_797,N_683);
or U1525 (N_1525,N_926,N_879);
nor U1526 (N_1526,N_795,N_636);
or U1527 (N_1527,N_905,N_671);
and U1528 (N_1528,N_718,N_610);
xor U1529 (N_1529,N_878,N_829);
nor U1530 (N_1530,N_742,N_778);
nor U1531 (N_1531,N_795,N_698);
nand U1532 (N_1532,N_730,N_1031);
or U1533 (N_1533,N_1069,N_723);
xor U1534 (N_1534,N_1084,N_1016);
xor U1535 (N_1535,N_861,N_890);
or U1536 (N_1536,N_1012,N_734);
and U1537 (N_1537,N_924,N_695);
or U1538 (N_1538,N_1181,N_952);
nor U1539 (N_1539,N_699,N_836);
and U1540 (N_1540,N_668,N_1114);
and U1541 (N_1541,N_822,N_950);
nand U1542 (N_1542,N_1103,N_857);
nor U1543 (N_1543,N_1094,N_831);
and U1544 (N_1544,N_1190,N_616);
or U1545 (N_1545,N_933,N_692);
nor U1546 (N_1546,N_759,N_1180);
nand U1547 (N_1547,N_802,N_605);
or U1548 (N_1548,N_853,N_1047);
or U1549 (N_1549,N_1045,N_895);
xnor U1550 (N_1550,N_690,N_778);
nand U1551 (N_1551,N_961,N_1123);
nand U1552 (N_1552,N_801,N_957);
and U1553 (N_1553,N_1037,N_1148);
nor U1554 (N_1554,N_1194,N_962);
xnor U1555 (N_1555,N_878,N_1042);
nor U1556 (N_1556,N_943,N_1058);
and U1557 (N_1557,N_1132,N_608);
nor U1558 (N_1558,N_820,N_1040);
nor U1559 (N_1559,N_658,N_1133);
xnor U1560 (N_1560,N_674,N_1036);
nor U1561 (N_1561,N_605,N_1013);
and U1562 (N_1562,N_703,N_1053);
nor U1563 (N_1563,N_644,N_886);
or U1564 (N_1564,N_1001,N_1119);
xor U1565 (N_1565,N_1119,N_644);
or U1566 (N_1566,N_810,N_1185);
or U1567 (N_1567,N_957,N_921);
nor U1568 (N_1568,N_989,N_815);
nor U1569 (N_1569,N_972,N_685);
or U1570 (N_1570,N_666,N_1037);
nor U1571 (N_1571,N_774,N_1020);
nor U1572 (N_1572,N_650,N_818);
nand U1573 (N_1573,N_610,N_1014);
or U1574 (N_1574,N_817,N_677);
nand U1575 (N_1575,N_835,N_799);
and U1576 (N_1576,N_1055,N_848);
or U1577 (N_1577,N_1110,N_607);
nor U1578 (N_1578,N_673,N_841);
nand U1579 (N_1579,N_942,N_933);
xor U1580 (N_1580,N_1047,N_707);
or U1581 (N_1581,N_1022,N_611);
or U1582 (N_1582,N_857,N_1154);
nor U1583 (N_1583,N_756,N_769);
and U1584 (N_1584,N_1151,N_1122);
and U1585 (N_1585,N_1061,N_1062);
xor U1586 (N_1586,N_1173,N_672);
nand U1587 (N_1587,N_686,N_978);
xnor U1588 (N_1588,N_1125,N_888);
or U1589 (N_1589,N_1155,N_1116);
nand U1590 (N_1590,N_1051,N_1154);
xnor U1591 (N_1591,N_687,N_686);
and U1592 (N_1592,N_801,N_841);
or U1593 (N_1593,N_1146,N_624);
xnor U1594 (N_1594,N_769,N_1106);
and U1595 (N_1595,N_769,N_973);
or U1596 (N_1596,N_742,N_801);
or U1597 (N_1597,N_1009,N_620);
or U1598 (N_1598,N_986,N_910);
and U1599 (N_1599,N_798,N_1024);
xnor U1600 (N_1600,N_735,N_1139);
nor U1601 (N_1601,N_1095,N_705);
nor U1602 (N_1602,N_822,N_790);
nand U1603 (N_1603,N_903,N_1144);
or U1604 (N_1604,N_712,N_981);
or U1605 (N_1605,N_1113,N_1046);
nor U1606 (N_1606,N_1073,N_1043);
nor U1607 (N_1607,N_833,N_970);
or U1608 (N_1608,N_977,N_944);
and U1609 (N_1609,N_619,N_889);
and U1610 (N_1610,N_1142,N_780);
nor U1611 (N_1611,N_612,N_1158);
nand U1612 (N_1612,N_1102,N_1110);
nand U1613 (N_1613,N_908,N_647);
nand U1614 (N_1614,N_726,N_648);
nand U1615 (N_1615,N_633,N_672);
nor U1616 (N_1616,N_1147,N_640);
or U1617 (N_1617,N_1146,N_1160);
or U1618 (N_1618,N_1001,N_1024);
and U1619 (N_1619,N_979,N_876);
and U1620 (N_1620,N_900,N_908);
nand U1621 (N_1621,N_809,N_768);
nor U1622 (N_1622,N_860,N_1030);
and U1623 (N_1623,N_1168,N_751);
nor U1624 (N_1624,N_1158,N_618);
and U1625 (N_1625,N_881,N_1056);
nand U1626 (N_1626,N_1099,N_998);
and U1627 (N_1627,N_1191,N_1070);
nor U1628 (N_1628,N_933,N_1021);
and U1629 (N_1629,N_1188,N_834);
nand U1630 (N_1630,N_955,N_1018);
or U1631 (N_1631,N_879,N_700);
or U1632 (N_1632,N_1129,N_882);
xnor U1633 (N_1633,N_764,N_1070);
nand U1634 (N_1634,N_1110,N_1169);
or U1635 (N_1635,N_1162,N_1072);
nor U1636 (N_1636,N_1023,N_1181);
nand U1637 (N_1637,N_1080,N_1070);
nor U1638 (N_1638,N_878,N_970);
nand U1639 (N_1639,N_1156,N_888);
nand U1640 (N_1640,N_636,N_1057);
nand U1641 (N_1641,N_732,N_861);
xor U1642 (N_1642,N_901,N_827);
or U1643 (N_1643,N_1047,N_1049);
and U1644 (N_1644,N_1085,N_1063);
or U1645 (N_1645,N_1025,N_671);
or U1646 (N_1646,N_884,N_1017);
nor U1647 (N_1647,N_989,N_1012);
and U1648 (N_1648,N_1137,N_1124);
and U1649 (N_1649,N_913,N_1033);
or U1650 (N_1650,N_1075,N_1082);
nor U1651 (N_1651,N_715,N_603);
and U1652 (N_1652,N_847,N_886);
and U1653 (N_1653,N_791,N_1145);
or U1654 (N_1654,N_994,N_1065);
nor U1655 (N_1655,N_985,N_824);
and U1656 (N_1656,N_1113,N_1168);
nor U1657 (N_1657,N_740,N_853);
or U1658 (N_1658,N_857,N_984);
nor U1659 (N_1659,N_840,N_1197);
nor U1660 (N_1660,N_885,N_668);
or U1661 (N_1661,N_798,N_1042);
or U1662 (N_1662,N_864,N_775);
and U1663 (N_1663,N_677,N_1195);
or U1664 (N_1664,N_1033,N_844);
or U1665 (N_1665,N_607,N_872);
and U1666 (N_1666,N_793,N_932);
and U1667 (N_1667,N_1196,N_908);
nor U1668 (N_1668,N_1074,N_861);
xnor U1669 (N_1669,N_1016,N_821);
and U1670 (N_1670,N_875,N_884);
and U1671 (N_1671,N_717,N_790);
or U1672 (N_1672,N_800,N_998);
nand U1673 (N_1673,N_853,N_652);
and U1674 (N_1674,N_610,N_979);
and U1675 (N_1675,N_659,N_603);
or U1676 (N_1676,N_731,N_760);
and U1677 (N_1677,N_874,N_1133);
or U1678 (N_1678,N_1048,N_949);
nand U1679 (N_1679,N_641,N_734);
and U1680 (N_1680,N_956,N_1156);
nand U1681 (N_1681,N_1178,N_760);
nor U1682 (N_1682,N_1189,N_1196);
and U1683 (N_1683,N_1078,N_1195);
and U1684 (N_1684,N_615,N_976);
nor U1685 (N_1685,N_795,N_858);
nand U1686 (N_1686,N_734,N_715);
xor U1687 (N_1687,N_1024,N_868);
xnor U1688 (N_1688,N_1151,N_1163);
and U1689 (N_1689,N_636,N_793);
or U1690 (N_1690,N_812,N_1171);
and U1691 (N_1691,N_909,N_1049);
nand U1692 (N_1692,N_908,N_1188);
nand U1693 (N_1693,N_1050,N_662);
or U1694 (N_1694,N_966,N_1132);
nand U1695 (N_1695,N_783,N_966);
nor U1696 (N_1696,N_1124,N_1158);
nand U1697 (N_1697,N_973,N_1113);
nor U1698 (N_1698,N_835,N_622);
and U1699 (N_1699,N_872,N_889);
nand U1700 (N_1700,N_620,N_740);
and U1701 (N_1701,N_1153,N_625);
or U1702 (N_1702,N_1140,N_1171);
nand U1703 (N_1703,N_809,N_709);
and U1704 (N_1704,N_635,N_896);
or U1705 (N_1705,N_1182,N_1119);
nor U1706 (N_1706,N_805,N_730);
nand U1707 (N_1707,N_1164,N_900);
nand U1708 (N_1708,N_1116,N_1055);
nand U1709 (N_1709,N_783,N_1194);
or U1710 (N_1710,N_1019,N_630);
nor U1711 (N_1711,N_956,N_1104);
nor U1712 (N_1712,N_1002,N_980);
and U1713 (N_1713,N_1111,N_1128);
or U1714 (N_1714,N_861,N_1136);
nor U1715 (N_1715,N_639,N_703);
or U1716 (N_1716,N_1114,N_1154);
or U1717 (N_1717,N_852,N_1091);
nor U1718 (N_1718,N_1017,N_1109);
nor U1719 (N_1719,N_1102,N_903);
or U1720 (N_1720,N_893,N_749);
or U1721 (N_1721,N_1136,N_975);
nor U1722 (N_1722,N_957,N_671);
or U1723 (N_1723,N_1187,N_694);
nor U1724 (N_1724,N_1138,N_1110);
nand U1725 (N_1725,N_779,N_1107);
or U1726 (N_1726,N_1061,N_763);
nand U1727 (N_1727,N_1001,N_1175);
nand U1728 (N_1728,N_754,N_822);
and U1729 (N_1729,N_703,N_685);
nand U1730 (N_1730,N_916,N_666);
nor U1731 (N_1731,N_970,N_1089);
nand U1732 (N_1732,N_1064,N_1027);
nand U1733 (N_1733,N_781,N_1157);
nor U1734 (N_1734,N_731,N_1119);
and U1735 (N_1735,N_920,N_861);
nand U1736 (N_1736,N_833,N_707);
or U1737 (N_1737,N_869,N_700);
or U1738 (N_1738,N_688,N_1105);
nand U1739 (N_1739,N_1081,N_830);
and U1740 (N_1740,N_992,N_666);
nand U1741 (N_1741,N_808,N_1120);
or U1742 (N_1742,N_1054,N_1052);
nor U1743 (N_1743,N_1039,N_1150);
nand U1744 (N_1744,N_942,N_1059);
xor U1745 (N_1745,N_614,N_825);
nand U1746 (N_1746,N_922,N_971);
nor U1747 (N_1747,N_676,N_620);
nand U1748 (N_1748,N_653,N_953);
xnor U1749 (N_1749,N_814,N_912);
or U1750 (N_1750,N_1086,N_682);
nand U1751 (N_1751,N_1064,N_675);
and U1752 (N_1752,N_1099,N_787);
nor U1753 (N_1753,N_1002,N_1122);
nor U1754 (N_1754,N_1069,N_1062);
nand U1755 (N_1755,N_774,N_1000);
nand U1756 (N_1756,N_617,N_850);
xnor U1757 (N_1757,N_850,N_842);
or U1758 (N_1758,N_832,N_890);
or U1759 (N_1759,N_910,N_613);
nand U1760 (N_1760,N_706,N_917);
xor U1761 (N_1761,N_926,N_1153);
xor U1762 (N_1762,N_1192,N_1105);
nand U1763 (N_1763,N_1029,N_700);
and U1764 (N_1764,N_886,N_784);
and U1765 (N_1765,N_975,N_670);
nand U1766 (N_1766,N_986,N_1129);
and U1767 (N_1767,N_926,N_834);
nor U1768 (N_1768,N_1056,N_991);
nand U1769 (N_1769,N_1048,N_716);
xor U1770 (N_1770,N_1151,N_797);
or U1771 (N_1771,N_745,N_727);
nand U1772 (N_1772,N_812,N_801);
nand U1773 (N_1773,N_683,N_1111);
and U1774 (N_1774,N_1129,N_906);
or U1775 (N_1775,N_704,N_884);
or U1776 (N_1776,N_815,N_1016);
nor U1777 (N_1777,N_1160,N_835);
nand U1778 (N_1778,N_625,N_976);
nand U1779 (N_1779,N_1063,N_961);
nand U1780 (N_1780,N_990,N_986);
nand U1781 (N_1781,N_788,N_625);
and U1782 (N_1782,N_1150,N_740);
nor U1783 (N_1783,N_764,N_685);
nor U1784 (N_1784,N_890,N_778);
and U1785 (N_1785,N_823,N_639);
nor U1786 (N_1786,N_816,N_1012);
nor U1787 (N_1787,N_1187,N_816);
or U1788 (N_1788,N_843,N_1147);
or U1789 (N_1789,N_1177,N_1060);
nor U1790 (N_1790,N_726,N_744);
nor U1791 (N_1791,N_655,N_815);
nor U1792 (N_1792,N_853,N_1089);
nor U1793 (N_1793,N_1125,N_923);
nor U1794 (N_1794,N_825,N_1114);
nor U1795 (N_1795,N_708,N_962);
nor U1796 (N_1796,N_606,N_1012);
and U1797 (N_1797,N_728,N_836);
xnor U1798 (N_1798,N_894,N_851);
nand U1799 (N_1799,N_796,N_700);
nor U1800 (N_1800,N_1768,N_1580);
and U1801 (N_1801,N_1358,N_1379);
xnor U1802 (N_1802,N_1417,N_1558);
or U1803 (N_1803,N_1633,N_1649);
or U1804 (N_1804,N_1583,N_1233);
xor U1805 (N_1805,N_1632,N_1458);
xnor U1806 (N_1806,N_1299,N_1241);
and U1807 (N_1807,N_1792,N_1711);
or U1808 (N_1808,N_1409,N_1537);
and U1809 (N_1809,N_1574,N_1582);
and U1810 (N_1810,N_1392,N_1466);
nand U1811 (N_1811,N_1626,N_1476);
and U1812 (N_1812,N_1706,N_1544);
or U1813 (N_1813,N_1664,N_1590);
and U1814 (N_1814,N_1290,N_1213);
or U1815 (N_1815,N_1346,N_1552);
nand U1816 (N_1816,N_1694,N_1521);
or U1817 (N_1817,N_1453,N_1545);
or U1818 (N_1818,N_1306,N_1645);
and U1819 (N_1819,N_1576,N_1553);
nor U1820 (N_1820,N_1204,N_1375);
or U1821 (N_1821,N_1469,N_1209);
and U1822 (N_1822,N_1651,N_1514);
or U1823 (N_1823,N_1389,N_1609);
and U1824 (N_1824,N_1765,N_1797);
nor U1825 (N_1825,N_1418,N_1620);
or U1826 (N_1826,N_1430,N_1349);
nor U1827 (N_1827,N_1762,N_1294);
nand U1828 (N_1828,N_1527,N_1281);
nor U1829 (N_1829,N_1634,N_1787);
nand U1830 (N_1830,N_1260,N_1266);
xor U1831 (N_1831,N_1619,N_1660);
or U1832 (N_1832,N_1330,N_1612);
xnor U1833 (N_1833,N_1665,N_1681);
or U1834 (N_1834,N_1309,N_1261);
nor U1835 (N_1835,N_1437,N_1723);
nand U1836 (N_1836,N_1699,N_1618);
nor U1837 (N_1837,N_1601,N_1473);
nor U1838 (N_1838,N_1311,N_1441);
nor U1839 (N_1839,N_1487,N_1411);
nor U1840 (N_1840,N_1229,N_1230);
and U1841 (N_1841,N_1408,N_1523);
nor U1842 (N_1842,N_1502,N_1220);
or U1843 (N_1843,N_1225,N_1308);
nor U1844 (N_1844,N_1697,N_1490);
or U1845 (N_1845,N_1368,N_1796);
xnor U1846 (N_1846,N_1231,N_1207);
xnor U1847 (N_1847,N_1508,N_1679);
and U1848 (N_1848,N_1273,N_1650);
nor U1849 (N_1849,N_1695,N_1313);
and U1850 (N_1850,N_1424,N_1480);
nor U1851 (N_1851,N_1530,N_1591);
nor U1852 (N_1852,N_1685,N_1572);
nand U1853 (N_1853,N_1485,N_1594);
xnor U1854 (N_1854,N_1596,N_1350);
nor U1855 (N_1855,N_1472,N_1690);
xor U1856 (N_1856,N_1321,N_1352);
or U1857 (N_1857,N_1775,N_1218);
nand U1858 (N_1858,N_1539,N_1267);
nor U1859 (N_1859,N_1735,N_1316);
and U1860 (N_1860,N_1746,N_1643);
or U1861 (N_1861,N_1464,N_1718);
nor U1862 (N_1862,N_1662,N_1646);
or U1863 (N_1863,N_1378,N_1394);
and U1864 (N_1864,N_1733,N_1743);
or U1865 (N_1865,N_1698,N_1211);
xnor U1866 (N_1866,N_1492,N_1438);
nor U1867 (N_1867,N_1784,N_1343);
and U1868 (N_1868,N_1700,N_1246);
nor U1869 (N_1869,N_1390,N_1707);
nand U1870 (N_1870,N_1377,N_1237);
xor U1871 (N_1871,N_1446,N_1513);
nor U1872 (N_1872,N_1728,N_1467);
and U1873 (N_1873,N_1372,N_1250);
and U1874 (N_1874,N_1658,N_1603);
or U1875 (N_1875,N_1347,N_1510);
nor U1876 (N_1876,N_1770,N_1624);
or U1877 (N_1877,N_1280,N_1630);
and U1878 (N_1878,N_1741,N_1341);
nor U1879 (N_1879,N_1327,N_1731);
or U1880 (N_1880,N_1355,N_1423);
and U1881 (N_1881,N_1400,N_1439);
nand U1882 (N_1882,N_1263,N_1406);
or U1883 (N_1883,N_1625,N_1428);
or U1884 (N_1884,N_1500,N_1274);
nor U1885 (N_1885,N_1791,N_1575);
nor U1886 (N_1886,N_1291,N_1286);
nor U1887 (N_1887,N_1676,N_1702);
and U1888 (N_1888,N_1564,N_1324);
nand U1889 (N_1889,N_1251,N_1482);
nor U1890 (N_1890,N_1614,N_1243);
or U1891 (N_1891,N_1738,N_1205);
nand U1892 (N_1892,N_1270,N_1647);
xor U1893 (N_1893,N_1318,N_1640);
or U1894 (N_1894,N_1226,N_1240);
or U1895 (N_1895,N_1786,N_1724);
and U1896 (N_1896,N_1616,N_1516);
or U1897 (N_1897,N_1666,N_1520);
nand U1898 (N_1898,N_1200,N_1669);
and U1899 (N_1899,N_1611,N_1714);
nor U1900 (N_1900,N_1440,N_1322);
nor U1901 (N_1901,N_1475,N_1203);
nand U1902 (N_1902,N_1344,N_1531);
or U1903 (N_1903,N_1568,N_1471);
or U1904 (N_1904,N_1479,N_1604);
nand U1905 (N_1905,N_1252,N_1444);
and U1906 (N_1906,N_1641,N_1518);
and U1907 (N_1907,N_1635,N_1317);
and U1908 (N_1908,N_1776,N_1675);
or U1909 (N_1909,N_1474,N_1283);
or U1910 (N_1910,N_1336,N_1592);
xor U1911 (N_1911,N_1534,N_1704);
nor U1912 (N_1912,N_1498,N_1692);
nand U1913 (N_1913,N_1259,N_1771);
nand U1914 (N_1914,N_1528,N_1331);
and U1915 (N_1915,N_1285,N_1570);
nor U1916 (N_1916,N_1405,N_1688);
and U1917 (N_1917,N_1566,N_1410);
and U1918 (N_1918,N_1247,N_1319);
or U1919 (N_1919,N_1427,N_1747);
nor U1920 (N_1920,N_1745,N_1454);
nor U1921 (N_1921,N_1465,N_1262);
and U1922 (N_1922,N_1452,N_1680);
nor U1923 (N_1923,N_1362,N_1788);
and U1924 (N_1924,N_1600,N_1223);
or U1925 (N_1925,N_1772,N_1555);
xor U1926 (N_1926,N_1351,N_1434);
and U1927 (N_1927,N_1238,N_1366);
nor U1928 (N_1928,N_1540,N_1538);
and U1929 (N_1929,N_1627,N_1505);
and U1930 (N_1930,N_1550,N_1637);
and U1931 (N_1931,N_1648,N_1754);
and U1932 (N_1932,N_1391,N_1468);
xor U1933 (N_1933,N_1329,N_1586);
nor U1934 (N_1934,N_1264,N_1753);
and U1935 (N_1935,N_1636,N_1774);
nand U1936 (N_1936,N_1388,N_1429);
or U1937 (N_1937,N_1345,N_1386);
xor U1938 (N_1938,N_1749,N_1760);
and U1939 (N_1939,N_1657,N_1548);
and U1940 (N_1940,N_1254,N_1461);
nor U1941 (N_1941,N_1216,N_1376);
nand U1942 (N_1942,N_1742,N_1668);
and U1943 (N_1943,N_1256,N_1551);
and U1944 (N_1944,N_1442,N_1393);
nand U1945 (N_1945,N_1224,N_1221);
nand U1946 (N_1946,N_1507,N_1549);
nor U1947 (N_1947,N_1701,N_1320);
or U1948 (N_1948,N_1210,N_1496);
and U1949 (N_1949,N_1484,N_1622);
nand U1950 (N_1950,N_1275,N_1597);
nand U1951 (N_1951,N_1790,N_1593);
or U1952 (N_1952,N_1374,N_1295);
or U1953 (N_1953,N_1232,N_1524);
nor U1954 (N_1954,N_1503,N_1310);
nand U1955 (N_1955,N_1638,N_1248);
nand U1956 (N_1956,N_1268,N_1778);
nor U1957 (N_1957,N_1677,N_1541);
nor U1958 (N_1958,N_1631,N_1412);
and U1959 (N_1959,N_1682,N_1559);
and U1960 (N_1960,N_1435,N_1615);
or U1961 (N_1961,N_1722,N_1421);
and U1962 (N_1962,N_1504,N_1323);
and U1963 (N_1963,N_1332,N_1269);
or U1964 (N_1964,N_1371,N_1721);
and U1965 (N_1965,N_1272,N_1739);
nand U1966 (N_1966,N_1312,N_1457);
and U1967 (N_1967,N_1511,N_1526);
or U1968 (N_1968,N_1659,N_1732);
or U1969 (N_1969,N_1342,N_1445);
nor U1970 (N_1970,N_1716,N_1562);
and U1971 (N_1971,N_1655,N_1613);
nand U1972 (N_1972,N_1767,N_1740);
or U1973 (N_1973,N_1509,N_1436);
and U1974 (N_1974,N_1258,N_1383);
nor U1975 (N_1975,N_1348,N_1585);
and U1976 (N_1976,N_1420,N_1443);
and U1977 (N_1977,N_1703,N_1307);
nor U1978 (N_1978,N_1470,N_1214);
nor U1979 (N_1979,N_1384,N_1696);
and U1980 (N_1980,N_1277,N_1244);
nand U1981 (N_1981,N_1654,N_1684);
or U1982 (N_1982,N_1397,N_1506);
nor U1983 (N_1983,N_1554,N_1486);
and U1984 (N_1984,N_1795,N_1799);
nand U1985 (N_1985,N_1414,N_1565);
or U1986 (N_1986,N_1426,N_1595);
nor U1987 (N_1987,N_1736,N_1517);
nor U1988 (N_1988,N_1305,N_1396);
or U1989 (N_1989,N_1756,N_1328);
or U1990 (N_1990,N_1380,N_1543);
nor U1991 (N_1991,N_1253,N_1673);
or U1992 (N_1992,N_1606,N_1292);
and U1993 (N_1993,N_1628,N_1720);
xnor U1994 (N_1994,N_1432,N_1413);
and U1995 (N_1995,N_1255,N_1717);
nand U1996 (N_1996,N_1278,N_1302);
or U1997 (N_1997,N_1757,N_1729);
nand U1998 (N_1998,N_1431,N_1367);
and U1999 (N_1999,N_1265,N_1661);
and U2000 (N_2000,N_1584,N_1569);
nand U2001 (N_2001,N_1573,N_1578);
or U2002 (N_2002,N_1782,N_1691);
and U2003 (N_2003,N_1556,N_1759);
or U2004 (N_2004,N_1338,N_1678);
and U2005 (N_2005,N_1712,N_1588);
nand U2006 (N_2006,N_1727,N_1547);
nand U2007 (N_2007,N_1354,N_1683);
or U2008 (N_2008,N_1755,N_1279);
and U2009 (N_2009,N_1215,N_1512);
nand U2010 (N_2010,N_1236,N_1610);
and U2011 (N_2011,N_1373,N_1361);
or U2012 (N_2012,N_1671,N_1402);
and U2013 (N_2013,N_1201,N_1644);
and U2014 (N_2014,N_1239,N_1730);
nor U2015 (N_2015,N_1687,N_1422);
nor U2016 (N_2016,N_1395,N_1761);
nand U2017 (N_2017,N_1663,N_1363);
and U2018 (N_2018,N_1744,N_1304);
nand U2019 (N_2019,N_1546,N_1623);
nand U2020 (N_2020,N_1710,N_1780);
and U2021 (N_2021,N_1777,N_1561);
nor U2022 (N_2022,N_1357,N_1222);
or U2023 (N_2023,N_1617,N_1370);
nand U2024 (N_2024,N_1621,N_1783);
and U2025 (N_2025,N_1288,N_1416);
or U2026 (N_2026,N_1491,N_1709);
nor U2027 (N_2027,N_1715,N_1581);
nand U2028 (N_2028,N_1401,N_1451);
or U2029 (N_2029,N_1672,N_1705);
nand U2030 (N_2030,N_1629,N_1748);
nand U2031 (N_2031,N_1202,N_1769);
nor U2032 (N_2032,N_1208,N_1462);
nand U2033 (N_2033,N_1234,N_1276);
and U2034 (N_2034,N_1257,N_1525);
xnor U2035 (N_2035,N_1497,N_1501);
nor U2036 (N_2036,N_1607,N_1608);
nor U2037 (N_2037,N_1382,N_1798);
nor U2038 (N_2038,N_1519,N_1535);
nand U2039 (N_2039,N_1488,N_1750);
nor U2040 (N_2040,N_1249,N_1766);
xnor U2041 (N_2041,N_1602,N_1404);
or U2042 (N_2042,N_1719,N_1653);
or U2043 (N_2043,N_1489,N_1340);
nand U2044 (N_2044,N_1477,N_1789);
nand U2045 (N_2045,N_1536,N_1301);
nor U2046 (N_2046,N_1334,N_1228);
xor U2047 (N_2047,N_1450,N_1642);
nand U2048 (N_2048,N_1781,N_1483);
xnor U2049 (N_2049,N_1693,N_1314);
nor U2050 (N_2050,N_1563,N_1785);
and U2051 (N_2051,N_1271,N_1300);
nand U2052 (N_2052,N_1571,N_1325);
nand U2053 (N_2053,N_1726,N_1577);
nor U2054 (N_2054,N_1763,N_1764);
nor U2055 (N_2055,N_1557,N_1656);
nand U2056 (N_2056,N_1708,N_1403);
and U2057 (N_2057,N_1326,N_1219);
or U2058 (N_2058,N_1407,N_1639);
or U2059 (N_2059,N_1399,N_1419);
nand U2060 (N_2060,N_1282,N_1449);
and U2061 (N_2061,N_1364,N_1289);
or U2062 (N_2062,N_1779,N_1455);
and U2063 (N_2063,N_1456,N_1293);
or U2064 (N_2064,N_1459,N_1359);
xor U2065 (N_2065,N_1460,N_1532);
and U2066 (N_2066,N_1560,N_1499);
nand U2067 (N_2067,N_1385,N_1734);
nor U2068 (N_2068,N_1758,N_1245);
nand U2069 (N_2069,N_1751,N_1533);
or U2070 (N_2070,N_1579,N_1433);
and U2071 (N_2071,N_1493,N_1713);
or U2072 (N_2072,N_1542,N_1478);
nand U2073 (N_2073,N_1737,N_1335);
or U2074 (N_2074,N_1587,N_1235);
nor U2075 (N_2075,N_1773,N_1353);
nor U2076 (N_2076,N_1315,N_1356);
xnor U2077 (N_2077,N_1674,N_1303);
or U2078 (N_2078,N_1689,N_1670);
nand U2079 (N_2079,N_1667,N_1598);
and U2080 (N_2080,N_1686,N_1337);
nand U2081 (N_2081,N_1481,N_1333);
and U2082 (N_2082,N_1387,N_1425);
and U2083 (N_2083,N_1339,N_1369);
nor U2084 (N_2084,N_1360,N_1447);
xor U2085 (N_2085,N_1752,N_1448);
nand U2086 (N_2086,N_1381,N_1242);
nand U2087 (N_2087,N_1463,N_1297);
nand U2088 (N_2088,N_1567,N_1522);
xnor U2089 (N_2089,N_1793,N_1515);
or U2090 (N_2090,N_1398,N_1206);
or U2091 (N_2091,N_1599,N_1494);
or U2092 (N_2092,N_1589,N_1296);
xnor U2093 (N_2093,N_1365,N_1212);
and U2094 (N_2094,N_1794,N_1227);
nand U2095 (N_2095,N_1298,N_1605);
xnor U2096 (N_2096,N_1495,N_1415);
nor U2097 (N_2097,N_1652,N_1287);
or U2098 (N_2098,N_1725,N_1529);
and U2099 (N_2099,N_1284,N_1217);
and U2100 (N_2100,N_1460,N_1463);
and U2101 (N_2101,N_1200,N_1753);
or U2102 (N_2102,N_1210,N_1582);
and U2103 (N_2103,N_1736,N_1274);
or U2104 (N_2104,N_1242,N_1470);
nor U2105 (N_2105,N_1248,N_1354);
nor U2106 (N_2106,N_1214,N_1382);
xnor U2107 (N_2107,N_1320,N_1589);
or U2108 (N_2108,N_1414,N_1786);
or U2109 (N_2109,N_1541,N_1455);
nor U2110 (N_2110,N_1355,N_1377);
nand U2111 (N_2111,N_1464,N_1463);
and U2112 (N_2112,N_1373,N_1433);
nand U2113 (N_2113,N_1451,N_1247);
and U2114 (N_2114,N_1590,N_1489);
and U2115 (N_2115,N_1211,N_1277);
and U2116 (N_2116,N_1294,N_1225);
nand U2117 (N_2117,N_1771,N_1688);
or U2118 (N_2118,N_1283,N_1675);
and U2119 (N_2119,N_1281,N_1761);
nor U2120 (N_2120,N_1722,N_1560);
nor U2121 (N_2121,N_1730,N_1426);
nor U2122 (N_2122,N_1399,N_1342);
or U2123 (N_2123,N_1216,N_1790);
nand U2124 (N_2124,N_1774,N_1567);
nand U2125 (N_2125,N_1430,N_1281);
nand U2126 (N_2126,N_1518,N_1281);
xor U2127 (N_2127,N_1683,N_1632);
nor U2128 (N_2128,N_1498,N_1777);
or U2129 (N_2129,N_1416,N_1455);
nor U2130 (N_2130,N_1487,N_1567);
nand U2131 (N_2131,N_1279,N_1329);
nand U2132 (N_2132,N_1304,N_1731);
nor U2133 (N_2133,N_1472,N_1722);
nor U2134 (N_2134,N_1227,N_1605);
or U2135 (N_2135,N_1709,N_1431);
or U2136 (N_2136,N_1359,N_1665);
nand U2137 (N_2137,N_1341,N_1597);
and U2138 (N_2138,N_1595,N_1318);
nor U2139 (N_2139,N_1292,N_1329);
nand U2140 (N_2140,N_1448,N_1354);
xnor U2141 (N_2141,N_1461,N_1355);
nor U2142 (N_2142,N_1351,N_1445);
or U2143 (N_2143,N_1627,N_1364);
nand U2144 (N_2144,N_1712,N_1378);
xnor U2145 (N_2145,N_1610,N_1776);
xnor U2146 (N_2146,N_1737,N_1777);
nor U2147 (N_2147,N_1357,N_1531);
or U2148 (N_2148,N_1215,N_1300);
nand U2149 (N_2149,N_1512,N_1601);
xor U2150 (N_2150,N_1483,N_1433);
and U2151 (N_2151,N_1390,N_1597);
and U2152 (N_2152,N_1744,N_1669);
xor U2153 (N_2153,N_1480,N_1529);
nand U2154 (N_2154,N_1270,N_1560);
and U2155 (N_2155,N_1621,N_1221);
nor U2156 (N_2156,N_1669,N_1761);
nor U2157 (N_2157,N_1224,N_1751);
nand U2158 (N_2158,N_1766,N_1469);
or U2159 (N_2159,N_1730,N_1223);
or U2160 (N_2160,N_1646,N_1764);
and U2161 (N_2161,N_1488,N_1698);
xor U2162 (N_2162,N_1573,N_1418);
and U2163 (N_2163,N_1567,N_1374);
and U2164 (N_2164,N_1247,N_1484);
nor U2165 (N_2165,N_1579,N_1489);
nor U2166 (N_2166,N_1748,N_1564);
nor U2167 (N_2167,N_1298,N_1545);
and U2168 (N_2168,N_1392,N_1495);
and U2169 (N_2169,N_1486,N_1736);
xor U2170 (N_2170,N_1682,N_1506);
and U2171 (N_2171,N_1225,N_1655);
or U2172 (N_2172,N_1483,N_1614);
nor U2173 (N_2173,N_1227,N_1466);
or U2174 (N_2174,N_1791,N_1733);
or U2175 (N_2175,N_1333,N_1461);
and U2176 (N_2176,N_1700,N_1556);
and U2177 (N_2177,N_1301,N_1256);
xor U2178 (N_2178,N_1471,N_1202);
or U2179 (N_2179,N_1581,N_1232);
nand U2180 (N_2180,N_1237,N_1388);
nor U2181 (N_2181,N_1495,N_1633);
xnor U2182 (N_2182,N_1279,N_1637);
xor U2183 (N_2183,N_1258,N_1321);
nor U2184 (N_2184,N_1671,N_1278);
nand U2185 (N_2185,N_1285,N_1302);
nor U2186 (N_2186,N_1721,N_1241);
nand U2187 (N_2187,N_1306,N_1618);
nor U2188 (N_2188,N_1688,N_1687);
nor U2189 (N_2189,N_1241,N_1300);
or U2190 (N_2190,N_1324,N_1606);
or U2191 (N_2191,N_1582,N_1441);
nand U2192 (N_2192,N_1685,N_1788);
and U2193 (N_2193,N_1610,N_1586);
and U2194 (N_2194,N_1271,N_1716);
nor U2195 (N_2195,N_1386,N_1243);
or U2196 (N_2196,N_1459,N_1590);
and U2197 (N_2197,N_1382,N_1418);
or U2198 (N_2198,N_1436,N_1336);
nor U2199 (N_2199,N_1540,N_1533);
or U2200 (N_2200,N_1324,N_1384);
or U2201 (N_2201,N_1564,N_1306);
or U2202 (N_2202,N_1699,N_1579);
nand U2203 (N_2203,N_1621,N_1719);
and U2204 (N_2204,N_1716,N_1397);
nor U2205 (N_2205,N_1203,N_1241);
and U2206 (N_2206,N_1738,N_1650);
nor U2207 (N_2207,N_1693,N_1222);
or U2208 (N_2208,N_1616,N_1795);
and U2209 (N_2209,N_1746,N_1535);
nand U2210 (N_2210,N_1544,N_1440);
xnor U2211 (N_2211,N_1540,N_1592);
nand U2212 (N_2212,N_1529,N_1647);
xor U2213 (N_2213,N_1235,N_1602);
or U2214 (N_2214,N_1370,N_1407);
nand U2215 (N_2215,N_1337,N_1601);
or U2216 (N_2216,N_1565,N_1659);
or U2217 (N_2217,N_1411,N_1700);
or U2218 (N_2218,N_1220,N_1363);
nand U2219 (N_2219,N_1773,N_1682);
or U2220 (N_2220,N_1655,N_1698);
nand U2221 (N_2221,N_1392,N_1213);
xor U2222 (N_2222,N_1743,N_1250);
nand U2223 (N_2223,N_1267,N_1487);
or U2224 (N_2224,N_1254,N_1419);
nor U2225 (N_2225,N_1679,N_1390);
and U2226 (N_2226,N_1386,N_1317);
nor U2227 (N_2227,N_1761,N_1379);
nand U2228 (N_2228,N_1510,N_1221);
and U2229 (N_2229,N_1542,N_1782);
nor U2230 (N_2230,N_1243,N_1404);
and U2231 (N_2231,N_1322,N_1668);
nand U2232 (N_2232,N_1257,N_1260);
and U2233 (N_2233,N_1579,N_1661);
or U2234 (N_2234,N_1582,N_1379);
xnor U2235 (N_2235,N_1322,N_1358);
or U2236 (N_2236,N_1680,N_1694);
xor U2237 (N_2237,N_1358,N_1720);
and U2238 (N_2238,N_1395,N_1327);
and U2239 (N_2239,N_1503,N_1383);
nor U2240 (N_2240,N_1589,N_1770);
and U2241 (N_2241,N_1566,N_1646);
and U2242 (N_2242,N_1401,N_1386);
nand U2243 (N_2243,N_1563,N_1520);
or U2244 (N_2244,N_1597,N_1455);
and U2245 (N_2245,N_1230,N_1221);
and U2246 (N_2246,N_1501,N_1745);
nand U2247 (N_2247,N_1582,N_1350);
nand U2248 (N_2248,N_1567,N_1410);
nor U2249 (N_2249,N_1228,N_1393);
or U2250 (N_2250,N_1509,N_1435);
nor U2251 (N_2251,N_1341,N_1443);
nor U2252 (N_2252,N_1392,N_1458);
or U2253 (N_2253,N_1478,N_1265);
nand U2254 (N_2254,N_1271,N_1574);
or U2255 (N_2255,N_1771,N_1303);
and U2256 (N_2256,N_1792,N_1247);
or U2257 (N_2257,N_1333,N_1272);
and U2258 (N_2258,N_1656,N_1625);
or U2259 (N_2259,N_1794,N_1760);
nand U2260 (N_2260,N_1551,N_1640);
nor U2261 (N_2261,N_1251,N_1232);
nand U2262 (N_2262,N_1291,N_1395);
nor U2263 (N_2263,N_1223,N_1639);
nor U2264 (N_2264,N_1491,N_1330);
xor U2265 (N_2265,N_1515,N_1334);
nor U2266 (N_2266,N_1779,N_1445);
and U2267 (N_2267,N_1594,N_1756);
nand U2268 (N_2268,N_1247,N_1772);
or U2269 (N_2269,N_1454,N_1384);
and U2270 (N_2270,N_1717,N_1212);
and U2271 (N_2271,N_1507,N_1641);
or U2272 (N_2272,N_1779,N_1410);
nor U2273 (N_2273,N_1458,N_1709);
nand U2274 (N_2274,N_1586,N_1342);
or U2275 (N_2275,N_1277,N_1300);
nand U2276 (N_2276,N_1683,N_1448);
and U2277 (N_2277,N_1235,N_1306);
nand U2278 (N_2278,N_1667,N_1671);
nor U2279 (N_2279,N_1714,N_1790);
nor U2280 (N_2280,N_1593,N_1266);
and U2281 (N_2281,N_1505,N_1649);
nor U2282 (N_2282,N_1496,N_1228);
nor U2283 (N_2283,N_1546,N_1481);
and U2284 (N_2284,N_1737,N_1695);
nand U2285 (N_2285,N_1739,N_1310);
nor U2286 (N_2286,N_1319,N_1209);
nand U2287 (N_2287,N_1739,N_1445);
nand U2288 (N_2288,N_1574,N_1475);
or U2289 (N_2289,N_1216,N_1435);
or U2290 (N_2290,N_1448,N_1420);
nand U2291 (N_2291,N_1383,N_1564);
nand U2292 (N_2292,N_1602,N_1524);
nand U2293 (N_2293,N_1681,N_1440);
or U2294 (N_2294,N_1462,N_1380);
nand U2295 (N_2295,N_1678,N_1296);
xor U2296 (N_2296,N_1499,N_1725);
nor U2297 (N_2297,N_1751,N_1400);
and U2298 (N_2298,N_1336,N_1779);
nand U2299 (N_2299,N_1498,N_1460);
or U2300 (N_2300,N_1693,N_1412);
nand U2301 (N_2301,N_1323,N_1635);
nor U2302 (N_2302,N_1764,N_1615);
nand U2303 (N_2303,N_1350,N_1484);
and U2304 (N_2304,N_1633,N_1380);
and U2305 (N_2305,N_1305,N_1386);
and U2306 (N_2306,N_1365,N_1568);
and U2307 (N_2307,N_1654,N_1466);
xnor U2308 (N_2308,N_1224,N_1668);
nand U2309 (N_2309,N_1529,N_1225);
and U2310 (N_2310,N_1723,N_1224);
or U2311 (N_2311,N_1259,N_1207);
nor U2312 (N_2312,N_1485,N_1237);
and U2313 (N_2313,N_1422,N_1629);
xnor U2314 (N_2314,N_1650,N_1711);
xor U2315 (N_2315,N_1410,N_1677);
nor U2316 (N_2316,N_1568,N_1763);
nand U2317 (N_2317,N_1338,N_1290);
and U2318 (N_2318,N_1762,N_1450);
nor U2319 (N_2319,N_1247,N_1273);
and U2320 (N_2320,N_1483,N_1311);
and U2321 (N_2321,N_1407,N_1424);
nor U2322 (N_2322,N_1550,N_1397);
and U2323 (N_2323,N_1369,N_1689);
and U2324 (N_2324,N_1545,N_1577);
xnor U2325 (N_2325,N_1317,N_1665);
nand U2326 (N_2326,N_1522,N_1596);
nor U2327 (N_2327,N_1584,N_1421);
nor U2328 (N_2328,N_1693,N_1700);
and U2329 (N_2329,N_1472,N_1670);
nand U2330 (N_2330,N_1408,N_1633);
nor U2331 (N_2331,N_1645,N_1487);
nor U2332 (N_2332,N_1756,N_1680);
or U2333 (N_2333,N_1251,N_1572);
and U2334 (N_2334,N_1758,N_1636);
or U2335 (N_2335,N_1379,N_1519);
or U2336 (N_2336,N_1388,N_1406);
and U2337 (N_2337,N_1418,N_1516);
or U2338 (N_2338,N_1510,N_1294);
nand U2339 (N_2339,N_1395,N_1383);
nor U2340 (N_2340,N_1733,N_1226);
nor U2341 (N_2341,N_1365,N_1368);
xnor U2342 (N_2342,N_1767,N_1291);
and U2343 (N_2343,N_1601,N_1631);
nand U2344 (N_2344,N_1703,N_1567);
nor U2345 (N_2345,N_1739,N_1722);
xor U2346 (N_2346,N_1473,N_1566);
and U2347 (N_2347,N_1771,N_1753);
and U2348 (N_2348,N_1526,N_1452);
nor U2349 (N_2349,N_1393,N_1519);
or U2350 (N_2350,N_1763,N_1405);
and U2351 (N_2351,N_1767,N_1694);
nor U2352 (N_2352,N_1244,N_1585);
nand U2353 (N_2353,N_1785,N_1442);
or U2354 (N_2354,N_1287,N_1741);
or U2355 (N_2355,N_1561,N_1634);
nand U2356 (N_2356,N_1351,N_1689);
or U2357 (N_2357,N_1342,N_1394);
and U2358 (N_2358,N_1489,N_1490);
or U2359 (N_2359,N_1307,N_1672);
and U2360 (N_2360,N_1550,N_1640);
nor U2361 (N_2361,N_1226,N_1747);
nand U2362 (N_2362,N_1580,N_1565);
and U2363 (N_2363,N_1518,N_1726);
nand U2364 (N_2364,N_1498,N_1290);
xor U2365 (N_2365,N_1709,N_1760);
or U2366 (N_2366,N_1690,N_1524);
nand U2367 (N_2367,N_1509,N_1259);
and U2368 (N_2368,N_1532,N_1381);
or U2369 (N_2369,N_1796,N_1441);
and U2370 (N_2370,N_1593,N_1350);
and U2371 (N_2371,N_1238,N_1223);
and U2372 (N_2372,N_1526,N_1784);
nor U2373 (N_2373,N_1235,N_1792);
nand U2374 (N_2374,N_1309,N_1389);
and U2375 (N_2375,N_1735,N_1381);
nand U2376 (N_2376,N_1592,N_1769);
and U2377 (N_2377,N_1711,N_1494);
or U2378 (N_2378,N_1669,N_1637);
or U2379 (N_2379,N_1614,N_1601);
or U2380 (N_2380,N_1752,N_1618);
nor U2381 (N_2381,N_1253,N_1365);
or U2382 (N_2382,N_1460,N_1386);
or U2383 (N_2383,N_1693,N_1616);
nor U2384 (N_2384,N_1346,N_1235);
nand U2385 (N_2385,N_1498,N_1392);
nor U2386 (N_2386,N_1442,N_1383);
nand U2387 (N_2387,N_1752,N_1507);
nand U2388 (N_2388,N_1565,N_1295);
and U2389 (N_2389,N_1454,N_1645);
or U2390 (N_2390,N_1673,N_1245);
and U2391 (N_2391,N_1376,N_1777);
nand U2392 (N_2392,N_1764,N_1219);
nand U2393 (N_2393,N_1656,N_1466);
nor U2394 (N_2394,N_1428,N_1296);
and U2395 (N_2395,N_1429,N_1629);
or U2396 (N_2396,N_1372,N_1252);
nand U2397 (N_2397,N_1634,N_1573);
or U2398 (N_2398,N_1377,N_1535);
xnor U2399 (N_2399,N_1229,N_1203);
xor U2400 (N_2400,N_1830,N_2064);
nand U2401 (N_2401,N_2335,N_2360);
or U2402 (N_2402,N_2254,N_2015);
or U2403 (N_2403,N_2204,N_2091);
nor U2404 (N_2404,N_2189,N_2282);
and U2405 (N_2405,N_1988,N_1881);
or U2406 (N_2406,N_2201,N_2279);
nand U2407 (N_2407,N_2365,N_2343);
and U2408 (N_2408,N_2021,N_2376);
nand U2409 (N_2409,N_2303,N_2008);
nor U2410 (N_2410,N_2146,N_1816);
or U2411 (N_2411,N_2144,N_1879);
or U2412 (N_2412,N_2242,N_1936);
or U2413 (N_2413,N_2097,N_1899);
or U2414 (N_2414,N_2224,N_2155);
or U2415 (N_2415,N_1984,N_1974);
and U2416 (N_2416,N_1860,N_2167);
and U2417 (N_2417,N_1803,N_1958);
nand U2418 (N_2418,N_2194,N_1950);
xor U2419 (N_2419,N_2361,N_2026);
nor U2420 (N_2420,N_2076,N_1996);
nand U2421 (N_2421,N_2328,N_2103);
or U2422 (N_2422,N_1983,N_2207);
and U2423 (N_2423,N_1859,N_1935);
nand U2424 (N_2424,N_2186,N_2142);
or U2425 (N_2425,N_1800,N_2330);
and U2426 (N_2426,N_2038,N_2288);
nor U2427 (N_2427,N_2210,N_2390);
and U2428 (N_2428,N_1833,N_2357);
nor U2429 (N_2429,N_2251,N_2171);
and U2430 (N_2430,N_1865,N_2252);
nand U2431 (N_2431,N_2320,N_2147);
xnor U2432 (N_2432,N_2043,N_2280);
xor U2433 (N_2433,N_2087,N_2096);
and U2434 (N_2434,N_2264,N_2336);
or U2435 (N_2435,N_2339,N_1907);
nor U2436 (N_2436,N_1912,N_2305);
nor U2437 (N_2437,N_2317,N_2300);
nand U2438 (N_2438,N_1910,N_2296);
xnor U2439 (N_2439,N_2215,N_1973);
or U2440 (N_2440,N_2106,N_2101);
and U2441 (N_2441,N_2246,N_1904);
nand U2442 (N_2442,N_2222,N_2318);
and U2443 (N_2443,N_2377,N_2397);
nor U2444 (N_2444,N_1819,N_1848);
and U2445 (N_2445,N_1853,N_2132);
xor U2446 (N_2446,N_2019,N_1869);
or U2447 (N_2447,N_2355,N_2152);
and U2448 (N_2448,N_2177,N_2205);
or U2449 (N_2449,N_1971,N_1832);
xor U2450 (N_2450,N_1801,N_2187);
nand U2451 (N_2451,N_1908,N_1858);
and U2452 (N_2452,N_2190,N_1995);
and U2453 (N_2453,N_1970,N_2089);
or U2454 (N_2454,N_1977,N_2206);
or U2455 (N_2455,N_2078,N_1813);
nor U2456 (N_2456,N_2306,N_1931);
or U2457 (N_2457,N_2050,N_2071);
xnor U2458 (N_2458,N_2009,N_2133);
nor U2459 (N_2459,N_2113,N_2145);
nand U2460 (N_2460,N_2114,N_2183);
or U2461 (N_2461,N_2291,N_2260);
or U2462 (N_2462,N_2202,N_2245);
nand U2463 (N_2463,N_2240,N_1992);
xor U2464 (N_2464,N_1829,N_1896);
nand U2465 (N_2465,N_2011,N_2121);
or U2466 (N_2466,N_2104,N_2322);
nand U2467 (N_2467,N_1962,N_1986);
nand U2468 (N_2468,N_2110,N_1878);
and U2469 (N_2469,N_2380,N_2378);
nand U2470 (N_2470,N_2182,N_2369);
and U2471 (N_2471,N_1849,N_2333);
xnor U2472 (N_2472,N_1981,N_2017);
or U2473 (N_2473,N_2081,N_2090);
xnor U2474 (N_2474,N_1978,N_1929);
nor U2475 (N_2475,N_2031,N_2368);
nor U2476 (N_2476,N_2338,N_2345);
nor U2477 (N_2477,N_1985,N_2267);
and U2478 (N_2478,N_2085,N_1890);
xor U2479 (N_2479,N_2178,N_2116);
or U2480 (N_2480,N_2272,N_2310);
nor U2481 (N_2481,N_1989,N_2072);
and U2482 (N_2482,N_1847,N_1812);
and U2483 (N_2483,N_1918,N_2118);
or U2484 (N_2484,N_2088,N_2023);
or U2485 (N_2485,N_1941,N_1954);
nand U2486 (N_2486,N_2065,N_2018);
and U2487 (N_2487,N_2354,N_2217);
nor U2488 (N_2488,N_2150,N_2080);
or U2489 (N_2489,N_2311,N_1979);
nand U2490 (N_2490,N_1825,N_2068);
nand U2491 (N_2491,N_2014,N_1898);
nand U2492 (N_2492,N_2093,N_2002);
or U2493 (N_2493,N_2062,N_1874);
and U2494 (N_2494,N_2129,N_2055);
and U2495 (N_2495,N_2346,N_1972);
nor U2496 (N_2496,N_2108,N_2006);
nor U2497 (N_2497,N_2332,N_1964);
and U2498 (N_2498,N_2229,N_2243);
nor U2499 (N_2499,N_1876,N_2176);
nor U2500 (N_2500,N_2079,N_2384);
and U2501 (N_2501,N_1947,N_1976);
nand U2502 (N_2502,N_2281,N_1834);
and U2503 (N_2503,N_2148,N_2124);
and U2504 (N_2504,N_2226,N_1915);
nand U2505 (N_2505,N_1822,N_2203);
and U2506 (N_2506,N_1946,N_1917);
nor U2507 (N_2507,N_2301,N_1961);
or U2508 (N_2508,N_2166,N_1938);
nor U2509 (N_2509,N_2175,N_1945);
nor U2510 (N_2510,N_2347,N_2052);
xor U2511 (N_2511,N_2373,N_2241);
nor U2512 (N_2512,N_2070,N_2214);
nor U2513 (N_2513,N_1914,N_1885);
nand U2514 (N_2514,N_2083,N_2063);
nor U2515 (N_2515,N_2061,N_2163);
or U2516 (N_2516,N_2351,N_1880);
xnor U2517 (N_2517,N_2004,N_2169);
nor U2518 (N_2518,N_2250,N_2273);
nor U2519 (N_2519,N_2294,N_2162);
nand U2520 (N_2520,N_1863,N_1894);
nor U2521 (N_2521,N_2197,N_2331);
and U2522 (N_2522,N_2234,N_1957);
or U2523 (N_2523,N_1844,N_2256);
xnor U2524 (N_2524,N_2225,N_2387);
or U2525 (N_2525,N_2125,N_2290);
nand U2526 (N_2526,N_2247,N_2117);
or U2527 (N_2527,N_1944,N_1905);
nor U2528 (N_2528,N_2033,N_2266);
nor U2529 (N_2529,N_2352,N_2341);
nand U2530 (N_2530,N_1921,N_1870);
nand U2531 (N_2531,N_1919,N_2131);
nand U2532 (N_2532,N_2134,N_2275);
or U2533 (N_2533,N_2048,N_2016);
nor U2534 (N_2534,N_1851,N_2151);
or U2535 (N_2535,N_2058,N_2153);
xnor U2536 (N_2536,N_1839,N_1933);
nand U2537 (N_2537,N_2040,N_1953);
or U2538 (N_2538,N_1866,N_1968);
nand U2539 (N_2539,N_2136,N_2027);
or U2540 (N_2540,N_2237,N_2299);
nand U2541 (N_2541,N_1903,N_1815);
or U2542 (N_2542,N_1930,N_2158);
or U2543 (N_2543,N_2156,N_2356);
and U2544 (N_2544,N_2265,N_1835);
and U2545 (N_2545,N_2379,N_1808);
nand U2546 (N_2546,N_1951,N_2286);
and U2547 (N_2547,N_2385,N_2054);
nand U2548 (N_2548,N_2003,N_2382);
nor U2549 (N_2549,N_2223,N_2013);
or U2550 (N_2550,N_2284,N_2321);
nor U2551 (N_2551,N_2139,N_2208);
xor U2552 (N_2552,N_2297,N_2375);
and U2553 (N_2553,N_2200,N_2302);
xor U2554 (N_2554,N_2025,N_2034);
or U2555 (N_2555,N_1886,N_2329);
xnor U2556 (N_2556,N_2107,N_2323);
or U2557 (N_2557,N_2277,N_1883);
nand U2558 (N_2558,N_1991,N_2137);
and U2559 (N_2559,N_2135,N_2358);
xnor U2560 (N_2560,N_2057,N_2289);
nand U2561 (N_2561,N_1932,N_2227);
or U2562 (N_2562,N_2024,N_2391);
xnor U2563 (N_2563,N_2313,N_2395);
xnor U2564 (N_2564,N_2193,N_2037);
and U2565 (N_2565,N_2199,N_2164);
xor U2566 (N_2566,N_2235,N_2278);
nand U2567 (N_2567,N_2389,N_2255);
nand U2568 (N_2568,N_2244,N_2367);
xnor U2569 (N_2569,N_2337,N_1854);
and U2570 (N_2570,N_1982,N_2334);
nand U2571 (N_2571,N_1891,N_1949);
and U2572 (N_2572,N_1925,N_2128);
and U2573 (N_2573,N_2039,N_2001);
or U2574 (N_2574,N_1850,N_2069);
and U2575 (N_2575,N_2271,N_2213);
and U2576 (N_2576,N_1804,N_1924);
nor U2577 (N_2577,N_2261,N_2073);
and U2578 (N_2578,N_1864,N_2074);
or U2579 (N_2579,N_2325,N_2269);
nand U2580 (N_2580,N_2010,N_2092);
nand U2581 (N_2581,N_1913,N_1852);
or U2582 (N_2582,N_1955,N_1952);
and U2583 (N_2583,N_2042,N_1873);
or U2584 (N_2584,N_2120,N_2059);
nand U2585 (N_2585,N_1809,N_2130);
nand U2586 (N_2586,N_2123,N_1855);
xnor U2587 (N_2587,N_1960,N_1810);
and U2588 (N_2588,N_1838,N_1916);
nand U2589 (N_2589,N_2398,N_1998);
and U2590 (N_2590,N_2259,N_2172);
or U2591 (N_2591,N_2324,N_2319);
nor U2592 (N_2592,N_1841,N_2198);
and U2593 (N_2593,N_2100,N_1887);
and U2594 (N_2594,N_1993,N_1943);
xnor U2595 (N_2595,N_2022,N_2253);
or U2596 (N_2596,N_2184,N_1821);
xor U2597 (N_2597,N_1867,N_1966);
xnor U2598 (N_2598,N_2180,N_2230);
and U2599 (N_2599,N_1857,N_1871);
and U2600 (N_2600,N_2188,N_1897);
nand U2601 (N_2601,N_2170,N_1927);
or U2602 (N_2602,N_2049,N_2105);
nand U2603 (N_2603,N_2374,N_2221);
nand U2604 (N_2604,N_2231,N_1828);
nand U2605 (N_2605,N_2095,N_1846);
or U2606 (N_2606,N_2349,N_2007);
nor U2607 (N_2607,N_1902,N_2053);
nand U2608 (N_2608,N_2233,N_2179);
and U2609 (N_2609,N_2394,N_2044);
xnor U2610 (N_2610,N_2258,N_1840);
and U2611 (N_2611,N_2056,N_2066);
nand U2612 (N_2612,N_1826,N_1948);
xnor U2613 (N_2613,N_2283,N_2191);
nand U2614 (N_2614,N_2115,N_2030);
nor U2615 (N_2615,N_2216,N_1882);
nand U2616 (N_2616,N_1817,N_1922);
and U2617 (N_2617,N_2036,N_2327);
xnor U2618 (N_2618,N_2126,N_1911);
nand U2619 (N_2619,N_2268,N_1893);
and U2620 (N_2620,N_2000,N_2046);
or U2621 (N_2621,N_2276,N_2168);
and U2622 (N_2622,N_2220,N_2262);
xnor U2623 (N_2623,N_1926,N_2141);
or U2624 (N_2624,N_1956,N_1934);
or U2625 (N_2625,N_1843,N_1802);
xnor U2626 (N_2626,N_2084,N_2154);
and U2627 (N_2627,N_2035,N_2287);
or U2628 (N_2628,N_2098,N_1999);
nand U2629 (N_2629,N_2238,N_2209);
nor U2630 (N_2630,N_2393,N_2370);
or U2631 (N_2631,N_1997,N_2316);
or U2632 (N_2632,N_2047,N_2344);
and U2633 (N_2633,N_1831,N_2138);
nor U2634 (N_2634,N_2236,N_2359);
and U2635 (N_2635,N_1856,N_2249);
or U2636 (N_2636,N_1965,N_2051);
and U2637 (N_2637,N_1940,N_1845);
nor U2638 (N_2638,N_2399,N_2174);
or U2639 (N_2639,N_2274,N_1823);
xor U2640 (N_2640,N_2307,N_1811);
and U2641 (N_2641,N_2012,N_2396);
nand U2642 (N_2642,N_2232,N_2181);
and U2643 (N_2643,N_2032,N_2228);
and U2644 (N_2644,N_2159,N_2315);
nor U2645 (N_2645,N_2075,N_2298);
or U2646 (N_2646,N_1836,N_2348);
and U2647 (N_2647,N_1862,N_2160);
nand U2648 (N_2648,N_2340,N_2028);
nand U2649 (N_2649,N_2364,N_1975);
or U2650 (N_2650,N_1889,N_2263);
and U2651 (N_2651,N_2308,N_2041);
nor U2652 (N_2652,N_2099,N_1827);
nand U2653 (N_2653,N_1877,N_2143);
or U2654 (N_2654,N_2102,N_2342);
and U2655 (N_2655,N_2392,N_2212);
nand U2656 (N_2656,N_2218,N_2388);
and U2657 (N_2657,N_1980,N_2293);
or U2658 (N_2658,N_1824,N_2295);
nand U2659 (N_2659,N_2020,N_2173);
and U2660 (N_2660,N_1814,N_1900);
and U2661 (N_2661,N_1990,N_2045);
nor U2662 (N_2662,N_1805,N_1942);
or U2663 (N_2663,N_2326,N_2309);
and U2664 (N_2664,N_1868,N_2140);
nand U2665 (N_2665,N_2292,N_1806);
nor U2666 (N_2666,N_2067,N_2270);
nand U2667 (N_2667,N_2157,N_2077);
or U2668 (N_2668,N_2372,N_2304);
nand U2669 (N_2669,N_1837,N_2086);
or U2670 (N_2670,N_2127,N_2112);
and U2671 (N_2671,N_1928,N_1959);
and U2672 (N_2672,N_2239,N_2285);
nor U2673 (N_2673,N_1872,N_1861);
and U2674 (N_2674,N_1895,N_2111);
or U2675 (N_2675,N_1937,N_1807);
xnor U2676 (N_2676,N_2257,N_2353);
or U2677 (N_2677,N_2196,N_2366);
and U2678 (N_2678,N_1994,N_2094);
xor U2679 (N_2679,N_2383,N_1875);
and U2680 (N_2680,N_2219,N_1967);
or U2681 (N_2681,N_2161,N_2192);
nand U2682 (N_2682,N_2362,N_2314);
xnor U2683 (N_2683,N_1923,N_2386);
nand U2684 (N_2684,N_2165,N_2119);
nand U2685 (N_2685,N_1888,N_1820);
nand U2686 (N_2686,N_2371,N_1987);
nor U2687 (N_2687,N_2005,N_2211);
or U2688 (N_2688,N_1939,N_1963);
and U2689 (N_2689,N_2185,N_1901);
or U2690 (N_2690,N_1884,N_1842);
or U2691 (N_2691,N_2248,N_1969);
and U2692 (N_2692,N_2029,N_1818);
and U2693 (N_2693,N_1906,N_2082);
or U2694 (N_2694,N_1920,N_2122);
or U2695 (N_2695,N_2109,N_2149);
nand U2696 (N_2696,N_2363,N_1909);
nor U2697 (N_2697,N_2060,N_2381);
nand U2698 (N_2698,N_2350,N_2195);
or U2699 (N_2699,N_1892,N_2312);
or U2700 (N_2700,N_1997,N_2177);
and U2701 (N_2701,N_1960,N_2172);
nor U2702 (N_2702,N_2109,N_2267);
xor U2703 (N_2703,N_2084,N_2333);
and U2704 (N_2704,N_2160,N_2020);
nor U2705 (N_2705,N_2305,N_2029);
nand U2706 (N_2706,N_2243,N_2347);
nor U2707 (N_2707,N_1997,N_2181);
and U2708 (N_2708,N_2041,N_1831);
nand U2709 (N_2709,N_1939,N_2165);
nand U2710 (N_2710,N_1858,N_2128);
and U2711 (N_2711,N_2042,N_2169);
or U2712 (N_2712,N_2199,N_1838);
xnor U2713 (N_2713,N_2106,N_2331);
nor U2714 (N_2714,N_1881,N_1814);
xnor U2715 (N_2715,N_1824,N_2030);
nand U2716 (N_2716,N_2330,N_2086);
and U2717 (N_2717,N_2205,N_1888);
nor U2718 (N_2718,N_2365,N_1813);
or U2719 (N_2719,N_1990,N_1819);
or U2720 (N_2720,N_2042,N_2055);
nor U2721 (N_2721,N_2361,N_2003);
xnor U2722 (N_2722,N_1976,N_1808);
nand U2723 (N_2723,N_2111,N_2287);
or U2724 (N_2724,N_2207,N_2050);
or U2725 (N_2725,N_2084,N_2041);
or U2726 (N_2726,N_2195,N_1835);
nor U2727 (N_2727,N_1988,N_1894);
nand U2728 (N_2728,N_2104,N_2258);
nor U2729 (N_2729,N_1913,N_2352);
and U2730 (N_2730,N_2240,N_2362);
xnor U2731 (N_2731,N_2172,N_2008);
and U2732 (N_2732,N_1907,N_2345);
and U2733 (N_2733,N_2046,N_2114);
and U2734 (N_2734,N_1913,N_2014);
nand U2735 (N_2735,N_2091,N_2325);
xnor U2736 (N_2736,N_1941,N_1819);
and U2737 (N_2737,N_1916,N_2331);
and U2738 (N_2738,N_2294,N_2065);
nor U2739 (N_2739,N_1829,N_2122);
or U2740 (N_2740,N_2236,N_2227);
and U2741 (N_2741,N_1942,N_2370);
or U2742 (N_2742,N_2083,N_2395);
nor U2743 (N_2743,N_2227,N_2081);
and U2744 (N_2744,N_2167,N_1951);
and U2745 (N_2745,N_2229,N_2319);
nand U2746 (N_2746,N_2070,N_2298);
or U2747 (N_2747,N_2256,N_2266);
xor U2748 (N_2748,N_2000,N_1838);
or U2749 (N_2749,N_1843,N_2282);
nand U2750 (N_2750,N_2266,N_1918);
and U2751 (N_2751,N_1960,N_2277);
nor U2752 (N_2752,N_2354,N_1866);
or U2753 (N_2753,N_2263,N_1870);
and U2754 (N_2754,N_1829,N_2226);
nand U2755 (N_2755,N_1980,N_2286);
xor U2756 (N_2756,N_2300,N_1848);
nand U2757 (N_2757,N_1953,N_2074);
nand U2758 (N_2758,N_2118,N_2167);
or U2759 (N_2759,N_2212,N_1898);
and U2760 (N_2760,N_2017,N_1865);
nand U2761 (N_2761,N_1826,N_2372);
nor U2762 (N_2762,N_1857,N_2121);
nand U2763 (N_2763,N_2359,N_1916);
or U2764 (N_2764,N_1844,N_2219);
or U2765 (N_2765,N_2332,N_1855);
nand U2766 (N_2766,N_1916,N_2297);
nor U2767 (N_2767,N_1823,N_1886);
and U2768 (N_2768,N_2365,N_2369);
nand U2769 (N_2769,N_2359,N_2309);
or U2770 (N_2770,N_2160,N_2261);
nand U2771 (N_2771,N_2254,N_2073);
or U2772 (N_2772,N_2271,N_1944);
nor U2773 (N_2773,N_2219,N_1811);
nor U2774 (N_2774,N_1887,N_1878);
and U2775 (N_2775,N_2192,N_2087);
nand U2776 (N_2776,N_2044,N_2362);
and U2777 (N_2777,N_2268,N_2161);
or U2778 (N_2778,N_2361,N_1857);
or U2779 (N_2779,N_1810,N_2053);
nand U2780 (N_2780,N_1897,N_2184);
nand U2781 (N_2781,N_2046,N_2123);
or U2782 (N_2782,N_2333,N_2224);
or U2783 (N_2783,N_1909,N_2374);
or U2784 (N_2784,N_1989,N_2298);
nand U2785 (N_2785,N_1929,N_2151);
or U2786 (N_2786,N_1841,N_2257);
and U2787 (N_2787,N_1974,N_1808);
xor U2788 (N_2788,N_2284,N_2006);
and U2789 (N_2789,N_2178,N_2235);
or U2790 (N_2790,N_2044,N_1924);
nor U2791 (N_2791,N_2162,N_2114);
xnor U2792 (N_2792,N_2114,N_2385);
xnor U2793 (N_2793,N_2151,N_1980);
nand U2794 (N_2794,N_1913,N_2037);
and U2795 (N_2795,N_2090,N_1989);
or U2796 (N_2796,N_2121,N_1842);
or U2797 (N_2797,N_1847,N_2133);
nand U2798 (N_2798,N_2386,N_2271);
or U2799 (N_2799,N_2350,N_2139);
nand U2800 (N_2800,N_1856,N_1803);
nand U2801 (N_2801,N_1897,N_2174);
and U2802 (N_2802,N_2279,N_2189);
and U2803 (N_2803,N_1882,N_2317);
nand U2804 (N_2804,N_2055,N_2238);
nor U2805 (N_2805,N_2277,N_1812);
and U2806 (N_2806,N_2224,N_2149);
nand U2807 (N_2807,N_1889,N_1868);
nand U2808 (N_2808,N_2303,N_1974);
xor U2809 (N_2809,N_2103,N_2096);
nor U2810 (N_2810,N_1905,N_2239);
or U2811 (N_2811,N_2257,N_2159);
and U2812 (N_2812,N_2374,N_2375);
nand U2813 (N_2813,N_1904,N_1837);
or U2814 (N_2814,N_2140,N_1996);
nand U2815 (N_2815,N_1932,N_2331);
nand U2816 (N_2816,N_1972,N_2252);
nor U2817 (N_2817,N_2292,N_2327);
and U2818 (N_2818,N_2369,N_2248);
and U2819 (N_2819,N_2109,N_1983);
nand U2820 (N_2820,N_1853,N_2099);
nor U2821 (N_2821,N_1954,N_2115);
xor U2822 (N_2822,N_1911,N_2173);
nand U2823 (N_2823,N_2318,N_2065);
nand U2824 (N_2824,N_1927,N_2265);
or U2825 (N_2825,N_2344,N_2150);
nand U2826 (N_2826,N_2175,N_1868);
nor U2827 (N_2827,N_2052,N_2094);
nor U2828 (N_2828,N_2370,N_2176);
nor U2829 (N_2829,N_1943,N_1879);
nand U2830 (N_2830,N_1893,N_2219);
nand U2831 (N_2831,N_2265,N_1952);
or U2832 (N_2832,N_2098,N_2133);
nand U2833 (N_2833,N_2256,N_1880);
nor U2834 (N_2834,N_2030,N_1928);
or U2835 (N_2835,N_2058,N_1944);
and U2836 (N_2836,N_2078,N_2386);
nor U2837 (N_2837,N_1954,N_2138);
nor U2838 (N_2838,N_1837,N_2223);
xnor U2839 (N_2839,N_2252,N_1930);
or U2840 (N_2840,N_2351,N_2348);
or U2841 (N_2841,N_1990,N_2120);
and U2842 (N_2842,N_1831,N_2351);
and U2843 (N_2843,N_2000,N_1997);
nand U2844 (N_2844,N_2293,N_1957);
xnor U2845 (N_2845,N_2176,N_1858);
or U2846 (N_2846,N_2381,N_2206);
nor U2847 (N_2847,N_1971,N_2249);
nor U2848 (N_2848,N_2294,N_2309);
nor U2849 (N_2849,N_2391,N_1838);
or U2850 (N_2850,N_2339,N_2318);
nor U2851 (N_2851,N_1887,N_2196);
nor U2852 (N_2852,N_2091,N_2005);
xor U2853 (N_2853,N_2377,N_1895);
nor U2854 (N_2854,N_2074,N_2060);
nand U2855 (N_2855,N_2366,N_1832);
and U2856 (N_2856,N_2300,N_2210);
or U2857 (N_2857,N_2147,N_2228);
nand U2858 (N_2858,N_2168,N_2073);
nand U2859 (N_2859,N_2306,N_1870);
and U2860 (N_2860,N_1873,N_2166);
xor U2861 (N_2861,N_1911,N_1895);
and U2862 (N_2862,N_2359,N_1887);
xor U2863 (N_2863,N_1915,N_2062);
nor U2864 (N_2864,N_2161,N_2341);
and U2865 (N_2865,N_1988,N_2239);
or U2866 (N_2866,N_1945,N_2346);
nand U2867 (N_2867,N_1822,N_1999);
nor U2868 (N_2868,N_2126,N_1807);
or U2869 (N_2869,N_2321,N_2208);
and U2870 (N_2870,N_1921,N_2116);
nor U2871 (N_2871,N_2228,N_1979);
and U2872 (N_2872,N_2109,N_2363);
nand U2873 (N_2873,N_2333,N_1819);
xor U2874 (N_2874,N_2210,N_1836);
or U2875 (N_2875,N_1816,N_2055);
nor U2876 (N_2876,N_1919,N_1841);
nand U2877 (N_2877,N_1919,N_2379);
nand U2878 (N_2878,N_2070,N_2073);
nor U2879 (N_2879,N_2297,N_2262);
and U2880 (N_2880,N_2226,N_2014);
or U2881 (N_2881,N_2028,N_1893);
or U2882 (N_2882,N_1862,N_1878);
nand U2883 (N_2883,N_1857,N_2099);
nor U2884 (N_2884,N_2180,N_2243);
or U2885 (N_2885,N_2282,N_2292);
nand U2886 (N_2886,N_1976,N_2371);
or U2887 (N_2887,N_2264,N_2369);
xnor U2888 (N_2888,N_2147,N_1869);
nor U2889 (N_2889,N_1993,N_2129);
nand U2890 (N_2890,N_1999,N_1927);
and U2891 (N_2891,N_1989,N_2371);
and U2892 (N_2892,N_2174,N_1882);
nand U2893 (N_2893,N_2165,N_2162);
nand U2894 (N_2894,N_2330,N_1814);
xnor U2895 (N_2895,N_1878,N_1957);
nor U2896 (N_2896,N_2157,N_1841);
nand U2897 (N_2897,N_2235,N_2289);
nand U2898 (N_2898,N_2097,N_2376);
nand U2899 (N_2899,N_1822,N_1832);
nor U2900 (N_2900,N_1906,N_1837);
or U2901 (N_2901,N_2300,N_2185);
and U2902 (N_2902,N_2309,N_1897);
nor U2903 (N_2903,N_2197,N_2344);
nand U2904 (N_2904,N_2286,N_1937);
xor U2905 (N_2905,N_1862,N_1884);
nor U2906 (N_2906,N_2117,N_1961);
nand U2907 (N_2907,N_2333,N_1899);
nand U2908 (N_2908,N_2370,N_2360);
and U2909 (N_2909,N_2229,N_2367);
xnor U2910 (N_2910,N_1990,N_2275);
xnor U2911 (N_2911,N_1881,N_1979);
nor U2912 (N_2912,N_2355,N_1937);
nor U2913 (N_2913,N_2335,N_2230);
nand U2914 (N_2914,N_2279,N_2153);
or U2915 (N_2915,N_2179,N_2074);
nand U2916 (N_2916,N_2287,N_2327);
or U2917 (N_2917,N_2173,N_1925);
nand U2918 (N_2918,N_2162,N_1933);
nand U2919 (N_2919,N_1860,N_2283);
nand U2920 (N_2920,N_2367,N_1964);
and U2921 (N_2921,N_1926,N_1807);
nand U2922 (N_2922,N_2222,N_2331);
nor U2923 (N_2923,N_2210,N_2204);
nor U2924 (N_2924,N_2019,N_2374);
or U2925 (N_2925,N_2330,N_2310);
and U2926 (N_2926,N_1822,N_2128);
xnor U2927 (N_2927,N_2119,N_1991);
nand U2928 (N_2928,N_2189,N_2024);
or U2929 (N_2929,N_1961,N_2147);
nor U2930 (N_2930,N_1817,N_1854);
nand U2931 (N_2931,N_1818,N_1904);
and U2932 (N_2932,N_2043,N_1998);
nand U2933 (N_2933,N_1821,N_1820);
or U2934 (N_2934,N_1809,N_1850);
nor U2935 (N_2935,N_2317,N_1849);
and U2936 (N_2936,N_2369,N_1950);
xnor U2937 (N_2937,N_2076,N_2033);
or U2938 (N_2938,N_2192,N_2046);
nand U2939 (N_2939,N_2095,N_2133);
nand U2940 (N_2940,N_2249,N_1822);
and U2941 (N_2941,N_2045,N_1825);
nand U2942 (N_2942,N_2064,N_1829);
nor U2943 (N_2943,N_2133,N_2158);
or U2944 (N_2944,N_2307,N_2355);
nand U2945 (N_2945,N_2005,N_2137);
and U2946 (N_2946,N_1861,N_1963);
xor U2947 (N_2947,N_1897,N_2227);
or U2948 (N_2948,N_1863,N_2242);
or U2949 (N_2949,N_2287,N_2043);
nand U2950 (N_2950,N_2140,N_1943);
nand U2951 (N_2951,N_2267,N_2376);
and U2952 (N_2952,N_1945,N_2213);
xnor U2953 (N_2953,N_1847,N_2065);
xor U2954 (N_2954,N_2280,N_2206);
or U2955 (N_2955,N_2288,N_2030);
or U2956 (N_2956,N_1874,N_2151);
nand U2957 (N_2957,N_2123,N_1992);
xor U2958 (N_2958,N_2311,N_2284);
and U2959 (N_2959,N_2389,N_2060);
nor U2960 (N_2960,N_1989,N_2323);
nand U2961 (N_2961,N_1898,N_2073);
nand U2962 (N_2962,N_1960,N_2134);
nand U2963 (N_2963,N_2202,N_2210);
or U2964 (N_2964,N_1907,N_2200);
or U2965 (N_2965,N_2184,N_2349);
nand U2966 (N_2966,N_2382,N_2179);
or U2967 (N_2967,N_1829,N_2386);
or U2968 (N_2968,N_1975,N_2190);
nor U2969 (N_2969,N_2178,N_2390);
nor U2970 (N_2970,N_2363,N_2252);
nor U2971 (N_2971,N_1946,N_2342);
or U2972 (N_2972,N_2169,N_2267);
nand U2973 (N_2973,N_2195,N_2102);
or U2974 (N_2974,N_2365,N_2394);
or U2975 (N_2975,N_2363,N_1980);
nand U2976 (N_2976,N_2039,N_2087);
or U2977 (N_2977,N_1963,N_1899);
or U2978 (N_2978,N_2281,N_2184);
nor U2979 (N_2979,N_1873,N_1985);
nor U2980 (N_2980,N_2254,N_2076);
xnor U2981 (N_2981,N_2355,N_2021);
nand U2982 (N_2982,N_2163,N_2139);
or U2983 (N_2983,N_2328,N_2108);
xnor U2984 (N_2984,N_1899,N_1891);
nand U2985 (N_2985,N_2299,N_1827);
and U2986 (N_2986,N_2350,N_1982);
xnor U2987 (N_2987,N_2273,N_2048);
or U2988 (N_2988,N_2062,N_2026);
or U2989 (N_2989,N_2229,N_1912);
nand U2990 (N_2990,N_2348,N_2036);
and U2991 (N_2991,N_1894,N_2365);
and U2992 (N_2992,N_1974,N_2158);
nand U2993 (N_2993,N_2294,N_1925);
nor U2994 (N_2994,N_2354,N_2009);
nand U2995 (N_2995,N_1956,N_2203);
and U2996 (N_2996,N_2043,N_2332);
and U2997 (N_2997,N_2250,N_2207);
nor U2998 (N_2998,N_2166,N_2387);
nand U2999 (N_2999,N_2101,N_2070);
and UO_0 (O_0,N_2782,N_2600);
or UO_1 (O_1,N_2781,N_2750);
or UO_2 (O_2,N_2854,N_2928);
xnor UO_3 (O_3,N_2649,N_2429);
nand UO_4 (O_4,N_2604,N_2775);
and UO_5 (O_5,N_2506,N_2425);
nand UO_6 (O_6,N_2763,N_2831);
nand UO_7 (O_7,N_2903,N_2812);
and UO_8 (O_8,N_2733,N_2578);
nand UO_9 (O_9,N_2704,N_2647);
and UO_10 (O_10,N_2746,N_2911);
xor UO_11 (O_11,N_2769,N_2748);
nand UO_12 (O_12,N_2939,N_2512);
or UO_13 (O_13,N_2980,N_2660);
and UO_14 (O_14,N_2848,N_2642);
nand UO_15 (O_15,N_2721,N_2910);
and UO_16 (O_16,N_2764,N_2666);
nand UO_17 (O_17,N_2577,N_2557);
nand UO_18 (O_18,N_2713,N_2899);
nor UO_19 (O_19,N_2561,N_2665);
nand UO_20 (O_20,N_2779,N_2460);
nor UO_21 (O_21,N_2857,N_2446);
and UO_22 (O_22,N_2679,N_2644);
or UO_23 (O_23,N_2596,N_2908);
nor UO_24 (O_24,N_2491,N_2637);
xor UO_25 (O_25,N_2450,N_2587);
nor UO_26 (O_26,N_2970,N_2631);
xnor UO_27 (O_27,N_2459,N_2437);
nor UO_28 (O_28,N_2796,N_2951);
or UO_29 (O_29,N_2950,N_2994);
and UO_30 (O_30,N_2946,N_2845);
nand UO_31 (O_31,N_2440,N_2747);
nand UO_32 (O_32,N_2580,N_2475);
nor UO_33 (O_33,N_2619,N_2919);
or UO_34 (O_34,N_2987,N_2489);
and UO_35 (O_35,N_2926,N_2916);
nand UO_36 (O_36,N_2653,N_2548);
and UO_37 (O_37,N_2873,N_2902);
nand UO_38 (O_38,N_2481,N_2958);
or UO_39 (O_39,N_2607,N_2757);
nand UO_40 (O_40,N_2530,N_2828);
or UO_41 (O_41,N_2770,N_2790);
and UO_42 (O_42,N_2671,N_2598);
nor UO_43 (O_43,N_2431,N_2803);
nor UO_44 (O_44,N_2420,N_2662);
nand UO_45 (O_45,N_2694,N_2984);
xor UO_46 (O_46,N_2710,N_2714);
nor UO_47 (O_47,N_2591,N_2936);
nand UO_48 (O_48,N_2488,N_2773);
or UO_49 (O_49,N_2435,N_2887);
xnor UO_50 (O_50,N_2687,N_2859);
and UO_51 (O_51,N_2808,N_2461);
nand UO_52 (O_52,N_2620,N_2403);
xor UO_53 (O_53,N_2675,N_2676);
nor UO_54 (O_54,N_2798,N_2978);
nor UO_55 (O_55,N_2406,N_2814);
and UO_56 (O_56,N_2641,N_2877);
nand UO_57 (O_57,N_2650,N_2457);
nor UO_58 (O_58,N_2633,N_2517);
and UO_59 (O_59,N_2989,N_2652);
or UO_60 (O_60,N_2473,N_2667);
nor UO_61 (O_61,N_2851,N_2906);
and UO_62 (O_62,N_2556,N_2863);
nand UO_63 (O_63,N_2504,N_2444);
and UO_64 (O_64,N_2449,N_2678);
or UO_65 (O_65,N_2510,N_2788);
nor UO_66 (O_66,N_2588,N_2719);
nor UO_67 (O_67,N_2836,N_2921);
and UO_68 (O_68,N_2526,N_2971);
nor UO_69 (O_69,N_2696,N_2811);
nor UO_70 (O_70,N_2819,N_2762);
or UO_71 (O_71,N_2981,N_2786);
and UO_72 (O_72,N_2486,N_2949);
nand UO_73 (O_73,N_2847,N_2458);
nand UO_74 (O_74,N_2944,N_2551);
nand UO_75 (O_75,N_2515,N_2691);
nand UO_76 (O_76,N_2521,N_2611);
or UO_77 (O_77,N_2527,N_2505);
or UO_78 (O_78,N_2472,N_2904);
nand UO_79 (O_79,N_2776,N_2953);
and UO_80 (O_80,N_2760,N_2617);
nor UO_81 (O_81,N_2560,N_2869);
nand UO_82 (O_82,N_2858,N_2448);
and UO_83 (O_83,N_2736,N_2988);
and UO_84 (O_84,N_2738,N_2948);
and UO_85 (O_85,N_2905,N_2842);
or UO_86 (O_86,N_2495,N_2659);
and UO_87 (O_87,N_2616,N_2998);
xor UO_88 (O_88,N_2547,N_2925);
or UO_89 (O_89,N_2780,N_2586);
xor UO_90 (O_90,N_2484,N_2592);
or UO_91 (O_91,N_2966,N_2913);
nor UO_92 (O_92,N_2840,N_2663);
and UO_93 (O_93,N_2879,N_2728);
xor UO_94 (O_94,N_2418,N_2477);
nor UO_95 (O_95,N_2933,N_2590);
and UO_96 (O_96,N_2542,N_2401);
or UO_97 (O_97,N_2576,N_2929);
nand UO_98 (O_98,N_2492,N_2534);
nor UO_99 (O_99,N_2683,N_2741);
or UO_100 (O_100,N_2638,N_2745);
nor UO_101 (O_101,N_2499,N_2882);
or UO_102 (O_102,N_2997,N_2940);
and UO_103 (O_103,N_2668,N_2648);
nand UO_104 (O_104,N_2955,N_2606);
and UO_105 (O_105,N_2729,N_2414);
nor UO_106 (O_106,N_2430,N_2661);
and UO_107 (O_107,N_2947,N_2417);
and UO_108 (O_108,N_2574,N_2570);
nand UO_109 (O_109,N_2875,N_2427);
nand UO_110 (O_110,N_2523,N_2471);
nand UO_111 (O_111,N_2680,N_2522);
or UO_112 (O_112,N_2669,N_2538);
or UO_113 (O_113,N_2800,N_2846);
or UO_114 (O_114,N_2563,N_2892);
or UO_115 (O_115,N_2476,N_2685);
nor UO_116 (O_116,N_2901,N_2708);
nor UO_117 (O_117,N_2500,N_2442);
nand UO_118 (O_118,N_2945,N_2732);
or UO_119 (O_119,N_2474,N_2829);
or UO_120 (O_120,N_2555,N_2549);
and UO_121 (O_121,N_2465,N_2802);
and UO_122 (O_122,N_2447,N_2524);
nand UO_123 (O_123,N_2428,N_2817);
and UO_124 (O_124,N_2843,N_2826);
nand UO_125 (O_125,N_2888,N_2751);
nand UO_126 (O_126,N_2756,N_2954);
nand UO_127 (O_127,N_2525,N_2885);
and UO_128 (O_128,N_2466,N_2795);
nand UO_129 (O_129,N_2407,N_2601);
xnor UO_130 (O_130,N_2503,N_2967);
nand UO_131 (O_131,N_2573,N_2402);
nand UO_132 (O_132,N_2868,N_2880);
and UO_133 (O_133,N_2884,N_2824);
or UO_134 (O_134,N_2799,N_2602);
nor UO_135 (O_135,N_2743,N_2640);
xnor UO_136 (O_136,N_2507,N_2864);
nand UO_137 (O_137,N_2546,N_2677);
or UO_138 (O_138,N_2927,N_2924);
and UO_139 (O_139,N_2720,N_2623);
or UO_140 (O_140,N_2479,N_2918);
or UO_141 (O_141,N_2722,N_2657);
and UO_142 (O_142,N_2862,N_2917);
or UO_143 (O_143,N_2451,N_2774);
nand UO_144 (O_144,N_2711,N_2454);
or UO_145 (O_145,N_2920,N_2895);
or UO_146 (O_146,N_2942,N_2636);
xnor UO_147 (O_147,N_2768,N_2584);
nand UO_148 (O_148,N_2866,N_2965);
or UO_149 (O_149,N_2532,N_2567);
and UO_150 (O_150,N_2702,N_2493);
nor UO_151 (O_151,N_2533,N_2935);
and UO_152 (O_152,N_2896,N_2835);
nor UO_153 (O_153,N_2583,N_2608);
nand UO_154 (O_154,N_2934,N_2985);
nand UO_155 (O_155,N_2634,N_2603);
nand UO_156 (O_156,N_2558,N_2566);
and UO_157 (O_157,N_2673,N_2830);
xor UO_158 (O_158,N_2618,N_2959);
nor UO_159 (O_159,N_2497,N_2412);
nand UO_160 (O_160,N_2872,N_2635);
nor UO_161 (O_161,N_2871,N_2737);
and UO_162 (O_162,N_2718,N_2571);
nand UO_163 (O_163,N_2852,N_2791);
or UO_164 (O_164,N_2700,N_2441);
and UO_165 (O_165,N_2595,N_2974);
or UO_166 (O_166,N_2681,N_2655);
xnor UO_167 (O_167,N_2498,N_2968);
and UO_168 (O_168,N_2597,N_2502);
nand UO_169 (O_169,N_2400,N_2575);
nor UO_170 (O_170,N_2629,N_2849);
nor UO_171 (O_171,N_2627,N_2893);
nor UO_172 (O_172,N_2579,N_2443);
and UO_173 (O_173,N_2801,N_2883);
or UO_174 (O_174,N_2931,N_2861);
or UO_175 (O_175,N_2421,N_2535);
nand UO_176 (O_176,N_2982,N_2469);
nor UO_177 (O_177,N_2979,N_2490);
or UO_178 (O_178,N_2529,N_2496);
or UO_179 (O_179,N_2411,N_2544);
nand UO_180 (O_180,N_2766,N_2463);
and UO_181 (O_181,N_2912,N_2664);
or UO_182 (O_182,N_2559,N_2754);
nand UO_183 (O_183,N_2881,N_2740);
nand UO_184 (O_184,N_2907,N_2509);
nor UO_185 (O_185,N_2876,N_2424);
nor UO_186 (O_186,N_2712,N_2519);
nand UO_187 (O_187,N_2996,N_2483);
or UO_188 (O_188,N_2975,N_2550);
or UO_189 (O_189,N_2821,N_2716);
or UO_190 (O_190,N_2426,N_2992);
nor UO_191 (O_191,N_2436,N_2531);
nand UO_192 (O_192,N_2438,N_2794);
nor UO_193 (O_193,N_2727,N_2609);
nand UO_194 (O_194,N_2964,N_2915);
nor UO_195 (O_195,N_2569,N_2993);
or UO_196 (O_196,N_2930,N_2742);
nand UO_197 (O_197,N_2581,N_2651);
nor UO_198 (O_198,N_2894,N_2914);
or UO_199 (O_199,N_2878,N_2839);
and UO_200 (O_200,N_2445,N_2815);
or UO_201 (O_201,N_2672,N_2784);
and UO_202 (O_202,N_2832,N_2897);
or UO_203 (O_203,N_2698,N_2957);
and UO_204 (O_204,N_2494,N_2889);
nor UO_205 (O_205,N_2804,N_2825);
xnor UO_206 (O_206,N_2639,N_2536);
and UO_207 (O_207,N_2612,N_2765);
nand UO_208 (O_208,N_2961,N_2886);
and UO_209 (O_209,N_2744,N_2416);
or UO_210 (O_210,N_2909,N_2991);
nand UO_211 (O_211,N_2514,N_2962);
nor UO_212 (O_212,N_2995,N_2543);
or UO_213 (O_213,N_2805,N_2455);
or UO_214 (O_214,N_2787,N_2865);
nand UO_215 (O_215,N_2844,N_2874);
or UO_216 (O_216,N_2856,N_2983);
or UO_217 (O_217,N_2772,N_2833);
and UO_218 (O_218,N_2943,N_2564);
xor UO_219 (O_219,N_2462,N_2761);
and UO_220 (O_220,N_2759,N_2478);
xor UO_221 (O_221,N_2562,N_2624);
nand UO_222 (O_222,N_2464,N_2870);
nor UO_223 (O_223,N_2599,N_2690);
or UO_224 (O_224,N_2482,N_2467);
nor UO_225 (O_225,N_2860,N_2572);
and UO_226 (O_226,N_2956,N_2963);
nor UO_227 (O_227,N_2777,N_2705);
nand UO_228 (O_228,N_2553,N_2969);
and UO_229 (O_229,N_2485,N_2793);
and UO_230 (O_230,N_2841,N_2941);
nand UO_231 (O_231,N_2594,N_2452);
nor UO_232 (O_232,N_2810,N_2990);
and UO_233 (O_233,N_2890,N_2709);
and UO_234 (O_234,N_2755,N_2837);
xor UO_235 (O_235,N_2827,N_2752);
or UO_236 (O_236,N_2726,N_2434);
or UO_237 (O_237,N_2568,N_2818);
xor UO_238 (O_238,N_2855,N_2646);
and UO_239 (O_239,N_2783,N_2614);
or UO_240 (O_240,N_2697,N_2986);
and UO_241 (O_241,N_2834,N_2593);
nand UO_242 (O_242,N_2735,N_2731);
xor UO_243 (O_243,N_2541,N_2518);
xor UO_244 (O_244,N_2701,N_2749);
and UO_245 (O_245,N_2820,N_2923);
and UO_246 (O_246,N_2898,N_2415);
and UO_247 (O_247,N_2409,N_2853);
nand UO_248 (O_248,N_2695,N_2707);
nor UO_249 (O_249,N_2423,N_2508);
nor UO_250 (O_250,N_2891,N_2552);
nor UO_251 (O_251,N_2582,N_2610);
nor UO_252 (O_252,N_2900,N_2758);
nand UO_253 (O_253,N_2806,N_2689);
or UO_254 (O_254,N_2626,N_2630);
and UO_255 (O_255,N_2932,N_2973);
nand UO_256 (O_256,N_2778,N_2554);
or UO_257 (O_257,N_2516,N_2405);
nor UO_258 (O_258,N_2976,N_2838);
xnor UO_259 (O_259,N_2537,N_2520);
xnor UO_260 (O_260,N_2809,N_2404);
or UO_261 (O_261,N_2419,N_2613);
nor UO_262 (O_262,N_2410,N_2674);
or UO_263 (O_263,N_2480,N_2682);
nor UO_264 (O_264,N_2977,N_2692);
xnor UO_265 (O_265,N_2703,N_2730);
and UO_266 (O_266,N_2565,N_2622);
xnor UO_267 (O_267,N_2456,N_2734);
nand UO_268 (O_268,N_2539,N_2433);
or UO_269 (O_269,N_2725,N_2408);
nor UO_270 (O_270,N_2501,N_2670);
nor UO_271 (O_271,N_2823,N_2589);
or UO_272 (O_272,N_2686,N_2816);
xor UO_273 (O_273,N_2487,N_2422);
nand UO_274 (O_274,N_2797,N_2771);
or UO_275 (O_275,N_2615,N_2922);
and UO_276 (O_276,N_2850,N_2767);
nor UO_277 (O_277,N_2605,N_2684);
and UO_278 (O_278,N_2432,N_2792);
nand UO_279 (O_279,N_2723,N_2688);
nand UO_280 (O_280,N_2470,N_2789);
xnor UO_281 (O_281,N_2513,N_2658);
or UO_282 (O_282,N_2867,N_2511);
nand UO_283 (O_283,N_2717,N_2625);
nor UO_284 (O_284,N_2952,N_2545);
nand UO_285 (O_285,N_2706,N_2413);
xor UO_286 (O_286,N_2528,N_2739);
nor UO_287 (O_287,N_2938,N_2645);
nand UO_288 (O_288,N_2628,N_2822);
and UO_289 (O_289,N_2972,N_2960);
xnor UO_290 (O_290,N_2785,N_2937);
or UO_291 (O_291,N_2715,N_2632);
and UO_292 (O_292,N_2999,N_2753);
or UO_293 (O_293,N_2724,N_2540);
and UO_294 (O_294,N_2621,N_2656);
and UO_295 (O_295,N_2439,N_2699);
or UO_296 (O_296,N_2807,N_2453);
and UO_297 (O_297,N_2693,N_2643);
nor UO_298 (O_298,N_2813,N_2468);
nand UO_299 (O_299,N_2585,N_2654);
or UO_300 (O_300,N_2987,N_2957);
xnor UO_301 (O_301,N_2449,N_2698);
nand UO_302 (O_302,N_2497,N_2466);
xnor UO_303 (O_303,N_2618,N_2642);
nor UO_304 (O_304,N_2951,N_2742);
and UO_305 (O_305,N_2740,N_2832);
or UO_306 (O_306,N_2613,N_2563);
nor UO_307 (O_307,N_2632,N_2975);
nor UO_308 (O_308,N_2990,N_2779);
or UO_309 (O_309,N_2688,N_2888);
or UO_310 (O_310,N_2831,N_2969);
nor UO_311 (O_311,N_2771,N_2744);
nor UO_312 (O_312,N_2717,N_2629);
nor UO_313 (O_313,N_2408,N_2811);
nand UO_314 (O_314,N_2681,N_2679);
and UO_315 (O_315,N_2638,N_2839);
nand UO_316 (O_316,N_2928,N_2817);
and UO_317 (O_317,N_2479,N_2797);
nor UO_318 (O_318,N_2566,N_2526);
nor UO_319 (O_319,N_2841,N_2575);
nor UO_320 (O_320,N_2493,N_2797);
and UO_321 (O_321,N_2842,N_2654);
xor UO_322 (O_322,N_2984,N_2709);
nand UO_323 (O_323,N_2886,N_2773);
or UO_324 (O_324,N_2978,N_2945);
nand UO_325 (O_325,N_2725,N_2799);
nor UO_326 (O_326,N_2442,N_2626);
or UO_327 (O_327,N_2737,N_2806);
nor UO_328 (O_328,N_2960,N_2434);
nand UO_329 (O_329,N_2631,N_2587);
or UO_330 (O_330,N_2413,N_2952);
nor UO_331 (O_331,N_2879,N_2701);
nor UO_332 (O_332,N_2519,N_2442);
or UO_333 (O_333,N_2855,N_2786);
nand UO_334 (O_334,N_2570,N_2901);
or UO_335 (O_335,N_2424,N_2735);
or UO_336 (O_336,N_2900,N_2880);
nand UO_337 (O_337,N_2490,N_2996);
nand UO_338 (O_338,N_2838,N_2411);
nor UO_339 (O_339,N_2858,N_2842);
and UO_340 (O_340,N_2813,N_2455);
nand UO_341 (O_341,N_2533,N_2961);
nor UO_342 (O_342,N_2781,N_2597);
and UO_343 (O_343,N_2967,N_2701);
nor UO_344 (O_344,N_2495,N_2812);
or UO_345 (O_345,N_2617,N_2555);
or UO_346 (O_346,N_2894,N_2674);
nor UO_347 (O_347,N_2426,N_2958);
nand UO_348 (O_348,N_2626,N_2418);
nor UO_349 (O_349,N_2752,N_2864);
xor UO_350 (O_350,N_2695,N_2820);
nand UO_351 (O_351,N_2489,N_2647);
nand UO_352 (O_352,N_2451,N_2464);
nor UO_353 (O_353,N_2659,N_2718);
nor UO_354 (O_354,N_2616,N_2555);
and UO_355 (O_355,N_2696,N_2458);
nand UO_356 (O_356,N_2516,N_2634);
nand UO_357 (O_357,N_2868,N_2581);
nand UO_358 (O_358,N_2666,N_2550);
nand UO_359 (O_359,N_2524,N_2463);
nand UO_360 (O_360,N_2970,N_2892);
and UO_361 (O_361,N_2611,N_2951);
and UO_362 (O_362,N_2784,N_2442);
nand UO_363 (O_363,N_2939,N_2714);
and UO_364 (O_364,N_2860,N_2650);
nand UO_365 (O_365,N_2804,N_2614);
and UO_366 (O_366,N_2792,N_2756);
nor UO_367 (O_367,N_2672,N_2970);
or UO_368 (O_368,N_2660,N_2443);
or UO_369 (O_369,N_2904,N_2829);
nand UO_370 (O_370,N_2518,N_2964);
nor UO_371 (O_371,N_2784,N_2774);
nand UO_372 (O_372,N_2941,N_2695);
and UO_373 (O_373,N_2642,N_2639);
and UO_374 (O_374,N_2908,N_2604);
and UO_375 (O_375,N_2779,N_2780);
and UO_376 (O_376,N_2675,N_2485);
nand UO_377 (O_377,N_2608,N_2919);
or UO_378 (O_378,N_2752,N_2740);
nor UO_379 (O_379,N_2731,N_2416);
or UO_380 (O_380,N_2838,N_2569);
or UO_381 (O_381,N_2517,N_2686);
nand UO_382 (O_382,N_2944,N_2799);
xnor UO_383 (O_383,N_2493,N_2849);
nand UO_384 (O_384,N_2679,N_2555);
xnor UO_385 (O_385,N_2651,N_2704);
nor UO_386 (O_386,N_2461,N_2930);
nand UO_387 (O_387,N_2887,N_2818);
nor UO_388 (O_388,N_2920,N_2523);
or UO_389 (O_389,N_2803,N_2611);
nand UO_390 (O_390,N_2526,N_2968);
or UO_391 (O_391,N_2774,N_2940);
nor UO_392 (O_392,N_2824,N_2563);
nor UO_393 (O_393,N_2421,N_2496);
nor UO_394 (O_394,N_2622,N_2433);
xor UO_395 (O_395,N_2718,N_2726);
and UO_396 (O_396,N_2755,N_2489);
and UO_397 (O_397,N_2464,N_2982);
and UO_398 (O_398,N_2406,N_2869);
or UO_399 (O_399,N_2912,N_2895);
and UO_400 (O_400,N_2891,N_2862);
nor UO_401 (O_401,N_2762,N_2803);
or UO_402 (O_402,N_2851,N_2862);
and UO_403 (O_403,N_2588,N_2669);
nand UO_404 (O_404,N_2585,N_2421);
and UO_405 (O_405,N_2578,N_2619);
xnor UO_406 (O_406,N_2458,N_2467);
and UO_407 (O_407,N_2940,N_2832);
and UO_408 (O_408,N_2900,N_2415);
nand UO_409 (O_409,N_2712,N_2617);
and UO_410 (O_410,N_2954,N_2832);
and UO_411 (O_411,N_2483,N_2920);
and UO_412 (O_412,N_2736,N_2858);
and UO_413 (O_413,N_2885,N_2828);
or UO_414 (O_414,N_2577,N_2490);
and UO_415 (O_415,N_2716,N_2525);
nand UO_416 (O_416,N_2574,N_2670);
nor UO_417 (O_417,N_2450,N_2942);
nand UO_418 (O_418,N_2572,N_2779);
or UO_419 (O_419,N_2893,N_2496);
xnor UO_420 (O_420,N_2665,N_2582);
nand UO_421 (O_421,N_2875,N_2661);
or UO_422 (O_422,N_2542,N_2446);
and UO_423 (O_423,N_2956,N_2453);
or UO_424 (O_424,N_2435,N_2616);
nand UO_425 (O_425,N_2493,N_2855);
and UO_426 (O_426,N_2774,N_2473);
nand UO_427 (O_427,N_2805,N_2984);
nor UO_428 (O_428,N_2522,N_2645);
and UO_429 (O_429,N_2491,N_2517);
nor UO_430 (O_430,N_2509,N_2755);
nor UO_431 (O_431,N_2777,N_2937);
nor UO_432 (O_432,N_2400,N_2817);
or UO_433 (O_433,N_2959,N_2987);
and UO_434 (O_434,N_2483,N_2761);
or UO_435 (O_435,N_2599,N_2834);
and UO_436 (O_436,N_2896,N_2560);
and UO_437 (O_437,N_2607,N_2775);
or UO_438 (O_438,N_2488,N_2497);
nand UO_439 (O_439,N_2879,N_2410);
nor UO_440 (O_440,N_2830,N_2534);
xor UO_441 (O_441,N_2884,N_2512);
and UO_442 (O_442,N_2623,N_2933);
nor UO_443 (O_443,N_2901,N_2752);
nand UO_444 (O_444,N_2553,N_2646);
or UO_445 (O_445,N_2629,N_2704);
nand UO_446 (O_446,N_2604,N_2887);
or UO_447 (O_447,N_2691,N_2850);
nand UO_448 (O_448,N_2427,N_2929);
or UO_449 (O_449,N_2815,N_2535);
and UO_450 (O_450,N_2825,N_2872);
nor UO_451 (O_451,N_2816,N_2990);
nor UO_452 (O_452,N_2880,N_2455);
xnor UO_453 (O_453,N_2942,N_2772);
nand UO_454 (O_454,N_2518,N_2423);
and UO_455 (O_455,N_2467,N_2965);
nand UO_456 (O_456,N_2589,N_2637);
and UO_457 (O_457,N_2563,N_2483);
nand UO_458 (O_458,N_2757,N_2865);
nand UO_459 (O_459,N_2474,N_2604);
or UO_460 (O_460,N_2699,N_2414);
nor UO_461 (O_461,N_2976,N_2743);
and UO_462 (O_462,N_2774,N_2492);
nand UO_463 (O_463,N_2799,N_2982);
or UO_464 (O_464,N_2625,N_2758);
nor UO_465 (O_465,N_2998,N_2933);
or UO_466 (O_466,N_2574,N_2697);
and UO_467 (O_467,N_2680,N_2977);
nor UO_468 (O_468,N_2585,N_2556);
xor UO_469 (O_469,N_2898,N_2518);
xnor UO_470 (O_470,N_2406,N_2610);
nor UO_471 (O_471,N_2446,N_2716);
nand UO_472 (O_472,N_2579,N_2437);
nand UO_473 (O_473,N_2439,N_2937);
nor UO_474 (O_474,N_2818,N_2722);
nand UO_475 (O_475,N_2717,N_2573);
nor UO_476 (O_476,N_2554,N_2713);
nand UO_477 (O_477,N_2677,N_2429);
nand UO_478 (O_478,N_2664,N_2429);
nand UO_479 (O_479,N_2507,N_2993);
or UO_480 (O_480,N_2862,N_2837);
or UO_481 (O_481,N_2475,N_2495);
nor UO_482 (O_482,N_2459,N_2879);
or UO_483 (O_483,N_2778,N_2501);
nor UO_484 (O_484,N_2419,N_2709);
and UO_485 (O_485,N_2648,N_2526);
or UO_486 (O_486,N_2822,N_2641);
xnor UO_487 (O_487,N_2867,N_2966);
or UO_488 (O_488,N_2433,N_2541);
xnor UO_489 (O_489,N_2538,N_2744);
or UO_490 (O_490,N_2763,N_2651);
nor UO_491 (O_491,N_2820,N_2968);
nor UO_492 (O_492,N_2629,N_2839);
xnor UO_493 (O_493,N_2841,N_2473);
nor UO_494 (O_494,N_2721,N_2404);
and UO_495 (O_495,N_2889,N_2720);
or UO_496 (O_496,N_2578,N_2966);
nand UO_497 (O_497,N_2586,N_2736);
nor UO_498 (O_498,N_2842,N_2981);
or UO_499 (O_499,N_2444,N_2965);
endmodule