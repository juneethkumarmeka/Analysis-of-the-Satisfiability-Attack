module basic_500_3000_500_30_levels_1xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_178,In_294);
or U1 (N_1,In_118,In_466);
nand U2 (N_2,In_91,In_205);
nand U3 (N_3,In_170,In_399);
and U4 (N_4,In_227,In_461);
or U5 (N_5,In_62,In_113);
nand U6 (N_6,In_224,In_330);
xor U7 (N_7,In_131,In_163);
nor U8 (N_8,In_384,In_428);
nor U9 (N_9,In_332,In_460);
nand U10 (N_10,In_183,In_284);
and U11 (N_11,In_124,In_499);
nand U12 (N_12,In_390,In_265);
or U13 (N_13,In_42,In_420);
and U14 (N_14,In_348,In_448);
or U15 (N_15,In_387,In_79);
and U16 (N_16,In_156,In_223);
nand U17 (N_17,In_167,In_446);
or U18 (N_18,In_68,In_482);
or U19 (N_19,In_288,In_371);
nor U20 (N_20,In_232,In_280);
nor U21 (N_21,In_145,In_203);
nor U22 (N_22,In_447,In_380);
nor U23 (N_23,In_308,In_12);
nand U24 (N_24,In_416,In_405);
and U25 (N_25,In_483,In_152);
nand U26 (N_26,In_426,In_339);
nor U27 (N_27,In_353,In_144);
nor U28 (N_28,In_396,In_327);
and U29 (N_29,In_52,In_293);
or U30 (N_30,In_86,In_143);
nor U31 (N_31,In_326,In_22);
and U32 (N_32,In_202,In_324);
or U33 (N_33,In_136,In_291);
and U34 (N_34,In_204,In_242);
nor U35 (N_35,In_254,In_243);
nand U36 (N_36,In_261,In_239);
nor U37 (N_37,In_322,In_382);
and U38 (N_38,In_320,In_153);
nand U39 (N_39,In_166,In_188);
or U40 (N_40,In_126,In_328);
and U41 (N_41,In_316,In_108);
nand U42 (N_42,In_484,In_295);
nand U43 (N_43,In_128,In_32);
or U44 (N_44,In_356,In_212);
and U45 (N_45,In_302,In_146);
nor U46 (N_46,In_459,In_278);
or U47 (N_47,In_38,In_341);
nand U48 (N_48,In_120,In_207);
and U49 (N_49,In_400,In_255);
and U50 (N_50,In_444,In_47);
or U51 (N_51,In_0,In_83);
or U52 (N_52,In_347,In_401);
nor U53 (N_53,In_192,In_365);
nor U54 (N_54,In_301,In_364);
nor U55 (N_55,In_236,In_479);
or U56 (N_56,In_422,In_84);
nand U57 (N_57,In_336,In_383);
or U58 (N_58,In_221,In_149);
and U59 (N_59,In_252,In_321);
or U60 (N_60,In_100,In_55);
and U61 (N_61,In_475,In_343);
and U62 (N_62,In_160,In_7);
or U63 (N_63,In_44,In_107);
or U64 (N_64,In_187,In_64);
or U65 (N_65,In_306,In_395);
nand U66 (N_66,In_6,In_331);
or U67 (N_67,In_51,In_218);
nand U68 (N_68,In_480,In_161);
or U69 (N_69,In_196,In_311);
nand U70 (N_70,In_184,In_436);
and U71 (N_71,In_61,In_282);
nand U72 (N_72,In_424,In_168);
nor U73 (N_73,In_429,In_344);
nor U74 (N_74,In_78,In_262);
or U75 (N_75,In_60,In_419);
or U76 (N_76,In_148,In_123);
nor U77 (N_77,In_50,In_18);
nor U78 (N_78,In_271,In_494);
nand U79 (N_79,In_93,In_171);
or U80 (N_80,In_317,In_299);
and U81 (N_81,In_125,In_25);
nor U82 (N_82,In_251,In_67);
nor U83 (N_83,In_24,In_338);
or U84 (N_84,In_437,In_442);
and U85 (N_85,In_443,In_240);
nand U86 (N_86,In_391,In_497);
or U87 (N_87,In_337,In_250);
and U88 (N_88,In_76,In_403);
or U89 (N_89,In_496,In_245);
or U90 (N_90,In_394,In_409);
nor U91 (N_91,In_69,In_412);
nand U92 (N_92,In_189,In_342);
nand U93 (N_93,In_57,In_375);
or U94 (N_94,In_290,In_367);
or U95 (N_95,In_427,In_346);
and U96 (N_96,In_440,In_111);
or U97 (N_97,In_402,In_358);
nand U98 (N_98,In_104,In_173);
nor U99 (N_99,In_267,In_374);
or U100 (N_100,In_457,In_281);
nand U101 (N_101,N_57,In_389);
or U102 (N_102,In_169,In_112);
nor U103 (N_103,In_435,In_49);
nand U104 (N_104,In_87,In_210);
nor U105 (N_105,N_32,In_28);
and U106 (N_106,In_360,In_115);
nor U107 (N_107,In_16,In_458);
or U108 (N_108,In_272,In_410);
nor U109 (N_109,In_190,In_398);
nor U110 (N_110,In_490,N_91);
nor U111 (N_111,In_425,In_200);
or U112 (N_112,In_355,In_119);
nand U113 (N_113,In_370,In_439);
nor U114 (N_114,N_59,In_135);
or U115 (N_115,In_368,In_88);
or U116 (N_116,In_415,In_63);
or U117 (N_117,N_58,In_154);
or U118 (N_118,In_27,In_274);
and U119 (N_119,In_477,In_372);
or U120 (N_120,N_25,In_433);
or U121 (N_121,N_82,In_40);
nand U122 (N_122,In_441,N_99);
nand U123 (N_123,N_98,In_417);
or U124 (N_124,In_13,In_90);
and U125 (N_125,In_231,In_286);
nor U126 (N_126,In_388,In_366);
or U127 (N_127,N_45,In_8);
nor U128 (N_128,In_77,In_462);
and U129 (N_129,N_92,In_305);
nand U130 (N_130,N_83,In_455);
nand U131 (N_131,In_33,In_48);
nor U132 (N_132,In_397,In_452);
and U133 (N_133,In_71,In_406);
nand U134 (N_134,In_206,N_16);
nand U135 (N_135,In_471,N_27);
and U136 (N_136,N_60,In_465);
nand U137 (N_137,N_70,In_139);
nand U138 (N_138,In_445,In_127);
nand U139 (N_139,N_11,In_414);
or U140 (N_140,N_67,In_185);
and U141 (N_141,N_35,N_81);
or U142 (N_142,N_75,In_379);
nand U143 (N_143,In_2,In_195);
nand U144 (N_144,In_359,In_408);
nor U145 (N_145,N_29,N_78);
or U146 (N_146,N_65,In_138);
nor U147 (N_147,In_208,N_97);
xnor U148 (N_148,N_6,In_101);
and U149 (N_149,In_14,In_489);
or U150 (N_150,In_323,In_109);
or U151 (N_151,In_335,In_85);
and U152 (N_152,N_76,N_49);
nand U153 (N_153,N_13,In_418);
or U154 (N_154,In_438,In_247);
or U155 (N_155,In_421,N_40);
nand U156 (N_156,In_319,In_46);
or U157 (N_157,In_469,In_373);
nand U158 (N_158,N_55,In_182);
or U159 (N_159,N_10,N_61);
and U160 (N_160,In_3,In_266);
and U161 (N_161,In_197,In_386);
nor U162 (N_162,N_63,In_357);
or U163 (N_163,In_31,N_14);
nor U164 (N_164,In_157,N_39);
nand U165 (N_165,N_7,N_12);
nor U166 (N_166,In_180,In_162);
and U167 (N_167,In_9,N_3);
nand U168 (N_168,In_434,In_130);
nand U169 (N_169,In_315,In_493);
nor U170 (N_170,In_292,In_256);
or U171 (N_171,In_492,In_34);
or U172 (N_172,In_26,In_334);
and U173 (N_173,In_222,N_62);
and U174 (N_174,In_423,N_77);
nor U175 (N_175,In_307,In_450);
and U176 (N_176,In_354,In_474);
or U177 (N_177,In_270,In_333);
nor U178 (N_178,In_211,In_468);
and U179 (N_179,In_404,In_228);
nor U180 (N_180,N_15,In_385);
and U181 (N_181,In_296,In_5);
nor U182 (N_182,In_476,N_74);
nor U183 (N_183,In_98,In_491);
nor U184 (N_184,In_407,In_129);
or U185 (N_185,In_392,N_71);
or U186 (N_186,In_4,In_45);
nor U187 (N_187,In_248,In_467);
nand U188 (N_188,In_472,N_0);
or U189 (N_189,N_88,In_485);
nand U190 (N_190,In_159,In_142);
or U191 (N_191,In_209,In_17);
or U192 (N_192,N_66,In_220);
nand U193 (N_193,N_42,N_87);
or U194 (N_194,N_22,In_451);
nor U195 (N_195,In_151,In_313);
and U196 (N_196,In_147,In_310);
nand U197 (N_197,In_340,N_50);
nor U198 (N_198,N_56,In_463);
or U199 (N_199,N_64,In_249);
nor U200 (N_200,N_151,N_107);
nand U201 (N_201,N_195,N_101);
nor U202 (N_202,N_47,In_81);
nand U203 (N_203,In_226,In_214);
nand U204 (N_204,In_275,In_241);
or U205 (N_205,N_147,N_20);
nor U206 (N_206,In_300,N_102);
nor U207 (N_207,In_20,N_181);
nor U208 (N_208,N_152,N_44);
or U209 (N_209,N_93,N_133);
and U210 (N_210,In_453,N_119);
and U211 (N_211,In_285,In_158);
nor U212 (N_212,N_145,In_133);
or U213 (N_213,In_481,N_121);
and U214 (N_214,N_54,In_54);
nor U215 (N_215,N_117,N_68);
and U216 (N_216,N_69,N_53);
nand U217 (N_217,In_141,In_89);
and U218 (N_218,In_413,N_183);
and U219 (N_219,In_96,N_85);
nand U220 (N_220,In_268,In_376);
and U221 (N_221,N_192,In_225);
nor U222 (N_222,In_478,N_72);
and U223 (N_223,In_276,In_174);
nor U224 (N_224,N_124,N_189);
nor U225 (N_225,N_161,In_488);
nand U226 (N_226,In_229,In_53);
or U227 (N_227,In_116,In_191);
nand U228 (N_228,N_100,N_33);
nand U229 (N_229,In_431,N_19);
or U230 (N_230,In_351,N_21);
or U231 (N_231,In_260,In_97);
nor U232 (N_232,N_95,In_36);
or U233 (N_233,N_163,In_257);
and U234 (N_234,In_110,In_94);
nor U235 (N_235,In_105,In_495);
nor U236 (N_236,In_273,N_169);
xor U237 (N_237,N_120,N_174);
or U238 (N_238,In_41,N_24);
nor U239 (N_239,In_114,In_219);
nor U240 (N_240,N_166,N_18);
nor U241 (N_241,In_198,In_325);
or U242 (N_242,N_106,In_70);
or U243 (N_243,N_94,N_104);
xor U244 (N_244,In_329,N_164);
nor U245 (N_245,In_92,N_197);
and U246 (N_246,In_473,In_362);
or U247 (N_247,In_264,N_118);
nand U248 (N_248,N_132,In_432);
and U249 (N_249,N_80,N_185);
nor U250 (N_250,N_129,In_186);
and U251 (N_251,N_148,In_121);
nand U252 (N_252,N_4,N_138);
and U253 (N_253,N_115,In_361);
nand U254 (N_254,N_79,In_309);
nand U255 (N_255,N_48,In_244);
and U256 (N_256,N_1,N_108);
nor U257 (N_257,In_289,In_263);
nand U258 (N_258,In_363,N_116);
nor U259 (N_259,N_127,In_132);
nor U260 (N_260,N_126,N_157);
or U261 (N_261,In_74,N_179);
nor U262 (N_262,In_75,In_140);
nand U263 (N_263,N_143,N_187);
nand U264 (N_264,In_381,N_162);
nor U265 (N_265,N_139,In_314);
and U266 (N_266,In_176,N_160);
and U267 (N_267,N_175,N_178);
nand U268 (N_268,In_377,N_158);
nand U269 (N_269,In_106,In_283);
and U270 (N_270,N_90,N_26);
nand U271 (N_271,N_86,In_175);
and U272 (N_272,In_82,N_41);
nor U273 (N_273,N_122,N_8);
and U274 (N_274,In_318,N_51);
nor U275 (N_275,N_173,N_111);
nand U276 (N_276,In_1,In_454);
or U277 (N_277,In_258,N_96);
nand U278 (N_278,N_168,N_105);
and U279 (N_279,N_171,In_179);
nand U280 (N_280,In_411,In_352);
nor U281 (N_281,N_130,N_114);
nor U282 (N_282,N_5,N_184);
nand U283 (N_283,In_449,In_164);
or U284 (N_284,In_11,In_134);
and U285 (N_285,N_176,In_269);
nand U286 (N_286,N_34,In_369);
and U287 (N_287,N_199,N_146);
nor U288 (N_288,N_155,N_123);
and U289 (N_289,N_196,In_102);
and U290 (N_290,In_43,In_30);
nand U291 (N_291,N_37,In_35);
or U292 (N_292,N_194,In_230);
or U293 (N_293,N_31,N_113);
and U294 (N_294,N_177,N_134);
nand U295 (N_295,N_89,In_464);
or U296 (N_296,In_312,N_186);
and U297 (N_297,In_287,In_378);
or U298 (N_298,In_172,In_345);
or U299 (N_299,In_193,In_29);
nand U300 (N_300,N_30,In_470);
and U301 (N_301,In_253,N_142);
and U302 (N_302,N_28,N_255);
or U303 (N_303,N_264,N_140);
nor U304 (N_304,N_207,In_73);
and U305 (N_305,N_219,In_297);
and U306 (N_306,N_188,N_46);
and U307 (N_307,In_72,N_43);
nor U308 (N_308,N_223,N_249);
and U309 (N_309,N_243,N_9);
and U310 (N_310,N_235,N_182);
and U311 (N_311,N_131,N_227);
nand U312 (N_312,N_222,N_204);
and U313 (N_313,N_190,N_218);
nor U314 (N_314,N_274,N_293);
nand U315 (N_315,N_220,In_277);
and U316 (N_316,In_201,N_286);
nor U317 (N_317,N_180,In_137);
or U318 (N_318,N_292,N_137);
nand U319 (N_319,In_215,In_298);
nor U320 (N_320,N_170,In_117);
and U321 (N_321,In_350,In_217);
or U322 (N_322,In_37,N_232);
and U323 (N_323,N_203,In_122);
or U324 (N_324,N_271,N_165);
nand U325 (N_325,In_246,N_245);
and U326 (N_326,N_298,N_150);
nand U327 (N_327,N_250,N_193);
nand U328 (N_328,N_210,N_266);
xor U329 (N_329,In_213,In_103);
nor U330 (N_330,In_237,N_228);
nor U331 (N_331,N_144,N_237);
and U332 (N_332,N_23,N_284);
nor U333 (N_333,In_216,In_165);
nand U334 (N_334,In_80,N_263);
or U335 (N_335,N_136,N_229);
or U336 (N_336,N_2,N_234);
or U337 (N_337,In_21,N_153);
or U338 (N_338,N_225,N_231);
and U339 (N_339,N_252,N_224);
nand U340 (N_340,N_251,N_110);
nand U341 (N_341,N_200,In_15);
nor U342 (N_342,N_276,N_247);
and U343 (N_343,N_212,N_275);
nor U344 (N_344,N_279,N_260);
nand U345 (N_345,In_194,In_238);
or U346 (N_346,N_135,N_84);
nor U347 (N_347,In_155,N_270);
nor U348 (N_348,N_209,In_430);
and U349 (N_349,In_349,N_283);
or U350 (N_350,N_278,N_282);
nor U351 (N_351,N_273,N_267);
and U352 (N_352,In_56,In_235);
and U353 (N_353,N_253,N_254);
or U354 (N_354,N_299,N_290);
and U355 (N_355,N_198,N_259);
nand U356 (N_356,In_181,In_150);
or U357 (N_357,N_272,In_393);
and U358 (N_358,N_36,N_141);
and U359 (N_359,N_230,In_303);
or U360 (N_360,N_156,In_498);
and U361 (N_361,N_17,N_221);
nand U362 (N_362,N_191,N_201);
or U363 (N_363,N_206,In_58);
or U364 (N_364,N_52,N_296);
nand U365 (N_365,In_486,N_295);
and U366 (N_366,N_159,N_280);
nand U367 (N_367,In_23,N_242);
nand U368 (N_368,N_233,N_246);
nor U369 (N_369,N_73,N_213);
and U370 (N_370,N_277,N_294);
nand U371 (N_371,N_205,N_208);
nand U372 (N_372,N_103,N_239);
nand U373 (N_373,N_240,N_241);
nor U374 (N_374,In_487,N_214);
and U375 (N_375,N_202,N_211);
nand U376 (N_376,In_59,In_19);
or U377 (N_377,N_258,N_149);
and U378 (N_378,N_287,In_99);
nand U379 (N_379,In_66,N_167);
and U380 (N_380,N_257,In_259);
or U381 (N_381,N_268,N_109);
nor U382 (N_382,N_112,N_248);
or U383 (N_383,In_199,N_217);
nand U384 (N_384,N_269,In_10);
or U385 (N_385,N_262,In_65);
nor U386 (N_386,N_297,N_236);
nor U387 (N_387,N_281,In_39);
and U388 (N_388,In_304,N_125);
or U389 (N_389,N_285,N_172);
and U390 (N_390,N_256,N_288);
and U391 (N_391,In_177,N_128);
nor U392 (N_392,In_233,N_215);
nand U393 (N_393,N_238,In_456);
and U394 (N_394,N_216,N_38);
nand U395 (N_395,In_279,N_289);
and U396 (N_396,In_234,N_261);
or U397 (N_397,N_291,N_244);
and U398 (N_398,N_265,N_154);
nor U399 (N_399,In_95,N_226);
and U400 (N_400,N_382,N_388);
or U401 (N_401,N_379,N_303);
and U402 (N_402,N_333,N_347);
and U403 (N_403,N_348,N_366);
nor U404 (N_404,N_384,N_367);
or U405 (N_405,N_370,N_316);
xnor U406 (N_406,N_377,N_322);
nor U407 (N_407,N_374,N_319);
and U408 (N_408,N_396,N_317);
or U409 (N_409,N_386,N_355);
and U410 (N_410,N_380,N_314);
nand U411 (N_411,N_369,N_346);
xor U412 (N_412,N_358,N_323);
or U413 (N_413,N_357,N_328);
nand U414 (N_414,N_387,N_373);
or U415 (N_415,N_308,N_307);
nand U416 (N_416,N_344,N_397);
nor U417 (N_417,N_350,N_310);
or U418 (N_418,N_371,N_375);
and U419 (N_419,N_364,N_385);
and U420 (N_420,N_338,N_311);
nor U421 (N_421,N_334,N_312);
nand U422 (N_422,N_330,N_362);
and U423 (N_423,N_327,N_325);
nor U424 (N_424,N_341,N_340);
nor U425 (N_425,N_393,N_352);
nand U426 (N_426,N_343,N_372);
and U427 (N_427,N_398,N_339);
or U428 (N_428,N_365,N_376);
or U429 (N_429,N_313,N_345);
or U430 (N_430,N_399,N_302);
and U431 (N_431,N_394,N_315);
or U432 (N_432,N_342,N_349);
nor U433 (N_433,N_363,N_337);
or U434 (N_434,N_301,N_356);
nor U435 (N_435,N_368,N_395);
xor U436 (N_436,N_354,N_360);
nand U437 (N_437,N_351,N_335);
or U438 (N_438,N_300,N_331);
xor U439 (N_439,N_321,N_320);
or U440 (N_440,N_383,N_353);
or U441 (N_441,N_332,N_304);
nand U442 (N_442,N_391,N_392);
nand U443 (N_443,N_390,N_305);
or U444 (N_444,N_378,N_336);
or U445 (N_445,N_326,N_389);
or U446 (N_446,N_324,N_318);
or U447 (N_447,N_359,N_309);
and U448 (N_448,N_329,N_361);
nor U449 (N_449,N_381,N_306);
nor U450 (N_450,N_300,N_309);
and U451 (N_451,N_308,N_311);
nor U452 (N_452,N_375,N_316);
nand U453 (N_453,N_395,N_376);
or U454 (N_454,N_332,N_348);
nand U455 (N_455,N_359,N_381);
nand U456 (N_456,N_359,N_363);
xnor U457 (N_457,N_327,N_398);
and U458 (N_458,N_319,N_331);
nand U459 (N_459,N_396,N_300);
nor U460 (N_460,N_322,N_306);
or U461 (N_461,N_322,N_376);
nand U462 (N_462,N_352,N_313);
and U463 (N_463,N_315,N_390);
nand U464 (N_464,N_384,N_346);
and U465 (N_465,N_334,N_335);
or U466 (N_466,N_305,N_301);
nand U467 (N_467,N_367,N_372);
xor U468 (N_468,N_336,N_371);
nor U469 (N_469,N_353,N_354);
or U470 (N_470,N_323,N_306);
nor U471 (N_471,N_347,N_309);
or U472 (N_472,N_383,N_372);
nand U473 (N_473,N_343,N_347);
nor U474 (N_474,N_346,N_381);
or U475 (N_475,N_328,N_398);
nor U476 (N_476,N_358,N_388);
or U477 (N_477,N_308,N_328);
and U478 (N_478,N_324,N_327);
nand U479 (N_479,N_301,N_379);
nand U480 (N_480,N_301,N_321);
nand U481 (N_481,N_372,N_369);
nor U482 (N_482,N_320,N_375);
or U483 (N_483,N_382,N_380);
nand U484 (N_484,N_336,N_370);
nor U485 (N_485,N_388,N_355);
nand U486 (N_486,N_358,N_387);
nand U487 (N_487,N_399,N_318);
nor U488 (N_488,N_377,N_337);
or U489 (N_489,N_358,N_367);
nand U490 (N_490,N_313,N_315);
or U491 (N_491,N_396,N_328);
nor U492 (N_492,N_386,N_312);
nand U493 (N_493,N_343,N_356);
and U494 (N_494,N_382,N_307);
and U495 (N_495,N_329,N_372);
and U496 (N_496,N_357,N_310);
nand U497 (N_497,N_371,N_308);
and U498 (N_498,N_388,N_317);
or U499 (N_499,N_344,N_348);
and U500 (N_500,N_484,N_441);
and U501 (N_501,N_477,N_492);
nor U502 (N_502,N_478,N_480);
nor U503 (N_503,N_467,N_428);
nor U504 (N_504,N_449,N_499);
nand U505 (N_505,N_405,N_498);
or U506 (N_506,N_496,N_485);
or U507 (N_507,N_490,N_414);
and U508 (N_508,N_447,N_440);
nor U509 (N_509,N_439,N_483);
nand U510 (N_510,N_495,N_486);
or U511 (N_511,N_443,N_413);
nand U512 (N_512,N_476,N_472);
nor U513 (N_513,N_434,N_451);
nor U514 (N_514,N_426,N_453);
or U515 (N_515,N_409,N_415);
nand U516 (N_516,N_444,N_423);
nand U517 (N_517,N_475,N_402);
nand U518 (N_518,N_456,N_494);
nor U519 (N_519,N_470,N_446);
nand U520 (N_520,N_433,N_429);
xor U521 (N_521,N_408,N_436);
nand U522 (N_522,N_421,N_400);
and U523 (N_523,N_407,N_489);
and U524 (N_524,N_454,N_469);
and U525 (N_525,N_458,N_459);
xnor U526 (N_526,N_497,N_487);
nor U527 (N_527,N_493,N_471);
or U528 (N_528,N_435,N_452);
nor U529 (N_529,N_468,N_406);
nand U530 (N_530,N_438,N_430);
nor U531 (N_531,N_466,N_411);
nor U532 (N_532,N_403,N_461);
nand U533 (N_533,N_442,N_473);
nand U534 (N_534,N_481,N_416);
and U535 (N_535,N_482,N_437);
or U536 (N_536,N_491,N_422);
nand U537 (N_537,N_457,N_445);
nand U538 (N_538,N_462,N_431);
nor U539 (N_539,N_412,N_460);
nand U540 (N_540,N_455,N_404);
or U541 (N_541,N_463,N_448);
or U542 (N_542,N_465,N_464);
nor U543 (N_543,N_417,N_401);
and U544 (N_544,N_419,N_474);
and U545 (N_545,N_479,N_425);
and U546 (N_546,N_427,N_488);
xnor U547 (N_547,N_432,N_424);
nor U548 (N_548,N_418,N_450);
and U549 (N_549,N_420,N_410);
or U550 (N_550,N_442,N_448);
and U551 (N_551,N_400,N_448);
or U552 (N_552,N_472,N_496);
and U553 (N_553,N_459,N_472);
and U554 (N_554,N_465,N_466);
and U555 (N_555,N_418,N_473);
or U556 (N_556,N_471,N_444);
and U557 (N_557,N_475,N_437);
and U558 (N_558,N_413,N_464);
or U559 (N_559,N_412,N_432);
nand U560 (N_560,N_467,N_487);
or U561 (N_561,N_466,N_492);
and U562 (N_562,N_410,N_479);
nor U563 (N_563,N_459,N_457);
nor U564 (N_564,N_428,N_435);
nor U565 (N_565,N_479,N_407);
nand U566 (N_566,N_418,N_426);
nor U567 (N_567,N_410,N_433);
nor U568 (N_568,N_428,N_484);
and U569 (N_569,N_437,N_451);
or U570 (N_570,N_488,N_418);
nand U571 (N_571,N_463,N_461);
or U572 (N_572,N_404,N_482);
nand U573 (N_573,N_444,N_459);
and U574 (N_574,N_474,N_494);
and U575 (N_575,N_420,N_479);
and U576 (N_576,N_417,N_481);
or U577 (N_577,N_474,N_411);
nand U578 (N_578,N_458,N_456);
and U579 (N_579,N_455,N_417);
and U580 (N_580,N_462,N_491);
nand U581 (N_581,N_429,N_481);
nor U582 (N_582,N_462,N_483);
nand U583 (N_583,N_488,N_456);
or U584 (N_584,N_489,N_415);
or U585 (N_585,N_428,N_447);
nor U586 (N_586,N_448,N_441);
and U587 (N_587,N_468,N_443);
nand U588 (N_588,N_408,N_456);
and U589 (N_589,N_472,N_423);
or U590 (N_590,N_445,N_498);
nor U591 (N_591,N_415,N_427);
or U592 (N_592,N_498,N_468);
or U593 (N_593,N_441,N_426);
nand U594 (N_594,N_432,N_454);
nand U595 (N_595,N_475,N_421);
nor U596 (N_596,N_493,N_441);
nor U597 (N_597,N_407,N_456);
or U598 (N_598,N_434,N_439);
or U599 (N_599,N_401,N_408);
and U600 (N_600,N_529,N_582);
and U601 (N_601,N_566,N_513);
and U602 (N_602,N_533,N_525);
nand U603 (N_603,N_593,N_548);
or U604 (N_604,N_505,N_550);
and U605 (N_605,N_547,N_549);
nor U606 (N_606,N_531,N_536);
or U607 (N_607,N_563,N_567);
nor U608 (N_608,N_517,N_576);
nand U609 (N_609,N_581,N_561);
nor U610 (N_610,N_503,N_569);
and U611 (N_611,N_542,N_575);
and U612 (N_612,N_577,N_580);
and U613 (N_613,N_526,N_532);
and U614 (N_614,N_565,N_589);
nor U615 (N_615,N_543,N_507);
nor U616 (N_616,N_516,N_506);
nor U617 (N_617,N_579,N_590);
nor U618 (N_618,N_524,N_508);
or U619 (N_619,N_596,N_521);
or U620 (N_620,N_553,N_591);
and U621 (N_621,N_594,N_538);
nor U622 (N_622,N_510,N_523);
or U623 (N_623,N_573,N_587);
xnor U624 (N_624,N_551,N_592);
xor U625 (N_625,N_520,N_546);
or U626 (N_626,N_501,N_555);
or U627 (N_627,N_530,N_583);
nor U628 (N_628,N_595,N_541);
and U629 (N_629,N_512,N_571);
and U630 (N_630,N_578,N_519);
and U631 (N_631,N_509,N_511);
nand U632 (N_632,N_544,N_557);
nand U633 (N_633,N_522,N_515);
nor U634 (N_634,N_554,N_570);
nand U635 (N_635,N_500,N_535);
and U636 (N_636,N_568,N_558);
nor U637 (N_637,N_504,N_540);
nor U638 (N_638,N_585,N_559);
and U639 (N_639,N_552,N_599);
nand U640 (N_640,N_572,N_534);
and U641 (N_641,N_597,N_584);
nor U642 (N_642,N_598,N_586);
and U643 (N_643,N_518,N_537);
nand U644 (N_644,N_562,N_545);
nor U645 (N_645,N_556,N_539);
and U646 (N_646,N_502,N_588);
and U647 (N_647,N_514,N_528);
nor U648 (N_648,N_564,N_574);
and U649 (N_649,N_560,N_527);
and U650 (N_650,N_573,N_537);
nor U651 (N_651,N_551,N_513);
or U652 (N_652,N_578,N_571);
or U653 (N_653,N_531,N_524);
nor U654 (N_654,N_576,N_560);
nor U655 (N_655,N_548,N_536);
nand U656 (N_656,N_513,N_565);
nand U657 (N_657,N_530,N_575);
nand U658 (N_658,N_586,N_566);
or U659 (N_659,N_528,N_538);
nand U660 (N_660,N_558,N_589);
and U661 (N_661,N_540,N_533);
or U662 (N_662,N_552,N_508);
nand U663 (N_663,N_516,N_543);
or U664 (N_664,N_582,N_519);
or U665 (N_665,N_569,N_570);
nand U666 (N_666,N_580,N_516);
nand U667 (N_667,N_521,N_586);
and U668 (N_668,N_570,N_558);
and U669 (N_669,N_508,N_550);
or U670 (N_670,N_599,N_541);
and U671 (N_671,N_524,N_537);
nor U672 (N_672,N_569,N_555);
nor U673 (N_673,N_564,N_593);
or U674 (N_674,N_580,N_506);
or U675 (N_675,N_560,N_570);
nand U676 (N_676,N_541,N_523);
nor U677 (N_677,N_525,N_557);
nand U678 (N_678,N_513,N_536);
nand U679 (N_679,N_540,N_550);
nand U680 (N_680,N_572,N_503);
and U681 (N_681,N_549,N_555);
nand U682 (N_682,N_560,N_526);
nand U683 (N_683,N_569,N_583);
or U684 (N_684,N_518,N_588);
nand U685 (N_685,N_532,N_579);
nor U686 (N_686,N_533,N_576);
nor U687 (N_687,N_586,N_559);
nor U688 (N_688,N_557,N_513);
nand U689 (N_689,N_543,N_560);
and U690 (N_690,N_552,N_597);
nor U691 (N_691,N_531,N_587);
nand U692 (N_692,N_594,N_548);
and U693 (N_693,N_535,N_541);
nor U694 (N_694,N_585,N_518);
and U695 (N_695,N_501,N_540);
or U696 (N_696,N_559,N_584);
nand U697 (N_697,N_543,N_596);
nand U698 (N_698,N_575,N_502);
nor U699 (N_699,N_524,N_513);
and U700 (N_700,N_697,N_612);
or U701 (N_701,N_638,N_661);
nand U702 (N_702,N_615,N_665);
or U703 (N_703,N_620,N_647);
or U704 (N_704,N_683,N_637);
nor U705 (N_705,N_660,N_698);
nand U706 (N_706,N_696,N_672);
or U707 (N_707,N_674,N_682);
nor U708 (N_708,N_684,N_602);
nor U709 (N_709,N_687,N_690);
or U710 (N_710,N_623,N_626);
nor U711 (N_711,N_613,N_617);
or U712 (N_712,N_654,N_633);
nor U713 (N_713,N_688,N_629);
nor U714 (N_714,N_656,N_607);
nor U715 (N_715,N_679,N_622);
and U716 (N_716,N_618,N_662);
nand U717 (N_717,N_643,N_680);
nor U718 (N_718,N_653,N_636);
and U719 (N_719,N_692,N_670);
or U720 (N_720,N_668,N_673);
and U721 (N_721,N_628,N_610);
or U722 (N_722,N_646,N_601);
or U723 (N_723,N_695,N_603);
nor U724 (N_724,N_663,N_664);
nor U725 (N_725,N_666,N_657);
and U726 (N_726,N_616,N_686);
nor U727 (N_727,N_675,N_651);
or U728 (N_728,N_650,N_625);
nor U729 (N_729,N_677,N_669);
or U730 (N_730,N_699,N_641);
and U731 (N_731,N_667,N_685);
nor U732 (N_732,N_635,N_606);
nand U733 (N_733,N_605,N_645);
and U734 (N_734,N_614,N_691);
nor U735 (N_735,N_604,N_678);
or U736 (N_736,N_640,N_648);
and U737 (N_737,N_639,N_611);
and U738 (N_738,N_658,N_642);
nand U739 (N_739,N_630,N_609);
nand U740 (N_740,N_608,N_649);
nor U741 (N_741,N_631,N_693);
nor U742 (N_742,N_621,N_634);
or U743 (N_743,N_689,N_681);
or U744 (N_744,N_694,N_652);
or U745 (N_745,N_671,N_659);
and U746 (N_746,N_600,N_644);
or U747 (N_747,N_632,N_627);
and U748 (N_748,N_619,N_655);
nor U749 (N_749,N_624,N_676);
nor U750 (N_750,N_660,N_642);
and U751 (N_751,N_628,N_682);
nand U752 (N_752,N_648,N_607);
or U753 (N_753,N_600,N_666);
or U754 (N_754,N_665,N_694);
nand U755 (N_755,N_630,N_685);
and U756 (N_756,N_692,N_653);
nor U757 (N_757,N_687,N_676);
nor U758 (N_758,N_612,N_686);
nand U759 (N_759,N_677,N_653);
nand U760 (N_760,N_633,N_615);
or U761 (N_761,N_666,N_632);
nand U762 (N_762,N_674,N_600);
and U763 (N_763,N_603,N_655);
and U764 (N_764,N_658,N_694);
nand U765 (N_765,N_643,N_687);
and U766 (N_766,N_657,N_662);
and U767 (N_767,N_687,N_689);
or U768 (N_768,N_625,N_662);
nor U769 (N_769,N_670,N_697);
or U770 (N_770,N_644,N_671);
xnor U771 (N_771,N_608,N_610);
or U772 (N_772,N_681,N_677);
nand U773 (N_773,N_631,N_639);
or U774 (N_774,N_614,N_641);
nand U775 (N_775,N_613,N_657);
or U776 (N_776,N_658,N_647);
nor U777 (N_777,N_672,N_642);
nand U778 (N_778,N_669,N_609);
and U779 (N_779,N_695,N_693);
xor U780 (N_780,N_639,N_669);
nor U781 (N_781,N_693,N_606);
or U782 (N_782,N_634,N_680);
nor U783 (N_783,N_673,N_661);
nand U784 (N_784,N_641,N_602);
nor U785 (N_785,N_680,N_636);
xnor U786 (N_786,N_630,N_694);
and U787 (N_787,N_669,N_666);
and U788 (N_788,N_648,N_674);
or U789 (N_789,N_668,N_608);
nor U790 (N_790,N_648,N_609);
and U791 (N_791,N_670,N_637);
and U792 (N_792,N_623,N_610);
nor U793 (N_793,N_691,N_625);
and U794 (N_794,N_627,N_634);
or U795 (N_795,N_662,N_659);
nor U796 (N_796,N_651,N_617);
nor U797 (N_797,N_678,N_631);
nand U798 (N_798,N_678,N_698);
nand U799 (N_799,N_679,N_654);
nand U800 (N_800,N_737,N_784);
or U801 (N_801,N_730,N_707);
or U802 (N_802,N_787,N_708);
nor U803 (N_803,N_755,N_791);
and U804 (N_804,N_709,N_714);
nand U805 (N_805,N_721,N_736);
and U806 (N_806,N_726,N_735);
nand U807 (N_807,N_754,N_780);
or U808 (N_808,N_706,N_744);
and U809 (N_809,N_731,N_774);
nor U810 (N_810,N_712,N_720);
and U811 (N_811,N_738,N_700);
nand U812 (N_812,N_777,N_782);
nand U813 (N_813,N_725,N_788);
and U814 (N_814,N_775,N_778);
nand U815 (N_815,N_749,N_747);
or U816 (N_816,N_770,N_794);
nand U817 (N_817,N_776,N_760);
nand U818 (N_818,N_757,N_727);
and U819 (N_819,N_773,N_789);
nand U820 (N_820,N_715,N_783);
or U821 (N_821,N_758,N_764);
or U822 (N_822,N_769,N_786);
and U823 (N_823,N_701,N_702);
nor U824 (N_824,N_723,N_753);
or U825 (N_825,N_761,N_740);
nor U826 (N_826,N_781,N_741);
and U827 (N_827,N_705,N_743);
nor U828 (N_828,N_797,N_713);
and U829 (N_829,N_768,N_745);
or U830 (N_830,N_722,N_739);
nand U831 (N_831,N_718,N_798);
and U832 (N_832,N_750,N_795);
nand U833 (N_833,N_762,N_742);
or U834 (N_834,N_704,N_759);
or U835 (N_835,N_711,N_796);
or U836 (N_836,N_729,N_703);
nand U837 (N_837,N_765,N_716);
nand U838 (N_838,N_746,N_724);
and U839 (N_839,N_717,N_751);
nand U840 (N_840,N_771,N_728);
nor U841 (N_841,N_799,N_734);
or U842 (N_842,N_733,N_779);
xnor U843 (N_843,N_767,N_772);
or U844 (N_844,N_792,N_785);
or U845 (N_845,N_766,N_756);
nand U846 (N_846,N_732,N_748);
nor U847 (N_847,N_719,N_793);
and U848 (N_848,N_763,N_790);
nand U849 (N_849,N_752,N_710);
or U850 (N_850,N_777,N_703);
nor U851 (N_851,N_727,N_783);
nor U852 (N_852,N_781,N_738);
or U853 (N_853,N_798,N_774);
nor U854 (N_854,N_776,N_747);
nor U855 (N_855,N_736,N_702);
and U856 (N_856,N_755,N_702);
xnor U857 (N_857,N_772,N_722);
nor U858 (N_858,N_796,N_710);
and U859 (N_859,N_728,N_726);
or U860 (N_860,N_719,N_760);
and U861 (N_861,N_743,N_797);
nor U862 (N_862,N_794,N_735);
or U863 (N_863,N_794,N_732);
nand U864 (N_864,N_782,N_773);
and U865 (N_865,N_789,N_754);
nand U866 (N_866,N_758,N_735);
nor U867 (N_867,N_778,N_709);
and U868 (N_868,N_761,N_722);
and U869 (N_869,N_788,N_700);
and U870 (N_870,N_722,N_727);
or U871 (N_871,N_773,N_779);
or U872 (N_872,N_709,N_724);
nand U873 (N_873,N_766,N_748);
and U874 (N_874,N_786,N_757);
nand U875 (N_875,N_718,N_788);
and U876 (N_876,N_782,N_738);
or U877 (N_877,N_739,N_782);
or U878 (N_878,N_701,N_758);
nor U879 (N_879,N_704,N_736);
nand U880 (N_880,N_744,N_778);
nand U881 (N_881,N_722,N_793);
and U882 (N_882,N_743,N_766);
and U883 (N_883,N_793,N_713);
nor U884 (N_884,N_720,N_739);
nand U885 (N_885,N_740,N_789);
and U886 (N_886,N_744,N_700);
or U887 (N_887,N_732,N_728);
nor U888 (N_888,N_739,N_715);
or U889 (N_889,N_701,N_754);
and U890 (N_890,N_715,N_794);
nor U891 (N_891,N_781,N_767);
or U892 (N_892,N_735,N_713);
nor U893 (N_893,N_789,N_795);
or U894 (N_894,N_741,N_703);
nor U895 (N_895,N_771,N_740);
or U896 (N_896,N_754,N_730);
nand U897 (N_897,N_704,N_744);
and U898 (N_898,N_711,N_740);
nor U899 (N_899,N_706,N_777);
and U900 (N_900,N_864,N_822);
nand U901 (N_901,N_895,N_891);
nand U902 (N_902,N_857,N_873);
or U903 (N_903,N_889,N_842);
and U904 (N_904,N_869,N_877);
nand U905 (N_905,N_893,N_820);
nor U906 (N_906,N_847,N_868);
and U907 (N_907,N_802,N_844);
nor U908 (N_908,N_801,N_882);
and U909 (N_909,N_828,N_848);
and U910 (N_910,N_858,N_826);
or U911 (N_911,N_843,N_841);
or U912 (N_912,N_852,N_897);
and U913 (N_913,N_839,N_890);
or U914 (N_914,N_871,N_845);
nand U915 (N_915,N_833,N_892);
nor U916 (N_916,N_836,N_837);
or U917 (N_917,N_888,N_816);
or U918 (N_918,N_886,N_814);
nand U919 (N_919,N_863,N_806);
or U920 (N_920,N_812,N_883);
xor U921 (N_921,N_887,N_832);
nand U922 (N_922,N_804,N_805);
nor U923 (N_923,N_808,N_870);
nand U924 (N_924,N_854,N_809);
or U925 (N_925,N_851,N_821);
or U926 (N_926,N_876,N_838);
and U927 (N_927,N_861,N_818);
and U928 (N_928,N_899,N_831);
or U929 (N_929,N_815,N_827);
nand U930 (N_930,N_803,N_894);
and U931 (N_931,N_829,N_866);
and U932 (N_932,N_855,N_862);
nand U933 (N_933,N_872,N_898);
and U934 (N_934,N_811,N_823);
nand U935 (N_935,N_819,N_834);
nand U936 (N_936,N_867,N_853);
and U937 (N_937,N_859,N_865);
nor U938 (N_938,N_896,N_846);
nor U939 (N_939,N_875,N_830);
nor U940 (N_940,N_813,N_824);
nor U941 (N_941,N_849,N_874);
nand U942 (N_942,N_880,N_881);
nand U943 (N_943,N_817,N_856);
nor U944 (N_944,N_807,N_825);
nand U945 (N_945,N_879,N_810);
nor U946 (N_946,N_878,N_860);
nor U947 (N_947,N_800,N_850);
nand U948 (N_948,N_885,N_835);
nand U949 (N_949,N_884,N_840);
nor U950 (N_950,N_820,N_808);
and U951 (N_951,N_890,N_860);
or U952 (N_952,N_859,N_863);
nor U953 (N_953,N_837,N_890);
nor U954 (N_954,N_863,N_891);
nand U955 (N_955,N_879,N_864);
nand U956 (N_956,N_829,N_824);
and U957 (N_957,N_838,N_880);
and U958 (N_958,N_870,N_801);
nor U959 (N_959,N_853,N_823);
nand U960 (N_960,N_868,N_846);
nor U961 (N_961,N_803,N_811);
and U962 (N_962,N_884,N_883);
nand U963 (N_963,N_867,N_859);
nand U964 (N_964,N_862,N_810);
and U965 (N_965,N_806,N_867);
nor U966 (N_966,N_811,N_889);
or U967 (N_967,N_882,N_842);
and U968 (N_968,N_825,N_809);
and U969 (N_969,N_827,N_831);
and U970 (N_970,N_885,N_880);
or U971 (N_971,N_844,N_800);
and U972 (N_972,N_855,N_817);
or U973 (N_973,N_867,N_817);
nor U974 (N_974,N_869,N_859);
and U975 (N_975,N_899,N_850);
and U976 (N_976,N_820,N_884);
and U977 (N_977,N_873,N_854);
nand U978 (N_978,N_838,N_800);
nor U979 (N_979,N_888,N_897);
and U980 (N_980,N_804,N_860);
nand U981 (N_981,N_834,N_803);
and U982 (N_982,N_824,N_850);
nand U983 (N_983,N_800,N_845);
nor U984 (N_984,N_884,N_800);
or U985 (N_985,N_830,N_854);
nand U986 (N_986,N_882,N_802);
nand U987 (N_987,N_843,N_893);
nand U988 (N_988,N_827,N_870);
nor U989 (N_989,N_866,N_805);
nand U990 (N_990,N_878,N_891);
or U991 (N_991,N_890,N_877);
nor U992 (N_992,N_860,N_855);
nand U993 (N_993,N_836,N_817);
and U994 (N_994,N_839,N_829);
nor U995 (N_995,N_868,N_845);
or U996 (N_996,N_861,N_866);
nor U997 (N_997,N_872,N_808);
xnor U998 (N_998,N_860,N_854);
and U999 (N_999,N_848,N_822);
or U1000 (N_1000,N_979,N_927);
nor U1001 (N_1001,N_956,N_904);
nand U1002 (N_1002,N_992,N_987);
nand U1003 (N_1003,N_953,N_900);
or U1004 (N_1004,N_912,N_950);
and U1005 (N_1005,N_917,N_994);
or U1006 (N_1006,N_942,N_935);
nand U1007 (N_1007,N_924,N_990);
and U1008 (N_1008,N_952,N_941);
and U1009 (N_1009,N_929,N_985);
nand U1010 (N_1010,N_939,N_969);
and U1011 (N_1011,N_978,N_991);
nand U1012 (N_1012,N_928,N_975);
nor U1013 (N_1013,N_993,N_937);
and U1014 (N_1014,N_946,N_998);
nor U1015 (N_1015,N_971,N_967);
or U1016 (N_1016,N_945,N_910);
and U1017 (N_1017,N_960,N_902);
or U1018 (N_1018,N_908,N_958);
or U1019 (N_1019,N_966,N_947);
and U1020 (N_1020,N_964,N_957);
nor U1021 (N_1021,N_954,N_988);
nand U1022 (N_1022,N_923,N_920);
nor U1023 (N_1023,N_948,N_918);
nor U1024 (N_1024,N_921,N_999);
nand U1025 (N_1025,N_911,N_905);
and U1026 (N_1026,N_933,N_949);
nor U1027 (N_1027,N_907,N_961);
or U1028 (N_1028,N_909,N_972);
nand U1029 (N_1029,N_915,N_903);
nand U1030 (N_1030,N_984,N_944);
nor U1031 (N_1031,N_932,N_973);
nor U1032 (N_1032,N_997,N_943);
or U1033 (N_1033,N_936,N_901);
nor U1034 (N_1034,N_919,N_968);
xnor U1035 (N_1035,N_938,N_989);
nand U1036 (N_1036,N_977,N_934);
or U1037 (N_1037,N_996,N_995);
or U1038 (N_1038,N_962,N_974);
and U1039 (N_1039,N_963,N_982);
nor U1040 (N_1040,N_930,N_940);
and U1041 (N_1041,N_955,N_906);
nor U1042 (N_1042,N_913,N_925);
and U1043 (N_1043,N_922,N_916);
or U1044 (N_1044,N_926,N_914);
nand U1045 (N_1045,N_980,N_951);
nor U1046 (N_1046,N_986,N_983);
nand U1047 (N_1047,N_965,N_931);
or U1048 (N_1048,N_970,N_959);
nand U1049 (N_1049,N_981,N_976);
nand U1050 (N_1050,N_978,N_920);
nor U1051 (N_1051,N_964,N_997);
and U1052 (N_1052,N_937,N_915);
and U1053 (N_1053,N_930,N_912);
nor U1054 (N_1054,N_999,N_928);
and U1055 (N_1055,N_900,N_967);
nand U1056 (N_1056,N_955,N_995);
nor U1057 (N_1057,N_976,N_923);
nor U1058 (N_1058,N_933,N_908);
or U1059 (N_1059,N_908,N_914);
or U1060 (N_1060,N_918,N_982);
and U1061 (N_1061,N_925,N_910);
nand U1062 (N_1062,N_904,N_903);
and U1063 (N_1063,N_995,N_982);
nor U1064 (N_1064,N_950,N_986);
nor U1065 (N_1065,N_915,N_923);
nor U1066 (N_1066,N_911,N_939);
and U1067 (N_1067,N_933,N_942);
nor U1068 (N_1068,N_957,N_995);
or U1069 (N_1069,N_985,N_941);
and U1070 (N_1070,N_960,N_936);
nand U1071 (N_1071,N_940,N_941);
nand U1072 (N_1072,N_928,N_909);
nor U1073 (N_1073,N_972,N_975);
nand U1074 (N_1074,N_919,N_979);
nor U1075 (N_1075,N_969,N_934);
nand U1076 (N_1076,N_930,N_962);
nand U1077 (N_1077,N_928,N_922);
and U1078 (N_1078,N_977,N_912);
nand U1079 (N_1079,N_930,N_925);
nor U1080 (N_1080,N_920,N_970);
nor U1081 (N_1081,N_948,N_999);
nand U1082 (N_1082,N_983,N_926);
or U1083 (N_1083,N_963,N_956);
nand U1084 (N_1084,N_936,N_942);
xnor U1085 (N_1085,N_986,N_978);
xnor U1086 (N_1086,N_953,N_985);
and U1087 (N_1087,N_934,N_961);
or U1088 (N_1088,N_948,N_949);
nor U1089 (N_1089,N_917,N_918);
nor U1090 (N_1090,N_936,N_934);
nor U1091 (N_1091,N_963,N_989);
nor U1092 (N_1092,N_940,N_938);
nand U1093 (N_1093,N_978,N_932);
nor U1094 (N_1094,N_908,N_962);
or U1095 (N_1095,N_986,N_908);
and U1096 (N_1096,N_990,N_902);
nor U1097 (N_1097,N_967,N_978);
or U1098 (N_1098,N_914,N_933);
nor U1099 (N_1099,N_976,N_999);
or U1100 (N_1100,N_1045,N_1055);
xnor U1101 (N_1101,N_1089,N_1094);
or U1102 (N_1102,N_1072,N_1048);
nand U1103 (N_1103,N_1076,N_1010);
nor U1104 (N_1104,N_1011,N_1033);
and U1105 (N_1105,N_1014,N_1073);
and U1106 (N_1106,N_1092,N_1084);
nor U1107 (N_1107,N_1025,N_1003);
nor U1108 (N_1108,N_1052,N_1082);
and U1109 (N_1109,N_1057,N_1016);
xor U1110 (N_1110,N_1059,N_1032);
nor U1111 (N_1111,N_1001,N_1031);
nor U1112 (N_1112,N_1026,N_1098);
or U1113 (N_1113,N_1077,N_1028);
or U1114 (N_1114,N_1008,N_1021);
nand U1115 (N_1115,N_1051,N_1054);
or U1116 (N_1116,N_1000,N_1038);
and U1117 (N_1117,N_1037,N_1058);
and U1118 (N_1118,N_1063,N_1060);
nand U1119 (N_1119,N_1086,N_1080);
or U1120 (N_1120,N_1056,N_1044);
nand U1121 (N_1121,N_1034,N_1066);
nor U1122 (N_1122,N_1009,N_1049);
or U1123 (N_1123,N_1039,N_1036);
nor U1124 (N_1124,N_1012,N_1071);
nor U1125 (N_1125,N_1046,N_1081);
or U1126 (N_1126,N_1015,N_1053);
or U1127 (N_1127,N_1043,N_1027);
and U1128 (N_1128,N_1020,N_1007);
nand U1129 (N_1129,N_1017,N_1042);
and U1130 (N_1130,N_1097,N_1040);
nor U1131 (N_1131,N_1022,N_1047);
or U1132 (N_1132,N_1024,N_1029);
nor U1133 (N_1133,N_1095,N_1041);
and U1134 (N_1134,N_1075,N_1013);
and U1135 (N_1135,N_1050,N_1078);
nand U1136 (N_1136,N_1064,N_1070);
nand U1137 (N_1137,N_1067,N_1090);
or U1138 (N_1138,N_1099,N_1096);
or U1139 (N_1139,N_1079,N_1083);
and U1140 (N_1140,N_1087,N_1023);
or U1141 (N_1141,N_1088,N_1068);
or U1142 (N_1142,N_1093,N_1062);
and U1143 (N_1143,N_1018,N_1061);
nor U1144 (N_1144,N_1002,N_1069);
or U1145 (N_1145,N_1074,N_1030);
or U1146 (N_1146,N_1005,N_1004);
or U1147 (N_1147,N_1091,N_1085);
nor U1148 (N_1148,N_1065,N_1006);
nand U1149 (N_1149,N_1019,N_1035);
or U1150 (N_1150,N_1020,N_1022);
and U1151 (N_1151,N_1087,N_1086);
or U1152 (N_1152,N_1059,N_1064);
nor U1153 (N_1153,N_1027,N_1034);
nand U1154 (N_1154,N_1044,N_1013);
nand U1155 (N_1155,N_1078,N_1028);
and U1156 (N_1156,N_1004,N_1024);
nand U1157 (N_1157,N_1069,N_1067);
and U1158 (N_1158,N_1050,N_1011);
nor U1159 (N_1159,N_1058,N_1098);
or U1160 (N_1160,N_1017,N_1020);
or U1161 (N_1161,N_1022,N_1076);
or U1162 (N_1162,N_1079,N_1098);
nand U1163 (N_1163,N_1054,N_1080);
nor U1164 (N_1164,N_1051,N_1057);
and U1165 (N_1165,N_1018,N_1087);
nor U1166 (N_1166,N_1037,N_1057);
or U1167 (N_1167,N_1095,N_1036);
nand U1168 (N_1168,N_1091,N_1071);
and U1169 (N_1169,N_1068,N_1096);
and U1170 (N_1170,N_1054,N_1034);
nor U1171 (N_1171,N_1077,N_1083);
nand U1172 (N_1172,N_1019,N_1029);
nor U1173 (N_1173,N_1063,N_1033);
and U1174 (N_1174,N_1024,N_1016);
or U1175 (N_1175,N_1079,N_1076);
or U1176 (N_1176,N_1072,N_1061);
nor U1177 (N_1177,N_1041,N_1069);
and U1178 (N_1178,N_1049,N_1012);
and U1179 (N_1179,N_1098,N_1027);
or U1180 (N_1180,N_1014,N_1041);
and U1181 (N_1181,N_1017,N_1043);
nand U1182 (N_1182,N_1022,N_1007);
and U1183 (N_1183,N_1027,N_1025);
and U1184 (N_1184,N_1053,N_1034);
or U1185 (N_1185,N_1046,N_1032);
nor U1186 (N_1186,N_1072,N_1051);
and U1187 (N_1187,N_1057,N_1095);
nor U1188 (N_1188,N_1027,N_1015);
nor U1189 (N_1189,N_1028,N_1027);
or U1190 (N_1190,N_1021,N_1098);
nand U1191 (N_1191,N_1009,N_1087);
or U1192 (N_1192,N_1024,N_1097);
nand U1193 (N_1193,N_1072,N_1082);
nor U1194 (N_1194,N_1073,N_1054);
nand U1195 (N_1195,N_1038,N_1081);
nand U1196 (N_1196,N_1039,N_1093);
nand U1197 (N_1197,N_1025,N_1009);
and U1198 (N_1198,N_1061,N_1050);
and U1199 (N_1199,N_1096,N_1034);
nor U1200 (N_1200,N_1111,N_1149);
and U1201 (N_1201,N_1141,N_1121);
or U1202 (N_1202,N_1129,N_1183);
and U1203 (N_1203,N_1194,N_1152);
nand U1204 (N_1204,N_1148,N_1184);
nand U1205 (N_1205,N_1124,N_1190);
or U1206 (N_1206,N_1117,N_1122);
and U1207 (N_1207,N_1134,N_1158);
or U1208 (N_1208,N_1116,N_1188);
or U1209 (N_1209,N_1176,N_1160);
nand U1210 (N_1210,N_1145,N_1123);
or U1211 (N_1211,N_1197,N_1139);
nor U1212 (N_1212,N_1171,N_1127);
and U1213 (N_1213,N_1196,N_1168);
nand U1214 (N_1214,N_1110,N_1164);
nor U1215 (N_1215,N_1104,N_1114);
and U1216 (N_1216,N_1172,N_1178);
nor U1217 (N_1217,N_1173,N_1137);
or U1218 (N_1218,N_1108,N_1159);
nand U1219 (N_1219,N_1130,N_1179);
and U1220 (N_1220,N_1199,N_1120);
or U1221 (N_1221,N_1140,N_1132);
and U1222 (N_1222,N_1103,N_1170);
or U1223 (N_1223,N_1192,N_1115);
nand U1224 (N_1224,N_1185,N_1175);
nor U1225 (N_1225,N_1156,N_1186);
nand U1226 (N_1226,N_1154,N_1151);
nand U1227 (N_1227,N_1131,N_1109);
nor U1228 (N_1228,N_1118,N_1112);
and U1229 (N_1229,N_1177,N_1138);
and U1230 (N_1230,N_1187,N_1163);
nor U1231 (N_1231,N_1143,N_1144);
nor U1232 (N_1232,N_1135,N_1198);
or U1233 (N_1233,N_1146,N_1155);
nand U1234 (N_1234,N_1100,N_1102);
or U1235 (N_1235,N_1101,N_1195);
nand U1236 (N_1236,N_1191,N_1128);
nand U1237 (N_1237,N_1107,N_1147);
and U1238 (N_1238,N_1189,N_1162);
and U1239 (N_1239,N_1133,N_1105);
nand U1240 (N_1240,N_1119,N_1181);
nor U1241 (N_1241,N_1166,N_1169);
nor U1242 (N_1242,N_1142,N_1150);
and U1243 (N_1243,N_1126,N_1180);
or U1244 (N_1244,N_1174,N_1167);
nand U1245 (N_1245,N_1157,N_1161);
and U1246 (N_1246,N_1106,N_1193);
nor U1247 (N_1247,N_1165,N_1113);
and U1248 (N_1248,N_1136,N_1182);
or U1249 (N_1249,N_1125,N_1153);
and U1250 (N_1250,N_1143,N_1124);
and U1251 (N_1251,N_1154,N_1175);
nand U1252 (N_1252,N_1148,N_1129);
nor U1253 (N_1253,N_1118,N_1176);
nand U1254 (N_1254,N_1139,N_1183);
nand U1255 (N_1255,N_1176,N_1183);
nor U1256 (N_1256,N_1151,N_1159);
nor U1257 (N_1257,N_1142,N_1126);
and U1258 (N_1258,N_1121,N_1134);
nand U1259 (N_1259,N_1158,N_1123);
nor U1260 (N_1260,N_1140,N_1116);
or U1261 (N_1261,N_1198,N_1188);
nand U1262 (N_1262,N_1139,N_1145);
or U1263 (N_1263,N_1107,N_1121);
xnor U1264 (N_1264,N_1175,N_1110);
nor U1265 (N_1265,N_1135,N_1101);
and U1266 (N_1266,N_1134,N_1116);
nand U1267 (N_1267,N_1146,N_1180);
or U1268 (N_1268,N_1184,N_1198);
nand U1269 (N_1269,N_1121,N_1118);
nand U1270 (N_1270,N_1146,N_1162);
nand U1271 (N_1271,N_1113,N_1171);
or U1272 (N_1272,N_1169,N_1104);
nand U1273 (N_1273,N_1172,N_1152);
and U1274 (N_1274,N_1109,N_1127);
and U1275 (N_1275,N_1184,N_1132);
or U1276 (N_1276,N_1118,N_1161);
nand U1277 (N_1277,N_1167,N_1112);
nand U1278 (N_1278,N_1188,N_1163);
and U1279 (N_1279,N_1191,N_1132);
nor U1280 (N_1280,N_1156,N_1170);
nor U1281 (N_1281,N_1109,N_1102);
nand U1282 (N_1282,N_1145,N_1165);
nor U1283 (N_1283,N_1193,N_1141);
nand U1284 (N_1284,N_1167,N_1155);
and U1285 (N_1285,N_1141,N_1172);
or U1286 (N_1286,N_1142,N_1183);
nand U1287 (N_1287,N_1163,N_1180);
nor U1288 (N_1288,N_1142,N_1122);
nand U1289 (N_1289,N_1147,N_1161);
or U1290 (N_1290,N_1120,N_1101);
nand U1291 (N_1291,N_1167,N_1188);
nor U1292 (N_1292,N_1134,N_1191);
nand U1293 (N_1293,N_1111,N_1145);
nand U1294 (N_1294,N_1142,N_1110);
nand U1295 (N_1295,N_1134,N_1125);
and U1296 (N_1296,N_1194,N_1177);
and U1297 (N_1297,N_1103,N_1118);
and U1298 (N_1298,N_1138,N_1131);
nor U1299 (N_1299,N_1184,N_1178);
nand U1300 (N_1300,N_1248,N_1244);
and U1301 (N_1301,N_1292,N_1275);
nand U1302 (N_1302,N_1206,N_1269);
nor U1303 (N_1303,N_1286,N_1231);
nor U1304 (N_1304,N_1213,N_1276);
or U1305 (N_1305,N_1280,N_1209);
or U1306 (N_1306,N_1237,N_1241);
and U1307 (N_1307,N_1258,N_1218);
or U1308 (N_1308,N_1225,N_1262);
and U1309 (N_1309,N_1203,N_1265);
nand U1310 (N_1310,N_1243,N_1205);
and U1311 (N_1311,N_1207,N_1268);
and U1312 (N_1312,N_1222,N_1297);
or U1313 (N_1313,N_1228,N_1247);
and U1314 (N_1314,N_1270,N_1226);
nor U1315 (N_1315,N_1261,N_1285);
and U1316 (N_1316,N_1236,N_1249);
nor U1317 (N_1317,N_1278,N_1293);
nor U1318 (N_1318,N_1257,N_1245);
and U1319 (N_1319,N_1284,N_1215);
and U1320 (N_1320,N_1252,N_1271);
nand U1321 (N_1321,N_1290,N_1251);
or U1322 (N_1322,N_1233,N_1201);
nand U1323 (N_1323,N_1224,N_1204);
or U1324 (N_1324,N_1277,N_1232);
nand U1325 (N_1325,N_1264,N_1240);
nand U1326 (N_1326,N_1294,N_1260);
nand U1327 (N_1327,N_1279,N_1229);
nand U1328 (N_1328,N_1230,N_1256);
nand U1329 (N_1329,N_1242,N_1223);
or U1330 (N_1330,N_1219,N_1239);
and U1331 (N_1331,N_1221,N_1298);
nand U1332 (N_1332,N_1235,N_1266);
and U1333 (N_1333,N_1212,N_1267);
or U1334 (N_1334,N_1289,N_1227);
or U1335 (N_1335,N_1255,N_1234);
nand U1336 (N_1336,N_1259,N_1210);
nand U1337 (N_1337,N_1272,N_1238);
and U1338 (N_1338,N_1214,N_1246);
or U1339 (N_1339,N_1217,N_1200);
nor U1340 (N_1340,N_1263,N_1208);
nand U1341 (N_1341,N_1211,N_1273);
nand U1342 (N_1342,N_1254,N_1250);
and U1343 (N_1343,N_1287,N_1202);
nand U1344 (N_1344,N_1274,N_1282);
or U1345 (N_1345,N_1283,N_1220);
or U1346 (N_1346,N_1216,N_1281);
or U1347 (N_1347,N_1288,N_1253);
and U1348 (N_1348,N_1295,N_1296);
nand U1349 (N_1349,N_1291,N_1299);
nor U1350 (N_1350,N_1239,N_1216);
or U1351 (N_1351,N_1250,N_1270);
nand U1352 (N_1352,N_1245,N_1265);
and U1353 (N_1353,N_1266,N_1257);
nor U1354 (N_1354,N_1282,N_1252);
nor U1355 (N_1355,N_1253,N_1257);
or U1356 (N_1356,N_1236,N_1267);
nor U1357 (N_1357,N_1268,N_1203);
or U1358 (N_1358,N_1251,N_1212);
or U1359 (N_1359,N_1256,N_1229);
or U1360 (N_1360,N_1246,N_1228);
and U1361 (N_1361,N_1261,N_1299);
or U1362 (N_1362,N_1232,N_1231);
or U1363 (N_1363,N_1260,N_1212);
nand U1364 (N_1364,N_1235,N_1287);
or U1365 (N_1365,N_1270,N_1256);
and U1366 (N_1366,N_1226,N_1227);
or U1367 (N_1367,N_1250,N_1261);
nor U1368 (N_1368,N_1227,N_1233);
nor U1369 (N_1369,N_1276,N_1203);
and U1370 (N_1370,N_1220,N_1221);
nor U1371 (N_1371,N_1238,N_1260);
nand U1372 (N_1372,N_1295,N_1262);
xnor U1373 (N_1373,N_1245,N_1205);
nand U1374 (N_1374,N_1241,N_1236);
nand U1375 (N_1375,N_1273,N_1233);
nand U1376 (N_1376,N_1237,N_1282);
nor U1377 (N_1377,N_1242,N_1258);
nor U1378 (N_1378,N_1212,N_1274);
nor U1379 (N_1379,N_1217,N_1221);
or U1380 (N_1380,N_1252,N_1258);
nand U1381 (N_1381,N_1205,N_1231);
nand U1382 (N_1382,N_1238,N_1297);
or U1383 (N_1383,N_1217,N_1202);
nor U1384 (N_1384,N_1252,N_1279);
and U1385 (N_1385,N_1268,N_1290);
and U1386 (N_1386,N_1265,N_1240);
nand U1387 (N_1387,N_1277,N_1249);
nand U1388 (N_1388,N_1230,N_1237);
or U1389 (N_1389,N_1206,N_1213);
nor U1390 (N_1390,N_1204,N_1220);
nor U1391 (N_1391,N_1269,N_1277);
and U1392 (N_1392,N_1252,N_1210);
nor U1393 (N_1393,N_1294,N_1218);
or U1394 (N_1394,N_1206,N_1280);
nor U1395 (N_1395,N_1248,N_1295);
and U1396 (N_1396,N_1205,N_1278);
or U1397 (N_1397,N_1295,N_1276);
or U1398 (N_1398,N_1275,N_1262);
nand U1399 (N_1399,N_1290,N_1266);
and U1400 (N_1400,N_1379,N_1374);
nand U1401 (N_1401,N_1331,N_1322);
and U1402 (N_1402,N_1300,N_1361);
nor U1403 (N_1403,N_1378,N_1317);
nor U1404 (N_1404,N_1351,N_1316);
nor U1405 (N_1405,N_1373,N_1313);
and U1406 (N_1406,N_1308,N_1346);
and U1407 (N_1407,N_1339,N_1325);
or U1408 (N_1408,N_1329,N_1356);
nor U1409 (N_1409,N_1323,N_1350);
and U1410 (N_1410,N_1375,N_1341);
or U1411 (N_1411,N_1337,N_1310);
nor U1412 (N_1412,N_1368,N_1314);
and U1413 (N_1413,N_1319,N_1393);
nand U1414 (N_1414,N_1396,N_1394);
or U1415 (N_1415,N_1342,N_1388);
and U1416 (N_1416,N_1301,N_1391);
or U1417 (N_1417,N_1304,N_1364);
and U1418 (N_1418,N_1399,N_1303);
and U1419 (N_1419,N_1354,N_1335);
and U1420 (N_1420,N_1305,N_1359);
nand U1421 (N_1421,N_1328,N_1372);
and U1422 (N_1422,N_1309,N_1343);
nand U1423 (N_1423,N_1380,N_1307);
nor U1424 (N_1424,N_1383,N_1320);
or U1425 (N_1425,N_1390,N_1384);
nor U1426 (N_1426,N_1367,N_1371);
nor U1427 (N_1427,N_1348,N_1397);
nand U1428 (N_1428,N_1336,N_1381);
or U1429 (N_1429,N_1318,N_1353);
nor U1430 (N_1430,N_1306,N_1355);
nor U1431 (N_1431,N_1334,N_1330);
nor U1432 (N_1432,N_1311,N_1338);
nand U1433 (N_1433,N_1370,N_1344);
nor U1434 (N_1434,N_1363,N_1321);
nor U1435 (N_1435,N_1340,N_1365);
or U1436 (N_1436,N_1362,N_1333);
or U1437 (N_1437,N_1315,N_1398);
nand U1438 (N_1438,N_1395,N_1358);
nor U1439 (N_1439,N_1357,N_1327);
or U1440 (N_1440,N_1376,N_1326);
nor U1441 (N_1441,N_1332,N_1386);
and U1442 (N_1442,N_1377,N_1352);
nand U1443 (N_1443,N_1345,N_1385);
nand U1444 (N_1444,N_1389,N_1382);
nand U1445 (N_1445,N_1347,N_1387);
or U1446 (N_1446,N_1312,N_1324);
or U1447 (N_1447,N_1366,N_1360);
or U1448 (N_1448,N_1302,N_1349);
xor U1449 (N_1449,N_1392,N_1369);
nor U1450 (N_1450,N_1336,N_1310);
or U1451 (N_1451,N_1366,N_1367);
nor U1452 (N_1452,N_1394,N_1374);
or U1453 (N_1453,N_1366,N_1323);
nor U1454 (N_1454,N_1321,N_1375);
nor U1455 (N_1455,N_1356,N_1319);
nor U1456 (N_1456,N_1302,N_1348);
nand U1457 (N_1457,N_1339,N_1397);
nor U1458 (N_1458,N_1306,N_1392);
or U1459 (N_1459,N_1382,N_1314);
nor U1460 (N_1460,N_1386,N_1372);
and U1461 (N_1461,N_1324,N_1305);
or U1462 (N_1462,N_1311,N_1360);
nor U1463 (N_1463,N_1316,N_1336);
nand U1464 (N_1464,N_1394,N_1373);
and U1465 (N_1465,N_1300,N_1389);
and U1466 (N_1466,N_1391,N_1300);
and U1467 (N_1467,N_1366,N_1306);
or U1468 (N_1468,N_1386,N_1347);
nand U1469 (N_1469,N_1346,N_1392);
nand U1470 (N_1470,N_1360,N_1333);
or U1471 (N_1471,N_1330,N_1310);
nor U1472 (N_1472,N_1381,N_1373);
or U1473 (N_1473,N_1345,N_1308);
nand U1474 (N_1474,N_1378,N_1377);
or U1475 (N_1475,N_1383,N_1385);
nor U1476 (N_1476,N_1330,N_1385);
and U1477 (N_1477,N_1304,N_1324);
nand U1478 (N_1478,N_1391,N_1373);
and U1479 (N_1479,N_1378,N_1353);
or U1480 (N_1480,N_1360,N_1389);
nor U1481 (N_1481,N_1397,N_1307);
or U1482 (N_1482,N_1398,N_1305);
or U1483 (N_1483,N_1351,N_1341);
nand U1484 (N_1484,N_1301,N_1378);
nor U1485 (N_1485,N_1352,N_1337);
and U1486 (N_1486,N_1383,N_1367);
nor U1487 (N_1487,N_1352,N_1304);
nand U1488 (N_1488,N_1300,N_1353);
nand U1489 (N_1489,N_1359,N_1397);
and U1490 (N_1490,N_1303,N_1332);
nand U1491 (N_1491,N_1336,N_1313);
or U1492 (N_1492,N_1330,N_1396);
nor U1493 (N_1493,N_1300,N_1324);
and U1494 (N_1494,N_1317,N_1380);
nand U1495 (N_1495,N_1377,N_1391);
and U1496 (N_1496,N_1393,N_1385);
nor U1497 (N_1497,N_1337,N_1331);
or U1498 (N_1498,N_1331,N_1338);
xnor U1499 (N_1499,N_1329,N_1308);
nand U1500 (N_1500,N_1461,N_1428);
nand U1501 (N_1501,N_1412,N_1401);
nand U1502 (N_1502,N_1487,N_1469);
and U1503 (N_1503,N_1402,N_1476);
nor U1504 (N_1504,N_1411,N_1429);
and U1505 (N_1505,N_1414,N_1456);
nor U1506 (N_1506,N_1408,N_1409);
or U1507 (N_1507,N_1484,N_1403);
nor U1508 (N_1508,N_1478,N_1448);
nor U1509 (N_1509,N_1489,N_1458);
or U1510 (N_1510,N_1445,N_1496);
and U1511 (N_1511,N_1497,N_1453);
or U1512 (N_1512,N_1450,N_1452);
and U1513 (N_1513,N_1420,N_1463);
or U1514 (N_1514,N_1439,N_1494);
nor U1515 (N_1515,N_1400,N_1483);
nor U1516 (N_1516,N_1443,N_1437);
xor U1517 (N_1517,N_1423,N_1466);
and U1518 (N_1518,N_1471,N_1481);
and U1519 (N_1519,N_1405,N_1488);
and U1520 (N_1520,N_1460,N_1413);
nand U1521 (N_1521,N_1486,N_1422);
and U1522 (N_1522,N_1457,N_1465);
nor U1523 (N_1523,N_1472,N_1490);
nor U1524 (N_1524,N_1426,N_1467);
nand U1525 (N_1525,N_1444,N_1455);
and U1526 (N_1526,N_1431,N_1415);
nand U1527 (N_1527,N_1482,N_1477);
or U1528 (N_1528,N_1462,N_1464);
and U1529 (N_1529,N_1427,N_1418);
nor U1530 (N_1530,N_1434,N_1449);
and U1531 (N_1531,N_1492,N_1485);
and U1532 (N_1532,N_1410,N_1451);
nand U1533 (N_1533,N_1407,N_1454);
and U1534 (N_1534,N_1480,N_1425);
nor U1535 (N_1535,N_1470,N_1491);
nand U1536 (N_1536,N_1417,N_1424);
nand U1537 (N_1537,N_1493,N_1499);
nand U1538 (N_1538,N_1430,N_1432);
and U1539 (N_1539,N_1441,N_1438);
nand U1540 (N_1540,N_1479,N_1419);
nor U1541 (N_1541,N_1421,N_1433);
nor U1542 (N_1542,N_1468,N_1416);
nor U1543 (N_1543,N_1406,N_1442);
or U1544 (N_1544,N_1447,N_1495);
or U1545 (N_1545,N_1446,N_1498);
nor U1546 (N_1546,N_1435,N_1473);
nand U1547 (N_1547,N_1459,N_1475);
nor U1548 (N_1548,N_1404,N_1440);
nand U1549 (N_1549,N_1436,N_1474);
nor U1550 (N_1550,N_1416,N_1444);
and U1551 (N_1551,N_1449,N_1457);
or U1552 (N_1552,N_1498,N_1495);
nand U1553 (N_1553,N_1431,N_1495);
or U1554 (N_1554,N_1485,N_1406);
or U1555 (N_1555,N_1428,N_1412);
or U1556 (N_1556,N_1460,N_1483);
nor U1557 (N_1557,N_1495,N_1485);
nand U1558 (N_1558,N_1457,N_1466);
nand U1559 (N_1559,N_1471,N_1426);
or U1560 (N_1560,N_1472,N_1480);
or U1561 (N_1561,N_1448,N_1454);
or U1562 (N_1562,N_1466,N_1437);
and U1563 (N_1563,N_1453,N_1419);
or U1564 (N_1564,N_1405,N_1469);
nand U1565 (N_1565,N_1460,N_1419);
nor U1566 (N_1566,N_1458,N_1424);
and U1567 (N_1567,N_1400,N_1438);
nor U1568 (N_1568,N_1478,N_1459);
nor U1569 (N_1569,N_1410,N_1486);
or U1570 (N_1570,N_1418,N_1444);
or U1571 (N_1571,N_1498,N_1499);
or U1572 (N_1572,N_1451,N_1453);
nor U1573 (N_1573,N_1409,N_1461);
xor U1574 (N_1574,N_1458,N_1423);
and U1575 (N_1575,N_1459,N_1463);
nor U1576 (N_1576,N_1416,N_1446);
nor U1577 (N_1577,N_1420,N_1478);
nand U1578 (N_1578,N_1449,N_1485);
xnor U1579 (N_1579,N_1469,N_1424);
nand U1580 (N_1580,N_1469,N_1429);
nor U1581 (N_1581,N_1486,N_1419);
and U1582 (N_1582,N_1472,N_1494);
and U1583 (N_1583,N_1436,N_1464);
or U1584 (N_1584,N_1443,N_1469);
nand U1585 (N_1585,N_1420,N_1450);
nor U1586 (N_1586,N_1427,N_1409);
and U1587 (N_1587,N_1429,N_1474);
nor U1588 (N_1588,N_1490,N_1456);
nor U1589 (N_1589,N_1491,N_1425);
nand U1590 (N_1590,N_1416,N_1438);
nor U1591 (N_1591,N_1483,N_1455);
nor U1592 (N_1592,N_1476,N_1449);
nand U1593 (N_1593,N_1458,N_1466);
nand U1594 (N_1594,N_1413,N_1431);
and U1595 (N_1595,N_1466,N_1445);
or U1596 (N_1596,N_1447,N_1428);
or U1597 (N_1597,N_1496,N_1495);
or U1598 (N_1598,N_1403,N_1485);
nor U1599 (N_1599,N_1410,N_1467);
nor U1600 (N_1600,N_1550,N_1596);
or U1601 (N_1601,N_1549,N_1580);
and U1602 (N_1602,N_1540,N_1534);
or U1603 (N_1603,N_1555,N_1538);
or U1604 (N_1604,N_1583,N_1515);
nor U1605 (N_1605,N_1514,N_1537);
or U1606 (N_1606,N_1510,N_1572);
nand U1607 (N_1607,N_1501,N_1552);
and U1608 (N_1608,N_1599,N_1513);
or U1609 (N_1609,N_1560,N_1563);
or U1610 (N_1610,N_1575,N_1532);
and U1611 (N_1611,N_1511,N_1567);
nand U1612 (N_1612,N_1526,N_1598);
or U1613 (N_1613,N_1566,N_1521);
and U1614 (N_1614,N_1504,N_1557);
nor U1615 (N_1615,N_1548,N_1582);
nand U1616 (N_1616,N_1553,N_1561);
nor U1617 (N_1617,N_1571,N_1525);
and U1618 (N_1618,N_1542,N_1589);
nand U1619 (N_1619,N_1528,N_1573);
nor U1620 (N_1620,N_1520,N_1586);
nand U1621 (N_1621,N_1595,N_1541);
or U1622 (N_1622,N_1591,N_1543);
and U1623 (N_1623,N_1593,N_1590);
nor U1624 (N_1624,N_1529,N_1564);
nor U1625 (N_1625,N_1544,N_1558);
nor U1626 (N_1626,N_1594,N_1502);
nand U1627 (N_1627,N_1505,N_1556);
and U1628 (N_1628,N_1577,N_1587);
or U1629 (N_1629,N_1546,N_1574);
or U1630 (N_1630,N_1506,N_1539);
or U1631 (N_1631,N_1535,N_1584);
or U1632 (N_1632,N_1518,N_1547);
and U1633 (N_1633,N_1576,N_1516);
nand U1634 (N_1634,N_1570,N_1530);
nand U1635 (N_1635,N_1517,N_1579);
nand U1636 (N_1636,N_1527,N_1585);
xor U1637 (N_1637,N_1508,N_1562);
and U1638 (N_1638,N_1512,N_1588);
nor U1639 (N_1639,N_1509,N_1592);
nand U1640 (N_1640,N_1545,N_1500);
or U1641 (N_1641,N_1568,N_1559);
or U1642 (N_1642,N_1524,N_1554);
nand U1643 (N_1643,N_1503,N_1581);
nor U1644 (N_1644,N_1531,N_1565);
nor U1645 (N_1645,N_1533,N_1536);
nand U1646 (N_1646,N_1519,N_1578);
and U1647 (N_1647,N_1522,N_1507);
and U1648 (N_1648,N_1551,N_1597);
and U1649 (N_1649,N_1569,N_1523);
nor U1650 (N_1650,N_1573,N_1530);
and U1651 (N_1651,N_1573,N_1538);
nand U1652 (N_1652,N_1539,N_1561);
nor U1653 (N_1653,N_1542,N_1518);
nor U1654 (N_1654,N_1509,N_1591);
nand U1655 (N_1655,N_1515,N_1577);
or U1656 (N_1656,N_1583,N_1517);
nor U1657 (N_1657,N_1571,N_1579);
nand U1658 (N_1658,N_1565,N_1593);
or U1659 (N_1659,N_1569,N_1591);
or U1660 (N_1660,N_1576,N_1550);
and U1661 (N_1661,N_1551,N_1579);
and U1662 (N_1662,N_1515,N_1548);
nand U1663 (N_1663,N_1507,N_1584);
nand U1664 (N_1664,N_1537,N_1527);
or U1665 (N_1665,N_1527,N_1595);
or U1666 (N_1666,N_1544,N_1561);
or U1667 (N_1667,N_1589,N_1586);
and U1668 (N_1668,N_1599,N_1541);
nor U1669 (N_1669,N_1500,N_1567);
nand U1670 (N_1670,N_1598,N_1585);
or U1671 (N_1671,N_1523,N_1530);
nor U1672 (N_1672,N_1556,N_1524);
nor U1673 (N_1673,N_1508,N_1516);
nand U1674 (N_1674,N_1597,N_1539);
nand U1675 (N_1675,N_1553,N_1525);
or U1676 (N_1676,N_1536,N_1557);
nand U1677 (N_1677,N_1547,N_1535);
nor U1678 (N_1678,N_1577,N_1576);
nor U1679 (N_1679,N_1518,N_1520);
nand U1680 (N_1680,N_1514,N_1505);
or U1681 (N_1681,N_1581,N_1572);
nand U1682 (N_1682,N_1560,N_1545);
and U1683 (N_1683,N_1519,N_1521);
nand U1684 (N_1684,N_1590,N_1536);
nand U1685 (N_1685,N_1517,N_1540);
nor U1686 (N_1686,N_1569,N_1549);
nor U1687 (N_1687,N_1548,N_1506);
nor U1688 (N_1688,N_1586,N_1532);
xnor U1689 (N_1689,N_1508,N_1502);
and U1690 (N_1690,N_1539,N_1599);
nor U1691 (N_1691,N_1512,N_1550);
and U1692 (N_1692,N_1515,N_1524);
nand U1693 (N_1693,N_1527,N_1522);
or U1694 (N_1694,N_1549,N_1529);
or U1695 (N_1695,N_1536,N_1519);
nor U1696 (N_1696,N_1513,N_1590);
and U1697 (N_1697,N_1581,N_1589);
nand U1698 (N_1698,N_1543,N_1563);
nand U1699 (N_1699,N_1542,N_1528);
and U1700 (N_1700,N_1609,N_1675);
nand U1701 (N_1701,N_1630,N_1623);
and U1702 (N_1702,N_1677,N_1681);
or U1703 (N_1703,N_1625,N_1617);
or U1704 (N_1704,N_1668,N_1671);
or U1705 (N_1705,N_1611,N_1624);
nor U1706 (N_1706,N_1697,N_1621);
nor U1707 (N_1707,N_1688,N_1615);
nor U1708 (N_1708,N_1620,N_1608);
and U1709 (N_1709,N_1629,N_1633);
xnor U1710 (N_1710,N_1626,N_1646);
and U1711 (N_1711,N_1665,N_1622);
or U1712 (N_1712,N_1647,N_1662);
nand U1713 (N_1713,N_1654,N_1627);
nand U1714 (N_1714,N_1696,N_1616);
and U1715 (N_1715,N_1689,N_1699);
and U1716 (N_1716,N_1602,N_1640);
nor U1717 (N_1717,N_1672,N_1601);
xor U1718 (N_1718,N_1658,N_1604);
nor U1719 (N_1719,N_1692,N_1632);
nor U1720 (N_1720,N_1679,N_1638);
or U1721 (N_1721,N_1631,N_1637);
nor U1722 (N_1722,N_1648,N_1683);
nor U1723 (N_1723,N_1669,N_1642);
or U1724 (N_1724,N_1603,N_1659);
nor U1725 (N_1725,N_1694,N_1641);
and U1726 (N_1726,N_1612,N_1639);
or U1727 (N_1727,N_1684,N_1693);
or U1728 (N_1728,N_1605,N_1698);
and U1729 (N_1729,N_1643,N_1655);
and U1730 (N_1730,N_1663,N_1682);
nand U1731 (N_1731,N_1687,N_1686);
nor U1732 (N_1732,N_1667,N_1656);
and U1733 (N_1733,N_1628,N_1664);
and U1734 (N_1734,N_1606,N_1690);
and U1735 (N_1735,N_1652,N_1614);
nand U1736 (N_1736,N_1651,N_1695);
nand U1737 (N_1737,N_1645,N_1661);
and U1738 (N_1738,N_1678,N_1649);
and U1739 (N_1739,N_1670,N_1636);
or U1740 (N_1740,N_1644,N_1657);
or U1741 (N_1741,N_1635,N_1610);
nor U1742 (N_1742,N_1673,N_1680);
and U1743 (N_1743,N_1618,N_1600);
nand U1744 (N_1744,N_1607,N_1674);
nor U1745 (N_1745,N_1653,N_1650);
nor U1746 (N_1746,N_1691,N_1676);
or U1747 (N_1747,N_1660,N_1613);
and U1748 (N_1748,N_1619,N_1634);
nand U1749 (N_1749,N_1666,N_1685);
nand U1750 (N_1750,N_1646,N_1632);
nand U1751 (N_1751,N_1634,N_1699);
or U1752 (N_1752,N_1688,N_1682);
and U1753 (N_1753,N_1667,N_1691);
nor U1754 (N_1754,N_1662,N_1617);
nor U1755 (N_1755,N_1609,N_1690);
or U1756 (N_1756,N_1606,N_1682);
nand U1757 (N_1757,N_1673,N_1646);
nand U1758 (N_1758,N_1642,N_1607);
nor U1759 (N_1759,N_1630,N_1603);
or U1760 (N_1760,N_1668,N_1694);
and U1761 (N_1761,N_1616,N_1604);
nand U1762 (N_1762,N_1664,N_1606);
and U1763 (N_1763,N_1652,N_1684);
nor U1764 (N_1764,N_1607,N_1688);
nand U1765 (N_1765,N_1668,N_1626);
nor U1766 (N_1766,N_1665,N_1654);
and U1767 (N_1767,N_1605,N_1660);
and U1768 (N_1768,N_1640,N_1658);
nand U1769 (N_1769,N_1612,N_1641);
or U1770 (N_1770,N_1641,N_1660);
nand U1771 (N_1771,N_1622,N_1661);
nor U1772 (N_1772,N_1687,N_1688);
or U1773 (N_1773,N_1638,N_1613);
and U1774 (N_1774,N_1657,N_1666);
and U1775 (N_1775,N_1691,N_1633);
nand U1776 (N_1776,N_1688,N_1696);
or U1777 (N_1777,N_1663,N_1655);
nor U1778 (N_1778,N_1665,N_1650);
nor U1779 (N_1779,N_1600,N_1659);
and U1780 (N_1780,N_1652,N_1632);
or U1781 (N_1781,N_1654,N_1637);
and U1782 (N_1782,N_1617,N_1639);
and U1783 (N_1783,N_1622,N_1662);
or U1784 (N_1784,N_1642,N_1647);
nand U1785 (N_1785,N_1688,N_1617);
nand U1786 (N_1786,N_1632,N_1621);
nor U1787 (N_1787,N_1638,N_1607);
and U1788 (N_1788,N_1668,N_1659);
or U1789 (N_1789,N_1619,N_1694);
and U1790 (N_1790,N_1693,N_1685);
nor U1791 (N_1791,N_1647,N_1608);
nor U1792 (N_1792,N_1670,N_1669);
nor U1793 (N_1793,N_1657,N_1658);
nor U1794 (N_1794,N_1699,N_1604);
and U1795 (N_1795,N_1624,N_1685);
nand U1796 (N_1796,N_1617,N_1668);
or U1797 (N_1797,N_1663,N_1674);
and U1798 (N_1798,N_1624,N_1634);
nand U1799 (N_1799,N_1675,N_1604);
and U1800 (N_1800,N_1710,N_1730);
and U1801 (N_1801,N_1760,N_1719);
nor U1802 (N_1802,N_1749,N_1791);
and U1803 (N_1803,N_1729,N_1778);
nand U1804 (N_1804,N_1787,N_1705);
nor U1805 (N_1805,N_1736,N_1789);
nor U1806 (N_1806,N_1738,N_1781);
or U1807 (N_1807,N_1782,N_1739);
and U1808 (N_1808,N_1776,N_1771);
and U1809 (N_1809,N_1766,N_1725);
and U1810 (N_1810,N_1751,N_1709);
xnor U1811 (N_1811,N_1775,N_1727);
nor U1812 (N_1812,N_1741,N_1745);
nand U1813 (N_1813,N_1770,N_1703);
and U1814 (N_1814,N_1732,N_1790);
nand U1815 (N_1815,N_1777,N_1714);
nand U1816 (N_1816,N_1759,N_1702);
xor U1817 (N_1817,N_1708,N_1720);
nand U1818 (N_1818,N_1704,N_1793);
and U1819 (N_1819,N_1780,N_1728);
or U1820 (N_1820,N_1752,N_1740);
or U1821 (N_1821,N_1707,N_1765);
and U1822 (N_1822,N_1769,N_1796);
or U1823 (N_1823,N_1735,N_1717);
nand U1824 (N_1824,N_1737,N_1700);
or U1825 (N_1825,N_1755,N_1754);
or U1826 (N_1826,N_1774,N_1773);
nor U1827 (N_1827,N_1706,N_1750);
nand U1828 (N_1828,N_1762,N_1767);
or U1829 (N_1829,N_1742,N_1733);
nor U1830 (N_1830,N_1763,N_1747);
nor U1831 (N_1831,N_1764,N_1713);
and U1832 (N_1832,N_1779,N_1743);
or U1833 (N_1833,N_1726,N_1731);
and U1834 (N_1834,N_1753,N_1711);
nor U1835 (N_1835,N_1786,N_1721);
and U1836 (N_1836,N_1792,N_1744);
and U1837 (N_1837,N_1718,N_1798);
and U1838 (N_1838,N_1722,N_1756);
nor U1839 (N_1839,N_1783,N_1757);
nor U1840 (N_1840,N_1785,N_1724);
nor U1841 (N_1841,N_1784,N_1758);
nand U1842 (N_1842,N_1748,N_1795);
or U1843 (N_1843,N_1799,N_1746);
nor U1844 (N_1844,N_1715,N_1761);
nand U1845 (N_1845,N_1716,N_1734);
and U1846 (N_1846,N_1768,N_1712);
nor U1847 (N_1847,N_1701,N_1723);
nand U1848 (N_1848,N_1794,N_1772);
or U1849 (N_1849,N_1788,N_1797);
nand U1850 (N_1850,N_1766,N_1734);
and U1851 (N_1851,N_1760,N_1728);
or U1852 (N_1852,N_1766,N_1754);
nor U1853 (N_1853,N_1746,N_1745);
or U1854 (N_1854,N_1756,N_1753);
nand U1855 (N_1855,N_1722,N_1772);
and U1856 (N_1856,N_1731,N_1765);
nor U1857 (N_1857,N_1795,N_1777);
or U1858 (N_1858,N_1792,N_1726);
nor U1859 (N_1859,N_1712,N_1731);
and U1860 (N_1860,N_1765,N_1794);
nand U1861 (N_1861,N_1741,N_1725);
or U1862 (N_1862,N_1788,N_1766);
nor U1863 (N_1863,N_1757,N_1767);
nor U1864 (N_1864,N_1755,N_1756);
nand U1865 (N_1865,N_1703,N_1789);
and U1866 (N_1866,N_1724,N_1766);
and U1867 (N_1867,N_1758,N_1708);
or U1868 (N_1868,N_1787,N_1796);
and U1869 (N_1869,N_1772,N_1756);
and U1870 (N_1870,N_1770,N_1750);
nand U1871 (N_1871,N_1775,N_1743);
or U1872 (N_1872,N_1773,N_1708);
nor U1873 (N_1873,N_1782,N_1738);
or U1874 (N_1874,N_1752,N_1729);
and U1875 (N_1875,N_1738,N_1731);
or U1876 (N_1876,N_1716,N_1711);
or U1877 (N_1877,N_1752,N_1719);
and U1878 (N_1878,N_1700,N_1780);
nor U1879 (N_1879,N_1703,N_1718);
nor U1880 (N_1880,N_1774,N_1771);
and U1881 (N_1881,N_1773,N_1742);
nand U1882 (N_1882,N_1719,N_1747);
xnor U1883 (N_1883,N_1714,N_1751);
nor U1884 (N_1884,N_1772,N_1788);
or U1885 (N_1885,N_1708,N_1709);
and U1886 (N_1886,N_1732,N_1713);
nor U1887 (N_1887,N_1705,N_1759);
and U1888 (N_1888,N_1729,N_1735);
nor U1889 (N_1889,N_1788,N_1781);
or U1890 (N_1890,N_1730,N_1739);
or U1891 (N_1891,N_1705,N_1712);
or U1892 (N_1892,N_1727,N_1778);
and U1893 (N_1893,N_1717,N_1741);
nor U1894 (N_1894,N_1782,N_1769);
or U1895 (N_1895,N_1789,N_1790);
nand U1896 (N_1896,N_1729,N_1727);
and U1897 (N_1897,N_1784,N_1770);
and U1898 (N_1898,N_1752,N_1784);
nor U1899 (N_1899,N_1773,N_1772);
or U1900 (N_1900,N_1829,N_1827);
or U1901 (N_1901,N_1845,N_1857);
or U1902 (N_1902,N_1805,N_1814);
nand U1903 (N_1903,N_1819,N_1820);
or U1904 (N_1904,N_1850,N_1824);
and U1905 (N_1905,N_1872,N_1866);
nor U1906 (N_1906,N_1854,N_1856);
and U1907 (N_1907,N_1852,N_1861);
and U1908 (N_1908,N_1892,N_1878);
and U1909 (N_1909,N_1891,N_1858);
nand U1910 (N_1910,N_1860,N_1868);
or U1911 (N_1911,N_1843,N_1801);
nor U1912 (N_1912,N_1890,N_1882);
nand U1913 (N_1913,N_1823,N_1804);
nand U1914 (N_1914,N_1886,N_1867);
and U1915 (N_1915,N_1803,N_1870);
nand U1916 (N_1916,N_1825,N_1822);
and U1917 (N_1917,N_1836,N_1821);
nand U1918 (N_1918,N_1853,N_1888);
nand U1919 (N_1919,N_1842,N_1806);
and U1920 (N_1920,N_1848,N_1818);
nand U1921 (N_1921,N_1826,N_1887);
and U1922 (N_1922,N_1830,N_1844);
and U1923 (N_1923,N_1883,N_1884);
nand U1924 (N_1924,N_1809,N_1881);
or U1925 (N_1925,N_1817,N_1834);
or U1926 (N_1926,N_1873,N_1895);
and U1927 (N_1927,N_1847,N_1835);
nor U1928 (N_1928,N_1889,N_1816);
nand U1929 (N_1929,N_1810,N_1871);
nor U1930 (N_1930,N_1837,N_1896);
nor U1931 (N_1931,N_1812,N_1863);
nor U1932 (N_1932,N_1808,N_1869);
and U1933 (N_1933,N_1862,N_1899);
and U1934 (N_1934,N_1838,N_1865);
nand U1935 (N_1935,N_1841,N_1879);
nand U1936 (N_1936,N_1864,N_1874);
and U1937 (N_1937,N_1840,N_1893);
nor U1938 (N_1938,N_1849,N_1839);
or U1939 (N_1939,N_1898,N_1828);
nand U1940 (N_1940,N_1876,N_1855);
and U1941 (N_1941,N_1813,N_1802);
nor U1942 (N_1942,N_1880,N_1859);
nor U1943 (N_1943,N_1800,N_1811);
nor U1944 (N_1944,N_1807,N_1877);
nor U1945 (N_1945,N_1851,N_1846);
or U1946 (N_1946,N_1894,N_1831);
and U1947 (N_1947,N_1815,N_1885);
and U1948 (N_1948,N_1875,N_1897);
or U1949 (N_1949,N_1832,N_1833);
and U1950 (N_1950,N_1833,N_1871);
xnor U1951 (N_1951,N_1860,N_1879);
and U1952 (N_1952,N_1897,N_1826);
nor U1953 (N_1953,N_1820,N_1878);
and U1954 (N_1954,N_1817,N_1828);
and U1955 (N_1955,N_1842,N_1813);
or U1956 (N_1956,N_1828,N_1879);
nor U1957 (N_1957,N_1889,N_1879);
and U1958 (N_1958,N_1828,N_1836);
and U1959 (N_1959,N_1896,N_1806);
and U1960 (N_1960,N_1895,N_1845);
or U1961 (N_1961,N_1869,N_1889);
nor U1962 (N_1962,N_1898,N_1823);
nor U1963 (N_1963,N_1854,N_1824);
and U1964 (N_1964,N_1894,N_1816);
or U1965 (N_1965,N_1820,N_1842);
nand U1966 (N_1966,N_1891,N_1880);
and U1967 (N_1967,N_1838,N_1889);
nor U1968 (N_1968,N_1864,N_1838);
or U1969 (N_1969,N_1813,N_1863);
or U1970 (N_1970,N_1817,N_1808);
nor U1971 (N_1971,N_1865,N_1836);
nor U1972 (N_1972,N_1822,N_1872);
nand U1973 (N_1973,N_1864,N_1882);
nand U1974 (N_1974,N_1885,N_1850);
and U1975 (N_1975,N_1842,N_1852);
nor U1976 (N_1976,N_1825,N_1891);
or U1977 (N_1977,N_1832,N_1829);
nor U1978 (N_1978,N_1897,N_1822);
nor U1979 (N_1979,N_1823,N_1840);
and U1980 (N_1980,N_1811,N_1866);
and U1981 (N_1981,N_1884,N_1825);
or U1982 (N_1982,N_1844,N_1869);
nand U1983 (N_1983,N_1824,N_1866);
or U1984 (N_1984,N_1892,N_1842);
nand U1985 (N_1985,N_1835,N_1814);
or U1986 (N_1986,N_1878,N_1810);
or U1987 (N_1987,N_1896,N_1854);
xnor U1988 (N_1988,N_1899,N_1898);
and U1989 (N_1989,N_1882,N_1887);
nand U1990 (N_1990,N_1898,N_1863);
and U1991 (N_1991,N_1829,N_1815);
nor U1992 (N_1992,N_1824,N_1811);
or U1993 (N_1993,N_1805,N_1827);
nand U1994 (N_1994,N_1846,N_1828);
or U1995 (N_1995,N_1804,N_1839);
nor U1996 (N_1996,N_1879,N_1853);
or U1997 (N_1997,N_1820,N_1838);
nor U1998 (N_1998,N_1839,N_1882);
or U1999 (N_1999,N_1815,N_1844);
nand U2000 (N_2000,N_1996,N_1970);
nand U2001 (N_2001,N_1900,N_1993);
nor U2002 (N_2002,N_1992,N_1951);
nand U2003 (N_2003,N_1958,N_1979);
nor U2004 (N_2004,N_1916,N_1976);
nor U2005 (N_2005,N_1918,N_1981);
nor U2006 (N_2006,N_1917,N_1956);
nand U2007 (N_2007,N_1931,N_1909);
nor U2008 (N_2008,N_1967,N_1945);
nand U2009 (N_2009,N_1930,N_1952);
or U2010 (N_2010,N_1986,N_1925);
or U2011 (N_2011,N_1995,N_1936);
nor U2012 (N_2012,N_1974,N_1908);
nor U2013 (N_2013,N_1988,N_1962);
nand U2014 (N_2014,N_1933,N_1934);
xnor U2015 (N_2015,N_1968,N_1921);
and U2016 (N_2016,N_1999,N_1928);
nand U2017 (N_2017,N_1957,N_1901);
nor U2018 (N_2018,N_1926,N_1991);
nor U2019 (N_2019,N_1915,N_1914);
or U2020 (N_2020,N_1903,N_1905);
nand U2021 (N_2021,N_1940,N_1972);
nor U2022 (N_2022,N_1997,N_1947);
and U2023 (N_2023,N_1938,N_1963);
and U2024 (N_2024,N_1971,N_1929);
nor U2025 (N_2025,N_1907,N_1944);
nand U2026 (N_2026,N_1982,N_1987);
nor U2027 (N_2027,N_1932,N_1911);
nand U2028 (N_2028,N_1984,N_1959);
nand U2029 (N_2029,N_1912,N_1990);
nor U2030 (N_2030,N_1953,N_1946);
xor U2031 (N_2031,N_1980,N_1973);
nand U2032 (N_2032,N_1969,N_1948);
or U2033 (N_2033,N_1913,N_1902);
or U2034 (N_2034,N_1961,N_1965);
nor U2035 (N_2035,N_1941,N_1927);
nand U2036 (N_2036,N_1920,N_1939);
xor U2037 (N_2037,N_1922,N_1955);
or U2038 (N_2038,N_1975,N_1919);
and U2039 (N_2039,N_1949,N_1966);
nand U2040 (N_2040,N_1924,N_1937);
nand U2041 (N_2041,N_1977,N_1910);
nand U2042 (N_2042,N_1983,N_1904);
nand U2043 (N_2043,N_1989,N_1998);
nor U2044 (N_2044,N_1960,N_1942);
xnor U2045 (N_2045,N_1950,N_1906);
and U2046 (N_2046,N_1943,N_1964);
nand U2047 (N_2047,N_1985,N_1954);
or U2048 (N_2048,N_1923,N_1978);
or U2049 (N_2049,N_1994,N_1935);
and U2050 (N_2050,N_1960,N_1976);
and U2051 (N_2051,N_1995,N_1906);
nand U2052 (N_2052,N_1964,N_1930);
nand U2053 (N_2053,N_1930,N_1948);
nor U2054 (N_2054,N_1968,N_1908);
or U2055 (N_2055,N_1932,N_1981);
or U2056 (N_2056,N_1959,N_1982);
and U2057 (N_2057,N_1977,N_1903);
nand U2058 (N_2058,N_1999,N_1927);
or U2059 (N_2059,N_1981,N_1994);
and U2060 (N_2060,N_1957,N_1971);
nand U2061 (N_2061,N_1942,N_1957);
and U2062 (N_2062,N_1961,N_1968);
nor U2063 (N_2063,N_1962,N_1948);
or U2064 (N_2064,N_1913,N_1931);
xor U2065 (N_2065,N_1973,N_1952);
and U2066 (N_2066,N_1930,N_1907);
nor U2067 (N_2067,N_1918,N_1980);
nor U2068 (N_2068,N_1933,N_1902);
or U2069 (N_2069,N_1954,N_1991);
or U2070 (N_2070,N_1925,N_1937);
or U2071 (N_2071,N_1967,N_1987);
and U2072 (N_2072,N_1989,N_1947);
nand U2073 (N_2073,N_1953,N_1932);
nand U2074 (N_2074,N_1989,N_1928);
and U2075 (N_2075,N_1920,N_1963);
nand U2076 (N_2076,N_1939,N_1982);
xnor U2077 (N_2077,N_1991,N_1949);
or U2078 (N_2078,N_1935,N_1986);
nand U2079 (N_2079,N_1921,N_1998);
nor U2080 (N_2080,N_1971,N_1998);
or U2081 (N_2081,N_1960,N_1930);
nor U2082 (N_2082,N_1956,N_1934);
nor U2083 (N_2083,N_1960,N_1966);
and U2084 (N_2084,N_1902,N_1993);
nand U2085 (N_2085,N_1922,N_1954);
nand U2086 (N_2086,N_1997,N_1903);
nand U2087 (N_2087,N_1983,N_1944);
and U2088 (N_2088,N_1918,N_1998);
nor U2089 (N_2089,N_1978,N_1982);
or U2090 (N_2090,N_1902,N_1909);
nor U2091 (N_2091,N_1962,N_1944);
and U2092 (N_2092,N_1935,N_1924);
nor U2093 (N_2093,N_1971,N_1991);
nor U2094 (N_2094,N_1943,N_1979);
nand U2095 (N_2095,N_1978,N_1950);
and U2096 (N_2096,N_1938,N_1968);
or U2097 (N_2097,N_1987,N_1979);
nand U2098 (N_2098,N_1943,N_1997);
or U2099 (N_2099,N_1958,N_1987);
or U2100 (N_2100,N_2092,N_2073);
nand U2101 (N_2101,N_2010,N_2008);
xor U2102 (N_2102,N_2090,N_2005);
and U2103 (N_2103,N_2039,N_2011);
and U2104 (N_2104,N_2002,N_2044);
or U2105 (N_2105,N_2022,N_2007);
or U2106 (N_2106,N_2009,N_2013);
xor U2107 (N_2107,N_2042,N_2041);
nand U2108 (N_2108,N_2015,N_2074);
nand U2109 (N_2109,N_2001,N_2077);
or U2110 (N_2110,N_2049,N_2069);
or U2111 (N_2111,N_2060,N_2068);
or U2112 (N_2112,N_2051,N_2081);
nor U2113 (N_2113,N_2033,N_2078);
nand U2114 (N_2114,N_2084,N_2083);
and U2115 (N_2115,N_2088,N_2097);
and U2116 (N_2116,N_2034,N_2093);
nor U2117 (N_2117,N_2095,N_2050);
nor U2118 (N_2118,N_2082,N_2038);
and U2119 (N_2119,N_2099,N_2059);
nand U2120 (N_2120,N_2094,N_2003);
nor U2121 (N_2121,N_2072,N_2036);
nand U2122 (N_2122,N_2058,N_2031);
nor U2123 (N_2123,N_2071,N_2062);
and U2124 (N_2124,N_2025,N_2032);
nand U2125 (N_2125,N_2021,N_2018);
nand U2126 (N_2126,N_2045,N_2080);
nand U2127 (N_2127,N_2024,N_2037);
nor U2128 (N_2128,N_2079,N_2043);
nand U2129 (N_2129,N_2035,N_2089);
or U2130 (N_2130,N_2056,N_2091);
and U2131 (N_2131,N_2014,N_2067);
or U2132 (N_2132,N_2057,N_2065);
nand U2133 (N_2133,N_2030,N_2053);
nor U2134 (N_2134,N_2004,N_2076);
or U2135 (N_2135,N_2016,N_2029);
and U2136 (N_2136,N_2040,N_2026);
nand U2137 (N_2137,N_2085,N_2012);
nor U2138 (N_2138,N_2064,N_2096);
and U2139 (N_2139,N_2098,N_2023);
and U2140 (N_2140,N_2020,N_2087);
or U2141 (N_2141,N_2046,N_2052);
and U2142 (N_2142,N_2054,N_2086);
and U2143 (N_2143,N_2006,N_2070);
and U2144 (N_2144,N_2075,N_2019);
nor U2145 (N_2145,N_2028,N_2063);
xor U2146 (N_2146,N_2027,N_2066);
nand U2147 (N_2147,N_2047,N_2048);
nand U2148 (N_2148,N_2017,N_2055);
nor U2149 (N_2149,N_2000,N_2061);
and U2150 (N_2150,N_2080,N_2079);
nor U2151 (N_2151,N_2082,N_2070);
and U2152 (N_2152,N_2039,N_2016);
nor U2153 (N_2153,N_2044,N_2033);
nor U2154 (N_2154,N_2072,N_2024);
or U2155 (N_2155,N_2008,N_2094);
or U2156 (N_2156,N_2063,N_2035);
nor U2157 (N_2157,N_2001,N_2060);
nand U2158 (N_2158,N_2096,N_2029);
nor U2159 (N_2159,N_2098,N_2046);
or U2160 (N_2160,N_2014,N_2035);
and U2161 (N_2161,N_2008,N_2011);
nand U2162 (N_2162,N_2008,N_2055);
nor U2163 (N_2163,N_2065,N_2005);
or U2164 (N_2164,N_2055,N_2015);
or U2165 (N_2165,N_2054,N_2019);
or U2166 (N_2166,N_2095,N_2025);
or U2167 (N_2167,N_2026,N_2049);
and U2168 (N_2168,N_2024,N_2031);
and U2169 (N_2169,N_2059,N_2057);
and U2170 (N_2170,N_2006,N_2004);
nand U2171 (N_2171,N_2059,N_2092);
and U2172 (N_2172,N_2022,N_2012);
nand U2173 (N_2173,N_2057,N_2094);
or U2174 (N_2174,N_2018,N_2085);
or U2175 (N_2175,N_2026,N_2047);
nand U2176 (N_2176,N_2033,N_2015);
or U2177 (N_2177,N_2077,N_2085);
or U2178 (N_2178,N_2028,N_2093);
nand U2179 (N_2179,N_2023,N_2090);
and U2180 (N_2180,N_2052,N_2017);
nor U2181 (N_2181,N_2005,N_2074);
nor U2182 (N_2182,N_2005,N_2047);
or U2183 (N_2183,N_2090,N_2038);
nor U2184 (N_2184,N_2014,N_2042);
nor U2185 (N_2185,N_2024,N_2091);
nor U2186 (N_2186,N_2036,N_2029);
nand U2187 (N_2187,N_2018,N_2074);
and U2188 (N_2188,N_2002,N_2048);
and U2189 (N_2189,N_2026,N_2051);
nand U2190 (N_2190,N_2099,N_2092);
and U2191 (N_2191,N_2020,N_2006);
or U2192 (N_2192,N_2072,N_2061);
nand U2193 (N_2193,N_2099,N_2075);
or U2194 (N_2194,N_2087,N_2082);
nand U2195 (N_2195,N_2072,N_2020);
and U2196 (N_2196,N_2098,N_2091);
nand U2197 (N_2197,N_2056,N_2017);
nand U2198 (N_2198,N_2082,N_2039);
and U2199 (N_2199,N_2045,N_2044);
nand U2200 (N_2200,N_2137,N_2145);
and U2201 (N_2201,N_2134,N_2122);
or U2202 (N_2202,N_2180,N_2150);
and U2203 (N_2203,N_2154,N_2155);
nand U2204 (N_2204,N_2172,N_2168);
nor U2205 (N_2205,N_2198,N_2162);
and U2206 (N_2206,N_2146,N_2175);
nor U2207 (N_2207,N_2114,N_2193);
and U2208 (N_2208,N_2124,N_2152);
or U2209 (N_2209,N_2121,N_2159);
nor U2210 (N_2210,N_2108,N_2165);
nor U2211 (N_2211,N_2129,N_2107);
nand U2212 (N_2212,N_2149,N_2197);
and U2213 (N_2213,N_2141,N_2139);
and U2214 (N_2214,N_2192,N_2167);
or U2215 (N_2215,N_2188,N_2183);
nand U2216 (N_2216,N_2181,N_2174);
and U2217 (N_2217,N_2195,N_2125);
and U2218 (N_2218,N_2102,N_2177);
nand U2219 (N_2219,N_2176,N_2173);
nor U2220 (N_2220,N_2190,N_2148);
nand U2221 (N_2221,N_2117,N_2113);
and U2222 (N_2222,N_2163,N_2170);
nor U2223 (N_2223,N_2158,N_2161);
nor U2224 (N_2224,N_2160,N_2106);
nor U2225 (N_2225,N_2123,N_2187);
nor U2226 (N_2226,N_2101,N_2132);
and U2227 (N_2227,N_2151,N_2110);
nor U2228 (N_2228,N_2112,N_2191);
nand U2229 (N_2229,N_2140,N_2105);
nand U2230 (N_2230,N_2189,N_2144);
nand U2231 (N_2231,N_2184,N_2127);
nand U2232 (N_2232,N_2128,N_2120);
nor U2233 (N_2233,N_2156,N_2169);
nand U2234 (N_2234,N_2131,N_2164);
or U2235 (N_2235,N_2100,N_2199);
or U2236 (N_2236,N_2194,N_2143);
and U2237 (N_2237,N_2118,N_2185);
and U2238 (N_2238,N_2111,N_2147);
or U2239 (N_2239,N_2157,N_2142);
nor U2240 (N_2240,N_2171,N_2135);
or U2241 (N_2241,N_2104,N_2136);
nor U2242 (N_2242,N_2126,N_2119);
nor U2243 (N_2243,N_2178,N_2166);
or U2244 (N_2244,N_2116,N_2153);
or U2245 (N_2245,N_2179,N_2115);
nand U2246 (N_2246,N_2130,N_2182);
and U2247 (N_2247,N_2103,N_2138);
or U2248 (N_2248,N_2186,N_2109);
nand U2249 (N_2249,N_2196,N_2133);
nor U2250 (N_2250,N_2196,N_2125);
and U2251 (N_2251,N_2122,N_2114);
or U2252 (N_2252,N_2156,N_2170);
nand U2253 (N_2253,N_2100,N_2183);
nor U2254 (N_2254,N_2146,N_2150);
nand U2255 (N_2255,N_2189,N_2126);
or U2256 (N_2256,N_2154,N_2108);
nor U2257 (N_2257,N_2173,N_2121);
nand U2258 (N_2258,N_2118,N_2129);
or U2259 (N_2259,N_2143,N_2170);
nand U2260 (N_2260,N_2161,N_2176);
and U2261 (N_2261,N_2136,N_2144);
nand U2262 (N_2262,N_2110,N_2180);
or U2263 (N_2263,N_2180,N_2172);
nand U2264 (N_2264,N_2182,N_2140);
or U2265 (N_2265,N_2194,N_2149);
and U2266 (N_2266,N_2171,N_2120);
nor U2267 (N_2267,N_2159,N_2138);
nand U2268 (N_2268,N_2118,N_2138);
nor U2269 (N_2269,N_2182,N_2147);
or U2270 (N_2270,N_2175,N_2147);
nor U2271 (N_2271,N_2141,N_2112);
or U2272 (N_2272,N_2118,N_2158);
and U2273 (N_2273,N_2113,N_2145);
and U2274 (N_2274,N_2128,N_2113);
nand U2275 (N_2275,N_2137,N_2182);
or U2276 (N_2276,N_2194,N_2129);
nand U2277 (N_2277,N_2110,N_2144);
or U2278 (N_2278,N_2164,N_2146);
nor U2279 (N_2279,N_2149,N_2164);
or U2280 (N_2280,N_2198,N_2130);
and U2281 (N_2281,N_2178,N_2182);
or U2282 (N_2282,N_2127,N_2181);
or U2283 (N_2283,N_2125,N_2114);
and U2284 (N_2284,N_2175,N_2172);
nor U2285 (N_2285,N_2107,N_2146);
and U2286 (N_2286,N_2107,N_2159);
nor U2287 (N_2287,N_2115,N_2149);
nor U2288 (N_2288,N_2112,N_2103);
nand U2289 (N_2289,N_2195,N_2162);
and U2290 (N_2290,N_2111,N_2112);
or U2291 (N_2291,N_2117,N_2128);
nand U2292 (N_2292,N_2112,N_2198);
nor U2293 (N_2293,N_2172,N_2196);
nand U2294 (N_2294,N_2126,N_2194);
and U2295 (N_2295,N_2121,N_2164);
or U2296 (N_2296,N_2100,N_2101);
and U2297 (N_2297,N_2179,N_2193);
and U2298 (N_2298,N_2173,N_2159);
and U2299 (N_2299,N_2104,N_2102);
nand U2300 (N_2300,N_2270,N_2252);
nand U2301 (N_2301,N_2235,N_2299);
and U2302 (N_2302,N_2246,N_2233);
nor U2303 (N_2303,N_2248,N_2258);
nor U2304 (N_2304,N_2204,N_2295);
nand U2305 (N_2305,N_2259,N_2228);
xnor U2306 (N_2306,N_2241,N_2226);
nor U2307 (N_2307,N_2216,N_2238);
nand U2308 (N_2308,N_2279,N_2232);
or U2309 (N_2309,N_2260,N_2280);
nand U2310 (N_2310,N_2288,N_2243);
nor U2311 (N_2311,N_2210,N_2234);
or U2312 (N_2312,N_2209,N_2206);
nor U2313 (N_2313,N_2253,N_2200);
and U2314 (N_2314,N_2278,N_2201);
nor U2315 (N_2315,N_2286,N_2267);
and U2316 (N_2316,N_2261,N_2297);
nand U2317 (N_2317,N_2285,N_2257);
nor U2318 (N_2318,N_2289,N_2237);
or U2319 (N_2319,N_2250,N_2236);
and U2320 (N_2320,N_2212,N_2249);
nand U2321 (N_2321,N_2293,N_2240);
and U2322 (N_2322,N_2298,N_2247);
and U2323 (N_2323,N_2291,N_2275);
nor U2324 (N_2324,N_2218,N_2290);
nand U2325 (N_2325,N_2273,N_2221);
nor U2326 (N_2326,N_2227,N_2203);
or U2327 (N_2327,N_2271,N_2276);
and U2328 (N_2328,N_2264,N_2224);
nor U2329 (N_2329,N_2255,N_2239);
nor U2330 (N_2330,N_2245,N_2287);
nand U2331 (N_2331,N_2283,N_2292);
or U2332 (N_2332,N_2277,N_2217);
or U2333 (N_2333,N_2208,N_2294);
nand U2334 (N_2334,N_2230,N_2220);
nand U2335 (N_2335,N_2254,N_2281);
nor U2336 (N_2336,N_2207,N_2266);
or U2337 (N_2337,N_2296,N_2213);
or U2338 (N_2338,N_2231,N_2225);
and U2339 (N_2339,N_2268,N_2215);
nand U2340 (N_2340,N_2219,N_2282);
and U2341 (N_2341,N_2251,N_2205);
or U2342 (N_2342,N_2263,N_2256);
or U2343 (N_2343,N_2214,N_2223);
or U2344 (N_2344,N_2274,N_2229);
and U2345 (N_2345,N_2269,N_2222);
or U2346 (N_2346,N_2284,N_2202);
and U2347 (N_2347,N_2244,N_2262);
nor U2348 (N_2348,N_2211,N_2242);
nand U2349 (N_2349,N_2265,N_2272);
nand U2350 (N_2350,N_2236,N_2291);
or U2351 (N_2351,N_2235,N_2293);
nand U2352 (N_2352,N_2209,N_2293);
nand U2353 (N_2353,N_2282,N_2283);
or U2354 (N_2354,N_2283,N_2231);
and U2355 (N_2355,N_2278,N_2211);
nor U2356 (N_2356,N_2268,N_2289);
nor U2357 (N_2357,N_2276,N_2218);
or U2358 (N_2358,N_2255,N_2200);
or U2359 (N_2359,N_2292,N_2299);
nand U2360 (N_2360,N_2237,N_2295);
or U2361 (N_2361,N_2228,N_2260);
nand U2362 (N_2362,N_2285,N_2274);
nor U2363 (N_2363,N_2293,N_2229);
or U2364 (N_2364,N_2255,N_2214);
nand U2365 (N_2365,N_2203,N_2201);
or U2366 (N_2366,N_2239,N_2284);
or U2367 (N_2367,N_2290,N_2226);
nand U2368 (N_2368,N_2298,N_2226);
nor U2369 (N_2369,N_2257,N_2253);
and U2370 (N_2370,N_2200,N_2266);
nor U2371 (N_2371,N_2263,N_2213);
or U2372 (N_2372,N_2281,N_2224);
or U2373 (N_2373,N_2214,N_2292);
and U2374 (N_2374,N_2227,N_2212);
nor U2375 (N_2375,N_2285,N_2273);
nand U2376 (N_2376,N_2292,N_2217);
and U2377 (N_2377,N_2217,N_2298);
or U2378 (N_2378,N_2277,N_2224);
nand U2379 (N_2379,N_2212,N_2204);
and U2380 (N_2380,N_2208,N_2262);
and U2381 (N_2381,N_2227,N_2254);
or U2382 (N_2382,N_2280,N_2261);
or U2383 (N_2383,N_2222,N_2251);
nor U2384 (N_2384,N_2281,N_2206);
or U2385 (N_2385,N_2250,N_2245);
or U2386 (N_2386,N_2214,N_2247);
or U2387 (N_2387,N_2203,N_2208);
nor U2388 (N_2388,N_2230,N_2272);
or U2389 (N_2389,N_2285,N_2256);
and U2390 (N_2390,N_2233,N_2272);
nand U2391 (N_2391,N_2240,N_2259);
nor U2392 (N_2392,N_2211,N_2258);
or U2393 (N_2393,N_2208,N_2246);
nand U2394 (N_2394,N_2251,N_2209);
or U2395 (N_2395,N_2294,N_2268);
nor U2396 (N_2396,N_2249,N_2208);
nor U2397 (N_2397,N_2261,N_2243);
or U2398 (N_2398,N_2291,N_2244);
nor U2399 (N_2399,N_2253,N_2245);
nand U2400 (N_2400,N_2337,N_2378);
nor U2401 (N_2401,N_2380,N_2318);
nand U2402 (N_2402,N_2373,N_2353);
and U2403 (N_2403,N_2398,N_2345);
nand U2404 (N_2404,N_2382,N_2308);
nand U2405 (N_2405,N_2311,N_2330);
or U2406 (N_2406,N_2374,N_2301);
nor U2407 (N_2407,N_2352,N_2320);
or U2408 (N_2408,N_2388,N_2393);
nand U2409 (N_2409,N_2384,N_2338);
and U2410 (N_2410,N_2346,N_2321);
or U2411 (N_2411,N_2343,N_2363);
nand U2412 (N_2412,N_2317,N_2376);
and U2413 (N_2413,N_2309,N_2340);
and U2414 (N_2414,N_2316,N_2359);
and U2415 (N_2415,N_2315,N_2314);
nor U2416 (N_2416,N_2325,N_2322);
nand U2417 (N_2417,N_2313,N_2344);
nand U2418 (N_2418,N_2377,N_2332);
or U2419 (N_2419,N_2327,N_2390);
and U2420 (N_2420,N_2306,N_2366);
and U2421 (N_2421,N_2333,N_2341);
nor U2422 (N_2422,N_2395,N_2372);
nand U2423 (N_2423,N_2328,N_2355);
nor U2424 (N_2424,N_2358,N_2368);
or U2425 (N_2425,N_2334,N_2370);
nand U2426 (N_2426,N_2369,N_2356);
or U2427 (N_2427,N_2385,N_2305);
or U2428 (N_2428,N_2361,N_2307);
nor U2429 (N_2429,N_2383,N_2324);
or U2430 (N_2430,N_2323,N_2381);
nor U2431 (N_2431,N_2300,N_2360);
nor U2432 (N_2432,N_2336,N_2389);
nor U2433 (N_2433,N_2347,N_2379);
nor U2434 (N_2434,N_2350,N_2302);
nor U2435 (N_2435,N_2357,N_2342);
or U2436 (N_2436,N_2394,N_2364);
nor U2437 (N_2437,N_2335,N_2351);
nor U2438 (N_2438,N_2399,N_2387);
or U2439 (N_2439,N_2310,N_2365);
or U2440 (N_2440,N_2375,N_2326);
and U2441 (N_2441,N_2362,N_2331);
or U2442 (N_2442,N_2396,N_2397);
or U2443 (N_2443,N_2349,N_2392);
or U2444 (N_2444,N_2354,N_2319);
nor U2445 (N_2445,N_2386,N_2303);
nand U2446 (N_2446,N_2329,N_2339);
or U2447 (N_2447,N_2348,N_2391);
or U2448 (N_2448,N_2367,N_2312);
or U2449 (N_2449,N_2371,N_2304);
nand U2450 (N_2450,N_2379,N_2312);
nand U2451 (N_2451,N_2395,N_2391);
nand U2452 (N_2452,N_2339,N_2326);
nand U2453 (N_2453,N_2377,N_2315);
or U2454 (N_2454,N_2328,N_2370);
nor U2455 (N_2455,N_2397,N_2373);
nor U2456 (N_2456,N_2383,N_2336);
or U2457 (N_2457,N_2316,N_2390);
or U2458 (N_2458,N_2383,N_2301);
nand U2459 (N_2459,N_2378,N_2349);
or U2460 (N_2460,N_2349,N_2332);
or U2461 (N_2461,N_2313,N_2377);
nand U2462 (N_2462,N_2318,N_2372);
nand U2463 (N_2463,N_2356,N_2315);
or U2464 (N_2464,N_2323,N_2319);
or U2465 (N_2465,N_2321,N_2335);
and U2466 (N_2466,N_2358,N_2316);
and U2467 (N_2467,N_2393,N_2323);
nor U2468 (N_2468,N_2335,N_2339);
or U2469 (N_2469,N_2313,N_2349);
and U2470 (N_2470,N_2361,N_2328);
nand U2471 (N_2471,N_2379,N_2310);
and U2472 (N_2472,N_2340,N_2322);
nand U2473 (N_2473,N_2355,N_2334);
or U2474 (N_2474,N_2307,N_2302);
nand U2475 (N_2475,N_2359,N_2307);
nor U2476 (N_2476,N_2330,N_2362);
and U2477 (N_2477,N_2320,N_2348);
and U2478 (N_2478,N_2311,N_2357);
nor U2479 (N_2479,N_2313,N_2335);
nor U2480 (N_2480,N_2383,N_2377);
nand U2481 (N_2481,N_2346,N_2396);
or U2482 (N_2482,N_2324,N_2308);
nand U2483 (N_2483,N_2387,N_2345);
or U2484 (N_2484,N_2309,N_2394);
nor U2485 (N_2485,N_2335,N_2364);
nor U2486 (N_2486,N_2370,N_2377);
nor U2487 (N_2487,N_2343,N_2388);
nor U2488 (N_2488,N_2357,N_2333);
or U2489 (N_2489,N_2355,N_2360);
and U2490 (N_2490,N_2360,N_2389);
or U2491 (N_2491,N_2342,N_2337);
nand U2492 (N_2492,N_2333,N_2338);
or U2493 (N_2493,N_2303,N_2317);
nand U2494 (N_2494,N_2365,N_2385);
xor U2495 (N_2495,N_2373,N_2343);
and U2496 (N_2496,N_2399,N_2335);
nor U2497 (N_2497,N_2382,N_2313);
nor U2498 (N_2498,N_2383,N_2372);
nand U2499 (N_2499,N_2354,N_2340);
nand U2500 (N_2500,N_2481,N_2459);
nand U2501 (N_2501,N_2435,N_2444);
or U2502 (N_2502,N_2454,N_2455);
and U2503 (N_2503,N_2452,N_2449);
or U2504 (N_2504,N_2410,N_2424);
or U2505 (N_2505,N_2470,N_2460);
nand U2506 (N_2506,N_2498,N_2485);
and U2507 (N_2507,N_2446,N_2417);
nand U2508 (N_2508,N_2490,N_2423);
nor U2509 (N_2509,N_2409,N_2489);
nor U2510 (N_2510,N_2432,N_2427);
nand U2511 (N_2511,N_2493,N_2422);
or U2512 (N_2512,N_2436,N_2406);
nand U2513 (N_2513,N_2407,N_2497);
nand U2514 (N_2514,N_2414,N_2491);
nand U2515 (N_2515,N_2492,N_2415);
nand U2516 (N_2516,N_2473,N_2472);
or U2517 (N_2517,N_2486,N_2428);
and U2518 (N_2518,N_2440,N_2411);
nand U2519 (N_2519,N_2457,N_2469);
or U2520 (N_2520,N_2462,N_2453);
nor U2521 (N_2521,N_2434,N_2403);
nor U2522 (N_2522,N_2448,N_2431);
and U2523 (N_2523,N_2447,N_2438);
and U2524 (N_2524,N_2476,N_2441);
nor U2525 (N_2525,N_2419,N_2404);
nor U2526 (N_2526,N_2445,N_2468);
and U2527 (N_2527,N_2477,N_2433);
nor U2528 (N_2528,N_2418,N_2412);
nor U2529 (N_2529,N_2458,N_2484);
nor U2530 (N_2530,N_2464,N_2416);
or U2531 (N_2531,N_2420,N_2437);
and U2532 (N_2532,N_2495,N_2465);
nand U2533 (N_2533,N_2478,N_2496);
or U2534 (N_2534,N_2400,N_2451);
nor U2535 (N_2535,N_2443,N_2421);
or U2536 (N_2536,N_2426,N_2430);
or U2537 (N_2537,N_2488,N_2405);
or U2538 (N_2538,N_2474,N_2401);
and U2539 (N_2539,N_2466,N_2479);
nand U2540 (N_2540,N_2499,N_2408);
nand U2541 (N_2541,N_2442,N_2429);
nor U2542 (N_2542,N_2480,N_2483);
nor U2543 (N_2543,N_2413,N_2471);
nor U2544 (N_2544,N_2402,N_2494);
and U2545 (N_2545,N_2461,N_2439);
xor U2546 (N_2546,N_2475,N_2487);
and U2547 (N_2547,N_2482,N_2425);
nand U2548 (N_2548,N_2450,N_2456);
nor U2549 (N_2549,N_2467,N_2463);
nor U2550 (N_2550,N_2462,N_2441);
or U2551 (N_2551,N_2478,N_2418);
nand U2552 (N_2552,N_2415,N_2469);
nor U2553 (N_2553,N_2464,N_2456);
or U2554 (N_2554,N_2414,N_2439);
nand U2555 (N_2555,N_2462,N_2468);
nand U2556 (N_2556,N_2426,N_2438);
nor U2557 (N_2557,N_2482,N_2432);
nor U2558 (N_2558,N_2412,N_2415);
and U2559 (N_2559,N_2430,N_2465);
nand U2560 (N_2560,N_2437,N_2484);
nand U2561 (N_2561,N_2476,N_2461);
nor U2562 (N_2562,N_2491,N_2446);
or U2563 (N_2563,N_2456,N_2432);
or U2564 (N_2564,N_2465,N_2429);
nand U2565 (N_2565,N_2412,N_2454);
or U2566 (N_2566,N_2406,N_2459);
or U2567 (N_2567,N_2400,N_2438);
or U2568 (N_2568,N_2403,N_2441);
nor U2569 (N_2569,N_2464,N_2433);
nor U2570 (N_2570,N_2469,N_2405);
nand U2571 (N_2571,N_2436,N_2459);
or U2572 (N_2572,N_2434,N_2402);
nor U2573 (N_2573,N_2462,N_2411);
and U2574 (N_2574,N_2466,N_2468);
xnor U2575 (N_2575,N_2425,N_2413);
nand U2576 (N_2576,N_2488,N_2428);
nor U2577 (N_2577,N_2400,N_2412);
and U2578 (N_2578,N_2497,N_2482);
nand U2579 (N_2579,N_2418,N_2435);
nand U2580 (N_2580,N_2449,N_2462);
nor U2581 (N_2581,N_2428,N_2431);
and U2582 (N_2582,N_2447,N_2442);
or U2583 (N_2583,N_2420,N_2435);
nor U2584 (N_2584,N_2476,N_2480);
nor U2585 (N_2585,N_2423,N_2488);
or U2586 (N_2586,N_2434,N_2419);
or U2587 (N_2587,N_2453,N_2419);
nor U2588 (N_2588,N_2471,N_2434);
nor U2589 (N_2589,N_2458,N_2456);
or U2590 (N_2590,N_2412,N_2421);
xor U2591 (N_2591,N_2432,N_2423);
nor U2592 (N_2592,N_2417,N_2418);
nand U2593 (N_2593,N_2438,N_2435);
or U2594 (N_2594,N_2456,N_2448);
or U2595 (N_2595,N_2499,N_2490);
nand U2596 (N_2596,N_2436,N_2463);
and U2597 (N_2597,N_2430,N_2408);
or U2598 (N_2598,N_2464,N_2470);
and U2599 (N_2599,N_2405,N_2414);
and U2600 (N_2600,N_2586,N_2562);
nor U2601 (N_2601,N_2571,N_2509);
nor U2602 (N_2602,N_2573,N_2503);
and U2603 (N_2603,N_2504,N_2595);
nor U2604 (N_2604,N_2560,N_2544);
nor U2605 (N_2605,N_2579,N_2512);
nand U2606 (N_2606,N_2572,N_2538);
and U2607 (N_2607,N_2556,N_2580);
nor U2608 (N_2608,N_2514,N_2505);
and U2609 (N_2609,N_2561,N_2546);
and U2610 (N_2610,N_2585,N_2536);
and U2611 (N_2611,N_2513,N_2549);
and U2612 (N_2612,N_2593,N_2576);
or U2613 (N_2613,N_2596,N_2592);
nand U2614 (N_2614,N_2526,N_2584);
nand U2615 (N_2615,N_2574,N_2589);
and U2616 (N_2616,N_2507,N_2559);
and U2617 (N_2617,N_2540,N_2570);
xor U2618 (N_2618,N_2598,N_2565);
nor U2619 (N_2619,N_2537,N_2558);
or U2620 (N_2620,N_2531,N_2582);
and U2621 (N_2621,N_2569,N_2588);
nor U2622 (N_2622,N_2522,N_2567);
and U2623 (N_2623,N_2506,N_2523);
or U2624 (N_2624,N_2518,N_2566);
and U2625 (N_2625,N_2568,N_2519);
or U2626 (N_2626,N_2581,N_2548);
nor U2627 (N_2627,N_2543,N_2500);
nor U2628 (N_2628,N_2590,N_2551);
nor U2629 (N_2629,N_2555,N_2510);
nor U2630 (N_2630,N_2516,N_2564);
nor U2631 (N_2631,N_2599,N_2502);
or U2632 (N_2632,N_2528,N_2553);
and U2633 (N_2633,N_2524,N_2578);
nor U2634 (N_2634,N_2515,N_2545);
and U2635 (N_2635,N_2508,N_2532);
or U2636 (N_2636,N_2535,N_2539);
nand U2637 (N_2637,N_2587,N_2554);
and U2638 (N_2638,N_2550,N_2517);
nand U2639 (N_2639,N_2541,N_2597);
or U2640 (N_2640,N_2557,N_2511);
and U2641 (N_2641,N_2520,N_2521);
or U2642 (N_2642,N_2591,N_2583);
and U2643 (N_2643,N_2501,N_2533);
or U2644 (N_2644,N_2529,N_2594);
or U2645 (N_2645,N_2527,N_2542);
nor U2646 (N_2646,N_2575,N_2552);
or U2647 (N_2647,N_2525,N_2534);
nor U2648 (N_2648,N_2530,N_2577);
and U2649 (N_2649,N_2563,N_2547);
nor U2650 (N_2650,N_2589,N_2556);
xnor U2651 (N_2651,N_2574,N_2536);
or U2652 (N_2652,N_2568,N_2554);
or U2653 (N_2653,N_2565,N_2544);
and U2654 (N_2654,N_2507,N_2587);
or U2655 (N_2655,N_2511,N_2533);
or U2656 (N_2656,N_2507,N_2522);
nor U2657 (N_2657,N_2529,N_2514);
nor U2658 (N_2658,N_2562,N_2500);
nand U2659 (N_2659,N_2525,N_2589);
and U2660 (N_2660,N_2577,N_2535);
or U2661 (N_2661,N_2591,N_2566);
and U2662 (N_2662,N_2591,N_2578);
or U2663 (N_2663,N_2507,N_2518);
or U2664 (N_2664,N_2509,N_2559);
nand U2665 (N_2665,N_2574,N_2514);
or U2666 (N_2666,N_2564,N_2562);
nand U2667 (N_2667,N_2547,N_2513);
or U2668 (N_2668,N_2549,N_2563);
and U2669 (N_2669,N_2555,N_2594);
nor U2670 (N_2670,N_2550,N_2537);
nor U2671 (N_2671,N_2563,N_2552);
nor U2672 (N_2672,N_2598,N_2593);
and U2673 (N_2673,N_2544,N_2590);
and U2674 (N_2674,N_2564,N_2507);
and U2675 (N_2675,N_2514,N_2524);
or U2676 (N_2676,N_2538,N_2586);
or U2677 (N_2677,N_2515,N_2598);
nor U2678 (N_2678,N_2546,N_2520);
nand U2679 (N_2679,N_2591,N_2505);
or U2680 (N_2680,N_2582,N_2591);
nand U2681 (N_2681,N_2565,N_2563);
and U2682 (N_2682,N_2500,N_2592);
or U2683 (N_2683,N_2528,N_2524);
nand U2684 (N_2684,N_2517,N_2555);
or U2685 (N_2685,N_2564,N_2523);
or U2686 (N_2686,N_2540,N_2579);
or U2687 (N_2687,N_2514,N_2569);
nand U2688 (N_2688,N_2571,N_2572);
or U2689 (N_2689,N_2562,N_2589);
nand U2690 (N_2690,N_2534,N_2579);
nand U2691 (N_2691,N_2568,N_2548);
and U2692 (N_2692,N_2560,N_2568);
or U2693 (N_2693,N_2531,N_2562);
nand U2694 (N_2694,N_2561,N_2539);
or U2695 (N_2695,N_2565,N_2552);
or U2696 (N_2696,N_2515,N_2508);
or U2697 (N_2697,N_2543,N_2513);
and U2698 (N_2698,N_2569,N_2583);
or U2699 (N_2699,N_2514,N_2538);
nand U2700 (N_2700,N_2698,N_2667);
or U2701 (N_2701,N_2603,N_2642);
or U2702 (N_2702,N_2614,N_2630);
or U2703 (N_2703,N_2690,N_2687);
nand U2704 (N_2704,N_2670,N_2602);
nor U2705 (N_2705,N_2638,N_2682);
or U2706 (N_2706,N_2649,N_2613);
and U2707 (N_2707,N_2622,N_2669);
nor U2708 (N_2708,N_2699,N_2612);
nor U2709 (N_2709,N_2627,N_2673);
and U2710 (N_2710,N_2607,N_2666);
nand U2711 (N_2711,N_2654,N_2668);
or U2712 (N_2712,N_2657,N_2691);
and U2713 (N_2713,N_2604,N_2647);
nor U2714 (N_2714,N_2631,N_2609);
nand U2715 (N_2715,N_2653,N_2623);
and U2716 (N_2716,N_2628,N_2674);
and U2717 (N_2717,N_2629,N_2662);
and U2718 (N_2718,N_2646,N_2635);
and U2719 (N_2719,N_2685,N_2681);
or U2720 (N_2720,N_2694,N_2651);
nor U2721 (N_2721,N_2655,N_2621);
nand U2722 (N_2722,N_2665,N_2688);
nor U2723 (N_2723,N_2624,N_2615);
nand U2724 (N_2724,N_2689,N_2640);
nand U2725 (N_2725,N_2697,N_2680);
nor U2726 (N_2726,N_2632,N_2679);
or U2727 (N_2727,N_2608,N_2606);
and U2728 (N_2728,N_2692,N_2671);
nand U2729 (N_2729,N_2634,N_2650);
nor U2730 (N_2730,N_2660,N_2611);
nor U2731 (N_2731,N_2663,N_2672);
and U2732 (N_2732,N_2616,N_2643);
nor U2733 (N_2733,N_2601,N_2678);
and U2734 (N_2734,N_2645,N_2625);
and U2735 (N_2735,N_2695,N_2617);
and U2736 (N_2736,N_2641,N_2610);
or U2737 (N_2737,N_2664,N_2659);
or U2738 (N_2738,N_2677,N_2658);
nor U2739 (N_2739,N_2639,N_2600);
nor U2740 (N_2740,N_2656,N_2693);
nand U2741 (N_2741,N_2648,N_2686);
nand U2742 (N_2742,N_2661,N_2684);
nor U2743 (N_2743,N_2626,N_2676);
or U2744 (N_2744,N_2675,N_2637);
nand U2745 (N_2745,N_2618,N_2683);
nand U2746 (N_2746,N_2652,N_2620);
and U2747 (N_2747,N_2633,N_2696);
or U2748 (N_2748,N_2619,N_2605);
nor U2749 (N_2749,N_2644,N_2636);
nor U2750 (N_2750,N_2677,N_2631);
or U2751 (N_2751,N_2625,N_2677);
or U2752 (N_2752,N_2636,N_2694);
and U2753 (N_2753,N_2653,N_2684);
and U2754 (N_2754,N_2666,N_2619);
nor U2755 (N_2755,N_2654,N_2633);
nor U2756 (N_2756,N_2644,N_2601);
nand U2757 (N_2757,N_2677,N_2607);
and U2758 (N_2758,N_2679,N_2651);
nor U2759 (N_2759,N_2609,N_2602);
or U2760 (N_2760,N_2674,N_2687);
nand U2761 (N_2761,N_2615,N_2643);
nand U2762 (N_2762,N_2621,N_2688);
and U2763 (N_2763,N_2656,N_2605);
and U2764 (N_2764,N_2657,N_2659);
nor U2765 (N_2765,N_2682,N_2601);
nor U2766 (N_2766,N_2635,N_2629);
nor U2767 (N_2767,N_2686,N_2679);
or U2768 (N_2768,N_2685,N_2641);
or U2769 (N_2769,N_2602,N_2612);
nand U2770 (N_2770,N_2638,N_2657);
or U2771 (N_2771,N_2672,N_2696);
nor U2772 (N_2772,N_2637,N_2652);
or U2773 (N_2773,N_2637,N_2670);
nand U2774 (N_2774,N_2615,N_2667);
nor U2775 (N_2775,N_2626,N_2678);
nor U2776 (N_2776,N_2630,N_2653);
or U2777 (N_2777,N_2617,N_2628);
and U2778 (N_2778,N_2606,N_2644);
or U2779 (N_2779,N_2661,N_2690);
nor U2780 (N_2780,N_2681,N_2614);
nor U2781 (N_2781,N_2673,N_2604);
nand U2782 (N_2782,N_2618,N_2625);
nor U2783 (N_2783,N_2634,N_2618);
and U2784 (N_2784,N_2676,N_2633);
nor U2785 (N_2785,N_2621,N_2604);
and U2786 (N_2786,N_2643,N_2655);
nor U2787 (N_2787,N_2648,N_2663);
or U2788 (N_2788,N_2638,N_2611);
or U2789 (N_2789,N_2602,N_2698);
and U2790 (N_2790,N_2676,N_2686);
nor U2791 (N_2791,N_2613,N_2678);
or U2792 (N_2792,N_2643,N_2618);
and U2793 (N_2793,N_2671,N_2648);
nor U2794 (N_2794,N_2632,N_2625);
nor U2795 (N_2795,N_2671,N_2651);
and U2796 (N_2796,N_2674,N_2640);
and U2797 (N_2797,N_2688,N_2662);
and U2798 (N_2798,N_2616,N_2651);
nor U2799 (N_2799,N_2640,N_2608);
nand U2800 (N_2800,N_2746,N_2751);
and U2801 (N_2801,N_2729,N_2760);
nor U2802 (N_2802,N_2745,N_2757);
xor U2803 (N_2803,N_2790,N_2771);
nor U2804 (N_2804,N_2780,N_2700);
xor U2805 (N_2805,N_2755,N_2766);
or U2806 (N_2806,N_2737,N_2794);
nand U2807 (N_2807,N_2748,N_2769);
or U2808 (N_2808,N_2708,N_2798);
nor U2809 (N_2809,N_2726,N_2709);
or U2810 (N_2810,N_2779,N_2725);
or U2811 (N_2811,N_2722,N_2759);
nor U2812 (N_2812,N_2735,N_2744);
nor U2813 (N_2813,N_2796,N_2784);
or U2814 (N_2814,N_2739,N_2753);
and U2815 (N_2815,N_2734,N_2789);
or U2816 (N_2816,N_2781,N_2707);
or U2817 (N_2817,N_2783,N_2791);
or U2818 (N_2818,N_2736,N_2711);
nand U2819 (N_2819,N_2742,N_2764);
nand U2820 (N_2820,N_2763,N_2733);
and U2821 (N_2821,N_2724,N_2799);
nor U2822 (N_2822,N_2717,N_2710);
or U2823 (N_2823,N_2773,N_2732);
and U2824 (N_2824,N_2728,N_2767);
nor U2825 (N_2825,N_2752,N_2718);
and U2826 (N_2826,N_2754,N_2721);
and U2827 (N_2827,N_2743,N_2740);
nor U2828 (N_2828,N_2793,N_2762);
and U2829 (N_2829,N_2730,N_2712);
and U2830 (N_2830,N_2705,N_2706);
nor U2831 (N_2831,N_2749,N_2788);
or U2832 (N_2832,N_2787,N_2731);
or U2833 (N_2833,N_2741,N_2756);
and U2834 (N_2834,N_2703,N_2797);
nor U2835 (N_2835,N_2785,N_2747);
nand U2836 (N_2836,N_2770,N_2782);
nand U2837 (N_2837,N_2778,N_2774);
or U2838 (N_2838,N_2704,N_2768);
nand U2839 (N_2839,N_2758,N_2723);
nand U2840 (N_2840,N_2750,N_2772);
or U2841 (N_2841,N_2713,N_2716);
or U2842 (N_2842,N_2719,N_2786);
nor U2843 (N_2843,N_2727,N_2777);
nor U2844 (N_2844,N_2775,N_2795);
xnor U2845 (N_2845,N_2720,N_2761);
or U2846 (N_2846,N_2776,N_2715);
and U2847 (N_2847,N_2701,N_2702);
nor U2848 (N_2848,N_2792,N_2765);
and U2849 (N_2849,N_2714,N_2738);
nor U2850 (N_2850,N_2753,N_2764);
and U2851 (N_2851,N_2732,N_2729);
and U2852 (N_2852,N_2722,N_2784);
nor U2853 (N_2853,N_2724,N_2788);
xor U2854 (N_2854,N_2772,N_2714);
and U2855 (N_2855,N_2775,N_2753);
and U2856 (N_2856,N_2729,N_2748);
nor U2857 (N_2857,N_2774,N_2751);
and U2858 (N_2858,N_2719,N_2724);
xnor U2859 (N_2859,N_2768,N_2707);
or U2860 (N_2860,N_2737,N_2722);
and U2861 (N_2861,N_2778,N_2784);
nor U2862 (N_2862,N_2769,N_2745);
nor U2863 (N_2863,N_2723,N_2782);
nor U2864 (N_2864,N_2758,N_2711);
and U2865 (N_2865,N_2738,N_2758);
or U2866 (N_2866,N_2787,N_2732);
nor U2867 (N_2867,N_2738,N_2769);
and U2868 (N_2868,N_2771,N_2727);
and U2869 (N_2869,N_2798,N_2796);
or U2870 (N_2870,N_2725,N_2723);
and U2871 (N_2871,N_2779,N_2746);
nand U2872 (N_2872,N_2775,N_2780);
or U2873 (N_2873,N_2736,N_2710);
nand U2874 (N_2874,N_2795,N_2704);
xnor U2875 (N_2875,N_2793,N_2722);
nor U2876 (N_2876,N_2731,N_2715);
xor U2877 (N_2877,N_2775,N_2762);
nor U2878 (N_2878,N_2716,N_2722);
and U2879 (N_2879,N_2798,N_2701);
or U2880 (N_2880,N_2701,N_2773);
nand U2881 (N_2881,N_2716,N_2789);
or U2882 (N_2882,N_2719,N_2742);
or U2883 (N_2883,N_2715,N_2785);
nor U2884 (N_2884,N_2785,N_2724);
or U2885 (N_2885,N_2743,N_2787);
nand U2886 (N_2886,N_2765,N_2797);
xnor U2887 (N_2887,N_2746,N_2711);
nand U2888 (N_2888,N_2735,N_2732);
and U2889 (N_2889,N_2720,N_2775);
or U2890 (N_2890,N_2775,N_2742);
nor U2891 (N_2891,N_2730,N_2770);
nand U2892 (N_2892,N_2773,N_2726);
or U2893 (N_2893,N_2766,N_2703);
and U2894 (N_2894,N_2744,N_2715);
nand U2895 (N_2895,N_2703,N_2770);
and U2896 (N_2896,N_2731,N_2708);
nand U2897 (N_2897,N_2714,N_2765);
nand U2898 (N_2898,N_2712,N_2764);
nor U2899 (N_2899,N_2728,N_2778);
xnor U2900 (N_2900,N_2836,N_2818);
nor U2901 (N_2901,N_2865,N_2857);
and U2902 (N_2902,N_2813,N_2819);
xor U2903 (N_2903,N_2812,N_2859);
nor U2904 (N_2904,N_2861,N_2827);
and U2905 (N_2905,N_2870,N_2806);
nand U2906 (N_2906,N_2872,N_2856);
nand U2907 (N_2907,N_2845,N_2850);
nor U2908 (N_2908,N_2863,N_2895);
or U2909 (N_2909,N_2860,N_2855);
or U2910 (N_2910,N_2893,N_2822);
nor U2911 (N_2911,N_2874,N_2887);
and U2912 (N_2912,N_2849,N_2864);
or U2913 (N_2913,N_2805,N_2815);
and U2914 (N_2914,N_2878,N_2837);
or U2915 (N_2915,N_2834,N_2880);
nor U2916 (N_2916,N_2840,N_2891);
or U2917 (N_2917,N_2897,N_2825);
nand U2918 (N_2918,N_2877,N_2810);
and U2919 (N_2919,N_2883,N_2885);
nand U2920 (N_2920,N_2809,N_2800);
nand U2921 (N_2921,N_2842,N_2811);
or U2922 (N_2922,N_2851,N_2826);
nand U2923 (N_2923,N_2816,N_2898);
and U2924 (N_2924,N_2831,N_2876);
or U2925 (N_2925,N_2833,N_2892);
nand U2926 (N_2926,N_2839,N_2890);
nor U2927 (N_2927,N_2888,N_2866);
nand U2928 (N_2928,N_2802,N_2828);
nand U2929 (N_2929,N_2801,N_2841);
and U2930 (N_2930,N_2830,N_2889);
or U2931 (N_2931,N_2896,N_2846);
nor U2932 (N_2932,N_2899,N_2852);
and U2933 (N_2933,N_2829,N_2853);
and U2934 (N_2934,N_2871,N_2808);
or U2935 (N_2935,N_2867,N_2879);
and U2936 (N_2936,N_2854,N_2847);
nor U2937 (N_2937,N_2821,N_2817);
and U2938 (N_2938,N_2814,N_2838);
nor U2939 (N_2939,N_2868,N_2881);
nand U2940 (N_2940,N_2894,N_2844);
nand U2941 (N_2941,N_2884,N_2804);
or U2942 (N_2942,N_2869,N_2843);
nor U2943 (N_2943,N_2832,N_2873);
nand U2944 (N_2944,N_2858,N_2824);
nor U2945 (N_2945,N_2886,N_2803);
nand U2946 (N_2946,N_2848,N_2807);
and U2947 (N_2947,N_2835,N_2823);
nand U2948 (N_2948,N_2862,N_2882);
nand U2949 (N_2949,N_2820,N_2875);
nor U2950 (N_2950,N_2877,N_2828);
nor U2951 (N_2951,N_2809,N_2829);
nand U2952 (N_2952,N_2846,N_2881);
nand U2953 (N_2953,N_2823,N_2872);
and U2954 (N_2954,N_2868,N_2871);
nor U2955 (N_2955,N_2823,N_2803);
or U2956 (N_2956,N_2863,N_2854);
and U2957 (N_2957,N_2857,N_2837);
or U2958 (N_2958,N_2851,N_2873);
nor U2959 (N_2959,N_2819,N_2889);
or U2960 (N_2960,N_2801,N_2846);
nor U2961 (N_2961,N_2807,N_2816);
or U2962 (N_2962,N_2836,N_2863);
nor U2963 (N_2963,N_2807,N_2812);
nor U2964 (N_2964,N_2820,N_2850);
and U2965 (N_2965,N_2892,N_2834);
nand U2966 (N_2966,N_2820,N_2825);
nor U2967 (N_2967,N_2807,N_2827);
nand U2968 (N_2968,N_2819,N_2803);
nor U2969 (N_2969,N_2885,N_2818);
nor U2970 (N_2970,N_2834,N_2879);
and U2971 (N_2971,N_2880,N_2807);
nand U2972 (N_2972,N_2874,N_2891);
and U2973 (N_2973,N_2857,N_2894);
or U2974 (N_2974,N_2859,N_2828);
nand U2975 (N_2975,N_2879,N_2856);
nor U2976 (N_2976,N_2858,N_2893);
and U2977 (N_2977,N_2871,N_2818);
nand U2978 (N_2978,N_2810,N_2849);
nor U2979 (N_2979,N_2809,N_2851);
and U2980 (N_2980,N_2858,N_2838);
nand U2981 (N_2981,N_2830,N_2807);
nor U2982 (N_2982,N_2867,N_2875);
or U2983 (N_2983,N_2841,N_2805);
nand U2984 (N_2984,N_2889,N_2880);
nand U2985 (N_2985,N_2874,N_2894);
and U2986 (N_2986,N_2871,N_2823);
nand U2987 (N_2987,N_2821,N_2857);
and U2988 (N_2988,N_2896,N_2800);
nor U2989 (N_2989,N_2818,N_2886);
nand U2990 (N_2990,N_2803,N_2835);
nor U2991 (N_2991,N_2838,N_2895);
nand U2992 (N_2992,N_2857,N_2853);
nand U2993 (N_2993,N_2830,N_2832);
and U2994 (N_2994,N_2888,N_2800);
or U2995 (N_2995,N_2843,N_2854);
nand U2996 (N_2996,N_2867,N_2899);
and U2997 (N_2997,N_2889,N_2817);
and U2998 (N_2998,N_2898,N_2841);
nand U2999 (N_2999,N_2863,N_2881);
and UO_0 (O_0,N_2908,N_2901);
and UO_1 (O_1,N_2973,N_2967);
nor UO_2 (O_2,N_2929,N_2955);
or UO_3 (O_3,N_2968,N_2945);
and UO_4 (O_4,N_2963,N_2910);
nor UO_5 (O_5,N_2966,N_2991);
nor UO_6 (O_6,N_2999,N_2972);
nor UO_7 (O_7,N_2950,N_2982);
or UO_8 (O_8,N_2949,N_2978);
or UO_9 (O_9,N_2917,N_2965);
nand UO_10 (O_10,N_2960,N_2934);
or UO_11 (O_11,N_2969,N_2971);
or UO_12 (O_12,N_2933,N_2995);
nand UO_13 (O_13,N_2947,N_2911);
and UO_14 (O_14,N_2948,N_2976);
nand UO_15 (O_15,N_2962,N_2957);
nand UO_16 (O_16,N_2935,N_2993);
nor UO_17 (O_17,N_2900,N_2970);
or UO_18 (O_18,N_2975,N_2919);
nand UO_19 (O_19,N_2939,N_2904);
nand UO_20 (O_20,N_2902,N_2918);
nor UO_21 (O_21,N_2997,N_2907);
and UO_22 (O_22,N_2928,N_2905);
or UO_23 (O_23,N_2938,N_2984);
nor UO_24 (O_24,N_2925,N_2914);
and UO_25 (O_25,N_2903,N_2959);
nor UO_26 (O_26,N_2921,N_2994);
and UO_27 (O_27,N_2942,N_2990);
and UO_28 (O_28,N_2927,N_2964);
and UO_29 (O_29,N_2977,N_2916);
nand UO_30 (O_30,N_2981,N_2913);
nor UO_31 (O_31,N_2952,N_2932);
and UO_32 (O_32,N_2909,N_2912);
nor UO_33 (O_33,N_2961,N_2958);
nor UO_34 (O_34,N_2954,N_2988);
nor UO_35 (O_35,N_2946,N_2941);
nor UO_36 (O_36,N_2937,N_2983);
and UO_37 (O_37,N_2980,N_2953);
nor UO_38 (O_38,N_2940,N_2936);
or UO_39 (O_39,N_2920,N_2985);
or UO_40 (O_40,N_2943,N_2956);
nand UO_41 (O_41,N_2989,N_2923);
nor UO_42 (O_42,N_2998,N_2979);
nor UO_43 (O_43,N_2996,N_2992);
or UO_44 (O_44,N_2987,N_2974);
nor UO_45 (O_45,N_2906,N_2915);
nor UO_46 (O_46,N_2951,N_2944);
nand UO_47 (O_47,N_2924,N_2930);
or UO_48 (O_48,N_2931,N_2926);
nor UO_49 (O_49,N_2986,N_2922);
nand UO_50 (O_50,N_2941,N_2908);
nand UO_51 (O_51,N_2927,N_2996);
nor UO_52 (O_52,N_2978,N_2933);
or UO_53 (O_53,N_2993,N_2913);
and UO_54 (O_54,N_2936,N_2969);
and UO_55 (O_55,N_2968,N_2939);
and UO_56 (O_56,N_2982,N_2903);
nand UO_57 (O_57,N_2998,N_2921);
and UO_58 (O_58,N_2939,N_2907);
nor UO_59 (O_59,N_2932,N_2981);
nand UO_60 (O_60,N_2990,N_2914);
nand UO_61 (O_61,N_2912,N_2908);
or UO_62 (O_62,N_2955,N_2952);
nor UO_63 (O_63,N_2996,N_2945);
nand UO_64 (O_64,N_2980,N_2910);
nand UO_65 (O_65,N_2927,N_2971);
or UO_66 (O_66,N_2900,N_2932);
and UO_67 (O_67,N_2938,N_2980);
nor UO_68 (O_68,N_2985,N_2990);
nand UO_69 (O_69,N_2988,N_2984);
nor UO_70 (O_70,N_2918,N_2989);
nor UO_71 (O_71,N_2956,N_2971);
and UO_72 (O_72,N_2962,N_2997);
nor UO_73 (O_73,N_2973,N_2907);
nand UO_74 (O_74,N_2905,N_2932);
nor UO_75 (O_75,N_2955,N_2944);
or UO_76 (O_76,N_2929,N_2976);
nor UO_77 (O_77,N_2939,N_2923);
nand UO_78 (O_78,N_2913,N_2939);
and UO_79 (O_79,N_2987,N_2958);
nand UO_80 (O_80,N_2962,N_2943);
nand UO_81 (O_81,N_2970,N_2977);
nor UO_82 (O_82,N_2933,N_2990);
nand UO_83 (O_83,N_2914,N_2955);
and UO_84 (O_84,N_2956,N_2923);
or UO_85 (O_85,N_2997,N_2935);
and UO_86 (O_86,N_2907,N_2920);
nand UO_87 (O_87,N_2929,N_2918);
nand UO_88 (O_88,N_2958,N_2960);
and UO_89 (O_89,N_2995,N_2991);
or UO_90 (O_90,N_2964,N_2966);
or UO_91 (O_91,N_2991,N_2904);
and UO_92 (O_92,N_2959,N_2977);
and UO_93 (O_93,N_2983,N_2954);
and UO_94 (O_94,N_2906,N_2968);
nor UO_95 (O_95,N_2989,N_2931);
nor UO_96 (O_96,N_2953,N_2928);
nor UO_97 (O_97,N_2963,N_2934);
nand UO_98 (O_98,N_2953,N_2975);
nand UO_99 (O_99,N_2973,N_2914);
nor UO_100 (O_100,N_2999,N_2932);
nand UO_101 (O_101,N_2915,N_2908);
nand UO_102 (O_102,N_2977,N_2952);
or UO_103 (O_103,N_2949,N_2956);
or UO_104 (O_104,N_2934,N_2935);
and UO_105 (O_105,N_2904,N_2943);
or UO_106 (O_106,N_2943,N_2991);
and UO_107 (O_107,N_2952,N_2931);
or UO_108 (O_108,N_2951,N_2952);
and UO_109 (O_109,N_2902,N_2994);
nand UO_110 (O_110,N_2987,N_2920);
or UO_111 (O_111,N_2903,N_2931);
and UO_112 (O_112,N_2996,N_2954);
nand UO_113 (O_113,N_2981,N_2966);
and UO_114 (O_114,N_2936,N_2922);
and UO_115 (O_115,N_2905,N_2999);
and UO_116 (O_116,N_2971,N_2957);
nand UO_117 (O_117,N_2934,N_2990);
nor UO_118 (O_118,N_2998,N_2960);
or UO_119 (O_119,N_2937,N_2992);
nand UO_120 (O_120,N_2966,N_2989);
and UO_121 (O_121,N_2985,N_2960);
or UO_122 (O_122,N_2959,N_2992);
nor UO_123 (O_123,N_2989,N_2902);
nor UO_124 (O_124,N_2975,N_2903);
or UO_125 (O_125,N_2953,N_2987);
nand UO_126 (O_126,N_2903,N_2964);
nor UO_127 (O_127,N_2995,N_2941);
nor UO_128 (O_128,N_2991,N_2950);
and UO_129 (O_129,N_2977,N_2966);
and UO_130 (O_130,N_2953,N_2999);
nor UO_131 (O_131,N_2999,N_2988);
or UO_132 (O_132,N_2995,N_2932);
nand UO_133 (O_133,N_2910,N_2990);
and UO_134 (O_134,N_2905,N_2979);
nor UO_135 (O_135,N_2949,N_2953);
nand UO_136 (O_136,N_2951,N_2912);
and UO_137 (O_137,N_2900,N_2907);
or UO_138 (O_138,N_2985,N_2971);
nor UO_139 (O_139,N_2925,N_2924);
xnor UO_140 (O_140,N_2937,N_2903);
and UO_141 (O_141,N_2963,N_2959);
or UO_142 (O_142,N_2917,N_2989);
or UO_143 (O_143,N_2986,N_2977);
nor UO_144 (O_144,N_2901,N_2925);
and UO_145 (O_145,N_2934,N_2941);
nand UO_146 (O_146,N_2904,N_2972);
or UO_147 (O_147,N_2985,N_2929);
and UO_148 (O_148,N_2956,N_2987);
nor UO_149 (O_149,N_2968,N_2914);
nand UO_150 (O_150,N_2927,N_2948);
and UO_151 (O_151,N_2964,N_2983);
and UO_152 (O_152,N_2962,N_2991);
nor UO_153 (O_153,N_2932,N_2985);
and UO_154 (O_154,N_2911,N_2967);
nor UO_155 (O_155,N_2933,N_2936);
nor UO_156 (O_156,N_2976,N_2912);
or UO_157 (O_157,N_2980,N_2909);
nand UO_158 (O_158,N_2945,N_2952);
nand UO_159 (O_159,N_2902,N_2922);
nor UO_160 (O_160,N_2934,N_2902);
nor UO_161 (O_161,N_2985,N_2931);
and UO_162 (O_162,N_2906,N_2971);
or UO_163 (O_163,N_2900,N_2961);
nor UO_164 (O_164,N_2955,N_2986);
xnor UO_165 (O_165,N_2944,N_2981);
nand UO_166 (O_166,N_2955,N_2946);
nand UO_167 (O_167,N_2984,N_2914);
nand UO_168 (O_168,N_2981,N_2933);
or UO_169 (O_169,N_2915,N_2911);
or UO_170 (O_170,N_2914,N_2963);
nor UO_171 (O_171,N_2942,N_2957);
or UO_172 (O_172,N_2947,N_2977);
or UO_173 (O_173,N_2990,N_2992);
or UO_174 (O_174,N_2914,N_2929);
or UO_175 (O_175,N_2941,N_2952);
nand UO_176 (O_176,N_2902,N_2935);
and UO_177 (O_177,N_2913,N_2945);
and UO_178 (O_178,N_2920,N_2943);
and UO_179 (O_179,N_2940,N_2909);
or UO_180 (O_180,N_2996,N_2978);
nand UO_181 (O_181,N_2988,N_2978);
nand UO_182 (O_182,N_2956,N_2936);
and UO_183 (O_183,N_2992,N_2910);
and UO_184 (O_184,N_2976,N_2913);
nand UO_185 (O_185,N_2900,N_2936);
nor UO_186 (O_186,N_2969,N_2955);
nand UO_187 (O_187,N_2999,N_2957);
nor UO_188 (O_188,N_2916,N_2964);
or UO_189 (O_189,N_2924,N_2903);
and UO_190 (O_190,N_2970,N_2972);
nor UO_191 (O_191,N_2996,N_2961);
and UO_192 (O_192,N_2900,N_2999);
or UO_193 (O_193,N_2965,N_2920);
nand UO_194 (O_194,N_2979,N_2954);
and UO_195 (O_195,N_2939,N_2964);
nand UO_196 (O_196,N_2933,N_2904);
or UO_197 (O_197,N_2916,N_2913);
and UO_198 (O_198,N_2916,N_2952);
nand UO_199 (O_199,N_2947,N_2994);
nor UO_200 (O_200,N_2970,N_2952);
and UO_201 (O_201,N_2908,N_2969);
nand UO_202 (O_202,N_2941,N_2932);
nor UO_203 (O_203,N_2955,N_2982);
or UO_204 (O_204,N_2981,N_2959);
and UO_205 (O_205,N_2983,N_2946);
nor UO_206 (O_206,N_2943,N_2972);
nor UO_207 (O_207,N_2994,N_2904);
and UO_208 (O_208,N_2962,N_2980);
and UO_209 (O_209,N_2923,N_2971);
nand UO_210 (O_210,N_2919,N_2968);
or UO_211 (O_211,N_2982,N_2914);
nand UO_212 (O_212,N_2990,N_2973);
or UO_213 (O_213,N_2958,N_2990);
or UO_214 (O_214,N_2930,N_2999);
or UO_215 (O_215,N_2995,N_2950);
or UO_216 (O_216,N_2942,N_2906);
nor UO_217 (O_217,N_2961,N_2931);
nor UO_218 (O_218,N_2912,N_2902);
and UO_219 (O_219,N_2980,N_2972);
or UO_220 (O_220,N_2936,N_2980);
nand UO_221 (O_221,N_2946,N_2969);
nand UO_222 (O_222,N_2903,N_2939);
and UO_223 (O_223,N_2985,N_2970);
or UO_224 (O_224,N_2961,N_2950);
nor UO_225 (O_225,N_2937,N_2918);
and UO_226 (O_226,N_2948,N_2929);
nand UO_227 (O_227,N_2985,N_2944);
and UO_228 (O_228,N_2904,N_2984);
nand UO_229 (O_229,N_2930,N_2920);
nand UO_230 (O_230,N_2950,N_2979);
nor UO_231 (O_231,N_2946,N_2981);
and UO_232 (O_232,N_2902,N_2917);
nand UO_233 (O_233,N_2973,N_2913);
nor UO_234 (O_234,N_2969,N_2963);
and UO_235 (O_235,N_2999,N_2979);
and UO_236 (O_236,N_2990,N_2903);
or UO_237 (O_237,N_2981,N_2928);
nand UO_238 (O_238,N_2995,N_2988);
nand UO_239 (O_239,N_2940,N_2990);
and UO_240 (O_240,N_2994,N_2901);
nand UO_241 (O_241,N_2940,N_2957);
nand UO_242 (O_242,N_2939,N_2915);
nor UO_243 (O_243,N_2912,N_2937);
nand UO_244 (O_244,N_2915,N_2933);
or UO_245 (O_245,N_2986,N_2960);
and UO_246 (O_246,N_2950,N_2919);
nand UO_247 (O_247,N_2920,N_2941);
and UO_248 (O_248,N_2933,N_2902);
nor UO_249 (O_249,N_2932,N_2940);
nand UO_250 (O_250,N_2979,N_2939);
and UO_251 (O_251,N_2905,N_2996);
nor UO_252 (O_252,N_2934,N_2968);
and UO_253 (O_253,N_2920,N_2974);
or UO_254 (O_254,N_2989,N_2912);
nor UO_255 (O_255,N_2937,N_2932);
xnor UO_256 (O_256,N_2949,N_2915);
or UO_257 (O_257,N_2917,N_2990);
nand UO_258 (O_258,N_2993,N_2946);
nor UO_259 (O_259,N_2965,N_2916);
and UO_260 (O_260,N_2918,N_2906);
nor UO_261 (O_261,N_2909,N_2959);
or UO_262 (O_262,N_2920,N_2975);
nor UO_263 (O_263,N_2900,N_2910);
or UO_264 (O_264,N_2944,N_2957);
and UO_265 (O_265,N_2988,N_2912);
nand UO_266 (O_266,N_2907,N_2956);
nor UO_267 (O_267,N_2913,N_2941);
nor UO_268 (O_268,N_2980,N_2994);
and UO_269 (O_269,N_2929,N_2970);
or UO_270 (O_270,N_2925,N_2997);
and UO_271 (O_271,N_2914,N_2952);
nand UO_272 (O_272,N_2953,N_2988);
nor UO_273 (O_273,N_2908,N_2911);
nor UO_274 (O_274,N_2949,N_2901);
nand UO_275 (O_275,N_2921,N_2922);
or UO_276 (O_276,N_2919,N_2967);
and UO_277 (O_277,N_2956,N_2988);
or UO_278 (O_278,N_2901,N_2989);
nor UO_279 (O_279,N_2969,N_2913);
or UO_280 (O_280,N_2975,N_2921);
nand UO_281 (O_281,N_2970,N_2920);
or UO_282 (O_282,N_2958,N_2985);
nor UO_283 (O_283,N_2993,N_2975);
nand UO_284 (O_284,N_2997,N_2920);
or UO_285 (O_285,N_2958,N_2914);
or UO_286 (O_286,N_2967,N_2990);
or UO_287 (O_287,N_2912,N_2973);
and UO_288 (O_288,N_2902,N_2976);
nand UO_289 (O_289,N_2992,N_2963);
or UO_290 (O_290,N_2971,N_2980);
nand UO_291 (O_291,N_2961,N_2924);
nor UO_292 (O_292,N_2980,N_2920);
and UO_293 (O_293,N_2958,N_2941);
or UO_294 (O_294,N_2999,N_2914);
nor UO_295 (O_295,N_2925,N_2960);
nand UO_296 (O_296,N_2986,N_2900);
nor UO_297 (O_297,N_2903,N_2965);
nand UO_298 (O_298,N_2989,N_2978);
and UO_299 (O_299,N_2916,N_2979);
or UO_300 (O_300,N_2952,N_2990);
nor UO_301 (O_301,N_2970,N_2958);
and UO_302 (O_302,N_2915,N_2991);
nor UO_303 (O_303,N_2900,N_2987);
or UO_304 (O_304,N_2935,N_2965);
and UO_305 (O_305,N_2933,N_2953);
nand UO_306 (O_306,N_2943,N_2937);
and UO_307 (O_307,N_2942,N_2993);
and UO_308 (O_308,N_2912,N_2964);
xnor UO_309 (O_309,N_2982,N_2971);
and UO_310 (O_310,N_2959,N_2929);
nand UO_311 (O_311,N_2932,N_2965);
nor UO_312 (O_312,N_2949,N_2910);
nor UO_313 (O_313,N_2982,N_2957);
and UO_314 (O_314,N_2919,N_2979);
and UO_315 (O_315,N_2911,N_2981);
or UO_316 (O_316,N_2963,N_2946);
and UO_317 (O_317,N_2916,N_2960);
or UO_318 (O_318,N_2935,N_2987);
or UO_319 (O_319,N_2955,N_2948);
or UO_320 (O_320,N_2960,N_2989);
and UO_321 (O_321,N_2978,N_2991);
or UO_322 (O_322,N_2910,N_2998);
or UO_323 (O_323,N_2916,N_2982);
and UO_324 (O_324,N_2906,N_2921);
nand UO_325 (O_325,N_2944,N_2920);
nor UO_326 (O_326,N_2914,N_2953);
nor UO_327 (O_327,N_2983,N_2944);
or UO_328 (O_328,N_2996,N_2919);
nand UO_329 (O_329,N_2909,N_2999);
nand UO_330 (O_330,N_2955,N_2915);
nor UO_331 (O_331,N_2928,N_2935);
and UO_332 (O_332,N_2979,N_2984);
and UO_333 (O_333,N_2988,N_2938);
nand UO_334 (O_334,N_2954,N_2962);
nand UO_335 (O_335,N_2994,N_2964);
and UO_336 (O_336,N_2931,N_2941);
nand UO_337 (O_337,N_2957,N_2997);
and UO_338 (O_338,N_2996,N_2974);
nand UO_339 (O_339,N_2918,N_2969);
nand UO_340 (O_340,N_2967,N_2915);
nand UO_341 (O_341,N_2912,N_2979);
nor UO_342 (O_342,N_2935,N_2921);
nand UO_343 (O_343,N_2942,N_2976);
and UO_344 (O_344,N_2944,N_2927);
nor UO_345 (O_345,N_2921,N_2963);
nand UO_346 (O_346,N_2982,N_2953);
and UO_347 (O_347,N_2971,N_2915);
nor UO_348 (O_348,N_2933,N_2962);
nor UO_349 (O_349,N_2968,N_2961);
or UO_350 (O_350,N_2947,N_2976);
or UO_351 (O_351,N_2979,N_2903);
or UO_352 (O_352,N_2979,N_2930);
nand UO_353 (O_353,N_2956,N_2986);
nor UO_354 (O_354,N_2915,N_2941);
or UO_355 (O_355,N_2974,N_2944);
and UO_356 (O_356,N_2960,N_2917);
nor UO_357 (O_357,N_2994,N_2985);
or UO_358 (O_358,N_2986,N_2940);
or UO_359 (O_359,N_2900,N_2956);
nor UO_360 (O_360,N_2993,N_2976);
and UO_361 (O_361,N_2962,N_2988);
nor UO_362 (O_362,N_2974,N_2976);
or UO_363 (O_363,N_2903,N_2976);
nor UO_364 (O_364,N_2967,N_2905);
and UO_365 (O_365,N_2961,N_2981);
nor UO_366 (O_366,N_2958,N_2933);
or UO_367 (O_367,N_2900,N_2924);
and UO_368 (O_368,N_2989,N_2955);
or UO_369 (O_369,N_2927,N_2917);
nand UO_370 (O_370,N_2967,N_2995);
nand UO_371 (O_371,N_2956,N_2919);
nand UO_372 (O_372,N_2920,N_2955);
or UO_373 (O_373,N_2954,N_2932);
nor UO_374 (O_374,N_2915,N_2962);
nor UO_375 (O_375,N_2998,N_2947);
nand UO_376 (O_376,N_2931,N_2954);
or UO_377 (O_377,N_2942,N_2929);
nor UO_378 (O_378,N_2968,N_2935);
or UO_379 (O_379,N_2938,N_2979);
nor UO_380 (O_380,N_2953,N_2947);
or UO_381 (O_381,N_2974,N_2909);
or UO_382 (O_382,N_2989,N_2920);
or UO_383 (O_383,N_2921,N_2942);
nor UO_384 (O_384,N_2963,N_2989);
or UO_385 (O_385,N_2900,N_2918);
nand UO_386 (O_386,N_2962,N_2995);
or UO_387 (O_387,N_2902,N_2936);
and UO_388 (O_388,N_2978,N_2903);
nand UO_389 (O_389,N_2961,N_2979);
and UO_390 (O_390,N_2924,N_2989);
nand UO_391 (O_391,N_2973,N_2941);
and UO_392 (O_392,N_2928,N_2948);
nor UO_393 (O_393,N_2956,N_2981);
or UO_394 (O_394,N_2933,N_2947);
nand UO_395 (O_395,N_2924,N_2968);
nor UO_396 (O_396,N_2970,N_2957);
and UO_397 (O_397,N_2940,N_2997);
and UO_398 (O_398,N_2969,N_2954);
and UO_399 (O_399,N_2949,N_2960);
nor UO_400 (O_400,N_2949,N_2930);
or UO_401 (O_401,N_2901,N_2943);
nand UO_402 (O_402,N_2910,N_2993);
or UO_403 (O_403,N_2960,N_2940);
and UO_404 (O_404,N_2925,N_2993);
nand UO_405 (O_405,N_2904,N_2900);
or UO_406 (O_406,N_2919,N_2980);
and UO_407 (O_407,N_2940,N_2991);
nor UO_408 (O_408,N_2936,N_2915);
and UO_409 (O_409,N_2917,N_2995);
or UO_410 (O_410,N_2997,N_2994);
and UO_411 (O_411,N_2958,N_2959);
nand UO_412 (O_412,N_2917,N_2925);
nor UO_413 (O_413,N_2908,N_2955);
nor UO_414 (O_414,N_2929,N_2989);
nand UO_415 (O_415,N_2936,N_2962);
and UO_416 (O_416,N_2999,N_2939);
nor UO_417 (O_417,N_2929,N_2966);
nor UO_418 (O_418,N_2907,N_2955);
nor UO_419 (O_419,N_2925,N_2948);
and UO_420 (O_420,N_2964,N_2956);
xnor UO_421 (O_421,N_2927,N_2961);
and UO_422 (O_422,N_2984,N_2970);
or UO_423 (O_423,N_2903,N_2922);
and UO_424 (O_424,N_2953,N_2917);
or UO_425 (O_425,N_2948,N_2972);
or UO_426 (O_426,N_2962,N_2927);
or UO_427 (O_427,N_2900,N_2902);
and UO_428 (O_428,N_2955,N_2963);
or UO_429 (O_429,N_2962,N_2913);
nor UO_430 (O_430,N_2951,N_2971);
or UO_431 (O_431,N_2908,N_2976);
nor UO_432 (O_432,N_2913,N_2998);
nand UO_433 (O_433,N_2932,N_2996);
or UO_434 (O_434,N_2967,N_2977);
nor UO_435 (O_435,N_2932,N_2959);
or UO_436 (O_436,N_2931,N_2947);
nor UO_437 (O_437,N_2953,N_2916);
nand UO_438 (O_438,N_2927,N_2919);
or UO_439 (O_439,N_2988,N_2942);
nand UO_440 (O_440,N_2939,N_2984);
or UO_441 (O_441,N_2972,N_2915);
nor UO_442 (O_442,N_2921,N_2934);
nor UO_443 (O_443,N_2946,N_2975);
nor UO_444 (O_444,N_2996,N_2930);
nand UO_445 (O_445,N_2945,N_2946);
or UO_446 (O_446,N_2970,N_2949);
and UO_447 (O_447,N_2991,N_2935);
nor UO_448 (O_448,N_2957,N_2992);
nor UO_449 (O_449,N_2993,N_2956);
and UO_450 (O_450,N_2973,N_2923);
nand UO_451 (O_451,N_2961,N_2942);
nor UO_452 (O_452,N_2943,N_2929);
nor UO_453 (O_453,N_2991,N_2921);
nand UO_454 (O_454,N_2934,N_2909);
or UO_455 (O_455,N_2981,N_2974);
nor UO_456 (O_456,N_2911,N_2982);
and UO_457 (O_457,N_2995,N_2944);
or UO_458 (O_458,N_2905,N_2985);
nand UO_459 (O_459,N_2992,N_2930);
or UO_460 (O_460,N_2939,N_2951);
nand UO_461 (O_461,N_2940,N_2999);
or UO_462 (O_462,N_2992,N_2953);
nand UO_463 (O_463,N_2966,N_2994);
and UO_464 (O_464,N_2932,N_2915);
and UO_465 (O_465,N_2960,N_2919);
or UO_466 (O_466,N_2958,N_2949);
or UO_467 (O_467,N_2959,N_2907);
or UO_468 (O_468,N_2965,N_2938);
nand UO_469 (O_469,N_2952,N_2981);
nor UO_470 (O_470,N_2927,N_2999);
nor UO_471 (O_471,N_2955,N_2959);
or UO_472 (O_472,N_2911,N_2953);
nand UO_473 (O_473,N_2913,N_2979);
or UO_474 (O_474,N_2985,N_2966);
nand UO_475 (O_475,N_2981,N_2903);
and UO_476 (O_476,N_2973,N_2926);
or UO_477 (O_477,N_2915,N_2954);
nand UO_478 (O_478,N_2906,N_2962);
nand UO_479 (O_479,N_2972,N_2975);
and UO_480 (O_480,N_2913,N_2959);
and UO_481 (O_481,N_2901,N_2970);
nand UO_482 (O_482,N_2901,N_2980);
or UO_483 (O_483,N_2982,N_2912);
nor UO_484 (O_484,N_2947,N_2984);
or UO_485 (O_485,N_2996,N_2976);
nand UO_486 (O_486,N_2981,N_2973);
and UO_487 (O_487,N_2940,N_2953);
nand UO_488 (O_488,N_2959,N_2925);
and UO_489 (O_489,N_2941,N_2974);
nand UO_490 (O_490,N_2948,N_2906);
or UO_491 (O_491,N_2912,N_2906);
and UO_492 (O_492,N_2990,N_2997);
nor UO_493 (O_493,N_2914,N_2992);
nor UO_494 (O_494,N_2976,N_2964);
and UO_495 (O_495,N_2929,N_2981);
nand UO_496 (O_496,N_2916,N_2920);
nor UO_497 (O_497,N_2931,N_2922);
or UO_498 (O_498,N_2958,N_2991);
nor UO_499 (O_499,N_2995,N_2971);
endmodule