module basic_500_3000_500_15_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_209,In_435);
nand U1 (N_1,In_470,In_412);
and U2 (N_2,In_87,In_193);
nand U3 (N_3,In_111,In_490);
nor U4 (N_4,In_370,In_171);
xnor U5 (N_5,In_186,In_420);
and U6 (N_6,In_141,In_244);
and U7 (N_7,In_16,In_320);
and U8 (N_8,In_20,In_97);
or U9 (N_9,In_486,In_433);
and U10 (N_10,In_173,In_31);
and U11 (N_11,In_450,In_15);
nand U12 (N_12,In_1,In_63);
nand U13 (N_13,In_106,In_135);
nor U14 (N_14,In_424,In_116);
and U15 (N_15,In_322,In_198);
nor U16 (N_16,In_384,In_45);
nor U17 (N_17,In_401,In_461);
and U18 (N_18,In_453,In_476);
nor U19 (N_19,In_249,In_441);
nand U20 (N_20,In_254,In_361);
nand U21 (N_21,In_301,In_287);
and U22 (N_22,In_324,In_313);
and U23 (N_23,In_346,In_274);
or U24 (N_24,In_245,In_76);
or U25 (N_25,In_277,In_146);
or U26 (N_26,In_165,In_280);
and U27 (N_27,In_419,In_284);
xnor U28 (N_28,In_493,In_91);
and U29 (N_29,In_283,In_119);
nand U30 (N_30,In_404,In_495);
nand U31 (N_31,In_491,In_93);
and U32 (N_32,In_469,In_482);
and U33 (N_33,In_43,In_485);
xnor U34 (N_34,In_72,In_204);
nor U35 (N_35,In_243,In_224);
and U36 (N_36,In_481,In_202);
xor U37 (N_37,In_457,In_19);
nor U38 (N_38,In_148,In_201);
nor U39 (N_39,In_238,In_108);
and U40 (N_40,In_377,In_321);
xnor U41 (N_41,In_257,In_154);
nor U42 (N_42,In_157,In_304);
and U43 (N_43,In_9,In_8);
and U44 (N_44,In_403,In_308);
nand U45 (N_45,In_399,In_475);
or U46 (N_46,In_300,In_84);
nand U47 (N_47,In_162,In_311);
and U48 (N_48,In_442,In_121);
and U49 (N_49,In_278,In_235);
nand U50 (N_50,In_448,In_328);
xnor U51 (N_51,In_139,In_223);
nor U52 (N_52,In_2,In_232);
or U53 (N_53,In_179,In_264);
nor U54 (N_54,In_151,In_187);
nor U55 (N_55,In_100,In_434);
or U56 (N_56,In_48,In_215);
nand U57 (N_57,In_85,In_68);
and U58 (N_58,In_227,In_89);
or U59 (N_59,In_14,In_467);
or U60 (N_60,In_26,In_423);
or U61 (N_61,In_6,In_410);
or U62 (N_62,In_71,In_340);
nor U63 (N_63,In_118,In_153);
nand U64 (N_64,In_364,In_421);
xor U65 (N_65,In_487,In_293);
nand U66 (N_66,In_234,In_360);
and U67 (N_67,In_488,In_443);
nand U68 (N_68,In_152,In_25);
nor U69 (N_69,In_417,In_411);
nor U70 (N_70,In_222,In_42);
and U71 (N_71,In_144,In_37);
xor U72 (N_72,In_58,In_344);
nand U73 (N_73,In_194,In_120);
or U74 (N_74,In_303,In_176);
or U75 (N_75,In_266,In_70);
and U76 (N_76,In_431,In_381);
or U77 (N_77,In_167,In_459);
nor U78 (N_78,In_241,In_53);
or U79 (N_79,In_110,In_231);
nor U80 (N_80,In_281,In_83);
nor U81 (N_81,In_21,In_253);
or U82 (N_82,In_279,In_126);
nand U83 (N_83,In_200,In_355);
nor U84 (N_84,In_378,In_214);
nor U85 (N_85,In_294,In_269);
and U86 (N_86,In_192,In_226);
nand U87 (N_87,In_79,In_205);
nor U88 (N_88,In_199,In_51);
or U89 (N_89,In_368,In_145);
nor U90 (N_90,In_50,In_77);
nor U91 (N_91,In_466,In_337);
nor U92 (N_92,In_317,In_455);
and U93 (N_93,In_221,In_252);
or U94 (N_94,In_286,In_142);
nor U95 (N_95,In_181,In_216);
or U96 (N_96,In_312,In_349);
nand U97 (N_97,In_496,In_465);
nor U98 (N_98,In_212,In_195);
or U99 (N_99,In_497,In_477);
and U100 (N_100,In_418,In_177);
nand U101 (N_101,In_348,In_471);
nor U102 (N_102,In_445,In_363);
and U103 (N_103,In_73,In_247);
nor U104 (N_104,In_333,In_124);
nor U105 (N_105,In_452,In_136);
nand U106 (N_106,In_271,In_387);
or U107 (N_107,In_75,In_468);
nand U108 (N_108,In_408,In_196);
and U109 (N_109,In_104,In_327);
nor U110 (N_110,In_422,In_65);
and U111 (N_111,In_147,In_62);
or U112 (N_112,In_81,In_331);
nor U113 (N_113,In_400,In_382);
nor U114 (N_114,In_66,In_402);
nor U115 (N_115,In_90,In_407);
nor U116 (N_116,In_207,In_432);
or U117 (N_117,In_131,In_449);
nand U118 (N_118,In_54,In_391);
or U119 (N_119,In_49,In_163);
nand U120 (N_120,In_101,In_127);
nand U121 (N_121,In_78,In_7);
or U122 (N_122,In_454,In_107);
and U123 (N_123,In_390,In_309);
nand U124 (N_124,In_140,In_319);
xnor U125 (N_125,In_255,In_260);
xor U126 (N_126,In_413,In_36);
nor U127 (N_127,In_302,In_12);
or U128 (N_128,In_392,In_183);
and U129 (N_129,In_463,In_158);
xnor U130 (N_130,In_5,In_270);
or U131 (N_131,In_155,In_64);
or U132 (N_132,In_123,In_296);
nor U133 (N_133,In_341,In_102);
nor U134 (N_134,In_330,In_233);
or U135 (N_135,In_460,In_347);
nand U136 (N_136,In_426,In_394);
and U137 (N_137,In_88,In_335);
and U138 (N_138,In_429,In_356);
and U139 (N_139,In_427,In_203);
or U140 (N_140,In_362,In_61);
nor U141 (N_141,In_342,In_57);
or U142 (N_142,In_11,In_275);
or U143 (N_143,In_109,In_166);
xnor U144 (N_144,In_210,In_339);
and U145 (N_145,In_354,In_440);
nor U146 (N_146,In_56,In_18);
nor U147 (N_147,In_369,In_30);
and U148 (N_148,In_32,In_379);
nand U149 (N_149,In_82,In_388);
nor U150 (N_150,In_246,In_197);
nor U151 (N_151,In_132,In_383);
nor U152 (N_152,In_288,In_456);
or U153 (N_153,In_251,In_315);
or U154 (N_154,In_473,In_98);
nor U155 (N_155,In_365,In_17);
nor U156 (N_156,In_67,In_299);
nand U157 (N_157,In_112,In_229);
nand U158 (N_158,In_334,In_86);
nand U159 (N_159,In_351,In_310);
nand U160 (N_160,In_298,In_24);
nand U161 (N_161,In_272,In_405);
nor U162 (N_162,In_80,In_323);
nor U163 (N_163,In_41,In_306);
and U164 (N_164,In_150,In_230);
or U165 (N_165,In_28,In_137);
xor U166 (N_166,In_430,In_375);
xnor U167 (N_167,In_217,In_479);
nor U168 (N_168,In_184,In_444);
and U169 (N_169,In_397,In_389);
nand U170 (N_170,In_34,In_492);
nand U171 (N_171,In_396,In_265);
xnor U172 (N_172,In_462,In_451);
or U173 (N_173,In_4,In_114);
and U174 (N_174,In_74,In_291);
nor U175 (N_175,In_182,In_168);
or U176 (N_176,In_117,In_329);
nand U177 (N_177,In_414,In_99);
nor U178 (N_178,In_267,In_55);
nand U179 (N_179,In_297,In_325);
nand U180 (N_180,In_160,In_95);
or U181 (N_181,In_164,In_393);
nor U182 (N_182,In_425,In_372);
or U183 (N_183,In_416,In_484);
or U184 (N_184,In_289,In_92);
nand U185 (N_185,In_105,In_237);
xnor U186 (N_186,In_38,In_191);
nor U187 (N_187,In_458,In_464);
xnor U188 (N_188,In_133,In_13);
and U189 (N_189,In_336,In_395);
nor U190 (N_190,In_273,In_386);
nand U191 (N_191,In_366,In_268);
nand U192 (N_192,In_409,In_474);
or U193 (N_193,In_282,In_256);
xor U194 (N_194,In_263,In_236);
nand U195 (N_195,In_295,In_318);
nand U196 (N_196,In_258,In_22);
and U197 (N_197,In_175,In_447);
nor U198 (N_198,In_138,In_314);
or U199 (N_199,In_316,In_113);
or U200 (N_200,N_5,N_50);
or U201 (N_201,In_373,In_220);
xor U202 (N_202,N_57,In_40);
or U203 (N_203,N_1,N_108);
xor U204 (N_204,N_48,In_290);
nor U205 (N_205,N_112,N_47);
nand U206 (N_206,N_179,N_148);
or U207 (N_207,N_20,In_345);
or U208 (N_208,N_144,In_385);
nand U209 (N_209,N_107,N_152);
and U210 (N_210,In_489,N_58);
or U211 (N_211,In_0,N_147);
nor U212 (N_212,N_80,In_174);
nand U213 (N_213,In_326,N_167);
nand U214 (N_214,In_380,N_109);
or U215 (N_215,N_18,In_415);
nor U216 (N_216,In_27,N_99);
and U217 (N_217,N_46,In_338);
nor U218 (N_218,N_117,N_195);
nor U219 (N_219,In_499,N_188);
nor U220 (N_220,N_73,In_428);
xnor U221 (N_221,In_357,N_161);
or U222 (N_222,N_126,N_71);
nor U223 (N_223,N_75,N_180);
nand U224 (N_224,N_190,In_39);
nand U225 (N_225,In_498,N_116);
and U226 (N_226,In_218,N_61);
and U227 (N_227,In_161,N_173);
nor U228 (N_228,In_343,N_26);
or U229 (N_229,N_2,N_157);
and U230 (N_230,In_44,N_184);
or U231 (N_231,N_121,N_87);
or U232 (N_232,N_102,N_186);
nand U233 (N_233,N_177,N_191);
or U234 (N_234,In_398,In_494);
nand U235 (N_235,In_367,In_180);
xnor U236 (N_236,In_96,In_103);
and U237 (N_237,N_42,N_65);
or U238 (N_238,N_111,In_439);
or U239 (N_239,N_90,N_77);
nand U240 (N_240,In_47,N_96);
nor U241 (N_241,N_29,N_92);
nand U242 (N_242,N_131,N_54);
and U243 (N_243,N_113,N_67);
and U244 (N_244,N_123,In_305);
and U245 (N_245,N_56,N_151);
nand U246 (N_246,N_9,In_225);
and U247 (N_247,N_154,In_129);
xor U248 (N_248,In_115,In_262);
nand U249 (N_249,N_8,N_53);
xnor U250 (N_250,N_6,In_228);
and U251 (N_251,In_33,N_66);
or U252 (N_252,N_181,N_27);
or U253 (N_253,In_29,In_248);
or U254 (N_254,In_35,In_10);
nor U255 (N_255,N_31,N_85);
xor U256 (N_256,N_10,N_72);
nand U257 (N_257,N_150,N_91);
xor U258 (N_258,N_159,N_63);
or U259 (N_259,N_21,N_138);
nand U260 (N_260,In_156,N_17);
nand U261 (N_261,N_15,In_59);
nor U262 (N_262,In_406,In_376);
and U263 (N_263,N_70,In_446);
and U264 (N_264,In_170,In_332);
xnor U265 (N_265,In_438,N_133);
nand U266 (N_266,In_69,N_0);
nand U267 (N_267,In_437,In_353);
or U268 (N_268,In_134,In_94);
nor U269 (N_269,N_139,In_125);
nand U270 (N_270,In_276,N_187);
nand U271 (N_271,In_242,In_159);
nor U272 (N_272,In_60,N_3);
or U273 (N_273,In_208,N_143);
nor U274 (N_274,N_88,In_350);
and U275 (N_275,N_127,N_45);
and U276 (N_276,N_97,N_120);
or U277 (N_277,N_162,In_178);
nand U278 (N_278,In_436,N_104);
nand U279 (N_279,N_52,N_101);
and U280 (N_280,N_94,N_93);
nor U281 (N_281,In_250,In_188);
or U282 (N_282,N_158,N_124);
and U283 (N_283,In_480,N_4);
nor U284 (N_284,N_137,N_193);
nand U285 (N_285,In_190,N_37);
nand U286 (N_286,N_16,N_134);
or U287 (N_287,N_197,In_359);
nand U288 (N_288,N_164,N_106);
or U289 (N_289,In_211,In_46);
nor U290 (N_290,In_239,N_156);
nor U291 (N_291,N_49,N_60);
and U292 (N_292,N_178,N_122);
nor U293 (N_293,In_219,N_160);
or U294 (N_294,N_136,N_55);
nand U295 (N_295,N_141,In_130);
or U296 (N_296,N_78,N_149);
or U297 (N_297,In_213,In_52);
and U298 (N_298,N_25,N_125);
or U299 (N_299,N_74,N_189);
xnor U300 (N_300,N_155,N_79);
nor U301 (N_301,In_189,N_33);
and U302 (N_302,N_142,N_100);
xnor U303 (N_303,N_36,N_198);
and U304 (N_304,N_185,N_69);
xor U305 (N_305,N_43,In_472);
nand U306 (N_306,N_114,N_38);
nor U307 (N_307,N_170,N_98);
nor U308 (N_308,N_23,N_140);
nor U309 (N_309,N_172,N_129);
nand U310 (N_310,N_196,In_122);
or U311 (N_311,In_358,N_30);
nand U312 (N_312,N_68,N_110);
nand U313 (N_313,N_59,In_172);
xnor U314 (N_314,N_103,N_168);
or U315 (N_315,N_34,N_130);
nor U316 (N_316,N_119,In_23);
or U317 (N_317,In_185,N_44);
xor U318 (N_318,N_13,N_28);
nand U319 (N_319,N_82,N_199);
nor U320 (N_320,In_128,N_183);
and U321 (N_321,N_135,N_22);
or U322 (N_322,N_165,N_86);
nand U323 (N_323,N_64,N_163);
or U324 (N_324,N_39,In_478);
nor U325 (N_325,N_118,N_182);
nor U326 (N_326,N_62,N_171);
and U327 (N_327,N_174,N_12);
nand U328 (N_328,In_352,N_41);
or U329 (N_329,In_374,N_19);
and U330 (N_330,In_483,N_35);
or U331 (N_331,N_175,N_51);
nand U332 (N_332,N_76,N_14);
and U333 (N_333,In_240,N_95);
xor U334 (N_334,N_166,In_261);
or U335 (N_335,In_371,N_81);
nand U336 (N_336,N_146,In_206);
nor U337 (N_337,N_11,In_149);
and U338 (N_338,In_292,N_115);
nor U339 (N_339,N_24,N_192);
and U340 (N_340,N_83,N_84);
and U341 (N_341,In_307,N_105);
and U342 (N_342,In_259,In_285);
nand U343 (N_343,N_132,N_40);
or U344 (N_344,N_153,N_169);
and U345 (N_345,N_89,In_3);
or U346 (N_346,In_143,N_32);
nor U347 (N_347,N_176,N_7);
nor U348 (N_348,In_169,N_145);
or U349 (N_349,N_194,N_128);
or U350 (N_350,In_436,N_167);
nor U351 (N_351,In_498,N_139);
or U352 (N_352,N_177,In_33);
xnor U353 (N_353,In_415,In_134);
xnor U354 (N_354,In_406,N_63);
nor U355 (N_355,N_176,In_211);
nand U356 (N_356,N_36,N_26);
or U357 (N_357,N_160,In_161);
nand U358 (N_358,N_176,N_95);
or U359 (N_359,N_31,N_71);
nor U360 (N_360,N_189,In_189);
and U361 (N_361,N_71,N_120);
and U362 (N_362,In_10,N_133);
nand U363 (N_363,N_110,In_46);
nor U364 (N_364,N_65,In_262);
nor U365 (N_365,In_218,N_97);
nand U366 (N_366,N_117,In_188);
and U367 (N_367,N_139,In_250);
nand U368 (N_368,N_76,In_446);
and U369 (N_369,In_343,N_77);
and U370 (N_370,N_155,N_25);
xnor U371 (N_371,N_95,N_195);
and U372 (N_372,N_44,N_103);
and U373 (N_373,N_146,N_50);
or U374 (N_374,N_36,In_371);
nor U375 (N_375,N_52,N_176);
and U376 (N_376,In_305,In_39);
nor U377 (N_377,N_136,N_4);
and U378 (N_378,In_446,N_147);
or U379 (N_379,N_165,N_178);
or U380 (N_380,N_136,In_307);
or U381 (N_381,N_154,N_85);
and U382 (N_382,N_164,N_3);
nand U383 (N_383,In_239,N_168);
nor U384 (N_384,N_166,In_206);
nand U385 (N_385,N_170,N_162);
and U386 (N_386,N_159,In_47);
nand U387 (N_387,N_87,N_141);
or U388 (N_388,In_115,N_155);
nand U389 (N_389,N_51,In_292);
nand U390 (N_390,N_51,N_12);
or U391 (N_391,In_242,N_2);
or U392 (N_392,N_112,In_446);
and U393 (N_393,N_85,In_149);
nand U394 (N_394,In_103,N_190);
or U395 (N_395,N_25,In_40);
or U396 (N_396,N_126,N_66);
xnor U397 (N_397,N_43,In_188);
nand U398 (N_398,N_194,N_58);
nand U399 (N_399,N_80,N_64);
and U400 (N_400,N_204,N_222);
nor U401 (N_401,N_203,N_280);
nor U402 (N_402,N_304,N_374);
xor U403 (N_403,N_309,N_265);
and U404 (N_404,N_334,N_209);
nor U405 (N_405,N_393,N_207);
nand U406 (N_406,N_262,N_398);
and U407 (N_407,N_353,N_223);
or U408 (N_408,N_298,N_357);
or U409 (N_409,N_384,N_253);
nor U410 (N_410,N_258,N_279);
nand U411 (N_411,N_387,N_231);
nor U412 (N_412,N_243,N_274);
or U413 (N_413,N_269,N_261);
nand U414 (N_414,N_399,N_378);
or U415 (N_415,N_317,N_234);
and U416 (N_416,N_268,N_368);
nand U417 (N_417,N_342,N_263);
and U418 (N_418,N_328,N_305);
and U419 (N_419,N_282,N_318);
and U420 (N_420,N_381,N_330);
and U421 (N_421,N_360,N_335);
nand U422 (N_422,N_237,N_362);
xnor U423 (N_423,N_386,N_345);
nor U424 (N_424,N_300,N_213);
nand U425 (N_425,N_316,N_354);
or U426 (N_426,N_296,N_249);
xnor U427 (N_427,N_264,N_214);
and U428 (N_428,N_232,N_240);
and U429 (N_429,N_370,N_239);
and U430 (N_430,N_329,N_247);
and U431 (N_431,N_392,N_211);
and U432 (N_432,N_358,N_217);
and U433 (N_433,N_385,N_397);
nor U434 (N_434,N_238,N_229);
and U435 (N_435,N_333,N_337);
nand U436 (N_436,N_295,N_285);
or U437 (N_437,N_355,N_291);
and U438 (N_438,N_272,N_289);
nor U439 (N_439,N_287,N_369);
xor U440 (N_440,N_202,N_270);
or U441 (N_441,N_303,N_308);
nor U442 (N_442,N_340,N_230);
and U443 (N_443,N_312,N_299);
or U444 (N_444,N_341,N_383);
or U445 (N_445,N_395,N_332);
xor U446 (N_446,N_376,N_322);
nor U447 (N_447,N_248,N_306);
and U448 (N_448,N_215,N_396);
and U449 (N_449,N_201,N_377);
nand U450 (N_450,N_361,N_365);
or U451 (N_451,N_391,N_311);
xnor U452 (N_452,N_244,N_346);
xnor U453 (N_453,N_338,N_284);
nand U454 (N_454,N_228,N_323);
or U455 (N_455,N_283,N_206);
or U456 (N_456,N_275,N_389);
nand U457 (N_457,N_326,N_200);
and U458 (N_458,N_367,N_325);
nand U459 (N_459,N_260,N_321);
nor U460 (N_460,N_221,N_314);
xor U461 (N_461,N_273,N_351);
nor U462 (N_462,N_349,N_315);
nor U463 (N_463,N_208,N_220);
nand U464 (N_464,N_366,N_218);
nand U465 (N_465,N_290,N_266);
and U466 (N_466,N_259,N_292);
nand U467 (N_467,N_394,N_388);
nand U468 (N_468,N_327,N_297);
nor U469 (N_469,N_294,N_278);
or U470 (N_470,N_271,N_359);
nand U471 (N_471,N_255,N_252);
nand U472 (N_472,N_319,N_233);
and U473 (N_473,N_331,N_372);
and U474 (N_474,N_236,N_224);
nand U475 (N_475,N_286,N_216);
and U476 (N_476,N_226,N_241);
and U477 (N_477,N_277,N_373);
nand U478 (N_478,N_254,N_288);
and U479 (N_479,N_371,N_281);
or U480 (N_480,N_205,N_352);
nand U481 (N_481,N_364,N_344);
or U482 (N_482,N_380,N_225);
and U483 (N_483,N_210,N_250);
or U484 (N_484,N_382,N_293);
nand U485 (N_485,N_320,N_276);
nor U486 (N_486,N_356,N_242);
nand U487 (N_487,N_348,N_336);
nor U488 (N_488,N_256,N_379);
or U489 (N_489,N_301,N_307);
nand U490 (N_490,N_347,N_219);
or U491 (N_491,N_313,N_246);
xor U492 (N_492,N_302,N_363);
nor U493 (N_493,N_227,N_339);
or U494 (N_494,N_390,N_257);
and U495 (N_495,N_350,N_245);
xor U496 (N_496,N_310,N_324);
nor U497 (N_497,N_212,N_343);
and U498 (N_498,N_251,N_267);
and U499 (N_499,N_235,N_375);
nor U500 (N_500,N_394,N_212);
nand U501 (N_501,N_269,N_313);
nor U502 (N_502,N_345,N_396);
nand U503 (N_503,N_206,N_305);
and U504 (N_504,N_395,N_251);
or U505 (N_505,N_241,N_311);
nor U506 (N_506,N_212,N_376);
xor U507 (N_507,N_306,N_376);
nand U508 (N_508,N_377,N_295);
xor U509 (N_509,N_361,N_346);
or U510 (N_510,N_249,N_258);
xnor U511 (N_511,N_239,N_330);
xnor U512 (N_512,N_263,N_367);
and U513 (N_513,N_325,N_265);
and U514 (N_514,N_325,N_342);
nand U515 (N_515,N_340,N_392);
or U516 (N_516,N_314,N_319);
and U517 (N_517,N_252,N_228);
nor U518 (N_518,N_258,N_228);
nand U519 (N_519,N_352,N_259);
nor U520 (N_520,N_382,N_304);
nor U521 (N_521,N_284,N_300);
nor U522 (N_522,N_298,N_257);
or U523 (N_523,N_252,N_279);
or U524 (N_524,N_324,N_224);
or U525 (N_525,N_250,N_304);
and U526 (N_526,N_387,N_377);
xnor U527 (N_527,N_306,N_340);
or U528 (N_528,N_322,N_229);
or U529 (N_529,N_276,N_282);
nand U530 (N_530,N_212,N_292);
and U531 (N_531,N_350,N_365);
or U532 (N_532,N_385,N_324);
nor U533 (N_533,N_259,N_277);
nand U534 (N_534,N_277,N_331);
nor U535 (N_535,N_252,N_207);
nor U536 (N_536,N_369,N_290);
nor U537 (N_537,N_214,N_332);
nor U538 (N_538,N_291,N_383);
nor U539 (N_539,N_336,N_366);
or U540 (N_540,N_345,N_218);
nor U541 (N_541,N_314,N_250);
or U542 (N_542,N_393,N_318);
nor U543 (N_543,N_393,N_309);
nor U544 (N_544,N_268,N_260);
or U545 (N_545,N_278,N_260);
nor U546 (N_546,N_390,N_282);
or U547 (N_547,N_264,N_385);
and U548 (N_548,N_396,N_305);
xor U549 (N_549,N_367,N_397);
and U550 (N_550,N_339,N_214);
and U551 (N_551,N_208,N_352);
or U552 (N_552,N_373,N_236);
xnor U553 (N_553,N_393,N_372);
xnor U554 (N_554,N_382,N_208);
nand U555 (N_555,N_325,N_344);
and U556 (N_556,N_325,N_388);
or U557 (N_557,N_248,N_347);
or U558 (N_558,N_249,N_267);
nand U559 (N_559,N_309,N_304);
and U560 (N_560,N_353,N_327);
xor U561 (N_561,N_257,N_231);
nand U562 (N_562,N_261,N_371);
or U563 (N_563,N_332,N_262);
xor U564 (N_564,N_238,N_273);
nor U565 (N_565,N_345,N_210);
nand U566 (N_566,N_381,N_396);
and U567 (N_567,N_253,N_335);
nand U568 (N_568,N_229,N_319);
nor U569 (N_569,N_388,N_314);
nand U570 (N_570,N_335,N_370);
nor U571 (N_571,N_357,N_220);
xnor U572 (N_572,N_240,N_239);
or U573 (N_573,N_390,N_320);
or U574 (N_574,N_358,N_268);
or U575 (N_575,N_346,N_252);
and U576 (N_576,N_350,N_324);
nor U577 (N_577,N_242,N_228);
nor U578 (N_578,N_316,N_265);
or U579 (N_579,N_367,N_225);
xnor U580 (N_580,N_235,N_209);
nand U581 (N_581,N_240,N_291);
xor U582 (N_582,N_327,N_239);
nand U583 (N_583,N_223,N_389);
nand U584 (N_584,N_346,N_366);
or U585 (N_585,N_379,N_230);
or U586 (N_586,N_362,N_345);
and U587 (N_587,N_310,N_209);
and U588 (N_588,N_351,N_243);
nor U589 (N_589,N_234,N_368);
xnor U590 (N_590,N_272,N_201);
nor U591 (N_591,N_263,N_229);
nor U592 (N_592,N_398,N_348);
or U593 (N_593,N_339,N_213);
nand U594 (N_594,N_337,N_279);
nor U595 (N_595,N_313,N_204);
or U596 (N_596,N_240,N_325);
and U597 (N_597,N_350,N_280);
and U598 (N_598,N_364,N_278);
nand U599 (N_599,N_333,N_334);
or U600 (N_600,N_428,N_526);
or U601 (N_601,N_542,N_481);
nand U602 (N_602,N_544,N_420);
xor U603 (N_603,N_437,N_495);
xnor U604 (N_604,N_571,N_511);
nand U605 (N_605,N_440,N_510);
nor U606 (N_606,N_546,N_450);
and U607 (N_607,N_489,N_592);
or U608 (N_608,N_568,N_549);
or U609 (N_609,N_468,N_446);
and U610 (N_610,N_404,N_453);
nand U611 (N_611,N_537,N_541);
nand U612 (N_612,N_540,N_506);
nand U613 (N_613,N_552,N_553);
nand U614 (N_614,N_480,N_458);
nand U615 (N_615,N_569,N_425);
and U616 (N_616,N_461,N_423);
or U617 (N_617,N_536,N_454);
nand U618 (N_618,N_561,N_488);
and U619 (N_619,N_523,N_421);
and U620 (N_620,N_572,N_433);
or U621 (N_621,N_528,N_470);
nand U622 (N_622,N_424,N_431);
nand U623 (N_623,N_460,N_406);
nand U624 (N_624,N_427,N_560);
nor U625 (N_625,N_533,N_418);
nor U626 (N_626,N_584,N_547);
and U627 (N_627,N_492,N_591);
or U628 (N_628,N_535,N_430);
xor U629 (N_629,N_409,N_442);
and U630 (N_630,N_590,N_550);
nand U631 (N_631,N_410,N_513);
and U632 (N_632,N_583,N_527);
nand U633 (N_633,N_518,N_562);
nor U634 (N_634,N_557,N_529);
xor U635 (N_635,N_509,N_574);
nor U636 (N_636,N_575,N_497);
nor U637 (N_637,N_545,N_429);
or U638 (N_638,N_556,N_416);
and U639 (N_639,N_465,N_567);
or U640 (N_640,N_548,N_448);
or U641 (N_641,N_598,N_405);
or U642 (N_642,N_554,N_525);
nor U643 (N_643,N_555,N_414);
xor U644 (N_644,N_474,N_594);
or U645 (N_645,N_596,N_482);
nor U646 (N_646,N_563,N_459);
and U647 (N_647,N_463,N_490);
nand U648 (N_648,N_508,N_499);
or U649 (N_649,N_521,N_524);
nor U650 (N_650,N_595,N_504);
nand U651 (N_651,N_500,N_402);
nand U652 (N_652,N_576,N_415);
xnor U653 (N_653,N_444,N_407);
nor U654 (N_654,N_457,N_438);
nor U655 (N_655,N_538,N_515);
or U656 (N_656,N_441,N_447);
xnor U657 (N_657,N_426,N_534);
nand U658 (N_658,N_516,N_413);
nor U659 (N_659,N_466,N_519);
nand U660 (N_660,N_597,N_491);
nor U661 (N_661,N_445,N_493);
or U662 (N_662,N_539,N_588);
or U663 (N_663,N_517,N_434);
or U664 (N_664,N_475,N_455);
xnor U665 (N_665,N_530,N_581);
nor U666 (N_666,N_471,N_412);
nand U667 (N_667,N_585,N_520);
nand U668 (N_668,N_473,N_559);
or U669 (N_669,N_472,N_551);
nand U670 (N_670,N_401,N_512);
and U671 (N_671,N_400,N_467);
nand U672 (N_672,N_570,N_496);
or U673 (N_673,N_531,N_514);
and U674 (N_674,N_579,N_505);
nor U675 (N_675,N_589,N_478);
nor U676 (N_676,N_435,N_593);
or U677 (N_677,N_494,N_578);
and U678 (N_678,N_487,N_469);
nor U679 (N_679,N_451,N_464);
or U680 (N_680,N_501,N_422);
nand U681 (N_681,N_449,N_443);
xor U682 (N_682,N_462,N_586);
nor U683 (N_683,N_439,N_483);
and U684 (N_684,N_452,N_477);
xnor U685 (N_685,N_507,N_417);
nand U686 (N_686,N_573,N_484);
or U687 (N_687,N_476,N_408);
nand U688 (N_688,N_479,N_543);
nor U689 (N_689,N_565,N_503);
nor U690 (N_690,N_564,N_587);
nand U691 (N_691,N_577,N_580);
nand U692 (N_692,N_522,N_566);
and U693 (N_693,N_419,N_432);
nor U694 (N_694,N_582,N_532);
nor U695 (N_695,N_485,N_436);
or U696 (N_696,N_403,N_599);
xnor U697 (N_697,N_456,N_558);
or U698 (N_698,N_498,N_502);
or U699 (N_699,N_411,N_486);
nor U700 (N_700,N_538,N_551);
and U701 (N_701,N_597,N_421);
and U702 (N_702,N_414,N_539);
nor U703 (N_703,N_499,N_419);
nand U704 (N_704,N_533,N_512);
nand U705 (N_705,N_463,N_565);
xnor U706 (N_706,N_483,N_433);
or U707 (N_707,N_571,N_472);
nor U708 (N_708,N_566,N_433);
nor U709 (N_709,N_546,N_488);
nor U710 (N_710,N_504,N_533);
nor U711 (N_711,N_473,N_470);
or U712 (N_712,N_411,N_551);
and U713 (N_713,N_498,N_493);
nand U714 (N_714,N_428,N_538);
nand U715 (N_715,N_495,N_519);
nor U716 (N_716,N_416,N_561);
and U717 (N_717,N_432,N_514);
nor U718 (N_718,N_401,N_425);
and U719 (N_719,N_432,N_473);
or U720 (N_720,N_441,N_548);
or U721 (N_721,N_474,N_576);
nand U722 (N_722,N_447,N_492);
xor U723 (N_723,N_554,N_418);
or U724 (N_724,N_478,N_567);
or U725 (N_725,N_420,N_428);
and U726 (N_726,N_457,N_532);
xor U727 (N_727,N_584,N_494);
and U728 (N_728,N_475,N_494);
nand U729 (N_729,N_580,N_568);
and U730 (N_730,N_470,N_550);
nor U731 (N_731,N_546,N_518);
and U732 (N_732,N_424,N_519);
or U733 (N_733,N_543,N_580);
xor U734 (N_734,N_599,N_589);
or U735 (N_735,N_471,N_401);
nand U736 (N_736,N_540,N_465);
and U737 (N_737,N_482,N_454);
or U738 (N_738,N_590,N_455);
and U739 (N_739,N_425,N_539);
and U740 (N_740,N_460,N_585);
xor U741 (N_741,N_516,N_595);
or U742 (N_742,N_420,N_504);
and U743 (N_743,N_588,N_501);
or U744 (N_744,N_468,N_421);
nand U745 (N_745,N_591,N_475);
nor U746 (N_746,N_432,N_575);
nand U747 (N_747,N_538,N_416);
nand U748 (N_748,N_514,N_590);
or U749 (N_749,N_508,N_464);
and U750 (N_750,N_549,N_463);
or U751 (N_751,N_584,N_524);
nand U752 (N_752,N_434,N_506);
and U753 (N_753,N_413,N_568);
and U754 (N_754,N_534,N_505);
nand U755 (N_755,N_526,N_536);
nor U756 (N_756,N_596,N_583);
or U757 (N_757,N_494,N_480);
nor U758 (N_758,N_477,N_475);
nor U759 (N_759,N_588,N_571);
nand U760 (N_760,N_416,N_478);
xnor U761 (N_761,N_592,N_507);
and U762 (N_762,N_428,N_573);
and U763 (N_763,N_462,N_452);
nor U764 (N_764,N_460,N_441);
or U765 (N_765,N_499,N_423);
xor U766 (N_766,N_404,N_533);
nand U767 (N_767,N_479,N_437);
xnor U768 (N_768,N_533,N_491);
nor U769 (N_769,N_473,N_444);
nor U770 (N_770,N_515,N_547);
xnor U771 (N_771,N_556,N_436);
or U772 (N_772,N_484,N_544);
nand U773 (N_773,N_447,N_533);
nand U774 (N_774,N_418,N_525);
nand U775 (N_775,N_514,N_549);
nor U776 (N_776,N_400,N_416);
nor U777 (N_777,N_470,N_543);
and U778 (N_778,N_482,N_426);
nand U779 (N_779,N_440,N_469);
nor U780 (N_780,N_572,N_523);
nand U781 (N_781,N_440,N_566);
nand U782 (N_782,N_556,N_400);
and U783 (N_783,N_584,N_510);
and U784 (N_784,N_556,N_419);
nor U785 (N_785,N_560,N_595);
nor U786 (N_786,N_520,N_588);
and U787 (N_787,N_583,N_494);
and U788 (N_788,N_569,N_410);
nor U789 (N_789,N_453,N_457);
nor U790 (N_790,N_562,N_458);
or U791 (N_791,N_488,N_423);
and U792 (N_792,N_448,N_442);
xor U793 (N_793,N_568,N_491);
or U794 (N_794,N_465,N_420);
nand U795 (N_795,N_513,N_558);
or U796 (N_796,N_552,N_500);
xor U797 (N_797,N_471,N_433);
or U798 (N_798,N_505,N_529);
nand U799 (N_799,N_560,N_542);
or U800 (N_800,N_730,N_799);
nor U801 (N_801,N_685,N_793);
nor U802 (N_802,N_625,N_798);
nand U803 (N_803,N_621,N_689);
and U804 (N_804,N_725,N_677);
or U805 (N_805,N_673,N_605);
nor U806 (N_806,N_781,N_687);
or U807 (N_807,N_751,N_622);
or U808 (N_808,N_679,N_702);
and U809 (N_809,N_697,N_768);
nand U810 (N_810,N_608,N_734);
nor U811 (N_811,N_766,N_646);
and U812 (N_812,N_660,N_795);
and U813 (N_813,N_729,N_669);
or U814 (N_814,N_694,N_645);
and U815 (N_815,N_770,N_789);
nand U816 (N_816,N_728,N_639);
nand U817 (N_817,N_736,N_754);
and U818 (N_818,N_632,N_790);
nor U819 (N_819,N_737,N_638);
and U820 (N_820,N_637,N_792);
and U821 (N_821,N_604,N_783);
and U822 (N_822,N_631,N_610);
or U823 (N_823,N_713,N_607);
and U824 (N_824,N_691,N_772);
or U825 (N_825,N_721,N_744);
nand U826 (N_826,N_603,N_714);
and U827 (N_827,N_726,N_747);
and U828 (N_828,N_735,N_708);
xnor U829 (N_829,N_627,N_650);
and U830 (N_830,N_620,N_681);
nand U831 (N_831,N_636,N_675);
and U832 (N_832,N_618,N_657);
nand U833 (N_833,N_743,N_680);
or U834 (N_834,N_753,N_665);
nand U835 (N_835,N_709,N_716);
nor U836 (N_836,N_676,N_794);
nand U837 (N_837,N_774,N_727);
or U838 (N_838,N_628,N_612);
nor U839 (N_839,N_600,N_630);
nor U840 (N_840,N_796,N_771);
nor U841 (N_841,N_769,N_760);
xor U842 (N_842,N_670,N_763);
or U843 (N_843,N_692,N_785);
nor U844 (N_844,N_649,N_664);
nor U845 (N_845,N_667,N_732);
or U846 (N_846,N_656,N_784);
nand U847 (N_847,N_663,N_723);
nand U848 (N_848,N_690,N_749);
nand U849 (N_849,N_658,N_672);
nor U850 (N_850,N_752,N_653);
and U851 (N_851,N_755,N_640);
or U852 (N_852,N_782,N_718);
or U853 (N_853,N_776,N_738);
or U854 (N_854,N_624,N_659);
and U855 (N_855,N_651,N_642);
and U856 (N_856,N_764,N_765);
nor U857 (N_857,N_750,N_602);
nand U858 (N_858,N_720,N_626);
and U859 (N_859,N_606,N_623);
nor U860 (N_860,N_775,N_715);
nor U861 (N_861,N_761,N_615);
and U862 (N_862,N_724,N_778);
xor U863 (N_863,N_731,N_787);
or U864 (N_864,N_683,N_698);
nor U865 (N_865,N_745,N_619);
and U866 (N_866,N_617,N_719);
and U867 (N_867,N_641,N_788);
xnor U868 (N_868,N_616,N_762);
and U869 (N_869,N_652,N_686);
or U870 (N_870,N_779,N_700);
xnor U871 (N_871,N_635,N_666);
xor U872 (N_872,N_759,N_647);
xnor U873 (N_873,N_654,N_678);
nand U874 (N_874,N_717,N_662);
and U875 (N_875,N_705,N_710);
nand U876 (N_876,N_739,N_701);
or U877 (N_877,N_741,N_614);
or U878 (N_878,N_711,N_671);
xnor U879 (N_879,N_633,N_742);
nand U880 (N_880,N_655,N_707);
xor U881 (N_881,N_757,N_722);
nand U882 (N_882,N_712,N_644);
nand U883 (N_883,N_746,N_634);
nand U884 (N_884,N_629,N_601);
xor U885 (N_885,N_693,N_611);
nor U886 (N_886,N_661,N_696);
and U887 (N_887,N_674,N_780);
nand U888 (N_888,N_609,N_773);
nor U889 (N_889,N_767,N_684);
nand U890 (N_890,N_703,N_791);
and U891 (N_891,N_695,N_777);
and U892 (N_892,N_613,N_758);
or U893 (N_893,N_688,N_733);
and U894 (N_894,N_699,N_682);
or U895 (N_895,N_648,N_756);
and U896 (N_896,N_748,N_740);
and U897 (N_897,N_797,N_668);
nor U898 (N_898,N_706,N_786);
nor U899 (N_899,N_643,N_704);
nand U900 (N_900,N_639,N_688);
and U901 (N_901,N_746,N_663);
or U902 (N_902,N_615,N_641);
nand U903 (N_903,N_698,N_721);
nor U904 (N_904,N_778,N_693);
or U905 (N_905,N_676,N_626);
nand U906 (N_906,N_748,N_725);
or U907 (N_907,N_741,N_650);
or U908 (N_908,N_783,N_772);
or U909 (N_909,N_683,N_607);
and U910 (N_910,N_687,N_618);
and U911 (N_911,N_789,N_646);
or U912 (N_912,N_745,N_618);
or U913 (N_913,N_662,N_652);
and U914 (N_914,N_664,N_602);
nand U915 (N_915,N_603,N_760);
nor U916 (N_916,N_736,N_689);
nand U917 (N_917,N_767,N_652);
and U918 (N_918,N_632,N_657);
xor U919 (N_919,N_605,N_774);
or U920 (N_920,N_664,N_612);
nor U921 (N_921,N_666,N_611);
xnor U922 (N_922,N_686,N_747);
nand U923 (N_923,N_736,N_681);
or U924 (N_924,N_683,N_668);
nor U925 (N_925,N_784,N_792);
nand U926 (N_926,N_734,N_765);
nand U927 (N_927,N_722,N_770);
and U928 (N_928,N_749,N_717);
nand U929 (N_929,N_714,N_757);
and U930 (N_930,N_715,N_690);
nor U931 (N_931,N_628,N_715);
nor U932 (N_932,N_778,N_716);
nor U933 (N_933,N_641,N_625);
nand U934 (N_934,N_643,N_600);
xnor U935 (N_935,N_640,N_703);
nand U936 (N_936,N_788,N_752);
and U937 (N_937,N_727,N_684);
nand U938 (N_938,N_631,N_697);
or U939 (N_939,N_656,N_603);
nand U940 (N_940,N_707,N_749);
nor U941 (N_941,N_773,N_746);
nand U942 (N_942,N_654,N_791);
and U943 (N_943,N_791,N_785);
nand U944 (N_944,N_790,N_608);
nor U945 (N_945,N_702,N_720);
xor U946 (N_946,N_673,N_760);
nor U947 (N_947,N_704,N_636);
or U948 (N_948,N_692,N_661);
or U949 (N_949,N_617,N_781);
or U950 (N_950,N_725,N_777);
nor U951 (N_951,N_658,N_713);
nor U952 (N_952,N_659,N_786);
or U953 (N_953,N_619,N_774);
nor U954 (N_954,N_664,N_606);
nor U955 (N_955,N_745,N_740);
or U956 (N_956,N_697,N_758);
xnor U957 (N_957,N_696,N_603);
or U958 (N_958,N_765,N_601);
and U959 (N_959,N_783,N_779);
nor U960 (N_960,N_629,N_645);
xnor U961 (N_961,N_689,N_799);
nor U962 (N_962,N_777,N_793);
nor U963 (N_963,N_619,N_760);
and U964 (N_964,N_678,N_618);
nand U965 (N_965,N_771,N_758);
or U966 (N_966,N_699,N_689);
nor U967 (N_967,N_791,N_761);
nor U968 (N_968,N_621,N_737);
or U969 (N_969,N_715,N_623);
nand U970 (N_970,N_615,N_645);
nor U971 (N_971,N_692,N_603);
nor U972 (N_972,N_635,N_647);
and U973 (N_973,N_734,N_761);
nand U974 (N_974,N_695,N_671);
nor U975 (N_975,N_783,N_726);
or U976 (N_976,N_623,N_683);
or U977 (N_977,N_664,N_670);
and U978 (N_978,N_723,N_626);
nor U979 (N_979,N_678,N_665);
nor U980 (N_980,N_709,N_670);
and U981 (N_981,N_686,N_785);
nand U982 (N_982,N_758,N_620);
nand U983 (N_983,N_700,N_727);
or U984 (N_984,N_739,N_748);
xor U985 (N_985,N_797,N_768);
or U986 (N_986,N_786,N_787);
and U987 (N_987,N_657,N_739);
and U988 (N_988,N_618,N_615);
or U989 (N_989,N_799,N_634);
nand U990 (N_990,N_655,N_777);
or U991 (N_991,N_660,N_615);
nand U992 (N_992,N_652,N_703);
nor U993 (N_993,N_784,N_699);
xnor U994 (N_994,N_602,N_639);
or U995 (N_995,N_605,N_701);
and U996 (N_996,N_787,N_626);
nand U997 (N_997,N_717,N_640);
nand U998 (N_998,N_738,N_775);
nand U999 (N_999,N_746,N_667);
nor U1000 (N_1000,N_947,N_922);
nor U1001 (N_1001,N_966,N_892);
nor U1002 (N_1002,N_965,N_817);
nor U1003 (N_1003,N_820,N_853);
nand U1004 (N_1004,N_992,N_878);
and U1005 (N_1005,N_875,N_864);
and U1006 (N_1006,N_842,N_818);
nand U1007 (N_1007,N_800,N_804);
nor U1008 (N_1008,N_995,N_830);
and U1009 (N_1009,N_928,N_975);
or U1010 (N_1010,N_998,N_913);
or U1011 (N_1011,N_857,N_968);
nor U1012 (N_1012,N_898,N_871);
nor U1013 (N_1013,N_921,N_969);
nand U1014 (N_1014,N_963,N_894);
xor U1015 (N_1015,N_930,N_927);
nor U1016 (N_1016,N_910,N_887);
nor U1017 (N_1017,N_891,N_845);
or U1018 (N_1018,N_955,N_885);
nor U1019 (N_1019,N_839,N_859);
xnor U1020 (N_1020,N_935,N_997);
nor U1021 (N_1021,N_941,N_999);
and U1022 (N_1022,N_843,N_976);
xor U1023 (N_1023,N_926,N_866);
and U1024 (N_1024,N_840,N_932);
nor U1025 (N_1025,N_942,N_906);
nor U1026 (N_1026,N_940,N_924);
nor U1027 (N_1027,N_879,N_987);
nor U1028 (N_1028,N_962,N_985);
xor U1029 (N_1029,N_849,N_824);
and U1030 (N_1030,N_972,N_909);
or U1031 (N_1031,N_893,N_851);
nand U1032 (N_1032,N_938,N_869);
or U1033 (N_1033,N_861,N_914);
nor U1034 (N_1034,N_990,N_948);
and U1035 (N_1035,N_929,N_946);
nor U1036 (N_1036,N_837,N_850);
or U1037 (N_1037,N_873,N_961);
or U1038 (N_1038,N_944,N_979);
nand U1039 (N_1039,N_970,N_958);
and U1040 (N_1040,N_826,N_952);
nand U1041 (N_1041,N_833,N_835);
or U1042 (N_1042,N_836,N_988);
nand U1043 (N_1043,N_899,N_986);
and U1044 (N_1044,N_889,N_828);
nand U1045 (N_1045,N_943,N_823);
or U1046 (N_1046,N_973,N_901);
or U1047 (N_1047,N_896,N_953);
or U1048 (N_1048,N_852,N_919);
nor U1049 (N_1049,N_862,N_888);
or U1050 (N_1050,N_980,N_829);
and U1051 (N_1051,N_874,N_827);
or U1052 (N_1052,N_960,N_884);
nand U1053 (N_1053,N_811,N_832);
or U1054 (N_1054,N_890,N_937);
nor U1055 (N_1055,N_847,N_814);
and U1056 (N_1056,N_971,N_933);
nand U1057 (N_1057,N_848,N_964);
xnor U1058 (N_1058,N_883,N_996);
nand U1059 (N_1059,N_865,N_900);
nor U1060 (N_1060,N_801,N_920);
or U1061 (N_1061,N_950,N_954);
nor U1062 (N_1062,N_974,N_802);
nand U1063 (N_1063,N_803,N_915);
nor U1064 (N_1064,N_905,N_831);
nand U1065 (N_1065,N_854,N_902);
nor U1066 (N_1066,N_816,N_880);
nand U1067 (N_1067,N_863,N_912);
nand U1068 (N_1068,N_925,N_834);
nor U1069 (N_1069,N_897,N_939);
nand U1070 (N_1070,N_978,N_807);
nand U1071 (N_1071,N_810,N_844);
and U1072 (N_1072,N_911,N_841);
or U1073 (N_1073,N_822,N_812);
nand U1074 (N_1074,N_918,N_886);
or U1075 (N_1075,N_959,N_945);
xnor U1076 (N_1076,N_882,N_956);
nand U1077 (N_1077,N_994,N_934);
or U1078 (N_1078,N_809,N_982);
or U1079 (N_1079,N_860,N_923);
or U1080 (N_1080,N_977,N_821);
or U1081 (N_1081,N_876,N_967);
and U1082 (N_1082,N_957,N_877);
xor U1083 (N_1083,N_858,N_819);
or U1084 (N_1084,N_989,N_936);
nand U1085 (N_1085,N_815,N_870);
nand U1086 (N_1086,N_903,N_806);
xnor U1087 (N_1087,N_904,N_917);
and U1088 (N_1088,N_855,N_808);
and U1089 (N_1089,N_951,N_907);
nand U1090 (N_1090,N_991,N_838);
xnor U1091 (N_1091,N_931,N_813);
and U1092 (N_1092,N_872,N_868);
nand U1093 (N_1093,N_993,N_856);
nor U1094 (N_1094,N_881,N_867);
or U1095 (N_1095,N_895,N_846);
and U1096 (N_1096,N_984,N_805);
nor U1097 (N_1097,N_908,N_983);
and U1098 (N_1098,N_916,N_981);
nand U1099 (N_1099,N_825,N_949);
and U1100 (N_1100,N_809,N_941);
nor U1101 (N_1101,N_864,N_845);
and U1102 (N_1102,N_850,N_921);
nor U1103 (N_1103,N_804,N_842);
and U1104 (N_1104,N_830,N_938);
nor U1105 (N_1105,N_854,N_838);
nor U1106 (N_1106,N_944,N_911);
nand U1107 (N_1107,N_879,N_882);
and U1108 (N_1108,N_852,N_875);
or U1109 (N_1109,N_989,N_806);
nand U1110 (N_1110,N_999,N_976);
nand U1111 (N_1111,N_963,N_981);
xnor U1112 (N_1112,N_803,N_910);
and U1113 (N_1113,N_870,N_939);
nor U1114 (N_1114,N_951,N_993);
nand U1115 (N_1115,N_985,N_848);
nor U1116 (N_1116,N_858,N_963);
or U1117 (N_1117,N_894,N_835);
and U1118 (N_1118,N_849,N_860);
nand U1119 (N_1119,N_852,N_944);
and U1120 (N_1120,N_815,N_882);
nand U1121 (N_1121,N_827,N_998);
or U1122 (N_1122,N_928,N_879);
nor U1123 (N_1123,N_964,N_842);
and U1124 (N_1124,N_813,N_926);
and U1125 (N_1125,N_814,N_878);
or U1126 (N_1126,N_941,N_995);
or U1127 (N_1127,N_871,N_996);
nor U1128 (N_1128,N_879,N_905);
or U1129 (N_1129,N_866,N_811);
nand U1130 (N_1130,N_931,N_889);
nand U1131 (N_1131,N_886,N_931);
and U1132 (N_1132,N_995,N_843);
or U1133 (N_1133,N_912,N_821);
nor U1134 (N_1134,N_980,N_938);
or U1135 (N_1135,N_911,N_913);
and U1136 (N_1136,N_921,N_882);
and U1137 (N_1137,N_987,N_906);
xnor U1138 (N_1138,N_892,N_993);
nor U1139 (N_1139,N_925,N_957);
xor U1140 (N_1140,N_899,N_945);
or U1141 (N_1141,N_927,N_850);
and U1142 (N_1142,N_931,N_976);
and U1143 (N_1143,N_939,N_800);
and U1144 (N_1144,N_802,N_986);
nor U1145 (N_1145,N_869,N_915);
or U1146 (N_1146,N_812,N_896);
nand U1147 (N_1147,N_837,N_947);
and U1148 (N_1148,N_826,N_869);
and U1149 (N_1149,N_885,N_941);
nor U1150 (N_1150,N_978,N_899);
and U1151 (N_1151,N_906,N_952);
and U1152 (N_1152,N_821,N_883);
nor U1153 (N_1153,N_961,N_848);
or U1154 (N_1154,N_885,N_873);
or U1155 (N_1155,N_904,N_908);
xnor U1156 (N_1156,N_964,N_863);
nor U1157 (N_1157,N_800,N_927);
nand U1158 (N_1158,N_834,N_993);
nor U1159 (N_1159,N_806,N_973);
and U1160 (N_1160,N_830,N_847);
nand U1161 (N_1161,N_987,N_845);
and U1162 (N_1162,N_860,N_835);
nor U1163 (N_1163,N_962,N_950);
nor U1164 (N_1164,N_953,N_843);
nand U1165 (N_1165,N_988,N_999);
or U1166 (N_1166,N_957,N_973);
nor U1167 (N_1167,N_844,N_819);
and U1168 (N_1168,N_831,N_931);
nand U1169 (N_1169,N_879,N_942);
nand U1170 (N_1170,N_984,N_827);
nand U1171 (N_1171,N_836,N_861);
or U1172 (N_1172,N_942,N_926);
nor U1173 (N_1173,N_829,N_805);
and U1174 (N_1174,N_989,N_934);
or U1175 (N_1175,N_850,N_923);
nor U1176 (N_1176,N_925,N_869);
or U1177 (N_1177,N_926,N_839);
or U1178 (N_1178,N_810,N_849);
or U1179 (N_1179,N_872,N_976);
nand U1180 (N_1180,N_886,N_917);
or U1181 (N_1181,N_937,N_941);
and U1182 (N_1182,N_990,N_944);
and U1183 (N_1183,N_852,N_840);
nor U1184 (N_1184,N_937,N_944);
and U1185 (N_1185,N_953,N_948);
or U1186 (N_1186,N_809,N_846);
nand U1187 (N_1187,N_801,N_883);
nor U1188 (N_1188,N_968,N_901);
or U1189 (N_1189,N_909,N_830);
nand U1190 (N_1190,N_830,N_841);
xor U1191 (N_1191,N_935,N_908);
and U1192 (N_1192,N_973,N_972);
or U1193 (N_1193,N_903,N_991);
and U1194 (N_1194,N_839,N_857);
or U1195 (N_1195,N_863,N_807);
nor U1196 (N_1196,N_903,N_945);
or U1197 (N_1197,N_956,N_868);
nor U1198 (N_1198,N_900,N_945);
and U1199 (N_1199,N_948,N_974);
nor U1200 (N_1200,N_1129,N_1160);
and U1201 (N_1201,N_1104,N_1062);
nand U1202 (N_1202,N_1007,N_1041);
nor U1203 (N_1203,N_1092,N_1055);
or U1204 (N_1204,N_1096,N_1037);
xnor U1205 (N_1205,N_1137,N_1027);
and U1206 (N_1206,N_1189,N_1122);
nor U1207 (N_1207,N_1118,N_1006);
nor U1208 (N_1208,N_1111,N_1143);
nor U1209 (N_1209,N_1176,N_1178);
xor U1210 (N_1210,N_1141,N_1126);
and U1211 (N_1211,N_1110,N_1063);
nor U1212 (N_1212,N_1073,N_1121);
xnor U1213 (N_1213,N_1167,N_1016);
nor U1214 (N_1214,N_1071,N_1149);
and U1215 (N_1215,N_1112,N_1172);
or U1216 (N_1216,N_1145,N_1010);
nor U1217 (N_1217,N_1087,N_1197);
and U1218 (N_1218,N_1161,N_1029);
xor U1219 (N_1219,N_1162,N_1072);
nor U1220 (N_1220,N_1101,N_1132);
or U1221 (N_1221,N_1181,N_1194);
nand U1222 (N_1222,N_1082,N_1198);
or U1223 (N_1223,N_1130,N_1075);
and U1224 (N_1224,N_1093,N_1183);
and U1225 (N_1225,N_1138,N_1155);
nand U1226 (N_1226,N_1025,N_1065);
nor U1227 (N_1227,N_1084,N_1020);
nor U1228 (N_1228,N_1159,N_1011);
and U1229 (N_1229,N_1128,N_1123);
xor U1230 (N_1230,N_1117,N_1085);
nor U1231 (N_1231,N_1195,N_1180);
xor U1232 (N_1232,N_1064,N_1100);
and U1233 (N_1233,N_1163,N_1186);
and U1234 (N_1234,N_1021,N_1050);
and U1235 (N_1235,N_1174,N_1151);
nand U1236 (N_1236,N_1142,N_1089);
or U1237 (N_1237,N_1033,N_1036);
nor U1238 (N_1238,N_1156,N_1177);
or U1239 (N_1239,N_1185,N_1059);
nand U1240 (N_1240,N_1135,N_1120);
or U1241 (N_1241,N_1031,N_1068);
or U1242 (N_1242,N_1106,N_1171);
and U1243 (N_1243,N_1049,N_1133);
and U1244 (N_1244,N_1125,N_1048);
nor U1245 (N_1245,N_1004,N_1045);
nor U1246 (N_1246,N_1191,N_1019);
or U1247 (N_1247,N_1067,N_1144);
and U1248 (N_1248,N_1192,N_1078);
or U1249 (N_1249,N_1146,N_1169);
xor U1250 (N_1250,N_1066,N_1152);
or U1251 (N_1251,N_1034,N_1001);
xor U1252 (N_1252,N_1090,N_1044);
or U1253 (N_1253,N_1088,N_1083);
nor U1254 (N_1254,N_1038,N_1051);
and U1255 (N_1255,N_1095,N_1168);
and U1256 (N_1256,N_1109,N_1052);
nor U1257 (N_1257,N_1103,N_1069);
nand U1258 (N_1258,N_1173,N_1182);
or U1259 (N_1259,N_1187,N_1000);
nor U1260 (N_1260,N_1165,N_1166);
or U1261 (N_1261,N_1193,N_1105);
nor U1262 (N_1262,N_1079,N_1077);
nand U1263 (N_1263,N_1074,N_1139);
nand U1264 (N_1264,N_1124,N_1008);
and U1265 (N_1265,N_1076,N_1119);
nor U1266 (N_1266,N_1115,N_1012);
and U1267 (N_1267,N_1184,N_1190);
nand U1268 (N_1268,N_1188,N_1170);
and U1269 (N_1269,N_1148,N_1153);
nand U1270 (N_1270,N_1042,N_1150);
xor U1271 (N_1271,N_1199,N_1017);
nor U1272 (N_1272,N_1023,N_1107);
and U1273 (N_1273,N_1081,N_1113);
nand U1274 (N_1274,N_1018,N_1058);
or U1275 (N_1275,N_1003,N_1039);
and U1276 (N_1276,N_1046,N_1099);
xor U1277 (N_1277,N_1005,N_1196);
nand U1278 (N_1278,N_1014,N_1022);
or U1279 (N_1279,N_1035,N_1056);
nor U1280 (N_1280,N_1009,N_1114);
or U1281 (N_1281,N_1030,N_1053);
nand U1282 (N_1282,N_1015,N_1097);
xor U1283 (N_1283,N_1013,N_1086);
or U1284 (N_1284,N_1043,N_1040);
nand U1285 (N_1285,N_1147,N_1154);
nor U1286 (N_1286,N_1164,N_1080);
and U1287 (N_1287,N_1057,N_1140);
nor U1288 (N_1288,N_1127,N_1175);
or U1289 (N_1289,N_1028,N_1026);
nor U1290 (N_1290,N_1070,N_1054);
nand U1291 (N_1291,N_1047,N_1098);
nand U1292 (N_1292,N_1131,N_1094);
or U1293 (N_1293,N_1024,N_1157);
xnor U1294 (N_1294,N_1032,N_1116);
nor U1295 (N_1295,N_1002,N_1136);
nand U1296 (N_1296,N_1158,N_1102);
nor U1297 (N_1297,N_1134,N_1108);
or U1298 (N_1298,N_1091,N_1061);
or U1299 (N_1299,N_1179,N_1060);
nand U1300 (N_1300,N_1153,N_1107);
nand U1301 (N_1301,N_1119,N_1148);
or U1302 (N_1302,N_1104,N_1056);
nor U1303 (N_1303,N_1134,N_1014);
and U1304 (N_1304,N_1079,N_1062);
and U1305 (N_1305,N_1075,N_1056);
nand U1306 (N_1306,N_1108,N_1115);
or U1307 (N_1307,N_1173,N_1091);
nand U1308 (N_1308,N_1170,N_1102);
nor U1309 (N_1309,N_1053,N_1075);
and U1310 (N_1310,N_1072,N_1061);
or U1311 (N_1311,N_1031,N_1188);
or U1312 (N_1312,N_1172,N_1168);
or U1313 (N_1313,N_1015,N_1119);
nand U1314 (N_1314,N_1044,N_1066);
nand U1315 (N_1315,N_1019,N_1193);
xnor U1316 (N_1316,N_1183,N_1159);
nor U1317 (N_1317,N_1101,N_1025);
or U1318 (N_1318,N_1032,N_1028);
and U1319 (N_1319,N_1106,N_1068);
or U1320 (N_1320,N_1002,N_1158);
nand U1321 (N_1321,N_1073,N_1188);
and U1322 (N_1322,N_1119,N_1009);
and U1323 (N_1323,N_1092,N_1041);
and U1324 (N_1324,N_1156,N_1055);
nor U1325 (N_1325,N_1133,N_1132);
nor U1326 (N_1326,N_1128,N_1065);
and U1327 (N_1327,N_1123,N_1108);
nor U1328 (N_1328,N_1084,N_1127);
or U1329 (N_1329,N_1125,N_1065);
nand U1330 (N_1330,N_1197,N_1139);
xnor U1331 (N_1331,N_1014,N_1034);
nor U1332 (N_1332,N_1186,N_1086);
nand U1333 (N_1333,N_1041,N_1033);
or U1334 (N_1334,N_1126,N_1111);
xor U1335 (N_1335,N_1077,N_1121);
nor U1336 (N_1336,N_1197,N_1186);
xnor U1337 (N_1337,N_1135,N_1098);
nor U1338 (N_1338,N_1159,N_1023);
and U1339 (N_1339,N_1030,N_1147);
and U1340 (N_1340,N_1017,N_1176);
or U1341 (N_1341,N_1098,N_1086);
nand U1342 (N_1342,N_1177,N_1180);
nand U1343 (N_1343,N_1176,N_1110);
nand U1344 (N_1344,N_1010,N_1018);
or U1345 (N_1345,N_1154,N_1160);
nand U1346 (N_1346,N_1125,N_1095);
and U1347 (N_1347,N_1171,N_1073);
or U1348 (N_1348,N_1136,N_1061);
and U1349 (N_1349,N_1083,N_1036);
xnor U1350 (N_1350,N_1053,N_1024);
or U1351 (N_1351,N_1079,N_1053);
and U1352 (N_1352,N_1052,N_1103);
or U1353 (N_1353,N_1167,N_1188);
nor U1354 (N_1354,N_1128,N_1172);
or U1355 (N_1355,N_1112,N_1093);
and U1356 (N_1356,N_1074,N_1066);
nor U1357 (N_1357,N_1153,N_1071);
nor U1358 (N_1358,N_1048,N_1016);
and U1359 (N_1359,N_1000,N_1194);
and U1360 (N_1360,N_1044,N_1184);
nor U1361 (N_1361,N_1024,N_1185);
xnor U1362 (N_1362,N_1007,N_1049);
nor U1363 (N_1363,N_1009,N_1140);
nor U1364 (N_1364,N_1102,N_1197);
xnor U1365 (N_1365,N_1086,N_1196);
or U1366 (N_1366,N_1004,N_1108);
xor U1367 (N_1367,N_1170,N_1000);
and U1368 (N_1368,N_1096,N_1115);
nor U1369 (N_1369,N_1135,N_1184);
or U1370 (N_1370,N_1191,N_1011);
and U1371 (N_1371,N_1097,N_1175);
nor U1372 (N_1372,N_1039,N_1007);
and U1373 (N_1373,N_1120,N_1007);
and U1374 (N_1374,N_1093,N_1193);
nand U1375 (N_1375,N_1015,N_1035);
nand U1376 (N_1376,N_1170,N_1149);
and U1377 (N_1377,N_1089,N_1049);
nand U1378 (N_1378,N_1166,N_1190);
nand U1379 (N_1379,N_1024,N_1115);
nor U1380 (N_1380,N_1065,N_1011);
and U1381 (N_1381,N_1020,N_1125);
nor U1382 (N_1382,N_1161,N_1009);
nor U1383 (N_1383,N_1116,N_1146);
and U1384 (N_1384,N_1122,N_1199);
or U1385 (N_1385,N_1043,N_1097);
xnor U1386 (N_1386,N_1112,N_1179);
and U1387 (N_1387,N_1165,N_1182);
or U1388 (N_1388,N_1007,N_1042);
nor U1389 (N_1389,N_1049,N_1073);
nand U1390 (N_1390,N_1119,N_1109);
nand U1391 (N_1391,N_1189,N_1118);
nor U1392 (N_1392,N_1197,N_1081);
nor U1393 (N_1393,N_1168,N_1013);
or U1394 (N_1394,N_1109,N_1190);
nor U1395 (N_1395,N_1188,N_1198);
nor U1396 (N_1396,N_1115,N_1022);
nor U1397 (N_1397,N_1085,N_1022);
or U1398 (N_1398,N_1095,N_1148);
or U1399 (N_1399,N_1165,N_1190);
nor U1400 (N_1400,N_1380,N_1320);
and U1401 (N_1401,N_1294,N_1267);
xor U1402 (N_1402,N_1384,N_1399);
nor U1403 (N_1403,N_1312,N_1393);
nand U1404 (N_1404,N_1271,N_1322);
or U1405 (N_1405,N_1369,N_1362);
or U1406 (N_1406,N_1217,N_1256);
nand U1407 (N_1407,N_1383,N_1232);
nor U1408 (N_1408,N_1261,N_1293);
xor U1409 (N_1409,N_1311,N_1325);
nand U1410 (N_1410,N_1373,N_1394);
nand U1411 (N_1411,N_1213,N_1389);
nand U1412 (N_1412,N_1370,N_1214);
and U1413 (N_1413,N_1318,N_1386);
nor U1414 (N_1414,N_1252,N_1249);
or U1415 (N_1415,N_1377,N_1228);
nand U1416 (N_1416,N_1255,N_1201);
nand U1417 (N_1417,N_1284,N_1301);
nand U1418 (N_1418,N_1203,N_1278);
nor U1419 (N_1419,N_1381,N_1305);
or U1420 (N_1420,N_1219,N_1210);
nand U1421 (N_1421,N_1266,N_1371);
nand U1422 (N_1422,N_1275,N_1287);
nor U1423 (N_1423,N_1243,N_1296);
or U1424 (N_1424,N_1215,N_1257);
or U1425 (N_1425,N_1277,N_1200);
nand U1426 (N_1426,N_1248,N_1388);
nand U1427 (N_1427,N_1205,N_1341);
nor U1428 (N_1428,N_1326,N_1361);
and U1429 (N_1429,N_1364,N_1289);
or U1430 (N_1430,N_1340,N_1374);
and U1431 (N_1431,N_1307,N_1390);
nand U1432 (N_1432,N_1297,N_1242);
xnor U1433 (N_1433,N_1358,N_1366);
nor U1434 (N_1434,N_1387,N_1230);
xor U1435 (N_1435,N_1259,N_1339);
and U1436 (N_1436,N_1246,N_1223);
nand U1437 (N_1437,N_1265,N_1395);
or U1438 (N_1438,N_1206,N_1338);
nor U1439 (N_1439,N_1220,N_1329);
nand U1440 (N_1440,N_1222,N_1349);
nor U1441 (N_1441,N_1333,N_1335);
nand U1442 (N_1442,N_1221,N_1225);
nor U1443 (N_1443,N_1254,N_1292);
and U1444 (N_1444,N_1218,N_1226);
nor U1445 (N_1445,N_1342,N_1309);
nor U1446 (N_1446,N_1283,N_1273);
or U1447 (N_1447,N_1328,N_1264);
xnor U1448 (N_1448,N_1291,N_1212);
and U1449 (N_1449,N_1321,N_1298);
and U1450 (N_1450,N_1348,N_1306);
nand U1451 (N_1451,N_1233,N_1238);
nor U1452 (N_1452,N_1279,N_1343);
and U1453 (N_1453,N_1241,N_1344);
or U1454 (N_1454,N_1351,N_1208);
nor U1455 (N_1455,N_1211,N_1276);
or U1456 (N_1456,N_1216,N_1270);
and U1457 (N_1457,N_1202,N_1239);
nand U1458 (N_1458,N_1245,N_1357);
or U1459 (N_1459,N_1355,N_1227);
and U1460 (N_1460,N_1234,N_1288);
and U1461 (N_1461,N_1237,N_1286);
or U1462 (N_1462,N_1379,N_1365);
nand U1463 (N_1463,N_1314,N_1398);
nand U1464 (N_1464,N_1319,N_1354);
nand U1465 (N_1465,N_1352,N_1209);
and U1466 (N_1466,N_1235,N_1269);
nand U1467 (N_1467,N_1290,N_1272);
nor U1468 (N_1468,N_1385,N_1375);
nand U1469 (N_1469,N_1300,N_1236);
or U1470 (N_1470,N_1397,N_1302);
and U1471 (N_1471,N_1347,N_1310);
xnor U1472 (N_1472,N_1372,N_1334);
xor U1473 (N_1473,N_1317,N_1244);
and U1474 (N_1474,N_1353,N_1376);
xnor U1475 (N_1475,N_1323,N_1240);
and U1476 (N_1476,N_1303,N_1345);
or U1477 (N_1477,N_1250,N_1396);
and U1478 (N_1478,N_1262,N_1324);
and U1479 (N_1479,N_1331,N_1327);
and U1480 (N_1480,N_1332,N_1392);
and U1481 (N_1481,N_1280,N_1336);
nand U1482 (N_1482,N_1391,N_1367);
or U1483 (N_1483,N_1282,N_1258);
nand U1484 (N_1484,N_1316,N_1281);
or U1485 (N_1485,N_1378,N_1315);
xnor U1486 (N_1486,N_1251,N_1274);
nand U1487 (N_1487,N_1346,N_1231);
or U1488 (N_1488,N_1304,N_1360);
or U1489 (N_1489,N_1268,N_1299);
and U1490 (N_1490,N_1337,N_1285);
xnor U1491 (N_1491,N_1308,N_1359);
or U1492 (N_1492,N_1207,N_1260);
and U1493 (N_1493,N_1356,N_1363);
nor U1494 (N_1494,N_1253,N_1368);
nor U1495 (N_1495,N_1204,N_1295);
nand U1496 (N_1496,N_1382,N_1330);
nand U1497 (N_1497,N_1247,N_1229);
or U1498 (N_1498,N_1263,N_1313);
or U1499 (N_1499,N_1350,N_1224);
and U1500 (N_1500,N_1241,N_1352);
and U1501 (N_1501,N_1231,N_1378);
nor U1502 (N_1502,N_1378,N_1262);
nand U1503 (N_1503,N_1396,N_1201);
xor U1504 (N_1504,N_1210,N_1251);
and U1505 (N_1505,N_1201,N_1308);
and U1506 (N_1506,N_1255,N_1244);
xor U1507 (N_1507,N_1382,N_1241);
nand U1508 (N_1508,N_1309,N_1373);
and U1509 (N_1509,N_1350,N_1204);
nor U1510 (N_1510,N_1347,N_1286);
nand U1511 (N_1511,N_1318,N_1205);
xnor U1512 (N_1512,N_1221,N_1222);
xnor U1513 (N_1513,N_1399,N_1274);
or U1514 (N_1514,N_1255,N_1378);
nand U1515 (N_1515,N_1266,N_1392);
and U1516 (N_1516,N_1265,N_1371);
or U1517 (N_1517,N_1355,N_1261);
and U1518 (N_1518,N_1242,N_1392);
and U1519 (N_1519,N_1215,N_1307);
nand U1520 (N_1520,N_1315,N_1252);
and U1521 (N_1521,N_1321,N_1344);
and U1522 (N_1522,N_1218,N_1381);
nor U1523 (N_1523,N_1257,N_1231);
and U1524 (N_1524,N_1317,N_1328);
or U1525 (N_1525,N_1249,N_1213);
nand U1526 (N_1526,N_1216,N_1313);
or U1527 (N_1527,N_1363,N_1370);
and U1528 (N_1528,N_1281,N_1341);
and U1529 (N_1529,N_1309,N_1266);
nand U1530 (N_1530,N_1337,N_1266);
nand U1531 (N_1531,N_1314,N_1263);
or U1532 (N_1532,N_1312,N_1338);
nand U1533 (N_1533,N_1363,N_1291);
and U1534 (N_1534,N_1285,N_1275);
nand U1535 (N_1535,N_1321,N_1324);
and U1536 (N_1536,N_1340,N_1228);
and U1537 (N_1537,N_1319,N_1231);
and U1538 (N_1538,N_1244,N_1265);
nand U1539 (N_1539,N_1244,N_1320);
and U1540 (N_1540,N_1347,N_1277);
and U1541 (N_1541,N_1250,N_1238);
and U1542 (N_1542,N_1386,N_1272);
nor U1543 (N_1543,N_1248,N_1267);
nand U1544 (N_1544,N_1368,N_1228);
nor U1545 (N_1545,N_1262,N_1373);
xor U1546 (N_1546,N_1289,N_1225);
and U1547 (N_1547,N_1347,N_1212);
or U1548 (N_1548,N_1338,N_1306);
or U1549 (N_1549,N_1362,N_1204);
and U1550 (N_1550,N_1399,N_1309);
nor U1551 (N_1551,N_1349,N_1337);
and U1552 (N_1552,N_1360,N_1397);
or U1553 (N_1553,N_1271,N_1254);
or U1554 (N_1554,N_1310,N_1384);
and U1555 (N_1555,N_1282,N_1379);
nand U1556 (N_1556,N_1323,N_1296);
and U1557 (N_1557,N_1382,N_1397);
or U1558 (N_1558,N_1343,N_1244);
or U1559 (N_1559,N_1242,N_1274);
and U1560 (N_1560,N_1303,N_1217);
nor U1561 (N_1561,N_1237,N_1334);
or U1562 (N_1562,N_1260,N_1369);
or U1563 (N_1563,N_1291,N_1241);
and U1564 (N_1564,N_1301,N_1269);
or U1565 (N_1565,N_1300,N_1233);
or U1566 (N_1566,N_1292,N_1280);
or U1567 (N_1567,N_1241,N_1201);
or U1568 (N_1568,N_1311,N_1249);
or U1569 (N_1569,N_1270,N_1218);
or U1570 (N_1570,N_1353,N_1364);
nor U1571 (N_1571,N_1385,N_1208);
or U1572 (N_1572,N_1214,N_1244);
nand U1573 (N_1573,N_1385,N_1364);
or U1574 (N_1574,N_1205,N_1229);
nor U1575 (N_1575,N_1242,N_1367);
nand U1576 (N_1576,N_1214,N_1315);
or U1577 (N_1577,N_1388,N_1263);
nand U1578 (N_1578,N_1267,N_1239);
xnor U1579 (N_1579,N_1352,N_1309);
or U1580 (N_1580,N_1331,N_1258);
nand U1581 (N_1581,N_1334,N_1296);
nor U1582 (N_1582,N_1303,N_1357);
nor U1583 (N_1583,N_1273,N_1382);
and U1584 (N_1584,N_1232,N_1280);
and U1585 (N_1585,N_1284,N_1348);
nand U1586 (N_1586,N_1351,N_1209);
nor U1587 (N_1587,N_1357,N_1387);
nor U1588 (N_1588,N_1398,N_1287);
and U1589 (N_1589,N_1355,N_1205);
or U1590 (N_1590,N_1284,N_1381);
nor U1591 (N_1591,N_1349,N_1202);
and U1592 (N_1592,N_1327,N_1200);
nor U1593 (N_1593,N_1316,N_1218);
and U1594 (N_1594,N_1284,N_1352);
nor U1595 (N_1595,N_1372,N_1201);
nor U1596 (N_1596,N_1350,N_1297);
nor U1597 (N_1597,N_1280,N_1356);
nor U1598 (N_1598,N_1288,N_1268);
or U1599 (N_1599,N_1365,N_1372);
nand U1600 (N_1600,N_1414,N_1546);
and U1601 (N_1601,N_1418,N_1486);
and U1602 (N_1602,N_1590,N_1447);
nor U1603 (N_1603,N_1407,N_1490);
or U1604 (N_1604,N_1599,N_1535);
nor U1605 (N_1605,N_1566,N_1503);
nor U1606 (N_1606,N_1428,N_1512);
xor U1607 (N_1607,N_1597,N_1579);
or U1608 (N_1608,N_1499,N_1526);
nor U1609 (N_1609,N_1523,N_1561);
or U1610 (N_1610,N_1554,N_1419);
and U1611 (N_1611,N_1400,N_1497);
or U1612 (N_1612,N_1464,N_1552);
nand U1613 (N_1613,N_1450,N_1459);
nor U1614 (N_1614,N_1514,N_1424);
or U1615 (N_1615,N_1462,N_1502);
nand U1616 (N_1616,N_1569,N_1433);
xnor U1617 (N_1617,N_1528,N_1427);
xor U1618 (N_1618,N_1513,N_1434);
nor U1619 (N_1619,N_1519,N_1417);
nor U1620 (N_1620,N_1518,N_1479);
nor U1621 (N_1621,N_1403,N_1507);
nand U1622 (N_1622,N_1422,N_1451);
xor U1623 (N_1623,N_1477,N_1525);
and U1624 (N_1624,N_1437,N_1409);
nand U1625 (N_1625,N_1574,N_1423);
nor U1626 (N_1626,N_1571,N_1556);
nand U1627 (N_1627,N_1544,N_1584);
nand U1628 (N_1628,N_1467,N_1588);
nand U1629 (N_1629,N_1402,N_1439);
nor U1630 (N_1630,N_1559,N_1530);
and U1631 (N_1631,N_1475,N_1411);
and U1632 (N_1632,N_1548,N_1442);
xnor U1633 (N_1633,N_1540,N_1468);
xor U1634 (N_1634,N_1443,N_1581);
nor U1635 (N_1635,N_1532,N_1465);
nor U1636 (N_1636,N_1553,N_1534);
nand U1637 (N_1637,N_1538,N_1496);
and U1638 (N_1638,N_1537,N_1586);
xnor U1639 (N_1639,N_1484,N_1458);
and U1640 (N_1640,N_1551,N_1408);
nand U1641 (N_1641,N_1539,N_1448);
or U1642 (N_1642,N_1598,N_1500);
or U1643 (N_1643,N_1431,N_1520);
nand U1644 (N_1644,N_1529,N_1406);
and U1645 (N_1645,N_1426,N_1436);
or U1646 (N_1646,N_1460,N_1470);
nor U1647 (N_1647,N_1515,N_1425);
or U1648 (N_1648,N_1405,N_1592);
and U1649 (N_1649,N_1582,N_1472);
and U1650 (N_1650,N_1541,N_1489);
xnor U1651 (N_1651,N_1488,N_1456);
nand U1652 (N_1652,N_1438,N_1570);
nor U1653 (N_1653,N_1522,N_1560);
or U1654 (N_1654,N_1483,N_1587);
and U1655 (N_1655,N_1536,N_1583);
nor U1656 (N_1656,N_1572,N_1412);
nand U1657 (N_1657,N_1567,N_1510);
and U1658 (N_1658,N_1430,N_1501);
or U1659 (N_1659,N_1481,N_1547);
or U1660 (N_1660,N_1454,N_1591);
or U1661 (N_1661,N_1533,N_1595);
nor U1662 (N_1662,N_1498,N_1485);
nand U1663 (N_1663,N_1446,N_1504);
or U1664 (N_1664,N_1480,N_1577);
and U1665 (N_1665,N_1463,N_1413);
nand U1666 (N_1666,N_1471,N_1473);
xnor U1667 (N_1667,N_1585,N_1404);
and U1668 (N_1668,N_1594,N_1568);
or U1669 (N_1669,N_1455,N_1492);
nand U1670 (N_1670,N_1573,N_1474);
or U1671 (N_1671,N_1495,N_1562);
nand U1672 (N_1672,N_1580,N_1478);
or U1673 (N_1673,N_1416,N_1415);
or U1674 (N_1674,N_1493,N_1543);
xnor U1675 (N_1675,N_1420,N_1593);
nor U1676 (N_1676,N_1457,N_1557);
nor U1677 (N_1677,N_1453,N_1527);
nand U1678 (N_1678,N_1509,N_1558);
nand U1679 (N_1679,N_1482,N_1441);
nor U1680 (N_1680,N_1516,N_1401);
or U1681 (N_1681,N_1508,N_1445);
or U1682 (N_1682,N_1511,N_1545);
nand U1683 (N_1683,N_1429,N_1596);
and U1684 (N_1684,N_1466,N_1549);
and U1685 (N_1685,N_1449,N_1589);
or U1686 (N_1686,N_1452,N_1578);
xnor U1687 (N_1687,N_1432,N_1421);
nand U1688 (N_1688,N_1505,N_1542);
nand U1689 (N_1689,N_1564,N_1555);
xor U1690 (N_1690,N_1521,N_1576);
and U1691 (N_1691,N_1487,N_1410);
xnor U1692 (N_1692,N_1517,N_1565);
nor U1693 (N_1693,N_1435,N_1461);
and U1694 (N_1694,N_1444,N_1563);
nand U1695 (N_1695,N_1440,N_1494);
nand U1696 (N_1696,N_1524,N_1531);
and U1697 (N_1697,N_1575,N_1476);
nor U1698 (N_1698,N_1469,N_1550);
or U1699 (N_1699,N_1506,N_1491);
and U1700 (N_1700,N_1553,N_1583);
nor U1701 (N_1701,N_1477,N_1474);
and U1702 (N_1702,N_1415,N_1467);
nor U1703 (N_1703,N_1403,N_1552);
and U1704 (N_1704,N_1430,N_1571);
nand U1705 (N_1705,N_1488,N_1528);
nor U1706 (N_1706,N_1560,N_1439);
and U1707 (N_1707,N_1560,N_1403);
xnor U1708 (N_1708,N_1456,N_1457);
nand U1709 (N_1709,N_1422,N_1529);
nor U1710 (N_1710,N_1400,N_1422);
nor U1711 (N_1711,N_1587,N_1454);
or U1712 (N_1712,N_1469,N_1437);
and U1713 (N_1713,N_1580,N_1472);
nand U1714 (N_1714,N_1449,N_1546);
and U1715 (N_1715,N_1561,N_1477);
nor U1716 (N_1716,N_1419,N_1450);
or U1717 (N_1717,N_1504,N_1435);
nor U1718 (N_1718,N_1589,N_1439);
and U1719 (N_1719,N_1492,N_1416);
xor U1720 (N_1720,N_1453,N_1587);
nor U1721 (N_1721,N_1490,N_1406);
and U1722 (N_1722,N_1585,N_1453);
xor U1723 (N_1723,N_1515,N_1482);
or U1724 (N_1724,N_1467,N_1560);
or U1725 (N_1725,N_1435,N_1462);
xnor U1726 (N_1726,N_1545,N_1553);
and U1727 (N_1727,N_1447,N_1461);
nand U1728 (N_1728,N_1458,N_1489);
nor U1729 (N_1729,N_1417,N_1571);
and U1730 (N_1730,N_1441,N_1454);
and U1731 (N_1731,N_1445,N_1482);
nor U1732 (N_1732,N_1539,N_1537);
and U1733 (N_1733,N_1403,N_1506);
nand U1734 (N_1734,N_1461,N_1547);
xor U1735 (N_1735,N_1433,N_1562);
nand U1736 (N_1736,N_1508,N_1585);
nand U1737 (N_1737,N_1476,N_1528);
and U1738 (N_1738,N_1475,N_1508);
and U1739 (N_1739,N_1550,N_1521);
nor U1740 (N_1740,N_1531,N_1508);
or U1741 (N_1741,N_1402,N_1526);
nand U1742 (N_1742,N_1531,N_1443);
or U1743 (N_1743,N_1442,N_1416);
and U1744 (N_1744,N_1542,N_1569);
nor U1745 (N_1745,N_1585,N_1496);
and U1746 (N_1746,N_1439,N_1408);
nand U1747 (N_1747,N_1492,N_1550);
and U1748 (N_1748,N_1458,N_1415);
nor U1749 (N_1749,N_1493,N_1429);
or U1750 (N_1750,N_1540,N_1534);
nand U1751 (N_1751,N_1444,N_1513);
and U1752 (N_1752,N_1574,N_1408);
and U1753 (N_1753,N_1502,N_1450);
or U1754 (N_1754,N_1567,N_1543);
nand U1755 (N_1755,N_1496,N_1415);
or U1756 (N_1756,N_1420,N_1491);
xor U1757 (N_1757,N_1503,N_1459);
nor U1758 (N_1758,N_1441,N_1422);
and U1759 (N_1759,N_1580,N_1513);
and U1760 (N_1760,N_1567,N_1430);
nor U1761 (N_1761,N_1557,N_1599);
nor U1762 (N_1762,N_1408,N_1545);
or U1763 (N_1763,N_1550,N_1584);
or U1764 (N_1764,N_1456,N_1573);
nor U1765 (N_1765,N_1482,N_1498);
nand U1766 (N_1766,N_1509,N_1560);
nor U1767 (N_1767,N_1491,N_1462);
nor U1768 (N_1768,N_1504,N_1513);
nand U1769 (N_1769,N_1580,N_1414);
or U1770 (N_1770,N_1542,N_1466);
nor U1771 (N_1771,N_1434,N_1550);
nor U1772 (N_1772,N_1572,N_1566);
xor U1773 (N_1773,N_1522,N_1570);
and U1774 (N_1774,N_1567,N_1492);
nand U1775 (N_1775,N_1461,N_1541);
nand U1776 (N_1776,N_1523,N_1509);
nor U1777 (N_1777,N_1556,N_1514);
and U1778 (N_1778,N_1441,N_1538);
nor U1779 (N_1779,N_1427,N_1517);
or U1780 (N_1780,N_1562,N_1540);
xor U1781 (N_1781,N_1577,N_1591);
nand U1782 (N_1782,N_1443,N_1518);
xnor U1783 (N_1783,N_1410,N_1567);
nor U1784 (N_1784,N_1500,N_1414);
xnor U1785 (N_1785,N_1515,N_1582);
xor U1786 (N_1786,N_1585,N_1560);
nand U1787 (N_1787,N_1504,N_1506);
or U1788 (N_1788,N_1519,N_1587);
or U1789 (N_1789,N_1542,N_1492);
nand U1790 (N_1790,N_1452,N_1514);
and U1791 (N_1791,N_1463,N_1582);
nand U1792 (N_1792,N_1483,N_1530);
xor U1793 (N_1793,N_1410,N_1596);
or U1794 (N_1794,N_1479,N_1580);
nand U1795 (N_1795,N_1402,N_1480);
nor U1796 (N_1796,N_1538,N_1587);
or U1797 (N_1797,N_1480,N_1584);
or U1798 (N_1798,N_1400,N_1434);
and U1799 (N_1799,N_1429,N_1438);
nor U1800 (N_1800,N_1712,N_1685);
or U1801 (N_1801,N_1680,N_1611);
and U1802 (N_1802,N_1700,N_1602);
and U1803 (N_1803,N_1672,N_1729);
nor U1804 (N_1804,N_1714,N_1688);
nor U1805 (N_1805,N_1662,N_1791);
xnor U1806 (N_1806,N_1728,N_1689);
or U1807 (N_1807,N_1620,N_1614);
nor U1808 (N_1808,N_1727,N_1656);
or U1809 (N_1809,N_1667,N_1780);
and U1810 (N_1810,N_1678,N_1610);
or U1811 (N_1811,N_1723,N_1710);
and U1812 (N_1812,N_1702,N_1642);
or U1813 (N_1813,N_1790,N_1601);
or U1814 (N_1814,N_1608,N_1766);
nor U1815 (N_1815,N_1600,N_1752);
or U1816 (N_1816,N_1622,N_1668);
xor U1817 (N_1817,N_1616,N_1634);
nor U1818 (N_1818,N_1701,N_1707);
or U1819 (N_1819,N_1736,N_1734);
nand U1820 (N_1820,N_1643,N_1756);
xor U1821 (N_1821,N_1648,N_1693);
and U1822 (N_1822,N_1740,N_1747);
and U1823 (N_1823,N_1695,N_1745);
nor U1824 (N_1824,N_1664,N_1730);
and U1825 (N_1825,N_1677,N_1794);
and U1826 (N_1826,N_1735,N_1731);
xnor U1827 (N_1827,N_1639,N_1606);
or U1828 (N_1828,N_1703,N_1787);
nand U1829 (N_1829,N_1719,N_1773);
nand U1830 (N_1830,N_1686,N_1632);
nand U1831 (N_1831,N_1673,N_1762);
and U1832 (N_1832,N_1647,N_1781);
nand U1833 (N_1833,N_1718,N_1690);
nor U1834 (N_1834,N_1692,N_1798);
and U1835 (N_1835,N_1792,N_1646);
nor U1836 (N_1836,N_1779,N_1774);
nor U1837 (N_1837,N_1708,N_1705);
xnor U1838 (N_1838,N_1706,N_1796);
nand U1839 (N_1839,N_1630,N_1759);
or U1840 (N_1840,N_1738,N_1741);
and U1841 (N_1841,N_1666,N_1783);
nand U1842 (N_1842,N_1755,N_1669);
or U1843 (N_1843,N_1742,N_1763);
or U1844 (N_1844,N_1627,N_1753);
nor U1845 (N_1845,N_1758,N_1623);
nand U1846 (N_1846,N_1699,N_1746);
nor U1847 (N_1847,N_1681,N_1644);
and U1848 (N_1848,N_1621,N_1604);
nor U1849 (N_1849,N_1612,N_1640);
and U1850 (N_1850,N_1785,N_1618);
nor U1851 (N_1851,N_1628,N_1613);
nand U1852 (N_1852,N_1776,N_1799);
nand U1853 (N_1853,N_1617,N_1754);
and U1854 (N_1854,N_1770,N_1625);
or U1855 (N_1855,N_1631,N_1637);
nand U1856 (N_1856,N_1725,N_1764);
or U1857 (N_1857,N_1657,N_1750);
nor U1858 (N_1858,N_1768,N_1733);
nor U1859 (N_1859,N_1769,N_1653);
xnor U1860 (N_1860,N_1713,N_1665);
nand U1861 (N_1861,N_1786,N_1715);
nand U1862 (N_1862,N_1603,N_1605);
and U1863 (N_1863,N_1626,N_1636);
and U1864 (N_1864,N_1615,N_1795);
and U1865 (N_1865,N_1743,N_1624);
nor U1866 (N_1866,N_1674,N_1697);
nand U1867 (N_1867,N_1749,N_1761);
nand U1868 (N_1868,N_1684,N_1757);
nand U1869 (N_1869,N_1760,N_1645);
and U1870 (N_1870,N_1651,N_1687);
nand U1871 (N_1871,N_1682,N_1732);
or U1872 (N_1872,N_1797,N_1691);
xnor U1873 (N_1873,N_1679,N_1619);
and U1874 (N_1874,N_1744,N_1661);
or U1875 (N_1875,N_1775,N_1654);
nand U1876 (N_1876,N_1777,N_1765);
nor U1877 (N_1877,N_1609,N_1683);
nand U1878 (N_1878,N_1771,N_1789);
and U1879 (N_1879,N_1670,N_1676);
nor U1880 (N_1880,N_1635,N_1629);
nand U1881 (N_1881,N_1767,N_1720);
nand U1882 (N_1882,N_1772,N_1782);
or U1883 (N_1883,N_1793,N_1694);
or U1884 (N_1884,N_1633,N_1739);
nand U1885 (N_1885,N_1641,N_1649);
nand U1886 (N_1886,N_1650,N_1709);
nand U1887 (N_1887,N_1737,N_1724);
or U1888 (N_1888,N_1721,N_1652);
or U1889 (N_1889,N_1607,N_1659);
or U1890 (N_1890,N_1660,N_1663);
and U1891 (N_1891,N_1716,N_1704);
nand U1892 (N_1892,N_1658,N_1711);
or U1893 (N_1893,N_1717,N_1726);
nor U1894 (N_1894,N_1784,N_1698);
and U1895 (N_1895,N_1748,N_1751);
or U1896 (N_1896,N_1696,N_1671);
nor U1897 (N_1897,N_1722,N_1788);
and U1898 (N_1898,N_1655,N_1675);
or U1899 (N_1899,N_1778,N_1638);
nor U1900 (N_1900,N_1692,N_1796);
nand U1901 (N_1901,N_1654,N_1688);
or U1902 (N_1902,N_1790,N_1710);
and U1903 (N_1903,N_1660,N_1647);
and U1904 (N_1904,N_1701,N_1760);
nand U1905 (N_1905,N_1659,N_1704);
or U1906 (N_1906,N_1700,N_1638);
and U1907 (N_1907,N_1663,N_1680);
nand U1908 (N_1908,N_1789,N_1751);
and U1909 (N_1909,N_1744,N_1673);
nor U1910 (N_1910,N_1656,N_1687);
and U1911 (N_1911,N_1792,N_1680);
nand U1912 (N_1912,N_1785,N_1637);
nand U1913 (N_1913,N_1672,N_1710);
nor U1914 (N_1914,N_1616,N_1775);
nor U1915 (N_1915,N_1708,N_1632);
xnor U1916 (N_1916,N_1650,N_1657);
nand U1917 (N_1917,N_1753,N_1775);
nand U1918 (N_1918,N_1779,N_1658);
nor U1919 (N_1919,N_1770,N_1664);
or U1920 (N_1920,N_1695,N_1682);
or U1921 (N_1921,N_1651,N_1767);
and U1922 (N_1922,N_1626,N_1752);
or U1923 (N_1923,N_1667,N_1729);
or U1924 (N_1924,N_1738,N_1689);
and U1925 (N_1925,N_1668,N_1695);
and U1926 (N_1926,N_1676,N_1681);
or U1927 (N_1927,N_1769,N_1618);
or U1928 (N_1928,N_1738,N_1760);
and U1929 (N_1929,N_1708,N_1653);
and U1930 (N_1930,N_1653,N_1685);
nand U1931 (N_1931,N_1790,N_1699);
and U1932 (N_1932,N_1715,N_1716);
nor U1933 (N_1933,N_1624,N_1771);
nand U1934 (N_1934,N_1707,N_1600);
nand U1935 (N_1935,N_1630,N_1699);
nand U1936 (N_1936,N_1640,N_1757);
nand U1937 (N_1937,N_1704,N_1782);
nor U1938 (N_1938,N_1752,N_1640);
nor U1939 (N_1939,N_1664,N_1639);
and U1940 (N_1940,N_1755,N_1651);
nand U1941 (N_1941,N_1755,N_1765);
xor U1942 (N_1942,N_1726,N_1706);
and U1943 (N_1943,N_1628,N_1747);
or U1944 (N_1944,N_1713,N_1642);
nor U1945 (N_1945,N_1753,N_1799);
xor U1946 (N_1946,N_1713,N_1721);
nor U1947 (N_1947,N_1698,N_1619);
nor U1948 (N_1948,N_1658,N_1661);
and U1949 (N_1949,N_1775,N_1670);
xnor U1950 (N_1950,N_1788,N_1798);
and U1951 (N_1951,N_1653,N_1661);
or U1952 (N_1952,N_1799,N_1700);
nand U1953 (N_1953,N_1659,N_1796);
nand U1954 (N_1954,N_1753,N_1738);
and U1955 (N_1955,N_1739,N_1799);
and U1956 (N_1956,N_1747,N_1618);
or U1957 (N_1957,N_1640,N_1670);
nand U1958 (N_1958,N_1628,N_1720);
nor U1959 (N_1959,N_1711,N_1769);
nand U1960 (N_1960,N_1684,N_1736);
nand U1961 (N_1961,N_1724,N_1615);
nand U1962 (N_1962,N_1654,N_1647);
nor U1963 (N_1963,N_1796,N_1684);
nor U1964 (N_1964,N_1764,N_1614);
nor U1965 (N_1965,N_1644,N_1791);
xor U1966 (N_1966,N_1625,N_1760);
or U1967 (N_1967,N_1642,N_1675);
or U1968 (N_1968,N_1778,N_1646);
nor U1969 (N_1969,N_1736,N_1757);
or U1970 (N_1970,N_1750,N_1605);
nor U1971 (N_1971,N_1718,N_1607);
and U1972 (N_1972,N_1609,N_1699);
nor U1973 (N_1973,N_1775,N_1689);
nor U1974 (N_1974,N_1774,N_1672);
and U1975 (N_1975,N_1658,N_1750);
and U1976 (N_1976,N_1687,N_1719);
xnor U1977 (N_1977,N_1633,N_1762);
nor U1978 (N_1978,N_1627,N_1691);
xor U1979 (N_1979,N_1681,N_1735);
xnor U1980 (N_1980,N_1603,N_1637);
and U1981 (N_1981,N_1716,N_1749);
nand U1982 (N_1982,N_1667,N_1617);
nand U1983 (N_1983,N_1770,N_1794);
and U1984 (N_1984,N_1700,N_1665);
nor U1985 (N_1985,N_1721,N_1671);
nand U1986 (N_1986,N_1654,N_1644);
and U1987 (N_1987,N_1668,N_1719);
nand U1988 (N_1988,N_1715,N_1612);
or U1989 (N_1989,N_1695,N_1754);
nand U1990 (N_1990,N_1615,N_1748);
and U1991 (N_1991,N_1646,N_1645);
or U1992 (N_1992,N_1771,N_1731);
and U1993 (N_1993,N_1782,N_1632);
and U1994 (N_1994,N_1604,N_1757);
or U1995 (N_1995,N_1700,N_1648);
nor U1996 (N_1996,N_1784,N_1749);
or U1997 (N_1997,N_1749,N_1620);
and U1998 (N_1998,N_1678,N_1674);
and U1999 (N_1999,N_1742,N_1609);
nor U2000 (N_2000,N_1879,N_1907);
or U2001 (N_2001,N_1980,N_1981);
and U2002 (N_2002,N_1903,N_1849);
nand U2003 (N_2003,N_1966,N_1833);
or U2004 (N_2004,N_1914,N_1825);
and U2005 (N_2005,N_1961,N_1979);
nor U2006 (N_2006,N_1852,N_1882);
or U2007 (N_2007,N_1856,N_1912);
nand U2008 (N_2008,N_1832,N_1843);
nor U2009 (N_2009,N_1908,N_1826);
nor U2010 (N_2010,N_1894,N_1904);
and U2011 (N_2011,N_1817,N_1801);
and U2012 (N_2012,N_1847,N_1804);
xor U2013 (N_2013,N_1997,N_1952);
nand U2014 (N_2014,N_1810,N_1866);
and U2015 (N_2015,N_1974,N_1800);
xor U2016 (N_2016,N_1870,N_1881);
xnor U2017 (N_2017,N_1965,N_1922);
nor U2018 (N_2018,N_1897,N_1996);
and U2019 (N_2019,N_1831,N_1850);
nor U2020 (N_2020,N_1948,N_1936);
and U2021 (N_2021,N_1943,N_1938);
or U2022 (N_2022,N_1932,N_1940);
and U2023 (N_2023,N_1975,N_1990);
nor U2024 (N_2024,N_1977,N_1900);
nor U2025 (N_2025,N_1955,N_1910);
and U2026 (N_2026,N_1830,N_1994);
nor U2027 (N_2027,N_1929,N_1877);
nor U2028 (N_2028,N_1998,N_1964);
nor U2029 (N_2029,N_1815,N_1916);
nor U2030 (N_2030,N_1814,N_1971);
nand U2031 (N_2031,N_1999,N_1803);
nor U2032 (N_2032,N_1919,N_1837);
or U2033 (N_2033,N_1845,N_1963);
or U2034 (N_2034,N_1834,N_1945);
and U2035 (N_2035,N_1973,N_1829);
nand U2036 (N_2036,N_1953,N_1868);
or U2037 (N_2037,N_1920,N_1958);
xor U2038 (N_2038,N_1935,N_1957);
nand U2039 (N_2039,N_1909,N_1836);
xnor U2040 (N_2040,N_1899,N_1853);
nand U2041 (N_2041,N_1988,N_1927);
nor U2042 (N_2042,N_1876,N_1923);
xnor U2043 (N_2043,N_1808,N_1861);
nor U2044 (N_2044,N_1928,N_1915);
nor U2045 (N_2045,N_1806,N_1887);
xor U2046 (N_2046,N_1802,N_1959);
nor U2047 (N_2047,N_1854,N_1895);
or U2048 (N_2048,N_1986,N_1993);
or U2049 (N_2049,N_1819,N_1872);
and U2050 (N_2050,N_1859,N_1931);
nand U2051 (N_2051,N_1883,N_1933);
and U2052 (N_2052,N_1946,N_1942);
or U2053 (N_2053,N_1823,N_1869);
nand U2054 (N_2054,N_1921,N_1969);
and U2055 (N_2055,N_1941,N_1867);
or U2056 (N_2056,N_1944,N_1820);
xnor U2057 (N_2057,N_1898,N_1924);
and U2058 (N_2058,N_1818,N_1913);
and U2059 (N_2059,N_1983,N_1937);
and U2060 (N_2060,N_1951,N_1805);
nand U2061 (N_2061,N_1930,N_1846);
nand U2062 (N_2062,N_1839,N_1934);
nor U2063 (N_2063,N_1809,N_1860);
xnor U2064 (N_2064,N_1967,N_1992);
and U2065 (N_2065,N_1811,N_1821);
xnor U2066 (N_2066,N_1890,N_1880);
and U2067 (N_2067,N_1851,N_1902);
or U2068 (N_2068,N_1970,N_1807);
nor U2069 (N_2069,N_1888,N_1989);
nor U2070 (N_2070,N_1855,N_1984);
or U2071 (N_2071,N_1835,N_1949);
nor U2072 (N_2072,N_1982,N_1873);
xor U2073 (N_2073,N_1862,N_1891);
nand U2074 (N_2074,N_1878,N_1842);
nand U2075 (N_2075,N_1885,N_1863);
xor U2076 (N_2076,N_1886,N_1812);
nand U2077 (N_2077,N_1871,N_1857);
nor U2078 (N_2078,N_1840,N_1906);
xor U2079 (N_2079,N_1917,N_1889);
and U2080 (N_2080,N_1874,N_1939);
or U2081 (N_2081,N_1968,N_1844);
nand U2082 (N_2082,N_1960,N_1858);
and U2083 (N_2083,N_1991,N_1925);
nor U2084 (N_2084,N_1978,N_1985);
or U2085 (N_2085,N_1841,N_1865);
nand U2086 (N_2086,N_1848,N_1893);
nor U2087 (N_2087,N_1947,N_1926);
or U2088 (N_2088,N_1954,N_1901);
nor U2089 (N_2089,N_1962,N_1827);
nor U2090 (N_2090,N_1864,N_1813);
and U2091 (N_2091,N_1918,N_1838);
and U2092 (N_2092,N_1892,N_1884);
nor U2093 (N_2093,N_1911,N_1822);
nor U2094 (N_2094,N_1976,N_1905);
nor U2095 (N_2095,N_1950,N_1987);
and U2096 (N_2096,N_1875,N_1816);
or U2097 (N_2097,N_1896,N_1828);
and U2098 (N_2098,N_1972,N_1956);
or U2099 (N_2099,N_1824,N_1995);
nor U2100 (N_2100,N_1833,N_1899);
nor U2101 (N_2101,N_1813,N_1861);
xnor U2102 (N_2102,N_1826,N_1871);
nand U2103 (N_2103,N_1930,N_1854);
and U2104 (N_2104,N_1869,N_1834);
or U2105 (N_2105,N_1848,N_1928);
and U2106 (N_2106,N_1952,N_1883);
nor U2107 (N_2107,N_1992,N_1970);
nor U2108 (N_2108,N_1959,N_1840);
nor U2109 (N_2109,N_1910,N_1883);
or U2110 (N_2110,N_1904,N_1820);
nor U2111 (N_2111,N_1886,N_1829);
or U2112 (N_2112,N_1911,N_1823);
or U2113 (N_2113,N_1833,N_1862);
or U2114 (N_2114,N_1803,N_1973);
nand U2115 (N_2115,N_1807,N_1814);
xor U2116 (N_2116,N_1817,N_1974);
xor U2117 (N_2117,N_1930,N_1843);
and U2118 (N_2118,N_1856,N_1971);
nand U2119 (N_2119,N_1860,N_1960);
nor U2120 (N_2120,N_1951,N_1935);
and U2121 (N_2121,N_1978,N_1896);
and U2122 (N_2122,N_1924,N_1911);
nor U2123 (N_2123,N_1915,N_1983);
and U2124 (N_2124,N_1901,N_1991);
and U2125 (N_2125,N_1946,N_1950);
nor U2126 (N_2126,N_1950,N_1804);
and U2127 (N_2127,N_1819,N_1805);
nor U2128 (N_2128,N_1898,N_1867);
nor U2129 (N_2129,N_1994,N_1876);
and U2130 (N_2130,N_1973,N_1933);
nand U2131 (N_2131,N_1932,N_1909);
and U2132 (N_2132,N_1947,N_1819);
nand U2133 (N_2133,N_1916,N_1920);
nand U2134 (N_2134,N_1834,N_1872);
and U2135 (N_2135,N_1806,N_1891);
or U2136 (N_2136,N_1891,N_1872);
nor U2137 (N_2137,N_1908,N_1972);
nand U2138 (N_2138,N_1849,N_1970);
or U2139 (N_2139,N_1887,N_1966);
nor U2140 (N_2140,N_1847,N_1914);
nand U2141 (N_2141,N_1879,N_1936);
nand U2142 (N_2142,N_1969,N_1927);
and U2143 (N_2143,N_1852,N_1821);
xor U2144 (N_2144,N_1930,N_1917);
or U2145 (N_2145,N_1889,N_1882);
xnor U2146 (N_2146,N_1884,N_1989);
nand U2147 (N_2147,N_1909,N_1859);
nand U2148 (N_2148,N_1987,N_1878);
and U2149 (N_2149,N_1937,N_1986);
or U2150 (N_2150,N_1966,N_1850);
and U2151 (N_2151,N_1886,N_1840);
or U2152 (N_2152,N_1844,N_1867);
and U2153 (N_2153,N_1876,N_1985);
nor U2154 (N_2154,N_1862,N_1844);
and U2155 (N_2155,N_1807,N_1927);
and U2156 (N_2156,N_1910,N_1808);
xnor U2157 (N_2157,N_1911,N_1887);
xnor U2158 (N_2158,N_1824,N_1815);
xor U2159 (N_2159,N_1918,N_1970);
nor U2160 (N_2160,N_1808,N_1906);
nand U2161 (N_2161,N_1939,N_1948);
or U2162 (N_2162,N_1969,N_1913);
xnor U2163 (N_2163,N_1873,N_1899);
or U2164 (N_2164,N_1937,N_1849);
and U2165 (N_2165,N_1982,N_1957);
nor U2166 (N_2166,N_1880,N_1921);
or U2167 (N_2167,N_1971,N_1886);
and U2168 (N_2168,N_1872,N_1807);
and U2169 (N_2169,N_1823,N_1815);
nor U2170 (N_2170,N_1912,N_1814);
nor U2171 (N_2171,N_1808,N_1938);
nand U2172 (N_2172,N_1997,N_1852);
nand U2173 (N_2173,N_1932,N_1964);
nor U2174 (N_2174,N_1829,N_1842);
nor U2175 (N_2175,N_1814,N_1990);
and U2176 (N_2176,N_1856,N_1882);
nor U2177 (N_2177,N_1945,N_1876);
nand U2178 (N_2178,N_1806,N_1923);
or U2179 (N_2179,N_1880,N_1898);
or U2180 (N_2180,N_1955,N_1862);
xnor U2181 (N_2181,N_1926,N_1964);
nand U2182 (N_2182,N_1889,N_1877);
or U2183 (N_2183,N_1923,N_1814);
nand U2184 (N_2184,N_1939,N_1867);
and U2185 (N_2185,N_1802,N_1948);
and U2186 (N_2186,N_1939,N_1877);
nor U2187 (N_2187,N_1852,N_1809);
nor U2188 (N_2188,N_1958,N_1895);
and U2189 (N_2189,N_1909,N_1808);
nor U2190 (N_2190,N_1805,N_1933);
nor U2191 (N_2191,N_1988,N_1808);
and U2192 (N_2192,N_1924,N_1854);
nor U2193 (N_2193,N_1812,N_1998);
and U2194 (N_2194,N_1926,N_1972);
and U2195 (N_2195,N_1961,N_1915);
nand U2196 (N_2196,N_1960,N_1935);
or U2197 (N_2197,N_1846,N_1958);
nand U2198 (N_2198,N_1993,N_1840);
or U2199 (N_2199,N_1963,N_1834);
xor U2200 (N_2200,N_2193,N_2076);
nand U2201 (N_2201,N_2088,N_2050);
nand U2202 (N_2202,N_2165,N_2077);
nor U2203 (N_2203,N_2096,N_2126);
xor U2204 (N_2204,N_2198,N_2093);
and U2205 (N_2205,N_2023,N_2079);
or U2206 (N_2206,N_2018,N_2045);
or U2207 (N_2207,N_2141,N_2176);
nand U2208 (N_2208,N_2075,N_2146);
nand U2209 (N_2209,N_2117,N_2154);
or U2210 (N_2210,N_2081,N_2190);
or U2211 (N_2211,N_2006,N_2056);
xnor U2212 (N_2212,N_2178,N_2001);
and U2213 (N_2213,N_2047,N_2175);
nor U2214 (N_2214,N_2010,N_2008);
nand U2215 (N_2215,N_2112,N_2014);
or U2216 (N_2216,N_2125,N_2149);
and U2217 (N_2217,N_2067,N_2105);
xor U2218 (N_2218,N_2034,N_2017);
and U2219 (N_2219,N_2061,N_2196);
nand U2220 (N_2220,N_2049,N_2156);
or U2221 (N_2221,N_2168,N_2054);
nor U2222 (N_2222,N_2015,N_2057);
or U2223 (N_2223,N_2084,N_2111);
and U2224 (N_2224,N_2072,N_2133);
nor U2225 (N_2225,N_2055,N_2065);
nor U2226 (N_2226,N_2058,N_2132);
nor U2227 (N_2227,N_2122,N_2129);
and U2228 (N_2228,N_2024,N_2043);
or U2229 (N_2229,N_2137,N_2027);
and U2230 (N_2230,N_2078,N_2103);
or U2231 (N_2231,N_2044,N_2127);
and U2232 (N_2232,N_2071,N_2036);
nand U2233 (N_2233,N_2091,N_2130);
or U2234 (N_2234,N_2086,N_2089);
and U2235 (N_2235,N_2134,N_2124);
xnor U2236 (N_2236,N_2032,N_2038);
nor U2237 (N_2237,N_2073,N_2094);
nor U2238 (N_2238,N_2082,N_2083);
and U2239 (N_2239,N_2119,N_2148);
or U2240 (N_2240,N_2114,N_2151);
nor U2241 (N_2241,N_2020,N_2025);
nor U2242 (N_2242,N_2185,N_2062);
or U2243 (N_2243,N_2157,N_2002);
and U2244 (N_2244,N_2192,N_2102);
or U2245 (N_2245,N_2195,N_2173);
or U2246 (N_2246,N_2187,N_2046);
nand U2247 (N_2247,N_2116,N_2182);
or U2248 (N_2248,N_2069,N_2121);
nand U2249 (N_2249,N_2120,N_2101);
nand U2250 (N_2250,N_2085,N_2042);
and U2251 (N_2251,N_2099,N_2090);
nand U2252 (N_2252,N_2033,N_2163);
nor U2253 (N_2253,N_2009,N_2186);
or U2254 (N_2254,N_2184,N_2109);
and U2255 (N_2255,N_2074,N_2092);
nor U2256 (N_2256,N_2097,N_2169);
xnor U2257 (N_2257,N_2098,N_2104);
nand U2258 (N_2258,N_2128,N_2022);
and U2259 (N_2259,N_2113,N_2164);
or U2260 (N_2260,N_2118,N_2011);
xor U2261 (N_2261,N_2030,N_2095);
nor U2262 (N_2262,N_2170,N_2189);
nand U2263 (N_2263,N_2140,N_2110);
nand U2264 (N_2264,N_2021,N_2037);
nor U2265 (N_2265,N_2035,N_2106);
nor U2266 (N_2266,N_2180,N_2166);
nand U2267 (N_2267,N_2108,N_2060);
and U2268 (N_2268,N_2161,N_2000);
nor U2269 (N_2269,N_2139,N_2158);
or U2270 (N_2270,N_2152,N_2028);
nand U2271 (N_2271,N_2145,N_2087);
or U2272 (N_2272,N_2142,N_2029);
or U2273 (N_2273,N_2153,N_2123);
nor U2274 (N_2274,N_2188,N_2026);
and U2275 (N_2275,N_2174,N_2031);
or U2276 (N_2276,N_2144,N_2167);
or U2277 (N_2277,N_2147,N_2150);
nand U2278 (N_2278,N_2181,N_2007);
nand U2279 (N_2279,N_2191,N_2136);
or U2280 (N_2280,N_2063,N_2066);
nand U2281 (N_2281,N_2039,N_2131);
and U2282 (N_2282,N_2059,N_2019);
or U2283 (N_2283,N_2183,N_2179);
nor U2284 (N_2284,N_2012,N_2041);
nand U2285 (N_2285,N_2177,N_2003);
or U2286 (N_2286,N_2070,N_2143);
nand U2287 (N_2287,N_2100,N_2138);
nor U2288 (N_2288,N_2040,N_2199);
xnor U2289 (N_2289,N_2155,N_2005);
and U2290 (N_2290,N_2172,N_2171);
nand U2291 (N_2291,N_2162,N_2068);
nand U2292 (N_2292,N_2160,N_2004);
nand U2293 (N_2293,N_2194,N_2197);
or U2294 (N_2294,N_2064,N_2053);
or U2295 (N_2295,N_2013,N_2051);
xnor U2296 (N_2296,N_2048,N_2016);
and U2297 (N_2297,N_2052,N_2107);
xnor U2298 (N_2298,N_2135,N_2115);
nand U2299 (N_2299,N_2080,N_2159);
or U2300 (N_2300,N_2020,N_2166);
and U2301 (N_2301,N_2040,N_2156);
and U2302 (N_2302,N_2098,N_2116);
and U2303 (N_2303,N_2076,N_2180);
nor U2304 (N_2304,N_2033,N_2192);
nor U2305 (N_2305,N_2039,N_2116);
nand U2306 (N_2306,N_2177,N_2048);
nor U2307 (N_2307,N_2010,N_2015);
or U2308 (N_2308,N_2120,N_2071);
xor U2309 (N_2309,N_2073,N_2178);
nor U2310 (N_2310,N_2021,N_2113);
nand U2311 (N_2311,N_2078,N_2079);
nand U2312 (N_2312,N_2025,N_2194);
or U2313 (N_2313,N_2002,N_2179);
or U2314 (N_2314,N_2095,N_2021);
or U2315 (N_2315,N_2048,N_2096);
nand U2316 (N_2316,N_2015,N_2119);
and U2317 (N_2317,N_2177,N_2106);
or U2318 (N_2318,N_2121,N_2153);
or U2319 (N_2319,N_2089,N_2031);
nand U2320 (N_2320,N_2165,N_2005);
or U2321 (N_2321,N_2006,N_2084);
xnor U2322 (N_2322,N_2022,N_2052);
nor U2323 (N_2323,N_2123,N_2064);
nor U2324 (N_2324,N_2067,N_2118);
nand U2325 (N_2325,N_2026,N_2174);
or U2326 (N_2326,N_2075,N_2089);
and U2327 (N_2327,N_2192,N_2094);
nor U2328 (N_2328,N_2002,N_2055);
and U2329 (N_2329,N_2003,N_2082);
and U2330 (N_2330,N_2068,N_2091);
or U2331 (N_2331,N_2171,N_2030);
nand U2332 (N_2332,N_2009,N_2133);
xor U2333 (N_2333,N_2013,N_2137);
and U2334 (N_2334,N_2056,N_2093);
xnor U2335 (N_2335,N_2133,N_2062);
or U2336 (N_2336,N_2101,N_2117);
or U2337 (N_2337,N_2094,N_2002);
and U2338 (N_2338,N_2069,N_2125);
or U2339 (N_2339,N_2081,N_2123);
and U2340 (N_2340,N_2020,N_2052);
and U2341 (N_2341,N_2186,N_2160);
or U2342 (N_2342,N_2030,N_2175);
nor U2343 (N_2343,N_2149,N_2195);
nand U2344 (N_2344,N_2033,N_2133);
xor U2345 (N_2345,N_2187,N_2148);
xnor U2346 (N_2346,N_2190,N_2107);
nand U2347 (N_2347,N_2173,N_2099);
or U2348 (N_2348,N_2017,N_2195);
or U2349 (N_2349,N_2106,N_2059);
or U2350 (N_2350,N_2123,N_2086);
and U2351 (N_2351,N_2080,N_2059);
nor U2352 (N_2352,N_2005,N_2087);
and U2353 (N_2353,N_2133,N_2088);
and U2354 (N_2354,N_2094,N_2147);
nor U2355 (N_2355,N_2059,N_2188);
nor U2356 (N_2356,N_2061,N_2058);
nor U2357 (N_2357,N_2150,N_2079);
or U2358 (N_2358,N_2054,N_2105);
nand U2359 (N_2359,N_2168,N_2185);
or U2360 (N_2360,N_2183,N_2194);
nand U2361 (N_2361,N_2102,N_2103);
nor U2362 (N_2362,N_2008,N_2131);
or U2363 (N_2363,N_2182,N_2066);
nand U2364 (N_2364,N_2113,N_2064);
nand U2365 (N_2365,N_2138,N_2145);
and U2366 (N_2366,N_2081,N_2005);
and U2367 (N_2367,N_2159,N_2158);
nor U2368 (N_2368,N_2071,N_2185);
or U2369 (N_2369,N_2197,N_2007);
nor U2370 (N_2370,N_2006,N_2031);
and U2371 (N_2371,N_2015,N_2120);
nand U2372 (N_2372,N_2175,N_2180);
nor U2373 (N_2373,N_2136,N_2066);
nand U2374 (N_2374,N_2001,N_2067);
and U2375 (N_2375,N_2048,N_2012);
or U2376 (N_2376,N_2182,N_2025);
nand U2377 (N_2377,N_2191,N_2107);
and U2378 (N_2378,N_2038,N_2118);
nand U2379 (N_2379,N_2085,N_2062);
nor U2380 (N_2380,N_2162,N_2017);
and U2381 (N_2381,N_2008,N_2145);
nand U2382 (N_2382,N_2080,N_2195);
nand U2383 (N_2383,N_2181,N_2197);
nand U2384 (N_2384,N_2116,N_2071);
nand U2385 (N_2385,N_2078,N_2177);
nand U2386 (N_2386,N_2007,N_2002);
nand U2387 (N_2387,N_2126,N_2161);
and U2388 (N_2388,N_2173,N_2189);
nor U2389 (N_2389,N_2192,N_2052);
and U2390 (N_2390,N_2117,N_2064);
or U2391 (N_2391,N_2095,N_2080);
and U2392 (N_2392,N_2016,N_2071);
nor U2393 (N_2393,N_2192,N_2007);
or U2394 (N_2394,N_2010,N_2065);
and U2395 (N_2395,N_2070,N_2026);
or U2396 (N_2396,N_2120,N_2173);
nand U2397 (N_2397,N_2035,N_2015);
and U2398 (N_2398,N_2130,N_2174);
and U2399 (N_2399,N_2073,N_2170);
nand U2400 (N_2400,N_2266,N_2250);
or U2401 (N_2401,N_2297,N_2257);
nor U2402 (N_2402,N_2332,N_2296);
nor U2403 (N_2403,N_2333,N_2331);
and U2404 (N_2404,N_2293,N_2281);
and U2405 (N_2405,N_2267,N_2279);
xnor U2406 (N_2406,N_2262,N_2208);
or U2407 (N_2407,N_2317,N_2213);
or U2408 (N_2408,N_2209,N_2248);
nor U2409 (N_2409,N_2367,N_2295);
xnor U2410 (N_2410,N_2339,N_2342);
xor U2411 (N_2411,N_2280,N_2382);
nand U2412 (N_2412,N_2299,N_2237);
and U2413 (N_2413,N_2277,N_2256);
and U2414 (N_2414,N_2230,N_2211);
and U2415 (N_2415,N_2320,N_2285);
nand U2416 (N_2416,N_2274,N_2329);
or U2417 (N_2417,N_2340,N_2228);
nand U2418 (N_2418,N_2217,N_2356);
or U2419 (N_2419,N_2222,N_2231);
and U2420 (N_2420,N_2380,N_2225);
and U2421 (N_2421,N_2328,N_2206);
or U2422 (N_2422,N_2304,N_2284);
or U2423 (N_2423,N_2303,N_2353);
nand U2424 (N_2424,N_2243,N_2319);
nand U2425 (N_2425,N_2330,N_2275);
and U2426 (N_2426,N_2210,N_2212);
nand U2427 (N_2427,N_2360,N_2252);
nor U2428 (N_2428,N_2325,N_2239);
nand U2429 (N_2429,N_2316,N_2207);
xor U2430 (N_2430,N_2387,N_2326);
nor U2431 (N_2431,N_2286,N_2246);
nor U2432 (N_2432,N_2273,N_2287);
nand U2433 (N_2433,N_2318,N_2364);
and U2434 (N_2434,N_2347,N_2323);
or U2435 (N_2435,N_2300,N_2288);
and U2436 (N_2436,N_2397,N_2346);
or U2437 (N_2437,N_2391,N_2254);
and U2438 (N_2438,N_2271,N_2334);
and U2439 (N_2439,N_2201,N_2311);
nor U2440 (N_2440,N_2388,N_2375);
or U2441 (N_2441,N_2392,N_2338);
and U2442 (N_2442,N_2224,N_2272);
or U2443 (N_2443,N_2242,N_2358);
and U2444 (N_2444,N_2363,N_2258);
or U2445 (N_2445,N_2255,N_2369);
xnor U2446 (N_2446,N_2355,N_2309);
nand U2447 (N_2447,N_2259,N_2386);
and U2448 (N_2448,N_2270,N_2384);
nor U2449 (N_2449,N_2261,N_2315);
nand U2450 (N_2450,N_2349,N_2322);
nor U2451 (N_2451,N_2200,N_2268);
nor U2452 (N_2452,N_2354,N_2241);
nand U2453 (N_2453,N_2378,N_2351);
xnor U2454 (N_2454,N_2381,N_2276);
nand U2455 (N_2455,N_2253,N_2232);
or U2456 (N_2456,N_2229,N_2389);
xor U2457 (N_2457,N_2306,N_2298);
xor U2458 (N_2458,N_2373,N_2362);
nand U2459 (N_2459,N_2219,N_2290);
and U2460 (N_2460,N_2289,N_2234);
nor U2461 (N_2461,N_2377,N_2366);
and U2462 (N_2462,N_2361,N_2383);
and U2463 (N_2463,N_2227,N_2305);
and U2464 (N_2464,N_2376,N_2269);
or U2465 (N_2465,N_2221,N_2370);
and U2466 (N_2466,N_2348,N_2240);
and U2467 (N_2467,N_2308,N_2283);
and U2468 (N_2468,N_2394,N_2327);
or U2469 (N_2469,N_2292,N_2226);
or U2470 (N_2470,N_2336,N_2359);
or U2471 (N_2471,N_2372,N_2282);
xor U2472 (N_2472,N_2236,N_2313);
or U2473 (N_2473,N_2278,N_2235);
nand U2474 (N_2474,N_2357,N_2310);
or U2475 (N_2475,N_2314,N_2345);
xnor U2476 (N_2476,N_2291,N_2205);
xor U2477 (N_2477,N_2220,N_2365);
nor U2478 (N_2478,N_2396,N_2245);
nand U2479 (N_2479,N_2264,N_2399);
nor U2480 (N_2480,N_2247,N_2218);
and U2481 (N_2481,N_2350,N_2335);
and U2482 (N_2482,N_2385,N_2249);
or U2483 (N_2483,N_2352,N_2265);
nor U2484 (N_2484,N_2301,N_2341);
and U2485 (N_2485,N_2368,N_2371);
or U2486 (N_2486,N_2343,N_2263);
and U2487 (N_2487,N_2214,N_2233);
and U2488 (N_2488,N_2393,N_2215);
nor U2489 (N_2489,N_2374,N_2216);
nand U2490 (N_2490,N_2260,N_2204);
nor U2491 (N_2491,N_2312,N_2294);
or U2492 (N_2492,N_2203,N_2307);
and U2493 (N_2493,N_2223,N_2202);
xor U2494 (N_2494,N_2344,N_2302);
and U2495 (N_2495,N_2251,N_2379);
or U2496 (N_2496,N_2238,N_2398);
nor U2497 (N_2497,N_2337,N_2390);
and U2498 (N_2498,N_2324,N_2321);
or U2499 (N_2499,N_2395,N_2244);
or U2500 (N_2500,N_2209,N_2233);
nor U2501 (N_2501,N_2300,N_2316);
xor U2502 (N_2502,N_2305,N_2353);
nor U2503 (N_2503,N_2357,N_2226);
and U2504 (N_2504,N_2234,N_2359);
and U2505 (N_2505,N_2384,N_2252);
or U2506 (N_2506,N_2303,N_2312);
and U2507 (N_2507,N_2243,N_2230);
xnor U2508 (N_2508,N_2224,N_2346);
or U2509 (N_2509,N_2221,N_2212);
xor U2510 (N_2510,N_2328,N_2205);
nand U2511 (N_2511,N_2229,N_2314);
xor U2512 (N_2512,N_2385,N_2332);
nor U2513 (N_2513,N_2219,N_2283);
nor U2514 (N_2514,N_2203,N_2303);
or U2515 (N_2515,N_2273,N_2266);
nor U2516 (N_2516,N_2299,N_2312);
or U2517 (N_2517,N_2395,N_2371);
xor U2518 (N_2518,N_2289,N_2363);
nor U2519 (N_2519,N_2377,N_2324);
xnor U2520 (N_2520,N_2295,N_2243);
nand U2521 (N_2521,N_2390,N_2292);
or U2522 (N_2522,N_2316,N_2387);
nor U2523 (N_2523,N_2297,N_2209);
and U2524 (N_2524,N_2392,N_2384);
and U2525 (N_2525,N_2242,N_2210);
and U2526 (N_2526,N_2273,N_2352);
nor U2527 (N_2527,N_2376,N_2201);
nand U2528 (N_2528,N_2252,N_2235);
or U2529 (N_2529,N_2352,N_2294);
or U2530 (N_2530,N_2361,N_2285);
or U2531 (N_2531,N_2286,N_2331);
nor U2532 (N_2532,N_2273,N_2394);
and U2533 (N_2533,N_2238,N_2227);
and U2534 (N_2534,N_2384,N_2309);
or U2535 (N_2535,N_2347,N_2215);
and U2536 (N_2536,N_2298,N_2302);
nor U2537 (N_2537,N_2367,N_2351);
or U2538 (N_2538,N_2229,N_2220);
nand U2539 (N_2539,N_2204,N_2295);
nor U2540 (N_2540,N_2306,N_2359);
or U2541 (N_2541,N_2387,N_2266);
nand U2542 (N_2542,N_2245,N_2287);
or U2543 (N_2543,N_2360,N_2328);
nor U2544 (N_2544,N_2354,N_2228);
or U2545 (N_2545,N_2344,N_2266);
and U2546 (N_2546,N_2226,N_2294);
xnor U2547 (N_2547,N_2373,N_2375);
nand U2548 (N_2548,N_2382,N_2391);
nand U2549 (N_2549,N_2224,N_2232);
and U2550 (N_2550,N_2296,N_2329);
and U2551 (N_2551,N_2245,N_2317);
and U2552 (N_2552,N_2375,N_2322);
nor U2553 (N_2553,N_2219,N_2368);
nor U2554 (N_2554,N_2349,N_2387);
xnor U2555 (N_2555,N_2249,N_2366);
nand U2556 (N_2556,N_2327,N_2211);
nand U2557 (N_2557,N_2264,N_2207);
nand U2558 (N_2558,N_2354,N_2244);
nor U2559 (N_2559,N_2263,N_2269);
nor U2560 (N_2560,N_2342,N_2334);
xor U2561 (N_2561,N_2345,N_2311);
nor U2562 (N_2562,N_2362,N_2291);
or U2563 (N_2563,N_2318,N_2377);
or U2564 (N_2564,N_2278,N_2307);
nor U2565 (N_2565,N_2228,N_2291);
xor U2566 (N_2566,N_2212,N_2308);
or U2567 (N_2567,N_2338,N_2305);
and U2568 (N_2568,N_2212,N_2311);
and U2569 (N_2569,N_2248,N_2308);
nand U2570 (N_2570,N_2256,N_2296);
or U2571 (N_2571,N_2329,N_2360);
and U2572 (N_2572,N_2231,N_2213);
or U2573 (N_2573,N_2242,N_2331);
nor U2574 (N_2574,N_2285,N_2343);
xor U2575 (N_2575,N_2344,N_2368);
and U2576 (N_2576,N_2304,N_2293);
and U2577 (N_2577,N_2382,N_2340);
xnor U2578 (N_2578,N_2345,N_2263);
or U2579 (N_2579,N_2239,N_2265);
and U2580 (N_2580,N_2341,N_2382);
nand U2581 (N_2581,N_2359,N_2322);
and U2582 (N_2582,N_2278,N_2214);
nand U2583 (N_2583,N_2372,N_2302);
nor U2584 (N_2584,N_2390,N_2247);
nor U2585 (N_2585,N_2258,N_2226);
nand U2586 (N_2586,N_2271,N_2329);
xnor U2587 (N_2587,N_2365,N_2212);
nand U2588 (N_2588,N_2281,N_2356);
nand U2589 (N_2589,N_2348,N_2230);
or U2590 (N_2590,N_2310,N_2359);
and U2591 (N_2591,N_2274,N_2238);
xor U2592 (N_2592,N_2246,N_2324);
nor U2593 (N_2593,N_2301,N_2256);
or U2594 (N_2594,N_2340,N_2270);
nor U2595 (N_2595,N_2370,N_2306);
and U2596 (N_2596,N_2367,N_2392);
nor U2597 (N_2597,N_2240,N_2243);
nand U2598 (N_2598,N_2205,N_2270);
or U2599 (N_2599,N_2369,N_2234);
nand U2600 (N_2600,N_2558,N_2514);
xnor U2601 (N_2601,N_2598,N_2527);
nand U2602 (N_2602,N_2465,N_2487);
and U2603 (N_2603,N_2435,N_2511);
and U2604 (N_2604,N_2588,N_2522);
or U2605 (N_2605,N_2587,N_2485);
and U2606 (N_2606,N_2592,N_2551);
or U2607 (N_2607,N_2515,N_2506);
or U2608 (N_2608,N_2599,N_2420);
and U2609 (N_2609,N_2484,N_2539);
or U2610 (N_2610,N_2561,N_2519);
xor U2611 (N_2611,N_2474,N_2579);
and U2612 (N_2612,N_2500,N_2569);
xor U2613 (N_2613,N_2548,N_2455);
nor U2614 (N_2614,N_2526,N_2491);
and U2615 (N_2615,N_2573,N_2497);
nand U2616 (N_2616,N_2477,N_2440);
or U2617 (N_2617,N_2401,N_2541);
and U2618 (N_2618,N_2415,N_2597);
nor U2619 (N_2619,N_2512,N_2595);
nand U2620 (N_2620,N_2517,N_2430);
nand U2621 (N_2621,N_2553,N_2467);
and U2622 (N_2622,N_2529,N_2534);
or U2623 (N_2623,N_2576,N_2594);
nor U2624 (N_2624,N_2505,N_2525);
nor U2625 (N_2625,N_2468,N_2499);
nor U2626 (N_2626,N_2549,N_2414);
and U2627 (N_2627,N_2501,N_2466);
nand U2628 (N_2628,N_2448,N_2483);
and U2629 (N_2629,N_2509,N_2585);
or U2630 (N_2630,N_2563,N_2432);
and U2631 (N_2631,N_2596,N_2584);
or U2632 (N_2632,N_2470,N_2535);
nand U2633 (N_2633,N_2403,N_2419);
or U2634 (N_2634,N_2575,N_2578);
nand U2635 (N_2635,N_2564,N_2580);
xnor U2636 (N_2636,N_2528,N_2533);
nand U2637 (N_2637,N_2425,N_2422);
and U2638 (N_2638,N_2591,N_2490);
or U2639 (N_2639,N_2445,N_2433);
or U2640 (N_2640,N_2482,N_2408);
and U2641 (N_2641,N_2498,N_2442);
nand U2642 (N_2642,N_2590,N_2418);
or U2643 (N_2643,N_2531,N_2547);
nand U2644 (N_2644,N_2568,N_2532);
nor U2645 (N_2645,N_2520,N_2550);
and U2646 (N_2646,N_2469,N_2554);
nor U2647 (N_2647,N_2446,N_2417);
or U2648 (N_2648,N_2503,N_2504);
and U2649 (N_2649,N_2404,N_2577);
nor U2650 (N_2650,N_2493,N_2513);
nand U2651 (N_2651,N_2582,N_2479);
nor U2652 (N_2652,N_2400,N_2431);
nand U2653 (N_2653,N_2492,N_2406);
nor U2654 (N_2654,N_2556,N_2447);
or U2655 (N_2655,N_2496,N_2586);
xor U2656 (N_2656,N_2544,N_2473);
or U2657 (N_2657,N_2495,N_2542);
or U2658 (N_2658,N_2540,N_2426);
and U2659 (N_2659,N_2502,N_2475);
or U2660 (N_2660,N_2508,N_2574);
or U2661 (N_2661,N_2530,N_2460);
nor U2662 (N_2662,N_2557,N_2565);
and U2663 (N_2663,N_2476,N_2507);
or U2664 (N_2664,N_2521,N_2518);
or U2665 (N_2665,N_2524,N_2489);
nand U2666 (N_2666,N_2413,N_2480);
nor U2667 (N_2667,N_2472,N_2444);
nand U2668 (N_2668,N_2428,N_2436);
nor U2669 (N_2669,N_2566,N_2571);
or U2670 (N_2670,N_2438,N_2562);
nand U2671 (N_2671,N_2464,N_2449);
and U2672 (N_2672,N_2461,N_2581);
or U2673 (N_2673,N_2516,N_2463);
nor U2674 (N_2674,N_2443,N_2452);
or U2675 (N_2675,N_2410,N_2416);
and U2676 (N_2676,N_2537,N_2421);
and U2677 (N_2677,N_2450,N_2481);
xor U2678 (N_2678,N_2546,N_2572);
and U2679 (N_2679,N_2462,N_2494);
and U2680 (N_2680,N_2429,N_2434);
and U2681 (N_2681,N_2589,N_2552);
nor U2682 (N_2682,N_2402,N_2543);
nand U2683 (N_2683,N_2453,N_2459);
nand U2684 (N_2684,N_2560,N_2471);
nand U2685 (N_2685,N_2458,N_2510);
nand U2686 (N_2686,N_2536,N_2457);
or U2687 (N_2687,N_2407,N_2570);
nor U2688 (N_2688,N_2454,N_2583);
or U2689 (N_2689,N_2456,N_2478);
or U2690 (N_2690,N_2545,N_2423);
nand U2691 (N_2691,N_2409,N_2555);
xnor U2692 (N_2692,N_2593,N_2412);
xor U2693 (N_2693,N_2424,N_2523);
or U2694 (N_2694,N_2441,N_2427);
nand U2695 (N_2695,N_2451,N_2405);
nor U2696 (N_2696,N_2567,N_2437);
nor U2697 (N_2697,N_2439,N_2559);
and U2698 (N_2698,N_2411,N_2486);
nor U2699 (N_2699,N_2538,N_2488);
nor U2700 (N_2700,N_2470,N_2486);
nand U2701 (N_2701,N_2518,N_2447);
nor U2702 (N_2702,N_2522,N_2568);
nand U2703 (N_2703,N_2566,N_2422);
and U2704 (N_2704,N_2585,N_2507);
xor U2705 (N_2705,N_2460,N_2579);
nand U2706 (N_2706,N_2567,N_2502);
or U2707 (N_2707,N_2571,N_2429);
xor U2708 (N_2708,N_2581,N_2574);
nand U2709 (N_2709,N_2557,N_2541);
or U2710 (N_2710,N_2535,N_2585);
nand U2711 (N_2711,N_2477,N_2566);
nor U2712 (N_2712,N_2474,N_2457);
and U2713 (N_2713,N_2476,N_2528);
or U2714 (N_2714,N_2551,N_2588);
or U2715 (N_2715,N_2553,N_2564);
or U2716 (N_2716,N_2579,N_2537);
nor U2717 (N_2717,N_2420,N_2598);
and U2718 (N_2718,N_2438,N_2452);
nand U2719 (N_2719,N_2478,N_2583);
or U2720 (N_2720,N_2407,N_2551);
nor U2721 (N_2721,N_2574,N_2457);
nor U2722 (N_2722,N_2413,N_2442);
xor U2723 (N_2723,N_2420,N_2500);
nand U2724 (N_2724,N_2443,N_2428);
nand U2725 (N_2725,N_2521,N_2487);
or U2726 (N_2726,N_2534,N_2527);
nand U2727 (N_2727,N_2569,N_2507);
or U2728 (N_2728,N_2504,N_2449);
xnor U2729 (N_2729,N_2569,N_2418);
nor U2730 (N_2730,N_2444,N_2572);
nand U2731 (N_2731,N_2430,N_2437);
or U2732 (N_2732,N_2412,N_2569);
xnor U2733 (N_2733,N_2510,N_2583);
or U2734 (N_2734,N_2454,N_2505);
and U2735 (N_2735,N_2541,N_2459);
xor U2736 (N_2736,N_2498,N_2552);
or U2737 (N_2737,N_2552,N_2508);
xor U2738 (N_2738,N_2583,N_2426);
nor U2739 (N_2739,N_2512,N_2590);
and U2740 (N_2740,N_2421,N_2538);
or U2741 (N_2741,N_2534,N_2593);
or U2742 (N_2742,N_2434,N_2422);
nor U2743 (N_2743,N_2405,N_2515);
nor U2744 (N_2744,N_2514,N_2498);
or U2745 (N_2745,N_2592,N_2571);
or U2746 (N_2746,N_2567,N_2538);
and U2747 (N_2747,N_2432,N_2480);
xor U2748 (N_2748,N_2484,N_2485);
and U2749 (N_2749,N_2570,N_2496);
nor U2750 (N_2750,N_2461,N_2584);
nand U2751 (N_2751,N_2546,N_2551);
xnor U2752 (N_2752,N_2584,N_2503);
xor U2753 (N_2753,N_2508,N_2408);
nor U2754 (N_2754,N_2546,N_2485);
nand U2755 (N_2755,N_2405,N_2445);
or U2756 (N_2756,N_2502,N_2554);
nor U2757 (N_2757,N_2504,N_2404);
and U2758 (N_2758,N_2594,N_2447);
and U2759 (N_2759,N_2479,N_2521);
and U2760 (N_2760,N_2545,N_2428);
and U2761 (N_2761,N_2457,N_2500);
and U2762 (N_2762,N_2471,N_2435);
and U2763 (N_2763,N_2497,N_2428);
or U2764 (N_2764,N_2490,N_2403);
nor U2765 (N_2765,N_2415,N_2503);
or U2766 (N_2766,N_2569,N_2553);
xor U2767 (N_2767,N_2594,N_2591);
and U2768 (N_2768,N_2459,N_2450);
or U2769 (N_2769,N_2454,N_2466);
and U2770 (N_2770,N_2568,N_2460);
nand U2771 (N_2771,N_2406,N_2532);
nand U2772 (N_2772,N_2473,N_2412);
and U2773 (N_2773,N_2450,N_2436);
nand U2774 (N_2774,N_2493,N_2550);
or U2775 (N_2775,N_2490,N_2527);
nor U2776 (N_2776,N_2591,N_2561);
or U2777 (N_2777,N_2582,N_2440);
nand U2778 (N_2778,N_2561,N_2481);
or U2779 (N_2779,N_2526,N_2420);
and U2780 (N_2780,N_2532,N_2492);
and U2781 (N_2781,N_2550,N_2480);
or U2782 (N_2782,N_2597,N_2402);
or U2783 (N_2783,N_2527,N_2465);
xnor U2784 (N_2784,N_2512,N_2526);
nor U2785 (N_2785,N_2441,N_2503);
xor U2786 (N_2786,N_2518,N_2568);
or U2787 (N_2787,N_2506,N_2413);
and U2788 (N_2788,N_2486,N_2537);
xor U2789 (N_2789,N_2401,N_2553);
and U2790 (N_2790,N_2442,N_2400);
nand U2791 (N_2791,N_2594,N_2518);
or U2792 (N_2792,N_2561,N_2535);
or U2793 (N_2793,N_2544,N_2434);
and U2794 (N_2794,N_2540,N_2490);
nand U2795 (N_2795,N_2553,N_2457);
and U2796 (N_2796,N_2524,N_2558);
or U2797 (N_2797,N_2546,N_2445);
nor U2798 (N_2798,N_2539,N_2435);
xor U2799 (N_2799,N_2596,N_2471);
and U2800 (N_2800,N_2778,N_2740);
nor U2801 (N_2801,N_2749,N_2707);
xnor U2802 (N_2802,N_2750,N_2670);
or U2803 (N_2803,N_2719,N_2773);
nand U2804 (N_2804,N_2678,N_2744);
nand U2805 (N_2805,N_2601,N_2632);
nor U2806 (N_2806,N_2709,N_2793);
nor U2807 (N_2807,N_2787,N_2761);
or U2808 (N_2808,N_2713,N_2722);
or U2809 (N_2809,N_2685,N_2792);
nand U2810 (N_2810,N_2731,N_2769);
nand U2811 (N_2811,N_2646,N_2635);
or U2812 (N_2812,N_2681,N_2779);
or U2813 (N_2813,N_2711,N_2768);
nand U2814 (N_2814,N_2715,N_2637);
nor U2815 (N_2815,N_2651,N_2694);
nor U2816 (N_2816,N_2746,N_2669);
nand U2817 (N_2817,N_2757,N_2683);
nor U2818 (N_2818,N_2727,N_2622);
nor U2819 (N_2819,N_2703,N_2643);
nand U2820 (N_2820,N_2755,N_2693);
nor U2821 (N_2821,N_2686,N_2777);
and U2822 (N_2822,N_2701,N_2605);
and U2823 (N_2823,N_2620,N_2742);
nor U2824 (N_2824,N_2760,N_2650);
nand U2825 (N_2825,N_2619,N_2795);
or U2826 (N_2826,N_2789,N_2763);
nand U2827 (N_2827,N_2663,N_2780);
or U2828 (N_2828,N_2790,N_2762);
nor U2829 (N_2829,N_2717,N_2676);
nor U2830 (N_2830,N_2700,N_2785);
and U2831 (N_2831,N_2626,N_2680);
and U2832 (N_2832,N_2614,N_2667);
or U2833 (N_2833,N_2736,N_2739);
nand U2834 (N_2834,N_2606,N_2775);
xnor U2835 (N_2835,N_2674,N_2774);
xor U2836 (N_2836,N_2788,N_2600);
and U2837 (N_2837,N_2690,N_2623);
and U2838 (N_2838,N_2672,N_2733);
and U2839 (N_2839,N_2689,N_2786);
nand U2840 (N_2840,N_2696,N_2721);
nand U2841 (N_2841,N_2756,N_2636);
nor U2842 (N_2842,N_2671,N_2603);
and U2843 (N_2843,N_2723,N_2714);
or U2844 (N_2844,N_2726,N_2611);
nor U2845 (N_2845,N_2615,N_2695);
nand U2846 (N_2846,N_2654,N_2638);
and U2847 (N_2847,N_2708,N_2698);
nor U2848 (N_2848,N_2630,N_2718);
nor U2849 (N_2849,N_2668,N_2642);
and U2850 (N_2850,N_2737,N_2675);
or U2851 (N_2851,N_2649,N_2662);
and U2852 (N_2852,N_2758,N_2791);
or U2853 (N_2853,N_2738,N_2627);
xnor U2854 (N_2854,N_2797,N_2647);
and U2855 (N_2855,N_2609,N_2652);
nor U2856 (N_2856,N_2765,N_2732);
nand U2857 (N_2857,N_2618,N_2759);
nor U2858 (N_2858,N_2604,N_2602);
nor U2859 (N_2859,N_2706,N_2613);
nand U2860 (N_2860,N_2608,N_2641);
or U2861 (N_2861,N_2659,N_2655);
or U2862 (N_2862,N_2702,N_2640);
or U2863 (N_2863,N_2741,N_2767);
nor U2864 (N_2864,N_2612,N_2782);
nor U2865 (N_2865,N_2661,N_2677);
or U2866 (N_2866,N_2682,N_2666);
nor U2867 (N_2867,N_2658,N_2625);
nor U2868 (N_2868,N_2783,N_2764);
or U2869 (N_2869,N_2631,N_2728);
and U2870 (N_2870,N_2617,N_2621);
or U2871 (N_2871,N_2716,N_2752);
nor U2872 (N_2872,N_2730,N_2624);
and U2873 (N_2873,N_2691,N_2634);
and U2874 (N_2874,N_2610,N_2616);
and U2875 (N_2875,N_2799,N_2705);
nand U2876 (N_2876,N_2697,N_2745);
nor U2877 (N_2877,N_2794,N_2771);
xor U2878 (N_2878,N_2665,N_2660);
xor U2879 (N_2879,N_2734,N_2781);
nor U2880 (N_2880,N_2729,N_2687);
nor U2881 (N_2881,N_2724,N_2710);
and U2882 (N_2882,N_2644,N_2754);
nand U2883 (N_2883,N_2657,N_2639);
or U2884 (N_2884,N_2679,N_2656);
or U2885 (N_2885,N_2673,N_2688);
and U2886 (N_2886,N_2692,N_2664);
nand U2887 (N_2887,N_2770,N_2648);
nor U2888 (N_2888,N_2776,N_2796);
and U2889 (N_2889,N_2753,N_2645);
or U2890 (N_2890,N_2747,N_2798);
nand U2891 (N_2891,N_2766,N_2607);
nor U2892 (N_2892,N_2725,N_2628);
nor U2893 (N_2893,N_2784,N_2712);
or U2894 (N_2894,N_2748,N_2704);
nand U2895 (N_2895,N_2699,N_2720);
or U2896 (N_2896,N_2772,N_2629);
nand U2897 (N_2897,N_2751,N_2684);
nor U2898 (N_2898,N_2743,N_2633);
nand U2899 (N_2899,N_2653,N_2735);
and U2900 (N_2900,N_2695,N_2771);
nand U2901 (N_2901,N_2782,N_2666);
nand U2902 (N_2902,N_2644,N_2640);
nor U2903 (N_2903,N_2697,N_2641);
or U2904 (N_2904,N_2682,N_2737);
nor U2905 (N_2905,N_2628,N_2621);
or U2906 (N_2906,N_2759,N_2704);
and U2907 (N_2907,N_2608,N_2633);
nand U2908 (N_2908,N_2717,N_2767);
xnor U2909 (N_2909,N_2633,N_2787);
xnor U2910 (N_2910,N_2794,N_2746);
xor U2911 (N_2911,N_2612,N_2794);
nand U2912 (N_2912,N_2630,N_2710);
nor U2913 (N_2913,N_2734,N_2648);
or U2914 (N_2914,N_2724,N_2696);
xor U2915 (N_2915,N_2612,N_2755);
nor U2916 (N_2916,N_2638,N_2775);
nand U2917 (N_2917,N_2693,N_2671);
nor U2918 (N_2918,N_2763,N_2798);
nor U2919 (N_2919,N_2714,N_2776);
nand U2920 (N_2920,N_2621,N_2743);
and U2921 (N_2921,N_2605,N_2774);
nor U2922 (N_2922,N_2691,N_2639);
nand U2923 (N_2923,N_2719,N_2758);
nor U2924 (N_2924,N_2628,N_2770);
nand U2925 (N_2925,N_2692,N_2716);
nor U2926 (N_2926,N_2726,N_2720);
and U2927 (N_2927,N_2698,N_2694);
nand U2928 (N_2928,N_2739,N_2701);
or U2929 (N_2929,N_2789,N_2708);
nor U2930 (N_2930,N_2784,N_2731);
nor U2931 (N_2931,N_2712,N_2659);
or U2932 (N_2932,N_2703,N_2686);
or U2933 (N_2933,N_2602,N_2638);
or U2934 (N_2934,N_2605,N_2699);
and U2935 (N_2935,N_2687,N_2737);
and U2936 (N_2936,N_2721,N_2708);
and U2937 (N_2937,N_2619,N_2693);
xor U2938 (N_2938,N_2660,N_2629);
and U2939 (N_2939,N_2780,N_2654);
nor U2940 (N_2940,N_2696,N_2781);
nor U2941 (N_2941,N_2759,N_2751);
nand U2942 (N_2942,N_2662,N_2624);
and U2943 (N_2943,N_2645,N_2791);
nor U2944 (N_2944,N_2628,N_2699);
and U2945 (N_2945,N_2717,N_2659);
nand U2946 (N_2946,N_2707,N_2741);
nand U2947 (N_2947,N_2693,N_2605);
xor U2948 (N_2948,N_2625,N_2797);
and U2949 (N_2949,N_2642,N_2766);
nor U2950 (N_2950,N_2719,N_2674);
nand U2951 (N_2951,N_2694,N_2667);
nor U2952 (N_2952,N_2733,N_2641);
nand U2953 (N_2953,N_2773,N_2699);
nand U2954 (N_2954,N_2658,N_2730);
nand U2955 (N_2955,N_2778,N_2795);
nand U2956 (N_2956,N_2775,N_2615);
or U2957 (N_2957,N_2704,N_2783);
xor U2958 (N_2958,N_2642,N_2719);
nand U2959 (N_2959,N_2706,N_2668);
nor U2960 (N_2960,N_2761,N_2615);
nand U2961 (N_2961,N_2741,N_2761);
or U2962 (N_2962,N_2711,N_2722);
nand U2963 (N_2963,N_2718,N_2763);
and U2964 (N_2964,N_2678,N_2604);
nor U2965 (N_2965,N_2789,N_2727);
and U2966 (N_2966,N_2707,N_2766);
and U2967 (N_2967,N_2694,N_2799);
nor U2968 (N_2968,N_2787,N_2788);
nor U2969 (N_2969,N_2777,N_2737);
nand U2970 (N_2970,N_2634,N_2614);
nor U2971 (N_2971,N_2660,N_2713);
and U2972 (N_2972,N_2787,N_2707);
nand U2973 (N_2973,N_2701,N_2646);
and U2974 (N_2974,N_2695,N_2693);
nand U2975 (N_2975,N_2785,N_2798);
or U2976 (N_2976,N_2650,N_2708);
nand U2977 (N_2977,N_2762,N_2722);
nor U2978 (N_2978,N_2616,N_2748);
nor U2979 (N_2979,N_2722,N_2790);
nand U2980 (N_2980,N_2645,N_2682);
and U2981 (N_2981,N_2615,N_2755);
nor U2982 (N_2982,N_2721,N_2774);
nand U2983 (N_2983,N_2669,N_2705);
nor U2984 (N_2984,N_2706,N_2705);
nor U2985 (N_2985,N_2620,N_2780);
nand U2986 (N_2986,N_2616,N_2604);
and U2987 (N_2987,N_2603,N_2798);
and U2988 (N_2988,N_2651,N_2681);
and U2989 (N_2989,N_2703,N_2603);
xor U2990 (N_2990,N_2792,N_2736);
and U2991 (N_2991,N_2793,N_2649);
nor U2992 (N_2992,N_2636,N_2616);
nand U2993 (N_2993,N_2744,N_2773);
nand U2994 (N_2994,N_2606,N_2760);
and U2995 (N_2995,N_2755,N_2670);
and U2996 (N_2996,N_2683,N_2695);
nor U2997 (N_2997,N_2687,N_2663);
or U2998 (N_2998,N_2625,N_2605);
or U2999 (N_2999,N_2789,N_2798);
or UO_0 (O_0,N_2951,N_2840);
nand UO_1 (O_1,N_2895,N_2893);
and UO_2 (O_2,N_2938,N_2833);
and UO_3 (O_3,N_2890,N_2891);
nand UO_4 (O_4,N_2942,N_2912);
or UO_5 (O_5,N_2920,N_2985);
nor UO_6 (O_6,N_2968,N_2998);
or UO_7 (O_7,N_2952,N_2929);
xnor UO_8 (O_8,N_2806,N_2991);
nor UO_9 (O_9,N_2953,N_2835);
or UO_10 (O_10,N_2902,N_2870);
nor UO_11 (O_11,N_2863,N_2831);
xor UO_12 (O_12,N_2880,N_2856);
nor UO_13 (O_13,N_2901,N_2868);
nor UO_14 (O_14,N_2958,N_2857);
nand UO_15 (O_15,N_2919,N_2913);
nand UO_16 (O_16,N_2839,N_2947);
xor UO_17 (O_17,N_2800,N_2842);
or UO_18 (O_18,N_2892,N_2841);
nor UO_19 (O_19,N_2972,N_2862);
nand UO_20 (O_20,N_2937,N_2943);
xor UO_21 (O_21,N_2871,N_2969);
nor UO_22 (O_22,N_2860,N_2996);
and UO_23 (O_23,N_2861,N_2818);
and UO_24 (O_24,N_2960,N_2925);
or UO_25 (O_25,N_2975,N_2944);
nand UO_26 (O_26,N_2829,N_2982);
xor UO_27 (O_27,N_2804,N_2986);
and UO_28 (O_28,N_2808,N_2810);
or UO_29 (O_29,N_2971,N_2956);
nand UO_30 (O_30,N_2801,N_2889);
nand UO_31 (O_31,N_2894,N_2917);
and UO_32 (O_32,N_2990,N_2916);
and UO_33 (O_33,N_2898,N_2957);
or UO_34 (O_34,N_2995,N_2845);
and UO_35 (O_35,N_2961,N_2907);
nand UO_36 (O_36,N_2979,N_2915);
and UO_37 (O_37,N_2906,N_2928);
nand UO_38 (O_38,N_2877,N_2876);
nor UO_39 (O_39,N_2843,N_2875);
and UO_40 (O_40,N_2934,N_2932);
and UO_41 (O_41,N_2993,N_2981);
and UO_42 (O_42,N_2984,N_2978);
nor UO_43 (O_43,N_2935,N_2983);
nor UO_44 (O_44,N_2814,N_2992);
nor UO_45 (O_45,N_2989,N_2970);
nor UO_46 (O_46,N_2930,N_2827);
xnor UO_47 (O_47,N_2834,N_2824);
and UO_48 (O_48,N_2900,N_2885);
or UO_49 (O_49,N_2830,N_2909);
and UO_50 (O_50,N_2816,N_2918);
xnor UO_51 (O_51,N_2936,N_2964);
and UO_52 (O_52,N_2948,N_2836);
xnor UO_53 (O_53,N_2850,N_2977);
xnor UO_54 (O_54,N_2897,N_2844);
nor UO_55 (O_55,N_2987,N_2976);
and UO_56 (O_56,N_2881,N_2832);
nor UO_57 (O_57,N_2858,N_2838);
and UO_58 (O_58,N_2869,N_2949);
and UO_59 (O_59,N_2966,N_2846);
or UO_60 (O_60,N_2945,N_2904);
xor UO_61 (O_61,N_2851,N_2809);
or UO_62 (O_62,N_2883,N_2820);
or UO_63 (O_63,N_2821,N_2813);
nand UO_64 (O_64,N_2973,N_2896);
nor UO_65 (O_65,N_2914,N_2852);
nor UO_66 (O_66,N_2803,N_2874);
nand UO_67 (O_67,N_2940,N_2997);
nand UO_68 (O_68,N_2980,N_2848);
nand UO_69 (O_69,N_2923,N_2926);
and UO_70 (O_70,N_2908,N_2805);
nor UO_71 (O_71,N_2886,N_2866);
and UO_72 (O_72,N_2922,N_2941);
nand UO_73 (O_73,N_2823,N_2802);
nand UO_74 (O_74,N_2879,N_2965);
nor UO_75 (O_75,N_2988,N_2819);
nor UO_76 (O_76,N_2884,N_2903);
nand UO_77 (O_77,N_2867,N_2967);
nor UO_78 (O_78,N_2878,N_2954);
nand UO_79 (O_79,N_2905,N_2837);
nand UO_80 (O_80,N_2853,N_2849);
or UO_81 (O_81,N_2873,N_2847);
nor UO_82 (O_82,N_2815,N_2826);
or UO_83 (O_83,N_2865,N_2933);
xnor UO_84 (O_84,N_2811,N_2812);
xor UO_85 (O_85,N_2822,N_2921);
nor UO_86 (O_86,N_2974,N_2817);
and UO_87 (O_87,N_2994,N_2955);
nor UO_88 (O_88,N_2887,N_2859);
and UO_89 (O_89,N_2959,N_2950);
nand UO_90 (O_90,N_2946,N_2963);
nand UO_91 (O_91,N_2854,N_2899);
and UO_92 (O_92,N_2825,N_2872);
and UO_93 (O_93,N_2882,N_2911);
or UO_94 (O_94,N_2864,N_2910);
or UO_95 (O_95,N_2888,N_2962);
or UO_96 (O_96,N_2927,N_2855);
and UO_97 (O_97,N_2939,N_2924);
xor UO_98 (O_98,N_2807,N_2828);
and UO_99 (O_99,N_2999,N_2931);
and UO_100 (O_100,N_2943,N_2988);
nor UO_101 (O_101,N_2952,N_2998);
or UO_102 (O_102,N_2861,N_2921);
and UO_103 (O_103,N_2909,N_2953);
nand UO_104 (O_104,N_2923,N_2874);
and UO_105 (O_105,N_2861,N_2940);
nor UO_106 (O_106,N_2907,N_2808);
nor UO_107 (O_107,N_2812,N_2966);
nor UO_108 (O_108,N_2902,N_2953);
and UO_109 (O_109,N_2863,N_2830);
and UO_110 (O_110,N_2947,N_2836);
nor UO_111 (O_111,N_2901,N_2878);
nand UO_112 (O_112,N_2929,N_2984);
xor UO_113 (O_113,N_2882,N_2944);
nor UO_114 (O_114,N_2894,N_2819);
and UO_115 (O_115,N_2813,N_2963);
xnor UO_116 (O_116,N_2854,N_2978);
nor UO_117 (O_117,N_2976,N_2878);
nand UO_118 (O_118,N_2941,N_2824);
or UO_119 (O_119,N_2894,N_2951);
nand UO_120 (O_120,N_2949,N_2806);
nand UO_121 (O_121,N_2944,N_2886);
and UO_122 (O_122,N_2887,N_2845);
and UO_123 (O_123,N_2867,N_2859);
nand UO_124 (O_124,N_2887,N_2901);
xnor UO_125 (O_125,N_2938,N_2937);
xnor UO_126 (O_126,N_2880,N_2867);
nor UO_127 (O_127,N_2870,N_2865);
or UO_128 (O_128,N_2899,N_2904);
nor UO_129 (O_129,N_2994,N_2855);
nor UO_130 (O_130,N_2978,N_2803);
and UO_131 (O_131,N_2814,N_2839);
or UO_132 (O_132,N_2933,N_2859);
and UO_133 (O_133,N_2800,N_2894);
and UO_134 (O_134,N_2948,N_2972);
xnor UO_135 (O_135,N_2893,N_2999);
nor UO_136 (O_136,N_2948,N_2848);
and UO_137 (O_137,N_2838,N_2820);
nor UO_138 (O_138,N_2993,N_2937);
and UO_139 (O_139,N_2911,N_2893);
or UO_140 (O_140,N_2947,N_2887);
nor UO_141 (O_141,N_2896,N_2967);
or UO_142 (O_142,N_2931,N_2843);
xor UO_143 (O_143,N_2843,N_2917);
and UO_144 (O_144,N_2909,N_2917);
nor UO_145 (O_145,N_2926,N_2911);
or UO_146 (O_146,N_2840,N_2890);
nor UO_147 (O_147,N_2926,N_2933);
and UO_148 (O_148,N_2936,N_2989);
nand UO_149 (O_149,N_2992,N_2833);
or UO_150 (O_150,N_2923,N_2870);
or UO_151 (O_151,N_2886,N_2869);
nor UO_152 (O_152,N_2814,N_2940);
or UO_153 (O_153,N_2858,N_2878);
nor UO_154 (O_154,N_2817,N_2865);
xor UO_155 (O_155,N_2817,N_2824);
xor UO_156 (O_156,N_2970,N_2927);
nor UO_157 (O_157,N_2925,N_2814);
or UO_158 (O_158,N_2801,N_2999);
and UO_159 (O_159,N_2802,N_2926);
or UO_160 (O_160,N_2906,N_2870);
nand UO_161 (O_161,N_2957,N_2823);
nand UO_162 (O_162,N_2837,N_2855);
nand UO_163 (O_163,N_2827,N_2841);
xnor UO_164 (O_164,N_2920,N_2826);
nand UO_165 (O_165,N_2946,N_2977);
or UO_166 (O_166,N_2995,N_2953);
or UO_167 (O_167,N_2828,N_2929);
nand UO_168 (O_168,N_2926,N_2804);
nand UO_169 (O_169,N_2965,N_2960);
nand UO_170 (O_170,N_2946,N_2806);
nor UO_171 (O_171,N_2972,N_2925);
and UO_172 (O_172,N_2841,N_2834);
or UO_173 (O_173,N_2991,N_2974);
nand UO_174 (O_174,N_2941,N_2994);
or UO_175 (O_175,N_2906,N_2848);
nand UO_176 (O_176,N_2932,N_2836);
nor UO_177 (O_177,N_2906,N_2879);
and UO_178 (O_178,N_2969,N_2904);
or UO_179 (O_179,N_2987,N_2805);
and UO_180 (O_180,N_2859,N_2855);
nand UO_181 (O_181,N_2821,N_2872);
nand UO_182 (O_182,N_2881,N_2987);
nand UO_183 (O_183,N_2825,N_2805);
nand UO_184 (O_184,N_2855,N_2810);
nor UO_185 (O_185,N_2973,N_2936);
nand UO_186 (O_186,N_2869,N_2836);
nor UO_187 (O_187,N_2812,N_2976);
and UO_188 (O_188,N_2940,N_2830);
nor UO_189 (O_189,N_2844,N_2997);
xor UO_190 (O_190,N_2854,N_2996);
xor UO_191 (O_191,N_2968,N_2960);
nor UO_192 (O_192,N_2956,N_2917);
nand UO_193 (O_193,N_2852,N_2814);
or UO_194 (O_194,N_2971,N_2917);
or UO_195 (O_195,N_2809,N_2998);
nand UO_196 (O_196,N_2973,N_2947);
xor UO_197 (O_197,N_2893,N_2931);
nor UO_198 (O_198,N_2869,N_2996);
nand UO_199 (O_199,N_2893,N_2849);
nand UO_200 (O_200,N_2939,N_2942);
xor UO_201 (O_201,N_2859,N_2846);
nand UO_202 (O_202,N_2936,N_2985);
or UO_203 (O_203,N_2933,N_2942);
or UO_204 (O_204,N_2867,N_2968);
nor UO_205 (O_205,N_2802,N_2909);
or UO_206 (O_206,N_2894,N_2905);
nand UO_207 (O_207,N_2964,N_2900);
nor UO_208 (O_208,N_2887,N_2815);
nor UO_209 (O_209,N_2914,N_2900);
nor UO_210 (O_210,N_2984,N_2975);
or UO_211 (O_211,N_2985,N_2821);
nand UO_212 (O_212,N_2872,N_2987);
nand UO_213 (O_213,N_2928,N_2831);
nor UO_214 (O_214,N_2806,N_2802);
nor UO_215 (O_215,N_2916,N_2909);
or UO_216 (O_216,N_2896,N_2940);
nand UO_217 (O_217,N_2979,N_2929);
nor UO_218 (O_218,N_2988,N_2958);
nor UO_219 (O_219,N_2993,N_2967);
xor UO_220 (O_220,N_2954,N_2949);
nand UO_221 (O_221,N_2911,N_2908);
nand UO_222 (O_222,N_2923,N_2967);
nor UO_223 (O_223,N_2924,N_2952);
or UO_224 (O_224,N_2930,N_2830);
or UO_225 (O_225,N_2982,N_2881);
nor UO_226 (O_226,N_2922,N_2993);
or UO_227 (O_227,N_2980,N_2925);
and UO_228 (O_228,N_2978,N_2844);
xnor UO_229 (O_229,N_2864,N_2952);
nor UO_230 (O_230,N_2800,N_2990);
or UO_231 (O_231,N_2899,N_2834);
nand UO_232 (O_232,N_2956,N_2810);
and UO_233 (O_233,N_2940,N_2905);
xor UO_234 (O_234,N_2809,N_2847);
or UO_235 (O_235,N_2935,N_2939);
nand UO_236 (O_236,N_2861,N_2851);
nor UO_237 (O_237,N_2832,N_2979);
and UO_238 (O_238,N_2904,N_2807);
nand UO_239 (O_239,N_2989,N_2881);
nor UO_240 (O_240,N_2816,N_2805);
nor UO_241 (O_241,N_2846,N_2942);
nand UO_242 (O_242,N_2869,N_2874);
and UO_243 (O_243,N_2883,N_2804);
or UO_244 (O_244,N_2981,N_2985);
and UO_245 (O_245,N_2922,N_2810);
and UO_246 (O_246,N_2810,N_2952);
and UO_247 (O_247,N_2842,N_2969);
nor UO_248 (O_248,N_2821,N_2808);
or UO_249 (O_249,N_2968,N_2804);
xor UO_250 (O_250,N_2868,N_2804);
and UO_251 (O_251,N_2854,N_2914);
and UO_252 (O_252,N_2843,N_2974);
nand UO_253 (O_253,N_2854,N_2930);
or UO_254 (O_254,N_2900,N_2832);
nand UO_255 (O_255,N_2939,N_2836);
and UO_256 (O_256,N_2985,N_2970);
xnor UO_257 (O_257,N_2822,N_2974);
nand UO_258 (O_258,N_2874,N_2850);
and UO_259 (O_259,N_2955,N_2854);
nor UO_260 (O_260,N_2825,N_2804);
nor UO_261 (O_261,N_2867,N_2987);
or UO_262 (O_262,N_2945,N_2975);
xor UO_263 (O_263,N_2987,N_2856);
or UO_264 (O_264,N_2954,N_2895);
and UO_265 (O_265,N_2918,N_2919);
or UO_266 (O_266,N_2990,N_2804);
nand UO_267 (O_267,N_2812,N_2920);
and UO_268 (O_268,N_2960,N_2985);
and UO_269 (O_269,N_2832,N_2813);
and UO_270 (O_270,N_2916,N_2845);
nor UO_271 (O_271,N_2897,N_2948);
nor UO_272 (O_272,N_2992,N_2924);
nand UO_273 (O_273,N_2813,N_2924);
and UO_274 (O_274,N_2979,N_2822);
and UO_275 (O_275,N_2873,N_2982);
or UO_276 (O_276,N_2906,N_2827);
xor UO_277 (O_277,N_2826,N_2860);
nor UO_278 (O_278,N_2837,N_2848);
or UO_279 (O_279,N_2892,N_2836);
and UO_280 (O_280,N_2978,N_2836);
or UO_281 (O_281,N_2859,N_2811);
or UO_282 (O_282,N_2855,N_2928);
and UO_283 (O_283,N_2860,N_2830);
nand UO_284 (O_284,N_2929,N_2871);
nor UO_285 (O_285,N_2931,N_2904);
nor UO_286 (O_286,N_2964,N_2996);
and UO_287 (O_287,N_2826,N_2862);
nand UO_288 (O_288,N_2872,N_2897);
nand UO_289 (O_289,N_2979,N_2909);
nand UO_290 (O_290,N_2949,N_2941);
and UO_291 (O_291,N_2994,N_2854);
and UO_292 (O_292,N_2880,N_2943);
or UO_293 (O_293,N_2995,N_2888);
nor UO_294 (O_294,N_2826,N_2803);
xnor UO_295 (O_295,N_2931,N_2985);
or UO_296 (O_296,N_2829,N_2957);
nand UO_297 (O_297,N_2965,N_2976);
xor UO_298 (O_298,N_2894,N_2982);
or UO_299 (O_299,N_2877,N_2860);
and UO_300 (O_300,N_2865,N_2876);
or UO_301 (O_301,N_2905,N_2959);
nor UO_302 (O_302,N_2826,N_2882);
nand UO_303 (O_303,N_2807,N_2930);
or UO_304 (O_304,N_2839,N_2831);
nand UO_305 (O_305,N_2878,N_2947);
or UO_306 (O_306,N_2895,N_2925);
nand UO_307 (O_307,N_2999,N_2979);
and UO_308 (O_308,N_2869,N_2955);
nor UO_309 (O_309,N_2920,N_2981);
or UO_310 (O_310,N_2850,N_2903);
or UO_311 (O_311,N_2965,N_2966);
nand UO_312 (O_312,N_2902,N_2905);
or UO_313 (O_313,N_2851,N_2979);
xor UO_314 (O_314,N_2937,N_2957);
or UO_315 (O_315,N_2952,N_2838);
or UO_316 (O_316,N_2827,N_2936);
and UO_317 (O_317,N_2950,N_2818);
or UO_318 (O_318,N_2855,N_2937);
and UO_319 (O_319,N_2871,N_2827);
or UO_320 (O_320,N_2937,N_2814);
xor UO_321 (O_321,N_2827,N_2993);
or UO_322 (O_322,N_2804,N_2888);
nand UO_323 (O_323,N_2964,N_2882);
or UO_324 (O_324,N_2998,N_2916);
nand UO_325 (O_325,N_2896,N_2815);
and UO_326 (O_326,N_2820,N_2949);
and UO_327 (O_327,N_2876,N_2850);
xnor UO_328 (O_328,N_2939,N_2902);
xor UO_329 (O_329,N_2865,N_2851);
or UO_330 (O_330,N_2829,N_2921);
or UO_331 (O_331,N_2806,N_2824);
nor UO_332 (O_332,N_2888,N_2822);
nor UO_333 (O_333,N_2860,N_2939);
or UO_334 (O_334,N_2832,N_2840);
nand UO_335 (O_335,N_2832,N_2982);
xor UO_336 (O_336,N_2906,N_2887);
nor UO_337 (O_337,N_2946,N_2918);
nand UO_338 (O_338,N_2889,N_2985);
or UO_339 (O_339,N_2894,N_2962);
xnor UO_340 (O_340,N_2806,N_2940);
nor UO_341 (O_341,N_2804,N_2865);
xor UO_342 (O_342,N_2903,N_2811);
and UO_343 (O_343,N_2940,N_2875);
xor UO_344 (O_344,N_2931,N_2965);
nor UO_345 (O_345,N_2960,N_2939);
nor UO_346 (O_346,N_2966,N_2862);
and UO_347 (O_347,N_2870,N_2910);
nand UO_348 (O_348,N_2993,N_2992);
nor UO_349 (O_349,N_2976,N_2910);
nor UO_350 (O_350,N_2961,N_2804);
or UO_351 (O_351,N_2988,N_2956);
nand UO_352 (O_352,N_2870,N_2835);
and UO_353 (O_353,N_2806,N_2968);
and UO_354 (O_354,N_2919,N_2845);
nand UO_355 (O_355,N_2931,N_2942);
and UO_356 (O_356,N_2864,N_2849);
xor UO_357 (O_357,N_2860,N_2987);
and UO_358 (O_358,N_2898,N_2966);
nand UO_359 (O_359,N_2841,N_2871);
or UO_360 (O_360,N_2908,N_2937);
and UO_361 (O_361,N_2805,N_2887);
and UO_362 (O_362,N_2829,N_2885);
nor UO_363 (O_363,N_2877,N_2935);
nor UO_364 (O_364,N_2864,N_2891);
nor UO_365 (O_365,N_2915,N_2923);
or UO_366 (O_366,N_2841,N_2850);
nor UO_367 (O_367,N_2854,N_2935);
xnor UO_368 (O_368,N_2981,N_2958);
nand UO_369 (O_369,N_2873,N_2892);
nand UO_370 (O_370,N_2816,N_2929);
nand UO_371 (O_371,N_2882,N_2920);
or UO_372 (O_372,N_2802,N_2889);
nor UO_373 (O_373,N_2830,N_2974);
and UO_374 (O_374,N_2881,N_2844);
and UO_375 (O_375,N_2992,N_2841);
nand UO_376 (O_376,N_2869,N_2915);
and UO_377 (O_377,N_2872,N_2847);
and UO_378 (O_378,N_2983,N_2802);
and UO_379 (O_379,N_2848,N_2963);
or UO_380 (O_380,N_2840,N_2847);
or UO_381 (O_381,N_2909,N_2901);
and UO_382 (O_382,N_2804,N_2987);
or UO_383 (O_383,N_2801,N_2882);
nand UO_384 (O_384,N_2948,N_2850);
nand UO_385 (O_385,N_2965,N_2888);
xnor UO_386 (O_386,N_2915,N_2902);
nor UO_387 (O_387,N_2958,N_2869);
or UO_388 (O_388,N_2923,N_2827);
or UO_389 (O_389,N_2851,N_2973);
xor UO_390 (O_390,N_2880,N_2865);
nand UO_391 (O_391,N_2869,N_2973);
and UO_392 (O_392,N_2978,N_2950);
or UO_393 (O_393,N_2800,N_2970);
nand UO_394 (O_394,N_2844,N_2884);
nor UO_395 (O_395,N_2918,N_2801);
and UO_396 (O_396,N_2880,N_2809);
and UO_397 (O_397,N_2851,N_2985);
nand UO_398 (O_398,N_2878,N_2840);
xnor UO_399 (O_399,N_2864,N_2846);
and UO_400 (O_400,N_2938,N_2874);
xor UO_401 (O_401,N_2943,N_2938);
and UO_402 (O_402,N_2896,N_2894);
nor UO_403 (O_403,N_2894,N_2809);
nor UO_404 (O_404,N_2896,N_2824);
and UO_405 (O_405,N_2841,N_2895);
nor UO_406 (O_406,N_2975,N_2946);
xnor UO_407 (O_407,N_2997,N_2906);
or UO_408 (O_408,N_2947,N_2864);
and UO_409 (O_409,N_2917,N_2847);
nand UO_410 (O_410,N_2964,N_2930);
xor UO_411 (O_411,N_2918,N_2910);
or UO_412 (O_412,N_2941,N_2960);
xor UO_413 (O_413,N_2817,N_2969);
nand UO_414 (O_414,N_2834,N_2959);
nor UO_415 (O_415,N_2825,N_2818);
xnor UO_416 (O_416,N_2888,N_2917);
and UO_417 (O_417,N_2876,N_2838);
or UO_418 (O_418,N_2888,N_2900);
nand UO_419 (O_419,N_2969,N_2959);
nand UO_420 (O_420,N_2801,N_2807);
nor UO_421 (O_421,N_2954,N_2976);
nor UO_422 (O_422,N_2873,N_2929);
nor UO_423 (O_423,N_2930,N_2944);
or UO_424 (O_424,N_2903,N_2820);
and UO_425 (O_425,N_2820,N_2826);
and UO_426 (O_426,N_2952,N_2858);
or UO_427 (O_427,N_2995,N_2923);
and UO_428 (O_428,N_2976,N_2964);
or UO_429 (O_429,N_2816,N_2847);
or UO_430 (O_430,N_2982,N_2904);
nand UO_431 (O_431,N_2985,N_2957);
or UO_432 (O_432,N_2811,N_2814);
and UO_433 (O_433,N_2853,N_2858);
nor UO_434 (O_434,N_2909,N_2817);
nand UO_435 (O_435,N_2834,N_2941);
and UO_436 (O_436,N_2982,N_2902);
and UO_437 (O_437,N_2922,N_2908);
xnor UO_438 (O_438,N_2979,N_2823);
or UO_439 (O_439,N_2968,N_2847);
or UO_440 (O_440,N_2887,N_2953);
or UO_441 (O_441,N_2924,N_2998);
nand UO_442 (O_442,N_2884,N_2955);
nor UO_443 (O_443,N_2946,N_2807);
nand UO_444 (O_444,N_2885,N_2856);
nor UO_445 (O_445,N_2969,N_2818);
xor UO_446 (O_446,N_2920,N_2992);
and UO_447 (O_447,N_2841,N_2975);
nor UO_448 (O_448,N_2952,N_2880);
nand UO_449 (O_449,N_2904,N_2939);
nand UO_450 (O_450,N_2811,N_2834);
or UO_451 (O_451,N_2942,N_2967);
nand UO_452 (O_452,N_2998,N_2872);
or UO_453 (O_453,N_2879,N_2869);
nor UO_454 (O_454,N_2817,N_2843);
nand UO_455 (O_455,N_2859,N_2988);
xnor UO_456 (O_456,N_2811,N_2887);
nand UO_457 (O_457,N_2949,N_2853);
nor UO_458 (O_458,N_2867,N_2981);
or UO_459 (O_459,N_2915,N_2969);
xor UO_460 (O_460,N_2978,N_2829);
nor UO_461 (O_461,N_2810,N_2837);
and UO_462 (O_462,N_2927,N_2851);
xnor UO_463 (O_463,N_2971,N_2823);
or UO_464 (O_464,N_2886,N_2844);
or UO_465 (O_465,N_2816,N_2852);
nor UO_466 (O_466,N_2832,N_2963);
nand UO_467 (O_467,N_2800,N_2992);
and UO_468 (O_468,N_2971,N_2891);
nand UO_469 (O_469,N_2993,N_2831);
or UO_470 (O_470,N_2815,N_2922);
nand UO_471 (O_471,N_2964,N_2800);
xor UO_472 (O_472,N_2829,N_2993);
nand UO_473 (O_473,N_2910,N_2911);
or UO_474 (O_474,N_2902,N_2948);
nand UO_475 (O_475,N_2805,N_2836);
or UO_476 (O_476,N_2864,N_2828);
nor UO_477 (O_477,N_2910,N_2986);
and UO_478 (O_478,N_2860,N_2837);
nand UO_479 (O_479,N_2882,N_2840);
and UO_480 (O_480,N_2973,N_2808);
nor UO_481 (O_481,N_2913,N_2918);
nor UO_482 (O_482,N_2971,N_2903);
nor UO_483 (O_483,N_2930,N_2987);
or UO_484 (O_484,N_2965,N_2841);
or UO_485 (O_485,N_2949,N_2973);
nand UO_486 (O_486,N_2875,N_2955);
and UO_487 (O_487,N_2802,N_2913);
or UO_488 (O_488,N_2888,N_2910);
or UO_489 (O_489,N_2953,N_2983);
nor UO_490 (O_490,N_2871,N_2898);
and UO_491 (O_491,N_2965,N_2954);
and UO_492 (O_492,N_2842,N_2917);
nand UO_493 (O_493,N_2871,N_2849);
or UO_494 (O_494,N_2890,N_2934);
nand UO_495 (O_495,N_2916,N_2962);
nand UO_496 (O_496,N_2916,N_2971);
nor UO_497 (O_497,N_2944,N_2864);
nand UO_498 (O_498,N_2952,N_2966);
and UO_499 (O_499,N_2842,N_2843);
endmodule