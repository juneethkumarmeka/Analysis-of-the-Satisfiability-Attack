module basic_1000_10000_1500_2_levels_1xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5001,N_5003,N_5004,N_5005,N_5006,N_5007,N_5009,N_5011,N_5012,N_5013,N_5014,N_5018,N_5019,N_5021,N_5022,N_5023,N_5026,N_5027,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5039,N_5040,N_5041,N_5043,N_5047,N_5048,N_5050,N_5053,N_5054,N_5055,N_5056,N_5058,N_5060,N_5068,N_5069,N_5070,N_5071,N_5073,N_5074,N_5075,N_5077,N_5078,N_5079,N_5080,N_5083,N_5087,N_5088,N_5089,N_5090,N_5093,N_5094,N_5095,N_5096,N_5098,N_5099,N_5100,N_5101,N_5104,N_5106,N_5109,N_5111,N_5115,N_5117,N_5119,N_5120,N_5122,N_5128,N_5130,N_5134,N_5137,N_5139,N_5140,N_5141,N_5144,N_5146,N_5147,N_5148,N_5150,N_5152,N_5153,N_5154,N_5155,N_5158,N_5159,N_5160,N_5162,N_5164,N_5165,N_5167,N_5168,N_5169,N_5171,N_5172,N_5173,N_5174,N_5175,N_5179,N_5184,N_5187,N_5188,N_5189,N_5190,N_5191,N_5193,N_5194,N_5197,N_5199,N_5200,N_5201,N_5203,N_5205,N_5209,N_5210,N_5211,N_5212,N_5213,N_5215,N_5216,N_5218,N_5221,N_5223,N_5225,N_5226,N_5227,N_5228,N_5230,N_5232,N_5233,N_5235,N_5239,N_5241,N_5243,N_5244,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5255,N_5258,N_5261,N_5263,N_5267,N_5268,N_5272,N_5275,N_5277,N_5279,N_5280,N_5281,N_5284,N_5286,N_5287,N_5289,N_5290,N_5291,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5304,N_5305,N_5309,N_5310,N_5312,N_5313,N_5314,N_5315,N_5317,N_5319,N_5321,N_5324,N_5325,N_5327,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5352,N_5355,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5367,N_5368,N_5370,N_5372,N_5374,N_5375,N_5376,N_5379,N_5380,N_5381,N_5385,N_5386,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5400,N_5402,N_5403,N_5404,N_5406,N_5408,N_5412,N_5413,N_5414,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5425,N_5426,N_5428,N_5432,N_5436,N_5437,N_5439,N_5441,N_5442,N_5443,N_5445,N_5446,N_5449,N_5450,N_5451,N_5452,N_5454,N_5457,N_5458,N_5459,N_5462,N_5463,N_5464,N_5465,N_5468,N_5469,N_5470,N_5471,N_5472,N_5476,N_5477,N_5478,N_5480,N_5483,N_5484,N_5485,N_5491,N_5493,N_5494,N_5496,N_5498,N_5499,N_5501,N_5506,N_5507,N_5508,N_5510,N_5513,N_5516,N_5517,N_5518,N_5519,N_5521,N_5522,N_5523,N_5526,N_5527,N_5530,N_5531,N_5532,N_5536,N_5539,N_5540,N_5541,N_5543,N_5544,N_5546,N_5548,N_5551,N_5552,N_5554,N_5555,N_5556,N_5557,N_5558,N_5561,N_5563,N_5565,N_5566,N_5567,N_5569,N_5573,N_5574,N_5575,N_5576,N_5578,N_5580,N_5581,N_5584,N_5587,N_5589,N_5590,N_5592,N_5594,N_5599,N_5600,N_5603,N_5605,N_5608,N_5609,N_5611,N_5612,N_5613,N_5614,N_5618,N_5621,N_5622,N_5623,N_5625,N_5627,N_5628,N_5630,N_5632,N_5634,N_5635,N_5639,N_5640,N_5641,N_5644,N_5645,N_5646,N_5647,N_5649,N_5650,N_5652,N_5654,N_5655,N_5656,N_5657,N_5658,N_5662,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5671,N_5677,N_5680,N_5682,N_5683,N_5684,N_5685,N_5686,N_5689,N_5690,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5710,N_5711,N_5713,N_5714,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5725,N_5726,N_5727,N_5729,N_5732,N_5733,N_5734,N_5735,N_5737,N_5738,N_5739,N_5741,N_5742,N_5743,N_5744,N_5749,N_5750,N_5752,N_5753,N_5754,N_5756,N_5761,N_5762,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5772,N_5775,N_5776,N_5777,N_5778,N_5779,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5789,N_5790,N_5791,N_5792,N_5794,N_5796,N_5797,N_5798,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5808,N_5809,N_5810,N_5811,N_5812,N_5814,N_5815,N_5817,N_5820,N_5821,N_5823,N_5824,N_5826,N_5827,N_5829,N_5831,N_5833,N_5834,N_5837,N_5839,N_5840,N_5842,N_5844,N_5846,N_5847,N_5848,N_5849,N_5850,N_5852,N_5856,N_5857,N_5858,N_5859,N_5860,N_5862,N_5863,N_5864,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5873,N_5874,N_5877,N_5878,N_5880,N_5881,N_5883,N_5885,N_5887,N_5888,N_5889,N_5891,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5901,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5911,N_5912,N_5913,N_5914,N_5916,N_5918,N_5919,N_5920,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5930,N_5931,N_5934,N_5935,N_5938,N_5939,N_5940,N_5942,N_5943,N_5947,N_5948,N_5949,N_5951,N_5952,N_5953,N_5954,N_5955,N_5958,N_5959,N_5960,N_5963,N_5965,N_5966,N_5969,N_5970,N_5971,N_5972,N_5973,N_5975,N_5979,N_5981,N_5983,N_5984,N_5985,N_5986,N_5988,N_5990,N_5991,N_5992,N_5995,N_5997,N_5998,N_5999,N_6000,N_6002,N_6003,N_6004,N_6005,N_6008,N_6009,N_6011,N_6014,N_6015,N_6016,N_6017,N_6018,N_6020,N_6021,N_6023,N_6026,N_6027,N_6029,N_6031,N_6033,N_6034,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6043,N_6049,N_6050,N_6051,N_6052,N_6056,N_6057,N_6059,N_6061,N_6062,N_6064,N_6067,N_6069,N_6070,N_6072,N_6075,N_6077,N_6078,N_6079,N_6083,N_6085,N_6086,N_6088,N_6089,N_6090,N_6092,N_6093,N_6095,N_6098,N_6099,N_6101,N_6102,N_6103,N_6104,N_6107,N_6108,N_6109,N_6110,N_6112,N_6114,N_6115,N_6118,N_6119,N_6121,N_6125,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6145,N_6146,N_6147,N_6148,N_6150,N_6153,N_6154,N_6155,N_6156,N_6159,N_6160,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6169,N_6170,N_6173,N_6175,N_6177,N_6178,N_6180,N_6183,N_6184,N_6185,N_6186,N_6188,N_6189,N_6191,N_6193,N_6194,N_6196,N_6197,N_6198,N_6199,N_6200,N_6203,N_6204,N_6205,N_6207,N_6208,N_6211,N_6212,N_6213,N_6216,N_6217,N_6218,N_6219,N_6221,N_6222,N_6224,N_6225,N_6226,N_6227,N_6228,N_6234,N_6238,N_6239,N_6240,N_6241,N_6243,N_6244,N_6245,N_6246,N_6247,N_6249,N_6250,N_6251,N_6252,N_6254,N_6255,N_6257,N_6260,N_6261,N_6262,N_6263,N_6266,N_6268,N_6270,N_6271,N_6272,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6282,N_6283,N_6285,N_6286,N_6287,N_6291,N_6293,N_6300,N_6304,N_6305,N_6306,N_6308,N_6310,N_6311,N_6312,N_6317,N_6318,N_6320,N_6322,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6335,N_6338,N_6339,N_6340,N_6342,N_6343,N_6345,N_6346,N_6347,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6359,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6369,N_6370,N_6373,N_6374,N_6375,N_6377,N_6381,N_6382,N_6385,N_6388,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6404,N_6406,N_6408,N_6409,N_6410,N_6412,N_6415,N_6416,N_6417,N_6418,N_6419,N_6421,N_6423,N_6425,N_6429,N_6431,N_6432,N_6436,N_6437,N_6440,N_6441,N_6444,N_6449,N_6450,N_6452,N_6454,N_6455,N_6457,N_6459,N_6461,N_6463,N_6464,N_6466,N_6468,N_6469,N_6470,N_6473,N_6474,N_6475,N_6476,N_6478,N_6483,N_6485,N_6486,N_6487,N_6489,N_6491,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6502,N_6503,N_6505,N_6507,N_6508,N_6509,N_6511,N_6512,N_6513,N_6514,N_6518,N_6520,N_6522,N_6523,N_6524,N_6525,N_6526,N_6528,N_6529,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6539,N_6540,N_6541,N_6542,N_6544,N_6548,N_6549,N_6550,N_6553,N_6555,N_6556,N_6559,N_6560,N_6562,N_6565,N_6567,N_6568,N_6569,N_6570,N_6572,N_6573,N_6575,N_6577,N_6580,N_6581,N_6582,N_6583,N_6585,N_6586,N_6588,N_6589,N_6590,N_6593,N_6594,N_6597,N_6601,N_6603,N_6604,N_6608,N_6609,N_6611,N_6612,N_6614,N_6615,N_6616,N_6617,N_6620,N_6623,N_6624,N_6625,N_6626,N_6629,N_6635,N_6637,N_6638,N_6640,N_6641,N_6642,N_6643,N_6647,N_6648,N_6649,N_6651,N_6652,N_6653,N_6656,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6666,N_6667,N_6668,N_6669,N_6671,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6680,N_6681,N_6682,N_6683,N_6684,N_6686,N_6687,N_6688,N_6689,N_6691,N_6692,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6703,N_6704,N_6705,N_6706,N_6708,N_6710,N_6711,N_6712,N_6717,N_6718,N_6719,N_6720,N_6724,N_6726,N_6728,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6737,N_6738,N_6739,N_6740,N_6741,N_6745,N_6746,N_6749,N_6751,N_6752,N_6753,N_6756,N_6763,N_6766,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6782,N_6783,N_6784,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6796,N_6797,N_6798,N_6799,N_6800,N_6806,N_6807,N_6808,N_6810,N_6811,N_6813,N_6815,N_6816,N_6817,N_6818,N_6820,N_6821,N_6822,N_6823,N_6825,N_6826,N_6827,N_6829,N_6830,N_6831,N_6833,N_6834,N_6835,N_6837,N_6839,N_6840,N_6841,N_6843,N_6846,N_6848,N_6849,N_6850,N_6851,N_6853,N_6856,N_6859,N_6860,N_6861,N_6863,N_6867,N_6868,N_6870,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6882,N_6887,N_6890,N_6892,N_6893,N_6894,N_6895,N_6897,N_6898,N_6899,N_6901,N_6902,N_6903,N_6905,N_6906,N_6907,N_6912,N_6913,N_6915,N_6916,N_6918,N_6920,N_6923,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6941,N_6947,N_6949,N_6952,N_6953,N_6954,N_6956,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6968,N_6970,N_6975,N_6976,N_6979,N_6982,N_6983,N_6985,N_6986,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6998,N_6999,N_7000,N_7003,N_7005,N_7007,N_7009,N_7012,N_7014,N_7016,N_7017,N_7020,N_7021,N_7023,N_7024,N_7026,N_7027,N_7028,N_7029,N_7033,N_7037,N_7038,N_7040,N_7041,N_7042,N_7044,N_7046,N_7047,N_7048,N_7049,N_7051,N_7053,N_7054,N_7055,N_7056,N_7058,N_7059,N_7060,N_7062,N_7067,N_7070,N_7072,N_7075,N_7078,N_7079,N_7080,N_7081,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7095,N_7096,N_7097,N_7098,N_7099,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7108,N_7112,N_7113,N_7115,N_7117,N_7119,N_7120,N_7123,N_7124,N_7126,N_7127,N_7128,N_7129,N_7131,N_7132,N_7134,N_7137,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7147,N_7150,N_7151,N_7152,N_7153,N_7154,N_7156,N_7159,N_7160,N_7162,N_7164,N_7165,N_7166,N_7168,N_7170,N_7171,N_7172,N_7174,N_7175,N_7176,N_7179,N_7181,N_7182,N_7184,N_7185,N_7187,N_7190,N_7191,N_7197,N_7203,N_7205,N_7206,N_7209,N_7210,N_7212,N_7213,N_7215,N_7216,N_7217,N_7221,N_7222,N_7223,N_7224,N_7226,N_7228,N_7232,N_7235,N_7236,N_7237,N_7239,N_7240,N_7242,N_7243,N_7246,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7270,N_7272,N_7275,N_7277,N_7278,N_7280,N_7281,N_7282,N_7284,N_7285,N_7288,N_7289,N_7290,N_7292,N_7293,N_7295,N_7296,N_7297,N_7298,N_7300,N_7303,N_7304,N_7308,N_7309,N_7312,N_7314,N_7318,N_7319,N_7320,N_7322,N_7323,N_7324,N_7325,N_7327,N_7330,N_7331,N_7332,N_7333,N_7336,N_7337,N_7338,N_7340,N_7342,N_7348,N_7349,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7364,N_7365,N_7367,N_7368,N_7369,N_7370,N_7372,N_7373,N_7374,N_7375,N_7376,N_7378,N_7379,N_7380,N_7384,N_7385,N_7390,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7399,N_7401,N_7403,N_7404,N_7406,N_7408,N_7409,N_7410,N_7412,N_7413,N_7415,N_7416,N_7417,N_7419,N_7421,N_7423,N_7424,N_7425,N_7427,N_7429,N_7431,N_7432,N_7433,N_7435,N_7436,N_7438,N_7441,N_7442,N_7443,N_7445,N_7446,N_7447,N_7448,N_7450,N_7452,N_7453,N_7454,N_7455,N_7457,N_7458,N_7459,N_7461,N_7463,N_7464,N_7472,N_7473,N_7474,N_7475,N_7476,N_7478,N_7479,N_7481,N_7482,N_7483,N_7484,N_7485,N_7487,N_7491,N_7492,N_7493,N_7494,N_7496,N_7500,N_7502,N_7503,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7514,N_7515,N_7516,N_7517,N_7518,N_7524,N_7525,N_7526,N_7528,N_7529,N_7530,N_7531,N_7533,N_7535,N_7536,N_7538,N_7540,N_7541,N_7542,N_7548,N_7551,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7564,N_7567,N_7570,N_7572,N_7574,N_7575,N_7577,N_7578,N_7580,N_7581,N_7582,N_7584,N_7587,N_7589,N_7592,N_7593,N_7594,N_7596,N_7597,N_7600,N_7601,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7616,N_7618,N_7620,N_7621,N_7622,N_7625,N_7627,N_7628,N_7629,N_7631,N_7635,N_7636,N_7638,N_7640,N_7641,N_7643,N_7644,N_7645,N_7646,N_7648,N_7650,N_7651,N_7652,N_7653,N_7654,N_7656,N_7658,N_7659,N_7660,N_7662,N_7663,N_7666,N_7667,N_7668,N_7670,N_7671,N_7673,N_7676,N_7677,N_7678,N_7679,N_7680,N_7685,N_7686,N_7688,N_7689,N_7690,N_7691,N_7694,N_7695,N_7696,N_7697,N_7699,N_7701,N_7702,N_7703,N_7706,N_7709,N_7710,N_7711,N_7712,N_7713,N_7716,N_7717,N_7718,N_7719,N_7720,N_7722,N_7723,N_7724,N_7725,N_7726,N_7728,N_7730,N_7734,N_7735,N_7737,N_7740,N_7742,N_7743,N_7744,N_7746,N_7750,N_7751,N_7752,N_7753,N_7754,N_7758,N_7763,N_7764,N_7765,N_7770,N_7773,N_7774,N_7775,N_7776,N_7778,N_7779,N_7780,N_7783,N_7785,N_7788,N_7790,N_7793,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7809,N_7810,N_7811,N_7814,N_7815,N_7816,N_7817,N_7818,N_7820,N_7822,N_7826,N_7830,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7842,N_7843,N_7846,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7860,N_7861,N_7864,N_7866,N_7867,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7878,N_7883,N_7885,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7896,N_7898,N_7901,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7913,N_7915,N_7918,N_7920,N_7922,N_7924,N_7925,N_7926,N_7927,N_7930,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7946,N_7951,N_7952,N_7954,N_7957,N_7958,N_7964,N_7965,N_7966,N_7967,N_7969,N_7970,N_7971,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7980,N_7981,N_7985,N_7986,N_7987,N_7988,N_7989,N_7991,N_7992,N_7993,N_7994,N_7997,N_7998,N_7999,N_8001,N_8004,N_8008,N_8011,N_8012,N_8013,N_8015,N_8017,N_8018,N_8019,N_8023,N_8024,N_8025,N_8027,N_8028,N_8029,N_8030,N_8032,N_8034,N_8035,N_8037,N_8038,N_8039,N_8040,N_8042,N_8043,N_8045,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8061,N_8063,N_8065,N_8066,N_8067,N_8069,N_8073,N_8074,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8091,N_8092,N_8093,N_8094,N_8101,N_8103,N_8104,N_8106,N_8107,N_8112,N_8113,N_8114,N_8116,N_8120,N_8121,N_8123,N_8124,N_8125,N_8128,N_8130,N_8132,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8144,N_8145,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8154,N_8156,N_8157,N_8158,N_8159,N_8160,N_8163,N_8166,N_8167,N_8168,N_8169,N_8171,N_8172,N_8173,N_8174,N_8177,N_8178,N_8180,N_8184,N_8185,N_8187,N_8189,N_8190,N_8192,N_8195,N_8196,N_8197,N_8198,N_8203,N_8204,N_8205,N_8206,N_8208,N_8209,N_8210,N_8211,N_8215,N_8216,N_8218,N_8219,N_8221,N_8222,N_8224,N_8225,N_8228,N_8230,N_8234,N_8235,N_8236,N_8242,N_8243,N_8245,N_8246,N_8248,N_8250,N_8251,N_8252,N_8255,N_8256,N_8257,N_8258,N_8262,N_8263,N_8264,N_8269,N_8272,N_8273,N_8275,N_8276,N_8277,N_8282,N_8283,N_8284,N_8285,N_8289,N_8290,N_8293,N_8295,N_8304,N_8305,N_8306,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8323,N_8324,N_8325,N_8326,N_8328,N_8329,N_8331,N_8332,N_8334,N_8340,N_8341,N_8342,N_8343,N_8347,N_8348,N_8349,N_8350,N_8351,N_8353,N_8354,N_8355,N_8357,N_8359,N_8360,N_8361,N_8362,N_8365,N_8366,N_8367,N_8368,N_8369,N_8372,N_8373,N_8375,N_8378,N_8379,N_8383,N_8385,N_8387,N_8388,N_8390,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8400,N_8401,N_8402,N_8403,N_8406,N_8408,N_8409,N_8410,N_8412,N_8413,N_8415,N_8416,N_8418,N_8420,N_8422,N_8424,N_8425,N_8426,N_8427,N_8428,N_8430,N_8431,N_8433,N_8435,N_8436,N_8439,N_8442,N_8443,N_8445,N_8446,N_8447,N_8448,N_8449,N_8452,N_8453,N_8455,N_8463,N_8464,N_8466,N_8467,N_8468,N_8469,N_8470,N_8475,N_8476,N_8478,N_8479,N_8480,N_8481,N_8483,N_8484,N_8487,N_8489,N_8492,N_8496,N_8499,N_8502,N_8503,N_8505,N_8506,N_8507,N_8508,N_8510,N_8511,N_8512,N_8513,N_8516,N_8518,N_8519,N_8520,N_8521,N_8525,N_8526,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8536,N_8537,N_8542,N_8543,N_8547,N_8550,N_8551,N_8552,N_8557,N_8562,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8576,N_8578,N_8580,N_8581,N_8584,N_8586,N_8587,N_8589,N_8595,N_8596,N_8601,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8611,N_8614,N_8615,N_8616,N_8617,N_8620,N_8621,N_8622,N_8624,N_8625,N_8629,N_8630,N_8633,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8646,N_8649,N_8650,N_8651,N_8655,N_8656,N_8660,N_8661,N_8663,N_8664,N_8665,N_8667,N_8669,N_8670,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8680,N_8681,N_8683,N_8685,N_8687,N_8688,N_8689,N_8690,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8709,N_8710,N_8714,N_8719,N_8720,N_8723,N_8725,N_8727,N_8729,N_8730,N_8732,N_8734,N_8735,N_8737,N_8738,N_8739,N_8740,N_8742,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8753,N_8754,N_8755,N_8757,N_8758,N_8759,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8771,N_8775,N_8776,N_8777,N_8779,N_8780,N_8783,N_8785,N_8787,N_8790,N_8791,N_8792,N_8793,N_8794,N_8796,N_8797,N_8798,N_8799,N_8800,N_8802,N_8804,N_8807,N_8812,N_8813,N_8815,N_8816,N_8819,N_8821,N_8823,N_8825,N_8830,N_8831,N_8833,N_8835,N_8836,N_8837,N_8839,N_8840,N_8842,N_8844,N_8845,N_8847,N_8848,N_8849,N_8853,N_8855,N_8856,N_8858,N_8859,N_8861,N_8862,N_8865,N_8867,N_8868,N_8869,N_8870,N_8873,N_8874,N_8876,N_8877,N_8880,N_8882,N_8883,N_8884,N_8885,N_8887,N_8888,N_8889,N_8890,N_8891,N_8894,N_8895,N_8896,N_8899,N_8900,N_8901,N_8905,N_8906,N_8907,N_8908,N_8909,N_8911,N_8912,N_8914,N_8915,N_8916,N_8917,N_8920,N_8921,N_8923,N_8924,N_8926,N_8931,N_8932,N_8934,N_8938,N_8940,N_8942,N_8946,N_8948,N_8949,N_8950,N_8951,N_8954,N_8956,N_8958,N_8959,N_8961,N_8963,N_8964,N_8965,N_8967,N_8969,N_8971,N_8976,N_8977,N_8979,N_8980,N_8981,N_8983,N_8984,N_8985,N_8986,N_8987,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_9000,N_9001,N_9003,N_9004,N_9007,N_9012,N_9014,N_9015,N_9016,N_9017,N_9023,N_9024,N_9025,N_9026,N_9027,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9045,N_9047,N_9048,N_9050,N_9051,N_9052,N_9053,N_9056,N_9058,N_9059,N_9060,N_9061,N_9064,N_9065,N_9067,N_9068,N_9071,N_9073,N_9076,N_9080,N_9084,N_9085,N_9086,N_9087,N_9089,N_9090,N_9091,N_9093,N_9094,N_9095,N_9097,N_9098,N_9099,N_9101,N_9102,N_9103,N_9104,N_9107,N_9109,N_9110,N_9112,N_9114,N_9116,N_9119,N_9124,N_9126,N_9127,N_9129,N_9131,N_9132,N_9133,N_9135,N_9136,N_9137,N_9143,N_9144,N_9145,N_9147,N_9149,N_9150,N_9152,N_9153,N_9155,N_9157,N_9159,N_9160,N_9163,N_9164,N_9168,N_9170,N_9171,N_9172,N_9175,N_9178,N_9179,N_9181,N_9182,N_9184,N_9185,N_9186,N_9189,N_9190,N_9191,N_9192,N_9194,N_9195,N_9196,N_9198,N_9201,N_9203,N_9204,N_9206,N_9207,N_9208,N_9209,N_9212,N_9213,N_9215,N_9216,N_9220,N_9221,N_9222,N_9224,N_9225,N_9227,N_9228,N_9229,N_9231,N_9232,N_9233,N_9235,N_9236,N_9239,N_9240,N_9242,N_9245,N_9246,N_9247,N_9248,N_9250,N_9251,N_9252,N_9253,N_9254,N_9256,N_9257,N_9260,N_9261,N_9262,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9272,N_9273,N_9274,N_9276,N_9277,N_9278,N_9281,N_9284,N_9285,N_9287,N_9288,N_9291,N_9293,N_9294,N_9296,N_9297,N_9298,N_9300,N_9301,N_9302,N_9304,N_9305,N_9306,N_9313,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9323,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9336,N_9337,N_9338,N_9340,N_9341,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9353,N_9354,N_9356,N_9358,N_9359,N_9360,N_9362,N_9363,N_9364,N_9368,N_9369,N_9371,N_9373,N_9375,N_9380,N_9383,N_9384,N_9385,N_9387,N_9388,N_9391,N_9392,N_9395,N_9396,N_9398,N_9399,N_9401,N_9402,N_9403,N_9404,N_9406,N_9409,N_9410,N_9411,N_9413,N_9415,N_9418,N_9419,N_9420,N_9423,N_9424,N_9425,N_9426,N_9429,N_9430,N_9433,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9443,N_9444,N_9448,N_9449,N_9451,N_9452,N_9453,N_9455,N_9456,N_9457,N_9458,N_9462,N_9463,N_9465,N_9467,N_9470,N_9471,N_9472,N_9473,N_9479,N_9480,N_9482,N_9483,N_9485,N_9487,N_9489,N_9490,N_9491,N_9492,N_9495,N_9497,N_9498,N_9500,N_9501,N_9502,N_9505,N_9506,N_9507,N_9508,N_9510,N_9513,N_9514,N_9516,N_9517,N_9518,N_9520,N_9524,N_9525,N_9526,N_9528,N_9529,N_9531,N_9532,N_9533,N_9534,N_9535,N_9537,N_9539,N_9542,N_9543,N_9544,N_9550,N_9551,N_9553,N_9556,N_9557,N_9558,N_9559,N_9560,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9570,N_9571,N_9574,N_9575,N_9576,N_9578,N_9581,N_9582,N_9583,N_9584,N_9587,N_9588,N_9589,N_9590,N_9592,N_9594,N_9595,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9607,N_9609,N_9611,N_9612,N_9613,N_9615,N_9616,N_9618,N_9619,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9628,N_9629,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9640,N_9641,N_9642,N_9643,N_9644,N_9646,N_9647,N_9649,N_9651,N_9652,N_9653,N_9658,N_9661,N_9662,N_9663,N_9664,N_9667,N_9668,N_9669,N_9670,N_9673,N_9675,N_9677,N_9679,N_9681,N_9682,N_9684,N_9685,N_9686,N_9689,N_9690,N_9692,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9706,N_9709,N_9711,N_9712,N_9716,N_9717,N_9719,N_9723,N_9727,N_9728,N_9730,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9739,N_9740,N_9741,N_9742,N_9746,N_9747,N_9749,N_9750,N_9751,N_9753,N_9756,N_9757,N_9758,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9770,N_9773,N_9774,N_9775,N_9776,N_9777,N_9779,N_9780,N_9782,N_9783,N_9784,N_9787,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9798,N_9799,N_9800,N_9802,N_9803,N_9804,N_9805,N_9808,N_9809,N_9810,N_9812,N_9813,N_9814,N_9820,N_9821,N_9822,N_9823,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9835,N_9837,N_9838,N_9840,N_9841,N_9844,N_9846,N_9850,N_9851,N_9853,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9862,N_9863,N_9864,N_9865,N_9866,N_9868,N_9869,N_9870,N_9873,N_9875,N_9877,N_9878,N_9879,N_9881,N_9882,N_9883,N_9885,N_9888,N_9889,N_9890,N_9894,N_9897,N_9899,N_9900,N_9901,N_9903,N_9904,N_9907,N_9908,N_9909,N_9910,N_9911,N_9914,N_9915,N_9916,N_9917,N_9921,N_9922,N_9924,N_9926,N_9927,N_9933,N_9934,N_9937,N_9938,N_9939,N_9940,N_9941,N_9943,N_9944,N_9945,N_9946,N_9949,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9958,N_9959,N_9960,N_9961,N_9964,N_9965,N_9966,N_9967,N_9968,N_9970,N_9971,N_9973,N_9976,N_9977,N_9979,N_9980,N_9982,N_9983,N_9985,N_9986,N_9989,N_9991,N_9992,N_9993,N_9994,N_9996,N_9998;
or U0 (N_0,In_466,In_510);
nor U1 (N_1,In_696,In_802);
and U2 (N_2,In_552,In_343);
or U3 (N_3,In_747,In_783);
or U4 (N_4,In_849,In_250);
and U5 (N_5,In_560,In_483);
nor U6 (N_6,In_206,In_470);
nand U7 (N_7,In_698,In_799);
nand U8 (N_8,In_681,In_272);
nor U9 (N_9,In_388,In_356);
nand U10 (N_10,In_716,In_439);
nor U11 (N_11,In_848,In_122);
nand U12 (N_12,In_894,In_803);
xor U13 (N_13,In_676,In_685);
nor U14 (N_14,In_966,In_455);
nand U15 (N_15,In_986,In_598);
and U16 (N_16,In_571,In_958);
nand U17 (N_17,In_807,In_130);
or U18 (N_18,In_96,In_48);
nand U19 (N_19,In_132,In_302);
nor U20 (N_20,In_509,In_754);
or U21 (N_21,In_298,In_666);
and U22 (N_22,In_69,In_850);
nor U23 (N_23,In_836,In_151);
or U24 (N_24,In_921,In_284);
nor U25 (N_25,In_713,In_394);
nor U26 (N_26,In_294,In_753);
and U27 (N_27,In_901,In_399);
nand U28 (N_28,In_533,In_594);
and U29 (N_29,In_451,In_27);
and U30 (N_30,In_977,In_464);
or U31 (N_31,In_965,In_621);
nand U32 (N_32,In_605,In_667);
nand U33 (N_33,In_175,In_715);
nor U34 (N_34,In_236,In_588);
nor U35 (N_35,In_665,In_818);
nand U36 (N_36,In_89,In_830);
and U37 (N_37,In_490,In_804);
nand U38 (N_38,In_903,In_992);
nor U39 (N_39,In_949,In_65);
and U40 (N_40,In_165,In_37);
nand U41 (N_41,In_309,In_609);
or U42 (N_42,In_936,In_817);
or U43 (N_43,In_253,In_25);
nand U44 (N_44,In_735,In_737);
nand U45 (N_45,In_819,In_290);
or U46 (N_46,In_264,In_307);
or U47 (N_47,In_756,In_242);
nand U48 (N_48,In_154,In_127);
or U49 (N_49,In_377,In_978);
nand U50 (N_50,In_796,In_422);
nor U51 (N_51,In_235,In_502);
nand U52 (N_52,In_520,In_960);
and U53 (N_53,In_327,In_380);
or U54 (N_54,In_390,In_941);
nand U55 (N_55,In_305,In_900);
and U56 (N_56,In_712,In_346);
nor U57 (N_57,In_318,In_207);
nor U58 (N_58,In_874,In_219);
and U59 (N_59,In_869,In_320);
nand U60 (N_60,In_927,In_959);
nand U61 (N_61,In_654,In_963);
and U62 (N_62,In_904,In_391);
xnor U63 (N_63,In_924,In_945);
and U64 (N_64,In_722,In_335);
and U65 (N_65,In_672,In_248);
or U66 (N_66,In_909,In_131);
xor U67 (N_67,In_24,In_762);
nand U68 (N_68,In_185,In_745);
or U69 (N_69,In_679,In_220);
nor U70 (N_70,In_263,In_825);
nor U71 (N_71,In_508,In_191);
and U72 (N_72,In_554,In_543);
or U73 (N_73,In_613,In_694);
nand U74 (N_74,In_315,In_984);
nor U75 (N_75,In_54,In_650);
or U76 (N_76,In_92,In_695);
nor U77 (N_77,In_771,In_763);
nand U78 (N_78,In_143,In_243);
nor U79 (N_79,In_761,In_480);
or U80 (N_80,In_943,In_720);
or U81 (N_81,In_604,In_8);
nor U82 (N_82,In_736,In_174);
and U83 (N_83,In_912,In_893);
or U84 (N_84,In_216,In_854);
nand U85 (N_85,In_177,In_425);
nand U86 (N_86,In_190,In_488);
or U87 (N_87,In_378,In_196);
nand U88 (N_88,In_164,In_922);
nor U89 (N_89,In_557,In_475);
and U90 (N_90,In_463,In_222);
nor U91 (N_91,In_252,In_682);
nand U92 (N_92,In_512,In_393);
nor U93 (N_93,In_52,In_226);
nor U94 (N_94,In_786,In_66);
nand U95 (N_95,In_11,In_10);
and U96 (N_96,In_968,In_435);
nor U97 (N_97,In_778,In_962);
nor U98 (N_98,In_7,In_266);
and U99 (N_99,In_148,In_370);
nor U100 (N_100,In_249,In_576);
nand U101 (N_101,In_701,In_368);
and U102 (N_102,In_873,In_946);
and U103 (N_103,In_246,In_999);
nor U104 (N_104,In_119,In_511);
nor U105 (N_105,In_234,In_271);
or U106 (N_106,In_410,In_957);
nand U107 (N_107,In_45,In_531);
and U108 (N_108,In_919,In_723);
nand U109 (N_109,In_70,In_532);
nor U110 (N_110,In_28,In_467);
nor U111 (N_111,In_627,In_592);
nand U112 (N_112,In_505,In_428);
nand U113 (N_113,In_767,In_141);
nor U114 (N_114,In_633,In_260);
or U115 (N_115,In_332,In_831);
nor U116 (N_116,In_71,In_529);
nor U117 (N_117,In_379,In_350);
nor U118 (N_118,In_485,In_201);
nor U119 (N_119,In_245,In_82);
xnor U120 (N_120,In_16,In_67);
or U121 (N_121,In_183,In_482);
and U122 (N_122,In_306,In_926);
nor U123 (N_123,In_147,In_74);
nor U124 (N_124,In_351,In_619);
xor U125 (N_125,In_348,In_653);
and U126 (N_126,In_556,In_997);
and U127 (N_127,In_628,In_4);
and U128 (N_128,In_765,In_292);
and U129 (N_129,In_856,In_935);
and U130 (N_130,In_342,In_504);
nand U131 (N_131,In_417,In_659);
and U132 (N_132,In_107,In_411);
nor U133 (N_133,In_213,In_282);
and U134 (N_134,In_801,In_44);
nand U135 (N_135,In_905,In_300);
nor U136 (N_136,In_822,In_103);
nor U137 (N_137,In_883,In_133);
or U138 (N_138,In_80,In_610);
nor U139 (N_139,In_404,In_114);
nand U140 (N_140,In_558,In_779);
and U141 (N_141,In_734,In_721);
nand U142 (N_142,In_275,In_397);
or U143 (N_143,In_642,In_738);
nor U144 (N_144,In_303,In_365);
nor U145 (N_145,In_383,In_469);
or U146 (N_146,In_432,In_217);
nand U147 (N_147,In_987,In_261);
or U148 (N_148,In_583,In_669);
nor U149 (N_149,In_436,In_325);
nand U150 (N_150,In_0,In_995);
or U151 (N_151,In_857,In_707);
nor U152 (N_152,In_702,In_430);
xor U153 (N_153,In_193,In_474);
or U154 (N_154,In_887,In_139);
or U155 (N_155,In_150,In_892);
nand U156 (N_156,In_443,In_159);
nor U157 (N_157,In_398,In_537);
or U158 (N_158,In_889,In_684);
or U159 (N_159,In_412,In_415);
or U160 (N_160,In_814,In_21);
and U161 (N_161,In_730,In_157);
nor U162 (N_162,In_810,In_834);
xnor U163 (N_163,In_539,In_648);
nor U164 (N_164,In_372,In_182);
nand U165 (N_165,In_116,In_145);
or U166 (N_166,In_321,In_200);
and U167 (N_167,In_956,In_79);
nor U168 (N_168,In_352,In_991);
nand U169 (N_169,In_395,In_823);
nor U170 (N_170,In_240,In_798);
nand U171 (N_171,In_884,In_929);
nand U172 (N_172,In_354,In_998);
nor U173 (N_173,In_714,In_496);
nor U174 (N_174,In_852,In_188);
or U175 (N_175,In_517,In_812);
nor U176 (N_176,In_36,In_471);
or U177 (N_177,In_13,In_573);
nand U178 (N_178,In_746,In_33);
nor U179 (N_179,In_575,In_457);
or U180 (N_180,In_751,In_846);
nor U181 (N_181,In_711,In_358);
and U182 (N_182,In_495,In_414);
and U183 (N_183,In_643,In_420);
and U184 (N_184,In_224,In_600);
nand U185 (N_185,In_46,In_705);
nand U186 (N_186,In_581,In_149);
nor U187 (N_187,In_908,In_741);
and U188 (N_188,In_331,In_408);
and U189 (N_189,In_385,In_255);
nand U190 (N_190,In_59,In_5);
or U191 (N_191,In_547,In_38);
or U192 (N_192,In_838,In_17);
nand U193 (N_193,In_35,In_550);
nor U194 (N_194,In_247,In_877);
or U195 (N_195,In_522,In_835);
or U196 (N_196,In_211,In_259);
nor U197 (N_197,In_155,In_112);
nor U198 (N_198,In_384,In_775);
nor U199 (N_199,In_915,In_228);
nand U200 (N_200,In_872,In_890);
nand U201 (N_201,In_400,In_981);
nand U202 (N_202,In_800,In_225);
nand U203 (N_203,In_280,In_62);
or U204 (N_204,In_757,In_523);
or U205 (N_205,In_797,In_421);
xnor U206 (N_206,In_3,In_611);
and U207 (N_207,In_452,In_406);
and U208 (N_208,In_210,In_584);
and U209 (N_209,In_56,In_766);
or U210 (N_210,In_494,In_258);
nor U211 (N_211,In_947,In_974);
and U212 (N_212,In_47,In_123);
and U213 (N_213,In_140,In_833);
and U214 (N_214,In_661,In_268);
nand U215 (N_215,In_914,In_983);
nor U216 (N_216,In_693,In_301);
nand U217 (N_217,In_597,In_238);
nand U218 (N_218,In_545,In_973);
nand U219 (N_219,In_572,In_885);
or U220 (N_220,In_376,In_178);
or U221 (N_221,In_780,In_29);
or U222 (N_222,In_832,In_160);
nand U223 (N_223,In_287,In_19);
and U224 (N_224,In_506,In_691);
and U225 (N_225,In_99,In_186);
nor U226 (N_226,In_204,In_652);
and U227 (N_227,In_184,In_386);
nor U228 (N_228,In_326,In_134);
nor U229 (N_229,In_446,In_618);
nand U230 (N_230,In_990,In_706);
and U231 (N_231,In_784,In_476);
and U232 (N_232,In_938,In_278);
and U233 (N_233,In_456,In_808);
and U234 (N_234,In_192,In_758);
nor U235 (N_235,In_953,In_262);
nand U236 (N_236,In_683,In_18);
or U237 (N_237,In_121,In_357);
nor U238 (N_238,In_189,In_590);
nand U239 (N_239,In_733,In_719);
and U240 (N_240,In_606,In_923);
and U241 (N_241,In_478,In_308);
nor U242 (N_242,In_413,In_891);
nand U243 (N_243,In_270,In_668);
nor U244 (N_244,In_530,In_144);
and U245 (N_245,In_88,In_330);
nand U246 (N_246,In_438,In_86);
nor U247 (N_247,In_83,In_975);
and U248 (N_248,In_646,In_907);
nand U249 (N_249,In_366,In_678);
or U250 (N_250,In_434,In_813);
nand U251 (N_251,In_988,In_60);
nand U252 (N_252,In_755,In_473);
nand U253 (N_253,In_640,In_793);
nor U254 (N_254,In_445,In_273);
nor U255 (N_255,In_624,In_349);
nor U256 (N_256,In_146,In_886);
and U257 (N_257,In_548,In_498);
and U258 (N_258,In_871,In_631);
nand U259 (N_259,In_657,In_536);
or U260 (N_260,In_172,In_39);
nor U261 (N_261,In_795,In_739);
or U262 (N_262,In_928,In_513);
or U263 (N_263,In_340,In_969);
and U264 (N_264,In_944,In_860);
nand U265 (N_265,In_615,In_269);
or U266 (N_266,In_447,In_84);
nand U267 (N_267,In_125,In_105);
and U268 (N_268,In_534,In_528);
nor U269 (N_269,In_769,In_970);
or U270 (N_270,In_879,In_329);
nor U271 (N_271,In_524,In_897);
nor U272 (N_272,In_310,In_641);
nand U273 (N_273,In_954,In_867);
or U274 (N_274,In_790,In_102);
and U275 (N_275,In_9,In_396);
or U276 (N_276,In_768,In_51);
or U277 (N_277,In_369,In_527);
nor U278 (N_278,In_12,In_239);
nand U279 (N_279,In_14,In_544);
and U280 (N_280,In_820,In_840);
nor U281 (N_281,In_203,In_317);
or U282 (N_282,In_78,In_634);
and U283 (N_283,In_847,In_50);
nor U284 (N_284,In_43,In_541);
nor U285 (N_285,In_491,In_567);
nor U286 (N_286,In_937,In_658);
or U287 (N_287,In_197,In_782);
nand U288 (N_288,In_30,In_792);
or U289 (N_289,In_816,In_855);
nand U290 (N_290,In_176,In_128);
or U291 (N_291,In_709,In_285);
nor U292 (N_292,In_355,In_842);
or U293 (N_293,In_95,In_468);
and U294 (N_294,In_586,In_333);
nand U295 (N_295,In_662,In_26);
nor U296 (N_296,In_251,In_374);
nand U297 (N_297,In_49,In_209);
or U298 (N_298,In_568,In_811);
nor U299 (N_299,In_500,In_221);
or U300 (N_300,In_231,In_656);
nand U301 (N_301,In_697,In_664);
or U302 (N_302,In_853,In_507);
nor U303 (N_303,In_161,In_72);
and U304 (N_304,In_23,In_129);
or U305 (N_305,In_612,In_97);
nor U306 (N_306,In_426,In_794);
and U307 (N_307,In_862,In_942);
or U308 (N_308,In_806,In_731);
and U309 (N_309,In_93,In_677);
and U310 (N_310,In_162,In_781);
nand U311 (N_311,In_651,In_163);
or U312 (N_312,In_345,In_324);
nand U313 (N_313,In_126,In_437);
and U314 (N_314,In_87,In_827);
nand U315 (N_315,In_109,In_644);
and U316 (N_316,In_663,In_645);
or U317 (N_317,In_138,In_880);
nand U318 (N_318,In_313,In_760);
nor U319 (N_319,In_865,In_982);
or U320 (N_320,In_791,In_996);
nand U321 (N_321,In_334,In_717);
and U322 (N_322,In_993,In_787);
nand U323 (N_323,In_902,In_323);
or U324 (N_324,In_939,In_839);
and U325 (N_325,In_913,In_311);
nor U326 (N_326,In_295,In_68);
nand U327 (N_327,In_347,In_789);
nor U328 (N_328,In_578,In_106);
and U329 (N_329,In_90,In_589);
or U330 (N_330,In_700,In_637);
nor U331 (N_331,In_626,In_967);
nand U332 (N_332,In_214,In_538);
or U333 (N_333,In_950,In_77);
and U334 (N_334,In_636,In_85);
and U335 (N_335,In_980,In_896);
and U336 (N_336,In_405,In_608);
or U337 (N_337,In_32,In_828);
or U338 (N_338,In_647,In_487);
or U339 (N_339,In_462,In_110);
nand U340 (N_340,In_418,In_519);
nor U341 (N_341,In_732,In_551);
nand U342 (N_342,In_603,In_289);
nor U343 (N_343,In_459,In_6);
nand U344 (N_344,In_770,In_158);
nand U345 (N_345,In_244,In_314);
nand U346 (N_346,In_764,In_387);
or U347 (N_347,In_288,In_256);
nand U348 (N_348,In_866,In_441);
and U349 (N_349,In_501,In_20);
or U350 (N_350,In_934,In_607);
or U351 (N_351,In_440,In_843);
nor U352 (N_352,In_740,In_57);
nand U353 (N_353,In_2,In_265);
nand U354 (N_354,In_166,In_373);
and U355 (N_355,In_363,In_424);
nand U356 (N_356,In_687,In_409);
nand U357 (N_357,In_622,In_427);
nand U358 (N_358,In_382,In_632);
nor U359 (N_359,In_574,In_194);
nand U360 (N_360,In_599,In_444);
and U361 (N_361,In_1,In_930);
and U362 (N_362,In_918,In_76);
nor U363 (N_363,In_171,In_955);
xor U364 (N_364,In_844,In_602);
or U365 (N_365,In_776,In_863);
nor U366 (N_366,In_108,In_774);
nor U367 (N_367,In_864,In_202);
nand U368 (N_368,In_458,In_895);
and U369 (N_369,In_861,In_948);
nand U370 (N_370,In_859,In_585);
and U371 (N_371,In_788,In_341);
or U372 (N_372,In_888,In_337);
nand U373 (N_373,In_403,In_195);
xor U374 (N_374,In_875,In_223);
and U375 (N_375,In_296,In_479);
nor U376 (N_376,In_858,In_199);
and U377 (N_377,In_136,In_638);
and U378 (N_378,In_925,In_392);
nand U379 (N_379,In_777,In_15);
and U380 (N_380,In_281,In_117);
and U381 (N_381,In_829,In_821);
nand U382 (N_382,In_596,In_499);
and U383 (N_383,In_339,In_381);
nand U384 (N_384,In_233,In_579);
nor U385 (N_385,In_559,In_81);
nand U386 (N_386,In_449,In_629);
nand U387 (N_387,In_994,In_153);
nand U388 (N_388,In_870,In_570);
nand U389 (N_389,In_359,In_727);
xor U390 (N_390,In_279,In_218);
and U391 (N_391,In_364,In_688);
and U392 (N_392,In_362,In_64);
or U393 (N_393,In_477,In_91);
or U394 (N_394,In_120,In_553);
nor U395 (N_395,In_749,In_743);
and U396 (N_396,In_932,In_595);
nor U397 (N_397,In_113,In_673);
or U398 (N_398,In_58,In_277);
nor U399 (N_399,In_526,In_450);
and U400 (N_400,In_845,In_625);
and U401 (N_401,In_639,In_293);
and U402 (N_402,In_728,In_111);
nor U403 (N_403,In_124,In_976);
nor U404 (N_404,In_173,In_419);
nor U405 (N_405,In_100,In_267);
or U406 (N_406,In_851,In_503);
nand U407 (N_407,In_916,In_569);
nor U408 (N_408,In_115,In_461);
nand U409 (N_409,In_360,In_229);
or U410 (N_410,In_55,In_961);
and U411 (N_411,In_484,In_232);
nor U412 (N_412,In_623,In_336);
and U413 (N_413,In_492,In_972);
nor U414 (N_414,In_481,In_906);
and U415 (N_415,In_489,In_227);
nor U416 (N_416,In_416,In_152);
nand U417 (N_417,In_911,In_367);
or U418 (N_418,In_179,In_617);
nor U419 (N_419,In_101,In_910);
nor U420 (N_420,In_655,In_718);
nand U421 (N_421,In_565,In_274);
nand U422 (N_422,In_431,In_692);
or U423 (N_423,In_167,In_725);
nand U424 (N_424,In_952,In_40);
nand U425 (N_425,In_297,In_555);
or U426 (N_426,In_22,In_205);
nand U427 (N_427,In_375,In_472);
nand U428 (N_428,In_675,In_561);
nor U429 (N_429,In_402,In_841);
or U430 (N_430,In_772,In_591);
nor U431 (N_431,In_42,In_442);
nor U432 (N_432,In_516,In_94);
nor U433 (N_433,In_299,In_989);
or U434 (N_434,In_286,In_423);
and U435 (N_435,In_542,In_971);
and U436 (N_436,In_389,In_407);
or U437 (N_437,In_878,In_815);
nand U438 (N_438,In_493,In_180);
nor U439 (N_439,In_429,In_899);
and U440 (N_440,In_41,In_601);
and U441 (N_441,In_951,In_34);
and U442 (N_442,In_876,In_549);
and U443 (N_443,In_104,In_254);
nand U444 (N_444,In_933,In_708);
or U445 (N_445,In_620,In_118);
nor U446 (N_446,In_587,In_212);
or U447 (N_447,In_31,In_344);
nor U448 (N_448,In_742,In_785);
nand U449 (N_449,In_353,In_614);
nor U450 (N_450,In_460,In_312);
nand U451 (N_451,In_540,In_241);
nor U452 (N_452,In_710,In_168);
nor U453 (N_453,In_169,In_316);
nor U454 (N_454,In_257,In_497);
nor U455 (N_455,In_181,In_304);
or U456 (N_456,In_837,In_371);
nor U457 (N_457,In_454,In_724);
nand U458 (N_458,In_680,In_525);
nor U459 (N_459,In_898,In_291);
and U460 (N_460,In_660,In_616);
or U461 (N_461,In_649,In_518);
nand U462 (N_462,In_546,In_917);
nand U463 (N_463,In_748,In_674);
nand U464 (N_464,In_338,In_75);
or U465 (N_465,In_319,In_448);
or U466 (N_466,In_63,In_73);
and U467 (N_467,In_577,In_752);
xnor U468 (N_468,In_671,In_593);
nor U469 (N_469,In_135,In_198);
and U470 (N_470,In_773,In_759);
xor U471 (N_471,In_142,In_562);
nand U472 (N_472,In_670,In_322);
nand U473 (N_473,In_750,In_535);
nor U474 (N_474,In_703,In_726);
or U475 (N_475,In_979,In_187);
and U476 (N_476,In_208,In_563);
nand U477 (N_477,In_486,In_433);
or U478 (N_478,In_465,In_940);
and U479 (N_479,In_689,In_156);
xor U480 (N_480,In_729,In_920);
or U481 (N_481,In_985,In_635);
xnor U482 (N_482,In_686,In_170);
nand U483 (N_483,In_521,In_514);
nand U484 (N_484,In_630,In_805);
nor U485 (N_485,In_361,In_98);
and U486 (N_486,In_328,In_401);
and U487 (N_487,In_215,In_580);
nand U488 (N_488,In_453,In_61);
or U489 (N_489,In_137,In_931);
and U490 (N_490,In_53,In_566);
nand U491 (N_491,In_276,In_826);
nand U492 (N_492,In_230,In_868);
nand U493 (N_493,In_690,In_515);
nor U494 (N_494,In_237,In_824);
and U495 (N_495,In_582,In_882);
or U496 (N_496,In_564,In_809);
nor U497 (N_497,In_283,In_704);
nor U498 (N_498,In_964,In_881);
nor U499 (N_499,In_699,In_744);
or U500 (N_500,In_342,In_410);
nor U501 (N_501,In_495,In_380);
nand U502 (N_502,In_980,In_696);
and U503 (N_503,In_624,In_715);
nand U504 (N_504,In_169,In_357);
xor U505 (N_505,In_130,In_348);
and U506 (N_506,In_268,In_889);
and U507 (N_507,In_539,In_817);
nor U508 (N_508,In_830,In_439);
nand U509 (N_509,In_649,In_225);
nand U510 (N_510,In_476,In_274);
nor U511 (N_511,In_956,In_374);
nand U512 (N_512,In_33,In_145);
nor U513 (N_513,In_810,In_386);
and U514 (N_514,In_128,In_653);
and U515 (N_515,In_897,In_466);
and U516 (N_516,In_703,In_372);
or U517 (N_517,In_962,In_681);
and U518 (N_518,In_922,In_491);
nor U519 (N_519,In_863,In_902);
nor U520 (N_520,In_991,In_924);
and U521 (N_521,In_400,In_979);
nor U522 (N_522,In_148,In_593);
or U523 (N_523,In_986,In_343);
nor U524 (N_524,In_965,In_310);
nand U525 (N_525,In_422,In_786);
nor U526 (N_526,In_578,In_844);
or U527 (N_527,In_935,In_340);
or U528 (N_528,In_677,In_100);
or U529 (N_529,In_463,In_816);
nand U530 (N_530,In_898,In_745);
and U531 (N_531,In_834,In_289);
or U532 (N_532,In_539,In_871);
nand U533 (N_533,In_991,In_167);
or U534 (N_534,In_265,In_334);
or U535 (N_535,In_263,In_630);
nand U536 (N_536,In_13,In_830);
xnor U537 (N_537,In_321,In_165);
xnor U538 (N_538,In_705,In_289);
and U539 (N_539,In_88,In_712);
nor U540 (N_540,In_56,In_209);
and U541 (N_541,In_832,In_139);
and U542 (N_542,In_805,In_747);
and U543 (N_543,In_614,In_750);
or U544 (N_544,In_248,In_915);
or U545 (N_545,In_625,In_881);
and U546 (N_546,In_250,In_819);
nand U547 (N_547,In_769,In_660);
nor U548 (N_548,In_57,In_584);
or U549 (N_549,In_328,In_393);
nor U550 (N_550,In_450,In_554);
nor U551 (N_551,In_167,In_339);
nor U552 (N_552,In_138,In_248);
nor U553 (N_553,In_642,In_771);
or U554 (N_554,In_864,In_493);
and U555 (N_555,In_661,In_818);
nor U556 (N_556,In_128,In_599);
nor U557 (N_557,In_460,In_232);
nor U558 (N_558,In_533,In_335);
and U559 (N_559,In_995,In_377);
nor U560 (N_560,In_551,In_816);
and U561 (N_561,In_708,In_205);
nand U562 (N_562,In_380,In_205);
nor U563 (N_563,In_904,In_483);
nand U564 (N_564,In_120,In_473);
nand U565 (N_565,In_713,In_223);
and U566 (N_566,In_213,In_564);
nor U567 (N_567,In_551,In_232);
nand U568 (N_568,In_152,In_289);
and U569 (N_569,In_547,In_147);
nor U570 (N_570,In_402,In_320);
nor U571 (N_571,In_844,In_791);
or U572 (N_572,In_888,In_163);
or U573 (N_573,In_111,In_635);
or U574 (N_574,In_166,In_947);
or U575 (N_575,In_496,In_612);
or U576 (N_576,In_385,In_991);
nand U577 (N_577,In_227,In_97);
nand U578 (N_578,In_576,In_873);
and U579 (N_579,In_894,In_150);
nor U580 (N_580,In_611,In_439);
or U581 (N_581,In_387,In_691);
nand U582 (N_582,In_302,In_100);
nor U583 (N_583,In_957,In_947);
nand U584 (N_584,In_598,In_641);
or U585 (N_585,In_592,In_385);
nand U586 (N_586,In_869,In_47);
nand U587 (N_587,In_127,In_519);
nand U588 (N_588,In_476,In_943);
nor U589 (N_589,In_971,In_154);
nand U590 (N_590,In_470,In_8);
nor U591 (N_591,In_505,In_487);
nand U592 (N_592,In_156,In_85);
nand U593 (N_593,In_799,In_628);
nor U594 (N_594,In_918,In_492);
or U595 (N_595,In_626,In_883);
nand U596 (N_596,In_501,In_189);
nor U597 (N_597,In_667,In_869);
nand U598 (N_598,In_784,In_980);
and U599 (N_599,In_898,In_932);
nor U600 (N_600,In_906,In_846);
and U601 (N_601,In_670,In_733);
or U602 (N_602,In_5,In_304);
nor U603 (N_603,In_867,In_362);
or U604 (N_604,In_711,In_314);
and U605 (N_605,In_174,In_839);
or U606 (N_606,In_150,In_336);
nand U607 (N_607,In_962,In_481);
and U608 (N_608,In_113,In_402);
and U609 (N_609,In_926,In_566);
nand U610 (N_610,In_971,In_338);
and U611 (N_611,In_619,In_333);
or U612 (N_612,In_813,In_271);
nor U613 (N_613,In_745,In_235);
or U614 (N_614,In_65,In_867);
and U615 (N_615,In_898,In_649);
nand U616 (N_616,In_591,In_266);
and U617 (N_617,In_944,In_134);
and U618 (N_618,In_22,In_302);
nand U619 (N_619,In_457,In_729);
and U620 (N_620,In_865,In_743);
nor U621 (N_621,In_450,In_78);
nand U622 (N_622,In_652,In_320);
nor U623 (N_623,In_958,In_466);
nor U624 (N_624,In_531,In_841);
and U625 (N_625,In_204,In_890);
xnor U626 (N_626,In_87,In_764);
and U627 (N_627,In_343,In_901);
or U628 (N_628,In_809,In_966);
and U629 (N_629,In_898,In_586);
nor U630 (N_630,In_564,In_908);
and U631 (N_631,In_664,In_606);
or U632 (N_632,In_289,In_166);
nand U633 (N_633,In_267,In_694);
nand U634 (N_634,In_86,In_904);
nand U635 (N_635,In_316,In_927);
or U636 (N_636,In_393,In_508);
nand U637 (N_637,In_273,In_829);
nor U638 (N_638,In_679,In_599);
nor U639 (N_639,In_511,In_261);
nor U640 (N_640,In_239,In_929);
and U641 (N_641,In_281,In_191);
nor U642 (N_642,In_804,In_637);
or U643 (N_643,In_963,In_505);
or U644 (N_644,In_407,In_71);
or U645 (N_645,In_14,In_886);
or U646 (N_646,In_578,In_298);
nand U647 (N_647,In_889,In_893);
or U648 (N_648,In_754,In_762);
and U649 (N_649,In_604,In_778);
nor U650 (N_650,In_854,In_361);
nand U651 (N_651,In_508,In_43);
and U652 (N_652,In_648,In_894);
and U653 (N_653,In_595,In_953);
nor U654 (N_654,In_201,In_63);
or U655 (N_655,In_429,In_924);
and U656 (N_656,In_528,In_97);
nor U657 (N_657,In_549,In_150);
and U658 (N_658,In_507,In_623);
or U659 (N_659,In_830,In_787);
nand U660 (N_660,In_931,In_510);
or U661 (N_661,In_655,In_143);
nand U662 (N_662,In_393,In_778);
nor U663 (N_663,In_235,In_303);
or U664 (N_664,In_16,In_207);
and U665 (N_665,In_141,In_145);
nand U666 (N_666,In_6,In_443);
and U667 (N_667,In_225,In_929);
nor U668 (N_668,In_524,In_440);
or U669 (N_669,In_691,In_149);
nand U670 (N_670,In_85,In_167);
nor U671 (N_671,In_833,In_613);
nand U672 (N_672,In_515,In_198);
or U673 (N_673,In_174,In_302);
and U674 (N_674,In_928,In_327);
or U675 (N_675,In_947,In_718);
and U676 (N_676,In_913,In_962);
nor U677 (N_677,In_707,In_68);
or U678 (N_678,In_950,In_716);
nand U679 (N_679,In_726,In_797);
nand U680 (N_680,In_584,In_787);
nand U681 (N_681,In_667,In_268);
nor U682 (N_682,In_764,In_449);
or U683 (N_683,In_67,In_316);
nand U684 (N_684,In_37,In_127);
nand U685 (N_685,In_573,In_903);
and U686 (N_686,In_362,In_337);
nor U687 (N_687,In_290,In_921);
nor U688 (N_688,In_356,In_521);
and U689 (N_689,In_184,In_232);
nor U690 (N_690,In_400,In_666);
and U691 (N_691,In_140,In_192);
nor U692 (N_692,In_743,In_863);
nand U693 (N_693,In_331,In_73);
nand U694 (N_694,In_833,In_477);
xor U695 (N_695,In_882,In_600);
or U696 (N_696,In_641,In_539);
or U697 (N_697,In_351,In_154);
and U698 (N_698,In_181,In_814);
or U699 (N_699,In_800,In_8);
nor U700 (N_700,In_345,In_549);
nor U701 (N_701,In_399,In_624);
nor U702 (N_702,In_227,In_924);
or U703 (N_703,In_961,In_786);
nand U704 (N_704,In_716,In_652);
nand U705 (N_705,In_312,In_159);
nand U706 (N_706,In_844,In_571);
and U707 (N_707,In_8,In_337);
or U708 (N_708,In_184,In_931);
nand U709 (N_709,In_381,In_669);
nand U710 (N_710,In_555,In_516);
and U711 (N_711,In_719,In_891);
nand U712 (N_712,In_648,In_497);
nor U713 (N_713,In_836,In_737);
nor U714 (N_714,In_683,In_227);
or U715 (N_715,In_295,In_709);
nor U716 (N_716,In_824,In_828);
or U717 (N_717,In_97,In_590);
nand U718 (N_718,In_126,In_424);
nand U719 (N_719,In_423,In_455);
nor U720 (N_720,In_319,In_442);
nand U721 (N_721,In_343,In_996);
nor U722 (N_722,In_816,In_395);
or U723 (N_723,In_763,In_118);
nand U724 (N_724,In_605,In_719);
nand U725 (N_725,In_610,In_541);
or U726 (N_726,In_475,In_889);
and U727 (N_727,In_130,In_855);
and U728 (N_728,In_650,In_475);
nor U729 (N_729,In_635,In_399);
and U730 (N_730,In_63,In_399);
and U731 (N_731,In_282,In_801);
or U732 (N_732,In_239,In_28);
nand U733 (N_733,In_33,In_438);
and U734 (N_734,In_906,In_274);
and U735 (N_735,In_285,In_630);
xnor U736 (N_736,In_852,In_800);
nand U737 (N_737,In_273,In_555);
or U738 (N_738,In_434,In_504);
and U739 (N_739,In_976,In_801);
or U740 (N_740,In_740,In_810);
and U741 (N_741,In_674,In_639);
nor U742 (N_742,In_148,In_902);
nand U743 (N_743,In_577,In_653);
or U744 (N_744,In_285,In_394);
nand U745 (N_745,In_55,In_586);
nor U746 (N_746,In_610,In_939);
or U747 (N_747,In_167,In_203);
xor U748 (N_748,In_627,In_280);
nor U749 (N_749,In_1,In_984);
and U750 (N_750,In_617,In_211);
and U751 (N_751,In_182,In_559);
or U752 (N_752,In_115,In_125);
nor U753 (N_753,In_863,In_592);
nand U754 (N_754,In_157,In_15);
and U755 (N_755,In_246,In_644);
nand U756 (N_756,In_122,In_783);
and U757 (N_757,In_471,In_98);
nor U758 (N_758,In_585,In_410);
nor U759 (N_759,In_771,In_947);
and U760 (N_760,In_785,In_22);
and U761 (N_761,In_360,In_325);
and U762 (N_762,In_699,In_870);
nor U763 (N_763,In_69,In_214);
nor U764 (N_764,In_897,In_962);
nor U765 (N_765,In_344,In_207);
and U766 (N_766,In_678,In_74);
or U767 (N_767,In_179,In_724);
or U768 (N_768,In_214,In_670);
nor U769 (N_769,In_232,In_829);
and U770 (N_770,In_133,In_23);
or U771 (N_771,In_337,In_508);
and U772 (N_772,In_858,In_580);
nor U773 (N_773,In_874,In_674);
nand U774 (N_774,In_15,In_356);
and U775 (N_775,In_36,In_940);
and U776 (N_776,In_669,In_45);
and U777 (N_777,In_419,In_562);
or U778 (N_778,In_190,In_883);
nand U779 (N_779,In_654,In_727);
nor U780 (N_780,In_352,In_866);
nand U781 (N_781,In_88,In_857);
or U782 (N_782,In_94,In_834);
nand U783 (N_783,In_385,In_940);
or U784 (N_784,In_562,In_867);
nor U785 (N_785,In_192,In_100);
nand U786 (N_786,In_20,In_972);
and U787 (N_787,In_943,In_233);
nor U788 (N_788,In_522,In_291);
nor U789 (N_789,In_663,In_263);
or U790 (N_790,In_600,In_866);
nand U791 (N_791,In_808,In_677);
nand U792 (N_792,In_628,In_752);
nand U793 (N_793,In_284,In_408);
nand U794 (N_794,In_847,In_17);
nand U795 (N_795,In_598,In_78);
nand U796 (N_796,In_712,In_742);
or U797 (N_797,In_949,In_92);
nand U798 (N_798,In_15,In_617);
and U799 (N_799,In_840,In_509);
nand U800 (N_800,In_845,In_633);
and U801 (N_801,In_950,In_580);
and U802 (N_802,In_485,In_650);
nand U803 (N_803,In_669,In_634);
nor U804 (N_804,In_975,In_851);
nand U805 (N_805,In_236,In_773);
nor U806 (N_806,In_851,In_50);
nor U807 (N_807,In_359,In_768);
nor U808 (N_808,In_440,In_391);
or U809 (N_809,In_963,In_101);
and U810 (N_810,In_420,In_282);
nor U811 (N_811,In_985,In_395);
nor U812 (N_812,In_219,In_977);
or U813 (N_813,In_402,In_14);
nor U814 (N_814,In_154,In_107);
or U815 (N_815,In_146,In_678);
and U816 (N_816,In_203,In_982);
or U817 (N_817,In_428,In_50);
nor U818 (N_818,In_507,In_399);
nor U819 (N_819,In_589,In_508);
and U820 (N_820,In_888,In_224);
or U821 (N_821,In_586,In_588);
or U822 (N_822,In_46,In_855);
and U823 (N_823,In_191,In_559);
nand U824 (N_824,In_156,In_650);
and U825 (N_825,In_432,In_580);
nand U826 (N_826,In_37,In_719);
nor U827 (N_827,In_401,In_667);
nor U828 (N_828,In_744,In_428);
and U829 (N_829,In_644,In_410);
nand U830 (N_830,In_636,In_231);
nand U831 (N_831,In_153,In_668);
or U832 (N_832,In_861,In_102);
and U833 (N_833,In_817,In_222);
nor U834 (N_834,In_783,In_594);
nor U835 (N_835,In_939,In_190);
or U836 (N_836,In_484,In_304);
and U837 (N_837,In_112,In_394);
and U838 (N_838,In_883,In_785);
nor U839 (N_839,In_662,In_577);
xor U840 (N_840,In_772,In_135);
nor U841 (N_841,In_817,In_745);
nor U842 (N_842,In_621,In_779);
nand U843 (N_843,In_250,In_103);
or U844 (N_844,In_55,In_247);
and U845 (N_845,In_224,In_13);
or U846 (N_846,In_991,In_903);
nor U847 (N_847,In_848,In_116);
and U848 (N_848,In_870,In_565);
xor U849 (N_849,In_449,In_179);
or U850 (N_850,In_137,In_907);
or U851 (N_851,In_529,In_627);
or U852 (N_852,In_897,In_181);
nor U853 (N_853,In_788,In_814);
and U854 (N_854,In_498,In_652);
xnor U855 (N_855,In_219,In_636);
xnor U856 (N_856,In_981,In_179);
nor U857 (N_857,In_647,In_0);
and U858 (N_858,In_310,In_477);
nand U859 (N_859,In_868,In_430);
nor U860 (N_860,In_231,In_410);
nand U861 (N_861,In_757,In_712);
and U862 (N_862,In_476,In_183);
and U863 (N_863,In_564,In_148);
and U864 (N_864,In_842,In_201);
and U865 (N_865,In_681,In_723);
or U866 (N_866,In_279,In_189);
nor U867 (N_867,In_230,In_452);
or U868 (N_868,In_604,In_492);
nor U869 (N_869,In_264,In_329);
nand U870 (N_870,In_333,In_894);
nor U871 (N_871,In_561,In_68);
or U872 (N_872,In_382,In_777);
and U873 (N_873,In_515,In_217);
nand U874 (N_874,In_967,In_52);
nand U875 (N_875,In_473,In_921);
nand U876 (N_876,In_319,In_343);
or U877 (N_877,In_591,In_824);
nand U878 (N_878,In_783,In_456);
and U879 (N_879,In_545,In_805);
and U880 (N_880,In_574,In_185);
nand U881 (N_881,In_15,In_289);
nor U882 (N_882,In_610,In_289);
nand U883 (N_883,In_27,In_860);
nand U884 (N_884,In_274,In_178);
nand U885 (N_885,In_731,In_224);
and U886 (N_886,In_764,In_885);
nor U887 (N_887,In_862,In_569);
or U888 (N_888,In_223,In_804);
and U889 (N_889,In_667,In_88);
nand U890 (N_890,In_181,In_343);
nand U891 (N_891,In_459,In_981);
nor U892 (N_892,In_317,In_567);
or U893 (N_893,In_803,In_60);
nand U894 (N_894,In_693,In_291);
nor U895 (N_895,In_93,In_536);
nor U896 (N_896,In_643,In_125);
nand U897 (N_897,In_486,In_808);
and U898 (N_898,In_561,In_893);
or U899 (N_899,In_865,In_838);
and U900 (N_900,In_137,In_175);
nor U901 (N_901,In_700,In_339);
nand U902 (N_902,In_310,In_692);
and U903 (N_903,In_257,In_65);
or U904 (N_904,In_240,In_750);
nand U905 (N_905,In_218,In_503);
nand U906 (N_906,In_298,In_690);
nand U907 (N_907,In_648,In_231);
and U908 (N_908,In_12,In_667);
and U909 (N_909,In_875,In_3);
nand U910 (N_910,In_709,In_873);
nand U911 (N_911,In_120,In_107);
nor U912 (N_912,In_203,In_113);
and U913 (N_913,In_839,In_118);
and U914 (N_914,In_508,In_338);
xnor U915 (N_915,In_675,In_957);
or U916 (N_916,In_922,In_707);
and U917 (N_917,In_157,In_126);
nor U918 (N_918,In_1,In_464);
and U919 (N_919,In_767,In_362);
nor U920 (N_920,In_837,In_372);
and U921 (N_921,In_299,In_393);
nor U922 (N_922,In_170,In_177);
nand U923 (N_923,In_214,In_499);
or U924 (N_924,In_335,In_164);
nor U925 (N_925,In_39,In_517);
and U926 (N_926,In_401,In_353);
or U927 (N_927,In_474,In_781);
or U928 (N_928,In_271,In_884);
nand U929 (N_929,In_112,In_252);
or U930 (N_930,In_625,In_846);
nand U931 (N_931,In_333,In_52);
or U932 (N_932,In_174,In_377);
and U933 (N_933,In_417,In_256);
nor U934 (N_934,In_833,In_176);
and U935 (N_935,In_342,In_487);
nor U936 (N_936,In_150,In_27);
nand U937 (N_937,In_904,In_702);
nor U938 (N_938,In_286,In_692);
and U939 (N_939,In_293,In_569);
nand U940 (N_940,In_625,In_879);
nor U941 (N_941,In_9,In_497);
and U942 (N_942,In_147,In_54);
or U943 (N_943,In_574,In_149);
nor U944 (N_944,In_386,In_542);
nand U945 (N_945,In_686,In_990);
and U946 (N_946,In_240,In_592);
and U947 (N_947,In_847,In_326);
nor U948 (N_948,In_733,In_58);
or U949 (N_949,In_974,In_817);
nand U950 (N_950,In_619,In_924);
or U951 (N_951,In_390,In_367);
nor U952 (N_952,In_21,In_970);
or U953 (N_953,In_671,In_624);
nor U954 (N_954,In_899,In_892);
and U955 (N_955,In_381,In_668);
and U956 (N_956,In_627,In_18);
and U957 (N_957,In_186,In_849);
nor U958 (N_958,In_32,In_685);
or U959 (N_959,In_114,In_251);
nand U960 (N_960,In_384,In_297);
nor U961 (N_961,In_454,In_168);
and U962 (N_962,In_756,In_802);
nand U963 (N_963,In_950,In_566);
and U964 (N_964,In_130,In_678);
and U965 (N_965,In_356,In_819);
or U966 (N_966,In_921,In_191);
and U967 (N_967,In_664,In_98);
nor U968 (N_968,In_999,In_788);
and U969 (N_969,In_350,In_329);
or U970 (N_970,In_629,In_263);
or U971 (N_971,In_173,In_60);
or U972 (N_972,In_489,In_226);
nand U973 (N_973,In_991,In_848);
or U974 (N_974,In_721,In_573);
nand U975 (N_975,In_765,In_819);
or U976 (N_976,In_832,In_300);
or U977 (N_977,In_993,In_917);
nand U978 (N_978,In_722,In_514);
nand U979 (N_979,In_730,In_430);
or U980 (N_980,In_846,In_142);
nor U981 (N_981,In_944,In_369);
or U982 (N_982,In_119,In_940);
nand U983 (N_983,In_827,In_994);
nand U984 (N_984,In_501,In_198);
or U985 (N_985,In_789,In_668);
or U986 (N_986,In_801,In_383);
nand U987 (N_987,In_552,In_215);
or U988 (N_988,In_688,In_2);
nor U989 (N_989,In_678,In_804);
nand U990 (N_990,In_563,In_597);
nand U991 (N_991,In_639,In_482);
nor U992 (N_992,In_693,In_819);
or U993 (N_993,In_802,In_614);
nand U994 (N_994,In_394,In_565);
and U995 (N_995,In_744,In_846);
and U996 (N_996,In_270,In_620);
xor U997 (N_997,In_739,In_911);
nand U998 (N_998,In_812,In_320);
nand U999 (N_999,In_112,In_524);
nand U1000 (N_1000,In_263,In_218);
or U1001 (N_1001,In_316,In_588);
or U1002 (N_1002,In_213,In_800);
or U1003 (N_1003,In_848,In_977);
and U1004 (N_1004,In_629,In_948);
nand U1005 (N_1005,In_988,In_454);
nand U1006 (N_1006,In_442,In_163);
nand U1007 (N_1007,In_262,In_835);
and U1008 (N_1008,In_791,In_572);
or U1009 (N_1009,In_135,In_220);
xnor U1010 (N_1010,In_244,In_472);
and U1011 (N_1011,In_545,In_688);
nand U1012 (N_1012,In_789,In_644);
or U1013 (N_1013,In_745,In_404);
nor U1014 (N_1014,In_468,In_699);
nand U1015 (N_1015,In_193,In_736);
nand U1016 (N_1016,In_598,In_975);
and U1017 (N_1017,In_945,In_677);
nor U1018 (N_1018,In_456,In_21);
nor U1019 (N_1019,In_830,In_38);
and U1020 (N_1020,In_74,In_1);
and U1021 (N_1021,In_873,In_812);
nor U1022 (N_1022,In_306,In_766);
xor U1023 (N_1023,In_375,In_320);
nand U1024 (N_1024,In_276,In_422);
nand U1025 (N_1025,In_376,In_281);
or U1026 (N_1026,In_337,In_447);
and U1027 (N_1027,In_478,In_189);
or U1028 (N_1028,In_415,In_759);
xnor U1029 (N_1029,In_691,In_620);
nor U1030 (N_1030,In_970,In_828);
nor U1031 (N_1031,In_645,In_648);
and U1032 (N_1032,In_77,In_271);
nand U1033 (N_1033,In_88,In_688);
nor U1034 (N_1034,In_606,In_14);
or U1035 (N_1035,In_444,In_417);
nor U1036 (N_1036,In_417,In_209);
nor U1037 (N_1037,In_861,In_680);
or U1038 (N_1038,In_745,In_881);
and U1039 (N_1039,In_583,In_753);
and U1040 (N_1040,In_83,In_413);
nand U1041 (N_1041,In_515,In_462);
nor U1042 (N_1042,In_913,In_409);
nand U1043 (N_1043,In_391,In_857);
or U1044 (N_1044,In_822,In_129);
and U1045 (N_1045,In_829,In_144);
and U1046 (N_1046,In_513,In_178);
nor U1047 (N_1047,In_474,In_175);
nor U1048 (N_1048,In_770,In_214);
nor U1049 (N_1049,In_773,In_893);
nor U1050 (N_1050,In_767,In_981);
and U1051 (N_1051,In_922,In_761);
and U1052 (N_1052,In_871,In_364);
nand U1053 (N_1053,In_753,In_399);
or U1054 (N_1054,In_624,In_447);
nand U1055 (N_1055,In_6,In_184);
nor U1056 (N_1056,In_82,In_761);
and U1057 (N_1057,In_390,In_705);
and U1058 (N_1058,In_636,In_853);
nor U1059 (N_1059,In_348,In_566);
nand U1060 (N_1060,In_575,In_949);
or U1061 (N_1061,In_289,In_928);
nor U1062 (N_1062,In_45,In_78);
and U1063 (N_1063,In_550,In_449);
or U1064 (N_1064,In_275,In_893);
nor U1065 (N_1065,In_799,In_160);
nor U1066 (N_1066,In_138,In_986);
nand U1067 (N_1067,In_759,In_780);
nor U1068 (N_1068,In_519,In_31);
nand U1069 (N_1069,In_305,In_472);
and U1070 (N_1070,In_162,In_400);
or U1071 (N_1071,In_840,In_537);
nor U1072 (N_1072,In_214,In_587);
and U1073 (N_1073,In_129,In_274);
and U1074 (N_1074,In_369,In_385);
nand U1075 (N_1075,In_727,In_89);
nand U1076 (N_1076,In_142,In_794);
or U1077 (N_1077,In_381,In_498);
and U1078 (N_1078,In_230,In_461);
and U1079 (N_1079,In_56,In_25);
nand U1080 (N_1080,In_197,In_168);
nor U1081 (N_1081,In_661,In_639);
and U1082 (N_1082,In_249,In_652);
nand U1083 (N_1083,In_73,In_848);
nor U1084 (N_1084,In_850,In_574);
nand U1085 (N_1085,In_125,In_865);
nand U1086 (N_1086,In_650,In_300);
or U1087 (N_1087,In_436,In_619);
nand U1088 (N_1088,In_123,In_144);
nand U1089 (N_1089,In_243,In_839);
and U1090 (N_1090,In_631,In_505);
and U1091 (N_1091,In_531,In_243);
or U1092 (N_1092,In_969,In_880);
and U1093 (N_1093,In_300,In_29);
nor U1094 (N_1094,In_84,In_911);
nand U1095 (N_1095,In_794,In_716);
and U1096 (N_1096,In_925,In_201);
or U1097 (N_1097,In_213,In_970);
nor U1098 (N_1098,In_96,In_387);
nand U1099 (N_1099,In_38,In_161);
nor U1100 (N_1100,In_234,In_151);
nand U1101 (N_1101,In_21,In_484);
or U1102 (N_1102,In_564,In_417);
or U1103 (N_1103,In_411,In_187);
nand U1104 (N_1104,In_274,In_731);
and U1105 (N_1105,In_853,In_548);
nand U1106 (N_1106,In_177,In_743);
nand U1107 (N_1107,In_671,In_302);
nor U1108 (N_1108,In_994,In_633);
nor U1109 (N_1109,In_46,In_231);
nand U1110 (N_1110,In_911,In_594);
nor U1111 (N_1111,In_61,In_809);
or U1112 (N_1112,In_217,In_420);
nand U1113 (N_1113,In_232,In_359);
nand U1114 (N_1114,In_57,In_530);
nor U1115 (N_1115,In_932,In_62);
nor U1116 (N_1116,In_354,In_740);
or U1117 (N_1117,In_347,In_623);
or U1118 (N_1118,In_439,In_349);
nand U1119 (N_1119,In_796,In_891);
and U1120 (N_1120,In_844,In_447);
nor U1121 (N_1121,In_502,In_396);
and U1122 (N_1122,In_361,In_67);
or U1123 (N_1123,In_285,In_287);
nor U1124 (N_1124,In_998,In_780);
or U1125 (N_1125,In_111,In_515);
or U1126 (N_1126,In_684,In_897);
or U1127 (N_1127,In_139,In_717);
and U1128 (N_1128,In_51,In_343);
and U1129 (N_1129,In_477,In_270);
nor U1130 (N_1130,In_624,In_945);
nand U1131 (N_1131,In_743,In_92);
nor U1132 (N_1132,In_559,In_533);
nand U1133 (N_1133,In_950,In_295);
and U1134 (N_1134,In_445,In_132);
or U1135 (N_1135,In_439,In_11);
or U1136 (N_1136,In_927,In_197);
nand U1137 (N_1137,In_825,In_18);
nor U1138 (N_1138,In_852,In_799);
or U1139 (N_1139,In_282,In_163);
nand U1140 (N_1140,In_271,In_149);
or U1141 (N_1141,In_272,In_85);
nor U1142 (N_1142,In_478,In_640);
nor U1143 (N_1143,In_774,In_255);
and U1144 (N_1144,In_868,In_563);
or U1145 (N_1145,In_59,In_411);
nor U1146 (N_1146,In_355,In_745);
and U1147 (N_1147,In_395,In_513);
nand U1148 (N_1148,In_503,In_293);
and U1149 (N_1149,In_82,In_647);
nand U1150 (N_1150,In_902,In_338);
nor U1151 (N_1151,In_88,In_803);
and U1152 (N_1152,In_879,In_367);
nor U1153 (N_1153,In_793,In_343);
nand U1154 (N_1154,In_277,In_983);
nor U1155 (N_1155,In_71,In_153);
nand U1156 (N_1156,In_44,In_995);
nor U1157 (N_1157,In_910,In_132);
nor U1158 (N_1158,In_797,In_599);
nand U1159 (N_1159,In_966,In_877);
nand U1160 (N_1160,In_688,In_949);
and U1161 (N_1161,In_610,In_152);
and U1162 (N_1162,In_629,In_217);
nand U1163 (N_1163,In_820,In_624);
nor U1164 (N_1164,In_513,In_30);
nand U1165 (N_1165,In_534,In_345);
and U1166 (N_1166,In_458,In_547);
nor U1167 (N_1167,In_674,In_336);
and U1168 (N_1168,In_550,In_851);
nor U1169 (N_1169,In_451,In_333);
or U1170 (N_1170,In_285,In_345);
nand U1171 (N_1171,In_539,In_982);
nor U1172 (N_1172,In_703,In_14);
nand U1173 (N_1173,In_866,In_836);
nor U1174 (N_1174,In_121,In_690);
and U1175 (N_1175,In_247,In_156);
nand U1176 (N_1176,In_809,In_980);
nand U1177 (N_1177,In_608,In_859);
nor U1178 (N_1178,In_692,In_921);
nor U1179 (N_1179,In_280,In_340);
and U1180 (N_1180,In_60,In_26);
nand U1181 (N_1181,In_939,In_134);
or U1182 (N_1182,In_876,In_795);
nand U1183 (N_1183,In_401,In_233);
nor U1184 (N_1184,In_333,In_317);
nor U1185 (N_1185,In_22,In_174);
and U1186 (N_1186,In_11,In_685);
nand U1187 (N_1187,In_126,In_211);
and U1188 (N_1188,In_523,In_137);
nor U1189 (N_1189,In_232,In_33);
nor U1190 (N_1190,In_967,In_537);
nand U1191 (N_1191,In_250,In_734);
and U1192 (N_1192,In_612,In_966);
or U1193 (N_1193,In_136,In_710);
and U1194 (N_1194,In_958,In_610);
or U1195 (N_1195,In_939,In_204);
nand U1196 (N_1196,In_237,In_453);
nor U1197 (N_1197,In_439,In_7);
or U1198 (N_1198,In_283,In_396);
or U1199 (N_1199,In_734,In_131);
or U1200 (N_1200,In_906,In_572);
nand U1201 (N_1201,In_416,In_442);
and U1202 (N_1202,In_258,In_883);
nand U1203 (N_1203,In_920,In_909);
or U1204 (N_1204,In_264,In_21);
and U1205 (N_1205,In_641,In_922);
or U1206 (N_1206,In_566,In_275);
or U1207 (N_1207,In_16,In_234);
or U1208 (N_1208,In_948,In_42);
or U1209 (N_1209,In_663,In_16);
and U1210 (N_1210,In_346,In_79);
nor U1211 (N_1211,In_342,In_709);
or U1212 (N_1212,In_387,In_366);
nand U1213 (N_1213,In_127,In_983);
nand U1214 (N_1214,In_552,In_407);
or U1215 (N_1215,In_480,In_194);
nand U1216 (N_1216,In_138,In_614);
or U1217 (N_1217,In_981,In_629);
or U1218 (N_1218,In_951,In_14);
nor U1219 (N_1219,In_720,In_898);
or U1220 (N_1220,In_651,In_210);
and U1221 (N_1221,In_989,In_624);
nand U1222 (N_1222,In_511,In_886);
nor U1223 (N_1223,In_448,In_776);
and U1224 (N_1224,In_204,In_656);
or U1225 (N_1225,In_738,In_970);
and U1226 (N_1226,In_842,In_545);
or U1227 (N_1227,In_735,In_343);
nor U1228 (N_1228,In_690,In_287);
nand U1229 (N_1229,In_782,In_342);
and U1230 (N_1230,In_77,In_800);
and U1231 (N_1231,In_208,In_845);
and U1232 (N_1232,In_666,In_493);
and U1233 (N_1233,In_747,In_953);
and U1234 (N_1234,In_981,In_592);
nand U1235 (N_1235,In_755,In_61);
and U1236 (N_1236,In_872,In_540);
and U1237 (N_1237,In_1,In_673);
or U1238 (N_1238,In_527,In_312);
nand U1239 (N_1239,In_891,In_327);
and U1240 (N_1240,In_998,In_235);
and U1241 (N_1241,In_783,In_612);
nor U1242 (N_1242,In_422,In_637);
nand U1243 (N_1243,In_802,In_547);
or U1244 (N_1244,In_269,In_722);
or U1245 (N_1245,In_798,In_466);
or U1246 (N_1246,In_757,In_132);
nand U1247 (N_1247,In_859,In_403);
nand U1248 (N_1248,In_419,In_108);
or U1249 (N_1249,In_709,In_16);
or U1250 (N_1250,In_312,In_592);
and U1251 (N_1251,In_66,In_77);
xor U1252 (N_1252,In_17,In_510);
nor U1253 (N_1253,In_216,In_903);
and U1254 (N_1254,In_980,In_353);
or U1255 (N_1255,In_220,In_243);
or U1256 (N_1256,In_197,In_558);
and U1257 (N_1257,In_492,In_258);
nor U1258 (N_1258,In_960,In_206);
and U1259 (N_1259,In_271,In_51);
nand U1260 (N_1260,In_196,In_853);
and U1261 (N_1261,In_593,In_169);
and U1262 (N_1262,In_673,In_802);
or U1263 (N_1263,In_915,In_879);
or U1264 (N_1264,In_468,In_845);
or U1265 (N_1265,In_952,In_797);
nand U1266 (N_1266,In_337,In_760);
nand U1267 (N_1267,In_931,In_551);
nor U1268 (N_1268,In_581,In_66);
nor U1269 (N_1269,In_60,In_935);
nand U1270 (N_1270,In_459,In_954);
or U1271 (N_1271,In_102,In_192);
and U1272 (N_1272,In_618,In_391);
or U1273 (N_1273,In_947,In_401);
nand U1274 (N_1274,In_94,In_851);
and U1275 (N_1275,In_488,In_452);
or U1276 (N_1276,In_892,In_408);
xnor U1277 (N_1277,In_989,In_508);
nand U1278 (N_1278,In_631,In_480);
nor U1279 (N_1279,In_953,In_993);
or U1280 (N_1280,In_559,In_448);
and U1281 (N_1281,In_516,In_981);
and U1282 (N_1282,In_284,In_507);
and U1283 (N_1283,In_195,In_606);
nor U1284 (N_1284,In_70,In_635);
and U1285 (N_1285,In_70,In_725);
and U1286 (N_1286,In_956,In_360);
nand U1287 (N_1287,In_614,In_593);
and U1288 (N_1288,In_258,In_971);
nor U1289 (N_1289,In_617,In_220);
and U1290 (N_1290,In_704,In_591);
or U1291 (N_1291,In_897,In_935);
or U1292 (N_1292,In_655,In_626);
nand U1293 (N_1293,In_456,In_430);
or U1294 (N_1294,In_93,In_465);
or U1295 (N_1295,In_89,In_321);
or U1296 (N_1296,In_400,In_153);
or U1297 (N_1297,In_479,In_620);
or U1298 (N_1298,In_607,In_198);
or U1299 (N_1299,In_504,In_622);
nand U1300 (N_1300,In_49,In_446);
and U1301 (N_1301,In_899,In_149);
nor U1302 (N_1302,In_692,In_972);
nand U1303 (N_1303,In_968,In_332);
or U1304 (N_1304,In_830,In_983);
or U1305 (N_1305,In_709,In_200);
xnor U1306 (N_1306,In_275,In_106);
or U1307 (N_1307,In_217,In_945);
and U1308 (N_1308,In_344,In_135);
nand U1309 (N_1309,In_186,In_708);
or U1310 (N_1310,In_195,In_584);
nor U1311 (N_1311,In_597,In_828);
nand U1312 (N_1312,In_748,In_142);
or U1313 (N_1313,In_399,In_426);
and U1314 (N_1314,In_124,In_468);
nand U1315 (N_1315,In_36,In_644);
and U1316 (N_1316,In_310,In_709);
nor U1317 (N_1317,In_454,In_815);
nor U1318 (N_1318,In_424,In_676);
and U1319 (N_1319,In_654,In_8);
or U1320 (N_1320,In_512,In_827);
or U1321 (N_1321,In_122,In_890);
or U1322 (N_1322,In_204,In_263);
or U1323 (N_1323,In_794,In_303);
nor U1324 (N_1324,In_19,In_289);
or U1325 (N_1325,In_166,In_137);
nor U1326 (N_1326,In_761,In_528);
and U1327 (N_1327,In_22,In_561);
nand U1328 (N_1328,In_875,In_69);
nor U1329 (N_1329,In_126,In_975);
and U1330 (N_1330,In_182,In_953);
nand U1331 (N_1331,In_687,In_16);
nand U1332 (N_1332,In_323,In_276);
or U1333 (N_1333,In_64,In_67);
nor U1334 (N_1334,In_636,In_612);
or U1335 (N_1335,In_690,In_604);
nor U1336 (N_1336,In_501,In_136);
nand U1337 (N_1337,In_9,In_306);
nand U1338 (N_1338,In_235,In_631);
and U1339 (N_1339,In_849,In_683);
and U1340 (N_1340,In_442,In_675);
and U1341 (N_1341,In_162,In_135);
or U1342 (N_1342,In_601,In_399);
nand U1343 (N_1343,In_484,In_606);
nand U1344 (N_1344,In_714,In_449);
and U1345 (N_1345,In_275,In_713);
nand U1346 (N_1346,In_741,In_958);
or U1347 (N_1347,In_992,In_73);
nor U1348 (N_1348,In_125,In_785);
nand U1349 (N_1349,In_942,In_902);
nand U1350 (N_1350,In_687,In_974);
or U1351 (N_1351,In_143,In_91);
nand U1352 (N_1352,In_722,In_256);
or U1353 (N_1353,In_841,In_878);
nor U1354 (N_1354,In_622,In_386);
nand U1355 (N_1355,In_261,In_0);
and U1356 (N_1356,In_100,In_788);
nand U1357 (N_1357,In_535,In_169);
nand U1358 (N_1358,In_908,In_785);
and U1359 (N_1359,In_520,In_114);
nand U1360 (N_1360,In_588,In_864);
nand U1361 (N_1361,In_106,In_758);
and U1362 (N_1362,In_267,In_209);
or U1363 (N_1363,In_457,In_566);
xnor U1364 (N_1364,In_25,In_427);
or U1365 (N_1365,In_169,In_948);
nor U1366 (N_1366,In_870,In_981);
xnor U1367 (N_1367,In_190,In_684);
nor U1368 (N_1368,In_164,In_286);
and U1369 (N_1369,In_160,In_203);
or U1370 (N_1370,In_991,In_59);
or U1371 (N_1371,In_28,In_628);
and U1372 (N_1372,In_882,In_655);
nor U1373 (N_1373,In_154,In_274);
nand U1374 (N_1374,In_623,In_555);
or U1375 (N_1375,In_562,In_218);
nor U1376 (N_1376,In_891,In_902);
and U1377 (N_1377,In_993,In_666);
and U1378 (N_1378,In_424,In_697);
or U1379 (N_1379,In_632,In_808);
nor U1380 (N_1380,In_491,In_679);
nor U1381 (N_1381,In_242,In_288);
nor U1382 (N_1382,In_285,In_864);
nand U1383 (N_1383,In_390,In_796);
or U1384 (N_1384,In_806,In_345);
or U1385 (N_1385,In_526,In_301);
and U1386 (N_1386,In_939,In_354);
and U1387 (N_1387,In_838,In_526);
nor U1388 (N_1388,In_747,In_695);
or U1389 (N_1389,In_52,In_82);
nand U1390 (N_1390,In_818,In_736);
or U1391 (N_1391,In_585,In_540);
nand U1392 (N_1392,In_355,In_645);
and U1393 (N_1393,In_395,In_598);
nand U1394 (N_1394,In_71,In_773);
or U1395 (N_1395,In_455,In_278);
nor U1396 (N_1396,In_932,In_53);
nand U1397 (N_1397,In_910,In_795);
nand U1398 (N_1398,In_177,In_204);
or U1399 (N_1399,In_660,In_424);
nand U1400 (N_1400,In_700,In_508);
nor U1401 (N_1401,In_944,In_356);
nand U1402 (N_1402,In_809,In_358);
and U1403 (N_1403,In_485,In_612);
and U1404 (N_1404,In_455,In_130);
and U1405 (N_1405,In_911,In_905);
nand U1406 (N_1406,In_979,In_104);
nor U1407 (N_1407,In_20,In_938);
nand U1408 (N_1408,In_710,In_517);
nand U1409 (N_1409,In_387,In_825);
and U1410 (N_1410,In_433,In_904);
nand U1411 (N_1411,In_608,In_861);
or U1412 (N_1412,In_550,In_772);
nor U1413 (N_1413,In_272,In_398);
or U1414 (N_1414,In_207,In_475);
or U1415 (N_1415,In_843,In_527);
nor U1416 (N_1416,In_30,In_111);
or U1417 (N_1417,In_360,In_528);
nand U1418 (N_1418,In_280,In_777);
nand U1419 (N_1419,In_179,In_396);
or U1420 (N_1420,In_631,In_321);
nor U1421 (N_1421,In_449,In_797);
nor U1422 (N_1422,In_371,In_624);
nand U1423 (N_1423,In_58,In_705);
nor U1424 (N_1424,In_225,In_237);
nand U1425 (N_1425,In_375,In_931);
nor U1426 (N_1426,In_28,In_272);
nand U1427 (N_1427,In_575,In_363);
and U1428 (N_1428,In_254,In_982);
nor U1429 (N_1429,In_284,In_435);
xor U1430 (N_1430,In_616,In_458);
and U1431 (N_1431,In_860,In_976);
and U1432 (N_1432,In_689,In_808);
nor U1433 (N_1433,In_37,In_474);
or U1434 (N_1434,In_684,In_636);
nand U1435 (N_1435,In_647,In_843);
nand U1436 (N_1436,In_458,In_636);
nand U1437 (N_1437,In_909,In_793);
nand U1438 (N_1438,In_601,In_813);
nor U1439 (N_1439,In_430,In_592);
and U1440 (N_1440,In_382,In_438);
nand U1441 (N_1441,In_397,In_254);
nor U1442 (N_1442,In_728,In_69);
and U1443 (N_1443,In_564,In_701);
and U1444 (N_1444,In_130,In_566);
or U1445 (N_1445,In_391,In_339);
or U1446 (N_1446,In_258,In_575);
nand U1447 (N_1447,In_142,In_331);
and U1448 (N_1448,In_130,In_51);
or U1449 (N_1449,In_704,In_997);
nand U1450 (N_1450,In_446,In_373);
nor U1451 (N_1451,In_183,In_767);
nand U1452 (N_1452,In_23,In_108);
nand U1453 (N_1453,In_667,In_464);
nand U1454 (N_1454,In_507,In_787);
or U1455 (N_1455,In_599,In_712);
nand U1456 (N_1456,In_996,In_446);
or U1457 (N_1457,In_940,In_554);
nor U1458 (N_1458,In_400,In_146);
nor U1459 (N_1459,In_925,In_345);
nor U1460 (N_1460,In_507,In_627);
and U1461 (N_1461,In_909,In_752);
nor U1462 (N_1462,In_456,In_645);
nand U1463 (N_1463,In_516,In_176);
nand U1464 (N_1464,In_101,In_649);
nor U1465 (N_1465,In_475,In_874);
and U1466 (N_1466,In_213,In_358);
or U1467 (N_1467,In_729,In_440);
nand U1468 (N_1468,In_154,In_857);
and U1469 (N_1469,In_623,In_228);
nand U1470 (N_1470,In_410,In_705);
and U1471 (N_1471,In_747,In_952);
and U1472 (N_1472,In_378,In_178);
or U1473 (N_1473,In_805,In_811);
or U1474 (N_1474,In_872,In_83);
nor U1475 (N_1475,In_222,In_525);
and U1476 (N_1476,In_191,In_396);
and U1477 (N_1477,In_846,In_182);
and U1478 (N_1478,In_904,In_261);
and U1479 (N_1479,In_605,In_335);
or U1480 (N_1480,In_962,In_986);
or U1481 (N_1481,In_259,In_814);
or U1482 (N_1482,In_678,In_178);
nand U1483 (N_1483,In_778,In_943);
nand U1484 (N_1484,In_99,In_910);
or U1485 (N_1485,In_33,In_350);
nand U1486 (N_1486,In_42,In_382);
or U1487 (N_1487,In_667,In_641);
nand U1488 (N_1488,In_48,In_197);
and U1489 (N_1489,In_446,In_155);
or U1490 (N_1490,In_797,In_842);
or U1491 (N_1491,In_314,In_909);
nor U1492 (N_1492,In_680,In_80);
and U1493 (N_1493,In_3,In_389);
nor U1494 (N_1494,In_217,In_989);
nor U1495 (N_1495,In_577,In_192);
or U1496 (N_1496,In_887,In_685);
and U1497 (N_1497,In_975,In_582);
or U1498 (N_1498,In_9,In_351);
nand U1499 (N_1499,In_617,In_521);
nor U1500 (N_1500,In_606,In_971);
nor U1501 (N_1501,In_823,In_979);
or U1502 (N_1502,In_869,In_530);
and U1503 (N_1503,In_116,In_650);
or U1504 (N_1504,In_861,In_635);
or U1505 (N_1505,In_799,In_420);
nor U1506 (N_1506,In_187,In_899);
or U1507 (N_1507,In_979,In_599);
and U1508 (N_1508,In_355,In_31);
or U1509 (N_1509,In_466,In_703);
nand U1510 (N_1510,In_818,In_475);
and U1511 (N_1511,In_670,In_437);
nand U1512 (N_1512,In_501,In_693);
and U1513 (N_1513,In_864,In_145);
and U1514 (N_1514,In_951,In_83);
and U1515 (N_1515,In_911,In_212);
or U1516 (N_1516,In_726,In_522);
or U1517 (N_1517,In_313,In_666);
or U1518 (N_1518,In_1,In_371);
nand U1519 (N_1519,In_995,In_840);
and U1520 (N_1520,In_476,In_239);
and U1521 (N_1521,In_269,In_63);
or U1522 (N_1522,In_330,In_824);
nor U1523 (N_1523,In_578,In_889);
nand U1524 (N_1524,In_599,In_318);
or U1525 (N_1525,In_769,In_674);
nor U1526 (N_1526,In_425,In_0);
nor U1527 (N_1527,In_448,In_222);
or U1528 (N_1528,In_230,In_41);
nand U1529 (N_1529,In_284,In_106);
and U1530 (N_1530,In_965,In_688);
nor U1531 (N_1531,In_123,In_971);
and U1532 (N_1532,In_388,In_151);
or U1533 (N_1533,In_852,In_87);
and U1534 (N_1534,In_362,In_907);
and U1535 (N_1535,In_82,In_861);
nand U1536 (N_1536,In_713,In_434);
and U1537 (N_1537,In_695,In_690);
or U1538 (N_1538,In_865,In_861);
nor U1539 (N_1539,In_594,In_468);
nand U1540 (N_1540,In_710,In_66);
nand U1541 (N_1541,In_139,In_796);
nor U1542 (N_1542,In_677,In_859);
nand U1543 (N_1543,In_880,In_74);
and U1544 (N_1544,In_151,In_11);
nand U1545 (N_1545,In_568,In_909);
and U1546 (N_1546,In_985,In_815);
or U1547 (N_1547,In_858,In_815);
xor U1548 (N_1548,In_543,In_733);
or U1549 (N_1549,In_264,In_994);
nor U1550 (N_1550,In_130,In_390);
nor U1551 (N_1551,In_701,In_688);
or U1552 (N_1552,In_465,In_991);
nand U1553 (N_1553,In_785,In_373);
and U1554 (N_1554,In_804,In_312);
and U1555 (N_1555,In_613,In_81);
or U1556 (N_1556,In_806,In_909);
and U1557 (N_1557,In_570,In_627);
and U1558 (N_1558,In_900,In_842);
nand U1559 (N_1559,In_803,In_431);
and U1560 (N_1560,In_59,In_191);
nor U1561 (N_1561,In_828,In_399);
and U1562 (N_1562,In_332,In_788);
nand U1563 (N_1563,In_456,In_618);
and U1564 (N_1564,In_110,In_376);
and U1565 (N_1565,In_681,In_315);
nor U1566 (N_1566,In_303,In_246);
nor U1567 (N_1567,In_193,In_387);
nand U1568 (N_1568,In_961,In_470);
nor U1569 (N_1569,In_490,In_71);
nand U1570 (N_1570,In_528,In_1);
or U1571 (N_1571,In_59,In_903);
and U1572 (N_1572,In_23,In_877);
nand U1573 (N_1573,In_837,In_13);
nor U1574 (N_1574,In_114,In_125);
and U1575 (N_1575,In_116,In_191);
or U1576 (N_1576,In_817,In_582);
nor U1577 (N_1577,In_717,In_578);
nor U1578 (N_1578,In_603,In_107);
nand U1579 (N_1579,In_42,In_274);
or U1580 (N_1580,In_412,In_99);
and U1581 (N_1581,In_15,In_141);
and U1582 (N_1582,In_755,In_324);
nor U1583 (N_1583,In_865,In_296);
nand U1584 (N_1584,In_159,In_521);
or U1585 (N_1585,In_204,In_382);
and U1586 (N_1586,In_262,In_137);
nor U1587 (N_1587,In_539,In_197);
nor U1588 (N_1588,In_499,In_408);
and U1589 (N_1589,In_612,In_188);
or U1590 (N_1590,In_384,In_651);
nor U1591 (N_1591,In_197,In_647);
or U1592 (N_1592,In_328,In_798);
nor U1593 (N_1593,In_759,In_354);
or U1594 (N_1594,In_444,In_827);
and U1595 (N_1595,In_788,In_437);
and U1596 (N_1596,In_868,In_283);
and U1597 (N_1597,In_453,In_437);
nor U1598 (N_1598,In_841,In_209);
or U1599 (N_1599,In_711,In_750);
or U1600 (N_1600,In_512,In_793);
nand U1601 (N_1601,In_983,In_398);
nor U1602 (N_1602,In_23,In_838);
or U1603 (N_1603,In_835,In_713);
and U1604 (N_1604,In_442,In_528);
nand U1605 (N_1605,In_508,In_607);
nand U1606 (N_1606,In_680,In_538);
and U1607 (N_1607,In_915,In_197);
and U1608 (N_1608,In_26,In_493);
nand U1609 (N_1609,In_947,In_344);
nand U1610 (N_1610,In_675,In_302);
and U1611 (N_1611,In_405,In_658);
nand U1612 (N_1612,In_3,In_386);
and U1613 (N_1613,In_152,In_745);
nand U1614 (N_1614,In_505,In_507);
nor U1615 (N_1615,In_131,In_713);
nor U1616 (N_1616,In_871,In_620);
nor U1617 (N_1617,In_674,In_478);
nand U1618 (N_1618,In_492,In_662);
nand U1619 (N_1619,In_685,In_568);
nand U1620 (N_1620,In_522,In_988);
nor U1621 (N_1621,In_554,In_208);
nor U1622 (N_1622,In_934,In_967);
nand U1623 (N_1623,In_53,In_73);
or U1624 (N_1624,In_428,In_624);
or U1625 (N_1625,In_19,In_627);
or U1626 (N_1626,In_800,In_960);
nor U1627 (N_1627,In_693,In_15);
nor U1628 (N_1628,In_60,In_437);
xnor U1629 (N_1629,In_849,In_847);
and U1630 (N_1630,In_933,In_696);
or U1631 (N_1631,In_730,In_723);
or U1632 (N_1632,In_145,In_659);
or U1633 (N_1633,In_848,In_922);
and U1634 (N_1634,In_997,In_638);
nor U1635 (N_1635,In_578,In_220);
nor U1636 (N_1636,In_685,In_622);
and U1637 (N_1637,In_422,In_901);
nand U1638 (N_1638,In_652,In_559);
nor U1639 (N_1639,In_211,In_578);
nand U1640 (N_1640,In_294,In_685);
or U1641 (N_1641,In_632,In_830);
nand U1642 (N_1642,In_668,In_681);
and U1643 (N_1643,In_585,In_997);
nand U1644 (N_1644,In_515,In_433);
nor U1645 (N_1645,In_250,In_813);
or U1646 (N_1646,In_712,In_682);
nor U1647 (N_1647,In_891,In_286);
and U1648 (N_1648,In_270,In_106);
nand U1649 (N_1649,In_103,In_727);
nor U1650 (N_1650,In_722,In_830);
and U1651 (N_1651,In_530,In_492);
and U1652 (N_1652,In_590,In_597);
or U1653 (N_1653,In_869,In_874);
nand U1654 (N_1654,In_554,In_892);
nor U1655 (N_1655,In_804,In_473);
nor U1656 (N_1656,In_883,In_385);
and U1657 (N_1657,In_701,In_521);
or U1658 (N_1658,In_13,In_209);
or U1659 (N_1659,In_621,In_222);
nand U1660 (N_1660,In_275,In_828);
or U1661 (N_1661,In_740,In_996);
and U1662 (N_1662,In_583,In_128);
nor U1663 (N_1663,In_937,In_651);
or U1664 (N_1664,In_588,In_461);
nor U1665 (N_1665,In_887,In_647);
or U1666 (N_1666,In_601,In_468);
and U1667 (N_1667,In_59,In_415);
and U1668 (N_1668,In_824,In_257);
nor U1669 (N_1669,In_330,In_508);
nor U1670 (N_1670,In_651,In_792);
nor U1671 (N_1671,In_31,In_688);
or U1672 (N_1672,In_61,In_138);
nand U1673 (N_1673,In_506,In_521);
or U1674 (N_1674,In_41,In_529);
nor U1675 (N_1675,In_567,In_279);
nand U1676 (N_1676,In_291,In_501);
and U1677 (N_1677,In_141,In_801);
or U1678 (N_1678,In_859,In_948);
or U1679 (N_1679,In_571,In_790);
nand U1680 (N_1680,In_719,In_310);
nand U1681 (N_1681,In_114,In_259);
and U1682 (N_1682,In_214,In_799);
and U1683 (N_1683,In_265,In_383);
nand U1684 (N_1684,In_610,In_521);
nor U1685 (N_1685,In_665,In_701);
or U1686 (N_1686,In_540,In_916);
nand U1687 (N_1687,In_128,In_487);
and U1688 (N_1688,In_480,In_125);
nor U1689 (N_1689,In_199,In_283);
nand U1690 (N_1690,In_218,In_89);
nor U1691 (N_1691,In_167,In_189);
nor U1692 (N_1692,In_823,In_481);
nand U1693 (N_1693,In_517,In_748);
and U1694 (N_1694,In_539,In_402);
nor U1695 (N_1695,In_66,In_845);
xor U1696 (N_1696,In_632,In_601);
or U1697 (N_1697,In_712,In_106);
nor U1698 (N_1698,In_158,In_15);
nand U1699 (N_1699,In_665,In_20);
nor U1700 (N_1700,In_47,In_258);
or U1701 (N_1701,In_633,In_426);
xor U1702 (N_1702,In_105,In_882);
nor U1703 (N_1703,In_49,In_53);
or U1704 (N_1704,In_743,In_573);
and U1705 (N_1705,In_565,In_825);
nand U1706 (N_1706,In_720,In_67);
nand U1707 (N_1707,In_463,In_330);
and U1708 (N_1708,In_766,In_224);
nand U1709 (N_1709,In_170,In_350);
nor U1710 (N_1710,In_985,In_217);
or U1711 (N_1711,In_942,In_17);
nor U1712 (N_1712,In_28,In_318);
and U1713 (N_1713,In_414,In_728);
or U1714 (N_1714,In_77,In_386);
nor U1715 (N_1715,In_718,In_95);
and U1716 (N_1716,In_863,In_313);
nand U1717 (N_1717,In_526,In_551);
or U1718 (N_1718,In_761,In_880);
nor U1719 (N_1719,In_881,In_991);
nor U1720 (N_1720,In_792,In_731);
xor U1721 (N_1721,In_982,In_172);
or U1722 (N_1722,In_881,In_924);
and U1723 (N_1723,In_850,In_24);
nor U1724 (N_1724,In_351,In_186);
or U1725 (N_1725,In_843,In_560);
or U1726 (N_1726,In_940,In_308);
nor U1727 (N_1727,In_476,In_848);
nand U1728 (N_1728,In_479,In_585);
nor U1729 (N_1729,In_468,In_863);
nand U1730 (N_1730,In_560,In_856);
nand U1731 (N_1731,In_126,In_448);
nand U1732 (N_1732,In_587,In_435);
and U1733 (N_1733,In_727,In_132);
nand U1734 (N_1734,In_177,In_888);
and U1735 (N_1735,In_85,In_286);
nand U1736 (N_1736,In_108,In_381);
and U1737 (N_1737,In_701,In_963);
nand U1738 (N_1738,In_775,In_456);
nor U1739 (N_1739,In_145,In_621);
and U1740 (N_1740,In_676,In_265);
or U1741 (N_1741,In_803,In_198);
or U1742 (N_1742,In_589,In_559);
nor U1743 (N_1743,In_932,In_598);
nand U1744 (N_1744,In_632,In_376);
and U1745 (N_1745,In_201,In_944);
nand U1746 (N_1746,In_201,In_359);
nor U1747 (N_1747,In_479,In_867);
nor U1748 (N_1748,In_605,In_732);
nor U1749 (N_1749,In_606,In_932);
and U1750 (N_1750,In_417,In_225);
nor U1751 (N_1751,In_856,In_768);
and U1752 (N_1752,In_470,In_824);
xnor U1753 (N_1753,In_756,In_19);
and U1754 (N_1754,In_156,In_526);
and U1755 (N_1755,In_624,In_602);
nand U1756 (N_1756,In_115,In_827);
and U1757 (N_1757,In_460,In_365);
nand U1758 (N_1758,In_939,In_750);
or U1759 (N_1759,In_308,In_966);
or U1760 (N_1760,In_471,In_864);
or U1761 (N_1761,In_737,In_825);
nor U1762 (N_1762,In_232,In_590);
or U1763 (N_1763,In_706,In_667);
and U1764 (N_1764,In_904,In_982);
and U1765 (N_1765,In_464,In_345);
nor U1766 (N_1766,In_537,In_272);
or U1767 (N_1767,In_441,In_324);
nand U1768 (N_1768,In_434,In_588);
or U1769 (N_1769,In_234,In_208);
nand U1770 (N_1770,In_653,In_702);
nand U1771 (N_1771,In_397,In_122);
or U1772 (N_1772,In_783,In_215);
and U1773 (N_1773,In_103,In_230);
or U1774 (N_1774,In_419,In_422);
nor U1775 (N_1775,In_700,In_642);
nor U1776 (N_1776,In_945,In_405);
and U1777 (N_1777,In_638,In_430);
and U1778 (N_1778,In_249,In_53);
and U1779 (N_1779,In_960,In_750);
or U1780 (N_1780,In_420,In_972);
or U1781 (N_1781,In_689,In_984);
nand U1782 (N_1782,In_94,In_287);
and U1783 (N_1783,In_787,In_321);
or U1784 (N_1784,In_497,In_804);
and U1785 (N_1785,In_114,In_323);
and U1786 (N_1786,In_898,In_558);
or U1787 (N_1787,In_647,In_403);
and U1788 (N_1788,In_96,In_904);
nand U1789 (N_1789,In_316,In_909);
and U1790 (N_1790,In_485,In_388);
or U1791 (N_1791,In_968,In_481);
or U1792 (N_1792,In_42,In_82);
nand U1793 (N_1793,In_894,In_787);
and U1794 (N_1794,In_472,In_451);
or U1795 (N_1795,In_294,In_282);
or U1796 (N_1796,In_207,In_172);
nor U1797 (N_1797,In_801,In_922);
nor U1798 (N_1798,In_885,In_756);
and U1799 (N_1799,In_252,In_115);
nor U1800 (N_1800,In_118,In_163);
or U1801 (N_1801,In_486,In_512);
nand U1802 (N_1802,In_422,In_16);
and U1803 (N_1803,In_410,In_769);
nor U1804 (N_1804,In_559,In_428);
and U1805 (N_1805,In_815,In_686);
nor U1806 (N_1806,In_429,In_906);
and U1807 (N_1807,In_445,In_188);
xnor U1808 (N_1808,In_345,In_682);
and U1809 (N_1809,In_559,In_491);
nand U1810 (N_1810,In_963,In_379);
nand U1811 (N_1811,In_864,In_846);
and U1812 (N_1812,In_921,In_981);
and U1813 (N_1813,In_715,In_551);
or U1814 (N_1814,In_140,In_967);
and U1815 (N_1815,In_921,In_330);
nor U1816 (N_1816,In_825,In_557);
nand U1817 (N_1817,In_729,In_748);
or U1818 (N_1818,In_339,In_454);
and U1819 (N_1819,In_28,In_402);
or U1820 (N_1820,In_755,In_757);
and U1821 (N_1821,In_484,In_764);
and U1822 (N_1822,In_448,In_987);
and U1823 (N_1823,In_969,In_356);
and U1824 (N_1824,In_998,In_220);
and U1825 (N_1825,In_389,In_927);
nand U1826 (N_1826,In_267,In_395);
nand U1827 (N_1827,In_585,In_296);
nand U1828 (N_1828,In_869,In_227);
and U1829 (N_1829,In_418,In_795);
or U1830 (N_1830,In_201,In_782);
nor U1831 (N_1831,In_591,In_679);
and U1832 (N_1832,In_938,In_862);
nor U1833 (N_1833,In_190,In_19);
nor U1834 (N_1834,In_343,In_9);
or U1835 (N_1835,In_461,In_245);
nor U1836 (N_1836,In_162,In_53);
or U1837 (N_1837,In_934,In_964);
and U1838 (N_1838,In_808,In_580);
or U1839 (N_1839,In_345,In_560);
nor U1840 (N_1840,In_399,In_424);
and U1841 (N_1841,In_312,In_10);
nor U1842 (N_1842,In_619,In_824);
nor U1843 (N_1843,In_956,In_378);
or U1844 (N_1844,In_587,In_693);
and U1845 (N_1845,In_137,In_40);
and U1846 (N_1846,In_420,In_763);
and U1847 (N_1847,In_94,In_517);
nand U1848 (N_1848,In_719,In_626);
or U1849 (N_1849,In_749,In_486);
nand U1850 (N_1850,In_839,In_698);
nor U1851 (N_1851,In_357,In_222);
nor U1852 (N_1852,In_884,In_640);
or U1853 (N_1853,In_391,In_458);
or U1854 (N_1854,In_287,In_408);
nand U1855 (N_1855,In_267,In_464);
xnor U1856 (N_1856,In_366,In_592);
nand U1857 (N_1857,In_614,In_758);
nand U1858 (N_1858,In_902,In_784);
xnor U1859 (N_1859,In_949,In_417);
or U1860 (N_1860,In_753,In_738);
or U1861 (N_1861,In_587,In_837);
or U1862 (N_1862,In_524,In_749);
nand U1863 (N_1863,In_723,In_154);
or U1864 (N_1864,In_174,In_566);
and U1865 (N_1865,In_364,In_634);
nor U1866 (N_1866,In_206,In_764);
or U1867 (N_1867,In_38,In_672);
nand U1868 (N_1868,In_76,In_480);
nor U1869 (N_1869,In_987,In_307);
or U1870 (N_1870,In_630,In_23);
nand U1871 (N_1871,In_67,In_595);
and U1872 (N_1872,In_51,In_26);
and U1873 (N_1873,In_106,In_983);
nand U1874 (N_1874,In_384,In_625);
or U1875 (N_1875,In_389,In_325);
nand U1876 (N_1876,In_818,In_459);
and U1877 (N_1877,In_901,In_652);
nand U1878 (N_1878,In_741,In_941);
nor U1879 (N_1879,In_743,In_227);
and U1880 (N_1880,In_243,In_705);
and U1881 (N_1881,In_710,In_217);
nor U1882 (N_1882,In_371,In_194);
nand U1883 (N_1883,In_540,In_366);
nor U1884 (N_1884,In_280,In_765);
nand U1885 (N_1885,In_931,In_808);
or U1886 (N_1886,In_204,In_536);
xor U1887 (N_1887,In_782,In_722);
nand U1888 (N_1888,In_315,In_699);
or U1889 (N_1889,In_539,In_757);
and U1890 (N_1890,In_112,In_517);
or U1891 (N_1891,In_878,In_644);
nor U1892 (N_1892,In_788,In_727);
or U1893 (N_1893,In_138,In_831);
and U1894 (N_1894,In_405,In_474);
nand U1895 (N_1895,In_963,In_177);
xnor U1896 (N_1896,In_913,In_575);
nand U1897 (N_1897,In_288,In_270);
nor U1898 (N_1898,In_4,In_285);
or U1899 (N_1899,In_19,In_177);
nor U1900 (N_1900,In_199,In_821);
nand U1901 (N_1901,In_454,In_694);
and U1902 (N_1902,In_78,In_511);
nor U1903 (N_1903,In_428,In_314);
nor U1904 (N_1904,In_900,In_463);
nand U1905 (N_1905,In_220,In_54);
nor U1906 (N_1906,In_499,In_616);
and U1907 (N_1907,In_471,In_263);
nand U1908 (N_1908,In_871,In_182);
and U1909 (N_1909,In_966,In_723);
nor U1910 (N_1910,In_134,In_490);
nor U1911 (N_1911,In_184,In_377);
and U1912 (N_1912,In_647,In_771);
and U1913 (N_1913,In_555,In_682);
or U1914 (N_1914,In_669,In_129);
nor U1915 (N_1915,In_747,In_659);
nor U1916 (N_1916,In_421,In_95);
nand U1917 (N_1917,In_732,In_470);
nand U1918 (N_1918,In_907,In_727);
and U1919 (N_1919,In_78,In_559);
nand U1920 (N_1920,In_419,In_567);
nand U1921 (N_1921,In_832,In_178);
and U1922 (N_1922,In_471,In_373);
or U1923 (N_1923,In_720,In_708);
or U1924 (N_1924,In_625,In_55);
nor U1925 (N_1925,In_203,In_173);
and U1926 (N_1926,In_790,In_171);
nand U1927 (N_1927,In_214,In_399);
nand U1928 (N_1928,In_56,In_665);
and U1929 (N_1929,In_527,In_206);
or U1930 (N_1930,In_234,In_754);
nand U1931 (N_1931,In_146,In_27);
and U1932 (N_1932,In_272,In_278);
nor U1933 (N_1933,In_599,In_265);
and U1934 (N_1934,In_461,In_562);
nor U1935 (N_1935,In_671,In_372);
or U1936 (N_1936,In_315,In_54);
nand U1937 (N_1937,In_36,In_792);
and U1938 (N_1938,In_247,In_91);
nand U1939 (N_1939,In_643,In_81);
nand U1940 (N_1940,In_175,In_837);
nor U1941 (N_1941,In_142,In_421);
nand U1942 (N_1942,In_365,In_899);
nor U1943 (N_1943,In_523,In_678);
nor U1944 (N_1944,In_29,In_330);
nand U1945 (N_1945,In_344,In_255);
or U1946 (N_1946,In_534,In_852);
and U1947 (N_1947,In_577,In_569);
or U1948 (N_1948,In_522,In_127);
and U1949 (N_1949,In_610,In_158);
nor U1950 (N_1950,In_329,In_676);
nor U1951 (N_1951,In_829,In_437);
or U1952 (N_1952,In_324,In_306);
nand U1953 (N_1953,In_383,In_796);
nor U1954 (N_1954,In_828,In_497);
or U1955 (N_1955,In_666,In_287);
or U1956 (N_1956,In_999,In_972);
xnor U1957 (N_1957,In_786,In_28);
nor U1958 (N_1958,In_649,In_812);
nand U1959 (N_1959,In_864,In_150);
nor U1960 (N_1960,In_865,In_251);
and U1961 (N_1961,In_474,In_973);
or U1962 (N_1962,In_697,In_194);
or U1963 (N_1963,In_958,In_533);
and U1964 (N_1964,In_400,In_832);
and U1965 (N_1965,In_161,In_697);
nand U1966 (N_1966,In_512,In_670);
and U1967 (N_1967,In_424,In_593);
xnor U1968 (N_1968,In_207,In_928);
nand U1969 (N_1969,In_184,In_421);
and U1970 (N_1970,In_549,In_429);
nand U1971 (N_1971,In_376,In_883);
xnor U1972 (N_1972,In_966,In_696);
and U1973 (N_1973,In_53,In_681);
nor U1974 (N_1974,In_478,In_579);
nand U1975 (N_1975,In_784,In_488);
or U1976 (N_1976,In_282,In_91);
and U1977 (N_1977,In_284,In_477);
or U1978 (N_1978,In_973,In_729);
nor U1979 (N_1979,In_897,In_760);
nor U1980 (N_1980,In_701,In_413);
and U1981 (N_1981,In_724,In_610);
nand U1982 (N_1982,In_156,In_251);
or U1983 (N_1983,In_246,In_201);
nand U1984 (N_1984,In_249,In_637);
nand U1985 (N_1985,In_600,In_830);
or U1986 (N_1986,In_179,In_923);
or U1987 (N_1987,In_254,In_178);
nand U1988 (N_1988,In_731,In_237);
and U1989 (N_1989,In_402,In_60);
nand U1990 (N_1990,In_380,In_564);
and U1991 (N_1991,In_500,In_343);
or U1992 (N_1992,In_298,In_341);
and U1993 (N_1993,In_597,In_880);
and U1994 (N_1994,In_365,In_437);
and U1995 (N_1995,In_624,In_130);
and U1996 (N_1996,In_807,In_416);
nand U1997 (N_1997,In_750,In_354);
or U1998 (N_1998,In_109,In_851);
or U1999 (N_1999,In_442,In_657);
and U2000 (N_2000,In_215,In_289);
and U2001 (N_2001,In_160,In_598);
nor U2002 (N_2002,In_678,In_232);
nor U2003 (N_2003,In_795,In_82);
nor U2004 (N_2004,In_446,In_178);
and U2005 (N_2005,In_121,In_672);
nand U2006 (N_2006,In_192,In_935);
nand U2007 (N_2007,In_830,In_719);
or U2008 (N_2008,In_569,In_796);
and U2009 (N_2009,In_654,In_478);
and U2010 (N_2010,In_529,In_308);
nor U2011 (N_2011,In_880,In_955);
nand U2012 (N_2012,In_481,In_100);
nand U2013 (N_2013,In_535,In_185);
nand U2014 (N_2014,In_474,In_11);
nor U2015 (N_2015,In_574,In_635);
nor U2016 (N_2016,In_882,In_496);
nor U2017 (N_2017,In_557,In_465);
or U2018 (N_2018,In_112,In_184);
nor U2019 (N_2019,In_705,In_469);
nor U2020 (N_2020,In_7,In_428);
or U2021 (N_2021,In_618,In_226);
or U2022 (N_2022,In_816,In_964);
nand U2023 (N_2023,In_190,In_912);
nand U2024 (N_2024,In_660,In_603);
or U2025 (N_2025,In_745,In_498);
and U2026 (N_2026,In_297,In_223);
nor U2027 (N_2027,In_674,In_220);
and U2028 (N_2028,In_358,In_539);
and U2029 (N_2029,In_175,In_554);
nor U2030 (N_2030,In_415,In_514);
or U2031 (N_2031,In_21,In_79);
and U2032 (N_2032,In_24,In_426);
and U2033 (N_2033,In_241,In_639);
nand U2034 (N_2034,In_676,In_323);
nor U2035 (N_2035,In_193,In_112);
and U2036 (N_2036,In_469,In_755);
or U2037 (N_2037,In_832,In_912);
nor U2038 (N_2038,In_917,In_960);
or U2039 (N_2039,In_945,In_802);
nand U2040 (N_2040,In_522,In_124);
or U2041 (N_2041,In_490,In_868);
and U2042 (N_2042,In_849,In_15);
or U2043 (N_2043,In_885,In_815);
nand U2044 (N_2044,In_283,In_471);
nand U2045 (N_2045,In_819,In_482);
and U2046 (N_2046,In_745,In_277);
or U2047 (N_2047,In_586,In_364);
nand U2048 (N_2048,In_299,In_275);
nor U2049 (N_2049,In_696,In_274);
nand U2050 (N_2050,In_48,In_973);
and U2051 (N_2051,In_374,In_38);
nor U2052 (N_2052,In_151,In_547);
nor U2053 (N_2053,In_473,In_765);
or U2054 (N_2054,In_418,In_82);
nand U2055 (N_2055,In_31,In_750);
nor U2056 (N_2056,In_289,In_663);
nor U2057 (N_2057,In_587,In_961);
nand U2058 (N_2058,In_96,In_187);
and U2059 (N_2059,In_24,In_461);
or U2060 (N_2060,In_170,In_606);
nor U2061 (N_2061,In_783,In_451);
nand U2062 (N_2062,In_244,In_308);
or U2063 (N_2063,In_259,In_257);
and U2064 (N_2064,In_513,In_93);
nor U2065 (N_2065,In_431,In_151);
nand U2066 (N_2066,In_944,In_731);
nand U2067 (N_2067,In_57,In_349);
nand U2068 (N_2068,In_998,In_666);
nor U2069 (N_2069,In_423,In_564);
and U2070 (N_2070,In_537,In_195);
or U2071 (N_2071,In_936,In_913);
nor U2072 (N_2072,In_792,In_256);
nand U2073 (N_2073,In_410,In_469);
nor U2074 (N_2074,In_923,In_459);
nand U2075 (N_2075,In_233,In_657);
nor U2076 (N_2076,In_22,In_156);
and U2077 (N_2077,In_276,In_669);
and U2078 (N_2078,In_240,In_675);
or U2079 (N_2079,In_578,In_105);
nand U2080 (N_2080,In_641,In_798);
or U2081 (N_2081,In_899,In_503);
and U2082 (N_2082,In_114,In_671);
or U2083 (N_2083,In_485,In_31);
nor U2084 (N_2084,In_735,In_42);
and U2085 (N_2085,In_415,In_360);
and U2086 (N_2086,In_676,In_830);
or U2087 (N_2087,In_817,In_76);
or U2088 (N_2088,In_391,In_207);
and U2089 (N_2089,In_618,In_208);
nand U2090 (N_2090,In_58,In_754);
and U2091 (N_2091,In_134,In_696);
and U2092 (N_2092,In_581,In_158);
nor U2093 (N_2093,In_764,In_183);
and U2094 (N_2094,In_337,In_305);
nor U2095 (N_2095,In_328,In_256);
nand U2096 (N_2096,In_35,In_937);
nand U2097 (N_2097,In_684,In_108);
and U2098 (N_2098,In_78,In_617);
nand U2099 (N_2099,In_543,In_7);
or U2100 (N_2100,In_688,In_919);
nand U2101 (N_2101,In_133,In_596);
nor U2102 (N_2102,In_145,In_344);
or U2103 (N_2103,In_255,In_467);
or U2104 (N_2104,In_682,In_582);
nand U2105 (N_2105,In_480,In_250);
and U2106 (N_2106,In_90,In_241);
and U2107 (N_2107,In_667,In_778);
or U2108 (N_2108,In_993,In_237);
nor U2109 (N_2109,In_985,In_286);
and U2110 (N_2110,In_172,In_376);
and U2111 (N_2111,In_737,In_395);
nand U2112 (N_2112,In_685,In_991);
and U2113 (N_2113,In_944,In_242);
and U2114 (N_2114,In_37,In_549);
nand U2115 (N_2115,In_650,In_202);
nand U2116 (N_2116,In_504,In_550);
or U2117 (N_2117,In_644,In_669);
nand U2118 (N_2118,In_306,In_185);
and U2119 (N_2119,In_591,In_649);
or U2120 (N_2120,In_112,In_194);
and U2121 (N_2121,In_37,In_925);
nand U2122 (N_2122,In_327,In_379);
and U2123 (N_2123,In_239,In_864);
nand U2124 (N_2124,In_668,In_436);
nand U2125 (N_2125,In_276,In_458);
or U2126 (N_2126,In_379,In_61);
and U2127 (N_2127,In_669,In_377);
or U2128 (N_2128,In_586,In_332);
and U2129 (N_2129,In_655,In_715);
and U2130 (N_2130,In_419,In_614);
nor U2131 (N_2131,In_179,In_566);
and U2132 (N_2132,In_265,In_441);
or U2133 (N_2133,In_345,In_869);
nand U2134 (N_2134,In_219,In_967);
or U2135 (N_2135,In_86,In_887);
nor U2136 (N_2136,In_714,In_709);
and U2137 (N_2137,In_749,In_504);
and U2138 (N_2138,In_949,In_775);
and U2139 (N_2139,In_375,In_84);
or U2140 (N_2140,In_556,In_743);
or U2141 (N_2141,In_593,In_242);
and U2142 (N_2142,In_340,In_483);
and U2143 (N_2143,In_347,In_863);
or U2144 (N_2144,In_476,In_482);
or U2145 (N_2145,In_417,In_384);
nand U2146 (N_2146,In_841,In_915);
and U2147 (N_2147,In_683,In_157);
nand U2148 (N_2148,In_547,In_475);
or U2149 (N_2149,In_518,In_48);
and U2150 (N_2150,In_338,In_670);
nor U2151 (N_2151,In_611,In_225);
nor U2152 (N_2152,In_363,In_853);
nor U2153 (N_2153,In_595,In_197);
and U2154 (N_2154,In_33,In_648);
and U2155 (N_2155,In_939,In_875);
or U2156 (N_2156,In_940,In_37);
or U2157 (N_2157,In_358,In_602);
and U2158 (N_2158,In_226,In_789);
or U2159 (N_2159,In_669,In_168);
nand U2160 (N_2160,In_156,In_283);
and U2161 (N_2161,In_922,In_719);
nor U2162 (N_2162,In_658,In_103);
or U2163 (N_2163,In_250,In_820);
nor U2164 (N_2164,In_753,In_445);
and U2165 (N_2165,In_217,In_714);
and U2166 (N_2166,In_621,In_326);
nor U2167 (N_2167,In_291,In_831);
or U2168 (N_2168,In_475,In_96);
nor U2169 (N_2169,In_938,In_64);
or U2170 (N_2170,In_221,In_660);
and U2171 (N_2171,In_129,In_735);
nand U2172 (N_2172,In_385,In_393);
nor U2173 (N_2173,In_455,In_885);
and U2174 (N_2174,In_987,In_166);
and U2175 (N_2175,In_54,In_40);
or U2176 (N_2176,In_423,In_179);
nor U2177 (N_2177,In_281,In_657);
nand U2178 (N_2178,In_577,In_395);
and U2179 (N_2179,In_715,In_29);
nand U2180 (N_2180,In_156,In_254);
nand U2181 (N_2181,In_868,In_895);
or U2182 (N_2182,In_260,In_795);
nand U2183 (N_2183,In_866,In_139);
and U2184 (N_2184,In_799,In_62);
and U2185 (N_2185,In_434,In_435);
nor U2186 (N_2186,In_351,In_747);
nor U2187 (N_2187,In_480,In_438);
nand U2188 (N_2188,In_916,In_873);
nor U2189 (N_2189,In_564,In_712);
nor U2190 (N_2190,In_101,In_194);
nor U2191 (N_2191,In_408,In_830);
nor U2192 (N_2192,In_217,In_489);
nor U2193 (N_2193,In_164,In_67);
and U2194 (N_2194,In_723,In_272);
and U2195 (N_2195,In_215,In_391);
or U2196 (N_2196,In_982,In_980);
and U2197 (N_2197,In_361,In_838);
or U2198 (N_2198,In_728,In_768);
nor U2199 (N_2199,In_443,In_936);
nand U2200 (N_2200,In_922,In_659);
nor U2201 (N_2201,In_365,In_918);
nand U2202 (N_2202,In_364,In_193);
nand U2203 (N_2203,In_765,In_230);
or U2204 (N_2204,In_978,In_803);
or U2205 (N_2205,In_519,In_505);
nand U2206 (N_2206,In_534,In_466);
nand U2207 (N_2207,In_724,In_699);
and U2208 (N_2208,In_551,In_914);
and U2209 (N_2209,In_930,In_557);
or U2210 (N_2210,In_754,In_331);
or U2211 (N_2211,In_607,In_677);
nand U2212 (N_2212,In_967,In_119);
and U2213 (N_2213,In_936,In_218);
nand U2214 (N_2214,In_963,In_267);
nand U2215 (N_2215,In_685,In_411);
nand U2216 (N_2216,In_42,In_986);
and U2217 (N_2217,In_641,In_986);
nor U2218 (N_2218,In_882,In_89);
and U2219 (N_2219,In_924,In_321);
nand U2220 (N_2220,In_238,In_894);
nand U2221 (N_2221,In_816,In_339);
nor U2222 (N_2222,In_270,In_611);
and U2223 (N_2223,In_382,In_364);
nand U2224 (N_2224,In_181,In_642);
or U2225 (N_2225,In_495,In_341);
nor U2226 (N_2226,In_303,In_963);
and U2227 (N_2227,In_509,In_959);
or U2228 (N_2228,In_19,In_142);
nand U2229 (N_2229,In_970,In_148);
and U2230 (N_2230,In_277,In_114);
nor U2231 (N_2231,In_29,In_912);
nand U2232 (N_2232,In_130,In_998);
nor U2233 (N_2233,In_840,In_760);
nor U2234 (N_2234,In_457,In_690);
and U2235 (N_2235,In_348,In_711);
nor U2236 (N_2236,In_49,In_400);
and U2237 (N_2237,In_683,In_300);
and U2238 (N_2238,In_551,In_407);
nor U2239 (N_2239,In_204,In_446);
nand U2240 (N_2240,In_485,In_970);
nand U2241 (N_2241,In_714,In_377);
nor U2242 (N_2242,In_84,In_962);
nand U2243 (N_2243,In_586,In_924);
nor U2244 (N_2244,In_65,In_33);
or U2245 (N_2245,In_659,In_71);
and U2246 (N_2246,In_46,In_860);
or U2247 (N_2247,In_990,In_364);
nand U2248 (N_2248,In_634,In_284);
or U2249 (N_2249,In_103,In_325);
nand U2250 (N_2250,In_967,In_638);
or U2251 (N_2251,In_276,In_697);
or U2252 (N_2252,In_839,In_559);
nand U2253 (N_2253,In_539,In_247);
nor U2254 (N_2254,In_164,In_387);
or U2255 (N_2255,In_671,In_286);
nand U2256 (N_2256,In_833,In_764);
nand U2257 (N_2257,In_241,In_362);
nand U2258 (N_2258,In_72,In_908);
nand U2259 (N_2259,In_332,In_358);
and U2260 (N_2260,In_645,In_259);
nand U2261 (N_2261,In_12,In_438);
nor U2262 (N_2262,In_394,In_522);
or U2263 (N_2263,In_920,In_664);
or U2264 (N_2264,In_658,In_41);
nand U2265 (N_2265,In_139,In_186);
xnor U2266 (N_2266,In_767,In_587);
or U2267 (N_2267,In_765,In_351);
or U2268 (N_2268,In_630,In_124);
or U2269 (N_2269,In_744,In_707);
and U2270 (N_2270,In_902,In_800);
nand U2271 (N_2271,In_197,In_345);
and U2272 (N_2272,In_882,In_673);
and U2273 (N_2273,In_524,In_369);
or U2274 (N_2274,In_276,In_299);
and U2275 (N_2275,In_178,In_471);
nand U2276 (N_2276,In_830,In_971);
nor U2277 (N_2277,In_920,In_814);
or U2278 (N_2278,In_701,In_837);
and U2279 (N_2279,In_882,In_34);
nand U2280 (N_2280,In_73,In_890);
nor U2281 (N_2281,In_149,In_717);
nor U2282 (N_2282,In_715,In_741);
nor U2283 (N_2283,In_683,In_212);
or U2284 (N_2284,In_992,In_190);
or U2285 (N_2285,In_641,In_512);
nor U2286 (N_2286,In_810,In_995);
and U2287 (N_2287,In_433,In_910);
or U2288 (N_2288,In_723,In_925);
or U2289 (N_2289,In_451,In_299);
and U2290 (N_2290,In_656,In_677);
or U2291 (N_2291,In_428,In_313);
or U2292 (N_2292,In_733,In_685);
and U2293 (N_2293,In_748,In_895);
and U2294 (N_2294,In_859,In_570);
nor U2295 (N_2295,In_847,In_843);
and U2296 (N_2296,In_237,In_575);
and U2297 (N_2297,In_111,In_411);
and U2298 (N_2298,In_953,In_453);
nand U2299 (N_2299,In_358,In_272);
or U2300 (N_2300,In_525,In_73);
nand U2301 (N_2301,In_718,In_499);
and U2302 (N_2302,In_199,In_238);
or U2303 (N_2303,In_439,In_989);
and U2304 (N_2304,In_17,In_836);
and U2305 (N_2305,In_772,In_663);
or U2306 (N_2306,In_987,In_500);
nand U2307 (N_2307,In_650,In_870);
and U2308 (N_2308,In_649,In_690);
and U2309 (N_2309,In_752,In_136);
nor U2310 (N_2310,In_722,In_19);
and U2311 (N_2311,In_225,In_836);
nand U2312 (N_2312,In_324,In_411);
nor U2313 (N_2313,In_398,In_497);
xnor U2314 (N_2314,In_372,In_766);
nand U2315 (N_2315,In_626,In_545);
nor U2316 (N_2316,In_28,In_537);
nor U2317 (N_2317,In_320,In_781);
and U2318 (N_2318,In_443,In_730);
nand U2319 (N_2319,In_128,In_384);
and U2320 (N_2320,In_695,In_637);
nor U2321 (N_2321,In_601,In_247);
or U2322 (N_2322,In_512,In_522);
and U2323 (N_2323,In_517,In_477);
nor U2324 (N_2324,In_61,In_883);
nand U2325 (N_2325,In_69,In_289);
nand U2326 (N_2326,In_189,In_846);
nand U2327 (N_2327,In_441,In_877);
nor U2328 (N_2328,In_338,In_67);
and U2329 (N_2329,In_805,In_552);
or U2330 (N_2330,In_735,In_354);
and U2331 (N_2331,In_242,In_537);
nor U2332 (N_2332,In_613,In_41);
and U2333 (N_2333,In_789,In_927);
nand U2334 (N_2334,In_609,In_87);
nand U2335 (N_2335,In_128,In_51);
nand U2336 (N_2336,In_654,In_222);
and U2337 (N_2337,In_635,In_62);
or U2338 (N_2338,In_886,In_81);
nand U2339 (N_2339,In_477,In_681);
and U2340 (N_2340,In_945,In_17);
or U2341 (N_2341,In_373,In_481);
nand U2342 (N_2342,In_100,In_460);
nand U2343 (N_2343,In_229,In_161);
nand U2344 (N_2344,In_316,In_83);
nand U2345 (N_2345,In_594,In_113);
nand U2346 (N_2346,In_690,In_345);
nand U2347 (N_2347,In_151,In_773);
nand U2348 (N_2348,In_484,In_116);
and U2349 (N_2349,In_556,In_627);
nor U2350 (N_2350,In_253,In_478);
or U2351 (N_2351,In_188,In_374);
nand U2352 (N_2352,In_450,In_907);
or U2353 (N_2353,In_495,In_191);
nor U2354 (N_2354,In_435,In_241);
nand U2355 (N_2355,In_308,In_407);
nand U2356 (N_2356,In_332,In_560);
nand U2357 (N_2357,In_682,In_226);
and U2358 (N_2358,In_690,In_425);
or U2359 (N_2359,In_967,In_427);
nand U2360 (N_2360,In_760,In_973);
nand U2361 (N_2361,In_310,In_930);
nor U2362 (N_2362,In_103,In_793);
or U2363 (N_2363,In_4,In_442);
and U2364 (N_2364,In_670,In_73);
or U2365 (N_2365,In_81,In_275);
or U2366 (N_2366,In_861,In_757);
or U2367 (N_2367,In_966,In_369);
and U2368 (N_2368,In_539,In_303);
nor U2369 (N_2369,In_140,In_144);
nor U2370 (N_2370,In_409,In_131);
nor U2371 (N_2371,In_925,In_211);
or U2372 (N_2372,In_19,In_473);
or U2373 (N_2373,In_818,In_709);
nor U2374 (N_2374,In_82,In_36);
and U2375 (N_2375,In_423,In_652);
nor U2376 (N_2376,In_622,In_983);
nor U2377 (N_2377,In_770,In_185);
nor U2378 (N_2378,In_699,In_154);
or U2379 (N_2379,In_369,In_956);
nor U2380 (N_2380,In_348,In_692);
or U2381 (N_2381,In_957,In_825);
nand U2382 (N_2382,In_384,In_284);
nand U2383 (N_2383,In_381,In_665);
nand U2384 (N_2384,In_851,In_160);
nand U2385 (N_2385,In_722,In_465);
and U2386 (N_2386,In_50,In_690);
or U2387 (N_2387,In_681,In_294);
xor U2388 (N_2388,In_916,In_814);
nor U2389 (N_2389,In_937,In_96);
nor U2390 (N_2390,In_537,In_466);
and U2391 (N_2391,In_192,In_67);
nor U2392 (N_2392,In_519,In_22);
and U2393 (N_2393,In_831,In_670);
nor U2394 (N_2394,In_225,In_657);
nor U2395 (N_2395,In_642,In_991);
nor U2396 (N_2396,In_892,In_395);
and U2397 (N_2397,In_639,In_838);
nor U2398 (N_2398,In_134,In_207);
nor U2399 (N_2399,In_451,In_99);
or U2400 (N_2400,In_174,In_587);
and U2401 (N_2401,In_312,In_734);
and U2402 (N_2402,In_625,In_277);
and U2403 (N_2403,In_838,In_614);
nand U2404 (N_2404,In_803,In_2);
xor U2405 (N_2405,In_334,In_103);
nand U2406 (N_2406,In_475,In_684);
nor U2407 (N_2407,In_256,In_314);
nor U2408 (N_2408,In_979,In_389);
nor U2409 (N_2409,In_767,In_323);
or U2410 (N_2410,In_993,In_672);
nor U2411 (N_2411,In_196,In_909);
or U2412 (N_2412,In_638,In_431);
nor U2413 (N_2413,In_996,In_386);
or U2414 (N_2414,In_487,In_823);
or U2415 (N_2415,In_688,In_614);
nor U2416 (N_2416,In_387,In_540);
nand U2417 (N_2417,In_696,In_765);
nand U2418 (N_2418,In_559,In_465);
and U2419 (N_2419,In_96,In_880);
nand U2420 (N_2420,In_261,In_58);
nor U2421 (N_2421,In_466,In_857);
or U2422 (N_2422,In_522,In_647);
and U2423 (N_2423,In_697,In_915);
nand U2424 (N_2424,In_517,In_8);
nor U2425 (N_2425,In_757,In_378);
nor U2426 (N_2426,In_301,In_587);
nor U2427 (N_2427,In_157,In_832);
nand U2428 (N_2428,In_320,In_181);
nor U2429 (N_2429,In_439,In_977);
and U2430 (N_2430,In_864,In_192);
nand U2431 (N_2431,In_349,In_19);
nand U2432 (N_2432,In_717,In_522);
nor U2433 (N_2433,In_183,In_658);
and U2434 (N_2434,In_558,In_376);
and U2435 (N_2435,In_50,In_598);
nor U2436 (N_2436,In_131,In_874);
or U2437 (N_2437,In_930,In_766);
nand U2438 (N_2438,In_436,In_844);
and U2439 (N_2439,In_206,In_445);
nand U2440 (N_2440,In_997,In_385);
or U2441 (N_2441,In_132,In_575);
and U2442 (N_2442,In_920,In_775);
nand U2443 (N_2443,In_748,In_118);
and U2444 (N_2444,In_80,In_706);
and U2445 (N_2445,In_341,In_864);
or U2446 (N_2446,In_602,In_295);
nand U2447 (N_2447,In_236,In_146);
and U2448 (N_2448,In_790,In_862);
and U2449 (N_2449,In_375,In_82);
nor U2450 (N_2450,In_132,In_638);
or U2451 (N_2451,In_536,In_244);
and U2452 (N_2452,In_351,In_897);
or U2453 (N_2453,In_523,In_241);
nand U2454 (N_2454,In_145,In_208);
or U2455 (N_2455,In_185,In_656);
nand U2456 (N_2456,In_625,In_127);
nand U2457 (N_2457,In_179,In_269);
and U2458 (N_2458,In_216,In_855);
nor U2459 (N_2459,In_931,In_541);
or U2460 (N_2460,In_450,In_444);
or U2461 (N_2461,In_251,In_738);
nor U2462 (N_2462,In_238,In_32);
nor U2463 (N_2463,In_894,In_518);
nor U2464 (N_2464,In_158,In_286);
and U2465 (N_2465,In_639,In_140);
nor U2466 (N_2466,In_519,In_804);
xnor U2467 (N_2467,In_418,In_562);
nor U2468 (N_2468,In_724,In_495);
nand U2469 (N_2469,In_482,In_744);
or U2470 (N_2470,In_893,In_884);
or U2471 (N_2471,In_648,In_160);
nor U2472 (N_2472,In_756,In_576);
nor U2473 (N_2473,In_991,In_53);
nand U2474 (N_2474,In_345,In_163);
or U2475 (N_2475,In_316,In_971);
or U2476 (N_2476,In_273,In_809);
or U2477 (N_2477,In_339,In_976);
or U2478 (N_2478,In_22,In_284);
and U2479 (N_2479,In_41,In_931);
nand U2480 (N_2480,In_919,In_63);
nor U2481 (N_2481,In_860,In_67);
nor U2482 (N_2482,In_418,In_185);
nand U2483 (N_2483,In_697,In_750);
or U2484 (N_2484,In_638,In_488);
or U2485 (N_2485,In_219,In_773);
or U2486 (N_2486,In_118,In_309);
and U2487 (N_2487,In_179,In_403);
and U2488 (N_2488,In_305,In_134);
nor U2489 (N_2489,In_517,In_462);
xnor U2490 (N_2490,In_220,In_718);
nor U2491 (N_2491,In_109,In_176);
and U2492 (N_2492,In_88,In_393);
nor U2493 (N_2493,In_13,In_831);
and U2494 (N_2494,In_611,In_478);
nor U2495 (N_2495,In_959,In_710);
and U2496 (N_2496,In_285,In_811);
nor U2497 (N_2497,In_711,In_444);
nand U2498 (N_2498,In_91,In_56);
nand U2499 (N_2499,In_969,In_461);
nand U2500 (N_2500,In_858,In_420);
nand U2501 (N_2501,In_617,In_696);
and U2502 (N_2502,In_260,In_736);
and U2503 (N_2503,In_805,In_153);
and U2504 (N_2504,In_185,In_181);
or U2505 (N_2505,In_693,In_51);
nand U2506 (N_2506,In_445,In_913);
nor U2507 (N_2507,In_508,In_840);
nand U2508 (N_2508,In_138,In_366);
nor U2509 (N_2509,In_517,In_829);
xnor U2510 (N_2510,In_491,In_659);
nor U2511 (N_2511,In_658,In_782);
nor U2512 (N_2512,In_814,In_190);
nor U2513 (N_2513,In_726,In_479);
nand U2514 (N_2514,In_568,In_730);
and U2515 (N_2515,In_594,In_206);
nand U2516 (N_2516,In_822,In_306);
and U2517 (N_2517,In_934,In_417);
or U2518 (N_2518,In_85,In_885);
nor U2519 (N_2519,In_562,In_62);
nand U2520 (N_2520,In_153,In_423);
nand U2521 (N_2521,In_259,In_540);
and U2522 (N_2522,In_354,In_140);
and U2523 (N_2523,In_189,In_648);
and U2524 (N_2524,In_997,In_126);
xnor U2525 (N_2525,In_446,In_646);
and U2526 (N_2526,In_130,In_210);
and U2527 (N_2527,In_55,In_507);
and U2528 (N_2528,In_975,In_267);
or U2529 (N_2529,In_115,In_848);
nand U2530 (N_2530,In_74,In_450);
nand U2531 (N_2531,In_868,In_747);
or U2532 (N_2532,In_435,In_957);
nor U2533 (N_2533,In_501,In_748);
or U2534 (N_2534,In_414,In_805);
or U2535 (N_2535,In_679,In_620);
nand U2536 (N_2536,In_133,In_46);
and U2537 (N_2537,In_630,In_208);
or U2538 (N_2538,In_689,In_314);
or U2539 (N_2539,In_992,In_698);
xor U2540 (N_2540,In_421,In_379);
and U2541 (N_2541,In_630,In_511);
nand U2542 (N_2542,In_82,In_680);
or U2543 (N_2543,In_270,In_936);
or U2544 (N_2544,In_761,In_924);
xnor U2545 (N_2545,In_570,In_902);
or U2546 (N_2546,In_462,In_188);
or U2547 (N_2547,In_459,In_318);
and U2548 (N_2548,In_36,In_335);
and U2549 (N_2549,In_137,In_93);
nand U2550 (N_2550,In_917,In_534);
or U2551 (N_2551,In_115,In_470);
or U2552 (N_2552,In_484,In_503);
or U2553 (N_2553,In_173,In_788);
and U2554 (N_2554,In_683,In_841);
nand U2555 (N_2555,In_905,In_295);
nand U2556 (N_2556,In_308,In_399);
or U2557 (N_2557,In_614,In_800);
and U2558 (N_2558,In_843,In_506);
or U2559 (N_2559,In_842,In_549);
or U2560 (N_2560,In_239,In_156);
nor U2561 (N_2561,In_659,In_341);
or U2562 (N_2562,In_726,In_463);
or U2563 (N_2563,In_147,In_451);
or U2564 (N_2564,In_126,In_952);
or U2565 (N_2565,In_348,In_603);
nor U2566 (N_2566,In_560,In_163);
nor U2567 (N_2567,In_791,In_732);
and U2568 (N_2568,In_966,In_957);
or U2569 (N_2569,In_768,In_796);
nor U2570 (N_2570,In_747,In_839);
or U2571 (N_2571,In_245,In_851);
nand U2572 (N_2572,In_334,In_132);
and U2573 (N_2573,In_992,In_635);
and U2574 (N_2574,In_144,In_990);
and U2575 (N_2575,In_785,In_12);
xnor U2576 (N_2576,In_180,In_810);
or U2577 (N_2577,In_589,In_190);
nor U2578 (N_2578,In_605,In_720);
nand U2579 (N_2579,In_481,In_95);
nand U2580 (N_2580,In_202,In_189);
or U2581 (N_2581,In_889,In_258);
or U2582 (N_2582,In_741,In_208);
and U2583 (N_2583,In_582,In_909);
and U2584 (N_2584,In_252,In_864);
and U2585 (N_2585,In_870,In_231);
nand U2586 (N_2586,In_102,In_557);
nand U2587 (N_2587,In_513,In_871);
nor U2588 (N_2588,In_144,In_728);
nor U2589 (N_2589,In_172,In_611);
and U2590 (N_2590,In_284,In_965);
nand U2591 (N_2591,In_562,In_198);
nand U2592 (N_2592,In_151,In_796);
nor U2593 (N_2593,In_206,In_522);
nor U2594 (N_2594,In_217,In_831);
and U2595 (N_2595,In_793,In_802);
nor U2596 (N_2596,In_567,In_918);
nand U2597 (N_2597,In_336,In_259);
and U2598 (N_2598,In_181,In_177);
or U2599 (N_2599,In_121,In_887);
nand U2600 (N_2600,In_695,In_953);
or U2601 (N_2601,In_943,In_96);
and U2602 (N_2602,In_560,In_522);
and U2603 (N_2603,In_696,In_570);
or U2604 (N_2604,In_151,In_103);
nand U2605 (N_2605,In_172,In_683);
and U2606 (N_2606,In_403,In_106);
nor U2607 (N_2607,In_9,In_77);
or U2608 (N_2608,In_766,In_927);
and U2609 (N_2609,In_961,In_82);
nand U2610 (N_2610,In_564,In_584);
nand U2611 (N_2611,In_131,In_625);
or U2612 (N_2612,In_419,In_706);
nand U2613 (N_2613,In_556,In_912);
nand U2614 (N_2614,In_641,In_285);
nand U2615 (N_2615,In_241,In_29);
or U2616 (N_2616,In_482,In_70);
nand U2617 (N_2617,In_372,In_154);
and U2618 (N_2618,In_680,In_832);
or U2619 (N_2619,In_673,In_317);
or U2620 (N_2620,In_153,In_69);
and U2621 (N_2621,In_326,In_518);
or U2622 (N_2622,In_543,In_53);
or U2623 (N_2623,In_870,In_537);
nor U2624 (N_2624,In_662,In_207);
nand U2625 (N_2625,In_478,In_583);
nor U2626 (N_2626,In_395,In_308);
and U2627 (N_2627,In_638,In_387);
nand U2628 (N_2628,In_851,In_960);
nand U2629 (N_2629,In_607,In_280);
nor U2630 (N_2630,In_409,In_667);
or U2631 (N_2631,In_446,In_724);
nand U2632 (N_2632,In_889,In_381);
nor U2633 (N_2633,In_274,In_369);
nor U2634 (N_2634,In_840,In_736);
nand U2635 (N_2635,In_807,In_882);
nor U2636 (N_2636,In_997,In_384);
or U2637 (N_2637,In_56,In_612);
and U2638 (N_2638,In_537,In_626);
nand U2639 (N_2639,In_654,In_959);
or U2640 (N_2640,In_521,In_434);
nor U2641 (N_2641,In_70,In_636);
nand U2642 (N_2642,In_822,In_387);
nor U2643 (N_2643,In_761,In_866);
nand U2644 (N_2644,In_922,In_969);
nand U2645 (N_2645,In_501,In_552);
nor U2646 (N_2646,In_680,In_967);
nand U2647 (N_2647,In_618,In_979);
nand U2648 (N_2648,In_864,In_906);
nor U2649 (N_2649,In_528,In_680);
and U2650 (N_2650,In_491,In_850);
and U2651 (N_2651,In_692,In_250);
nand U2652 (N_2652,In_69,In_676);
nand U2653 (N_2653,In_120,In_194);
or U2654 (N_2654,In_490,In_676);
and U2655 (N_2655,In_917,In_295);
and U2656 (N_2656,In_45,In_163);
nor U2657 (N_2657,In_92,In_38);
and U2658 (N_2658,In_683,In_415);
nor U2659 (N_2659,In_959,In_830);
or U2660 (N_2660,In_377,In_612);
or U2661 (N_2661,In_445,In_825);
nor U2662 (N_2662,In_841,In_106);
nor U2663 (N_2663,In_662,In_801);
nand U2664 (N_2664,In_223,In_664);
and U2665 (N_2665,In_944,In_999);
and U2666 (N_2666,In_359,In_134);
or U2667 (N_2667,In_312,In_180);
and U2668 (N_2668,In_130,In_646);
nand U2669 (N_2669,In_139,In_260);
or U2670 (N_2670,In_249,In_465);
or U2671 (N_2671,In_54,In_765);
or U2672 (N_2672,In_128,In_953);
nand U2673 (N_2673,In_313,In_182);
nor U2674 (N_2674,In_873,In_568);
and U2675 (N_2675,In_603,In_279);
nand U2676 (N_2676,In_347,In_422);
or U2677 (N_2677,In_860,In_353);
and U2678 (N_2678,In_69,In_342);
nand U2679 (N_2679,In_36,In_46);
and U2680 (N_2680,In_135,In_237);
or U2681 (N_2681,In_913,In_192);
nand U2682 (N_2682,In_855,In_515);
nand U2683 (N_2683,In_747,In_116);
nor U2684 (N_2684,In_299,In_503);
nor U2685 (N_2685,In_571,In_476);
nor U2686 (N_2686,In_320,In_521);
and U2687 (N_2687,In_56,In_533);
nand U2688 (N_2688,In_184,In_810);
nand U2689 (N_2689,In_95,In_13);
xor U2690 (N_2690,In_246,In_777);
and U2691 (N_2691,In_433,In_63);
nor U2692 (N_2692,In_790,In_712);
nor U2693 (N_2693,In_712,In_320);
nor U2694 (N_2694,In_38,In_391);
nor U2695 (N_2695,In_940,In_478);
nor U2696 (N_2696,In_610,In_165);
nor U2697 (N_2697,In_152,In_237);
nor U2698 (N_2698,In_755,In_955);
nor U2699 (N_2699,In_137,In_540);
or U2700 (N_2700,In_601,In_365);
or U2701 (N_2701,In_395,In_517);
nor U2702 (N_2702,In_536,In_645);
or U2703 (N_2703,In_931,In_579);
nand U2704 (N_2704,In_730,In_190);
nand U2705 (N_2705,In_337,In_786);
or U2706 (N_2706,In_570,In_977);
and U2707 (N_2707,In_445,In_494);
and U2708 (N_2708,In_199,In_405);
nand U2709 (N_2709,In_366,In_458);
or U2710 (N_2710,In_600,In_529);
or U2711 (N_2711,In_657,In_98);
and U2712 (N_2712,In_505,In_180);
and U2713 (N_2713,In_899,In_906);
and U2714 (N_2714,In_81,In_524);
and U2715 (N_2715,In_756,In_789);
and U2716 (N_2716,In_109,In_849);
nor U2717 (N_2717,In_335,In_714);
and U2718 (N_2718,In_241,In_477);
nand U2719 (N_2719,In_799,In_810);
nor U2720 (N_2720,In_138,In_748);
or U2721 (N_2721,In_458,In_159);
or U2722 (N_2722,In_97,In_508);
nand U2723 (N_2723,In_551,In_132);
nor U2724 (N_2724,In_128,In_546);
and U2725 (N_2725,In_942,In_674);
or U2726 (N_2726,In_967,In_38);
nand U2727 (N_2727,In_938,In_729);
nor U2728 (N_2728,In_200,In_825);
and U2729 (N_2729,In_880,In_713);
nand U2730 (N_2730,In_705,In_594);
nand U2731 (N_2731,In_832,In_816);
or U2732 (N_2732,In_671,In_786);
and U2733 (N_2733,In_731,In_580);
nor U2734 (N_2734,In_984,In_10);
nand U2735 (N_2735,In_239,In_157);
xnor U2736 (N_2736,In_539,In_893);
or U2737 (N_2737,In_755,In_583);
or U2738 (N_2738,In_656,In_555);
or U2739 (N_2739,In_420,In_19);
or U2740 (N_2740,In_85,In_803);
nand U2741 (N_2741,In_687,In_342);
or U2742 (N_2742,In_130,In_829);
and U2743 (N_2743,In_986,In_868);
or U2744 (N_2744,In_273,In_503);
nor U2745 (N_2745,In_540,In_446);
or U2746 (N_2746,In_463,In_691);
or U2747 (N_2747,In_315,In_801);
and U2748 (N_2748,In_295,In_113);
nand U2749 (N_2749,In_373,In_65);
or U2750 (N_2750,In_954,In_81);
nor U2751 (N_2751,In_843,In_601);
nand U2752 (N_2752,In_792,In_764);
nand U2753 (N_2753,In_603,In_806);
nand U2754 (N_2754,In_750,In_470);
and U2755 (N_2755,In_253,In_504);
nand U2756 (N_2756,In_696,In_217);
or U2757 (N_2757,In_801,In_444);
nor U2758 (N_2758,In_769,In_230);
or U2759 (N_2759,In_141,In_995);
and U2760 (N_2760,In_838,In_901);
or U2761 (N_2761,In_755,In_575);
and U2762 (N_2762,In_90,In_252);
nor U2763 (N_2763,In_714,In_734);
and U2764 (N_2764,In_963,In_741);
and U2765 (N_2765,In_437,In_743);
or U2766 (N_2766,In_492,In_723);
nand U2767 (N_2767,In_901,In_238);
and U2768 (N_2768,In_439,In_503);
nor U2769 (N_2769,In_364,In_75);
or U2770 (N_2770,In_634,In_496);
nor U2771 (N_2771,In_184,In_590);
nor U2772 (N_2772,In_416,In_353);
or U2773 (N_2773,In_124,In_889);
nand U2774 (N_2774,In_840,In_614);
nand U2775 (N_2775,In_732,In_742);
nor U2776 (N_2776,In_518,In_606);
nand U2777 (N_2777,In_796,In_844);
nor U2778 (N_2778,In_689,In_64);
or U2779 (N_2779,In_375,In_259);
and U2780 (N_2780,In_645,In_145);
or U2781 (N_2781,In_997,In_68);
and U2782 (N_2782,In_916,In_617);
nand U2783 (N_2783,In_321,In_848);
or U2784 (N_2784,In_12,In_923);
and U2785 (N_2785,In_986,In_943);
nor U2786 (N_2786,In_812,In_920);
nand U2787 (N_2787,In_108,In_727);
and U2788 (N_2788,In_462,In_838);
nor U2789 (N_2789,In_709,In_814);
or U2790 (N_2790,In_412,In_997);
nor U2791 (N_2791,In_753,In_473);
nand U2792 (N_2792,In_289,In_99);
and U2793 (N_2793,In_88,In_202);
nor U2794 (N_2794,In_245,In_790);
nand U2795 (N_2795,In_777,In_465);
nand U2796 (N_2796,In_863,In_524);
nor U2797 (N_2797,In_888,In_314);
and U2798 (N_2798,In_470,In_664);
or U2799 (N_2799,In_721,In_402);
or U2800 (N_2800,In_868,In_941);
nor U2801 (N_2801,In_22,In_469);
or U2802 (N_2802,In_246,In_331);
and U2803 (N_2803,In_1,In_342);
or U2804 (N_2804,In_710,In_682);
and U2805 (N_2805,In_711,In_800);
and U2806 (N_2806,In_906,In_848);
or U2807 (N_2807,In_883,In_418);
nor U2808 (N_2808,In_216,In_617);
and U2809 (N_2809,In_608,In_498);
xnor U2810 (N_2810,In_820,In_522);
nor U2811 (N_2811,In_808,In_16);
nand U2812 (N_2812,In_30,In_444);
nand U2813 (N_2813,In_863,In_784);
or U2814 (N_2814,In_163,In_845);
and U2815 (N_2815,In_196,In_416);
nor U2816 (N_2816,In_130,In_750);
nand U2817 (N_2817,In_724,In_443);
and U2818 (N_2818,In_778,In_597);
or U2819 (N_2819,In_172,In_174);
nand U2820 (N_2820,In_629,In_569);
and U2821 (N_2821,In_642,In_370);
nand U2822 (N_2822,In_453,In_927);
or U2823 (N_2823,In_722,In_495);
and U2824 (N_2824,In_987,In_678);
nor U2825 (N_2825,In_824,In_854);
or U2826 (N_2826,In_136,In_607);
nand U2827 (N_2827,In_3,In_268);
and U2828 (N_2828,In_774,In_98);
or U2829 (N_2829,In_790,In_710);
nor U2830 (N_2830,In_161,In_817);
and U2831 (N_2831,In_963,In_82);
or U2832 (N_2832,In_996,In_607);
nand U2833 (N_2833,In_597,In_306);
and U2834 (N_2834,In_232,In_570);
or U2835 (N_2835,In_545,In_119);
nand U2836 (N_2836,In_590,In_877);
nand U2837 (N_2837,In_371,In_357);
or U2838 (N_2838,In_818,In_617);
nor U2839 (N_2839,In_778,In_47);
and U2840 (N_2840,In_273,In_784);
or U2841 (N_2841,In_911,In_405);
nand U2842 (N_2842,In_409,In_966);
nand U2843 (N_2843,In_344,In_59);
nand U2844 (N_2844,In_964,In_204);
and U2845 (N_2845,In_119,In_182);
nand U2846 (N_2846,In_292,In_202);
or U2847 (N_2847,In_513,In_879);
nor U2848 (N_2848,In_710,In_355);
or U2849 (N_2849,In_72,In_567);
nand U2850 (N_2850,In_914,In_499);
or U2851 (N_2851,In_159,In_339);
and U2852 (N_2852,In_548,In_149);
or U2853 (N_2853,In_500,In_220);
and U2854 (N_2854,In_184,In_690);
or U2855 (N_2855,In_782,In_17);
nand U2856 (N_2856,In_750,In_458);
nand U2857 (N_2857,In_940,In_648);
nand U2858 (N_2858,In_474,In_492);
nor U2859 (N_2859,In_672,In_496);
or U2860 (N_2860,In_451,In_165);
and U2861 (N_2861,In_363,In_459);
nor U2862 (N_2862,In_605,In_598);
nand U2863 (N_2863,In_376,In_967);
nor U2864 (N_2864,In_992,In_606);
and U2865 (N_2865,In_268,In_310);
nor U2866 (N_2866,In_985,In_805);
nor U2867 (N_2867,In_292,In_898);
or U2868 (N_2868,In_373,In_927);
nand U2869 (N_2869,In_828,In_76);
and U2870 (N_2870,In_190,In_721);
or U2871 (N_2871,In_441,In_452);
nand U2872 (N_2872,In_366,In_483);
or U2873 (N_2873,In_309,In_20);
nand U2874 (N_2874,In_475,In_788);
xnor U2875 (N_2875,In_276,In_551);
nand U2876 (N_2876,In_133,In_80);
or U2877 (N_2877,In_157,In_257);
or U2878 (N_2878,In_786,In_506);
and U2879 (N_2879,In_995,In_561);
nor U2880 (N_2880,In_612,In_281);
or U2881 (N_2881,In_557,In_292);
and U2882 (N_2882,In_177,In_290);
or U2883 (N_2883,In_446,In_52);
nor U2884 (N_2884,In_651,In_17);
nand U2885 (N_2885,In_631,In_735);
and U2886 (N_2886,In_627,In_316);
and U2887 (N_2887,In_956,In_153);
and U2888 (N_2888,In_579,In_433);
or U2889 (N_2889,In_719,In_721);
nand U2890 (N_2890,In_925,In_770);
nand U2891 (N_2891,In_90,In_412);
nand U2892 (N_2892,In_978,In_258);
nand U2893 (N_2893,In_306,In_128);
nand U2894 (N_2894,In_77,In_689);
nand U2895 (N_2895,In_487,In_191);
nand U2896 (N_2896,In_31,In_289);
nand U2897 (N_2897,In_546,In_195);
and U2898 (N_2898,In_364,In_320);
and U2899 (N_2899,In_278,In_750);
or U2900 (N_2900,In_594,In_778);
nor U2901 (N_2901,In_3,In_494);
and U2902 (N_2902,In_418,In_817);
nor U2903 (N_2903,In_20,In_213);
nand U2904 (N_2904,In_180,In_584);
or U2905 (N_2905,In_681,In_596);
nor U2906 (N_2906,In_519,In_146);
and U2907 (N_2907,In_288,In_259);
and U2908 (N_2908,In_479,In_512);
and U2909 (N_2909,In_461,In_364);
nand U2910 (N_2910,In_817,In_97);
and U2911 (N_2911,In_565,In_945);
nand U2912 (N_2912,In_320,In_816);
and U2913 (N_2913,In_648,In_393);
nor U2914 (N_2914,In_559,In_532);
or U2915 (N_2915,In_129,In_554);
nor U2916 (N_2916,In_430,In_8);
nand U2917 (N_2917,In_876,In_313);
and U2918 (N_2918,In_219,In_264);
nand U2919 (N_2919,In_551,In_828);
or U2920 (N_2920,In_135,In_762);
and U2921 (N_2921,In_808,In_762);
nand U2922 (N_2922,In_499,In_471);
or U2923 (N_2923,In_624,In_104);
and U2924 (N_2924,In_260,In_579);
or U2925 (N_2925,In_161,In_281);
nor U2926 (N_2926,In_157,In_982);
nor U2927 (N_2927,In_523,In_399);
nand U2928 (N_2928,In_676,In_812);
nand U2929 (N_2929,In_264,In_39);
or U2930 (N_2930,In_40,In_168);
and U2931 (N_2931,In_778,In_843);
or U2932 (N_2932,In_532,In_47);
or U2933 (N_2933,In_153,In_890);
or U2934 (N_2934,In_106,In_588);
nor U2935 (N_2935,In_680,In_179);
nor U2936 (N_2936,In_18,In_942);
and U2937 (N_2937,In_995,In_542);
nand U2938 (N_2938,In_914,In_378);
or U2939 (N_2939,In_783,In_786);
or U2940 (N_2940,In_81,In_394);
or U2941 (N_2941,In_968,In_5);
and U2942 (N_2942,In_339,In_144);
nor U2943 (N_2943,In_974,In_913);
nand U2944 (N_2944,In_920,In_169);
nand U2945 (N_2945,In_806,In_298);
nand U2946 (N_2946,In_238,In_104);
and U2947 (N_2947,In_316,In_249);
nand U2948 (N_2948,In_189,In_768);
and U2949 (N_2949,In_468,In_241);
nor U2950 (N_2950,In_472,In_398);
nor U2951 (N_2951,In_716,In_249);
and U2952 (N_2952,In_983,In_60);
nand U2953 (N_2953,In_566,In_186);
or U2954 (N_2954,In_260,In_711);
or U2955 (N_2955,In_223,In_40);
nor U2956 (N_2956,In_977,In_731);
or U2957 (N_2957,In_502,In_78);
or U2958 (N_2958,In_317,In_242);
nand U2959 (N_2959,In_252,In_542);
and U2960 (N_2960,In_473,In_68);
nand U2961 (N_2961,In_961,In_158);
nand U2962 (N_2962,In_780,In_510);
nor U2963 (N_2963,In_155,In_382);
nor U2964 (N_2964,In_592,In_665);
nor U2965 (N_2965,In_957,In_249);
nand U2966 (N_2966,In_336,In_96);
nand U2967 (N_2967,In_164,In_462);
and U2968 (N_2968,In_209,In_350);
and U2969 (N_2969,In_378,In_973);
nand U2970 (N_2970,In_640,In_261);
and U2971 (N_2971,In_956,In_858);
nor U2972 (N_2972,In_159,In_879);
and U2973 (N_2973,In_274,In_679);
nand U2974 (N_2974,In_213,In_418);
nand U2975 (N_2975,In_930,In_475);
nor U2976 (N_2976,In_930,In_940);
nor U2977 (N_2977,In_410,In_898);
and U2978 (N_2978,In_872,In_305);
nor U2979 (N_2979,In_481,In_214);
nand U2980 (N_2980,In_968,In_521);
nand U2981 (N_2981,In_895,In_260);
nand U2982 (N_2982,In_633,In_770);
and U2983 (N_2983,In_104,In_845);
and U2984 (N_2984,In_337,In_236);
or U2985 (N_2985,In_485,In_615);
or U2986 (N_2986,In_536,In_538);
or U2987 (N_2987,In_714,In_574);
nand U2988 (N_2988,In_569,In_592);
or U2989 (N_2989,In_66,In_785);
nand U2990 (N_2990,In_819,In_568);
nand U2991 (N_2991,In_192,In_425);
and U2992 (N_2992,In_103,In_557);
nor U2993 (N_2993,In_218,In_990);
or U2994 (N_2994,In_521,In_608);
nor U2995 (N_2995,In_390,In_279);
or U2996 (N_2996,In_143,In_938);
or U2997 (N_2997,In_119,In_653);
nand U2998 (N_2998,In_994,In_51);
or U2999 (N_2999,In_711,In_726);
and U3000 (N_3000,In_542,In_715);
nand U3001 (N_3001,In_458,In_453);
nor U3002 (N_3002,In_866,In_216);
and U3003 (N_3003,In_496,In_775);
nor U3004 (N_3004,In_432,In_569);
nor U3005 (N_3005,In_877,In_738);
and U3006 (N_3006,In_288,In_547);
nand U3007 (N_3007,In_339,In_838);
nor U3008 (N_3008,In_204,In_872);
or U3009 (N_3009,In_787,In_134);
nor U3010 (N_3010,In_816,In_187);
xor U3011 (N_3011,In_591,In_176);
and U3012 (N_3012,In_105,In_287);
nor U3013 (N_3013,In_169,In_966);
nand U3014 (N_3014,In_430,In_334);
nor U3015 (N_3015,In_592,In_141);
or U3016 (N_3016,In_158,In_578);
nor U3017 (N_3017,In_10,In_49);
or U3018 (N_3018,In_924,In_594);
and U3019 (N_3019,In_11,In_554);
or U3020 (N_3020,In_201,In_505);
nor U3021 (N_3021,In_373,In_348);
and U3022 (N_3022,In_213,In_18);
and U3023 (N_3023,In_722,In_630);
and U3024 (N_3024,In_685,In_898);
nor U3025 (N_3025,In_376,In_761);
nor U3026 (N_3026,In_949,In_487);
nor U3027 (N_3027,In_820,In_114);
nor U3028 (N_3028,In_347,In_515);
nand U3029 (N_3029,In_117,In_239);
nand U3030 (N_3030,In_297,In_434);
nand U3031 (N_3031,In_11,In_201);
or U3032 (N_3032,In_487,In_161);
and U3033 (N_3033,In_476,In_849);
nor U3034 (N_3034,In_85,In_221);
nor U3035 (N_3035,In_277,In_749);
nor U3036 (N_3036,In_320,In_196);
nand U3037 (N_3037,In_819,In_965);
nor U3038 (N_3038,In_762,In_790);
and U3039 (N_3039,In_991,In_474);
nor U3040 (N_3040,In_338,In_894);
nor U3041 (N_3041,In_930,In_377);
or U3042 (N_3042,In_982,In_154);
and U3043 (N_3043,In_695,In_216);
nand U3044 (N_3044,In_647,In_461);
nand U3045 (N_3045,In_892,In_414);
and U3046 (N_3046,In_757,In_734);
nor U3047 (N_3047,In_838,In_724);
and U3048 (N_3048,In_693,In_224);
nor U3049 (N_3049,In_725,In_874);
or U3050 (N_3050,In_334,In_312);
nand U3051 (N_3051,In_678,In_721);
and U3052 (N_3052,In_972,In_995);
nor U3053 (N_3053,In_301,In_73);
or U3054 (N_3054,In_976,In_118);
nand U3055 (N_3055,In_855,In_664);
nand U3056 (N_3056,In_63,In_176);
and U3057 (N_3057,In_952,In_307);
and U3058 (N_3058,In_235,In_966);
and U3059 (N_3059,In_559,In_656);
or U3060 (N_3060,In_441,In_290);
nor U3061 (N_3061,In_15,In_687);
or U3062 (N_3062,In_174,In_670);
nand U3063 (N_3063,In_175,In_541);
nand U3064 (N_3064,In_974,In_420);
nor U3065 (N_3065,In_564,In_539);
or U3066 (N_3066,In_60,In_262);
nand U3067 (N_3067,In_646,In_613);
and U3068 (N_3068,In_684,In_384);
nand U3069 (N_3069,In_481,In_538);
nand U3070 (N_3070,In_680,In_892);
or U3071 (N_3071,In_990,In_76);
or U3072 (N_3072,In_282,In_868);
or U3073 (N_3073,In_895,In_999);
nor U3074 (N_3074,In_287,In_888);
and U3075 (N_3075,In_560,In_673);
nand U3076 (N_3076,In_950,In_101);
nor U3077 (N_3077,In_805,In_653);
or U3078 (N_3078,In_436,In_766);
xor U3079 (N_3079,In_833,In_905);
or U3080 (N_3080,In_445,In_121);
or U3081 (N_3081,In_877,In_399);
xor U3082 (N_3082,In_647,In_515);
nand U3083 (N_3083,In_611,In_451);
nand U3084 (N_3084,In_776,In_787);
or U3085 (N_3085,In_688,In_860);
or U3086 (N_3086,In_348,In_762);
nand U3087 (N_3087,In_716,In_347);
nor U3088 (N_3088,In_381,In_591);
and U3089 (N_3089,In_878,In_220);
and U3090 (N_3090,In_131,In_541);
nor U3091 (N_3091,In_94,In_225);
nand U3092 (N_3092,In_326,In_521);
and U3093 (N_3093,In_316,In_653);
or U3094 (N_3094,In_616,In_973);
nand U3095 (N_3095,In_187,In_442);
nor U3096 (N_3096,In_594,In_895);
nand U3097 (N_3097,In_558,In_859);
nor U3098 (N_3098,In_13,In_298);
and U3099 (N_3099,In_840,In_893);
nand U3100 (N_3100,In_829,In_258);
or U3101 (N_3101,In_510,In_425);
nand U3102 (N_3102,In_582,In_70);
or U3103 (N_3103,In_169,In_1);
nor U3104 (N_3104,In_693,In_690);
and U3105 (N_3105,In_150,In_101);
or U3106 (N_3106,In_259,In_203);
nand U3107 (N_3107,In_261,In_733);
and U3108 (N_3108,In_36,In_410);
or U3109 (N_3109,In_300,In_889);
nand U3110 (N_3110,In_856,In_527);
nand U3111 (N_3111,In_473,In_149);
or U3112 (N_3112,In_696,In_800);
and U3113 (N_3113,In_909,In_944);
nand U3114 (N_3114,In_219,In_929);
and U3115 (N_3115,In_258,In_852);
and U3116 (N_3116,In_287,In_400);
nand U3117 (N_3117,In_876,In_400);
nor U3118 (N_3118,In_642,In_397);
and U3119 (N_3119,In_181,In_535);
nand U3120 (N_3120,In_368,In_238);
nand U3121 (N_3121,In_652,In_180);
nor U3122 (N_3122,In_190,In_680);
and U3123 (N_3123,In_579,In_452);
nand U3124 (N_3124,In_131,In_328);
and U3125 (N_3125,In_256,In_320);
and U3126 (N_3126,In_612,In_702);
or U3127 (N_3127,In_647,In_419);
nor U3128 (N_3128,In_232,In_750);
nand U3129 (N_3129,In_311,In_911);
nor U3130 (N_3130,In_51,In_102);
nand U3131 (N_3131,In_716,In_829);
or U3132 (N_3132,In_730,In_651);
nor U3133 (N_3133,In_834,In_119);
nor U3134 (N_3134,In_871,In_55);
nand U3135 (N_3135,In_326,In_419);
or U3136 (N_3136,In_58,In_544);
or U3137 (N_3137,In_922,In_876);
and U3138 (N_3138,In_390,In_181);
nand U3139 (N_3139,In_662,In_20);
and U3140 (N_3140,In_36,In_145);
and U3141 (N_3141,In_248,In_712);
nand U3142 (N_3142,In_360,In_526);
or U3143 (N_3143,In_799,In_533);
or U3144 (N_3144,In_284,In_648);
nor U3145 (N_3145,In_968,In_278);
and U3146 (N_3146,In_495,In_463);
and U3147 (N_3147,In_600,In_482);
nor U3148 (N_3148,In_409,In_833);
and U3149 (N_3149,In_200,In_367);
nand U3150 (N_3150,In_870,In_28);
or U3151 (N_3151,In_118,In_144);
and U3152 (N_3152,In_798,In_39);
and U3153 (N_3153,In_332,In_784);
nor U3154 (N_3154,In_553,In_152);
or U3155 (N_3155,In_37,In_197);
nand U3156 (N_3156,In_157,In_516);
nor U3157 (N_3157,In_110,In_187);
or U3158 (N_3158,In_389,In_81);
nand U3159 (N_3159,In_727,In_620);
nor U3160 (N_3160,In_424,In_738);
nor U3161 (N_3161,In_680,In_498);
nand U3162 (N_3162,In_449,In_92);
or U3163 (N_3163,In_403,In_927);
or U3164 (N_3164,In_681,In_924);
or U3165 (N_3165,In_783,In_859);
and U3166 (N_3166,In_19,In_268);
nand U3167 (N_3167,In_636,In_360);
or U3168 (N_3168,In_46,In_876);
or U3169 (N_3169,In_497,In_518);
nor U3170 (N_3170,In_880,In_439);
nand U3171 (N_3171,In_598,In_144);
and U3172 (N_3172,In_310,In_657);
or U3173 (N_3173,In_496,In_588);
nand U3174 (N_3174,In_909,In_556);
or U3175 (N_3175,In_535,In_257);
nor U3176 (N_3176,In_840,In_482);
and U3177 (N_3177,In_446,In_894);
nor U3178 (N_3178,In_73,In_151);
or U3179 (N_3179,In_263,In_77);
nor U3180 (N_3180,In_942,In_610);
or U3181 (N_3181,In_930,In_540);
or U3182 (N_3182,In_232,In_4);
nor U3183 (N_3183,In_198,In_573);
nand U3184 (N_3184,In_697,In_802);
nand U3185 (N_3185,In_992,In_932);
nor U3186 (N_3186,In_401,In_253);
nor U3187 (N_3187,In_296,In_455);
or U3188 (N_3188,In_397,In_227);
or U3189 (N_3189,In_377,In_265);
and U3190 (N_3190,In_312,In_430);
and U3191 (N_3191,In_693,In_309);
or U3192 (N_3192,In_79,In_812);
or U3193 (N_3193,In_922,In_425);
nor U3194 (N_3194,In_297,In_433);
and U3195 (N_3195,In_543,In_62);
nor U3196 (N_3196,In_962,In_811);
nand U3197 (N_3197,In_547,In_836);
nand U3198 (N_3198,In_768,In_985);
or U3199 (N_3199,In_388,In_692);
and U3200 (N_3200,In_648,In_989);
and U3201 (N_3201,In_3,In_790);
and U3202 (N_3202,In_968,In_309);
nand U3203 (N_3203,In_489,In_70);
or U3204 (N_3204,In_8,In_105);
nor U3205 (N_3205,In_293,In_619);
or U3206 (N_3206,In_245,In_126);
nand U3207 (N_3207,In_20,In_657);
or U3208 (N_3208,In_266,In_259);
nor U3209 (N_3209,In_116,In_890);
nand U3210 (N_3210,In_454,In_725);
or U3211 (N_3211,In_657,In_311);
or U3212 (N_3212,In_885,In_235);
nand U3213 (N_3213,In_498,In_542);
and U3214 (N_3214,In_63,In_244);
or U3215 (N_3215,In_989,In_592);
and U3216 (N_3216,In_368,In_592);
nand U3217 (N_3217,In_711,In_354);
nor U3218 (N_3218,In_828,In_109);
nor U3219 (N_3219,In_532,In_530);
or U3220 (N_3220,In_722,In_598);
and U3221 (N_3221,In_651,In_804);
and U3222 (N_3222,In_402,In_731);
or U3223 (N_3223,In_950,In_65);
nand U3224 (N_3224,In_889,In_850);
nor U3225 (N_3225,In_861,In_127);
nor U3226 (N_3226,In_555,In_206);
nand U3227 (N_3227,In_544,In_673);
and U3228 (N_3228,In_796,In_658);
nor U3229 (N_3229,In_625,In_335);
and U3230 (N_3230,In_146,In_443);
and U3231 (N_3231,In_743,In_29);
nand U3232 (N_3232,In_50,In_376);
or U3233 (N_3233,In_427,In_134);
nand U3234 (N_3234,In_267,In_344);
or U3235 (N_3235,In_186,In_134);
or U3236 (N_3236,In_586,In_116);
or U3237 (N_3237,In_711,In_68);
or U3238 (N_3238,In_890,In_55);
nor U3239 (N_3239,In_992,In_718);
and U3240 (N_3240,In_623,In_496);
nor U3241 (N_3241,In_725,In_175);
nand U3242 (N_3242,In_246,In_868);
nor U3243 (N_3243,In_578,In_586);
nand U3244 (N_3244,In_190,In_837);
or U3245 (N_3245,In_508,In_768);
or U3246 (N_3246,In_91,In_102);
nand U3247 (N_3247,In_555,In_404);
nor U3248 (N_3248,In_901,In_920);
nand U3249 (N_3249,In_445,In_539);
nor U3250 (N_3250,In_615,In_728);
nor U3251 (N_3251,In_466,In_584);
nor U3252 (N_3252,In_459,In_725);
or U3253 (N_3253,In_94,In_793);
or U3254 (N_3254,In_804,In_502);
or U3255 (N_3255,In_403,In_111);
nand U3256 (N_3256,In_960,In_465);
nor U3257 (N_3257,In_319,In_309);
nor U3258 (N_3258,In_719,In_144);
nand U3259 (N_3259,In_256,In_219);
or U3260 (N_3260,In_491,In_125);
nor U3261 (N_3261,In_973,In_67);
nand U3262 (N_3262,In_57,In_133);
or U3263 (N_3263,In_342,In_547);
and U3264 (N_3264,In_758,In_437);
nor U3265 (N_3265,In_761,In_609);
or U3266 (N_3266,In_959,In_415);
or U3267 (N_3267,In_569,In_439);
or U3268 (N_3268,In_770,In_431);
nor U3269 (N_3269,In_179,In_349);
and U3270 (N_3270,In_330,In_797);
nor U3271 (N_3271,In_142,In_935);
or U3272 (N_3272,In_437,In_830);
or U3273 (N_3273,In_150,In_210);
nor U3274 (N_3274,In_251,In_785);
and U3275 (N_3275,In_882,In_733);
nor U3276 (N_3276,In_471,In_107);
xnor U3277 (N_3277,In_750,In_927);
or U3278 (N_3278,In_601,In_113);
or U3279 (N_3279,In_166,In_611);
and U3280 (N_3280,In_692,In_846);
nand U3281 (N_3281,In_365,In_618);
or U3282 (N_3282,In_577,In_407);
nor U3283 (N_3283,In_859,In_557);
or U3284 (N_3284,In_898,In_312);
and U3285 (N_3285,In_866,In_508);
nand U3286 (N_3286,In_156,In_387);
or U3287 (N_3287,In_347,In_841);
nand U3288 (N_3288,In_836,In_988);
nor U3289 (N_3289,In_411,In_999);
nor U3290 (N_3290,In_391,In_40);
or U3291 (N_3291,In_997,In_246);
or U3292 (N_3292,In_831,In_642);
nor U3293 (N_3293,In_630,In_157);
or U3294 (N_3294,In_872,In_247);
and U3295 (N_3295,In_192,In_619);
and U3296 (N_3296,In_931,In_217);
and U3297 (N_3297,In_691,In_494);
or U3298 (N_3298,In_87,In_351);
nand U3299 (N_3299,In_743,In_845);
nand U3300 (N_3300,In_208,In_671);
nor U3301 (N_3301,In_802,In_308);
nor U3302 (N_3302,In_369,In_247);
nand U3303 (N_3303,In_98,In_930);
and U3304 (N_3304,In_321,In_156);
nand U3305 (N_3305,In_896,In_817);
nor U3306 (N_3306,In_694,In_261);
nand U3307 (N_3307,In_269,In_136);
and U3308 (N_3308,In_39,In_866);
nor U3309 (N_3309,In_322,In_439);
or U3310 (N_3310,In_717,In_631);
and U3311 (N_3311,In_688,In_548);
nor U3312 (N_3312,In_837,In_770);
nor U3313 (N_3313,In_113,In_264);
nor U3314 (N_3314,In_659,In_955);
or U3315 (N_3315,In_208,In_85);
nand U3316 (N_3316,In_735,In_521);
and U3317 (N_3317,In_821,In_896);
nand U3318 (N_3318,In_576,In_154);
nor U3319 (N_3319,In_326,In_905);
nand U3320 (N_3320,In_946,In_350);
or U3321 (N_3321,In_795,In_984);
or U3322 (N_3322,In_928,In_854);
nand U3323 (N_3323,In_477,In_33);
nand U3324 (N_3324,In_681,In_539);
nand U3325 (N_3325,In_983,In_248);
nor U3326 (N_3326,In_960,In_251);
nand U3327 (N_3327,In_692,In_226);
and U3328 (N_3328,In_292,In_875);
and U3329 (N_3329,In_183,In_980);
nand U3330 (N_3330,In_874,In_195);
or U3331 (N_3331,In_699,In_257);
nor U3332 (N_3332,In_960,In_429);
and U3333 (N_3333,In_183,In_955);
nand U3334 (N_3334,In_917,In_387);
and U3335 (N_3335,In_58,In_994);
and U3336 (N_3336,In_856,In_381);
and U3337 (N_3337,In_941,In_151);
and U3338 (N_3338,In_785,In_845);
or U3339 (N_3339,In_107,In_966);
and U3340 (N_3340,In_522,In_637);
nand U3341 (N_3341,In_739,In_522);
nor U3342 (N_3342,In_79,In_292);
nand U3343 (N_3343,In_573,In_834);
or U3344 (N_3344,In_760,In_885);
nor U3345 (N_3345,In_762,In_641);
and U3346 (N_3346,In_615,In_947);
nand U3347 (N_3347,In_529,In_940);
and U3348 (N_3348,In_974,In_767);
nand U3349 (N_3349,In_693,In_371);
and U3350 (N_3350,In_489,In_88);
or U3351 (N_3351,In_237,In_498);
or U3352 (N_3352,In_236,In_151);
nand U3353 (N_3353,In_465,In_772);
or U3354 (N_3354,In_760,In_611);
and U3355 (N_3355,In_748,In_551);
or U3356 (N_3356,In_131,In_301);
and U3357 (N_3357,In_26,In_18);
nor U3358 (N_3358,In_623,In_379);
or U3359 (N_3359,In_820,In_8);
xnor U3360 (N_3360,In_866,In_835);
or U3361 (N_3361,In_43,In_426);
or U3362 (N_3362,In_145,In_366);
or U3363 (N_3363,In_371,In_738);
nor U3364 (N_3364,In_762,In_654);
nand U3365 (N_3365,In_552,In_844);
and U3366 (N_3366,In_516,In_109);
nand U3367 (N_3367,In_74,In_42);
nand U3368 (N_3368,In_908,In_410);
or U3369 (N_3369,In_799,In_745);
nor U3370 (N_3370,In_34,In_795);
nor U3371 (N_3371,In_66,In_116);
and U3372 (N_3372,In_438,In_258);
and U3373 (N_3373,In_340,In_446);
xor U3374 (N_3374,In_50,In_758);
and U3375 (N_3375,In_620,In_317);
and U3376 (N_3376,In_483,In_62);
and U3377 (N_3377,In_404,In_241);
nor U3378 (N_3378,In_452,In_605);
or U3379 (N_3379,In_305,In_857);
or U3380 (N_3380,In_820,In_220);
nor U3381 (N_3381,In_321,In_282);
nand U3382 (N_3382,In_148,In_469);
nor U3383 (N_3383,In_631,In_957);
or U3384 (N_3384,In_51,In_228);
and U3385 (N_3385,In_672,In_447);
nand U3386 (N_3386,In_52,In_488);
nor U3387 (N_3387,In_866,In_659);
nor U3388 (N_3388,In_307,In_161);
nor U3389 (N_3389,In_273,In_979);
nor U3390 (N_3390,In_837,In_930);
nand U3391 (N_3391,In_400,In_765);
and U3392 (N_3392,In_884,In_239);
and U3393 (N_3393,In_468,In_155);
or U3394 (N_3394,In_299,In_174);
or U3395 (N_3395,In_96,In_455);
nand U3396 (N_3396,In_179,In_984);
nand U3397 (N_3397,In_767,In_234);
nor U3398 (N_3398,In_319,In_816);
and U3399 (N_3399,In_857,In_874);
or U3400 (N_3400,In_171,In_161);
and U3401 (N_3401,In_302,In_544);
and U3402 (N_3402,In_543,In_492);
or U3403 (N_3403,In_101,In_842);
nor U3404 (N_3404,In_240,In_398);
nand U3405 (N_3405,In_418,In_690);
nand U3406 (N_3406,In_756,In_171);
and U3407 (N_3407,In_499,In_534);
and U3408 (N_3408,In_752,In_793);
or U3409 (N_3409,In_923,In_741);
nor U3410 (N_3410,In_390,In_731);
and U3411 (N_3411,In_179,In_307);
or U3412 (N_3412,In_661,In_602);
or U3413 (N_3413,In_555,In_622);
and U3414 (N_3414,In_664,In_615);
and U3415 (N_3415,In_381,In_367);
nor U3416 (N_3416,In_181,In_847);
nor U3417 (N_3417,In_730,In_33);
and U3418 (N_3418,In_888,In_294);
nor U3419 (N_3419,In_532,In_572);
and U3420 (N_3420,In_794,In_849);
nor U3421 (N_3421,In_118,In_83);
or U3422 (N_3422,In_724,In_445);
nand U3423 (N_3423,In_709,In_269);
and U3424 (N_3424,In_812,In_721);
and U3425 (N_3425,In_100,In_646);
or U3426 (N_3426,In_608,In_120);
nor U3427 (N_3427,In_406,In_67);
and U3428 (N_3428,In_866,In_114);
xnor U3429 (N_3429,In_925,In_85);
or U3430 (N_3430,In_392,In_27);
and U3431 (N_3431,In_968,In_174);
and U3432 (N_3432,In_990,In_105);
nor U3433 (N_3433,In_462,In_710);
or U3434 (N_3434,In_152,In_615);
nand U3435 (N_3435,In_551,In_26);
or U3436 (N_3436,In_210,In_927);
and U3437 (N_3437,In_82,In_434);
nand U3438 (N_3438,In_454,In_463);
or U3439 (N_3439,In_476,In_70);
and U3440 (N_3440,In_368,In_741);
nand U3441 (N_3441,In_48,In_272);
nand U3442 (N_3442,In_6,In_573);
nand U3443 (N_3443,In_161,In_969);
or U3444 (N_3444,In_427,In_307);
and U3445 (N_3445,In_816,In_49);
nor U3446 (N_3446,In_594,In_834);
nor U3447 (N_3447,In_104,In_965);
nor U3448 (N_3448,In_146,In_772);
nand U3449 (N_3449,In_643,In_484);
nor U3450 (N_3450,In_198,In_123);
and U3451 (N_3451,In_771,In_583);
or U3452 (N_3452,In_986,In_349);
nor U3453 (N_3453,In_869,In_457);
and U3454 (N_3454,In_145,In_193);
or U3455 (N_3455,In_326,In_91);
and U3456 (N_3456,In_949,In_687);
nand U3457 (N_3457,In_490,In_453);
nand U3458 (N_3458,In_903,In_156);
and U3459 (N_3459,In_380,In_356);
xnor U3460 (N_3460,In_19,In_246);
and U3461 (N_3461,In_517,In_551);
or U3462 (N_3462,In_712,In_802);
nand U3463 (N_3463,In_398,In_987);
nand U3464 (N_3464,In_534,In_640);
and U3465 (N_3465,In_516,In_573);
nor U3466 (N_3466,In_554,In_556);
nand U3467 (N_3467,In_969,In_897);
nor U3468 (N_3468,In_115,In_153);
or U3469 (N_3469,In_459,In_366);
or U3470 (N_3470,In_944,In_759);
nor U3471 (N_3471,In_965,In_110);
nor U3472 (N_3472,In_164,In_504);
or U3473 (N_3473,In_421,In_392);
or U3474 (N_3474,In_78,In_464);
and U3475 (N_3475,In_345,In_362);
and U3476 (N_3476,In_199,In_757);
nand U3477 (N_3477,In_680,In_939);
nand U3478 (N_3478,In_567,In_485);
or U3479 (N_3479,In_674,In_678);
or U3480 (N_3480,In_344,In_76);
nand U3481 (N_3481,In_614,In_416);
and U3482 (N_3482,In_656,In_100);
and U3483 (N_3483,In_900,In_467);
or U3484 (N_3484,In_331,In_51);
or U3485 (N_3485,In_736,In_899);
or U3486 (N_3486,In_626,In_121);
nor U3487 (N_3487,In_518,In_842);
or U3488 (N_3488,In_343,In_262);
and U3489 (N_3489,In_14,In_473);
and U3490 (N_3490,In_146,In_842);
nand U3491 (N_3491,In_988,In_233);
and U3492 (N_3492,In_836,In_417);
nor U3493 (N_3493,In_108,In_542);
xnor U3494 (N_3494,In_665,In_402);
or U3495 (N_3495,In_705,In_244);
and U3496 (N_3496,In_441,In_303);
nand U3497 (N_3497,In_226,In_944);
nor U3498 (N_3498,In_759,In_465);
or U3499 (N_3499,In_540,In_505);
nand U3500 (N_3500,In_258,In_794);
or U3501 (N_3501,In_935,In_243);
and U3502 (N_3502,In_730,In_121);
nand U3503 (N_3503,In_444,In_650);
nand U3504 (N_3504,In_650,In_740);
nor U3505 (N_3505,In_523,In_908);
nand U3506 (N_3506,In_877,In_721);
or U3507 (N_3507,In_732,In_101);
nor U3508 (N_3508,In_525,In_83);
nor U3509 (N_3509,In_54,In_92);
nand U3510 (N_3510,In_85,In_91);
nand U3511 (N_3511,In_219,In_267);
nand U3512 (N_3512,In_683,In_410);
nand U3513 (N_3513,In_267,In_358);
nor U3514 (N_3514,In_579,In_236);
nor U3515 (N_3515,In_62,In_686);
nand U3516 (N_3516,In_487,In_91);
nor U3517 (N_3517,In_225,In_492);
nand U3518 (N_3518,In_540,In_177);
nand U3519 (N_3519,In_583,In_147);
nand U3520 (N_3520,In_166,In_296);
xor U3521 (N_3521,In_592,In_199);
nand U3522 (N_3522,In_624,In_865);
and U3523 (N_3523,In_244,In_292);
and U3524 (N_3524,In_708,In_910);
nor U3525 (N_3525,In_282,In_818);
and U3526 (N_3526,In_671,In_336);
nor U3527 (N_3527,In_245,In_507);
and U3528 (N_3528,In_175,In_429);
nand U3529 (N_3529,In_102,In_56);
and U3530 (N_3530,In_906,In_175);
or U3531 (N_3531,In_977,In_796);
nor U3532 (N_3532,In_832,In_627);
nor U3533 (N_3533,In_757,In_666);
nor U3534 (N_3534,In_541,In_555);
or U3535 (N_3535,In_755,In_894);
and U3536 (N_3536,In_824,In_309);
nor U3537 (N_3537,In_313,In_3);
and U3538 (N_3538,In_132,In_966);
or U3539 (N_3539,In_845,In_830);
and U3540 (N_3540,In_432,In_282);
or U3541 (N_3541,In_306,In_477);
and U3542 (N_3542,In_528,In_63);
nand U3543 (N_3543,In_845,In_42);
or U3544 (N_3544,In_610,In_432);
nor U3545 (N_3545,In_624,In_949);
and U3546 (N_3546,In_111,In_617);
and U3547 (N_3547,In_655,In_930);
nor U3548 (N_3548,In_601,In_670);
or U3549 (N_3549,In_94,In_782);
or U3550 (N_3550,In_393,In_885);
or U3551 (N_3551,In_364,In_599);
nor U3552 (N_3552,In_267,In_972);
or U3553 (N_3553,In_969,In_888);
nand U3554 (N_3554,In_437,In_380);
or U3555 (N_3555,In_508,In_715);
nand U3556 (N_3556,In_341,In_709);
or U3557 (N_3557,In_80,In_167);
and U3558 (N_3558,In_631,In_108);
and U3559 (N_3559,In_2,In_657);
nor U3560 (N_3560,In_109,In_945);
and U3561 (N_3561,In_276,In_156);
nand U3562 (N_3562,In_543,In_701);
or U3563 (N_3563,In_723,In_313);
and U3564 (N_3564,In_838,In_477);
nor U3565 (N_3565,In_812,In_943);
or U3566 (N_3566,In_16,In_954);
and U3567 (N_3567,In_964,In_676);
and U3568 (N_3568,In_351,In_93);
or U3569 (N_3569,In_315,In_766);
nor U3570 (N_3570,In_975,In_430);
nor U3571 (N_3571,In_818,In_547);
nor U3572 (N_3572,In_981,In_542);
nand U3573 (N_3573,In_10,In_451);
and U3574 (N_3574,In_810,In_159);
nand U3575 (N_3575,In_323,In_656);
and U3576 (N_3576,In_217,In_122);
nand U3577 (N_3577,In_364,In_915);
nor U3578 (N_3578,In_412,In_947);
or U3579 (N_3579,In_801,In_674);
nor U3580 (N_3580,In_605,In_843);
and U3581 (N_3581,In_892,In_956);
or U3582 (N_3582,In_538,In_589);
and U3583 (N_3583,In_339,In_565);
and U3584 (N_3584,In_305,In_180);
nor U3585 (N_3585,In_896,In_951);
or U3586 (N_3586,In_318,In_813);
or U3587 (N_3587,In_522,In_205);
nor U3588 (N_3588,In_600,In_377);
nand U3589 (N_3589,In_617,In_304);
nor U3590 (N_3590,In_345,In_140);
nor U3591 (N_3591,In_72,In_118);
nand U3592 (N_3592,In_846,In_347);
nor U3593 (N_3593,In_537,In_746);
or U3594 (N_3594,In_529,In_101);
nor U3595 (N_3595,In_848,In_330);
and U3596 (N_3596,In_760,In_189);
nor U3597 (N_3597,In_28,In_5);
xor U3598 (N_3598,In_103,In_729);
or U3599 (N_3599,In_776,In_879);
and U3600 (N_3600,In_981,In_993);
or U3601 (N_3601,In_266,In_809);
nand U3602 (N_3602,In_517,In_80);
or U3603 (N_3603,In_639,In_516);
nand U3604 (N_3604,In_218,In_809);
nor U3605 (N_3605,In_505,In_797);
or U3606 (N_3606,In_609,In_974);
nor U3607 (N_3607,In_267,In_134);
and U3608 (N_3608,In_163,In_521);
and U3609 (N_3609,In_992,In_636);
and U3610 (N_3610,In_545,In_157);
or U3611 (N_3611,In_551,In_143);
or U3612 (N_3612,In_40,In_811);
and U3613 (N_3613,In_560,In_817);
and U3614 (N_3614,In_693,In_781);
and U3615 (N_3615,In_690,In_834);
or U3616 (N_3616,In_922,In_962);
and U3617 (N_3617,In_441,In_354);
or U3618 (N_3618,In_269,In_182);
and U3619 (N_3619,In_878,In_61);
nand U3620 (N_3620,In_204,In_648);
nor U3621 (N_3621,In_985,In_280);
and U3622 (N_3622,In_65,In_240);
or U3623 (N_3623,In_344,In_885);
nor U3624 (N_3624,In_259,In_960);
nor U3625 (N_3625,In_886,In_595);
or U3626 (N_3626,In_961,In_744);
or U3627 (N_3627,In_609,In_420);
or U3628 (N_3628,In_342,In_893);
and U3629 (N_3629,In_809,In_747);
and U3630 (N_3630,In_837,In_737);
nor U3631 (N_3631,In_634,In_334);
nor U3632 (N_3632,In_920,In_407);
and U3633 (N_3633,In_919,In_616);
nand U3634 (N_3634,In_374,In_253);
nand U3635 (N_3635,In_773,In_197);
nand U3636 (N_3636,In_947,In_956);
nor U3637 (N_3637,In_610,In_950);
nand U3638 (N_3638,In_259,In_813);
and U3639 (N_3639,In_132,In_351);
nor U3640 (N_3640,In_969,In_773);
and U3641 (N_3641,In_254,In_837);
nand U3642 (N_3642,In_692,In_455);
and U3643 (N_3643,In_573,In_275);
or U3644 (N_3644,In_262,In_916);
or U3645 (N_3645,In_714,In_540);
or U3646 (N_3646,In_528,In_998);
nand U3647 (N_3647,In_813,In_6);
nor U3648 (N_3648,In_905,In_78);
or U3649 (N_3649,In_990,In_393);
nor U3650 (N_3650,In_67,In_293);
nor U3651 (N_3651,In_838,In_226);
nor U3652 (N_3652,In_83,In_527);
nor U3653 (N_3653,In_739,In_871);
and U3654 (N_3654,In_175,In_267);
or U3655 (N_3655,In_935,In_555);
nand U3656 (N_3656,In_872,In_700);
or U3657 (N_3657,In_319,In_476);
nand U3658 (N_3658,In_650,In_445);
nor U3659 (N_3659,In_927,In_672);
and U3660 (N_3660,In_427,In_252);
nor U3661 (N_3661,In_968,In_504);
and U3662 (N_3662,In_450,In_252);
nor U3663 (N_3663,In_922,In_437);
and U3664 (N_3664,In_999,In_434);
nand U3665 (N_3665,In_173,In_272);
and U3666 (N_3666,In_932,In_362);
and U3667 (N_3667,In_408,In_505);
and U3668 (N_3668,In_574,In_193);
nand U3669 (N_3669,In_19,In_654);
and U3670 (N_3670,In_681,In_15);
and U3671 (N_3671,In_673,In_504);
nor U3672 (N_3672,In_928,In_738);
or U3673 (N_3673,In_856,In_581);
or U3674 (N_3674,In_86,In_645);
nor U3675 (N_3675,In_341,In_979);
nand U3676 (N_3676,In_124,In_711);
nand U3677 (N_3677,In_548,In_923);
nand U3678 (N_3678,In_537,In_669);
and U3679 (N_3679,In_235,In_617);
or U3680 (N_3680,In_321,In_672);
or U3681 (N_3681,In_246,In_127);
nor U3682 (N_3682,In_138,In_320);
nand U3683 (N_3683,In_714,In_562);
or U3684 (N_3684,In_387,In_757);
nor U3685 (N_3685,In_640,In_529);
nand U3686 (N_3686,In_12,In_370);
or U3687 (N_3687,In_973,In_819);
or U3688 (N_3688,In_943,In_191);
nor U3689 (N_3689,In_554,In_593);
nand U3690 (N_3690,In_622,In_420);
nand U3691 (N_3691,In_178,In_44);
nor U3692 (N_3692,In_209,In_912);
nand U3693 (N_3693,In_330,In_233);
or U3694 (N_3694,In_925,In_657);
nand U3695 (N_3695,In_972,In_226);
nand U3696 (N_3696,In_753,In_931);
nor U3697 (N_3697,In_250,In_993);
nor U3698 (N_3698,In_999,In_493);
and U3699 (N_3699,In_578,In_783);
nand U3700 (N_3700,In_691,In_982);
and U3701 (N_3701,In_529,In_82);
and U3702 (N_3702,In_360,In_744);
and U3703 (N_3703,In_242,In_293);
and U3704 (N_3704,In_634,In_722);
nor U3705 (N_3705,In_590,In_591);
and U3706 (N_3706,In_475,In_310);
and U3707 (N_3707,In_965,In_162);
and U3708 (N_3708,In_228,In_206);
or U3709 (N_3709,In_889,In_81);
or U3710 (N_3710,In_145,In_420);
or U3711 (N_3711,In_857,In_625);
or U3712 (N_3712,In_973,In_984);
and U3713 (N_3713,In_591,In_155);
nand U3714 (N_3714,In_464,In_488);
and U3715 (N_3715,In_654,In_778);
and U3716 (N_3716,In_236,In_988);
and U3717 (N_3717,In_48,In_807);
and U3718 (N_3718,In_203,In_613);
or U3719 (N_3719,In_757,In_152);
nand U3720 (N_3720,In_803,In_257);
and U3721 (N_3721,In_975,In_329);
and U3722 (N_3722,In_381,In_440);
nor U3723 (N_3723,In_961,In_332);
or U3724 (N_3724,In_73,In_736);
xnor U3725 (N_3725,In_276,In_308);
nor U3726 (N_3726,In_607,In_408);
nor U3727 (N_3727,In_994,In_457);
or U3728 (N_3728,In_832,In_206);
and U3729 (N_3729,In_677,In_363);
and U3730 (N_3730,In_870,In_711);
or U3731 (N_3731,In_297,In_337);
or U3732 (N_3732,In_647,In_240);
and U3733 (N_3733,In_697,In_975);
nand U3734 (N_3734,In_918,In_277);
or U3735 (N_3735,In_959,In_172);
nand U3736 (N_3736,In_150,In_472);
nand U3737 (N_3737,In_394,In_486);
nor U3738 (N_3738,In_58,In_18);
nand U3739 (N_3739,In_470,In_347);
or U3740 (N_3740,In_474,In_995);
nor U3741 (N_3741,In_191,In_42);
nand U3742 (N_3742,In_541,In_361);
and U3743 (N_3743,In_482,In_41);
nand U3744 (N_3744,In_44,In_715);
or U3745 (N_3745,In_349,In_170);
nand U3746 (N_3746,In_332,In_512);
or U3747 (N_3747,In_242,In_921);
nor U3748 (N_3748,In_789,In_958);
nand U3749 (N_3749,In_310,In_939);
and U3750 (N_3750,In_258,In_496);
nor U3751 (N_3751,In_414,In_212);
nor U3752 (N_3752,In_155,In_603);
and U3753 (N_3753,In_429,In_310);
nor U3754 (N_3754,In_891,In_80);
or U3755 (N_3755,In_298,In_403);
nor U3756 (N_3756,In_384,In_142);
nand U3757 (N_3757,In_787,In_521);
and U3758 (N_3758,In_164,In_935);
and U3759 (N_3759,In_6,In_905);
and U3760 (N_3760,In_983,In_566);
and U3761 (N_3761,In_551,In_986);
nor U3762 (N_3762,In_550,In_655);
or U3763 (N_3763,In_751,In_410);
nor U3764 (N_3764,In_655,In_21);
nor U3765 (N_3765,In_422,In_931);
nor U3766 (N_3766,In_923,In_219);
nand U3767 (N_3767,In_875,In_982);
nand U3768 (N_3768,In_804,In_520);
xnor U3769 (N_3769,In_435,In_673);
nor U3770 (N_3770,In_391,In_634);
nand U3771 (N_3771,In_581,In_678);
nand U3772 (N_3772,In_292,In_62);
nor U3773 (N_3773,In_794,In_928);
nor U3774 (N_3774,In_914,In_694);
nand U3775 (N_3775,In_711,In_251);
or U3776 (N_3776,In_660,In_271);
nand U3777 (N_3777,In_935,In_358);
nand U3778 (N_3778,In_353,In_131);
or U3779 (N_3779,In_69,In_734);
or U3780 (N_3780,In_19,In_350);
nor U3781 (N_3781,In_896,In_398);
nor U3782 (N_3782,In_656,In_531);
and U3783 (N_3783,In_738,In_831);
nor U3784 (N_3784,In_675,In_312);
nand U3785 (N_3785,In_760,In_55);
or U3786 (N_3786,In_608,In_385);
nor U3787 (N_3787,In_682,In_365);
nor U3788 (N_3788,In_970,In_778);
nor U3789 (N_3789,In_413,In_328);
or U3790 (N_3790,In_189,In_371);
nor U3791 (N_3791,In_755,In_233);
nand U3792 (N_3792,In_50,In_719);
or U3793 (N_3793,In_334,In_381);
and U3794 (N_3794,In_706,In_496);
nand U3795 (N_3795,In_478,In_901);
and U3796 (N_3796,In_368,In_105);
or U3797 (N_3797,In_124,In_232);
nor U3798 (N_3798,In_328,In_683);
and U3799 (N_3799,In_175,In_39);
or U3800 (N_3800,In_402,In_53);
nand U3801 (N_3801,In_850,In_466);
nor U3802 (N_3802,In_46,In_738);
or U3803 (N_3803,In_653,In_418);
or U3804 (N_3804,In_862,In_301);
or U3805 (N_3805,In_720,In_254);
nand U3806 (N_3806,In_976,In_356);
or U3807 (N_3807,In_714,In_528);
nor U3808 (N_3808,In_621,In_124);
nor U3809 (N_3809,In_561,In_459);
nand U3810 (N_3810,In_948,In_555);
nand U3811 (N_3811,In_610,In_584);
and U3812 (N_3812,In_374,In_991);
or U3813 (N_3813,In_190,In_293);
nor U3814 (N_3814,In_647,In_397);
nand U3815 (N_3815,In_619,In_135);
and U3816 (N_3816,In_72,In_96);
nor U3817 (N_3817,In_232,In_87);
and U3818 (N_3818,In_544,In_310);
nor U3819 (N_3819,In_436,In_233);
or U3820 (N_3820,In_150,In_60);
and U3821 (N_3821,In_335,In_862);
nand U3822 (N_3822,In_180,In_732);
and U3823 (N_3823,In_516,In_9);
and U3824 (N_3824,In_618,In_716);
and U3825 (N_3825,In_807,In_872);
and U3826 (N_3826,In_264,In_792);
nor U3827 (N_3827,In_38,In_942);
or U3828 (N_3828,In_391,In_338);
and U3829 (N_3829,In_348,In_268);
or U3830 (N_3830,In_425,In_300);
nand U3831 (N_3831,In_379,In_351);
nand U3832 (N_3832,In_551,In_513);
nor U3833 (N_3833,In_881,In_414);
and U3834 (N_3834,In_95,In_322);
nand U3835 (N_3835,In_904,In_838);
and U3836 (N_3836,In_830,In_128);
and U3837 (N_3837,In_573,In_684);
or U3838 (N_3838,In_150,In_36);
nor U3839 (N_3839,In_758,In_540);
nor U3840 (N_3840,In_228,In_938);
nand U3841 (N_3841,In_467,In_806);
and U3842 (N_3842,In_138,In_20);
nand U3843 (N_3843,In_947,In_522);
xor U3844 (N_3844,In_528,In_409);
nand U3845 (N_3845,In_479,In_988);
nor U3846 (N_3846,In_146,In_636);
and U3847 (N_3847,In_312,In_139);
or U3848 (N_3848,In_15,In_669);
or U3849 (N_3849,In_374,In_497);
nor U3850 (N_3850,In_545,In_934);
and U3851 (N_3851,In_48,In_168);
and U3852 (N_3852,In_385,In_247);
nand U3853 (N_3853,In_951,In_771);
nor U3854 (N_3854,In_914,In_630);
nor U3855 (N_3855,In_441,In_991);
nand U3856 (N_3856,In_734,In_723);
and U3857 (N_3857,In_353,In_569);
and U3858 (N_3858,In_479,In_686);
or U3859 (N_3859,In_439,In_293);
or U3860 (N_3860,In_8,In_64);
nand U3861 (N_3861,In_919,In_611);
nand U3862 (N_3862,In_291,In_139);
nor U3863 (N_3863,In_406,In_669);
or U3864 (N_3864,In_360,In_546);
nor U3865 (N_3865,In_28,In_118);
and U3866 (N_3866,In_920,In_163);
or U3867 (N_3867,In_228,In_976);
nor U3868 (N_3868,In_934,In_853);
and U3869 (N_3869,In_463,In_402);
nand U3870 (N_3870,In_318,In_536);
or U3871 (N_3871,In_489,In_714);
nand U3872 (N_3872,In_240,In_71);
or U3873 (N_3873,In_585,In_101);
and U3874 (N_3874,In_762,In_371);
and U3875 (N_3875,In_427,In_26);
and U3876 (N_3876,In_862,In_646);
or U3877 (N_3877,In_267,In_872);
and U3878 (N_3878,In_789,In_338);
or U3879 (N_3879,In_722,In_972);
nand U3880 (N_3880,In_750,In_436);
nand U3881 (N_3881,In_200,In_214);
nor U3882 (N_3882,In_281,In_936);
or U3883 (N_3883,In_830,In_702);
nor U3884 (N_3884,In_861,In_796);
and U3885 (N_3885,In_359,In_567);
nand U3886 (N_3886,In_297,In_845);
and U3887 (N_3887,In_917,In_544);
and U3888 (N_3888,In_15,In_374);
nor U3889 (N_3889,In_94,In_709);
or U3890 (N_3890,In_748,In_625);
nand U3891 (N_3891,In_513,In_715);
nand U3892 (N_3892,In_713,In_89);
nand U3893 (N_3893,In_278,In_869);
nor U3894 (N_3894,In_339,In_25);
or U3895 (N_3895,In_627,In_582);
and U3896 (N_3896,In_896,In_737);
or U3897 (N_3897,In_373,In_623);
nor U3898 (N_3898,In_622,In_314);
nor U3899 (N_3899,In_153,In_3);
and U3900 (N_3900,In_144,In_53);
nand U3901 (N_3901,In_461,In_650);
and U3902 (N_3902,In_401,In_247);
nor U3903 (N_3903,In_436,In_262);
nand U3904 (N_3904,In_683,In_807);
or U3905 (N_3905,In_185,In_698);
nor U3906 (N_3906,In_762,In_564);
nand U3907 (N_3907,In_358,In_707);
nor U3908 (N_3908,In_549,In_600);
nand U3909 (N_3909,In_971,In_372);
nand U3910 (N_3910,In_429,In_802);
nor U3911 (N_3911,In_85,In_4);
nand U3912 (N_3912,In_458,In_669);
or U3913 (N_3913,In_124,In_772);
xor U3914 (N_3914,In_279,In_288);
nor U3915 (N_3915,In_664,In_771);
or U3916 (N_3916,In_178,In_746);
nor U3917 (N_3917,In_879,In_939);
and U3918 (N_3918,In_284,In_540);
nand U3919 (N_3919,In_476,In_128);
xnor U3920 (N_3920,In_343,In_254);
and U3921 (N_3921,In_530,In_747);
nor U3922 (N_3922,In_307,In_143);
nand U3923 (N_3923,In_243,In_730);
nor U3924 (N_3924,In_973,In_903);
nand U3925 (N_3925,In_376,In_151);
nand U3926 (N_3926,In_885,In_984);
or U3927 (N_3927,In_301,In_657);
and U3928 (N_3928,In_336,In_404);
and U3929 (N_3929,In_84,In_569);
xnor U3930 (N_3930,In_679,In_762);
nand U3931 (N_3931,In_920,In_78);
nor U3932 (N_3932,In_723,In_320);
nand U3933 (N_3933,In_408,In_242);
nand U3934 (N_3934,In_880,In_513);
nor U3935 (N_3935,In_458,In_482);
nand U3936 (N_3936,In_282,In_639);
nor U3937 (N_3937,In_105,In_428);
nor U3938 (N_3938,In_470,In_784);
or U3939 (N_3939,In_956,In_815);
or U3940 (N_3940,In_531,In_116);
nand U3941 (N_3941,In_451,In_325);
or U3942 (N_3942,In_988,In_725);
and U3943 (N_3943,In_280,In_604);
nor U3944 (N_3944,In_951,In_365);
or U3945 (N_3945,In_199,In_716);
and U3946 (N_3946,In_501,In_965);
nand U3947 (N_3947,In_648,In_545);
and U3948 (N_3948,In_717,In_718);
or U3949 (N_3949,In_267,In_228);
nor U3950 (N_3950,In_556,In_906);
or U3951 (N_3951,In_162,In_810);
nand U3952 (N_3952,In_898,In_830);
nor U3953 (N_3953,In_321,In_891);
or U3954 (N_3954,In_508,In_472);
and U3955 (N_3955,In_899,In_7);
nor U3956 (N_3956,In_616,In_892);
or U3957 (N_3957,In_857,In_939);
and U3958 (N_3958,In_563,In_917);
nor U3959 (N_3959,In_230,In_331);
and U3960 (N_3960,In_77,In_334);
nand U3961 (N_3961,In_672,In_314);
and U3962 (N_3962,In_941,In_37);
or U3963 (N_3963,In_373,In_379);
and U3964 (N_3964,In_490,In_695);
nor U3965 (N_3965,In_283,In_815);
nor U3966 (N_3966,In_898,In_395);
or U3967 (N_3967,In_28,In_566);
nand U3968 (N_3968,In_507,In_596);
nand U3969 (N_3969,In_17,In_529);
or U3970 (N_3970,In_915,In_134);
or U3971 (N_3971,In_790,In_670);
or U3972 (N_3972,In_460,In_889);
or U3973 (N_3973,In_664,In_969);
or U3974 (N_3974,In_490,In_622);
and U3975 (N_3975,In_588,In_492);
and U3976 (N_3976,In_246,In_15);
nor U3977 (N_3977,In_598,In_822);
nor U3978 (N_3978,In_500,In_657);
or U3979 (N_3979,In_121,In_228);
nor U3980 (N_3980,In_157,In_768);
nand U3981 (N_3981,In_147,In_979);
nand U3982 (N_3982,In_986,In_148);
or U3983 (N_3983,In_206,In_761);
nor U3984 (N_3984,In_981,In_950);
nand U3985 (N_3985,In_102,In_907);
or U3986 (N_3986,In_467,In_70);
nand U3987 (N_3987,In_221,In_441);
or U3988 (N_3988,In_309,In_838);
and U3989 (N_3989,In_612,In_328);
nand U3990 (N_3990,In_615,In_26);
nand U3991 (N_3991,In_663,In_155);
nor U3992 (N_3992,In_759,In_763);
or U3993 (N_3993,In_124,In_814);
nor U3994 (N_3994,In_414,In_522);
nor U3995 (N_3995,In_774,In_415);
and U3996 (N_3996,In_717,In_271);
nor U3997 (N_3997,In_118,In_757);
nand U3998 (N_3998,In_176,In_472);
or U3999 (N_3999,In_345,In_779);
or U4000 (N_4000,In_164,In_295);
or U4001 (N_4001,In_715,In_833);
or U4002 (N_4002,In_258,In_77);
and U4003 (N_4003,In_507,In_411);
nor U4004 (N_4004,In_608,In_503);
nor U4005 (N_4005,In_957,In_492);
nand U4006 (N_4006,In_941,In_410);
nor U4007 (N_4007,In_426,In_684);
and U4008 (N_4008,In_303,In_260);
nand U4009 (N_4009,In_963,In_279);
nor U4010 (N_4010,In_778,In_721);
nand U4011 (N_4011,In_5,In_605);
or U4012 (N_4012,In_602,In_752);
and U4013 (N_4013,In_847,In_127);
and U4014 (N_4014,In_800,In_535);
nor U4015 (N_4015,In_614,In_94);
nor U4016 (N_4016,In_224,In_850);
nand U4017 (N_4017,In_444,In_138);
nand U4018 (N_4018,In_39,In_167);
and U4019 (N_4019,In_228,In_965);
and U4020 (N_4020,In_220,In_397);
nand U4021 (N_4021,In_990,In_632);
nand U4022 (N_4022,In_750,In_248);
nand U4023 (N_4023,In_629,In_267);
and U4024 (N_4024,In_798,In_339);
nor U4025 (N_4025,In_608,In_448);
nor U4026 (N_4026,In_575,In_801);
and U4027 (N_4027,In_36,In_268);
and U4028 (N_4028,In_801,In_510);
and U4029 (N_4029,In_503,In_124);
nand U4030 (N_4030,In_327,In_497);
nand U4031 (N_4031,In_211,In_263);
and U4032 (N_4032,In_55,In_651);
nand U4033 (N_4033,In_918,In_307);
nand U4034 (N_4034,In_870,In_753);
xnor U4035 (N_4035,In_95,In_904);
nand U4036 (N_4036,In_721,In_440);
and U4037 (N_4037,In_883,In_253);
nor U4038 (N_4038,In_507,In_992);
nand U4039 (N_4039,In_188,In_381);
and U4040 (N_4040,In_108,In_623);
nor U4041 (N_4041,In_125,In_968);
nor U4042 (N_4042,In_11,In_336);
nand U4043 (N_4043,In_988,In_976);
nand U4044 (N_4044,In_248,In_325);
and U4045 (N_4045,In_845,In_507);
nor U4046 (N_4046,In_858,In_971);
nand U4047 (N_4047,In_496,In_767);
or U4048 (N_4048,In_335,In_992);
nand U4049 (N_4049,In_386,In_958);
nor U4050 (N_4050,In_342,In_250);
or U4051 (N_4051,In_936,In_13);
or U4052 (N_4052,In_714,In_514);
or U4053 (N_4053,In_853,In_111);
and U4054 (N_4054,In_466,In_631);
and U4055 (N_4055,In_367,In_68);
and U4056 (N_4056,In_609,In_744);
and U4057 (N_4057,In_810,In_857);
or U4058 (N_4058,In_39,In_828);
and U4059 (N_4059,In_499,In_373);
nor U4060 (N_4060,In_990,In_159);
and U4061 (N_4061,In_518,In_949);
nor U4062 (N_4062,In_300,In_9);
and U4063 (N_4063,In_32,In_387);
nand U4064 (N_4064,In_723,In_765);
nor U4065 (N_4065,In_425,In_356);
and U4066 (N_4066,In_965,In_419);
and U4067 (N_4067,In_766,In_233);
or U4068 (N_4068,In_42,In_244);
nor U4069 (N_4069,In_525,In_491);
nand U4070 (N_4070,In_496,In_222);
nand U4071 (N_4071,In_784,In_487);
nand U4072 (N_4072,In_896,In_823);
nand U4073 (N_4073,In_710,In_449);
nor U4074 (N_4074,In_714,In_488);
nand U4075 (N_4075,In_355,In_215);
and U4076 (N_4076,In_694,In_757);
nor U4077 (N_4077,In_904,In_420);
nor U4078 (N_4078,In_329,In_481);
nand U4079 (N_4079,In_274,In_916);
and U4080 (N_4080,In_418,In_93);
or U4081 (N_4081,In_628,In_239);
nor U4082 (N_4082,In_888,In_387);
and U4083 (N_4083,In_551,In_159);
or U4084 (N_4084,In_838,In_10);
and U4085 (N_4085,In_173,In_398);
nor U4086 (N_4086,In_287,In_277);
or U4087 (N_4087,In_686,In_202);
and U4088 (N_4088,In_57,In_375);
nand U4089 (N_4089,In_413,In_155);
nand U4090 (N_4090,In_793,In_858);
nor U4091 (N_4091,In_803,In_305);
nor U4092 (N_4092,In_318,In_127);
nor U4093 (N_4093,In_786,In_310);
and U4094 (N_4094,In_974,In_866);
nand U4095 (N_4095,In_448,In_408);
and U4096 (N_4096,In_235,In_125);
and U4097 (N_4097,In_717,In_835);
nand U4098 (N_4098,In_338,In_704);
or U4099 (N_4099,In_605,In_100);
nor U4100 (N_4100,In_499,In_699);
and U4101 (N_4101,In_790,In_39);
or U4102 (N_4102,In_674,In_318);
and U4103 (N_4103,In_209,In_801);
and U4104 (N_4104,In_623,In_688);
and U4105 (N_4105,In_672,In_886);
nand U4106 (N_4106,In_286,In_456);
nand U4107 (N_4107,In_697,In_343);
nor U4108 (N_4108,In_711,In_297);
and U4109 (N_4109,In_659,In_983);
and U4110 (N_4110,In_542,In_578);
or U4111 (N_4111,In_813,In_681);
and U4112 (N_4112,In_71,In_197);
and U4113 (N_4113,In_592,In_918);
and U4114 (N_4114,In_475,In_501);
and U4115 (N_4115,In_948,In_364);
xnor U4116 (N_4116,In_757,In_334);
nand U4117 (N_4117,In_630,In_142);
and U4118 (N_4118,In_116,In_332);
nor U4119 (N_4119,In_870,In_847);
nand U4120 (N_4120,In_814,In_675);
or U4121 (N_4121,In_947,In_618);
nor U4122 (N_4122,In_582,In_770);
and U4123 (N_4123,In_237,In_492);
or U4124 (N_4124,In_191,In_86);
or U4125 (N_4125,In_221,In_579);
nor U4126 (N_4126,In_663,In_406);
and U4127 (N_4127,In_887,In_663);
nor U4128 (N_4128,In_468,In_826);
or U4129 (N_4129,In_337,In_98);
and U4130 (N_4130,In_110,In_386);
or U4131 (N_4131,In_331,In_377);
nand U4132 (N_4132,In_362,In_156);
or U4133 (N_4133,In_370,In_555);
or U4134 (N_4134,In_850,In_672);
and U4135 (N_4135,In_147,In_505);
or U4136 (N_4136,In_940,In_292);
nand U4137 (N_4137,In_137,In_66);
nand U4138 (N_4138,In_581,In_264);
and U4139 (N_4139,In_2,In_610);
or U4140 (N_4140,In_814,In_614);
nor U4141 (N_4141,In_788,In_496);
nand U4142 (N_4142,In_379,In_769);
and U4143 (N_4143,In_318,In_625);
xnor U4144 (N_4144,In_380,In_608);
and U4145 (N_4145,In_153,In_406);
and U4146 (N_4146,In_326,In_150);
or U4147 (N_4147,In_308,In_972);
or U4148 (N_4148,In_138,In_821);
nor U4149 (N_4149,In_870,In_519);
or U4150 (N_4150,In_650,In_994);
nand U4151 (N_4151,In_286,In_318);
nand U4152 (N_4152,In_75,In_797);
nor U4153 (N_4153,In_650,In_674);
and U4154 (N_4154,In_664,In_708);
or U4155 (N_4155,In_386,In_263);
or U4156 (N_4156,In_912,In_59);
and U4157 (N_4157,In_459,In_867);
nand U4158 (N_4158,In_520,In_435);
nor U4159 (N_4159,In_950,In_944);
or U4160 (N_4160,In_649,In_498);
nand U4161 (N_4161,In_48,In_289);
nand U4162 (N_4162,In_676,In_324);
nor U4163 (N_4163,In_350,In_732);
nor U4164 (N_4164,In_768,In_910);
or U4165 (N_4165,In_391,In_935);
nand U4166 (N_4166,In_498,In_954);
nand U4167 (N_4167,In_617,In_758);
nor U4168 (N_4168,In_292,In_139);
or U4169 (N_4169,In_919,In_55);
and U4170 (N_4170,In_832,In_998);
nand U4171 (N_4171,In_762,In_819);
and U4172 (N_4172,In_783,In_561);
nor U4173 (N_4173,In_85,In_805);
nor U4174 (N_4174,In_995,In_397);
nand U4175 (N_4175,In_982,In_851);
nor U4176 (N_4176,In_285,In_802);
nand U4177 (N_4177,In_336,In_378);
nand U4178 (N_4178,In_730,In_382);
or U4179 (N_4179,In_1,In_200);
nor U4180 (N_4180,In_235,In_120);
nand U4181 (N_4181,In_562,In_614);
nor U4182 (N_4182,In_357,In_884);
or U4183 (N_4183,In_175,In_316);
nor U4184 (N_4184,In_910,In_853);
nor U4185 (N_4185,In_66,In_697);
or U4186 (N_4186,In_897,In_306);
nor U4187 (N_4187,In_144,In_429);
or U4188 (N_4188,In_633,In_545);
or U4189 (N_4189,In_251,In_202);
or U4190 (N_4190,In_564,In_870);
nor U4191 (N_4191,In_15,In_678);
nor U4192 (N_4192,In_930,In_296);
or U4193 (N_4193,In_595,In_836);
nor U4194 (N_4194,In_435,In_881);
nor U4195 (N_4195,In_943,In_447);
nand U4196 (N_4196,In_228,In_218);
nand U4197 (N_4197,In_36,In_999);
or U4198 (N_4198,In_912,In_685);
or U4199 (N_4199,In_835,In_65);
nand U4200 (N_4200,In_458,In_388);
or U4201 (N_4201,In_549,In_612);
nand U4202 (N_4202,In_577,In_529);
nand U4203 (N_4203,In_546,In_167);
and U4204 (N_4204,In_655,In_754);
and U4205 (N_4205,In_406,In_34);
and U4206 (N_4206,In_568,In_635);
and U4207 (N_4207,In_650,In_727);
nor U4208 (N_4208,In_985,In_957);
and U4209 (N_4209,In_873,In_987);
nand U4210 (N_4210,In_978,In_781);
nor U4211 (N_4211,In_392,In_14);
nor U4212 (N_4212,In_84,In_606);
and U4213 (N_4213,In_233,In_632);
or U4214 (N_4214,In_295,In_98);
and U4215 (N_4215,In_871,In_221);
nand U4216 (N_4216,In_827,In_615);
nor U4217 (N_4217,In_816,In_694);
nand U4218 (N_4218,In_982,In_714);
nand U4219 (N_4219,In_424,In_542);
and U4220 (N_4220,In_144,In_393);
and U4221 (N_4221,In_9,In_258);
and U4222 (N_4222,In_285,In_974);
nor U4223 (N_4223,In_883,In_877);
nor U4224 (N_4224,In_895,In_732);
or U4225 (N_4225,In_356,In_652);
nand U4226 (N_4226,In_525,In_580);
nand U4227 (N_4227,In_932,In_973);
nor U4228 (N_4228,In_436,In_264);
and U4229 (N_4229,In_896,In_109);
nand U4230 (N_4230,In_899,In_508);
and U4231 (N_4231,In_169,In_38);
nand U4232 (N_4232,In_635,In_951);
nand U4233 (N_4233,In_428,In_616);
and U4234 (N_4234,In_495,In_689);
and U4235 (N_4235,In_810,In_210);
nor U4236 (N_4236,In_665,In_912);
nor U4237 (N_4237,In_852,In_715);
or U4238 (N_4238,In_219,In_228);
and U4239 (N_4239,In_454,In_188);
nor U4240 (N_4240,In_749,In_666);
nand U4241 (N_4241,In_463,In_502);
and U4242 (N_4242,In_897,In_25);
nor U4243 (N_4243,In_697,In_31);
nand U4244 (N_4244,In_428,In_597);
and U4245 (N_4245,In_303,In_866);
and U4246 (N_4246,In_972,In_604);
nand U4247 (N_4247,In_599,In_685);
nand U4248 (N_4248,In_248,In_856);
and U4249 (N_4249,In_387,In_751);
nand U4250 (N_4250,In_715,In_935);
nand U4251 (N_4251,In_839,In_789);
nand U4252 (N_4252,In_261,In_728);
nor U4253 (N_4253,In_69,In_752);
and U4254 (N_4254,In_251,In_146);
or U4255 (N_4255,In_582,In_86);
and U4256 (N_4256,In_210,In_73);
or U4257 (N_4257,In_108,In_647);
nand U4258 (N_4258,In_246,In_417);
or U4259 (N_4259,In_915,In_66);
nand U4260 (N_4260,In_503,In_153);
nor U4261 (N_4261,In_590,In_939);
nand U4262 (N_4262,In_214,In_362);
and U4263 (N_4263,In_706,In_304);
and U4264 (N_4264,In_255,In_224);
or U4265 (N_4265,In_76,In_747);
nor U4266 (N_4266,In_576,In_982);
nand U4267 (N_4267,In_784,In_941);
nor U4268 (N_4268,In_469,In_576);
nor U4269 (N_4269,In_247,In_993);
and U4270 (N_4270,In_789,In_795);
nand U4271 (N_4271,In_842,In_837);
nor U4272 (N_4272,In_346,In_178);
nor U4273 (N_4273,In_974,In_820);
and U4274 (N_4274,In_808,In_192);
nand U4275 (N_4275,In_331,In_279);
and U4276 (N_4276,In_459,In_383);
nand U4277 (N_4277,In_900,In_55);
nand U4278 (N_4278,In_245,In_101);
nor U4279 (N_4279,In_914,In_801);
or U4280 (N_4280,In_869,In_332);
nand U4281 (N_4281,In_932,In_915);
nor U4282 (N_4282,In_504,In_502);
nor U4283 (N_4283,In_70,In_28);
nor U4284 (N_4284,In_227,In_648);
nand U4285 (N_4285,In_488,In_737);
xor U4286 (N_4286,In_975,In_613);
nor U4287 (N_4287,In_424,In_168);
nand U4288 (N_4288,In_470,In_706);
nand U4289 (N_4289,In_883,In_513);
nor U4290 (N_4290,In_411,In_472);
nor U4291 (N_4291,In_799,In_954);
nand U4292 (N_4292,In_899,In_534);
nand U4293 (N_4293,In_942,In_921);
and U4294 (N_4294,In_490,In_8);
nor U4295 (N_4295,In_318,In_436);
or U4296 (N_4296,In_419,In_216);
nor U4297 (N_4297,In_162,In_952);
nand U4298 (N_4298,In_150,In_542);
and U4299 (N_4299,In_765,In_754);
and U4300 (N_4300,In_797,In_618);
or U4301 (N_4301,In_290,In_992);
or U4302 (N_4302,In_199,In_93);
and U4303 (N_4303,In_658,In_876);
nor U4304 (N_4304,In_692,In_201);
nor U4305 (N_4305,In_877,In_382);
or U4306 (N_4306,In_690,In_228);
or U4307 (N_4307,In_414,In_683);
or U4308 (N_4308,In_173,In_391);
or U4309 (N_4309,In_465,In_585);
and U4310 (N_4310,In_469,In_192);
nor U4311 (N_4311,In_858,In_888);
and U4312 (N_4312,In_215,In_446);
nand U4313 (N_4313,In_886,In_288);
and U4314 (N_4314,In_100,In_365);
nand U4315 (N_4315,In_232,In_591);
or U4316 (N_4316,In_616,In_958);
nand U4317 (N_4317,In_432,In_182);
nand U4318 (N_4318,In_999,In_534);
nor U4319 (N_4319,In_961,In_977);
nor U4320 (N_4320,In_378,In_581);
or U4321 (N_4321,In_392,In_783);
or U4322 (N_4322,In_411,In_803);
and U4323 (N_4323,In_10,In_492);
and U4324 (N_4324,In_494,In_208);
nor U4325 (N_4325,In_487,In_204);
nand U4326 (N_4326,In_50,In_718);
and U4327 (N_4327,In_794,In_982);
or U4328 (N_4328,In_623,In_974);
nor U4329 (N_4329,In_555,In_479);
nand U4330 (N_4330,In_576,In_205);
xnor U4331 (N_4331,In_442,In_930);
nor U4332 (N_4332,In_579,In_691);
nand U4333 (N_4333,In_218,In_178);
nand U4334 (N_4334,In_149,In_276);
or U4335 (N_4335,In_50,In_81);
nand U4336 (N_4336,In_838,In_63);
nor U4337 (N_4337,In_800,In_426);
or U4338 (N_4338,In_351,In_848);
nand U4339 (N_4339,In_625,In_528);
or U4340 (N_4340,In_586,In_889);
nand U4341 (N_4341,In_958,In_662);
or U4342 (N_4342,In_333,In_705);
and U4343 (N_4343,In_425,In_458);
nor U4344 (N_4344,In_789,In_275);
nand U4345 (N_4345,In_155,In_629);
and U4346 (N_4346,In_520,In_16);
nor U4347 (N_4347,In_946,In_700);
or U4348 (N_4348,In_366,In_132);
and U4349 (N_4349,In_913,In_123);
or U4350 (N_4350,In_676,In_699);
and U4351 (N_4351,In_423,In_531);
nand U4352 (N_4352,In_49,In_721);
or U4353 (N_4353,In_359,In_850);
nand U4354 (N_4354,In_522,In_690);
and U4355 (N_4355,In_185,In_156);
nand U4356 (N_4356,In_998,In_886);
and U4357 (N_4357,In_511,In_498);
nor U4358 (N_4358,In_740,In_4);
nor U4359 (N_4359,In_83,In_744);
and U4360 (N_4360,In_783,In_492);
nor U4361 (N_4361,In_475,In_133);
nand U4362 (N_4362,In_872,In_702);
or U4363 (N_4363,In_969,In_412);
nor U4364 (N_4364,In_401,In_547);
nor U4365 (N_4365,In_820,In_817);
nor U4366 (N_4366,In_296,In_856);
and U4367 (N_4367,In_78,In_42);
or U4368 (N_4368,In_297,In_437);
nand U4369 (N_4369,In_151,In_881);
or U4370 (N_4370,In_175,In_856);
or U4371 (N_4371,In_717,In_7);
nor U4372 (N_4372,In_656,In_293);
or U4373 (N_4373,In_518,In_150);
nor U4374 (N_4374,In_501,In_78);
nor U4375 (N_4375,In_251,In_788);
nand U4376 (N_4376,In_571,In_822);
or U4377 (N_4377,In_234,In_36);
nor U4378 (N_4378,In_797,In_795);
nor U4379 (N_4379,In_616,In_381);
and U4380 (N_4380,In_275,In_533);
and U4381 (N_4381,In_762,In_893);
or U4382 (N_4382,In_788,In_848);
nor U4383 (N_4383,In_465,In_609);
and U4384 (N_4384,In_379,In_906);
or U4385 (N_4385,In_56,In_30);
or U4386 (N_4386,In_604,In_135);
or U4387 (N_4387,In_115,In_786);
nand U4388 (N_4388,In_109,In_500);
nand U4389 (N_4389,In_177,In_781);
nor U4390 (N_4390,In_356,In_339);
or U4391 (N_4391,In_333,In_822);
or U4392 (N_4392,In_449,In_334);
nor U4393 (N_4393,In_699,In_97);
nor U4394 (N_4394,In_202,In_518);
nor U4395 (N_4395,In_804,In_461);
nand U4396 (N_4396,In_914,In_42);
and U4397 (N_4397,In_538,In_163);
nand U4398 (N_4398,In_385,In_835);
nand U4399 (N_4399,In_861,In_760);
nor U4400 (N_4400,In_532,In_213);
or U4401 (N_4401,In_548,In_577);
nand U4402 (N_4402,In_167,In_331);
nor U4403 (N_4403,In_386,In_786);
nand U4404 (N_4404,In_224,In_127);
nand U4405 (N_4405,In_466,In_136);
or U4406 (N_4406,In_867,In_457);
nand U4407 (N_4407,In_103,In_102);
and U4408 (N_4408,In_766,In_439);
or U4409 (N_4409,In_737,In_299);
and U4410 (N_4410,In_583,In_44);
nand U4411 (N_4411,In_853,In_63);
nand U4412 (N_4412,In_235,In_49);
nand U4413 (N_4413,In_497,In_667);
and U4414 (N_4414,In_251,In_482);
and U4415 (N_4415,In_22,In_90);
or U4416 (N_4416,In_8,In_314);
xor U4417 (N_4417,In_50,In_883);
nand U4418 (N_4418,In_161,In_148);
xnor U4419 (N_4419,In_512,In_838);
nor U4420 (N_4420,In_988,In_760);
or U4421 (N_4421,In_20,In_735);
and U4422 (N_4422,In_491,In_183);
and U4423 (N_4423,In_732,In_162);
or U4424 (N_4424,In_925,In_710);
and U4425 (N_4425,In_274,In_520);
nor U4426 (N_4426,In_375,In_234);
and U4427 (N_4427,In_421,In_708);
nand U4428 (N_4428,In_847,In_852);
or U4429 (N_4429,In_161,In_512);
or U4430 (N_4430,In_346,In_870);
nor U4431 (N_4431,In_937,In_795);
and U4432 (N_4432,In_289,In_281);
or U4433 (N_4433,In_432,In_629);
nor U4434 (N_4434,In_793,In_731);
or U4435 (N_4435,In_524,In_958);
nand U4436 (N_4436,In_781,In_614);
and U4437 (N_4437,In_143,In_319);
and U4438 (N_4438,In_954,In_495);
nand U4439 (N_4439,In_131,In_478);
or U4440 (N_4440,In_395,In_401);
or U4441 (N_4441,In_534,In_421);
and U4442 (N_4442,In_940,In_267);
or U4443 (N_4443,In_219,In_905);
or U4444 (N_4444,In_139,In_723);
nor U4445 (N_4445,In_546,In_27);
nor U4446 (N_4446,In_795,In_8);
or U4447 (N_4447,In_25,In_289);
and U4448 (N_4448,In_260,In_771);
or U4449 (N_4449,In_617,In_684);
and U4450 (N_4450,In_616,In_635);
and U4451 (N_4451,In_32,In_84);
nand U4452 (N_4452,In_910,In_91);
and U4453 (N_4453,In_443,In_590);
or U4454 (N_4454,In_632,In_964);
and U4455 (N_4455,In_436,In_371);
nand U4456 (N_4456,In_494,In_620);
and U4457 (N_4457,In_857,In_350);
or U4458 (N_4458,In_629,In_812);
and U4459 (N_4459,In_172,In_90);
nand U4460 (N_4460,In_791,In_855);
and U4461 (N_4461,In_466,In_764);
nand U4462 (N_4462,In_619,In_461);
and U4463 (N_4463,In_272,In_982);
or U4464 (N_4464,In_578,In_250);
or U4465 (N_4465,In_950,In_686);
and U4466 (N_4466,In_934,In_123);
nand U4467 (N_4467,In_273,In_912);
nand U4468 (N_4468,In_654,In_954);
or U4469 (N_4469,In_319,In_379);
or U4470 (N_4470,In_248,In_688);
nor U4471 (N_4471,In_712,In_61);
nand U4472 (N_4472,In_140,In_565);
nor U4473 (N_4473,In_889,In_571);
and U4474 (N_4474,In_543,In_829);
nor U4475 (N_4475,In_890,In_169);
and U4476 (N_4476,In_543,In_233);
nand U4477 (N_4477,In_609,In_292);
xnor U4478 (N_4478,In_163,In_748);
xor U4479 (N_4479,In_83,In_569);
or U4480 (N_4480,In_867,In_620);
nor U4481 (N_4481,In_925,In_544);
and U4482 (N_4482,In_302,In_307);
or U4483 (N_4483,In_575,In_799);
nor U4484 (N_4484,In_735,In_122);
and U4485 (N_4485,In_799,In_862);
nand U4486 (N_4486,In_707,In_180);
and U4487 (N_4487,In_386,In_225);
nor U4488 (N_4488,In_830,In_367);
nand U4489 (N_4489,In_892,In_889);
and U4490 (N_4490,In_96,In_68);
nand U4491 (N_4491,In_485,In_619);
nor U4492 (N_4492,In_183,In_418);
and U4493 (N_4493,In_774,In_724);
nor U4494 (N_4494,In_430,In_124);
nand U4495 (N_4495,In_564,In_486);
nor U4496 (N_4496,In_403,In_952);
nand U4497 (N_4497,In_298,In_299);
or U4498 (N_4498,In_605,In_859);
nand U4499 (N_4499,In_668,In_706);
nand U4500 (N_4500,In_222,In_733);
nor U4501 (N_4501,In_955,In_424);
or U4502 (N_4502,In_520,In_224);
nor U4503 (N_4503,In_171,In_515);
nor U4504 (N_4504,In_216,In_154);
nor U4505 (N_4505,In_880,In_816);
nor U4506 (N_4506,In_741,In_901);
nor U4507 (N_4507,In_217,In_730);
nand U4508 (N_4508,In_579,In_381);
nor U4509 (N_4509,In_749,In_251);
nor U4510 (N_4510,In_415,In_379);
nor U4511 (N_4511,In_683,In_169);
nand U4512 (N_4512,In_92,In_61);
or U4513 (N_4513,In_612,In_227);
and U4514 (N_4514,In_719,In_598);
nand U4515 (N_4515,In_13,In_862);
or U4516 (N_4516,In_827,In_885);
nand U4517 (N_4517,In_106,In_269);
nand U4518 (N_4518,In_495,In_319);
or U4519 (N_4519,In_967,In_397);
nor U4520 (N_4520,In_96,In_407);
nand U4521 (N_4521,In_66,In_159);
nor U4522 (N_4522,In_234,In_520);
or U4523 (N_4523,In_979,In_899);
and U4524 (N_4524,In_43,In_14);
nor U4525 (N_4525,In_520,In_647);
nor U4526 (N_4526,In_913,In_634);
nor U4527 (N_4527,In_419,In_435);
nand U4528 (N_4528,In_56,In_927);
nor U4529 (N_4529,In_417,In_535);
and U4530 (N_4530,In_595,In_796);
nor U4531 (N_4531,In_377,In_75);
nor U4532 (N_4532,In_62,In_298);
or U4533 (N_4533,In_331,In_769);
nor U4534 (N_4534,In_923,In_823);
and U4535 (N_4535,In_744,In_745);
nand U4536 (N_4536,In_559,In_227);
and U4537 (N_4537,In_424,In_166);
and U4538 (N_4538,In_67,In_320);
nor U4539 (N_4539,In_272,In_343);
nand U4540 (N_4540,In_41,In_412);
or U4541 (N_4541,In_236,In_641);
nor U4542 (N_4542,In_883,In_630);
nor U4543 (N_4543,In_11,In_383);
nand U4544 (N_4544,In_646,In_30);
and U4545 (N_4545,In_650,In_713);
and U4546 (N_4546,In_490,In_802);
nor U4547 (N_4547,In_263,In_622);
or U4548 (N_4548,In_315,In_317);
nor U4549 (N_4549,In_693,In_600);
nor U4550 (N_4550,In_512,In_839);
and U4551 (N_4551,In_108,In_480);
nor U4552 (N_4552,In_876,In_632);
and U4553 (N_4553,In_486,In_156);
and U4554 (N_4554,In_737,In_580);
and U4555 (N_4555,In_291,In_334);
and U4556 (N_4556,In_316,In_450);
nand U4557 (N_4557,In_255,In_762);
nand U4558 (N_4558,In_51,In_621);
nand U4559 (N_4559,In_962,In_188);
nor U4560 (N_4560,In_874,In_339);
nor U4561 (N_4561,In_978,In_243);
and U4562 (N_4562,In_240,In_855);
and U4563 (N_4563,In_743,In_234);
nor U4564 (N_4564,In_347,In_396);
nor U4565 (N_4565,In_751,In_118);
nand U4566 (N_4566,In_544,In_206);
and U4567 (N_4567,In_462,In_127);
or U4568 (N_4568,In_131,In_15);
nand U4569 (N_4569,In_9,In_894);
nor U4570 (N_4570,In_641,In_182);
and U4571 (N_4571,In_134,In_929);
nand U4572 (N_4572,In_194,In_96);
nand U4573 (N_4573,In_593,In_688);
nand U4574 (N_4574,In_138,In_629);
or U4575 (N_4575,In_325,In_191);
or U4576 (N_4576,In_844,In_795);
or U4577 (N_4577,In_125,In_301);
nor U4578 (N_4578,In_557,In_425);
nand U4579 (N_4579,In_793,In_195);
nor U4580 (N_4580,In_786,In_949);
nor U4581 (N_4581,In_94,In_456);
or U4582 (N_4582,In_202,In_669);
nand U4583 (N_4583,In_766,In_932);
and U4584 (N_4584,In_977,In_337);
nand U4585 (N_4585,In_900,In_634);
or U4586 (N_4586,In_760,In_502);
or U4587 (N_4587,In_199,In_157);
nor U4588 (N_4588,In_976,In_81);
nor U4589 (N_4589,In_727,In_767);
nor U4590 (N_4590,In_882,In_412);
nand U4591 (N_4591,In_119,In_448);
and U4592 (N_4592,In_838,In_666);
nand U4593 (N_4593,In_44,In_268);
and U4594 (N_4594,In_491,In_580);
nor U4595 (N_4595,In_217,In_439);
and U4596 (N_4596,In_208,In_735);
or U4597 (N_4597,In_128,In_218);
and U4598 (N_4598,In_820,In_348);
and U4599 (N_4599,In_173,In_186);
or U4600 (N_4600,In_996,In_76);
nor U4601 (N_4601,In_700,In_694);
nor U4602 (N_4602,In_476,In_311);
or U4603 (N_4603,In_14,In_324);
and U4604 (N_4604,In_116,In_671);
nor U4605 (N_4605,In_145,In_95);
nand U4606 (N_4606,In_834,In_942);
nor U4607 (N_4607,In_627,In_952);
nor U4608 (N_4608,In_588,In_134);
nor U4609 (N_4609,In_415,In_467);
nand U4610 (N_4610,In_733,In_109);
nor U4611 (N_4611,In_634,In_549);
nand U4612 (N_4612,In_90,In_119);
or U4613 (N_4613,In_500,In_13);
or U4614 (N_4614,In_894,In_213);
or U4615 (N_4615,In_708,In_703);
or U4616 (N_4616,In_806,In_969);
and U4617 (N_4617,In_833,In_322);
and U4618 (N_4618,In_218,In_924);
or U4619 (N_4619,In_836,In_762);
nor U4620 (N_4620,In_727,In_444);
nand U4621 (N_4621,In_738,In_870);
nor U4622 (N_4622,In_454,In_326);
and U4623 (N_4623,In_105,In_359);
nand U4624 (N_4624,In_272,In_284);
nand U4625 (N_4625,In_704,In_539);
and U4626 (N_4626,In_400,In_788);
or U4627 (N_4627,In_605,In_24);
xnor U4628 (N_4628,In_16,In_595);
and U4629 (N_4629,In_132,In_187);
nor U4630 (N_4630,In_512,In_403);
or U4631 (N_4631,In_735,In_15);
and U4632 (N_4632,In_790,In_566);
nor U4633 (N_4633,In_346,In_331);
nand U4634 (N_4634,In_145,In_253);
nor U4635 (N_4635,In_370,In_293);
or U4636 (N_4636,In_666,In_413);
and U4637 (N_4637,In_995,In_939);
nand U4638 (N_4638,In_364,In_226);
or U4639 (N_4639,In_921,In_956);
nor U4640 (N_4640,In_162,In_655);
nor U4641 (N_4641,In_658,In_398);
or U4642 (N_4642,In_894,In_633);
nand U4643 (N_4643,In_275,In_748);
nand U4644 (N_4644,In_195,In_175);
or U4645 (N_4645,In_663,In_59);
nand U4646 (N_4646,In_853,In_832);
nor U4647 (N_4647,In_625,In_8);
and U4648 (N_4648,In_67,In_210);
nand U4649 (N_4649,In_390,In_764);
nor U4650 (N_4650,In_65,In_425);
and U4651 (N_4651,In_906,In_149);
nand U4652 (N_4652,In_256,In_808);
or U4653 (N_4653,In_267,In_581);
or U4654 (N_4654,In_376,In_991);
and U4655 (N_4655,In_394,In_531);
nor U4656 (N_4656,In_734,In_978);
nor U4657 (N_4657,In_996,In_524);
nand U4658 (N_4658,In_601,In_403);
and U4659 (N_4659,In_887,In_454);
and U4660 (N_4660,In_869,In_652);
nand U4661 (N_4661,In_212,In_324);
or U4662 (N_4662,In_519,In_493);
nor U4663 (N_4663,In_417,In_791);
nand U4664 (N_4664,In_654,In_882);
nand U4665 (N_4665,In_266,In_904);
nand U4666 (N_4666,In_674,In_893);
and U4667 (N_4667,In_204,In_47);
nor U4668 (N_4668,In_133,In_60);
nand U4669 (N_4669,In_584,In_243);
or U4670 (N_4670,In_192,In_95);
or U4671 (N_4671,In_825,In_96);
or U4672 (N_4672,In_12,In_43);
nor U4673 (N_4673,In_92,In_823);
or U4674 (N_4674,In_830,In_155);
nor U4675 (N_4675,In_504,In_477);
nor U4676 (N_4676,In_712,In_818);
nand U4677 (N_4677,In_749,In_740);
nor U4678 (N_4678,In_190,In_804);
and U4679 (N_4679,In_909,In_130);
nand U4680 (N_4680,In_10,In_456);
or U4681 (N_4681,In_998,In_620);
or U4682 (N_4682,In_71,In_514);
or U4683 (N_4683,In_761,In_508);
and U4684 (N_4684,In_763,In_162);
or U4685 (N_4685,In_121,In_67);
nor U4686 (N_4686,In_265,In_217);
nor U4687 (N_4687,In_350,In_585);
or U4688 (N_4688,In_333,In_504);
nand U4689 (N_4689,In_849,In_14);
and U4690 (N_4690,In_103,In_192);
nand U4691 (N_4691,In_598,In_609);
and U4692 (N_4692,In_925,In_284);
or U4693 (N_4693,In_582,In_636);
nor U4694 (N_4694,In_207,In_433);
and U4695 (N_4695,In_469,In_467);
or U4696 (N_4696,In_561,In_880);
or U4697 (N_4697,In_544,In_496);
nand U4698 (N_4698,In_981,In_455);
and U4699 (N_4699,In_203,In_816);
nand U4700 (N_4700,In_678,In_752);
nand U4701 (N_4701,In_396,In_810);
nand U4702 (N_4702,In_186,In_720);
and U4703 (N_4703,In_253,In_483);
or U4704 (N_4704,In_384,In_75);
and U4705 (N_4705,In_119,In_234);
and U4706 (N_4706,In_342,In_646);
nand U4707 (N_4707,In_489,In_998);
and U4708 (N_4708,In_288,In_735);
nor U4709 (N_4709,In_280,In_845);
or U4710 (N_4710,In_517,In_144);
nand U4711 (N_4711,In_581,In_943);
nor U4712 (N_4712,In_564,In_157);
nand U4713 (N_4713,In_756,In_614);
nand U4714 (N_4714,In_789,In_555);
or U4715 (N_4715,In_973,In_29);
nand U4716 (N_4716,In_55,In_925);
nand U4717 (N_4717,In_637,In_423);
nor U4718 (N_4718,In_718,In_133);
or U4719 (N_4719,In_687,In_414);
or U4720 (N_4720,In_689,In_163);
nor U4721 (N_4721,In_840,In_672);
nand U4722 (N_4722,In_671,In_230);
nor U4723 (N_4723,In_8,In_755);
or U4724 (N_4724,In_577,In_789);
nor U4725 (N_4725,In_59,In_932);
and U4726 (N_4726,In_46,In_423);
or U4727 (N_4727,In_115,In_296);
xnor U4728 (N_4728,In_110,In_589);
and U4729 (N_4729,In_605,In_649);
and U4730 (N_4730,In_132,In_358);
nor U4731 (N_4731,In_109,In_441);
nor U4732 (N_4732,In_506,In_410);
and U4733 (N_4733,In_576,In_765);
and U4734 (N_4734,In_150,In_591);
and U4735 (N_4735,In_271,In_759);
or U4736 (N_4736,In_605,In_602);
and U4737 (N_4737,In_112,In_708);
and U4738 (N_4738,In_281,In_217);
or U4739 (N_4739,In_305,In_858);
or U4740 (N_4740,In_150,In_774);
and U4741 (N_4741,In_483,In_120);
and U4742 (N_4742,In_341,In_962);
nand U4743 (N_4743,In_462,In_496);
nand U4744 (N_4744,In_576,In_750);
or U4745 (N_4745,In_810,In_476);
and U4746 (N_4746,In_250,In_209);
or U4747 (N_4747,In_948,In_840);
or U4748 (N_4748,In_700,In_756);
nand U4749 (N_4749,In_429,In_439);
and U4750 (N_4750,In_771,In_475);
or U4751 (N_4751,In_973,In_361);
nand U4752 (N_4752,In_296,In_580);
nand U4753 (N_4753,In_559,In_605);
and U4754 (N_4754,In_965,In_542);
or U4755 (N_4755,In_330,In_992);
nor U4756 (N_4756,In_386,In_202);
and U4757 (N_4757,In_94,In_1);
or U4758 (N_4758,In_250,In_984);
nor U4759 (N_4759,In_670,In_882);
nand U4760 (N_4760,In_120,In_477);
and U4761 (N_4761,In_886,In_244);
or U4762 (N_4762,In_121,In_981);
nor U4763 (N_4763,In_253,In_748);
and U4764 (N_4764,In_201,In_689);
or U4765 (N_4765,In_168,In_739);
nor U4766 (N_4766,In_750,In_66);
nand U4767 (N_4767,In_123,In_522);
and U4768 (N_4768,In_213,In_814);
nand U4769 (N_4769,In_700,In_16);
or U4770 (N_4770,In_320,In_308);
nand U4771 (N_4771,In_578,In_907);
and U4772 (N_4772,In_572,In_450);
nor U4773 (N_4773,In_607,In_269);
nor U4774 (N_4774,In_394,In_935);
nor U4775 (N_4775,In_306,In_674);
nor U4776 (N_4776,In_420,In_194);
and U4777 (N_4777,In_845,In_799);
nand U4778 (N_4778,In_246,In_263);
or U4779 (N_4779,In_940,In_606);
nor U4780 (N_4780,In_466,In_201);
or U4781 (N_4781,In_690,In_947);
and U4782 (N_4782,In_4,In_794);
and U4783 (N_4783,In_394,In_880);
or U4784 (N_4784,In_866,In_614);
or U4785 (N_4785,In_550,In_902);
or U4786 (N_4786,In_970,In_640);
or U4787 (N_4787,In_697,In_716);
nand U4788 (N_4788,In_773,In_471);
and U4789 (N_4789,In_62,In_58);
nand U4790 (N_4790,In_236,In_174);
nand U4791 (N_4791,In_312,In_40);
and U4792 (N_4792,In_796,In_177);
or U4793 (N_4793,In_693,In_891);
and U4794 (N_4794,In_165,In_79);
and U4795 (N_4795,In_122,In_819);
and U4796 (N_4796,In_215,In_343);
nor U4797 (N_4797,In_871,In_635);
nand U4798 (N_4798,In_9,In_296);
or U4799 (N_4799,In_338,In_163);
nand U4800 (N_4800,In_374,In_650);
and U4801 (N_4801,In_248,In_366);
and U4802 (N_4802,In_717,In_350);
and U4803 (N_4803,In_318,In_254);
nand U4804 (N_4804,In_450,In_348);
nor U4805 (N_4805,In_96,In_512);
or U4806 (N_4806,In_146,In_79);
nor U4807 (N_4807,In_618,In_795);
nor U4808 (N_4808,In_297,In_180);
or U4809 (N_4809,In_587,In_397);
or U4810 (N_4810,In_944,In_149);
or U4811 (N_4811,In_672,In_616);
or U4812 (N_4812,In_187,In_58);
xnor U4813 (N_4813,In_94,In_127);
nand U4814 (N_4814,In_678,In_450);
nor U4815 (N_4815,In_528,In_485);
xor U4816 (N_4816,In_768,In_965);
nor U4817 (N_4817,In_660,In_871);
and U4818 (N_4818,In_213,In_524);
or U4819 (N_4819,In_296,In_523);
nand U4820 (N_4820,In_590,In_826);
nand U4821 (N_4821,In_354,In_696);
nor U4822 (N_4822,In_4,In_369);
nor U4823 (N_4823,In_888,In_983);
xor U4824 (N_4824,In_406,In_825);
and U4825 (N_4825,In_948,In_8);
xnor U4826 (N_4826,In_445,In_196);
nand U4827 (N_4827,In_476,In_836);
and U4828 (N_4828,In_162,In_511);
nor U4829 (N_4829,In_445,In_69);
and U4830 (N_4830,In_237,In_440);
or U4831 (N_4831,In_809,In_69);
and U4832 (N_4832,In_470,In_75);
or U4833 (N_4833,In_94,In_438);
and U4834 (N_4834,In_877,In_268);
nor U4835 (N_4835,In_103,In_380);
nor U4836 (N_4836,In_839,In_588);
nand U4837 (N_4837,In_314,In_794);
or U4838 (N_4838,In_304,In_813);
nor U4839 (N_4839,In_347,In_124);
and U4840 (N_4840,In_583,In_539);
or U4841 (N_4841,In_11,In_756);
nand U4842 (N_4842,In_770,In_91);
and U4843 (N_4843,In_825,In_253);
or U4844 (N_4844,In_867,In_176);
and U4845 (N_4845,In_443,In_481);
nor U4846 (N_4846,In_784,In_911);
nor U4847 (N_4847,In_771,In_198);
nand U4848 (N_4848,In_614,In_791);
nand U4849 (N_4849,In_966,In_903);
nor U4850 (N_4850,In_521,In_138);
and U4851 (N_4851,In_329,In_883);
and U4852 (N_4852,In_339,In_260);
nand U4853 (N_4853,In_856,In_905);
and U4854 (N_4854,In_835,In_498);
xor U4855 (N_4855,In_710,In_52);
or U4856 (N_4856,In_77,In_700);
and U4857 (N_4857,In_33,In_282);
or U4858 (N_4858,In_101,In_44);
or U4859 (N_4859,In_236,In_809);
nand U4860 (N_4860,In_87,In_440);
and U4861 (N_4861,In_334,In_667);
nand U4862 (N_4862,In_426,In_637);
nor U4863 (N_4863,In_106,In_323);
nor U4864 (N_4864,In_444,In_577);
nor U4865 (N_4865,In_810,In_296);
nand U4866 (N_4866,In_929,In_279);
nand U4867 (N_4867,In_613,In_672);
and U4868 (N_4868,In_495,In_11);
nand U4869 (N_4869,In_490,In_964);
nor U4870 (N_4870,In_279,In_684);
and U4871 (N_4871,In_131,In_148);
and U4872 (N_4872,In_73,In_35);
nand U4873 (N_4873,In_494,In_497);
or U4874 (N_4874,In_131,In_732);
or U4875 (N_4875,In_960,In_705);
nor U4876 (N_4876,In_491,In_582);
nor U4877 (N_4877,In_557,In_914);
or U4878 (N_4878,In_551,In_187);
nand U4879 (N_4879,In_652,In_936);
nor U4880 (N_4880,In_846,In_730);
and U4881 (N_4881,In_159,In_412);
or U4882 (N_4882,In_654,In_670);
and U4883 (N_4883,In_721,In_922);
or U4884 (N_4884,In_380,In_919);
or U4885 (N_4885,In_803,In_734);
and U4886 (N_4886,In_139,In_226);
or U4887 (N_4887,In_132,In_123);
or U4888 (N_4888,In_698,In_215);
and U4889 (N_4889,In_568,In_25);
or U4890 (N_4890,In_932,In_188);
or U4891 (N_4891,In_712,In_797);
nor U4892 (N_4892,In_822,In_119);
nor U4893 (N_4893,In_537,In_311);
xnor U4894 (N_4894,In_349,In_881);
nor U4895 (N_4895,In_650,In_105);
or U4896 (N_4896,In_284,In_729);
and U4897 (N_4897,In_735,In_985);
and U4898 (N_4898,In_281,In_957);
nand U4899 (N_4899,In_51,In_967);
nand U4900 (N_4900,In_908,In_86);
and U4901 (N_4901,In_167,In_683);
nand U4902 (N_4902,In_301,In_975);
and U4903 (N_4903,In_884,In_21);
and U4904 (N_4904,In_867,In_189);
nand U4905 (N_4905,In_764,In_995);
nor U4906 (N_4906,In_983,In_682);
nor U4907 (N_4907,In_339,In_324);
nor U4908 (N_4908,In_595,In_940);
and U4909 (N_4909,In_184,In_833);
nand U4910 (N_4910,In_242,In_549);
nand U4911 (N_4911,In_952,In_667);
and U4912 (N_4912,In_640,In_650);
or U4913 (N_4913,In_289,In_694);
or U4914 (N_4914,In_812,In_696);
or U4915 (N_4915,In_996,In_206);
and U4916 (N_4916,In_18,In_62);
xor U4917 (N_4917,In_314,In_894);
nand U4918 (N_4918,In_995,In_242);
nand U4919 (N_4919,In_384,In_705);
and U4920 (N_4920,In_127,In_210);
nand U4921 (N_4921,In_856,In_302);
and U4922 (N_4922,In_507,In_615);
or U4923 (N_4923,In_862,In_685);
or U4924 (N_4924,In_830,In_493);
nor U4925 (N_4925,In_918,In_287);
and U4926 (N_4926,In_879,In_986);
nand U4927 (N_4927,In_1,In_394);
and U4928 (N_4928,In_643,In_584);
nand U4929 (N_4929,In_319,In_981);
nand U4930 (N_4930,In_981,In_24);
or U4931 (N_4931,In_583,In_48);
or U4932 (N_4932,In_732,In_469);
nor U4933 (N_4933,In_752,In_838);
nand U4934 (N_4934,In_62,In_220);
nand U4935 (N_4935,In_196,In_913);
nor U4936 (N_4936,In_414,In_222);
nor U4937 (N_4937,In_27,In_42);
nand U4938 (N_4938,In_816,In_210);
nor U4939 (N_4939,In_207,In_664);
and U4940 (N_4940,In_658,In_217);
nor U4941 (N_4941,In_587,In_329);
or U4942 (N_4942,In_246,In_619);
or U4943 (N_4943,In_359,In_654);
nor U4944 (N_4944,In_366,In_117);
and U4945 (N_4945,In_209,In_773);
and U4946 (N_4946,In_767,In_742);
nand U4947 (N_4947,In_761,In_474);
and U4948 (N_4948,In_459,In_785);
or U4949 (N_4949,In_383,In_222);
nand U4950 (N_4950,In_277,In_327);
and U4951 (N_4951,In_152,In_677);
nor U4952 (N_4952,In_467,In_510);
nor U4953 (N_4953,In_91,In_829);
and U4954 (N_4954,In_67,In_732);
nor U4955 (N_4955,In_322,In_564);
and U4956 (N_4956,In_569,In_869);
nor U4957 (N_4957,In_660,In_933);
and U4958 (N_4958,In_230,In_752);
and U4959 (N_4959,In_955,In_989);
nand U4960 (N_4960,In_519,In_900);
nor U4961 (N_4961,In_911,In_396);
xnor U4962 (N_4962,In_209,In_839);
or U4963 (N_4963,In_374,In_548);
and U4964 (N_4964,In_11,In_258);
nand U4965 (N_4965,In_505,In_930);
or U4966 (N_4966,In_181,In_673);
or U4967 (N_4967,In_475,In_591);
and U4968 (N_4968,In_916,In_658);
or U4969 (N_4969,In_499,In_3);
nand U4970 (N_4970,In_567,In_834);
or U4971 (N_4971,In_364,In_998);
nor U4972 (N_4972,In_785,In_108);
or U4973 (N_4973,In_960,In_603);
nand U4974 (N_4974,In_871,In_296);
nand U4975 (N_4975,In_67,In_633);
nand U4976 (N_4976,In_501,In_70);
nor U4977 (N_4977,In_866,In_751);
nand U4978 (N_4978,In_422,In_493);
or U4979 (N_4979,In_854,In_754);
or U4980 (N_4980,In_188,In_165);
or U4981 (N_4981,In_698,In_393);
or U4982 (N_4982,In_85,In_473);
nor U4983 (N_4983,In_662,In_933);
nor U4984 (N_4984,In_596,In_45);
nor U4985 (N_4985,In_199,In_63);
or U4986 (N_4986,In_750,In_734);
or U4987 (N_4987,In_84,In_797);
or U4988 (N_4988,In_268,In_651);
nor U4989 (N_4989,In_776,In_728);
nand U4990 (N_4990,In_419,In_752);
and U4991 (N_4991,In_620,In_41);
nand U4992 (N_4992,In_261,In_334);
or U4993 (N_4993,In_327,In_267);
or U4994 (N_4994,In_161,In_417);
or U4995 (N_4995,In_39,In_710);
nand U4996 (N_4996,In_348,In_187);
or U4997 (N_4997,In_964,In_971);
xor U4998 (N_4998,In_445,In_649);
nor U4999 (N_4999,In_841,In_752);
nand U5000 (N_5000,N_722,N_4404);
and U5001 (N_5001,N_3419,N_1995);
nand U5002 (N_5002,N_227,N_230);
nor U5003 (N_5003,N_1828,N_4765);
nor U5004 (N_5004,N_542,N_1623);
nor U5005 (N_5005,N_3301,N_2611);
nor U5006 (N_5006,N_1080,N_2529);
nand U5007 (N_5007,N_82,N_4696);
nand U5008 (N_5008,N_2169,N_289);
or U5009 (N_5009,N_506,N_1233);
nand U5010 (N_5010,N_684,N_411);
or U5011 (N_5011,N_2860,N_2936);
and U5012 (N_5012,N_2202,N_2621);
and U5013 (N_5013,N_40,N_1700);
or U5014 (N_5014,N_1257,N_2285);
nand U5015 (N_5015,N_2708,N_2219);
and U5016 (N_5016,N_2438,N_3441);
and U5017 (N_5017,N_1895,N_3006);
nand U5018 (N_5018,N_4542,N_394);
nor U5019 (N_5019,N_3411,N_486);
nand U5020 (N_5020,N_1315,N_2259);
or U5021 (N_5021,N_832,N_256);
nor U5022 (N_5022,N_4116,N_866);
and U5023 (N_5023,N_4079,N_1903);
or U5024 (N_5024,N_4844,N_71);
nand U5025 (N_5025,N_2674,N_2363);
nand U5026 (N_5026,N_2516,N_3068);
or U5027 (N_5027,N_3726,N_2849);
nor U5028 (N_5028,N_2535,N_4094);
or U5029 (N_5029,N_1775,N_1920);
and U5030 (N_5030,N_2176,N_3947);
or U5031 (N_5031,N_4881,N_4572);
or U5032 (N_5032,N_4208,N_2852);
nor U5033 (N_5033,N_3921,N_701);
nor U5034 (N_5034,N_4521,N_881);
nor U5035 (N_5035,N_673,N_1583);
and U5036 (N_5036,N_3599,N_3474);
nor U5037 (N_5037,N_3048,N_4221);
nor U5038 (N_5038,N_3970,N_1224);
and U5039 (N_5039,N_1928,N_1516);
and U5040 (N_5040,N_149,N_3230);
or U5041 (N_5041,N_3362,N_91);
nand U5042 (N_5042,N_1880,N_2778);
or U5043 (N_5043,N_333,N_1591);
nor U5044 (N_5044,N_4308,N_1353);
and U5045 (N_5045,N_2972,N_3330);
nand U5046 (N_5046,N_4742,N_4201);
nor U5047 (N_5047,N_492,N_3909);
and U5048 (N_5048,N_1253,N_1944);
and U5049 (N_5049,N_2262,N_2079);
nand U5050 (N_5050,N_4279,N_3566);
and U5051 (N_5051,N_1898,N_51);
or U5052 (N_5052,N_2297,N_1105);
and U5053 (N_5053,N_4135,N_2098);
or U5054 (N_5054,N_3002,N_315);
or U5055 (N_5055,N_4974,N_4200);
nand U5056 (N_5056,N_1184,N_2080);
and U5057 (N_5057,N_4351,N_3359);
nand U5058 (N_5058,N_283,N_2786);
and U5059 (N_5059,N_3174,N_4719);
and U5060 (N_5060,N_2802,N_824);
nand U5061 (N_5061,N_2105,N_2833);
nor U5062 (N_5062,N_3737,N_4724);
nor U5063 (N_5063,N_4140,N_4868);
and U5064 (N_5064,N_1753,N_347);
and U5065 (N_5065,N_1457,N_1242);
nor U5066 (N_5066,N_682,N_549);
and U5067 (N_5067,N_4539,N_4027);
nand U5068 (N_5068,N_1128,N_167);
nand U5069 (N_5069,N_401,N_2389);
and U5070 (N_5070,N_1280,N_2942);
nor U5071 (N_5071,N_3029,N_780);
and U5072 (N_5072,N_4635,N_3437);
nor U5073 (N_5073,N_1857,N_2827);
nand U5074 (N_5074,N_2247,N_4893);
and U5075 (N_5075,N_233,N_2814);
xor U5076 (N_5076,N_3616,N_1476);
or U5077 (N_5077,N_4908,N_4268);
nand U5078 (N_5078,N_1447,N_1470);
nand U5079 (N_5079,N_766,N_3024);
nand U5080 (N_5080,N_4357,N_1258);
or U5081 (N_5081,N_893,N_4008);
and U5082 (N_5082,N_4360,N_4016);
nor U5083 (N_5083,N_4468,N_2911);
nand U5084 (N_5084,N_4904,N_3856);
or U5085 (N_5085,N_4128,N_925);
and U5086 (N_5086,N_1567,N_3932);
or U5087 (N_5087,N_1384,N_3762);
and U5088 (N_5088,N_1617,N_309);
nand U5089 (N_5089,N_1374,N_3548);
nand U5090 (N_5090,N_4647,N_480);
nand U5091 (N_5091,N_1252,N_4217);
nor U5092 (N_5092,N_4501,N_2239);
and U5093 (N_5093,N_1788,N_85);
and U5094 (N_5094,N_1714,N_4843);
or U5095 (N_5095,N_108,N_238);
nand U5096 (N_5096,N_2561,N_2891);
xnor U5097 (N_5097,N_1207,N_4356);
nor U5098 (N_5098,N_63,N_4512);
nand U5099 (N_5099,N_4957,N_2109);
nand U5100 (N_5100,N_3687,N_3070);
or U5101 (N_5101,N_1984,N_4414);
nor U5102 (N_5102,N_226,N_2783);
or U5103 (N_5103,N_4388,N_635);
and U5104 (N_5104,N_584,N_1621);
and U5105 (N_5105,N_792,N_3235);
nor U5106 (N_5106,N_397,N_1862);
or U5107 (N_5107,N_3078,N_1445);
nor U5108 (N_5108,N_1906,N_1912);
and U5109 (N_5109,N_4232,N_3335);
nand U5110 (N_5110,N_3018,N_4629);
and U5111 (N_5111,N_4456,N_214);
and U5112 (N_5112,N_209,N_15);
nor U5113 (N_5113,N_580,N_675);
nor U5114 (N_5114,N_2213,N_1795);
or U5115 (N_5115,N_1355,N_236);
nand U5116 (N_5116,N_243,N_2836);
and U5117 (N_5117,N_2792,N_3483);
or U5118 (N_5118,N_3770,N_1245);
or U5119 (N_5119,N_1217,N_2075);
nor U5120 (N_5120,N_1138,N_2043);
or U5121 (N_5121,N_61,N_4144);
and U5122 (N_5122,N_3169,N_2515);
nor U5123 (N_5123,N_3735,N_4337);
nand U5124 (N_5124,N_4259,N_4364);
or U5125 (N_5125,N_1879,N_3505);
nand U5126 (N_5126,N_3473,N_2492);
and U5127 (N_5127,N_2279,N_1902);
and U5128 (N_5128,N_2137,N_1405);
nor U5129 (N_5129,N_4828,N_3692);
and U5130 (N_5130,N_679,N_3738);
or U5131 (N_5131,N_4523,N_2397);
nor U5132 (N_5132,N_2083,N_1295);
nor U5133 (N_5133,N_1861,N_4601);
nand U5134 (N_5134,N_939,N_3279);
nand U5135 (N_5135,N_1216,N_3630);
nor U5136 (N_5136,N_2918,N_280);
and U5137 (N_5137,N_468,N_1799);
nor U5138 (N_5138,N_1129,N_3944);
or U5139 (N_5139,N_2152,N_3775);
or U5140 (N_5140,N_693,N_406);
nand U5141 (N_5141,N_3847,N_1218);
or U5142 (N_5142,N_84,N_2995);
nand U5143 (N_5143,N_4177,N_3522);
nand U5144 (N_5144,N_3972,N_2038);
or U5145 (N_5145,N_2121,N_4444);
or U5146 (N_5146,N_4980,N_647);
nand U5147 (N_5147,N_2633,N_1663);
and U5148 (N_5148,N_3284,N_417);
and U5149 (N_5149,N_357,N_253);
or U5150 (N_5150,N_1602,N_450);
nand U5151 (N_5151,N_1026,N_1488);
nand U5152 (N_5152,N_29,N_36);
or U5153 (N_5153,N_2551,N_3826);
nor U5154 (N_5154,N_1084,N_4538);
nand U5155 (N_5155,N_1446,N_1502);
or U5156 (N_5156,N_93,N_1744);
and U5157 (N_5157,N_1115,N_1812);
and U5158 (N_5158,N_4049,N_3644);
or U5159 (N_5159,N_546,N_3128);
nand U5160 (N_5160,N_1691,N_3067);
nor U5161 (N_5161,N_4657,N_799);
or U5162 (N_5162,N_3189,N_3447);
and U5163 (N_5163,N_306,N_1001);
nand U5164 (N_5164,N_64,N_307);
and U5165 (N_5165,N_2634,N_4085);
and U5166 (N_5166,N_2823,N_14);
nor U5167 (N_5167,N_4443,N_4431);
nand U5168 (N_5168,N_4046,N_586);
nor U5169 (N_5169,N_3240,N_3171);
and U5170 (N_5170,N_2355,N_1041);
and U5171 (N_5171,N_3310,N_3297);
or U5172 (N_5172,N_4889,N_1655);
nand U5173 (N_5173,N_3320,N_2930);
nand U5174 (N_5174,N_2673,N_3998);
and U5175 (N_5175,N_706,N_1509);
nor U5176 (N_5176,N_2686,N_332);
and U5177 (N_5177,N_2116,N_4557);
nor U5178 (N_5178,N_3901,N_1342);
nand U5179 (N_5179,N_1222,N_3443);
nand U5180 (N_5180,N_1859,N_4391);
and U5181 (N_5181,N_2653,N_2971);
nand U5182 (N_5182,N_3269,N_1779);
and U5183 (N_5183,N_537,N_3044);
and U5184 (N_5184,N_3400,N_694);
nand U5185 (N_5185,N_982,N_1133);
or U5186 (N_5186,N_2520,N_451);
and U5187 (N_5187,N_4457,N_4579);
nor U5188 (N_5188,N_2587,N_4568);
nor U5189 (N_5189,N_190,N_2504);
nand U5190 (N_5190,N_1734,N_3224);
or U5191 (N_5191,N_4888,N_259);
nor U5192 (N_5192,N_4989,N_2395);
and U5193 (N_5193,N_1275,N_2073);
nand U5194 (N_5194,N_2908,N_155);
nor U5195 (N_5195,N_2089,N_3165);
and U5196 (N_5196,N_2224,N_3794);
and U5197 (N_5197,N_793,N_4979);
nor U5198 (N_5198,N_589,N_3129);
or U5199 (N_5199,N_4303,N_4172);
and U5200 (N_5200,N_1586,N_2409);
or U5201 (N_5201,N_2639,N_3654);
nand U5202 (N_5202,N_2149,N_2555);
nor U5203 (N_5203,N_3621,N_1843);
xor U5204 (N_5204,N_1540,N_2939);
or U5205 (N_5205,N_1597,N_2312);
and U5206 (N_5206,N_1251,N_1611);
nand U5207 (N_5207,N_1420,N_1800);
nand U5208 (N_5208,N_3523,N_2052);
nand U5209 (N_5209,N_1177,N_1225);
nor U5210 (N_5210,N_1936,N_3296);
nor U5211 (N_5211,N_1571,N_4193);
or U5212 (N_5212,N_3047,N_2484);
or U5213 (N_5213,N_1176,N_2097);
nor U5214 (N_5214,N_908,N_1182);
or U5215 (N_5215,N_403,N_1229);
or U5216 (N_5216,N_3436,N_3990);
or U5217 (N_5217,N_2789,N_4389);
and U5218 (N_5218,N_1035,N_2145);
nand U5219 (N_5219,N_877,N_663);
and U5220 (N_5220,N_4118,N_2984);
and U5221 (N_5221,N_2842,N_3346);
and U5222 (N_5222,N_1599,N_3575);
or U5223 (N_5223,N_871,N_1208);
and U5224 (N_5224,N_498,N_4341);
or U5225 (N_5225,N_2134,N_4277);
and U5226 (N_5226,N_4614,N_2607);
nor U5227 (N_5227,N_4628,N_4358);
and U5228 (N_5228,N_3118,N_2615);
nor U5229 (N_5229,N_355,N_453);
and U5230 (N_5230,N_3595,N_721);
and U5231 (N_5231,N_775,N_4921);
nor U5232 (N_5232,N_2877,N_1338);
nand U5233 (N_5233,N_1768,N_1822);
nor U5234 (N_5234,N_3622,N_505);
and U5235 (N_5235,N_4660,N_2457);
nand U5236 (N_5236,N_4339,N_3699);
and U5237 (N_5237,N_3102,N_2528);
or U5238 (N_5238,N_418,N_3210);
and U5239 (N_5239,N_4237,N_1034);
or U5240 (N_5240,N_2315,N_2273);
nand U5241 (N_5241,N_2595,N_4439);
nand U5242 (N_5242,N_3625,N_3053);
nor U5243 (N_5243,N_2039,N_3767);
nor U5244 (N_5244,N_1410,N_2147);
or U5245 (N_5245,N_1747,N_1475);
nor U5246 (N_5246,N_494,N_1722);
and U5247 (N_5247,N_590,N_3456);
nor U5248 (N_5248,N_4879,N_1300);
and U5249 (N_5249,N_2072,N_4331);
or U5250 (N_5250,N_4694,N_4772);
nand U5251 (N_5251,N_2710,N_4990);
and U5252 (N_5252,N_2254,N_2980);
xor U5253 (N_5253,N_111,N_2549);
or U5254 (N_5254,N_4771,N_2030);
nor U5255 (N_5255,N_330,N_1578);
nor U5256 (N_5256,N_4190,N_1652);
and U5257 (N_5257,N_1842,N_4595);
or U5258 (N_5258,N_605,N_1926);
and U5259 (N_5259,N_2195,N_3912);
and U5260 (N_5260,N_2525,N_1283);
and U5261 (N_5261,N_3464,N_717);
or U5262 (N_5262,N_4065,N_2862);
or U5263 (N_5263,N_3401,N_3058);
nand U5264 (N_5264,N_3842,N_1919);
and U5265 (N_5265,N_2976,N_2923);
xor U5266 (N_5266,N_3977,N_4226);
and U5267 (N_5267,N_1570,N_2288);
nand U5268 (N_5268,N_363,N_1407);
or U5269 (N_5269,N_4996,N_1441);
and U5270 (N_5270,N_1847,N_2875);
or U5271 (N_5271,N_1726,N_2948);
nand U5272 (N_5272,N_1894,N_178);
and U5273 (N_5273,N_3969,N_4096);
or U5274 (N_5274,N_1288,N_2664);
nor U5275 (N_5275,N_3779,N_3117);
or U5276 (N_5276,N_1520,N_2157);
or U5277 (N_5277,N_1318,N_652);
nor U5278 (N_5278,N_1977,N_2831);
xor U5279 (N_5279,N_2135,N_3881);
nand U5280 (N_5280,N_602,N_2122);
or U5281 (N_5281,N_1230,N_3529);
nand U5282 (N_5282,N_748,N_420);
nand U5283 (N_5283,N_3648,N_3509);
or U5284 (N_5284,N_3982,N_835);
nor U5285 (N_5285,N_2441,N_291);
nor U5286 (N_5286,N_1750,N_20);
nor U5287 (N_5287,N_593,N_1631);
or U5288 (N_5288,N_4048,N_142);
nor U5289 (N_5289,N_4154,N_944);
nand U5290 (N_5290,N_1990,N_445);
nand U5291 (N_5291,N_4463,N_317);
and U5292 (N_5292,N_206,N_3431);
or U5293 (N_5293,N_1131,N_4690);
and U5294 (N_5294,N_999,N_3163);
nand U5295 (N_5295,N_1416,N_1363);
or U5296 (N_5296,N_4835,N_3711);
or U5297 (N_5297,N_2377,N_4415);
and U5298 (N_5298,N_2829,N_2882);
nand U5299 (N_5299,N_3403,N_3094);
and U5300 (N_5300,N_3217,N_1007);
or U5301 (N_5301,N_4064,N_4795);
nand U5302 (N_5302,N_2205,N_1062);
or U5303 (N_5303,N_141,N_4914);
and U5304 (N_5304,N_2503,N_4864);
nor U5305 (N_5305,N_2959,N_2846);
nor U5306 (N_5306,N_3634,N_4361);
or U5307 (N_5307,N_4711,N_1945);
and U5308 (N_5308,N_1169,N_2482);
nand U5309 (N_5309,N_2330,N_2008);
nor U5310 (N_5310,N_4440,N_2021);
and U5311 (N_5311,N_3023,N_3175);
nand U5312 (N_5312,N_1680,N_4832);
or U5313 (N_5313,N_714,N_2489);
nand U5314 (N_5314,N_3409,N_4878);
and U5315 (N_5315,N_718,N_4746);
or U5316 (N_5316,N_1885,N_1739);
nand U5317 (N_5317,N_2758,N_3781);
nand U5318 (N_5318,N_4345,N_2820);
nand U5319 (N_5319,N_3334,N_2767);
nor U5320 (N_5320,N_3476,N_115);
nand U5321 (N_5321,N_2667,N_2818);
nor U5322 (N_5322,N_1530,N_3710);
nor U5323 (N_5323,N_3484,N_3827);
nand U5324 (N_5324,N_3375,N_4098);
nand U5325 (N_5325,N_4802,N_4805);
nor U5326 (N_5326,N_1029,N_81);
nand U5327 (N_5327,N_405,N_159);
or U5328 (N_5328,N_3000,N_2426);
nor U5329 (N_5329,N_765,N_250);
or U5330 (N_5330,N_820,N_1019);
and U5331 (N_5331,N_2850,N_2016);
nand U5332 (N_5332,N_3590,N_3724);
nor U5333 (N_5333,N_4040,N_2593);
and U5334 (N_5334,N_3949,N_4932);
and U5335 (N_5335,N_4618,N_3818);
and U5336 (N_5336,N_692,N_349);
and U5337 (N_5337,N_2935,N_4067);
and U5338 (N_5338,N_517,N_491);
nand U5339 (N_5339,N_1145,N_127);
nand U5340 (N_5340,N_1314,N_4276);
nor U5341 (N_5341,N_4449,N_4166);
nor U5342 (N_5342,N_922,N_1336);
or U5343 (N_5343,N_3577,N_3323);
nand U5344 (N_5344,N_4739,N_4503);
nor U5345 (N_5345,N_3507,N_2553);
or U5346 (N_5346,N_487,N_763);
nand U5347 (N_5347,N_1918,N_4428);
nor U5348 (N_5348,N_3553,N_1999);
nor U5349 (N_5349,N_3142,N_3394);
nor U5350 (N_5350,N_4516,N_819);
nand U5351 (N_5351,N_1627,N_2234);
nand U5352 (N_5352,N_3588,N_3745);
or U5353 (N_5353,N_4109,N_621);
or U5354 (N_5354,N_4862,N_4338);
nor U5355 (N_5355,N_1962,N_3515);
and U5356 (N_5356,N_1266,N_3931);
and U5357 (N_5357,N_1524,N_2910);
and U5358 (N_5358,N_4336,N_162);
nor U5359 (N_5359,N_1046,N_1913);
nand U5360 (N_5360,N_449,N_1042);
nor U5361 (N_5361,N_642,N_990);
and U5362 (N_5362,N_3110,N_929);
and U5363 (N_5363,N_4225,N_755);
or U5364 (N_5364,N_676,N_2937);
nand U5365 (N_5365,N_3228,N_4876);
nor U5366 (N_5366,N_2221,N_3558);
and U5367 (N_5367,N_1517,N_4622);
nand U5368 (N_5368,N_1908,N_4235);
or U5369 (N_5369,N_2699,N_2393);
and U5370 (N_5370,N_564,N_2180);
or U5371 (N_5371,N_619,N_3686);
and U5372 (N_5372,N_2407,N_2546);
nand U5373 (N_5373,N_876,N_1905);
or U5374 (N_5374,N_4569,N_2428);
nand U5375 (N_5375,N_1942,N_1770);
and U5376 (N_5376,N_1616,N_2559);
nand U5377 (N_5377,N_540,N_786);
nor U5378 (N_5378,N_345,N_2696);
nand U5379 (N_5379,N_1093,N_4682);
nand U5380 (N_5380,N_3404,N_1006);
nand U5381 (N_5381,N_1681,N_2624);
or U5382 (N_5382,N_4875,N_1151);
nand U5383 (N_5383,N_3039,N_3983);
and U5384 (N_5384,N_2,N_4106);
nand U5385 (N_5385,N_2283,N_3199);
nand U5386 (N_5386,N_3698,N_3088);
or U5387 (N_5387,N_2659,N_1204);
nor U5388 (N_5388,N_1254,N_4924);
nor U5389 (N_5389,N_4555,N_4986);
and U5390 (N_5390,N_862,N_4323);
or U5391 (N_5391,N_2126,N_3056);
nor U5392 (N_5392,N_4769,N_2928);
nor U5393 (N_5393,N_4681,N_2068);
nor U5394 (N_5394,N_2220,N_1625);
nand U5395 (N_5395,N_1486,N_1883);
or U5396 (N_5396,N_4204,N_4400);
nor U5397 (N_5397,N_1250,N_1816);
nand U5398 (N_5398,N_4344,N_1988);
or U5399 (N_5399,N_3657,N_2750);
and U5400 (N_5400,N_3064,N_1400);
and U5401 (N_5401,N_2537,N_4540);
nor U5402 (N_5402,N_770,N_751);
or U5403 (N_5403,N_2352,N_4821);
or U5404 (N_5404,N_396,N_1430);
nand U5405 (N_5405,N_1900,N_1626);
and U5406 (N_5406,N_844,N_4346);
nand U5407 (N_5407,N_3673,N_628);
and U5408 (N_5408,N_2400,N_3229);
nor U5409 (N_5409,N_3683,N_4708);
nand U5410 (N_5410,N_2851,N_1805);
nand U5411 (N_5411,N_4104,N_2319);
nand U5412 (N_5412,N_4214,N_4465);
and U5413 (N_5413,N_1651,N_2385);
or U5414 (N_5414,N_367,N_1994);
or U5415 (N_5415,N_2878,N_4426);
nand U5416 (N_5416,N_4231,N_4978);
and U5417 (N_5417,N_1555,N_3267);
or U5418 (N_5418,N_4811,N_4);
or U5419 (N_5419,N_207,N_1272);
or U5420 (N_5420,N_976,N_7);
xor U5421 (N_5421,N_185,N_8);
nor U5422 (N_5422,N_3559,N_3173);
or U5423 (N_5423,N_1732,N_2841);
nor U5424 (N_5424,N_3902,N_1649);
or U5425 (N_5425,N_1507,N_1426);
and U5426 (N_5426,N_614,N_2444);
nand U5427 (N_5427,N_754,N_202);
and U5428 (N_5428,N_1071,N_3481);
and U5429 (N_5429,N_458,N_1239);
or U5430 (N_5430,N_607,N_4670);
nand U5431 (N_5431,N_2651,N_803);
or U5432 (N_5432,N_3860,N_1143);
nand U5433 (N_5433,N_1986,N_2408);
nor U5434 (N_5434,N_57,N_2804);
and U5435 (N_5435,N_1855,N_4766);
nand U5436 (N_5436,N_1674,N_4298);
or U5437 (N_5437,N_4091,N_3627);
and U5438 (N_5438,N_954,N_3156);
nor U5439 (N_5439,N_430,N_4935);
or U5440 (N_5440,N_2893,N_3578);
and U5441 (N_5441,N_1480,N_668);
or U5442 (N_5442,N_4056,N_2679);
nor U5443 (N_5443,N_4384,N_2583);
nand U5444 (N_5444,N_4625,N_3572);
nor U5445 (N_5445,N_3384,N_3573);
nand U5446 (N_5446,N_2168,N_4038);
and U5447 (N_5447,N_3255,N_4830);
nor U5448 (N_5448,N_4671,N_1562);
nor U5449 (N_5449,N_3223,N_3337);
nor U5450 (N_5450,N_18,N_1180);
and U5451 (N_5451,N_2227,N_1201);
nand U5452 (N_5452,N_3073,N_3785);
or U5453 (N_5453,N_1116,N_4866);
nor U5454 (N_5454,N_4162,N_4877);
nand U5455 (N_5455,N_981,N_2320);
and U5456 (N_5456,N_4535,N_1576);
or U5457 (N_5457,N_4630,N_3886);
nor U5458 (N_5458,N_556,N_774);
or U5459 (N_5459,N_2230,N_4152);
and U5460 (N_5460,N_4011,N_4915);
and U5461 (N_5461,N_4939,N_2532);
and U5462 (N_5462,N_3442,N_1801);
or U5463 (N_5463,N_4134,N_1063);
or U5464 (N_5464,N_2103,N_2446);
nor U5465 (N_5465,N_4581,N_2643);
nor U5466 (N_5466,N_3342,N_4438);
nor U5467 (N_5467,N_600,N_3571);
nand U5468 (N_5468,N_1877,N_1973);
nor U5469 (N_5469,N_4913,N_932);
and U5470 (N_5470,N_1109,N_4649);
and U5471 (N_5471,N_1868,N_4840);
nor U5472 (N_5472,N_2774,N_471);
nor U5473 (N_5473,N_2287,N_1411);
nand U5474 (N_5474,N_4349,N_4236);
or U5475 (N_5475,N_861,N_1479);
or U5476 (N_5476,N_3327,N_828);
and U5477 (N_5477,N_1552,N_416);
or U5478 (N_5478,N_3396,N_3782);
nor U5479 (N_5479,N_4591,N_2597);
or U5480 (N_5480,N_4510,N_667);
nor U5481 (N_5481,N_4290,N_1505);
or U5482 (N_5482,N_2382,N_4774);
nand U5483 (N_5483,N_2258,N_4695);
and U5484 (N_5484,N_1574,N_854);
nand U5485 (N_5485,N_4002,N_3541);
or U5486 (N_5486,N_359,N_3307);
nand U5487 (N_5487,N_2588,N_234);
nand U5488 (N_5488,N_1741,N_4894);
nand U5489 (N_5489,N_3453,N_2460);
or U5490 (N_5490,N_2200,N_114);
and U5491 (N_5491,N_4368,N_4229);
nand U5492 (N_5492,N_597,N_1381);
or U5493 (N_5493,N_3167,N_3871);
nand U5494 (N_5494,N_2396,N_489);
nor U5495 (N_5495,N_4329,N_1467);
or U5496 (N_5496,N_577,N_2617);
and U5497 (N_5497,N_1553,N_4069);
or U5498 (N_5498,N_2580,N_2100);
and U5499 (N_5499,N_199,N_1156);
nand U5500 (N_5500,N_808,N_1090);
or U5501 (N_5501,N_768,N_2442);
nand U5502 (N_5502,N_2945,N_3137);
and U5503 (N_5503,N_3542,N_2256);
nor U5504 (N_5504,N_2006,N_2264);
nand U5505 (N_5505,N_4944,N_273);
nand U5506 (N_5506,N_220,N_2749);
nor U5507 (N_5507,N_978,N_3867);
and U5508 (N_5508,N_4926,N_2729);
or U5509 (N_5509,N_2307,N_2118);
nand U5510 (N_5510,N_942,N_1163);
nor U5511 (N_5511,N_4301,N_4195);
or U5512 (N_5512,N_3214,N_4754);
and U5513 (N_5513,N_4283,N_4778);
and U5514 (N_5514,N_3777,N_3448);
nor U5515 (N_5515,N_2599,N_2088);
or U5516 (N_5516,N_4975,N_1506);
nor U5517 (N_5517,N_1628,N_2133);
xor U5518 (N_5518,N_1539,N_514);
or U5519 (N_5519,N_2001,N_3879);
nor U5520 (N_5520,N_4819,N_1704);
or U5521 (N_5521,N_3598,N_1832);
and U5522 (N_5522,N_4107,N_1587);
nor U5523 (N_5523,N_3428,N_737);
and U5524 (N_5524,N_4959,N_671);
and U5525 (N_5525,N_344,N_2023);
nor U5526 (N_5526,N_4886,N_1308);
nand U5527 (N_5527,N_2119,N_242);
or U5528 (N_5528,N_3825,N_393);
nand U5529 (N_5529,N_433,N_4454);
nor U5530 (N_5530,N_2826,N_3817);
nand U5531 (N_5531,N_2045,N_659);
nand U5532 (N_5532,N_3200,N_1957);
nor U5533 (N_5533,N_120,N_2678);
nor U5534 (N_5534,N_1699,N_12);
and U5535 (N_5535,N_2175,N_475);
nand U5536 (N_5536,N_3126,N_641);
xnor U5537 (N_5537,N_814,N_3552);
or U5538 (N_5538,N_3466,N_3034);
and U5539 (N_5539,N_3046,N_1072);
nand U5540 (N_5540,N_3646,N_4946);
nor U5541 (N_5541,N_4717,N_1290);
and U5542 (N_5542,N_4224,N_9);
and U5543 (N_5543,N_2509,N_2629);
nor U5544 (N_5544,N_2991,N_940);
nor U5545 (N_5545,N_1548,N_69);
and U5546 (N_5546,N_4136,N_4083);
nand U5547 (N_5547,N_203,N_1504);
nor U5548 (N_5548,N_2677,N_496);
or U5549 (N_5549,N_2563,N_1473);
and U5550 (N_5550,N_2158,N_2403);
nor U5551 (N_5551,N_738,N_4621);
or U5552 (N_5552,N_4583,N_1341);
and U5553 (N_5553,N_4037,N_459);
or U5554 (N_5554,N_3424,N_4963);
and U5555 (N_5555,N_2199,N_1096);
or U5556 (N_5556,N_1434,N_2104);
nor U5557 (N_5557,N_4305,N_4692);
and U5558 (N_5558,N_3719,N_4267);
and U5559 (N_5559,N_228,N_60);
or U5560 (N_5560,N_3135,N_2500);
nand U5561 (N_5561,N_3786,N_336);
nor U5562 (N_5562,N_2974,N_4420);
or U5563 (N_5563,N_4704,N_3557);
or U5564 (N_5564,N_3769,N_2856);
nand U5565 (N_5565,N_1159,N_398);
nor U5566 (N_5566,N_3600,N_2946);
or U5567 (N_5567,N_3740,N_534);
nor U5568 (N_5568,N_3429,N_2998);
and U5569 (N_5569,N_1022,N_1249);
and U5570 (N_5570,N_1644,N_4665);
or U5571 (N_5571,N_4714,N_611);
or U5572 (N_5572,N_402,N_2358);
and U5573 (N_5573,N_4018,N_1692);
and U5574 (N_5574,N_3520,N_4192);
or U5575 (N_5575,N_646,N_1015);
and U5576 (N_5576,N_630,N_2086);
or U5577 (N_5577,N_4520,N_28);
or U5578 (N_5578,N_4078,N_3922);
or U5579 (N_5579,N_2415,N_4327);
or U5580 (N_5580,N_2568,N_2453);
or U5581 (N_5581,N_1002,N_3455);
and U5582 (N_5582,N_3966,N_294);
or U5583 (N_5583,N_3934,N_2556);
and U5584 (N_5584,N_1876,N_1396);
or U5585 (N_5585,N_2832,N_2853);
or U5586 (N_5586,N_4683,N_4750);
nor U5587 (N_5587,N_2432,N_2751);
nor U5588 (N_5588,N_3888,N_4870);
nor U5589 (N_5589,N_3266,N_3193);
and U5590 (N_5590,N_3162,N_2170);
and U5591 (N_5591,N_1526,N_4310);
nor U5592 (N_5592,N_3940,N_2331);
and U5593 (N_5593,N_2115,N_3059);
and U5594 (N_5594,N_2187,N_3722);
or U5595 (N_5595,N_3734,N_4767);
or U5596 (N_5596,N_4489,N_2920);
and U5597 (N_5597,N_1469,N_3620);
nor U5598 (N_5598,N_1189,N_4552);
or U5599 (N_5599,N_3205,N_1767);
nand U5600 (N_5600,N_4369,N_4291);
nor U5601 (N_5601,N_4003,N_4072);
or U5602 (N_5602,N_4131,N_2970);
nand U5603 (N_5603,N_194,N_2165);
xor U5604 (N_5604,N_4196,N_2071);
nand U5605 (N_5605,N_4860,N_3604);
or U5606 (N_5606,N_2476,N_3347);
nand U5607 (N_5607,N_463,N_50);
nand U5608 (N_5608,N_2867,N_4350);
or U5609 (N_5609,N_4220,N_4242);
and U5610 (N_5610,N_4257,N_2269);
nor U5611 (N_5611,N_4917,N_1596);
or U5612 (N_5612,N_2968,N_4567);
or U5613 (N_5613,N_3531,N_455);
and U5614 (N_5614,N_4150,N_2735);
and U5615 (N_5615,N_3812,N_3227);
or U5616 (N_5616,N_3257,N_601);
nand U5617 (N_5617,N_3166,N_1299);
nor U5618 (N_5618,N_2728,N_262);
nor U5619 (N_5619,N_1858,N_2485);
and U5620 (N_5620,N_1735,N_4253);
or U5621 (N_5621,N_899,N_2299);
or U5622 (N_5622,N_1260,N_553);
nand U5623 (N_5623,N_1594,N_4060);
nand U5624 (N_5624,N_4968,N_2543);
or U5625 (N_5625,N_1709,N_4176);
or U5626 (N_5626,N_2569,N_3209);
and U5627 (N_5627,N_3570,N_4922);
nor U5628 (N_5628,N_4851,N_1048);
nor U5629 (N_5629,N_3123,N_4789);
nor U5630 (N_5630,N_4859,N_3181);
nor U5631 (N_5631,N_2669,N_4164);
and U5632 (N_5632,N_1455,N_4703);
nand U5633 (N_5633,N_235,N_3695);
nor U5634 (N_5634,N_1364,N_900);
and U5635 (N_5635,N_2477,N_2334);
nand U5636 (N_5636,N_3801,N_4112);
nor U5637 (N_5637,N_903,N_2364);
and U5638 (N_5638,N_3611,N_2026);
nor U5639 (N_5639,N_2552,N_4473);
nor U5640 (N_5640,N_2257,N_337);
or U5641 (N_5641,N_4780,N_895);
and U5642 (N_5642,N_2069,N_3916);
and U5643 (N_5643,N_2566,N_2876);
nand U5644 (N_5644,N_4010,N_2756);
and U5645 (N_5645,N_2095,N_538);
nor U5646 (N_5646,N_62,N_1117);
or U5647 (N_5647,N_3844,N_4478);
and U5648 (N_5648,N_3744,N_3596);
nor U5649 (N_5649,N_4509,N_4119);
nor U5650 (N_5650,N_4386,N_2399);
and U5651 (N_5651,N_4122,N_2024);
nor U5652 (N_5652,N_665,N_613);
or U5653 (N_5653,N_3731,N_1347);
and U5654 (N_5654,N_956,N_2161);
or U5655 (N_5655,N_2034,N_3677);
nand U5656 (N_5656,N_4477,N_3340);
or U5657 (N_5657,N_1796,N_4161);
nor U5658 (N_5658,N_1113,N_3811);
nor U5659 (N_5659,N_3304,N_707);
nor U5660 (N_5660,N_4009,N_1191);
nand U5661 (N_5661,N_1172,N_2725);
or U5662 (N_5662,N_1803,N_662);
and U5663 (N_5663,N_4139,N_975);
nor U5664 (N_5664,N_2388,N_1719);
and U5665 (N_5665,N_2695,N_848);
or U5666 (N_5666,N_2208,N_3514);
or U5667 (N_5667,N_3547,N_1228);
nor U5668 (N_5668,N_1397,N_2934);
nand U5669 (N_5669,N_2838,N_541);
or U5670 (N_5670,N_3784,N_1044);
nand U5671 (N_5671,N_4004,N_3610);
and U5672 (N_5672,N_1738,N_2229);
nor U5673 (N_5673,N_1461,N_752);
nor U5674 (N_5674,N_1559,N_2602);
xnor U5675 (N_5675,N_847,N_4585);
nand U5676 (N_5676,N_624,N_423);
nor U5677 (N_5677,N_3194,N_2890);
nor U5678 (N_5678,N_2093,N_2365);
nor U5679 (N_5679,N_4184,N_3935);
and U5680 (N_5680,N_497,N_1666);
or U5681 (N_5681,N_1683,N_4451);
nor U5682 (N_5682,N_241,N_2275);
and U5683 (N_5683,N_2724,N_2356);
nor U5684 (N_5684,N_2326,N_2029);
nand U5685 (N_5685,N_964,N_3170);
and U5686 (N_5686,N_2763,N_4123);
nor U5687 (N_5687,N_3368,N_2652);
or U5688 (N_5688,N_4088,N_3467);
nand U5689 (N_5689,N_2816,N_2662);
and U5690 (N_5690,N_2630,N_1529);
nor U5691 (N_5691,N_4912,N_2654);
nor U5692 (N_5692,N_3642,N_1521);
nand U5693 (N_5693,N_1056,N_1487);
or U5694 (N_5694,N_381,N_2670);
xor U5695 (N_5695,N_1050,N_1409);
or U5696 (N_5696,N_1436,N_1328);
nor U5697 (N_5697,N_2251,N_1593);
nor U5698 (N_5698,N_3387,N_1120);
nand U5699 (N_5699,N_4594,N_4702);
nor U5700 (N_5700,N_4210,N_104);
and U5701 (N_5701,N_3765,N_1921);
nor U5702 (N_5702,N_327,N_4281);
or U5703 (N_5703,N_3721,N_3348);
and U5704 (N_5704,N_3955,N_1040);
or U5705 (N_5705,N_1863,N_4713);
nand U5706 (N_5706,N_0,N_4981);
nand U5707 (N_5707,N_3533,N_4410);
and U5708 (N_5708,N_1620,N_4117);
or U5709 (N_5709,N_3846,N_3360);
and U5710 (N_5710,N_153,N_419);
and U5711 (N_5711,N_2268,N_4263);
and U5712 (N_5712,N_1604,N_2869);
nor U5713 (N_5713,N_521,N_4920);
or U5714 (N_5714,N_121,N_3016);
nor U5715 (N_5715,N_2562,N_1813);
nor U5716 (N_5716,N_366,N_2201);
and U5717 (N_5717,N_4554,N_1878);
or U5718 (N_5718,N_2644,N_1373);
nand U5719 (N_5719,N_267,N_119);
and U5720 (N_5720,N_2092,N_1819);
or U5721 (N_5721,N_192,N_796);
nor U5722 (N_5722,N_4800,N_3501);
nor U5723 (N_5723,N_67,N_34);
xnor U5724 (N_5724,N_4299,N_2123);
nand U5725 (N_5725,N_4565,N_3152);
or U5726 (N_5726,N_1095,N_252);
and U5727 (N_5727,N_1634,N_3823);
nor U5728 (N_5728,N_4171,N_4447);
or U5729 (N_5729,N_1874,N_4379);
or U5730 (N_5730,N_3534,N_3796);
nand U5731 (N_5731,N_3115,N_148);
nand U5732 (N_5732,N_3277,N_1985);
or U5733 (N_5733,N_439,N_4149);
nand U5734 (N_5734,N_2022,N_175);
nand U5735 (N_5735,N_962,N_3497);
nand U5736 (N_5736,N_351,N_3145);
nand U5737 (N_5737,N_3131,N_3975);
nand U5738 (N_5738,N_4380,N_408);
nor U5739 (N_5739,N_3180,N_4383);
nor U5740 (N_5740,N_3543,N_3187);
nor U5741 (N_5741,N_493,N_3042);
nand U5742 (N_5742,N_1794,N_4395);
or U5743 (N_5743,N_1271,N_3768);
nor U5744 (N_5744,N_1869,N_1243);
nand U5745 (N_5745,N_1969,N_4320);
and U5746 (N_5746,N_3080,N_3603);
or U5747 (N_5747,N_1641,N_361);
and U5748 (N_5748,N_123,N_3104);
and U5749 (N_5749,N_3890,N_4833);
nor U5750 (N_5750,N_4464,N_4146);
and U5751 (N_5751,N_3416,N_1439);
nor U5752 (N_5752,N_2738,N_254);
or U5753 (N_5753,N_5,N_1851);
nand U5754 (N_5754,N_3421,N_4544);
nand U5755 (N_5755,N_2999,N_1303);
nor U5756 (N_5756,N_2637,N_4937);
and U5757 (N_5757,N_1997,N_269);
nor U5758 (N_5758,N_368,N_4883);
or U5759 (N_5759,N_2622,N_2341);
nand U5760 (N_5760,N_3226,N_3119);
or U5761 (N_5761,N_3196,N_3213);
nor U5762 (N_5762,N_3305,N_3212);
nand U5763 (N_5763,N_502,N_92);
or U5764 (N_5764,N_4574,N_499);
nor U5765 (N_5765,N_712,N_1351);
nor U5766 (N_5766,N_1478,N_2292);
and U5767 (N_5767,N_4275,N_3756);
or U5768 (N_5768,N_3318,N_4311);
nand U5769 (N_5769,N_778,N_1246);
nand U5770 (N_5770,N_3215,N_2301);
or U5771 (N_5771,N_4497,N_746);
nor U5772 (N_5772,N_1789,N_3402);
or U5773 (N_5773,N_3276,N_2947);
or U5774 (N_5774,N_1573,N_1535);
xnor U5775 (N_5775,N_2143,N_4928);
nand U5776 (N_5776,N_2815,N_276);
and U5777 (N_5777,N_4626,N_215);
or U5778 (N_5778,N_1992,N_4007);
nor U5779 (N_5779,N_733,N_2907);
or U5780 (N_5780,N_4730,N_1955);
xor U5781 (N_5781,N_3539,N_4304);
and U5782 (N_5782,N_295,N_2215);
or U5783 (N_5783,N_1797,N_4051);
and U5784 (N_5784,N_3748,N_2855);
nand U5785 (N_5785,N_2317,N_874);
or U5786 (N_5786,N_3292,N_686);
and U5787 (N_5787,N_4015,N_2153);
nand U5788 (N_5788,N_2090,N_3851);
nand U5789 (N_5789,N_3863,N_1181);
or U5790 (N_5790,N_585,N_3766);
and U5791 (N_5791,N_958,N_2730);
nor U5792 (N_5792,N_1638,N_3946);
and U5793 (N_5793,N_945,N_3465);
and U5794 (N_5794,N_3052,N_1483);
nand U5795 (N_5795,N_231,N_3143);
and U5796 (N_5796,N_1852,N_2726);
nand U5797 (N_5797,N_2545,N_784);
and U5798 (N_5798,N_2745,N_1371);
and U5799 (N_5799,N_4590,N_937);
nand U5800 (N_5800,N_919,N_3252);
nor U5801 (N_5801,N_4992,N_3788);
nor U5802 (N_5802,N_1897,N_2064);
and U5803 (N_5803,N_2265,N_2421);
and U5804 (N_5804,N_3184,N_1198);
nand U5805 (N_5805,N_3702,N_1317);
nor U5806 (N_5806,N_4836,N_1178);
or U5807 (N_5807,N_973,N_948);
nand U5808 (N_5808,N_4616,N_1361);
nand U5809 (N_5809,N_700,N_3282);
and U5810 (N_5810,N_2305,N_2081);
and U5811 (N_5811,N_2909,N_431);
or U5812 (N_5812,N_1934,N_3874);
nor U5813 (N_5813,N_110,N_3415);
nor U5814 (N_5814,N_4852,N_3757);
nand U5815 (N_5815,N_4869,N_4994);
nor U5816 (N_5816,N_4317,N_4296);
or U5817 (N_5817,N_1632,N_4958);
or U5818 (N_5818,N_364,N_4764);
nand U5819 (N_5819,N_282,N_4133);
nor U5820 (N_5820,N_1004,N_1825);
xnor U5821 (N_5821,N_1760,N_687);
nand U5822 (N_5822,N_1462,N_2997);
and U5823 (N_5823,N_77,N_2938);
or U5824 (N_5824,N_1387,N_3458);
nand U5825 (N_5825,N_1640,N_3662);
and U5826 (N_5826,N_1932,N_3750);
and U5827 (N_5827,N_3729,N_2181);
nand U5828 (N_5828,N_2983,N_3357);
or U5829 (N_5829,N_4399,N_3449);
and U5830 (N_5830,N_469,N_1772);
or U5831 (N_5831,N_3095,N_869);
and U5832 (N_5832,N_1099,N_2564);
nor U5833 (N_5833,N_320,N_2881);
and U5834 (N_5834,N_2329,N_33);
nor U5835 (N_5835,N_797,N_1687);
and U5836 (N_5836,N_761,N_4905);
nor U5837 (N_5837,N_3147,N_2495);
nor U5838 (N_5838,N_3278,N_4254);
nor U5839 (N_5839,N_3242,N_2057);
and U5840 (N_5840,N_2612,N_98);
nor U5841 (N_5841,N_3417,N_4971);
nand U5842 (N_5842,N_739,N_422);
nand U5843 (N_5843,N_1533,N_2585);
nand U5844 (N_5844,N_1717,N_2744);
nor U5845 (N_5845,N_1319,N_2337);
nand U5846 (N_5846,N_3637,N_4788);
and U5847 (N_5847,N_68,N_1460);
nand U5848 (N_5848,N_237,N_3422);
nand U5849 (N_5849,N_1311,N_3619);
nor U5850 (N_5850,N_840,N_3528);
nor U5851 (N_5851,N_285,N_3040);
nand U5852 (N_5852,N_3928,N_2839);
nor U5853 (N_5853,N_2210,N_3693);
nor U5854 (N_5854,N_1970,N_4167);
nor U5855 (N_5855,N_2128,N_1136);
and U5856 (N_5856,N_4000,N_3701);
nand U5857 (N_5857,N_2941,N_4264);
and U5858 (N_5858,N_4736,N_1543);
nor U5859 (N_5859,N_97,N_1654);
and U5860 (N_5860,N_1684,N_1437);
nor U5861 (N_5861,N_38,N_2214);
nor U5862 (N_5862,N_3669,N_960);
nand U5863 (N_5863,N_3979,N_4720);
and U5864 (N_5864,N_4553,N_4942);
or U5865 (N_5865,N_4306,N_2919);
and U5866 (N_5866,N_2688,N_4398);
and U5867 (N_5867,N_1368,N_4728);
or U5868 (N_5868,N_4743,N_1277);
and U5869 (N_5869,N_879,N_2958);
nor U5870 (N_5870,N_1743,N_4543);
and U5871 (N_5871,N_4498,N_4218);
or U5872 (N_5872,N_1952,N_4634);
and U5873 (N_5873,N_3499,N_2311);
or U5874 (N_5874,N_1882,N_126);
nor U5875 (N_5875,N_1173,N_1468);
and U5876 (N_5876,N_1025,N_2192);
or U5877 (N_5877,N_1648,N_255);
xor U5878 (N_5878,N_4960,N_4058);
nand U5879 (N_5879,N_1785,N_1196);
or U5880 (N_5880,N_2747,N_892);
nor U5881 (N_5881,N_186,N_3965);
or U5882 (N_5882,N_3936,N_1592);
nor U5883 (N_5883,N_2734,N_734);
and U5884 (N_5884,N_1268,N_2732);
nor U5885 (N_5885,N_4753,N_3589);
xnor U5886 (N_5886,N_2140,N_1378);
nor U5887 (N_5887,N_554,N_2423);
nor U5888 (N_5888,N_822,N_2880);
nand U5889 (N_5889,N_4365,N_1589);
nand U5890 (N_5890,N_3771,N_2222);
nor U5891 (N_5891,N_3633,N_2427);
and U5892 (N_5892,N_4103,N_1689);
or U5893 (N_5893,N_810,N_1933);
or U5894 (N_5894,N_3525,N_1255);
or U5895 (N_5895,N_4325,N_4834);
nand U5896 (N_5896,N_143,N_3300);
and U5897 (N_5897,N_2085,N_4159);
and U5898 (N_5898,N_1907,N_3063);
and U5899 (N_5899,N_2835,N_467);
and U5900 (N_5900,N_1135,N_4951);
or U5901 (N_5901,N_3195,N_1971);
and U5902 (N_5902,N_827,N_2940);
or U5903 (N_5903,N_3858,N_328);
or U5904 (N_5904,N_4316,N_4111);
and U5905 (N_5905,N_66,N_3343);
and U5906 (N_5906,N_3349,N_991);
and U5907 (N_5907,N_817,N_2286);
and U5908 (N_5908,N_3057,N_1761);
and U5909 (N_5909,N_2340,N_3316);
or U5910 (N_5910,N_4370,N_1508);
nand U5911 (N_5911,N_3105,N_440);
nand U5912 (N_5912,N_4962,N_2573);
nand U5913 (N_5913,N_1211,N_503);
nand U5914 (N_5914,N_2987,N_510);
nor U5915 (N_5915,N_1450,N_239);
nand U5916 (N_5916,N_2277,N_1421);
nor U5917 (N_5917,N_1827,N_3291);
or U5918 (N_5918,N_689,N_3077);
and U5919 (N_5919,N_1306,N_757);
and U5920 (N_5920,N_2926,N_2589);
and U5921 (N_5921,N_1406,N_2955);
or U5922 (N_5922,N_2702,N_4848);
nor U5923 (N_5923,N_1937,N_4087);
nand U5924 (N_5924,N_4933,N_842);
or U5925 (N_5925,N_3741,N_2687);
nor U5926 (N_5926,N_461,N_1494);
or U5927 (N_5927,N_3198,N_4013);
and U5928 (N_5928,N_1348,N_3028);
or U5929 (N_5929,N_181,N_3390);
or U5930 (N_5930,N_350,N_3706);
nand U5931 (N_5931,N_1606,N_428);
nor U5932 (N_5932,N_917,N_2582);
and U5933 (N_5933,N_3395,N_838);
or U5934 (N_5934,N_3287,N_867);
and U5935 (N_5935,N_787,N_2591);
and U5936 (N_5936,N_2716,N_2795);
and U5937 (N_5937,N_2130,N_48);
or U5938 (N_5938,N_4394,N_4577);
nand U5939 (N_5939,N_993,N_2102);
nor U5940 (N_5940,N_1061,N_4001);
and U5941 (N_5941,N_1670,N_1636);
or U5942 (N_5942,N_4511,N_1577);
nor U5943 (N_5943,N_1840,N_637);
nand U5944 (N_5944,N_4524,N_2697);
and U5945 (N_5945,N_3774,N_2665);
nand U5946 (N_5946,N_3852,N_1991);
and U5947 (N_5947,N_1575,N_2015);
nor U5948 (N_5948,N_409,N_1016);
nand U5949 (N_5949,N_809,N_2967);
nor U5950 (N_5950,N_4648,N_2473);
nor U5951 (N_5951,N_4631,N_1845);
or U5952 (N_5952,N_1580,N_3624);
nor U5953 (N_5953,N_1346,N_4315);
or U5954 (N_5954,N_833,N_3651);
and U5955 (N_5955,N_959,N_3606);
and U5956 (N_5956,N_4138,N_4280);
nand U5957 (N_5957,N_2526,N_1864);
nand U5958 (N_5958,N_1231,N_4309);
or U5959 (N_5959,N_3690,N_22);
nand U5960 (N_5960,N_1399,N_3010);
or U5961 (N_5961,N_4198,N_2904);
nor U5962 (N_5962,N_3355,N_1212);
nand U5963 (N_5963,N_132,N_2191);
or U5964 (N_5964,N_1009,N_4801);
or U5965 (N_5965,N_4424,N_2386);
and U5966 (N_5966,N_1264,N_3153);
nor U5967 (N_5967,N_4374,N_2209);
or U5968 (N_5968,N_2733,N_2055);
or U5969 (N_5969,N_4953,N_968);
nand U5970 (N_5970,N_3302,N_2070);
or U5971 (N_5971,N_1017,N_1982);
or U5972 (N_5972,N_3489,N_4619);
nor U5973 (N_5973,N_1028,N_4900);
and U5974 (N_5974,N_4651,N_2430);
nand U5975 (N_5975,N_1193,N_1682);
and U5976 (N_5976,N_3386,N_1525);
xor U5977 (N_5977,N_1513,N_2694);
and U5978 (N_5978,N_1220,N_1088);
and U5979 (N_5979,N_552,N_1309);
and U5980 (N_5980,N_4188,N_2318);
nand U5981 (N_5981,N_4620,N_972);
nor U5982 (N_5982,N_3430,N_2596);
and U5983 (N_5983,N_1234,N_4243);
or U5984 (N_5984,N_1333,N_4412);
nor U5985 (N_5985,N_2226,N_279);
and U5986 (N_5986,N_1005,N_901);
nand U5987 (N_5987,N_3875,N_2718);
nand U5988 (N_5988,N_2975,N_1901);
or U5989 (N_5989,N_1829,N_4781);
nand U5990 (N_5990,N_1357,N_338);
nand U5991 (N_5991,N_415,N_1481);
nor U5992 (N_5992,N_3670,N_4599);
or U5993 (N_5993,N_65,N_4121);
nor U5994 (N_5994,N_2866,N_790);
nor U5995 (N_5995,N_2779,N_3151);
nor U5996 (N_5996,N_335,N_3555);
and U5997 (N_5997,N_4603,N_888);
nor U5998 (N_5998,N_3090,N_372);
or U5999 (N_5999,N_4573,N_4312);
or U6000 (N_6000,N_3685,N_565);
nand U6001 (N_6001,N_579,N_1523);
or U6002 (N_6002,N_1866,N_4502);
and U6003 (N_6003,N_208,N_281);
or U6004 (N_6004,N_4950,N_974);
or U6005 (N_6005,N_4940,N_387);
and U6006 (N_6006,N_4055,N_342);
nor U6007 (N_6007,N_4664,N_4934);
or U6008 (N_6008,N_3661,N_946);
and U6009 (N_6009,N_310,N_52);
and U6010 (N_6010,N_1727,N_4227);
or U6011 (N_6011,N_532,N_4863);
or U6012 (N_6012,N_4999,N_1622);
and U6013 (N_6013,N_4493,N_3364);
nor U6014 (N_6014,N_558,N_4297);
and U6015 (N_6015,N_3418,N_697);
nand U6016 (N_6016,N_3082,N_2420);
and U6017 (N_6017,N_3306,N_1998);
nand U6018 (N_6018,N_727,N_4155);
nor U6019 (N_6019,N_2082,N_4328);
and U6020 (N_6020,N_4163,N_2900);
nor U6021 (N_6021,N_2371,N_1953);
and U6022 (N_6022,N_3179,N_4672);
and U6023 (N_6023,N_4729,N_557);
nor U6024 (N_6024,N_217,N_1938);
or U6025 (N_6025,N_191,N_3248);
nor U6026 (N_6026,N_1464,N_2993);
nand U6027 (N_6027,N_804,N_1987);
or U6028 (N_6028,N_293,N_736);
xnor U6029 (N_6029,N_3218,N_4491);
nor U6030 (N_6030,N_3241,N_3388);
nor U6031 (N_6031,N_3508,N_1875);
nor U6032 (N_6032,N_4637,N_530);
and U6033 (N_6033,N_2493,N_2506);
nor U6034 (N_6034,N_4307,N_2194);
xor U6035 (N_6035,N_2302,N_2534);
and U6036 (N_6036,N_4784,N_4677);
or U6037 (N_6037,N_3491,N_2387);
nor U6038 (N_6038,N_4429,N_997);
and U6039 (N_6039,N_4197,N_4401);
nor U6040 (N_6040,N_3751,N_857);
nand U6041 (N_6041,N_76,N_1292);
nor U6042 (N_6042,N_1188,N_4486);
nand U6043 (N_6043,N_4804,N_4282);
nand U6044 (N_6044,N_699,N_1297);
nand U6045 (N_6045,N_4533,N_3281);
nor U6046 (N_6046,N_4678,N_2261);
nand U6047 (N_6047,N_609,N_2770);
nor U6048 (N_6048,N_4406,N_391);
and U6049 (N_6049,N_2004,N_257);
and U6050 (N_6050,N_3319,N_4090);
nand U6051 (N_6051,N_4470,N_4028);
nor U6052 (N_6052,N_1304,N_2803);
and U6053 (N_6053,N_740,N_182);
or U6054 (N_6054,N_2467,N_4173);
nor U6055 (N_6055,N_3154,N_4348);
or U6056 (N_6056,N_348,N_240);
nand U6057 (N_6057,N_4892,N_2372);
and U6058 (N_6058,N_10,N_380);
or U6059 (N_6059,N_4022,N_3211);
or U6060 (N_6060,N_3120,N_3530);
or U6061 (N_6061,N_930,N_2469);
and U6062 (N_6062,N_1241,N_811);
and U6063 (N_6063,N_560,N_4615);
nand U6064 (N_6064,N_3628,N_4995);
nor U6065 (N_6065,N_3178,N_1202);
or U6066 (N_6066,N_3933,N_2603);
or U6067 (N_6067,N_1854,N_545);
xor U6068 (N_6068,N_2479,N_168);
nand U6069 (N_6069,N_3708,N_4347);
nand U6070 (N_6070,N_3013,N_1463);
and U6071 (N_6071,N_4831,N_3072);
and U6072 (N_6072,N_151,N_72);
and U6073 (N_6073,N_1168,N_4527);
and U6074 (N_6074,N_2700,N_2263);
nor U6075 (N_6075,N_4700,N_3783);
or U6076 (N_6076,N_2772,N_3631);
nor U6077 (N_6077,N_1150,N_3204);
or U6078 (N_6078,N_966,N_2542);
or U6079 (N_6079,N_2193,N_212);
or U6080 (N_6080,N_4265,N_4673);
and U6081 (N_6081,N_1959,N_3688);
nor U6082 (N_6082,N_2771,N_3261);
nand U6083 (N_6083,N_2042,N_680);
or U6084 (N_6084,N_300,N_1981);
and U6085 (N_6085,N_2009,N_3883);
and U6086 (N_6086,N_3545,N_4528);
or U6087 (N_6087,N_1783,N_1296);
and U6088 (N_6088,N_3314,N_4861);
nor U6089 (N_6089,N_1890,N_4047);
and U6090 (N_6090,N_3739,N_1492);
nand U6091 (N_6091,N_1064,N_2144);
nor U6092 (N_6092,N_2527,N_3759);
nor U6093 (N_6093,N_1612,N_2290);
and U6094 (N_6094,N_886,N_744);
nor U6095 (N_6095,N_4715,N_3615);
nand U6096 (N_6096,N_4558,N_2754);
nand U6097 (N_6097,N_2775,N_1043);
nand U6098 (N_6098,N_1352,N_2461);
and U6099 (N_6099,N_2106,N_432);
nor U6100 (N_6100,N_1126,N_2830);
nand U6101 (N_6101,N_4659,N_340);
and U6102 (N_6102,N_1706,N_2289);
nor U6103 (N_6103,N_201,N_1337);
and U6104 (N_6104,N_1731,N_3632);
and U6105 (N_6105,N_2915,N_1142);
or U6106 (N_6106,N_4045,N_650);
nor U6107 (N_6107,N_898,N_3772);
nand U6108 (N_6108,N_4541,N_816);
nand U6109 (N_6109,N_912,N_1261);
or U6110 (N_6110,N_625,N_323);
nor U6111 (N_6111,N_2895,N_610);
or U6112 (N_6112,N_4442,N_2886);
or U6113 (N_6113,N_2577,N_2472);
nand U6114 (N_6114,N_3258,N_2796);
nand U6115 (N_6115,N_3127,N_3582);
nor U6116 (N_6116,N_574,N_2178);
or U6117 (N_6117,N_96,N_3800);
or U6118 (N_6118,N_4806,N_2378);
and U6119 (N_6119,N_2087,N_3370);
nor U6120 (N_6120,N_1466,N_2518);
and U6121 (N_6121,N_1943,N_3587);
and U6122 (N_6122,N_1456,N_1358);
nor U6123 (N_6123,N_1764,N_3815);
xor U6124 (N_6124,N_205,N_2447);
or U6125 (N_6125,N_2243,N_1053);
nand U6126 (N_6126,N_4460,N_4517);
or U6127 (N_6127,N_2332,N_3454);
and U6128 (N_6128,N_933,N_3076);
nor U6129 (N_6129,N_473,N_594);
nor U6130 (N_6130,N_4450,N_3848);
or U6131 (N_6131,N_2296,N_4761);
or U6132 (N_6132,N_2741,N_4274);
nor U6133 (N_6133,N_3103,N_2120);
nand U6134 (N_6134,N_1301,N_2253);
and U6135 (N_6135,N_2383,N_2244);
nor U6136 (N_6136,N_4156,N_715);
or U6137 (N_6137,N_3838,N_371);
xor U6138 (N_6138,N_1566,N_3714);
or U6139 (N_6139,N_1091,N_1679);
or U6140 (N_6140,N_3993,N_4108);
or U6141 (N_6141,N_2463,N_2047);
or U6142 (N_6142,N_1427,N_3071);
nor U6143 (N_6143,N_331,N_2781);
or U6144 (N_6144,N_1323,N_915);
and U6145 (N_6145,N_3503,N_3309);
or U6146 (N_6146,N_1030,N_2951);
and U6147 (N_6147,N_1676,N_2626);
or U6148 (N_6148,N_3918,N_1435);
nand U6149 (N_6149,N_2019,N_2510);
nand U6150 (N_6150,N_2164,N_298);
nand U6151 (N_6151,N_425,N_4891);
and U6152 (N_6152,N_3253,N_938);
nand U6153 (N_6153,N_1076,N_1765);
nand U6154 (N_6154,N_504,N_3190);
nand U6155 (N_6155,N_1278,N_4006);
or U6156 (N_6156,N_1889,N_4488);
nor U6157 (N_6157,N_3492,N_4191);
nand U6158 (N_6158,N_3780,N_4287);
nor U6159 (N_6159,N_764,N_2246);
nor U6160 (N_6160,N_2655,N_4741);
and U6161 (N_6161,N_3629,N_781);
nand U6162 (N_6162,N_1850,N_4588);
nor U6163 (N_6163,N_218,N_4407);
or U6164 (N_6164,N_1771,N_157);
nand U6165 (N_6165,N_4084,N_2693);
nand U6166 (N_6166,N_4988,N_4919);
nor U6167 (N_6167,N_2760,N_821);
nand U6168 (N_6168,N_1608,N_3371);
nor U6169 (N_6169,N_3155,N_612);
and U6170 (N_6170,N_2717,N_1581);
nor U6171 (N_6171,N_2231,N_4612);
nand U6172 (N_6172,N_4102,N_2723);
nor U6173 (N_6173,N_4748,N_4923);
or U6174 (N_6174,N_4518,N_2985);
or U6175 (N_6175,N_41,N_758);
nand U6176 (N_6176,N_4293,N_4239);
or U6177 (N_6177,N_2828,N_4895);
and U6178 (N_6178,N_272,N_2953);
nor U6179 (N_6179,N_4658,N_3957);
or U6180 (N_6180,N_1716,N_853);
nand U6181 (N_6181,N_4288,N_527);
or U6182 (N_6182,N_2455,N_3864);
or U6183 (N_6183,N_4645,N_698);
nand U6184 (N_6184,N_759,N_2517);
or U6185 (N_6185,N_4822,N_1289);
nor U6186 (N_6186,N_3917,N_4562);
nand U6187 (N_6187,N_3551,N_952);
or U6188 (N_6188,N_1321,N_466);
or U6189 (N_6189,N_3322,N_4636);
or U6190 (N_6190,N_3379,N_695);
nor U6191 (N_6191,N_523,N_3066);
and U6192 (N_6192,N_913,N_4480);
and U6193 (N_6193,N_3012,N_2471);
or U6194 (N_6194,N_2303,N_2146);
and U6195 (N_6195,N_823,N_1815);
and U6196 (N_6196,N_2060,N_4183);
and U6197 (N_6197,N_3107,N_4397);
nor U6198 (N_6198,N_979,N_356);
or U6199 (N_6199,N_4033,N_3506);
nand U6200 (N_6200,N_3617,N_1391);
or U6201 (N_6201,N_3329,N_3495);
and U6202 (N_6202,N_1037,N_1345);
or U6203 (N_6203,N_329,N_2903);
and U6204 (N_6204,N_1390,N_910);
nand U6205 (N_6205,N_164,N_2619);
and U6206 (N_6206,N_2418,N_2044);
nand U6207 (N_6207,N_2766,N_4073);
nand U6208 (N_6208,N_2512,N_4827);
and U6209 (N_6209,N_4716,N_3964);
nor U6210 (N_6210,N_3828,N_4777);
nand U6211 (N_6211,N_3822,N_2376);
or U6212 (N_6212,N_1327,N_2398);
and U6213 (N_6213,N_2906,N_4376);
or U6214 (N_6214,N_1956,N_524);
and U6215 (N_6215,N_219,N_3280);
or U6216 (N_6216,N_4059,N_1281);
or U6217 (N_6217,N_286,N_3820);
nor U6218 (N_6218,N_1560,N_1284);
nor U6219 (N_6219,N_3925,N_3254);
and U6220 (N_6220,N_4479,N_187);
nand U6221 (N_6221,N_2335,N_3452);
and U6222 (N_6222,N_719,N_2884);
or U6223 (N_6223,N_1330,N_4285);
or U6224 (N_6224,N_1376,N_1698);
or U6225 (N_6225,N_3463,N_4213);
nand U6226 (N_6226,N_2605,N_4598);
or U6227 (N_6227,N_849,N_3580);
or U6228 (N_6228,N_2076,N_731);
nor U6229 (N_6229,N_3233,N_4853);
nand U6230 (N_6230,N_4791,N_1111);
and U6231 (N_6231,N_1154,N_2037);
nor U6232 (N_6232,N_3262,N_4402);
nand U6233 (N_6233,N_1069,N_470);
nor U6234 (N_6234,N_55,N_260);
or U6235 (N_6235,N_4050,N_488);
nor U6236 (N_6236,N_1448,N_4901);
nand U6237 (N_6237,N_2218,N_4829);
nand U6238 (N_6238,N_2053,N_4733);
nor U6239 (N_6239,N_1032,N_2381);
nor U6240 (N_6240,N_1010,N_2349);
nor U6241 (N_6241,N_2931,N_596);
nor U6242 (N_6242,N_454,N_4377);
xnor U6243 (N_6243,N_1746,N_4586);
and U6244 (N_6244,N_2581,N_2666);
and U6245 (N_6245,N_3675,N_3148);
nor U6246 (N_6246,N_4143,N_1658);
nor U6247 (N_6247,N_4168,N_3961);
nor U6248 (N_6248,N_4110,N_3197);
nand U6249 (N_6249,N_3504,N_2294);
and U6250 (N_6250,N_669,N_27);
nand U6251 (N_6251,N_2921,N_1424);
and U6252 (N_6252,N_2650,N_4699);
or U6253 (N_6253,N_2041,N_144);
nor U6254 (N_6254,N_79,N_843);
and U6255 (N_6255,N_3808,N_4898);
nor U6256 (N_6256,N_305,N_1329);
or U6257 (N_6257,N_535,N_2113);
and U6258 (N_6258,N_1263,N_4897);
and U6259 (N_6259,N_2005,N_225);
or U6260 (N_6260,N_1055,N_3638);
nor U6261 (N_6261,N_1045,N_934);
or U6262 (N_6262,N_2274,N_615);
nor U6263 (N_6263,N_4906,N_1291);
and U6264 (N_6264,N_4556,N_3891);
nand U6265 (N_6265,N_4284,N_1870);
and U6266 (N_6266,N_321,N_4124);
and U6267 (N_6267,N_4525,N_2188);
nor U6268 (N_6268,N_3397,N_2136);
nor U6269 (N_6269,N_992,N_664);
nor U6270 (N_6270,N_3157,N_4505);
nor U6271 (N_6271,N_2709,N_724);
or U6272 (N_6272,N_297,N_2521);
and U6273 (N_6273,N_4014,N_3399);
or U6274 (N_6274,N_3853,N_3344);
nor U6275 (N_6275,N_2308,N_32);
and U6276 (N_6276,N_3350,N_1083);
nand U6277 (N_6277,N_1749,N_1510);
and U6278 (N_6278,N_3391,N_4993);
or U6279 (N_6279,N_2031,N_1227);
or U6280 (N_6280,N_3408,N_271);
nand U6281 (N_6281,N_1707,N_3696);
and U6282 (N_6282,N_539,N_4031);
and U6283 (N_6283,N_1568,N_1031);
and U6284 (N_6284,N_2392,N_3899);
nand U6285 (N_6285,N_4593,N_550);
nand U6286 (N_6286,N_3003,N_2857);
or U6287 (N_6287,N_3840,N_4873);
and U6288 (N_6288,N_3439,N_4300);
or U6289 (N_6289,N_677,N_1070);
nand U6290 (N_6290,N_1534,N_4039);
or U6291 (N_6291,N_3987,N_4846);
and U6292 (N_6292,N_3907,N_2431);
and U6293 (N_6293,N_3500,N_2606);
nand U6294 (N_6294,N_2740,N_518);
or U6295 (N_6295,N_618,N_3723);
or U6296 (N_6296,N_2189,N_2497);
and U6297 (N_6297,N_1817,N_4245);
nand U6298 (N_6298,N_3845,N_708);
nor U6299 (N_6299,N_3065,N_4669);
or U6300 (N_6300,N_998,N_2413);
nor U6301 (N_6301,N_3813,N_4571);
nor U6302 (N_6302,N_1673,N_4638);
nand U6303 (N_6303,N_4271,N_529);
or U6304 (N_6304,N_1810,N_170);
and U6305 (N_6305,N_1472,N_1958);
nand U6306 (N_6306,N_4787,N_1499);
nand U6307 (N_6307,N_1219,N_3009);
nand U6308 (N_6308,N_4575,N_4247);
nor U6309 (N_6309,N_3793,N_794);
and U6310 (N_6310,N_4931,N_1392);
or U6311 (N_6311,N_1541,N_4698);
nor U6312 (N_6312,N_270,N_3832);
or U6313 (N_6313,N_490,N_2350);
and U6314 (N_6314,N_4602,N_278);
nand U6315 (N_6315,N_4550,N_2584);
and U6316 (N_6316,N_520,N_3716);
and U6317 (N_6317,N_2018,N_4326);
or U6318 (N_6318,N_3967,N_941);
or U6319 (N_6319,N_4817,N_1588);
nor U6320 (N_6320,N_4998,N_3124);
nor U6321 (N_6321,N_1214,N_3540);
and U6322 (N_6322,N_3221,N_3996);
nand U6323 (N_6323,N_1036,N_3954);
or U6324 (N_6324,N_2010,N_4770);
nor U6325 (N_6325,N_1911,N_413);
nand U6326 (N_6326,N_3778,N_4948);
and U6327 (N_6327,N_1482,N_1379);
nor U6328 (N_6328,N_2755,N_1269);
and U6329 (N_6329,N_957,N_2868);
or U6330 (N_6330,N_4153,N_1695);
nor U6331 (N_6331,N_474,N_4234);
nand U6332 (N_6332,N_870,N_1429);
nand U6333 (N_6333,N_4244,N_3482);
and U6334 (N_6334,N_312,N_1979);
and U6335 (N_6335,N_2994,N_35);
nor U6336 (N_6336,N_1074,N_1931);
nor U6337 (N_6337,N_583,N_1954);
or U6338 (N_6338,N_681,N_4723);
or U6339 (N_6339,N_936,N_887);
nor U6340 (N_6340,N_1349,N_3988);
nor U6341 (N_6341,N_4872,N_805);
or U6342 (N_6342,N_1141,N_970);
nand U6343 (N_6343,N_362,N_4680);
and U6344 (N_6344,N_4373,N_526);
nand U6345 (N_6345,N_1844,N_2932);
nand U6346 (N_6346,N_654,N_2731);
or U6347 (N_6347,N_1657,N_4151);
nor U6348 (N_6348,N_3561,N_742);
and U6349 (N_6349,N_3877,N_4475);
nand U6350 (N_6350,N_3569,N_2452);
nor U6351 (N_6351,N_2474,N_1215);
nor U6352 (N_6352,N_4476,N_2295);
nand U6353 (N_6353,N_777,N_3134);
nor U6354 (N_6354,N_788,N_4294);
or U6355 (N_6355,N_1820,N_555);
nand U6356 (N_6356,N_2316,N_1023);
nand U6357 (N_6357,N_462,N_3333);
and U6358 (N_6358,N_1585,N_931);
or U6359 (N_6359,N_184,N_3315);
nand U6360 (N_6360,N_3462,N_3096);
or U6361 (N_6361,N_3426,N_4005);
or U6362 (N_6362,N_863,N_2969);
and U6363 (N_6363,N_2373,N_1477);
nand U6364 (N_6364,N_2360,N_4726);
nand U6365 (N_6365,N_4911,N_1279);
or U6366 (N_6366,N_2040,N_4776);
nand U6367 (N_6367,N_3238,N_2059);
or U6368 (N_6368,N_4684,N_2162);
and U6369 (N_6369,N_4441,N_2824);
nand U6370 (N_6370,N_2663,N_4816);
and U6371 (N_6371,N_476,N_251);
or U6372 (N_6372,N_377,N_3081);
or U6373 (N_6373,N_313,N_1192);
and U6374 (N_6374,N_1350,N_4434);
nand U6375 (N_6375,N_1690,N_4181);
and U6376 (N_6376,N_4857,N_263);
or U6377 (N_6377,N_3208,N_3914);
nor U6378 (N_6378,N_3425,N_3789);
nand U6379 (N_6379,N_3787,N_3083);
nor U6380 (N_6380,N_1872,N_4956);
nor U6381 (N_6381,N_4219,N_3446);
nor U6382 (N_6382,N_581,N_2739);
and U6383 (N_6383,N_1,N_2228);
nand U6384 (N_6384,N_4458,N_500);
nor U6385 (N_6385,N_2712,N_841);
nor U6386 (N_6386,N_4925,N_3203);
nand U6387 (N_6387,N_4354,N_1367);
and U6388 (N_6388,N_370,N_3650);
nor U6389 (N_6389,N_4487,N_2291);
and U6390 (N_6390,N_3790,N_4411);
and U6391 (N_6391,N_2033,N_3250);
or U6392 (N_6392,N_3671,N_4982);
and U6393 (N_6393,N_154,N_1125);
nand U6394 (N_6394,N_4216,N_1404);
and U6395 (N_6395,N_4970,N_3146);
nor U6396 (N_6396,N_1360,N_4481);
nand U6397 (N_6397,N_2896,N_188);
nand U6398 (N_6398,N_2698,N_1190);
and U6399 (N_6399,N_4492,N_4757);
nor U6400 (N_6400,N_4624,N_3367);
nor U6401 (N_6401,N_4093,N_4530);
nand U6402 (N_6402,N_1112,N_3122);
nand U6403 (N_6403,N_3268,N_949);
or U6404 (N_6404,N_2167,N_2362);
and U6405 (N_6405,N_568,N_4471);
and U6406 (N_6406,N_2216,N_1240);
nor U6407 (N_6407,N_2017,N_3889);
or U6408 (N_6408,N_2902,N_399);
nor U6409 (N_6409,N_352,N_1740);
nor U6410 (N_6410,N_2151,N_2159);
or U6411 (N_6411,N_435,N_2924);
nand U6412 (N_6412,N_1881,N_3293);
nand U6413 (N_6413,N_4890,N_3030);
and U6414 (N_6414,N_1910,N_3331);
or U6415 (N_6415,N_4578,N_1153);
and U6416 (N_6416,N_3697,N_1826);
or U6417 (N_6417,N_324,N_1860);
and U6418 (N_6418,N_3007,N_587);
nand U6419 (N_6419,N_2405,N_4408);
and U6420 (N_6420,N_1629,N_4654);
nand U6421 (N_6421,N_1059,N_2462);
nor U6422 (N_6422,N_99,N_2353);
nand U6423 (N_6423,N_767,N_815);
and U6424 (N_6424,N_249,N_2366);
and U6425 (N_6425,N_4779,N_2099);
nor U6426 (N_6426,N_1165,N_4580);
and U6427 (N_6427,N_2809,N_3366);
nand U6428 (N_6428,N_3251,N_3810);
or U6429 (N_6429,N_2822,N_3365);
nand U6430 (N_6430,N_4295,N_1778);
nand U6431 (N_6431,N_1733,N_3239);
or U6432 (N_6432,N_3336,N_389);
nand U6433 (N_6433,N_4663,N_1551);
nor U6434 (N_6434,N_3953,N_709);
nor U6435 (N_6435,N_1186,N_4043);
nand U6436 (N_6436,N_2117,N_1848);
nand U6437 (N_6437,N_636,N_346);
nand U6438 (N_6438,N_1720,N_872);
or U6439 (N_6439,N_1282,N_1511);
nor U6440 (N_6440,N_4343,N_1519);
nor U6441 (N_6441,N_424,N_4653);
and U6442 (N_6442,N_1564,N_1849);
and U6443 (N_6443,N_446,N_3263);
nand U6444 (N_6444,N_1948,N_985);
or U6445 (N_6445,N_448,N_2586);
nand U6446 (N_6446,N_3385,N_4032);
nand U6447 (N_6447,N_2384,N_4850);
nand U6448 (N_6448,N_509,N_1546);
nand U6449 (N_6449,N_2343,N_3369);
nand U6450 (N_6450,N_3298,N_1873);
and U6451 (N_6451,N_325,N_4074);
and U6452 (N_6452,N_4623,N_434);
or U6453 (N_6453,N_2270,N_1708);
and U6454 (N_6454,N_37,N_1887);
or U6455 (N_6455,N_3728,N_1027);
or U6456 (N_6456,N_2616,N_47);
and U6457 (N_6457,N_935,N_4496);
and U6458 (N_6458,N_3639,N_4608);
nor U6459 (N_6459,N_2613,N_2488);
nor U6460 (N_6460,N_392,N_651);
nor U6461 (N_6461,N_174,N_3014);
nand U6462 (N_6462,N_2689,N_1235);
or U6463 (N_6463,N_287,N_813);
nand U6464 (N_6464,N_4017,N_4113);
nand U6465 (N_6465,N_3461,N_54);
and U6466 (N_6466,N_3995,N_4041);
or U6467 (N_6467,N_3727,N_1531);
nor U6468 (N_6468,N_3618,N_4722);
nand U6469 (N_6469,N_3910,N_4519);
nor U6470 (N_6470,N_2894,N_1838);
and U6471 (N_6471,N_2404,N_245);
or U6472 (N_6472,N_2424,N_4375);
and U6473 (N_6473,N_78,N_800);
nor U6474 (N_6474,N_2858,N_3564);
or U6475 (N_6475,N_4302,N_3591);
or U6476 (N_6476,N_3679,N_3243);
or U6477 (N_6477,N_3183,N_705);
nand U6478 (N_6478,N_4790,N_292);
and U6479 (N_6479,N_4114,N_1888);
nor U6480 (N_6480,N_31,N_2142);
and U6481 (N_6481,N_2922,N_4248);
nor U6482 (N_6482,N_3445,N_2914);
or U6483 (N_6483,N_1394,N_1605);
or U6484 (N_6484,N_4095,N_1667);
and U6485 (N_6485,N_3857,N_2703);
nor U6486 (N_6486,N_2610,N_4867);
or U6487 (N_6487,N_4880,N_1183);
or U6488 (N_6488,N_3868,N_3601);
and U6489 (N_6489,N_1503,N_2036);
or U6490 (N_6490,N_3893,N_2885);
or U6491 (N_6491,N_977,N_2727);
nor U6492 (N_6492,N_4061,N_2530);
nand U6493 (N_6493,N_2054,N_859);
or U6494 (N_6494,N_3398,N_2656);
and U6495 (N_6495,N_109,N_1386);
or U6496 (N_6496,N_3689,N_4194);
nor U6497 (N_6497,N_1185,N_1639);
and U6498 (N_6498,N_4824,N_1630);
nor U6499 (N_6499,N_1660,N_284);
nand U6500 (N_6500,N_2127,N_678);
or U6501 (N_6501,N_125,N_785);
and U6502 (N_6502,N_1619,N_3681);
nor U6503 (N_6503,N_3440,N_3485);
nand U6504 (N_6504,N_2782,N_1941);
nor U6505 (N_6505,N_1021,N_1637);
nand U6506 (N_6506,N_3085,N_2916);
or U6507 (N_6507,N_543,N_4141);
nand U6508 (N_6508,N_3517,N_2380);
nor U6509 (N_6509,N_3079,N_386);
nand U6510 (N_6510,N_4983,N_73);
nor U6511 (N_6511,N_1393,N_2439);
or U6512 (N_6512,N_578,N_3438);
or U6513 (N_6513,N_4185,N_2719);
or U6514 (N_6514,N_789,N_2293);
nand U6515 (N_6515,N_1000,N_4885);
nor U6516 (N_6516,N_2807,N_3008);
and U6517 (N_6517,N_2314,N_4086);
and U6518 (N_6518,N_2248,N_4826);
or U6519 (N_6519,N_1104,N_3378);
nand U6520 (N_6520,N_2183,N_4490);
or U6521 (N_6521,N_4916,N_4613);
nand U6522 (N_6522,N_1939,N_632);
nand U6523 (N_6523,N_3649,N_4446);
nand U6524 (N_6524,N_1966,N_2481);
or U6525 (N_6525,N_2785,N_2711);
nor U6526 (N_6526,N_244,N_1033);
and U6527 (N_6527,N_567,N_1947);
and U6528 (N_6528,N_216,N_1975);
nand U6529 (N_6529,N_1601,N_2989);
and U6530 (N_6530,N_1431,N_1453);
and U6531 (N_6531,N_943,N_2715);
nor U6532 (N_6532,N_2647,N_2468);
nand U6533 (N_6533,N_452,N_1248);
nor U6534 (N_6534,N_1024,N_1532);
nand U6535 (N_6535,N_914,N_3177);
and U6536 (N_6536,N_2272,N_3906);
and U6537 (N_6537,N_137,N_4430);
nand U6538 (N_6538,N_290,N_3919);
nand U6539 (N_6539,N_75,N_649);
nor U6540 (N_6540,N_3674,N_1935);
or U6541 (N_6541,N_3911,N_3958);
or U6542 (N_6542,N_4686,N_2375);
or U6543 (N_6543,N_2374,N_4529);
or U6544 (N_6544,N_1356,N_3477);
or U6545 (N_6545,N_19,N_1891);
and U6546 (N_6546,N_839,N_3937);
nand U6547 (N_6547,N_1814,N_2567);
or U6548 (N_6548,N_1974,N_3855);
and U6549 (N_6549,N_4705,N_2973);
nand U6550 (N_6550,N_2278,N_180);
or U6551 (N_6551,N_3974,N_2690);
and U6552 (N_6552,N_4054,N_2177);
nand U6553 (N_6553,N_4035,N_4792);
nor U6554 (N_6554,N_3353,N_2179);
nor U6555 (N_6555,N_3850,N_3160);
nor U6556 (N_6556,N_873,N_2777);
and U6557 (N_6557,N_4147,N_2722);
or U6558 (N_6558,N_3201,N_533);
nand U6559 (N_6559,N_3773,N_4137);
and U6560 (N_6560,N_716,N_1320);
and U6561 (N_6561,N_3470,N_45);
nand U6562 (N_6562,N_2746,N_2800);
nand U6563 (N_6563,N_2486,N_1762);
and U6564 (N_6564,N_878,N_3876);
or U6565 (N_6565,N_3668,N_3380);
or U6566 (N_6566,N_3,N_1624);
and U6567 (N_6567,N_4984,N_322);
and U6568 (N_6568,N_2348,N_1993);
nand U6569 (N_6569,N_2623,N_210);
or U6570 (N_6570,N_4068,N_2267);
and U6571 (N_6571,N_4500,N_147);
nor U6572 (N_6572,N_3259,N_3614);
and U6573 (N_6573,N_4432,N_1550);
or U6574 (N_6574,N_2657,N_3705);
nor U6575 (N_6575,N_1718,N_2166);
nor U6576 (N_6576,N_196,N_3020);
nand U6577 (N_6577,N_2609,N_3703);
nand U6578 (N_6578,N_1124,N_2544);
nor U6579 (N_6579,N_353,N_1118);
nand U6580 (N_6580,N_3392,N_750);
nor U6581 (N_6581,N_4130,N_1287);
or U6582 (N_6582,N_3583,N_2929);
nand U6583 (N_6583,N_3653,N_2306);
or U6584 (N_6584,N_3519,N_4175);
nand U6585 (N_6585,N_2648,N_1871);
nor U6586 (N_6586,N_1432,N_2011);
nand U6587 (N_6587,N_1725,N_3272);
and U6588 (N_6588,N_4029,N_1824);
and U6589 (N_6589,N_3011,N_1316);
or U6590 (N_6590,N_4362,N_3985);
and U6591 (N_6591,N_421,N_4605);
or U6592 (N_6592,N_608,N_1514);
nor U6593 (N_6593,N_1442,N_1238);
or U6594 (N_6594,N_571,N_43);
nor U6595 (N_6595,N_2713,N_1537);
nand U6596 (N_6596,N_1972,N_1711);
nor U6597 (N_6597,N_1792,N_4314);
nor U6598 (N_6598,N_666,N_2425);
or U6599 (N_6599,N_4170,N_544);
and U6600 (N_6600,N_4532,N_1703);
or U6601 (N_6601,N_1697,N_2977);
and U6602 (N_6602,N_436,N_1265);
nor U6603 (N_6603,N_2949,N_2845);
or U6604 (N_6604,N_896,N_2844);
and U6605 (N_6605,N_2840,N_4318);
nand U6606 (N_6606,N_3658,N_1757);
nand U6607 (N_6607,N_4019,N_1008);
and U6608 (N_6608,N_1174,N_4142);
and U6609 (N_6609,N_3764,N_1106);
and U6610 (N_6610,N_2402,N_3069);
nor U6611 (N_6611,N_3908,N_747);
xor U6612 (N_6612,N_3795,N_2682);
or U6613 (N_6613,N_756,N_1012);
and U6614 (N_6614,N_3819,N_1831);
or U6615 (N_6615,N_4127,N_3562);
nand U6616 (N_6616,N_3887,N_2107);
and U6617 (N_6617,N_626,N_622);
nand U6618 (N_6618,N_3037,N_711);
nand U6619 (N_6619,N_4537,N_3130);
or U6620 (N_6620,N_884,N_1417);
nor U6621 (N_6621,N_4551,N_3667);
nand U6622 (N_6622,N_4053,N_656);
or U6623 (N_6623,N_3244,N_623);
or U6624 (N_6624,N_4985,N_4515);
and U6625 (N_6625,N_783,N_1821);
and U6626 (N_6626,N_3612,N_2575);
nor U6627 (N_6627,N_4367,N_3372);
nor U6628 (N_6628,N_4759,N_2345);
or U6629 (N_6629,N_2284,N_1713);
nand U6630 (N_6630,N_4640,N_3490);
or U6631 (N_6631,N_3927,N_1098);
and U6632 (N_6632,N_1989,N_3406);
or U6633 (N_6633,N_760,N_369);
nand U6634 (N_6634,N_3527,N_4082);
nand U6635 (N_6635,N_1784,N_2821);
nand U6636 (N_6636,N_4710,N_967);
nor U6637 (N_6637,N_616,N_1051);
or U6638 (N_6638,N_2514,N_3511);
and U6639 (N_6639,N_1209,N_1380);
and U6640 (N_6640,N_1413,N_2513);
or U6641 (N_6641,N_4453,N_442);
or U6642 (N_6642,N_4949,N_801);
and U6643 (N_6643,N_1776,N_3432);
or U6644 (N_6644,N_987,N_1167);
nand U6645 (N_6645,N_4472,N_3859);
nor U6646 (N_6646,N_702,N_4057);
nand U6647 (N_6647,N_266,N_2237);
nand U6648 (N_6648,N_4378,N_3676);
nand U6649 (N_6649,N_2793,N_1170);
or U6650 (N_6650,N_1471,N_743);
or U6651 (N_6651,N_4355,N_3986);
nand U6652 (N_6652,N_883,N_1451);
and U6653 (N_6653,N_2154,N_3164);
nand U6654 (N_6654,N_2007,N_3895);
and U6655 (N_6655,N_1598,N_2578);
xnor U6656 (N_6656,N_4707,N_633);
and U6657 (N_6657,N_4187,N_195);
nor U6658 (N_6658,N_3607,N_3526);
nor U6659 (N_6659,N_1140,N_2944);
and U6660 (N_6660,N_1833,N_2805);
nor U6661 (N_6661,N_4882,N_2359);
xor U6662 (N_6662,N_4910,N_2594);
and U6663 (N_6663,N_3512,N_4617);
nand U6664 (N_6664,N_3672,N_2344);
or U6665 (N_6665,N_1899,N_2704);
nand U6666 (N_6666,N_4215,N_1114);
and U6667 (N_6667,N_4818,N_1187);
and U6668 (N_6668,N_4546,N_2642);
nor U6669 (N_6669,N_3991,N_21);
or U6670 (N_6670,N_4206,N_1497);
and U6671 (N_6671,N_3050,N_3984);
and U6672 (N_6672,N_2035,N_4165);
nor U6673 (N_6673,N_1068,N_4977);
nor U6674 (N_6674,N_916,N_3613);
and U6675 (N_6675,N_3831,N_460);
nand U6676 (N_6676,N_3086,N_3656);
and U6677 (N_6677,N_1756,N_1256);
nor U6678 (N_6678,N_551,N_1157);
or U6679 (N_6679,N_3172,N_4735);
and U6680 (N_6680,N_1837,N_1149);
nand U6681 (N_6681,N_89,N_582);
or U6682 (N_6682,N_3487,N_1375);
and U6683 (N_6683,N_4392,N_1929);
and U6684 (N_6684,N_261,N_3274);
and U6685 (N_6685,N_44,N_3478);
nor U6686 (N_6686,N_4976,N_890);
and U6687 (N_6687,N_383,N_4052);
nand U6688 (N_6688,N_481,N_465);
or U6689 (N_6689,N_4474,N_1693);
nor U6690 (N_6690,N_3435,N_4604);
nand U6691 (N_6691,N_3978,N_951);
nor U6692 (N_6692,N_850,N_311);
or U6693 (N_6693,N_2817,N_1383);
nand U6694 (N_6694,N_1175,N_4838);
nand U6695 (N_6695,N_3222,N_4794);
nand U6696 (N_6696,N_2370,N_2912);
and U6697 (N_6697,N_2883,N_1148);
nor U6698 (N_6698,N_2339,N_4495);
nor U6699 (N_6699,N_1305,N_885);
and U6700 (N_6700,N_1020,N_2925);
nand U6701 (N_6701,N_1656,N_4101);
or U6702 (N_6702,N_4737,N_4943);
nor U6703 (N_6703,N_1147,N_3206);
or U6704 (N_6704,N_3755,N_4642);
or U6705 (N_6705,N_955,N_1976);
nand U6706 (N_6706,N_171,N_1960);
or U6707 (N_6707,N_1489,N_2061);
or U6708 (N_6708,N_2101,N_3678);
or U6709 (N_6709,N_969,N_176);
or U6710 (N_6710,N_1786,N_2519);
nand U6711 (N_6711,N_911,N_1065);
nand U6712 (N_6712,N_2764,N_2174);
or U6713 (N_6713,N_2401,N_1671);
and U6714 (N_6714,N_2155,N_4178);
or U6715 (N_6715,N_3903,N_2978);
nor U6716 (N_6716,N_1925,N_4273);
and U6717 (N_6717,N_1459,N_2752);
nor U6718 (N_6718,N_2110,N_2250);
nand U6719 (N_6719,N_135,N_376);
nand U6720 (N_6720,N_4203,N_4725);
nor U6721 (N_6721,N_2917,N_2013);
nor U6722 (N_6722,N_3753,N_1613);
nor U6723 (N_6723,N_4662,N_3989);
or U6724 (N_6724,N_836,N_13);
and U6725 (N_6725,N_3835,N_1121);
and U6726 (N_6726,N_591,N_3186);
or U6727 (N_6727,N_1590,N_1343);
or U6728 (N_6728,N_2813,N_2066);
nand U6729 (N_6729,N_1865,N_3752);
or U6730 (N_6730,N_3089,N_3518);
nand U6731 (N_6731,N_4513,N_1276);
and U6732 (N_6732,N_570,N_1139);
nand U6733 (N_6733,N_3659,N_927);
nor U6734 (N_6734,N_25,N_288);
or U6735 (N_6735,N_1054,N_1362);
nor U6736 (N_6736,N_4740,N_318);
nand U6737 (N_6737,N_4972,N_56);
and U6738 (N_6738,N_2863,N_3943);
nand U6739 (N_6739,N_4814,N_268);
or U6740 (N_6740,N_3383,N_1759);
nor U6741 (N_6741,N_3026,N_3502);
nand U6742 (N_6742,N_1490,N_4105);
and U6743 (N_6743,N_3356,N_963);
nand U6744 (N_6744,N_2558,N_3968);
nor U6745 (N_6745,N_4758,N_2429);
nor U6746 (N_6746,N_1401,N_4169);
nor U6747 (N_6747,N_1914,N_58);
or U6748 (N_6748,N_1179,N_851);
and U6749 (N_6749,N_3816,N_536);
and U6750 (N_6750,N_4266,N_1665);
and U6751 (N_6751,N_1331,N_4751);
nor U6752 (N_6752,N_4448,N_275);
and U6753 (N_6753,N_3275,N_516);
or U6754 (N_6754,N_464,N_572);
and U6755 (N_6755,N_4148,N_1038);
and U6756 (N_6756,N_200,N_1653);
and U6757 (N_6757,N_3956,N_124);
nor U6758 (N_6758,N_2000,N_1221);
and U6759 (N_6759,N_1607,N_4548);
or U6760 (N_6760,N_2966,N_2466);
nand U6761 (N_6761,N_4126,N_1664);
or U6762 (N_6762,N_2539,N_2027);
and U6763 (N_6763,N_3420,N_441);
nand U6764 (N_6764,N_3216,N_1755);
nand U6765 (N_6765,N_4522,N_4258);
nand U6766 (N_6766,N_4452,N_1402);
nor U6767 (N_6767,N_3192,N_4927);
and U6768 (N_6768,N_3041,N_4044);
nor U6769 (N_6769,N_90,N_4545);
and U6770 (N_6770,N_4661,N_24);
or U6771 (N_6771,N_858,N_1339);
nor U6772 (N_6772,N_599,N_4467);
and U6773 (N_6773,N_53,N_4607);
nor U6774 (N_6774,N_1079,N_2736);
or U6775 (N_6775,N_4783,N_1097);
or U6776 (N_6776,N_4030,N_3433);
nor U6777 (N_6777,N_2981,N_3923);
or U6778 (N_6778,N_3776,N_3125);
nand U6779 (N_6779,N_4189,N_3339);
nand U6780 (N_6780,N_316,N_4793);
or U6781 (N_6781,N_1286,N_80);
or U6782 (N_6782,N_852,N_4132);
or U6783 (N_6783,N_3665,N_1232);
nand U6784 (N_6784,N_3576,N_798);
and U6785 (N_6785,N_1818,N_1669);
and U6786 (N_6786,N_1595,N_2645);
nor U6787 (N_6787,N_4504,N_2508);
nor U6788 (N_6788,N_213,N_4494);
nand U6789 (N_6789,N_989,N_2658);
or U6790 (N_6790,N_2204,N_2003);
and U6791 (N_6791,N_2661,N_3338);
nor U6792 (N_6792,N_2887,N_2058);
nor U6793 (N_6793,N_1949,N_1556);
nor U6794 (N_6794,N_2541,N_690);
xor U6795 (N_6795,N_2410,N_2417);
or U6796 (N_6796,N_444,N_4526);
and U6797 (N_6797,N_812,N_299);
nand U6798 (N_6798,N_1206,N_1856);
nor U6799 (N_6799,N_1161,N_1195);
nor U6800 (N_6800,N_4592,N_158);
nand U6801 (N_6801,N_1210,N_2451);
nor U6802 (N_6802,N_3556,N_395);
nand U6803 (N_6803,N_3407,N_1310);
nand U6804 (N_6804,N_4421,N_3121);
and U6805 (N_6805,N_2600,N_2346);
nor U6806 (N_6806,N_4655,N_4319);
nand U6807 (N_6807,N_1066,N_1458);
and U6808 (N_6808,N_4352,N_1197);
nand U6809 (N_6809,N_131,N_1395);
nor U6810 (N_6810,N_3535,N_1226);
and U6811 (N_6811,N_3017,N_4679);
and U6812 (N_6812,N_2281,N_4066);
or U6813 (N_6813,N_3814,N_484);
nand U6814 (N_6814,N_4390,N_753);
and U6815 (N_6815,N_4261,N_2049);
nor U6816 (N_6816,N_4991,N_501);
and U6817 (N_6817,N_3475,N_1643);
or U6818 (N_6818,N_1542,N_4745);
nor U6819 (N_6819,N_1968,N_4955);
and U6820 (N_6820,N_4129,N_2720);
and U6821 (N_6821,N_2536,N_106);
nand U6822 (N_6822,N_3836,N_749);
and U6823 (N_6823,N_3938,N_732);
or U6824 (N_6824,N_2548,N_3799);
nand U6825 (N_6825,N_1618,N_2310);
nand U6826 (N_6826,N_2854,N_1223);
and U6827 (N_6827,N_1806,N_4709);
and U6828 (N_6828,N_1428,N_414);
nor U6829 (N_6829,N_2996,N_1285);
nor U6830 (N_6830,N_1057,N_4967);
or U6831 (N_6831,N_1419,N_723);
nand U6832 (N_6832,N_1600,N_4023);
and U6833 (N_6833,N_3038,N_1052);
and U6834 (N_6834,N_3746,N_2478);
nand U6835 (N_6835,N_3736,N_4584);
or U6836 (N_6836,N_3393,N_2706);
and U6837 (N_6837,N_103,N_161);
nand U6838 (N_6838,N_1536,N_1635);
and U6839 (N_6839,N_4587,N_2207);
nor U6840 (N_6840,N_3597,N_343);
nor U6841 (N_6841,N_1452,N_1927);
and U6842 (N_6842,N_1846,N_1793);
or U6843 (N_6843,N_4092,N_3682);
and U6844 (N_6844,N_1701,N_1408);
nor U6845 (N_6845,N_3313,N_2096);
and U6846 (N_6846,N_3075,N_2450);
nor U6847 (N_6847,N_140,N_3324);
nand U6848 (N_6848,N_128,N_1443);
nand U6849 (N_6849,N_889,N_2791);
nand U6850 (N_6850,N_3459,N_2705);
or U6851 (N_6851,N_2960,N_726);
nor U6852 (N_6852,N_378,N_4762);
or U6853 (N_6853,N_1924,N_4508);
or U6854 (N_6854,N_1565,N_4403);
nor U6855 (N_6855,N_1160,N_3898);
nor U6856 (N_6856,N_926,N_2714);
or U6857 (N_6857,N_2986,N_4899);
or U6858 (N_6858,N_3524,N_4952);
nand U6859 (N_6859,N_74,N_87);
or U6860 (N_6860,N_1752,N_3220);
nor U6861 (N_6861,N_3022,N_1672);
nand U6862 (N_6862,N_1964,N_3479);
nor U6863 (N_6863,N_2806,N_4785);
and U6864 (N_6864,N_4997,N_1544);
or U6865 (N_6865,N_1325,N_1923);
nand U6866 (N_6866,N_1018,N_4752);
nor U6867 (N_6867,N_2743,N_1123);
and U6868 (N_6868,N_2964,N_3303);
nand U6869 (N_6869,N_508,N_2091);
nand U6870 (N_6870,N_528,N_3700);
or U6871 (N_6871,N_264,N_4782);
nand U6872 (N_6872,N_2271,N_308);
and U6873 (N_6873,N_136,N_2681);
and U6874 (N_6874,N_3930,N_1365);
or U6875 (N_6875,N_2483,N_1582);
nand U6876 (N_6876,N_4202,N_3882);
and U6877 (N_6877,N_4547,N_4125);
nand U6878 (N_6878,N_1075,N_2238);
nor U6879 (N_6879,N_1802,N_1798);
and U6880 (N_6880,N_2063,N_2494);
and U6881 (N_6881,N_3158,N_1603);
xnor U6882 (N_6882,N_4081,N_2956);
or U6883 (N_6883,N_729,N_4230);
nor U6884 (N_6884,N_3031,N_1712);
or U6885 (N_6885,N_1930,N_3264);
and U6886 (N_6886,N_2198,N_4020);
and U6887 (N_6887,N_4174,N_3704);
nor U6888 (N_6888,N_1963,N_782);
and U6889 (N_6889,N_3635,N_3707);
or U6890 (N_6890,N_4371,N_1162);
or U6891 (N_6891,N_4157,N_2801);
or U6892 (N_6892,N_3623,N_485);
and U6893 (N_6893,N_146,N_3093);
or U6894 (N_6894,N_1491,N_4849);
and U6895 (N_6895,N_4459,N_4961);
nand U6896 (N_6896,N_4810,N_4887);
or U6897 (N_6897,N_2422,N_3494);
nand U6898 (N_6898,N_2641,N_1086);
and U6899 (N_6899,N_1965,N_223);
and U6900 (N_6900,N_1137,N_4076);
or U6901 (N_6901,N_645,N_3427);
or U6902 (N_6902,N_2550,N_2524);
and U6903 (N_6903,N_4483,N_2141);
nand U6904 (N_6904,N_4858,N_3809);
nor U6905 (N_6905,N_3997,N_3950);
or U6906 (N_6906,N_2540,N_3804);
or U6907 (N_6907,N_2848,N_4251);
and U6908 (N_6908,N_4333,N_117);
or U6909 (N_6909,N_4255,N_606);
nand U6910 (N_6910,N_3345,N_2861);
or U6911 (N_6911,N_562,N_906);
or U6912 (N_6912,N_3709,N_4381);
nand U6913 (N_6913,N_3807,N_904);
nand U6914 (N_6914,N_3328,N_894);
nor U6915 (N_6915,N_4773,N_559);
and U6916 (N_6916,N_4507,N_1996);
nor U6917 (N_6917,N_846,N_4652);
nand U6918 (N_6918,N_4718,N_2232);
and U6919 (N_6919,N_3176,N_1547);
or U6920 (N_6920,N_4738,N_1100);
and U6921 (N_6921,N_2604,N_4732);
or U6922 (N_6922,N_3905,N_4796);
xnor U6923 (N_6923,N_314,N_447);
or U6924 (N_6924,N_4874,N_4973);
and U6925 (N_6925,N_3894,N_2721);
nor U6926 (N_6926,N_4419,N_456);
nor U6927 (N_6927,N_1449,N_2465);
or U6928 (N_6928,N_4756,N_3594);
and U6929 (N_6929,N_4482,N_2084);
nand U6930 (N_6930,N_513,N_4042);
and U6931 (N_6931,N_2952,N_2825);
and U6932 (N_6932,N_2475,N_1980);
and U6933 (N_6933,N_4918,N_112);
and U6934 (N_6934,N_2676,N_703);
and U6935 (N_6935,N_2992,N_3256);
nor U6936 (N_6936,N_3830,N_704);
nor U6937 (N_6937,N_2837,N_2186);
nor U6938 (N_6938,N_2768,N_4182);
nor U6939 (N_6939,N_3099,N_2810);
xnor U6940 (N_6940,N_1498,N_3951);
and U6941 (N_6941,N_3132,N_2625);
and U6942 (N_6942,N_222,N_918);
or U6943 (N_6943,N_4099,N_2298);
or U6944 (N_6944,N_3992,N_4597);
nor U6945 (N_6945,N_769,N_2572);
and U6946 (N_6946,N_2433,N_4034);
nor U6947 (N_6947,N_2203,N_2456);
nor U6948 (N_6948,N_2394,N_1662);
or U6949 (N_6949,N_4240,N_3655);
nand U6950 (N_6950,N_3839,N_2235);
or U6951 (N_6951,N_4689,N_4445);
nand U6952 (N_6952,N_17,N_139);
or U6953 (N_6953,N_482,N_4359);
nand U6954 (N_6954,N_2309,N_1273);
nand U6955 (N_6955,N_4561,N_2131);
nor U6956 (N_6956,N_548,N_2173);
nand U6957 (N_6957,N_1961,N_1647);
and U6958 (N_6958,N_1122,N_2249);
or U6959 (N_6959,N_2304,N_339);
nand U6960 (N_6960,N_3720,N_426);
nand U6961 (N_6961,N_3161,N_531);
nand U6962 (N_6962,N_1422,N_2990);
xor U6963 (N_6963,N_4763,N_2212);
and U6964 (N_6964,N_3100,N_1528);
and U6965 (N_6965,N_2570,N_2787);
or U6966 (N_6966,N_3149,N_4674);
nor U6967 (N_6967,N_189,N_2480);
or U6968 (N_6968,N_4798,N_3691);
nor U6969 (N_6969,N_868,N_745);
nand U6970 (N_6970,N_2701,N_384);
nand U6971 (N_6971,N_3663,N_2685);
and U6972 (N_6972,N_3805,N_2627);
or U6973 (N_6973,N_4820,N_3854);
and U6974 (N_6974,N_277,N_3265);
nor U6975 (N_6975,N_2692,N_3325);
and U6976 (N_6976,N_2242,N_4627);
nor U6977 (N_6977,N_4856,N_1403);
or U6978 (N_6978,N_1324,N_1294);
nand U6979 (N_6979,N_947,N_880);
nor U6980 (N_6980,N_2241,N_3880);
nand U6981 (N_6981,N_165,N_3413);
and U6982 (N_6982,N_4945,N_2196);
nor U6983 (N_6983,N_2280,N_1645);
and U6984 (N_6984,N_2799,N_1769);
and U6985 (N_6985,N_2276,N_980);
nor U6986 (N_6986,N_3593,N_1094);
and U6987 (N_6987,N_830,N_4610);
nand U6988 (N_6988,N_374,N_795);
or U6989 (N_6989,N_3112,N_379);
nand U6990 (N_6990,N_229,N_2458);
and U6991 (N_6991,N_2954,N_3568);
nand U6992 (N_6992,N_6,N_221);
nand U6993 (N_6993,N_4668,N_4589);
or U6994 (N_6994,N_1444,N_1579);
nor U6995 (N_6995,N_3862,N_3760);
nand U6996 (N_6996,N_2533,N_183);
nor U6997 (N_6997,N_3098,N_634);
nand U6998 (N_6998,N_2988,N_3821);
nand U6999 (N_6999,N_3581,N_2094);
nand U7000 (N_7000,N_1766,N_2560);
and U7001 (N_7001,N_3247,N_3290);
nor U7002 (N_7002,N_776,N_2391);
nor U7003 (N_7003,N_4393,N_691);
nor U7004 (N_7004,N_2982,N_713);
or U7005 (N_7005,N_2913,N_304);
nor U7006 (N_7006,N_2808,N_4484);
or U7007 (N_7007,N_4656,N_2025);
nand U7008 (N_7008,N_4340,N_145);
nand U7009 (N_7009,N_2574,N_3311);
nand U7010 (N_7010,N_3471,N_1751);
nor U7011 (N_7011,N_3019,N_4803);
and U7012 (N_7012,N_2618,N_2843);
or U7013 (N_7013,N_902,N_1811);
or U7014 (N_7014,N_984,N_3074);
and U7015 (N_7015,N_2684,N_3295);
and U7016 (N_7016,N_4466,N_2470);
nor U7017 (N_7017,N_773,N_855);
or U7018 (N_7018,N_3049,N_457);
and U7019 (N_7019,N_2683,N_4270);
nand U7020 (N_7020,N_1807,N_3091);
nor U7021 (N_7021,N_3579,N_2020);
or U7022 (N_7022,N_1440,N_172);
and U7023 (N_7023,N_3246,N_4675);
and U7024 (N_7024,N_3742,N_4842);
nand U7025 (N_7025,N_477,N_905);
nand U7026 (N_7026,N_26,N_4436);
and U7027 (N_7027,N_2874,N_3640);
and U7028 (N_7028,N_2342,N_3609);
nor U7029 (N_7029,N_4600,N_2449);
and U7030 (N_7030,N_4423,N_3260);
or U7031 (N_7031,N_2445,N_4747);
nor U7032 (N_7032,N_3939,N_3994);
and U7033 (N_7033,N_3843,N_1646);
nor U7034 (N_7034,N_2635,N_3942);
nand U7035 (N_7035,N_4687,N_4209);
or U7036 (N_7036,N_3884,N_4896);
nor U7037 (N_7037,N_3498,N_4120);
nor U7038 (N_7038,N_495,N_133);
nand U7039 (N_7039,N_101,N_688);
or U7040 (N_7040,N_1668,N_4233);
or U7041 (N_7041,N_1893,N_3973);
nor U7042 (N_7042,N_2748,N_4841);
nand U7043 (N_7043,N_2933,N_3486);
or U7044 (N_7044,N_4278,N_1484);
nand U7045 (N_7045,N_4570,N_3870);
xor U7046 (N_7046,N_1896,N_3021);
nand U7047 (N_7047,N_1518,N_4160);
nor U7048 (N_7048,N_2171,N_1742);
or U7049 (N_7049,N_3684,N_4909);
and U7050 (N_7050,N_3231,N_1344);
nor U7051 (N_7051,N_2150,N_627);
nand U7052 (N_7052,N_4902,N_102);
and U7053 (N_7053,N_1946,N_258);
nand U7054 (N_7054,N_1609,N_4272);
nor U7055 (N_7055,N_472,N_3289);
nor U7056 (N_7056,N_2707,N_735);
or U7057 (N_7057,N_1774,N_1496);
or U7058 (N_7058,N_4024,N_4097);
nor U7059 (N_7059,N_1244,N_1236);
or U7060 (N_7060,N_2327,N_1841);
or U7061 (N_7061,N_3873,N_1377);
and U7062 (N_7062,N_1685,N_2217);
and U7063 (N_7063,N_576,N_4966);
and U7064 (N_7064,N_3138,N_2892);
nand U7065 (N_7065,N_923,N_3758);
nor U7066 (N_7066,N_2324,N_2411);
or U7067 (N_7067,N_49,N_3381);
and U7068 (N_7068,N_3513,N_950);
nor U7069 (N_7069,N_658,N_4799);
nand U7070 (N_7070,N_1418,N_3717);
nand U7071 (N_7071,N_2901,N_1003);
and U7072 (N_7072,N_1867,N_3087);
and U7073 (N_7073,N_88,N_2502);
or U7074 (N_7074,N_4324,N_224);
nor U7075 (N_7075,N_129,N_1545);
or U7076 (N_7076,N_86,N_4387);
and U7077 (N_7077,N_1369,N_1389);
nand U7078 (N_7078,N_3450,N_2871);
or U7079 (N_7079,N_365,N_11);
nor U7080 (N_7080,N_4260,N_2898);
nor U7081 (N_7081,N_2074,N_2282);
or U7082 (N_7082,N_802,N_1688);
nand U7083 (N_7083,N_3414,N_211);
and U7084 (N_7084,N_1781,N_3389);
nor U7085 (N_7085,N_334,N_3285);
and U7086 (N_7086,N_3605,N_3062);
nand U7087 (N_7087,N_3423,N_2321);
and U7088 (N_7088,N_3412,N_2211);
or U7089 (N_7089,N_4422,N_326);
nand U7090 (N_7090,N_3054,N_826);
nor U7091 (N_7091,N_3713,N_3111);
nor U7092 (N_7092,N_4633,N_2788);
nor U7093 (N_7093,N_2206,N_3608);
nor U7094 (N_7094,N_3554,N_130);
or U7095 (N_7095,N_358,N_2313);
nand U7096 (N_7096,N_3033,N_1950);
nor U7097 (N_7097,N_648,N_341);
and U7098 (N_7098,N_152,N_3444);
and U7099 (N_7099,N_4330,N_1836);
or U7100 (N_7100,N_4611,N_2927);
and U7101 (N_7101,N_4199,N_427);
nor U7102 (N_7102,N_638,N_1830);
nor U7103 (N_7103,N_1171,N_1495);
and U7104 (N_7104,N_3792,N_2361);
nor U7105 (N_7105,N_2236,N_2336);
nor U7106 (N_7106,N_1388,N_4335);
nand U7107 (N_7107,N_4036,N_660);
and U7108 (N_7108,N_4418,N_3005);
and U7109 (N_7109,N_1572,N_2576);
nor U7110 (N_7110,N_2437,N_696);
and U7111 (N_7111,N_3920,N_2197);
or U7112 (N_7112,N_3829,N_1892);
and U7113 (N_7113,N_2245,N_961);
or U7114 (N_7114,N_2369,N_2233);
and U7115 (N_7115,N_4366,N_3798);
nor U7116 (N_7116,N_2225,N_2125);
and U7117 (N_7117,N_177,N_4566);
or U7118 (N_7118,N_39,N_2501);
nor U7119 (N_7119,N_2067,N_2062);
and U7120 (N_7120,N_511,N_1721);
or U7121 (N_7121,N_2671,N_95);
nand U7122 (N_7122,N_412,N_860);
nand U7123 (N_7123,N_23,N_4727);
or U7124 (N_7124,N_2565,N_1144);
or U7125 (N_7125,N_1332,N_3232);
nand U7126 (N_7126,N_655,N_1415);
and U7127 (N_7127,N_4797,N_1729);
nand U7128 (N_7128,N_2046,N_1777);
nand U7129 (N_7129,N_375,N_3113);
or U7130 (N_7130,N_1089,N_2223);
nor U7131 (N_7131,N_547,N_1780);
and U7132 (N_7132,N_4930,N_3666);
or U7133 (N_7133,N_3374,N_4437);
nand U7134 (N_7134,N_741,N_4969);
nand U7135 (N_7135,N_2834,N_204);
nor U7136 (N_7136,N_3712,N_4749);
nand U7137 (N_7137,N_3926,N_639);
or U7138 (N_7138,N_2538,N_1694);
nand U7139 (N_7139,N_1398,N_4405);
nand U7140 (N_7140,N_653,N_4286);
nand U7141 (N_7141,N_1423,N_3245);
or U7142 (N_7142,N_1835,N_791);
nand U7143 (N_7143,N_2138,N_1916);
nor U7144 (N_7144,N_4812,N_3097);
nor U7145 (N_7145,N_3321,N_2979);
nand U7146 (N_7146,N_3549,N_2051);
nor U7147 (N_7147,N_107,N_725);
nor U7148 (N_7148,N_4596,N_3602);
or U7149 (N_7149,N_2592,N_3061);
or U7150 (N_7150,N_4212,N_3563);
nor U7151 (N_7151,N_2638,N_3106);
or U7152 (N_7152,N_710,N_3532);
nand U7153 (N_7153,N_3457,N_3036);
nand U7154 (N_7154,N_2077,N_4071);
and U7155 (N_7155,N_2322,N_3032);
nor U7156 (N_7156,N_1474,N_1262);
or U7157 (N_7157,N_156,N_2114);
nor U7158 (N_7158,N_4639,N_3546);
or U7159 (N_7159,N_1790,N_3732);
nand U7160 (N_7160,N_1354,N_1791);
nor U7161 (N_7161,N_2646,N_3948);
nand U7162 (N_7162,N_2014,N_2870);
nand U7163 (N_7163,N_3652,N_897);
xor U7164 (N_7164,N_2762,N_2668);
nor U7165 (N_7165,N_3878,N_1915);
or U7166 (N_7166,N_274,N_2865);
nand U7167 (N_7167,N_3377,N_640);
nand U7168 (N_7168,N_4115,N_4823);
and U7169 (N_7169,N_631,N_1205);
nand U7170 (N_7170,N_4321,N_1237);
nor U7171 (N_7171,N_2416,N_1293);
nand U7172 (N_7172,N_4179,N_2812);
nor U7173 (N_7173,N_2608,N_4211);
nand U7174 (N_7174,N_2491,N_4667);
or U7175 (N_7175,N_4026,N_988);
nor U7176 (N_7176,N_1758,N_604);
or U7177 (N_7177,N_1512,N_3060);
nor U7178 (N_7178,N_2797,N_1723);
nor U7179 (N_7179,N_94,N_818);
nor U7180 (N_7180,N_3791,N_4564);
and U7181 (N_7181,N_617,N_2108);
or U7182 (N_7182,N_232,N_437);
nor U7183 (N_7183,N_2367,N_2390);
nand U7184 (N_7184,N_1659,N_2499);
xnor U7185 (N_7185,N_4205,N_856);
nand U7186 (N_7186,N_3434,N_2357);
or U7187 (N_7187,N_3718,N_588);
nor U7188 (N_7188,N_920,N_197);
nand U7189 (N_7189,N_4531,N_3092);
and U7190 (N_7190,N_3574,N_3680);
nor U7191 (N_7191,N_772,N_720);
and U7192 (N_7192,N_762,N_1194);
nand U7193 (N_7193,N_2598,N_1465);
or U7194 (N_7194,N_994,N_2897);
nor U7195 (N_7195,N_3763,N_1270);
and U7196 (N_7196,N_507,N_2571);
nor U7197 (N_7197,N_1642,N_3249);
and U7198 (N_7198,N_2255,N_2859);
nor U7199 (N_7199,N_2790,N_2351);
nand U7200 (N_7200,N_302,N_2078);
nor U7201 (N_7201,N_2769,N_4186);
nor U7202 (N_7202,N_1633,N_3150);
or U7203 (N_7203,N_198,N_2773);
nand U7204 (N_7204,N_1334,N_1060);
and U7205 (N_7205,N_986,N_1372);
nand U7206 (N_7206,N_2260,N_1922);
nor U7207 (N_7207,N_3114,N_4691);
and U7208 (N_7208,N_3521,N_4760);
or U7209 (N_7209,N_1940,N_1737);
and U7210 (N_7210,N_4606,N_4534);
nand U7211 (N_7211,N_3833,N_4644);
or U7212 (N_7212,N_3869,N_4865);
nor U7213 (N_7213,N_891,N_875);
and U7214 (N_7214,N_4938,N_2620);
or U7215 (N_7215,N_1103,N_865);
or U7216 (N_7216,N_644,N_4334);
nand U7217 (N_7217,N_563,N_2496);
and U7218 (N_7218,N_3108,N_3834);
nor U7219 (N_7219,N_1705,N_373);
nand U7220 (N_7220,N_1247,N_2776);
nor U7221 (N_7221,N_1839,N_728);
nand U7222 (N_7222,N_2012,N_2957);
nor U7223 (N_7223,N_3803,N_3004);
nor U7224 (N_7224,N_3236,N_105);
or U7225 (N_7225,N_4768,N_3382);
nand U7226 (N_7226,N_303,N_3237);
and U7227 (N_7227,N_4222,N_4786);
nor U7228 (N_7228,N_4641,N_4941);
nand U7229 (N_7229,N_1259,N_3202);
xnor U7230 (N_7230,N_4021,N_4559);
nor U7231 (N_7231,N_683,N_3537);
nand U7232 (N_7232,N_672,N_2522);
xnor U7233 (N_7233,N_1563,N_1614);
or U7234 (N_7234,N_2354,N_1515);
nand U7235 (N_7235,N_390,N_3841);
xor U7236 (N_7236,N_4839,N_1049);
nand U7237 (N_7237,N_1728,N_522);
or U7238 (N_7238,N_4461,N_2050);
nand U7239 (N_7239,N_2065,N_4871);
nor U7240 (N_7240,N_1561,N_2368);
and U7241 (N_7241,N_1313,N_2889);
and U7242 (N_7242,N_2888,N_2505);
and U7243 (N_7243,N_30,N_2660);
and U7244 (N_7244,N_2129,N_1359);
nor U7245 (N_7245,N_1013,N_4417);
or U7246 (N_7246,N_3159,N_1438);
nand U7247 (N_7247,N_3133,N_2798);
or U7248 (N_7248,N_4425,N_907);
nand U7249 (N_7249,N_3636,N_2111);
or U7250 (N_7250,N_443,N_319);
or U7251 (N_7251,N_3981,N_771);
nand U7252 (N_7252,N_4207,N_561);
and U7253 (N_7253,N_4025,N_2899);
and U7254 (N_7254,N_983,N_882);
nand U7255 (N_7255,N_1335,N_2252);
or U7256 (N_7256,N_4413,N_1549);
nor U7257 (N_7257,N_4688,N_3332);
nor U7258 (N_7258,N_1696,N_4809);
nor U7259 (N_7259,N_1558,N_4372);
nand U7260 (N_7260,N_100,N_1917);
and U7261 (N_7261,N_166,N_3544);
or U7262 (N_7262,N_1678,N_4965);
and U7263 (N_7263,N_3219,N_4929);
and U7264 (N_7264,N_2680,N_4070);
or U7265 (N_7265,N_1158,N_3892);
nand U7266 (N_7266,N_3747,N_3271);
nand U7267 (N_7267,N_831,N_3660);
or U7268 (N_7268,N_4947,N_4632);
nand U7269 (N_7269,N_2056,N_1382);
nor U7270 (N_7270,N_1493,N_2412);
nand U7271 (N_7271,N_1307,N_4685);
nand U7272 (N_7272,N_3270,N_3027);
and U7273 (N_7273,N_1702,N_4269);
nor U7274 (N_7274,N_2498,N_1134);
and U7275 (N_7275,N_4353,N_3308);
nand U7276 (N_7276,N_4609,N_2325);
or U7277 (N_7277,N_629,N_3743);
and U7278 (N_7278,N_2112,N_2185);
and U7279 (N_7279,N_483,N_3861);
nor U7280 (N_7280,N_3849,N_685);
or U7281 (N_7281,N_1340,N_410);
nor U7282 (N_7282,N_2511,N_4435);
nand U7283 (N_7283,N_4063,N_3715);
nand U7284 (N_7284,N_2590,N_3567);
or U7285 (N_7285,N_2961,N_4427);
or U7286 (N_7286,N_3664,N_4499);
nor U7287 (N_7287,N_3001,N_429);
and U7288 (N_7288,N_179,N_1909);
or U7289 (N_7289,N_3896,N_4062);
nor U7290 (N_7290,N_3352,N_4907);
or U7291 (N_7291,N_1557,N_479);
nand U7292 (N_7292,N_3312,N_4322);
or U7293 (N_7293,N_3915,N_2266);
nand U7294 (N_7294,N_3051,N_2759);
or U7295 (N_7295,N_1014,N_1754);
nand U7296 (N_7296,N_4292,N_2160);
nand U7297 (N_7297,N_674,N_3109);
nor U7298 (N_7298,N_928,N_3645);
nor U7299 (N_7299,N_4813,N_3363);
or U7300 (N_7300,N_3140,N_4396);
or U7301 (N_7301,N_4256,N_4903);
or U7302 (N_7302,N_3960,N_4145);
and U7303 (N_7303,N_1661,N_2184);
nor U7304 (N_7304,N_3480,N_301);
and U7305 (N_7305,N_113,N_3234);
nand U7306 (N_7306,N_2240,N_4536);
nand U7307 (N_7307,N_1748,N_2406);
or U7308 (N_7308,N_1302,N_2640);
nor U7309 (N_7309,N_4382,N_1425);
nor U7310 (N_7310,N_1152,N_2672);
and U7311 (N_7311,N_2454,N_2579);
nand U7312 (N_7312,N_4241,N_3376);
or U7313 (N_7313,N_3999,N_3897);
or U7314 (N_7314,N_1164,N_1834);
nor U7315 (N_7315,N_385,N_2636);
and U7316 (N_7316,N_3865,N_1569);
nor U7317 (N_7317,N_3565,N_1274);
nor U7318 (N_7318,N_3538,N_4077);
and U7319 (N_7319,N_4560,N_2872);
or U7320 (N_7320,N_1082,N_2905);
nor U7321 (N_7321,N_3550,N_1808);
nand U7322 (N_7322,N_1073,N_837);
and U7323 (N_7323,N_2139,N_2780);
and U7324 (N_7324,N_4693,N_46);
or U7325 (N_7325,N_1203,N_1370);
nor U7326 (N_7326,N_1078,N_3806);
nand U7327 (N_7327,N_1500,N_1110);
and U7328 (N_7328,N_150,N_3225);
or U7329 (N_7329,N_70,N_1102);
nor U7330 (N_7330,N_1715,N_4775);
nand U7331 (N_7331,N_4289,N_3469);
and U7332 (N_7332,N_4721,N_3945);
nor U7333 (N_7333,N_404,N_1615);
and U7334 (N_7334,N_3191,N_1155);
or U7335 (N_7335,N_3373,N_3592);
nand U7336 (N_7336,N_3451,N_42);
nand U7337 (N_7337,N_3586,N_1675);
nor U7338 (N_7338,N_388,N_3188);
nand U7339 (N_7339,N_2737,N_4936);
or U7340 (N_7340,N_248,N_3288);
or U7341 (N_7341,N_4080,N_3802);
and U7342 (N_7342,N_246,N_2628);
and U7343 (N_7343,N_1787,N_1686);
nand U7344 (N_7344,N_1092,N_2691);
nand U7345 (N_7345,N_1522,N_265);
or U7346 (N_7346,N_845,N_1773);
and U7347 (N_7347,N_1433,N_138);
nor U7348 (N_7348,N_160,N_163);
and U7349 (N_7349,N_3641,N_3797);
nand U7350 (N_7350,N_1132,N_1782);
nor U7351 (N_7351,N_4807,N_806);
nor U7352 (N_7352,N_3405,N_3962);
nand U7353 (N_7353,N_3460,N_1326);
nand U7354 (N_7354,N_2765,N_2163);
or U7355 (N_7355,N_2347,N_1085);
or U7356 (N_7356,N_4223,N_1967);
and U7357 (N_7357,N_2448,N_2338);
and U7358 (N_7358,N_953,N_3976);
nand U7359 (N_7359,N_3294,N_1823);
or U7360 (N_7360,N_3144,N_1485);
nand U7361 (N_7361,N_3872,N_3351);
nor U7362 (N_7362,N_1710,N_4744);
nand U7363 (N_7363,N_1322,N_3025);
or U7364 (N_7364,N_924,N_3141);
and U7365 (N_7365,N_3341,N_730);
nor U7366 (N_7366,N_620,N_4089);
and U7367 (N_7367,N_3900,N_2507);
nor U7368 (N_7368,N_4964,N_2323);
nor U7369 (N_7369,N_1745,N_3326);
nor U7370 (N_7370,N_3496,N_3963);
or U7371 (N_7371,N_643,N_4409);
or U7372 (N_7372,N_3754,N_2048);
and U7373 (N_7373,N_2601,N_4712);
nor U7374 (N_7374,N_1081,N_4462);
nor U7375 (N_7375,N_657,N_3730);
nor U7376 (N_7376,N_2434,N_1650);
nand U7377 (N_7377,N_829,N_4332);
nor U7378 (N_7378,N_1809,N_1011);
nor U7379 (N_7379,N_2557,N_2435);
and U7380 (N_7380,N_3585,N_573);
nand U7381 (N_7381,N_598,N_1951);
nor U7382 (N_7382,N_921,N_4731);
or U7383 (N_7383,N_4847,N_1584);
nor U7384 (N_7384,N_4250,N_515);
nor U7385 (N_7385,N_3472,N_4363);
and U7386 (N_7386,N_995,N_247);
nor U7387 (N_7387,N_169,N_4228);
or U7388 (N_7388,N_779,N_407);
nor U7389 (N_7389,N_4676,N_4854);
and U7390 (N_7390,N_4643,N_2333);
or U7391 (N_7391,N_4954,N_575);
nand U7392 (N_7392,N_3904,N_1763);
or U7393 (N_7393,N_1978,N_2965);
and U7394 (N_7394,N_4884,N_2794);
nor U7395 (N_7395,N_971,N_965);
and U7396 (N_7396,N_2487,N_1804);
nor U7397 (N_7397,N_1119,N_4701);
and U7398 (N_7398,N_4238,N_3959);
or U7399 (N_7399,N_1554,N_512);
or U7400 (N_7400,N_3185,N_1736);
or U7401 (N_7401,N_2443,N_2419);
nand U7402 (N_7402,N_864,N_1087);
nor U7403 (N_7403,N_4646,N_1199);
and U7404 (N_7404,N_566,N_59);
and U7405 (N_7405,N_1884,N_3283);
nand U7406 (N_7406,N_360,N_3168);
nor U7407 (N_7407,N_3410,N_525);
nor U7408 (N_7408,N_3824,N_3045);
nor U7409 (N_7409,N_1730,N_1724);
nand U7410 (N_7410,N_3733,N_3516);
nand U7411 (N_7411,N_3101,N_2440);
or U7412 (N_7412,N_3749,N_2614);
and U7413 (N_7413,N_382,N_3358);
and U7414 (N_7414,N_1047,N_4563);
nor U7415 (N_7415,N_2950,N_2554);
nor U7416 (N_7416,N_909,N_4808);
nand U7417 (N_7417,N_1108,N_2757);
nor U7418 (N_7418,N_2962,N_3924);
and U7419 (N_7419,N_4262,N_2631);
or U7420 (N_7420,N_1414,N_173);
xor U7421 (N_7421,N_2414,N_3885);
nor U7422 (N_7422,N_2547,N_834);
nand U7423 (N_7423,N_354,N_1213);
and U7424 (N_7424,N_4855,N_3980);
nor U7425 (N_7425,N_478,N_2943);
or U7426 (N_7426,N_4576,N_595);
and U7427 (N_7427,N_670,N_438);
nor U7428 (N_7428,N_1904,N_2632);
nor U7429 (N_7429,N_592,N_4706);
nand U7430 (N_7430,N_3139,N_4485);
nor U7431 (N_7431,N_2156,N_1107);
and U7432 (N_7432,N_4549,N_3493);
and U7433 (N_7433,N_2028,N_3035);
and U7434 (N_7434,N_1130,N_3837);
and U7435 (N_7435,N_1385,N_2300);
and U7436 (N_7436,N_1538,N_2002);
nand U7437 (N_7437,N_3560,N_3725);
nor U7438 (N_7438,N_3913,N_134);
and U7439 (N_7439,N_519,N_4342);
nand U7440 (N_7440,N_2879,N_16);
nand U7441 (N_7441,N_4252,N_4837);
or U7442 (N_7442,N_2811,N_3488);
or U7443 (N_7443,N_3043,N_4433);
or U7444 (N_7444,N_1039,N_1101);
nor U7445 (N_7445,N_2523,N_4650);
and U7446 (N_7446,N_1312,N_2328);
and U7447 (N_7447,N_3626,N_4506);
and U7448 (N_7448,N_1454,N_4416);
nor U7449 (N_7449,N_1200,N_3015);
and U7450 (N_7450,N_1077,N_603);
and U7451 (N_7451,N_3510,N_1166);
nor U7452 (N_7452,N_3971,N_116);
nor U7453 (N_7453,N_2742,N_2182);
or U7454 (N_7454,N_1412,N_996);
and U7455 (N_7455,N_3941,N_2675);
nand U7456 (N_7456,N_825,N_3317);
nand U7457 (N_7457,N_1146,N_3952);
and U7458 (N_7458,N_1067,N_2819);
and U7459 (N_7459,N_1366,N_296);
nor U7460 (N_7460,N_4582,N_569);
or U7461 (N_7461,N_3536,N_4385);
or U7462 (N_7462,N_3643,N_2649);
nand U7463 (N_7463,N_4100,N_1501);
nand U7464 (N_7464,N_1610,N_83);
nand U7465 (N_7465,N_4469,N_4249);
or U7466 (N_7466,N_2190,N_3207);
and U7467 (N_7467,N_3136,N_3116);
nand U7468 (N_7468,N_2864,N_4012);
nand U7469 (N_7469,N_661,N_2379);
nand U7470 (N_7470,N_3866,N_2124);
nor U7471 (N_7471,N_4666,N_2132);
or U7472 (N_7472,N_1127,N_1058);
or U7473 (N_7473,N_3361,N_4455);
or U7474 (N_7474,N_3182,N_2963);
nor U7475 (N_7475,N_4514,N_4755);
nand U7476 (N_7476,N_3286,N_4825);
nor U7477 (N_7477,N_1853,N_2873);
nand U7478 (N_7478,N_1983,N_3647);
nor U7479 (N_7479,N_193,N_2761);
nand U7480 (N_7480,N_3584,N_1527);
and U7481 (N_7481,N_3273,N_807);
nor U7482 (N_7482,N_400,N_2784);
or U7483 (N_7483,N_4987,N_4313);
and U7484 (N_7484,N_2464,N_3468);
and U7485 (N_7485,N_2172,N_3084);
nor U7486 (N_7486,N_2531,N_4180);
nand U7487 (N_7487,N_1677,N_2490);
nor U7488 (N_7488,N_1886,N_3299);
and U7489 (N_7489,N_4734,N_3055);
nor U7490 (N_7490,N_4845,N_4158);
and U7491 (N_7491,N_1298,N_2032);
nor U7492 (N_7492,N_122,N_2847);
nor U7493 (N_7493,N_4246,N_2753);
and U7494 (N_7494,N_3694,N_4697);
or U7495 (N_7495,N_3929,N_3761);
and U7496 (N_7496,N_2148,N_1267);
nand U7497 (N_7497,N_2436,N_4075);
or U7498 (N_7498,N_118,N_2459);
nand U7499 (N_7499,N_4815,N_3354);
and U7500 (N_7500,N_2349,N_4751);
nand U7501 (N_7501,N_629,N_638);
nor U7502 (N_7502,N_3513,N_1786);
and U7503 (N_7503,N_2397,N_4587);
and U7504 (N_7504,N_13,N_1722);
or U7505 (N_7505,N_3061,N_443);
nand U7506 (N_7506,N_1703,N_1863);
xnor U7507 (N_7507,N_2625,N_3514);
nand U7508 (N_7508,N_827,N_4494);
and U7509 (N_7509,N_2050,N_839);
nand U7510 (N_7510,N_1372,N_4422);
and U7511 (N_7511,N_2217,N_4377);
or U7512 (N_7512,N_4992,N_4943);
and U7513 (N_7513,N_1124,N_1759);
and U7514 (N_7514,N_458,N_4267);
nor U7515 (N_7515,N_2182,N_4014);
nand U7516 (N_7516,N_1723,N_3462);
nor U7517 (N_7517,N_264,N_4764);
nor U7518 (N_7518,N_566,N_2295);
and U7519 (N_7519,N_190,N_523);
and U7520 (N_7520,N_4616,N_382);
nor U7521 (N_7521,N_149,N_702);
and U7522 (N_7522,N_4484,N_188);
and U7523 (N_7523,N_363,N_3928);
nand U7524 (N_7524,N_3390,N_3200);
and U7525 (N_7525,N_1256,N_65);
and U7526 (N_7526,N_3735,N_2540);
or U7527 (N_7527,N_4955,N_4591);
nand U7528 (N_7528,N_3685,N_2292);
nor U7529 (N_7529,N_356,N_1974);
nor U7530 (N_7530,N_3560,N_4150);
and U7531 (N_7531,N_3889,N_1804);
or U7532 (N_7532,N_1496,N_3187);
and U7533 (N_7533,N_2671,N_113);
or U7534 (N_7534,N_464,N_4210);
xor U7535 (N_7535,N_4642,N_4110);
nor U7536 (N_7536,N_2459,N_516);
and U7537 (N_7537,N_1023,N_2516);
nor U7538 (N_7538,N_4218,N_2062);
nand U7539 (N_7539,N_4324,N_2662);
nor U7540 (N_7540,N_271,N_1298);
nor U7541 (N_7541,N_2724,N_2010);
nor U7542 (N_7542,N_2149,N_1908);
nand U7543 (N_7543,N_4514,N_1031);
nand U7544 (N_7544,N_4513,N_4191);
nor U7545 (N_7545,N_1546,N_2131);
nand U7546 (N_7546,N_826,N_978);
or U7547 (N_7547,N_1946,N_3911);
nor U7548 (N_7548,N_3795,N_302);
or U7549 (N_7549,N_1369,N_1880);
or U7550 (N_7550,N_4083,N_3100);
nor U7551 (N_7551,N_902,N_745);
or U7552 (N_7552,N_2132,N_1124);
nor U7553 (N_7553,N_3114,N_4974);
and U7554 (N_7554,N_4932,N_4987);
nor U7555 (N_7555,N_2898,N_2722);
nand U7556 (N_7556,N_4276,N_2596);
and U7557 (N_7557,N_3512,N_4390);
or U7558 (N_7558,N_1229,N_3263);
nand U7559 (N_7559,N_369,N_2562);
nand U7560 (N_7560,N_676,N_1706);
nor U7561 (N_7561,N_4918,N_2400);
or U7562 (N_7562,N_185,N_3507);
nand U7563 (N_7563,N_3838,N_1944);
nand U7564 (N_7564,N_2944,N_865);
and U7565 (N_7565,N_3258,N_3448);
nor U7566 (N_7566,N_765,N_2653);
or U7567 (N_7567,N_3612,N_4197);
and U7568 (N_7568,N_2626,N_3877);
and U7569 (N_7569,N_115,N_1127);
nor U7570 (N_7570,N_3037,N_4131);
or U7571 (N_7571,N_1488,N_3776);
nor U7572 (N_7572,N_2592,N_4551);
nand U7573 (N_7573,N_2552,N_3936);
or U7574 (N_7574,N_3729,N_1477);
nor U7575 (N_7575,N_1591,N_3054);
nor U7576 (N_7576,N_2619,N_401);
nand U7577 (N_7577,N_1018,N_1835);
and U7578 (N_7578,N_2363,N_4578);
nor U7579 (N_7579,N_1158,N_2316);
or U7580 (N_7580,N_4151,N_4254);
nor U7581 (N_7581,N_3880,N_3353);
nand U7582 (N_7582,N_2032,N_1512);
nor U7583 (N_7583,N_2226,N_1047);
nand U7584 (N_7584,N_943,N_1766);
nor U7585 (N_7585,N_2292,N_2464);
and U7586 (N_7586,N_1231,N_474);
or U7587 (N_7587,N_2533,N_2687);
nor U7588 (N_7588,N_4928,N_182);
nor U7589 (N_7589,N_2624,N_38);
or U7590 (N_7590,N_3519,N_2772);
and U7591 (N_7591,N_3855,N_1665);
nor U7592 (N_7592,N_3879,N_179);
or U7593 (N_7593,N_2298,N_3390);
and U7594 (N_7594,N_2461,N_895);
nor U7595 (N_7595,N_3481,N_1648);
nor U7596 (N_7596,N_4641,N_133);
nand U7597 (N_7597,N_207,N_1551);
or U7598 (N_7598,N_1642,N_2788);
or U7599 (N_7599,N_4554,N_2968);
and U7600 (N_7600,N_2166,N_1944);
nand U7601 (N_7601,N_4534,N_714);
or U7602 (N_7602,N_3278,N_173);
or U7603 (N_7603,N_1685,N_2913);
nand U7604 (N_7604,N_2806,N_4272);
and U7605 (N_7605,N_2561,N_4963);
and U7606 (N_7606,N_4184,N_2773);
nor U7607 (N_7607,N_2703,N_3579);
and U7608 (N_7608,N_1692,N_2303);
nor U7609 (N_7609,N_2917,N_2157);
or U7610 (N_7610,N_3795,N_3629);
nor U7611 (N_7611,N_4052,N_1317);
or U7612 (N_7612,N_2544,N_3208);
and U7613 (N_7613,N_3347,N_4440);
and U7614 (N_7614,N_1198,N_4113);
nor U7615 (N_7615,N_3011,N_1318);
and U7616 (N_7616,N_1906,N_2396);
or U7617 (N_7617,N_1761,N_4414);
and U7618 (N_7618,N_128,N_4150);
and U7619 (N_7619,N_4498,N_4930);
or U7620 (N_7620,N_2596,N_4261);
nand U7621 (N_7621,N_4162,N_3908);
nand U7622 (N_7622,N_368,N_1786);
and U7623 (N_7623,N_1670,N_3634);
and U7624 (N_7624,N_3471,N_245);
nor U7625 (N_7625,N_731,N_2119);
and U7626 (N_7626,N_3246,N_2922);
and U7627 (N_7627,N_4674,N_2180);
nand U7628 (N_7628,N_3215,N_4819);
and U7629 (N_7629,N_4126,N_3694);
and U7630 (N_7630,N_3640,N_3742);
and U7631 (N_7631,N_3282,N_2883);
nand U7632 (N_7632,N_1613,N_3558);
or U7633 (N_7633,N_197,N_1483);
and U7634 (N_7634,N_3382,N_1862);
or U7635 (N_7635,N_3646,N_4976);
and U7636 (N_7636,N_1481,N_1644);
nand U7637 (N_7637,N_2089,N_4417);
nand U7638 (N_7638,N_2078,N_1961);
nand U7639 (N_7639,N_3538,N_4361);
and U7640 (N_7640,N_4002,N_1082);
or U7641 (N_7641,N_2039,N_254);
nor U7642 (N_7642,N_3465,N_641);
nor U7643 (N_7643,N_1260,N_4860);
nor U7644 (N_7644,N_4501,N_230);
nand U7645 (N_7645,N_4994,N_4263);
and U7646 (N_7646,N_2200,N_2315);
nand U7647 (N_7647,N_748,N_4942);
and U7648 (N_7648,N_4369,N_3555);
and U7649 (N_7649,N_2440,N_1059);
or U7650 (N_7650,N_2523,N_1540);
or U7651 (N_7651,N_906,N_694);
xor U7652 (N_7652,N_2210,N_2261);
nand U7653 (N_7653,N_3119,N_3122);
and U7654 (N_7654,N_940,N_1695);
nor U7655 (N_7655,N_3727,N_4984);
nor U7656 (N_7656,N_83,N_517);
or U7657 (N_7657,N_3708,N_2946);
or U7658 (N_7658,N_2327,N_4421);
nand U7659 (N_7659,N_2232,N_3669);
nor U7660 (N_7660,N_3172,N_766);
nor U7661 (N_7661,N_3030,N_259);
nor U7662 (N_7662,N_3736,N_3115);
and U7663 (N_7663,N_423,N_2193);
and U7664 (N_7664,N_2035,N_2958);
nand U7665 (N_7665,N_1955,N_2411);
or U7666 (N_7666,N_3735,N_727);
nor U7667 (N_7667,N_2394,N_4964);
nand U7668 (N_7668,N_3055,N_231);
or U7669 (N_7669,N_2938,N_2516);
nand U7670 (N_7670,N_4217,N_1655);
and U7671 (N_7671,N_4205,N_997);
nor U7672 (N_7672,N_3539,N_3521);
nand U7673 (N_7673,N_524,N_4450);
nor U7674 (N_7674,N_4361,N_1058);
and U7675 (N_7675,N_3451,N_4304);
nand U7676 (N_7676,N_1779,N_3500);
nand U7677 (N_7677,N_2106,N_4969);
nand U7678 (N_7678,N_625,N_2701);
or U7679 (N_7679,N_3252,N_1202);
or U7680 (N_7680,N_1504,N_2680);
and U7681 (N_7681,N_4375,N_2052);
or U7682 (N_7682,N_1972,N_2412);
nand U7683 (N_7683,N_248,N_1352);
or U7684 (N_7684,N_1107,N_434);
or U7685 (N_7685,N_1050,N_4259);
nor U7686 (N_7686,N_3241,N_2418);
nand U7687 (N_7687,N_874,N_4135);
nand U7688 (N_7688,N_971,N_3440);
nand U7689 (N_7689,N_1573,N_2198);
nor U7690 (N_7690,N_1055,N_2853);
nor U7691 (N_7691,N_1408,N_3816);
nand U7692 (N_7692,N_3437,N_3251);
xnor U7693 (N_7693,N_696,N_2884);
nor U7694 (N_7694,N_1356,N_4740);
nor U7695 (N_7695,N_4830,N_4664);
xnor U7696 (N_7696,N_4620,N_4036);
or U7697 (N_7697,N_3351,N_1788);
and U7698 (N_7698,N_4170,N_2551);
nand U7699 (N_7699,N_1284,N_3326);
nor U7700 (N_7700,N_1388,N_2491);
and U7701 (N_7701,N_4885,N_3610);
or U7702 (N_7702,N_3949,N_4439);
nor U7703 (N_7703,N_421,N_4079);
or U7704 (N_7704,N_3747,N_2765);
nor U7705 (N_7705,N_1059,N_50);
and U7706 (N_7706,N_2851,N_2802);
and U7707 (N_7707,N_4441,N_3381);
nand U7708 (N_7708,N_4800,N_4330);
or U7709 (N_7709,N_2456,N_1079);
nand U7710 (N_7710,N_3097,N_2508);
and U7711 (N_7711,N_1966,N_3227);
nor U7712 (N_7712,N_3196,N_524);
and U7713 (N_7713,N_3369,N_3083);
nand U7714 (N_7714,N_3513,N_4307);
and U7715 (N_7715,N_1015,N_2513);
nand U7716 (N_7716,N_4284,N_135);
nand U7717 (N_7717,N_4237,N_1992);
and U7718 (N_7718,N_372,N_3582);
and U7719 (N_7719,N_1343,N_779);
nor U7720 (N_7720,N_3969,N_3856);
nor U7721 (N_7721,N_4586,N_3435);
nor U7722 (N_7722,N_1231,N_2991);
and U7723 (N_7723,N_3970,N_4316);
and U7724 (N_7724,N_1846,N_4330);
nand U7725 (N_7725,N_13,N_3051);
nand U7726 (N_7726,N_925,N_4050);
and U7727 (N_7727,N_605,N_3214);
nor U7728 (N_7728,N_1253,N_1274);
and U7729 (N_7729,N_4224,N_4552);
nor U7730 (N_7730,N_908,N_2336);
nor U7731 (N_7731,N_3077,N_2282);
nand U7732 (N_7732,N_3635,N_3207);
or U7733 (N_7733,N_3315,N_1708);
nand U7734 (N_7734,N_187,N_250);
nor U7735 (N_7735,N_4236,N_2624);
and U7736 (N_7736,N_2656,N_1096);
nor U7737 (N_7737,N_1219,N_3454);
nand U7738 (N_7738,N_2514,N_490);
nor U7739 (N_7739,N_3006,N_469);
or U7740 (N_7740,N_3183,N_3962);
and U7741 (N_7741,N_1999,N_2263);
nand U7742 (N_7742,N_2809,N_2801);
nor U7743 (N_7743,N_3102,N_64);
nand U7744 (N_7744,N_101,N_492);
nand U7745 (N_7745,N_2019,N_118);
or U7746 (N_7746,N_2675,N_4181);
nand U7747 (N_7747,N_2313,N_1835);
nor U7748 (N_7748,N_24,N_4191);
or U7749 (N_7749,N_1609,N_162);
nand U7750 (N_7750,N_2147,N_2954);
nand U7751 (N_7751,N_3401,N_2361);
nor U7752 (N_7752,N_3179,N_1975);
and U7753 (N_7753,N_2353,N_4563);
or U7754 (N_7754,N_80,N_4583);
and U7755 (N_7755,N_3031,N_1059);
or U7756 (N_7756,N_1333,N_1386);
or U7757 (N_7757,N_3613,N_678);
or U7758 (N_7758,N_760,N_1374);
or U7759 (N_7759,N_4384,N_4594);
or U7760 (N_7760,N_963,N_3087);
nand U7761 (N_7761,N_2856,N_937);
and U7762 (N_7762,N_915,N_1538);
or U7763 (N_7763,N_4804,N_3882);
nand U7764 (N_7764,N_131,N_368);
nand U7765 (N_7765,N_2825,N_956);
nor U7766 (N_7766,N_2608,N_2942);
nor U7767 (N_7767,N_3541,N_868);
or U7768 (N_7768,N_907,N_1958);
or U7769 (N_7769,N_2757,N_2818);
or U7770 (N_7770,N_2846,N_4240);
nor U7771 (N_7771,N_4788,N_772);
and U7772 (N_7772,N_1419,N_1435);
and U7773 (N_7773,N_3378,N_2682);
and U7774 (N_7774,N_1455,N_3623);
nor U7775 (N_7775,N_2505,N_3509);
and U7776 (N_7776,N_2798,N_2353);
nor U7777 (N_7777,N_2175,N_2159);
nor U7778 (N_7778,N_2589,N_3730);
xnor U7779 (N_7779,N_232,N_1757);
nand U7780 (N_7780,N_3686,N_480);
nor U7781 (N_7781,N_1906,N_1407);
or U7782 (N_7782,N_658,N_39);
nand U7783 (N_7783,N_2071,N_742);
nand U7784 (N_7784,N_779,N_3844);
nand U7785 (N_7785,N_3592,N_3134);
nor U7786 (N_7786,N_1638,N_1631);
and U7787 (N_7787,N_387,N_3736);
nor U7788 (N_7788,N_1505,N_4923);
nand U7789 (N_7789,N_3455,N_4222);
nand U7790 (N_7790,N_3153,N_4076);
or U7791 (N_7791,N_1440,N_390);
and U7792 (N_7792,N_4974,N_3151);
or U7793 (N_7793,N_220,N_1354);
nand U7794 (N_7794,N_4027,N_1916);
nor U7795 (N_7795,N_3166,N_3368);
nand U7796 (N_7796,N_1683,N_4940);
and U7797 (N_7797,N_2111,N_356);
nand U7798 (N_7798,N_1967,N_1642);
and U7799 (N_7799,N_1959,N_3459);
and U7800 (N_7800,N_4478,N_1388);
nor U7801 (N_7801,N_3405,N_2581);
nand U7802 (N_7802,N_3670,N_2407);
nor U7803 (N_7803,N_356,N_3151);
and U7804 (N_7804,N_2480,N_972);
nor U7805 (N_7805,N_181,N_3614);
and U7806 (N_7806,N_2512,N_1588);
nand U7807 (N_7807,N_4096,N_3250);
or U7808 (N_7808,N_759,N_629);
nand U7809 (N_7809,N_3712,N_3658);
or U7810 (N_7810,N_2805,N_2310);
and U7811 (N_7811,N_3706,N_1421);
and U7812 (N_7812,N_1281,N_3022);
nor U7813 (N_7813,N_3483,N_2064);
and U7814 (N_7814,N_368,N_2268);
xor U7815 (N_7815,N_2965,N_2654);
nand U7816 (N_7816,N_2825,N_3160);
or U7817 (N_7817,N_4309,N_4227);
or U7818 (N_7818,N_940,N_855);
and U7819 (N_7819,N_359,N_2204);
nor U7820 (N_7820,N_1569,N_2343);
and U7821 (N_7821,N_1306,N_1640);
nand U7822 (N_7822,N_658,N_3133);
and U7823 (N_7823,N_4718,N_4563);
nand U7824 (N_7824,N_257,N_4747);
nor U7825 (N_7825,N_2735,N_4512);
nand U7826 (N_7826,N_4254,N_1810);
or U7827 (N_7827,N_4927,N_1466);
or U7828 (N_7828,N_3254,N_4243);
nor U7829 (N_7829,N_850,N_2435);
nand U7830 (N_7830,N_3748,N_1466);
nor U7831 (N_7831,N_4382,N_4065);
or U7832 (N_7832,N_194,N_560);
or U7833 (N_7833,N_4096,N_2487);
or U7834 (N_7834,N_1558,N_4377);
or U7835 (N_7835,N_18,N_3070);
or U7836 (N_7836,N_2793,N_909);
nor U7837 (N_7837,N_3511,N_1749);
nor U7838 (N_7838,N_4579,N_1598);
or U7839 (N_7839,N_964,N_4515);
or U7840 (N_7840,N_3578,N_1248);
nand U7841 (N_7841,N_1735,N_1056);
or U7842 (N_7842,N_1801,N_4789);
nand U7843 (N_7843,N_61,N_3925);
nand U7844 (N_7844,N_4127,N_4354);
nand U7845 (N_7845,N_1517,N_2833);
nor U7846 (N_7846,N_4602,N_1118);
nor U7847 (N_7847,N_951,N_903);
nor U7848 (N_7848,N_1341,N_853);
and U7849 (N_7849,N_1587,N_1557);
nor U7850 (N_7850,N_1333,N_1330);
nor U7851 (N_7851,N_1726,N_67);
or U7852 (N_7852,N_4736,N_1325);
nand U7853 (N_7853,N_3622,N_2207);
nand U7854 (N_7854,N_3265,N_2728);
or U7855 (N_7855,N_608,N_2353);
and U7856 (N_7856,N_691,N_4131);
nor U7857 (N_7857,N_1371,N_2043);
nand U7858 (N_7858,N_668,N_617);
or U7859 (N_7859,N_1941,N_4262);
nor U7860 (N_7860,N_4804,N_283);
nor U7861 (N_7861,N_2277,N_1876);
and U7862 (N_7862,N_2762,N_2231);
and U7863 (N_7863,N_3917,N_4384);
or U7864 (N_7864,N_1656,N_610);
nor U7865 (N_7865,N_972,N_1783);
and U7866 (N_7866,N_2112,N_409);
nand U7867 (N_7867,N_1937,N_4071);
nor U7868 (N_7868,N_4012,N_4886);
and U7869 (N_7869,N_3007,N_2196);
and U7870 (N_7870,N_3090,N_4663);
and U7871 (N_7871,N_1500,N_4496);
nand U7872 (N_7872,N_1538,N_701);
nand U7873 (N_7873,N_245,N_728);
and U7874 (N_7874,N_298,N_3778);
nand U7875 (N_7875,N_1273,N_3015);
nor U7876 (N_7876,N_3785,N_1744);
nor U7877 (N_7877,N_4738,N_2148);
nand U7878 (N_7878,N_4077,N_4656);
or U7879 (N_7879,N_4349,N_39);
nor U7880 (N_7880,N_412,N_4627);
nand U7881 (N_7881,N_4108,N_4473);
nand U7882 (N_7882,N_1457,N_1844);
or U7883 (N_7883,N_2330,N_4127);
and U7884 (N_7884,N_2570,N_1456);
nor U7885 (N_7885,N_3738,N_962);
or U7886 (N_7886,N_2540,N_2181);
nand U7887 (N_7887,N_2074,N_1169);
or U7888 (N_7888,N_557,N_1305);
or U7889 (N_7889,N_604,N_2177);
and U7890 (N_7890,N_919,N_1321);
and U7891 (N_7891,N_3339,N_789);
or U7892 (N_7892,N_757,N_3621);
nor U7893 (N_7893,N_1964,N_2342);
nor U7894 (N_7894,N_2595,N_141);
or U7895 (N_7895,N_4585,N_4419);
nor U7896 (N_7896,N_2846,N_2303);
and U7897 (N_7897,N_2253,N_935);
or U7898 (N_7898,N_4556,N_2071);
nor U7899 (N_7899,N_807,N_817);
nand U7900 (N_7900,N_4039,N_4290);
nand U7901 (N_7901,N_1944,N_2617);
nand U7902 (N_7902,N_2207,N_834);
nor U7903 (N_7903,N_2525,N_4792);
and U7904 (N_7904,N_3239,N_1182);
nor U7905 (N_7905,N_2670,N_2313);
and U7906 (N_7906,N_3176,N_2433);
or U7907 (N_7907,N_988,N_4526);
or U7908 (N_7908,N_4996,N_4482);
nand U7909 (N_7909,N_2869,N_3013);
or U7910 (N_7910,N_64,N_4809);
nor U7911 (N_7911,N_1540,N_4279);
or U7912 (N_7912,N_265,N_3719);
nor U7913 (N_7913,N_221,N_3541);
nand U7914 (N_7914,N_1395,N_1867);
nor U7915 (N_7915,N_2741,N_225);
nand U7916 (N_7916,N_1710,N_114);
nand U7917 (N_7917,N_800,N_3726);
nor U7918 (N_7918,N_475,N_692);
or U7919 (N_7919,N_173,N_4967);
or U7920 (N_7920,N_548,N_4538);
nand U7921 (N_7921,N_2593,N_1667);
and U7922 (N_7922,N_4182,N_868);
nor U7923 (N_7923,N_4953,N_3354);
nand U7924 (N_7924,N_4878,N_2869);
nor U7925 (N_7925,N_4783,N_4156);
and U7926 (N_7926,N_1435,N_656);
nor U7927 (N_7927,N_3247,N_637);
and U7928 (N_7928,N_2444,N_2655);
nor U7929 (N_7929,N_1719,N_1112);
nor U7930 (N_7930,N_2834,N_1880);
or U7931 (N_7931,N_1315,N_2620);
xor U7932 (N_7932,N_2038,N_2192);
or U7933 (N_7933,N_4253,N_4731);
nand U7934 (N_7934,N_581,N_3189);
nor U7935 (N_7935,N_1915,N_3750);
and U7936 (N_7936,N_3799,N_3870);
nand U7937 (N_7937,N_3075,N_206);
or U7938 (N_7938,N_1235,N_2885);
nor U7939 (N_7939,N_1349,N_1213);
or U7940 (N_7940,N_1162,N_1893);
nor U7941 (N_7941,N_995,N_3763);
nor U7942 (N_7942,N_3506,N_2074);
or U7943 (N_7943,N_4108,N_736);
or U7944 (N_7944,N_230,N_3355);
and U7945 (N_7945,N_506,N_4602);
nand U7946 (N_7946,N_1087,N_3784);
xor U7947 (N_7947,N_3100,N_1297);
and U7948 (N_7948,N_322,N_931);
or U7949 (N_7949,N_326,N_984);
nand U7950 (N_7950,N_3264,N_746);
nand U7951 (N_7951,N_167,N_1070);
or U7952 (N_7952,N_1070,N_4220);
nor U7953 (N_7953,N_272,N_427);
nand U7954 (N_7954,N_1399,N_955);
or U7955 (N_7955,N_1018,N_281);
or U7956 (N_7956,N_3801,N_2805);
nor U7957 (N_7957,N_4711,N_4328);
nand U7958 (N_7958,N_1664,N_1151);
nor U7959 (N_7959,N_3031,N_3126);
or U7960 (N_7960,N_755,N_611);
and U7961 (N_7961,N_4347,N_3431);
nand U7962 (N_7962,N_125,N_3672);
nor U7963 (N_7963,N_819,N_1465);
nand U7964 (N_7964,N_4569,N_1283);
or U7965 (N_7965,N_4002,N_3669);
or U7966 (N_7966,N_3893,N_26);
nor U7967 (N_7967,N_2949,N_3704);
or U7968 (N_7968,N_1343,N_1623);
nor U7969 (N_7969,N_1487,N_2326);
nand U7970 (N_7970,N_3541,N_2614);
nand U7971 (N_7971,N_1454,N_4206);
and U7972 (N_7972,N_3187,N_681);
nor U7973 (N_7973,N_3041,N_1723);
or U7974 (N_7974,N_2963,N_2538);
and U7975 (N_7975,N_2089,N_3951);
or U7976 (N_7976,N_2088,N_580);
nand U7977 (N_7977,N_4827,N_1182);
or U7978 (N_7978,N_1485,N_2366);
nor U7979 (N_7979,N_3811,N_4457);
and U7980 (N_7980,N_2216,N_1180);
and U7981 (N_7981,N_414,N_1716);
nand U7982 (N_7982,N_2646,N_3288);
or U7983 (N_7983,N_1282,N_660);
or U7984 (N_7984,N_2871,N_3774);
and U7985 (N_7985,N_3070,N_3778);
and U7986 (N_7986,N_690,N_1875);
and U7987 (N_7987,N_1046,N_3294);
or U7988 (N_7988,N_1874,N_1033);
nand U7989 (N_7989,N_1185,N_3813);
or U7990 (N_7990,N_3367,N_4994);
and U7991 (N_7991,N_1734,N_4769);
or U7992 (N_7992,N_2810,N_3467);
nand U7993 (N_7993,N_3066,N_1841);
nor U7994 (N_7994,N_1340,N_4656);
nand U7995 (N_7995,N_2169,N_3731);
nand U7996 (N_7996,N_2499,N_3770);
nor U7997 (N_7997,N_1216,N_4632);
or U7998 (N_7998,N_3315,N_3558);
and U7999 (N_7999,N_1639,N_1853);
and U8000 (N_8000,N_422,N_302);
nand U8001 (N_8001,N_2912,N_3443);
or U8002 (N_8002,N_4222,N_1294);
nand U8003 (N_8003,N_2808,N_2691);
or U8004 (N_8004,N_401,N_748);
nor U8005 (N_8005,N_1322,N_4751);
nand U8006 (N_8006,N_3707,N_986);
and U8007 (N_8007,N_551,N_656);
and U8008 (N_8008,N_566,N_1822);
nand U8009 (N_8009,N_2519,N_2057);
and U8010 (N_8010,N_2850,N_4786);
and U8011 (N_8011,N_1864,N_465);
and U8012 (N_8012,N_3874,N_2958);
and U8013 (N_8013,N_3916,N_929);
nor U8014 (N_8014,N_1490,N_3441);
and U8015 (N_8015,N_2961,N_1463);
or U8016 (N_8016,N_74,N_1720);
nand U8017 (N_8017,N_1624,N_1566);
or U8018 (N_8018,N_2515,N_1616);
nand U8019 (N_8019,N_2717,N_4365);
and U8020 (N_8020,N_671,N_4987);
and U8021 (N_8021,N_838,N_3745);
nor U8022 (N_8022,N_4119,N_4393);
nor U8023 (N_8023,N_990,N_3930);
nand U8024 (N_8024,N_4651,N_393);
nand U8025 (N_8025,N_4207,N_596);
nor U8026 (N_8026,N_3218,N_3391);
and U8027 (N_8027,N_9,N_3768);
nor U8028 (N_8028,N_4625,N_710);
and U8029 (N_8029,N_169,N_572);
nor U8030 (N_8030,N_1035,N_3125);
and U8031 (N_8031,N_4211,N_2507);
nor U8032 (N_8032,N_1204,N_558);
nand U8033 (N_8033,N_3361,N_2595);
or U8034 (N_8034,N_4595,N_3802);
and U8035 (N_8035,N_3024,N_1050);
or U8036 (N_8036,N_2753,N_2367);
nor U8037 (N_8037,N_2949,N_3715);
nor U8038 (N_8038,N_4061,N_3276);
and U8039 (N_8039,N_2422,N_31);
nor U8040 (N_8040,N_2231,N_1387);
nand U8041 (N_8041,N_4295,N_3034);
and U8042 (N_8042,N_3604,N_2131);
nor U8043 (N_8043,N_913,N_800);
or U8044 (N_8044,N_2337,N_3605);
nand U8045 (N_8045,N_2494,N_433);
nor U8046 (N_8046,N_2195,N_2783);
nand U8047 (N_8047,N_1732,N_4493);
and U8048 (N_8048,N_1713,N_2082);
and U8049 (N_8049,N_3165,N_1733);
or U8050 (N_8050,N_1459,N_3584);
nor U8051 (N_8051,N_4677,N_304);
nor U8052 (N_8052,N_957,N_4809);
nand U8053 (N_8053,N_3307,N_3224);
nor U8054 (N_8054,N_377,N_195);
and U8055 (N_8055,N_4390,N_2426);
nand U8056 (N_8056,N_231,N_2686);
and U8057 (N_8057,N_4683,N_2347);
nor U8058 (N_8058,N_1618,N_3158);
nand U8059 (N_8059,N_4656,N_3481);
and U8060 (N_8060,N_473,N_3809);
or U8061 (N_8061,N_96,N_1214);
or U8062 (N_8062,N_3773,N_1009);
nand U8063 (N_8063,N_4895,N_4084);
nor U8064 (N_8064,N_4269,N_3010);
or U8065 (N_8065,N_348,N_197);
and U8066 (N_8066,N_1341,N_1372);
xor U8067 (N_8067,N_2155,N_1556);
nand U8068 (N_8068,N_1762,N_4464);
nand U8069 (N_8069,N_2995,N_1680);
or U8070 (N_8070,N_3296,N_4429);
and U8071 (N_8071,N_3556,N_3533);
xnor U8072 (N_8072,N_4545,N_2941);
nand U8073 (N_8073,N_4924,N_4074);
and U8074 (N_8074,N_2319,N_3504);
nand U8075 (N_8075,N_1,N_3331);
nand U8076 (N_8076,N_1330,N_1420);
or U8077 (N_8077,N_1577,N_3620);
or U8078 (N_8078,N_2417,N_4255);
and U8079 (N_8079,N_3461,N_3542);
nor U8080 (N_8080,N_664,N_147);
nand U8081 (N_8081,N_949,N_2767);
nand U8082 (N_8082,N_4003,N_4143);
or U8083 (N_8083,N_934,N_3563);
and U8084 (N_8084,N_4499,N_1843);
or U8085 (N_8085,N_2413,N_1152);
or U8086 (N_8086,N_212,N_3021);
and U8087 (N_8087,N_806,N_3495);
or U8088 (N_8088,N_3981,N_2148);
and U8089 (N_8089,N_1544,N_1922);
nand U8090 (N_8090,N_3069,N_2876);
nor U8091 (N_8091,N_2206,N_913);
nand U8092 (N_8092,N_3955,N_2294);
nor U8093 (N_8093,N_1034,N_2261);
and U8094 (N_8094,N_114,N_1468);
and U8095 (N_8095,N_2540,N_1435);
or U8096 (N_8096,N_1587,N_3662);
nand U8097 (N_8097,N_4057,N_2421);
and U8098 (N_8098,N_3038,N_947);
nand U8099 (N_8099,N_512,N_4941);
or U8100 (N_8100,N_1419,N_1651);
nand U8101 (N_8101,N_1127,N_2493);
nor U8102 (N_8102,N_2261,N_902);
and U8103 (N_8103,N_2747,N_1259);
nand U8104 (N_8104,N_1994,N_412);
nor U8105 (N_8105,N_4824,N_28);
nor U8106 (N_8106,N_2619,N_4756);
nor U8107 (N_8107,N_1433,N_4114);
nand U8108 (N_8108,N_1040,N_3883);
and U8109 (N_8109,N_3936,N_3280);
nand U8110 (N_8110,N_1465,N_2244);
xnor U8111 (N_8111,N_1182,N_3693);
or U8112 (N_8112,N_297,N_1770);
nand U8113 (N_8113,N_522,N_4079);
and U8114 (N_8114,N_3909,N_1434);
and U8115 (N_8115,N_2237,N_3085);
or U8116 (N_8116,N_2311,N_2711);
nand U8117 (N_8117,N_2799,N_384);
and U8118 (N_8118,N_875,N_3197);
or U8119 (N_8119,N_2950,N_3473);
and U8120 (N_8120,N_3906,N_4494);
nor U8121 (N_8121,N_2381,N_2171);
nand U8122 (N_8122,N_4367,N_3519);
nand U8123 (N_8123,N_1894,N_3001);
nand U8124 (N_8124,N_107,N_1487);
or U8125 (N_8125,N_1483,N_4030);
nand U8126 (N_8126,N_4442,N_4120);
nand U8127 (N_8127,N_66,N_1793);
and U8128 (N_8128,N_820,N_2775);
nor U8129 (N_8129,N_4731,N_1903);
nand U8130 (N_8130,N_2041,N_1124);
nand U8131 (N_8131,N_3714,N_268);
nor U8132 (N_8132,N_3764,N_4094);
nand U8133 (N_8133,N_1386,N_18);
and U8134 (N_8134,N_1705,N_2331);
nand U8135 (N_8135,N_1678,N_1390);
nand U8136 (N_8136,N_512,N_2161);
nand U8137 (N_8137,N_1245,N_1913);
nand U8138 (N_8138,N_2212,N_2121);
and U8139 (N_8139,N_2794,N_4268);
nor U8140 (N_8140,N_815,N_3174);
and U8141 (N_8141,N_3773,N_4820);
nor U8142 (N_8142,N_2021,N_3530);
and U8143 (N_8143,N_1998,N_2214);
nor U8144 (N_8144,N_1556,N_4969);
or U8145 (N_8145,N_1461,N_3975);
and U8146 (N_8146,N_2173,N_2240);
or U8147 (N_8147,N_2011,N_2543);
and U8148 (N_8148,N_4617,N_4808);
or U8149 (N_8149,N_3293,N_4887);
or U8150 (N_8150,N_655,N_1049);
nand U8151 (N_8151,N_808,N_4208);
or U8152 (N_8152,N_440,N_4172);
and U8153 (N_8153,N_2901,N_4732);
nand U8154 (N_8154,N_1388,N_990);
or U8155 (N_8155,N_3257,N_2575);
nand U8156 (N_8156,N_3421,N_707);
nor U8157 (N_8157,N_3427,N_172);
nand U8158 (N_8158,N_1211,N_90);
nor U8159 (N_8159,N_880,N_3448);
or U8160 (N_8160,N_4529,N_3962);
or U8161 (N_8161,N_618,N_1177);
nand U8162 (N_8162,N_4714,N_4816);
nor U8163 (N_8163,N_4097,N_2981);
nor U8164 (N_8164,N_4870,N_4799);
and U8165 (N_8165,N_3463,N_3547);
and U8166 (N_8166,N_1527,N_3634);
nand U8167 (N_8167,N_2802,N_366);
nand U8168 (N_8168,N_2476,N_3929);
nor U8169 (N_8169,N_823,N_3866);
nor U8170 (N_8170,N_2871,N_3729);
nor U8171 (N_8171,N_3054,N_4607);
or U8172 (N_8172,N_2754,N_998);
nand U8173 (N_8173,N_3898,N_2234);
nor U8174 (N_8174,N_318,N_4570);
nor U8175 (N_8175,N_3855,N_1567);
and U8176 (N_8176,N_3770,N_1796);
nor U8177 (N_8177,N_1497,N_1654);
nand U8178 (N_8178,N_2833,N_249);
or U8179 (N_8179,N_1970,N_740);
xnor U8180 (N_8180,N_1172,N_164);
nor U8181 (N_8181,N_1841,N_2653);
nand U8182 (N_8182,N_3850,N_1865);
and U8183 (N_8183,N_1588,N_4139);
nor U8184 (N_8184,N_2553,N_16);
nand U8185 (N_8185,N_2054,N_132);
and U8186 (N_8186,N_1137,N_4005);
or U8187 (N_8187,N_288,N_3749);
and U8188 (N_8188,N_4023,N_2158);
and U8189 (N_8189,N_3203,N_3134);
xnor U8190 (N_8190,N_4491,N_2721);
and U8191 (N_8191,N_287,N_4370);
or U8192 (N_8192,N_641,N_4714);
nor U8193 (N_8193,N_4656,N_61);
or U8194 (N_8194,N_783,N_779);
or U8195 (N_8195,N_932,N_2952);
nor U8196 (N_8196,N_2290,N_1414);
nand U8197 (N_8197,N_4498,N_1568);
nand U8198 (N_8198,N_3427,N_2128);
and U8199 (N_8199,N_445,N_3719);
or U8200 (N_8200,N_1956,N_1288);
nor U8201 (N_8201,N_1079,N_3566);
and U8202 (N_8202,N_4908,N_636);
nand U8203 (N_8203,N_4014,N_3474);
nand U8204 (N_8204,N_4829,N_3378);
and U8205 (N_8205,N_1028,N_516);
and U8206 (N_8206,N_537,N_1630);
nand U8207 (N_8207,N_1854,N_2093);
and U8208 (N_8208,N_1962,N_4152);
nor U8209 (N_8209,N_2151,N_3173);
nor U8210 (N_8210,N_4085,N_3113);
or U8211 (N_8211,N_3236,N_774);
and U8212 (N_8212,N_4468,N_534);
and U8213 (N_8213,N_1644,N_1198);
nand U8214 (N_8214,N_3433,N_2761);
nor U8215 (N_8215,N_532,N_300);
nor U8216 (N_8216,N_1057,N_2794);
or U8217 (N_8217,N_4856,N_3487);
nand U8218 (N_8218,N_4570,N_1627);
nand U8219 (N_8219,N_2695,N_1667);
nand U8220 (N_8220,N_4440,N_2937);
and U8221 (N_8221,N_1289,N_363);
or U8222 (N_8222,N_927,N_3590);
nand U8223 (N_8223,N_2734,N_483);
and U8224 (N_8224,N_3675,N_4608);
nor U8225 (N_8225,N_793,N_2096);
or U8226 (N_8226,N_4476,N_3961);
nor U8227 (N_8227,N_2195,N_1856);
nand U8228 (N_8228,N_4187,N_716);
and U8229 (N_8229,N_4534,N_2149);
nor U8230 (N_8230,N_1694,N_342);
or U8231 (N_8231,N_733,N_4402);
or U8232 (N_8232,N_3492,N_584);
and U8233 (N_8233,N_3222,N_1308);
or U8234 (N_8234,N_1272,N_4939);
nand U8235 (N_8235,N_3747,N_3098);
nor U8236 (N_8236,N_3081,N_1529);
or U8237 (N_8237,N_4483,N_3983);
nor U8238 (N_8238,N_1562,N_2049);
and U8239 (N_8239,N_1685,N_4043);
or U8240 (N_8240,N_4022,N_2601);
nor U8241 (N_8241,N_4295,N_1173);
and U8242 (N_8242,N_1101,N_702);
and U8243 (N_8243,N_3094,N_4975);
and U8244 (N_8244,N_4438,N_2431);
nand U8245 (N_8245,N_449,N_723);
or U8246 (N_8246,N_4467,N_2961);
or U8247 (N_8247,N_3861,N_2604);
or U8248 (N_8248,N_4987,N_4482);
or U8249 (N_8249,N_3540,N_1189);
nor U8250 (N_8250,N_3898,N_4820);
nand U8251 (N_8251,N_1692,N_460);
nor U8252 (N_8252,N_1178,N_3121);
nor U8253 (N_8253,N_3122,N_4439);
nand U8254 (N_8254,N_2502,N_1018);
and U8255 (N_8255,N_116,N_221);
and U8256 (N_8256,N_2578,N_4316);
or U8257 (N_8257,N_845,N_3603);
and U8258 (N_8258,N_2660,N_1456);
and U8259 (N_8259,N_3979,N_1829);
nor U8260 (N_8260,N_4644,N_2691);
nand U8261 (N_8261,N_2327,N_4906);
nand U8262 (N_8262,N_4609,N_3700);
and U8263 (N_8263,N_100,N_2602);
nor U8264 (N_8264,N_3503,N_1752);
or U8265 (N_8265,N_3284,N_898);
and U8266 (N_8266,N_1939,N_1245);
nor U8267 (N_8267,N_4256,N_4314);
or U8268 (N_8268,N_3074,N_2889);
nor U8269 (N_8269,N_2229,N_1021);
and U8270 (N_8270,N_454,N_4929);
and U8271 (N_8271,N_4924,N_3420);
nand U8272 (N_8272,N_2776,N_4230);
and U8273 (N_8273,N_3541,N_701);
nor U8274 (N_8274,N_2074,N_2358);
and U8275 (N_8275,N_14,N_3578);
nor U8276 (N_8276,N_3293,N_3857);
nor U8277 (N_8277,N_4642,N_2654);
nor U8278 (N_8278,N_2555,N_2773);
nor U8279 (N_8279,N_3521,N_439);
nand U8280 (N_8280,N_1609,N_839);
or U8281 (N_8281,N_1935,N_1953);
nand U8282 (N_8282,N_2036,N_3001);
or U8283 (N_8283,N_920,N_4639);
nor U8284 (N_8284,N_661,N_3909);
and U8285 (N_8285,N_2141,N_1693);
and U8286 (N_8286,N_1246,N_3057);
nor U8287 (N_8287,N_686,N_3644);
or U8288 (N_8288,N_532,N_3482);
or U8289 (N_8289,N_1357,N_1215);
nor U8290 (N_8290,N_768,N_1080);
nor U8291 (N_8291,N_922,N_834);
or U8292 (N_8292,N_4520,N_4020);
nand U8293 (N_8293,N_1771,N_1860);
or U8294 (N_8294,N_4471,N_3788);
nand U8295 (N_8295,N_4934,N_2820);
nand U8296 (N_8296,N_2923,N_4499);
nand U8297 (N_8297,N_699,N_238);
nand U8298 (N_8298,N_2026,N_2644);
and U8299 (N_8299,N_4477,N_766);
or U8300 (N_8300,N_1937,N_4731);
or U8301 (N_8301,N_1766,N_3797);
nor U8302 (N_8302,N_466,N_540);
or U8303 (N_8303,N_452,N_2441);
nor U8304 (N_8304,N_3086,N_2352);
nor U8305 (N_8305,N_3046,N_4491);
or U8306 (N_8306,N_1578,N_2172);
or U8307 (N_8307,N_1989,N_1164);
nand U8308 (N_8308,N_432,N_4294);
nor U8309 (N_8309,N_4476,N_709);
nand U8310 (N_8310,N_2052,N_4366);
nand U8311 (N_8311,N_1309,N_4616);
and U8312 (N_8312,N_3875,N_4164);
nand U8313 (N_8313,N_30,N_1246);
nand U8314 (N_8314,N_491,N_3991);
nor U8315 (N_8315,N_2427,N_2655);
or U8316 (N_8316,N_3910,N_3887);
nor U8317 (N_8317,N_1719,N_2876);
nor U8318 (N_8318,N_3250,N_4470);
or U8319 (N_8319,N_638,N_2228);
nand U8320 (N_8320,N_4578,N_4494);
and U8321 (N_8321,N_974,N_4341);
and U8322 (N_8322,N_2333,N_4531);
and U8323 (N_8323,N_1860,N_4257);
and U8324 (N_8324,N_2196,N_893);
nand U8325 (N_8325,N_809,N_3431);
and U8326 (N_8326,N_291,N_2874);
nand U8327 (N_8327,N_2539,N_2196);
xnor U8328 (N_8328,N_1669,N_1146);
nor U8329 (N_8329,N_4477,N_391);
or U8330 (N_8330,N_254,N_1400);
nor U8331 (N_8331,N_3472,N_1439);
and U8332 (N_8332,N_650,N_4900);
nand U8333 (N_8333,N_360,N_675);
and U8334 (N_8334,N_2473,N_2051);
nor U8335 (N_8335,N_4367,N_1509);
xnor U8336 (N_8336,N_4665,N_1686);
nor U8337 (N_8337,N_2221,N_4636);
and U8338 (N_8338,N_4143,N_4660);
nand U8339 (N_8339,N_536,N_2576);
and U8340 (N_8340,N_2246,N_1759);
and U8341 (N_8341,N_946,N_3675);
nor U8342 (N_8342,N_3301,N_2521);
xor U8343 (N_8343,N_3980,N_2886);
nor U8344 (N_8344,N_2997,N_749);
nand U8345 (N_8345,N_858,N_872);
or U8346 (N_8346,N_4910,N_702);
and U8347 (N_8347,N_1910,N_3688);
or U8348 (N_8348,N_962,N_3310);
nor U8349 (N_8349,N_443,N_4553);
or U8350 (N_8350,N_1918,N_2507);
or U8351 (N_8351,N_1521,N_21);
or U8352 (N_8352,N_274,N_154);
and U8353 (N_8353,N_758,N_4761);
and U8354 (N_8354,N_1465,N_4965);
and U8355 (N_8355,N_567,N_4468);
or U8356 (N_8356,N_1309,N_3058);
nand U8357 (N_8357,N_4815,N_1706);
nand U8358 (N_8358,N_2355,N_2535);
nand U8359 (N_8359,N_619,N_3788);
or U8360 (N_8360,N_2887,N_2158);
nor U8361 (N_8361,N_1632,N_1022);
nand U8362 (N_8362,N_1642,N_2003);
and U8363 (N_8363,N_3389,N_3831);
nor U8364 (N_8364,N_4196,N_1371);
or U8365 (N_8365,N_4925,N_1806);
and U8366 (N_8366,N_4029,N_117);
and U8367 (N_8367,N_3304,N_3131);
nor U8368 (N_8368,N_3147,N_4589);
or U8369 (N_8369,N_1296,N_2130);
nor U8370 (N_8370,N_2685,N_3882);
and U8371 (N_8371,N_3634,N_3004);
and U8372 (N_8372,N_4287,N_4893);
xor U8373 (N_8373,N_3622,N_2489);
and U8374 (N_8374,N_541,N_2228);
nor U8375 (N_8375,N_792,N_4727);
and U8376 (N_8376,N_4289,N_112);
or U8377 (N_8377,N_2424,N_1615);
or U8378 (N_8378,N_2829,N_4867);
or U8379 (N_8379,N_1524,N_4547);
nor U8380 (N_8380,N_3400,N_1493);
nor U8381 (N_8381,N_1521,N_1577);
nand U8382 (N_8382,N_86,N_2420);
or U8383 (N_8383,N_2011,N_4611);
or U8384 (N_8384,N_1667,N_2030);
and U8385 (N_8385,N_540,N_3746);
nand U8386 (N_8386,N_3962,N_4909);
nor U8387 (N_8387,N_1480,N_236);
nor U8388 (N_8388,N_221,N_458);
nand U8389 (N_8389,N_2182,N_4101);
xnor U8390 (N_8390,N_713,N_3090);
nor U8391 (N_8391,N_551,N_617);
nand U8392 (N_8392,N_3296,N_289);
nand U8393 (N_8393,N_228,N_1425);
and U8394 (N_8394,N_2236,N_3230);
nand U8395 (N_8395,N_2921,N_2239);
nor U8396 (N_8396,N_953,N_4938);
nor U8397 (N_8397,N_541,N_3049);
or U8398 (N_8398,N_498,N_3228);
or U8399 (N_8399,N_1159,N_1914);
nor U8400 (N_8400,N_673,N_3454);
or U8401 (N_8401,N_4108,N_4057);
or U8402 (N_8402,N_2616,N_986);
or U8403 (N_8403,N_583,N_4129);
nor U8404 (N_8404,N_4003,N_2966);
nor U8405 (N_8405,N_3328,N_53);
and U8406 (N_8406,N_4722,N_4521);
xor U8407 (N_8407,N_2148,N_3324);
and U8408 (N_8408,N_4938,N_4417);
and U8409 (N_8409,N_155,N_1946);
nand U8410 (N_8410,N_709,N_2245);
nand U8411 (N_8411,N_2543,N_1883);
and U8412 (N_8412,N_1001,N_3560);
and U8413 (N_8413,N_2478,N_628);
or U8414 (N_8414,N_1906,N_2212);
nand U8415 (N_8415,N_1057,N_3315);
nor U8416 (N_8416,N_3492,N_1605);
or U8417 (N_8417,N_2539,N_4735);
nor U8418 (N_8418,N_4132,N_3017);
and U8419 (N_8419,N_4849,N_115);
nor U8420 (N_8420,N_953,N_1208);
nand U8421 (N_8421,N_2808,N_2065);
and U8422 (N_8422,N_2208,N_4492);
or U8423 (N_8423,N_480,N_3823);
and U8424 (N_8424,N_3949,N_2334);
nor U8425 (N_8425,N_2651,N_1684);
and U8426 (N_8426,N_1101,N_695);
nand U8427 (N_8427,N_602,N_4911);
nor U8428 (N_8428,N_3985,N_2397);
nand U8429 (N_8429,N_632,N_3886);
nor U8430 (N_8430,N_4696,N_2383);
nand U8431 (N_8431,N_129,N_245);
or U8432 (N_8432,N_353,N_1074);
nor U8433 (N_8433,N_4603,N_1830);
or U8434 (N_8434,N_833,N_2093);
nor U8435 (N_8435,N_1271,N_1461);
and U8436 (N_8436,N_1330,N_3869);
or U8437 (N_8437,N_1365,N_2176);
nand U8438 (N_8438,N_923,N_409);
or U8439 (N_8439,N_3688,N_4693);
xor U8440 (N_8440,N_217,N_4905);
nand U8441 (N_8441,N_3245,N_2121);
and U8442 (N_8442,N_4280,N_68);
and U8443 (N_8443,N_4530,N_4572);
nor U8444 (N_8444,N_3693,N_3562);
and U8445 (N_8445,N_1678,N_2190);
and U8446 (N_8446,N_455,N_1896);
or U8447 (N_8447,N_15,N_1049);
nand U8448 (N_8448,N_4724,N_2575);
xor U8449 (N_8449,N_3474,N_1001);
or U8450 (N_8450,N_4494,N_2368);
or U8451 (N_8451,N_4596,N_1391);
nor U8452 (N_8452,N_4369,N_3331);
and U8453 (N_8453,N_438,N_855);
nand U8454 (N_8454,N_3938,N_4389);
or U8455 (N_8455,N_3395,N_2692);
nand U8456 (N_8456,N_560,N_4659);
or U8457 (N_8457,N_4674,N_4388);
nand U8458 (N_8458,N_1520,N_288);
or U8459 (N_8459,N_4356,N_2847);
or U8460 (N_8460,N_415,N_355);
or U8461 (N_8461,N_3444,N_1821);
or U8462 (N_8462,N_3817,N_2123);
and U8463 (N_8463,N_469,N_1355);
nor U8464 (N_8464,N_2714,N_1197);
and U8465 (N_8465,N_4345,N_816);
and U8466 (N_8466,N_145,N_2430);
xnor U8467 (N_8467,N_1827,N_1672);
or U8468 (N_8468,N_2115,N_464);
nand U8469 (N_8469,N_3614,N_246);
and U8470 (N_8470,N_4695,N_554);
or U8471 (N_8471,N_2221,N_4433);
nand U8472 (N_8472,N_973,N_3515);
and U8473 (N_8473,N_4989,N_3491);
nor U8474 (N_8474,N_983,N_2036);
and U8475 (N_8475,N_809,N_81);
or U8476 (N_8476,N_1188,N_982);
nand U8477 (N_8477,N_2192,N_890);
nor U8478 (N_8478,N_4887,N_2215);
nand U8479 (N_8479,N_2499,N_1630);
nor U8480 (N_8480,N_470,N_4020);
nand U8481 (N_8481,N_1652,N_2309);
nand U8482 (N_8482,N_3372,N_988);
and U8483 (N_8483,N_1991,N_1144);
nand U8484 (N_8484,N_792,N_2045);
and U8485 (N_8485,N_3623,N_404);
and U8486 (N_8486,N_858,N_4520);
nand U8487 (N_8487,N_1227,N_415);
and U8488 (N_8488,N_3485,N_3656);
nor U8489 (N_8489,N_2336,N_2363);
and U8490 (N_8490,N_2081,N_1444);
nand U8491 (N_8491,N_3974,N_323);
and U8492 (N_8492,N_2780,N_2832);
nand U8493 (N_8493,N_1852,N_4788);
or U8494 (N_8494,N_4914,N_3258);
nor U8495 (N_8495,N_2917,N_1667);
and U8496 (N_8496,N_4852,N_4856);
or U8497 (N_8497,N_72,N_350);
xnor U8498 (N_8498,N_3309,N_1387);
nor U8499 (N_8499,N_3428,N_70);
and U8500 (N_8500,N_330,N_4020);
and U8501 (N_8501,N_2296,N_4312);
nand U8502 (N_8502,N_4963,N_2500);
nor U8503 (N_8503,N_4874,N_830);
and U8504 (N_8504,N_1297,N_89);
and U8505 (N_8505,N_4812,N_1198);
and U8506 (N_8506,N_3450,N_3763);
nand U8507 (N_8507,N_1894,N_2115);
and U8508 (N_8508,N_3649,N_1546);
nor U8509 (N_8509,N_1672,N_895);
or U8510 (N_8510,N_714,N_83);
nand U8511 (N_8511,N_2004,N_4369);
nor U8512 (N_8512,N_1902,N_3500);
and U8513 (N_8513,N_562,N_1725);
and U8514 (N_8514,N_2742,N_3226);
and U8515 (N_8515,N_2746,N_3174);
nor U8516 (N_8516,N_1858,N_3649);
or U8517 (N_8517,N_318,N_238);
nand U8518 (N_8518,N_4592,N_690);
nor U8519 (N_8519,N_3511,N_1049);
nand U8520 (N_8520,N_1806,N_4188);
nor U8521 (N_8521,N_4270,N_187);
nor U8522 (N_8522,N_721,N_2229);
and U8523 (N_8523,N_1722,N_1082);
or U8524 (N_8524,N_4222,N_4814);
or U8525 (N_8525,N_3846,N_4484);
and U8526 (N_8526,N_827,N_2068);
nor U8527 (N_8527,N_671,N_4977);
nor U8528 (N_8528,N_729,N_2541);
and U8529 (N_8529,N_2517,N_2418);
and U8530 (N_8530,N_3432,N_1819);
and U8531 (N_8531,N_3148,N_3309);
nor U8532 (N_8532,N_1962,N_4694);
and U8533 (N_8533,N_479,N_2201);
nand U8534 (N_8534,N_437,N_1197);
or U8535 (N_8535,N_172,N_316);
or U8536 (N_8536,N_3458,N_3376);
nand U8537 (N_8537,N_3546,N_2659);
or U8538 (N_8538,N_337,N_215);
nor U8539 (N_8539,N_1034,N_4287);
nand U8540 (N_8540,N_3598,N_4558);
nand U8541 (N_8541,N_4957,N_1926);
nand U8542 (N_8542,N_2784,N_2704);
or U8543 (N_8543,N_4742,N_3112);
nand U8544 (N_8544,N_1388,N_866);
nand U8545 (N_8545,N_3340,N_111);
and U8546 (N_8546,N_457,N_1882);
nor U8547 (N_8547,N_1694,N_821);
and U8548 (N_8548,N_2919,N_4817);
nand U8549 (N_8549,N_4316,N_4471);
nor U8550 (N_8550,N_2993,N_779);
nor U8551 (N_8551,N_2835,N_1705);
and U8552 (N_8552,N_1,N_4415);
and U8553 (N_8553,N_2566,N_376);
nand U8554 (N_8554,N_4739,N_1209);
and U8555 (N_8555,N_2897,N_2539);
or U8556 (N_8556,N_3771,N_766);
and U8557 (N_8557,N_2396,N_1351);
or U8558 (N_8558,N_1527,N_1458);
and U8559 (N_8559,N_3513,N_1014);
nand U8560 (N_8560,N_371,N_22);
or U8561 (N_8561,N_4318,N_1262);
and U8562 (N_8562,N_4776,N_4761);
and U8563 (N_8563,N_1459,N_3284);
nor U8564 (N_8564,N_426,N_1461);
nand U8565 (N_8565,N_3892,N_2758);
nor U8566 (N_8566,N_498,N_4568);
and U8567 (N_8567,N_3265,N_181);
nor U8568 (N_8568,N_63,N_2020);
nand U8569 (N_8569,N_2091,N_435);
or U8570 (N_8570,N_51,N_3644);
and U8571 (N_8571,N_4417,N_229);
nand U8572 (N_8572,N_2130,N_1363);
or U8573 (N_8573,N_2170,N_4447);
nor U8574 (N_8574,N_3452,N_3170);
or U8575 (N_8575,N_4091,N_2588);
nand U8576 (N_8576,N_2694,N_2212);
nand U8577 (N_8577,N_2172,N_1462);
or U8578 (N_8578,N_4010,N_866);
or U8579 (N_8579,N_3955,N_4858);
and U8580 (N_8580,N_1397,N_1356);
nand U8581 (N_8581,N_1193,N_276);
nand U8582 (N_8582,N_700,N_4471);
nand U8583 (N_8583,N_2370,N_4445);
nor U8584 (N_8584,N_443,N_2831);
nand U8585 (N_8585,N_3809,N_2942);
nor U8586 (N_8586,N_3864,N_4964);
nand U8587 (N_8587,N_2143,N_1850);
or U8588 (N_8588,N_3483,N_1415);
nand U8589 (N_8589,N_1378,N_527);
nand U8590 (N_8590,N_1527,N_2062);
and U8591 (N_8591,N_3292,N_1132);
nand U8592 (N_8592,N_2702,N_1271);
and U8593 (N_8593,N_3472,N_2206);
nand U8594 (N_8594,N_4443,N_3487);
nor U8595 (N_8595,N_811,N_4063);
or U8596 (N_8596,N_87,N_693);
nand U8597 (N_8597,N_4252,N_446);
and U8598 (N_8598,N_2007,N_2966);
nor U8599 (N_8599,N_4118,N_364);
or U8600 (N_8600,N_3050,N_691);
nand U8601 (N_8601,N_2376,N_1417);
nand U8602 (N_8602,N_4074,N_4218);
nor U8603 (N_8603,N_3751,N_1083);
nor U8604 (N_8604,N_68,N_4056);
or U8605 (N_8605,N_4576,N_4323);
nand U8606 (N_8606,N_3740,N_3401);
or U8607 (N_8607,N_264,N_708);
nand U8608 (N_8608,N_1708,N_3596);
or U8609 (N_8609,N_2724,N_2455);
nand U8610 (N_8610,N_1494,N_1818);
nand U8611 (N_8611,N_3104,N_3913);
and U8612 (N_8612,N_1766,N_104);
and U8613 (N_8613,N_3104,N_2280);
nor U8614 (N_8614,N_834,N_4853);
nand U8615 (N_8615,N_3644,N_2115);
nand U8616 (N_8616,N_2286,N_2475);
or U8617 (N_8617,N_3312,N_4459);
nand U8618 (N_8618,N_1772,N_1943);
nand U8619 (N_8619,N_123,N_3668);
nand U8620 (N_8620,N_1088,N_463);
and U8621 (N_8621,N_3587,N_4789);
and U8622 (N_8622,N_4183,N_4362);
or U8623 (N_8623,N_3408,N_4304);
nand U8624 (N_8624,N_1835,N_4650);
nand U8625 (N_8625,N_4988,N_1100);
and U8626 (N_8626,N_976,N_4497);
and U8627 (N_8627,N_4790,N_4282);
nand U8628 (N_8628,N_493,N_3845);
and U8629 (N_8629,N_4054,N_3252);
nand U8630 (N_8630,N_3342,N_384);
and U8631 (N_8631,N_4229,N_3586);
nand U8632 (N_8632,N_1289,N_4091);
nor U8633 (N_8633,N_2845,N_507);
and U8634 (N_8634,N_283,N_4304);
or U8635 (N_8635,N_1069,N_4969);
nor U8636 (N_8636,N_2168,N_1852);
nor U8637 (N_8637,N_4463,N_4263);
or U8638 (N_8638,N_2427,N_4544);
nand U8639 (N_8639,N_2027,N_4376);
or U8640 (N_8640,N_1862,N_344);
or U8641 (N_8641,N_2837,N_136);
nor U8642 (N_8642,N_2294,N_2488);
nor U8643 (N_8643,N_3061,N_3378);
nand U8644 (N_8644,N_3630,N_2826);
and U8645 (N_8645,N_1421,N_366);
nand U8646 (N_8646,N_4266,N_1904);
and U8647 (N_8647,N_1337,N_2027);
nor U8648 (N_8648,N_2683,N_4263);
and U8649 (N_8649,N_2300,N_1723);
nor U8650 (N_8650,N_112,N_3333);
or U8651 (N_8651,N_496,N_3359);
nor U8652 (N_8652,N_1051,N_1115);
or U8653 (N_8653,N_12,N_1172);
nand U8654 (N_8654,N_4132,N_3614);
or U8655 (N_8655,N_4347,N_1621);
nand U8656 (N_8656,N_4190,N_1318);
nor U8657 (N_8657,N_2375,N_1285);
or U8658 (N_8658,N_1661,N_3213);
or U8659 (N_8659,N_2241,N_269);
and U8660 (N_8660,N_1619,N_3971);
nor U8661 (N_8661,N_4074,N_3269);
and U8662 (N_8662,N_4926,N_3463);
or U8663 (N_8663,N_2022,N_115);
nor U8664 (N_8664,N_568,N_3671);
and U8665 (N_8665,N_1016,N_3340);
nand U8666 (N_8666,N_45,N_124);
nand U8667 (N_8667,N_2255,N_2302);
or U8668 (N_8668,N_4444,N_4259);
nor U8669 (N_8669,N_2499,N_3230);
and U8670 (N_8670,N_3756,N_4234);
and U8671 (N_8671,N_4247,N_3354);
nand U8672 (N_8672,N_514,N_2236);
nor U8673 (N_8673,N_2246,N_3382);
and U8674 (N_8674,N_2979,N_2630);
nor U8675 (N_8675,N_2957,N_2524);
and U8676 (N_8676,N_4037,N_1228);
and U8677 (N_8677,N_3807,N_3153);
nor U8678 (N_8678,N_2905,N_673);
nand U8679 (N_8679,N_3844,N_711);
or U8680 (N_8680,N_3324,N_4980);
nand U8681 (N_8681,N_3727,N_1667);
nand U8682 (N_8682,N_1094,N_2146);
nand U8683 (N_8683,N_817,N_4171);
nand U8684 (N_8684,N_3601,N_2982);
or U8685 (N_8685,N_3440,N_3202);
and U8686 (N_8686,N_3684,N_2864);
or U8687 (N_8687,N_2457,N_698);
nand U8688 (N_8688,N_714,N_3983);
xnor U8689 (N_8689,N_1927,N_3870);
or U8690 (N_8690,N_1603,N_4509);
nand U8691 (N_8691,N_4812,N_4719);
xnor U8692 (N_8692,N_1299,N_4076);
or U8693 (N_8693,N_4231,N_1744);
nor U8694 (N_8694,N_1072,N_4478);
nor U8695 (N_8695,N_2679,N_1546);
nand U8696 (N_8696,N_3710,N_1036);
nor U8697 (N_8697,N_4332,N_3609);
and U8698 (N_8698,N_1306,N_776);
nand U8699 (N_8699,N_1803,N_3306);
nand U8700 (N_8700,N_2544,N_1065);
nand U8701 (N_8701,N_322,N_914);
nand U8702 (N_8702,N_2297,N_1345);
or U8703 (N_8703,N_787,N_2016);
or U8704 (N_8704,N_4693,N_2079);
nor U8705 (N_8705,N_1626,N_1095);
nor U8706 (N_8706,N_2433,N_1872);
nand U8707 (N_8707,N_3511,N_4083);
or U8708 (N_8708,N_2774,N_3720);
or U8709 (N_8709,N_2464,N_4447);
and U8710 (N_8710,N_3034,N_2493);
nor U8711 (N_8711,N_1477,N_1442);
nor U8712 (N_8712,N_2715,N_4783);
and U8713 (N_8713,N_3307,N_2335);
or U8714 (N_8714,N_3165,N_1774);
or U8715 (N_8715,N_3304,N_2066);
nand U8716 (N_8716,N_4140,N_752);
nand U8717 (N_8717,N_2220,N_2984);
or U8718 (N_8718,N_1369,N_935);
and U8719 (N_8719,N_524,N_3350);
nor U8720 (N_8720,N_1968,N_2627);
nand U8721 (N_8721,N_4432,N_2648);
and U8722 (N_8722,N_4061,N_1178);
or U8723 (N_8723,N_4201,N_2421);
xnor U8724 (N_8724,N_1354,N_2073);
nand U8725 (N_8725,N_1532,N_750);
or U8726 (N_8726,N_1636,N_2707);
nand U8727 (N_8727,N_2858,N_999);
or U8728 (N_8728,N_4503,N_3464);
and U8729 (N_8729,N_475,N_2468);
nor U8730 (N_8730,N_1498,N_80);
or U8731 (N_8731,N_3787,N_4664);
or U8732 (N_8732,N_2167,N_4781);
nor U8733 (N_8733,N_4912,N_3709);
nor U8734 (N_8734,N_647,N_4476);
or U8735 (N_8735,N_2969,N_2480);
nor U8736 (N_8736,N_805,N_3672);
or U8737 (N_8737,N_2061,N_806);
and U8738 (N_8738,N_3485,N_2921);
or U8739 (N_8739,N_1557,N_4578);
and U8740 (N_8740,N_2511,N_230);
nor U8741 (N_8741,N_4224,N_3237);
nor U8742 (N_8742,N_1305,N_141);
and U8743 (N_8743,N_3107,N_1848);
nand U8744 (N_8744,N_234,N_3085);
nand U8745 (N_8745,N_2660,N_2434);
nand U8746 (N_8746,N_1203,N_1649);
nand U8747 (N_8747,N_4058,N_2967);
nand U8748 (N_8748,N_2275,N_678);
nand U8749 (N_8749,N_4738,N_192);
nand U8750 (N_8750,N_4628,N_2696);
or U8751 (N_8751,N_1926,N_2284);
nand U8752 (N_8752,N_3752,N_971);
and U8753 (N_8753,N_3099,N_4404);
or U8754 (N_8754,N_1438,N_4949);
nand U8755 (N_8755,N_4215,N_957);
nand U8756 (N_8756,N_3981,N_4392);
nand U8757 (N_8757,N_2233,N_2026);
or U8758 (N_8758,N_332,N_94);
or U8759 (N_8759,N_2173,N_450);
or U8760 (N_8760,N_3321,N_2256);
nand U8761 (N_8761,N_4881,N_4473);
or U8762 (N_8762,N_4035,N_2335);
nor U8763 (N_8763,N_1128,N_2593);
and U8764 (N_8764,N_3691,N_138);
or U8765 (N_8765,N_103,N_841);
and U8766 (N_8766,N_1138,N_4715);
nor U8767 (N_8767,N_4408,N_1118);
nand U8768 (N_8768,N_4025,N_217);
nand U8769 (N_8769,N_2997,N_4366);
nor U8770 (N_8770,N_980,N_1560);
and U8771 (N_8771,N_3184,N_254);
and U8772 (N_8772,N_1250,N_1306);
or U8773 (N_8773,N_3118,N_2342);
and U8774 (N_8774,N_2033,N_1094);
nand U8775 (N_8775,N_1343,N_868);
or U8776 (N_8776,N_2903,N_3845);
or U8777 (N_8777,N_3999,N_4087);
or U8778 (N_8778,N_1919,N_1583);
nand U8779 (N_8779,N_2636,N_3138);
nand U8780 (N_8780,N_1924,N_472);
and U8781 (N_8781,N_1575,N_1745);
nor U8782 (N_8782,N_3586,N_2769);
nand U8783 (N_8783,N_1693,N_614);
nand U8784 (N_8784,N_3827,N_4602);
nor U8785 (N_8785,N_750,N_2643);
or U8786 (N_8786,N_3992,N_3987);
and U8787 (N_8787,N_4874,N_3511);
nor U8788 (N_8788,N_4676,N_2848);
nor U8789 (N_8789,N_4980,N_1069);
or U8790 (N_8790,N_4564,N_4421);
or U8791 (N_8791,N_825,N_2994);
nand U8792 (N_8792,N_2945,N_736);
or U8793 (N_8793,N_3536,N_2161);
nor U8794 (N_8794,N_2619,N_2103);
and U8795 (N_8795,N_2813,N_3497);
or U8796 (N_8796,N_2411,N_1293);
or U8797 (N_8797,N_4586,N_1161);
nor U8798 (N_8798,N_4137,N_4689);
and U8799 (N_8799,N_1695,N_2508);
and U8800 (N_8800,N_2364,N_2819);
or U8801 (N_8801,N_2754,N_3659);
nand U8802 (N_8802,N_850,N_2054);
nor U8803 (N_8803,N_4616,N_2090);
nand U8804 (N_8804,N_1090,N_98);
and U8805 (N_8805,N_3620,N_2953);
and U8806 (N_8806,N_691,N_4885);
nand U8807 (N_8807,N_4517,N_179);
or U8808 (N_8808,N_4530,N_2364);
nor U8809 (N_8809,N_877,N_1909);
nand U8810 (N_8810,N_4685,N_3157);
and U8811 (N_8811,N_3947,N_1331);
and U8812 (N_8812,N_571,N_2299);
nand U8813 (N_8813,N_4048,N_1979);
nand U8814 (N_8814,N_1943,N_1025);
or U8815 (N_8815,N_2732,N_807);
or U8816 (N_8816,N_4688,N_1603);
and U8817 (N_8817,N_2622,N_2021);
and U8818 (N_8818,N_2342,N_4789);
nor U8819 (N_8819,N_2422,N_4048);
nor U8820 (N_8820,N_2409,N_3457);
nand U8821 (N_8821,N_2673,N_3693);
or U8822 (N_8822,N_4500,N_1516);
and U8823 (N_8823,N_4251,N_4359);
or U8824 (N_8824,N_2930,N_3635);
nand U8825 (N_8825,N_1536,N_4678);
and U8826 (N_8826,N_203,N_4637);
or U8827 (N_8827,N_1358,N_631);
nor U8828 (N_8828,N_3649,N_931);
and U8829 (N_8829,N_744,N_3925);
xor U8830 (N_8830,N_2257,N_261);
nand U8831 (N_8831,N_3806,N_3098);
nor U8832 (N_8832,N_450,N_4180);
nand U8833 (N_8833,N_3300,N_2148);
nand U8834 (N_8834,N_2018,N_2206);
and U8835 (N_8835,N_3128,N_1766);
nand U8836 (N_8836,N_1916,N_1320);
and U8837 (N_8837,N_2611,N_153);
nor U8838 (N_8838,N_2718,N_1419);
nor U8839 (N_8839,N_2461,N_1366);
or U8840 (N_8840,N_3600,N_4425);
nor U8841 (N_8841,N_4549,N_3247);
and U8842 (N_8842,N_1912,N_4137);
nand U8843 (N_8843,N_1281,N_2291);
nor U8844 (N_8844,N_4845,N_2164);
nand U8845 (N_8845,N_2301,N_3734);
and U8846 (N_8846,N_1021,N_1836);
nand U8847 (N_8847,N_430,N_1674);
and U8848 (N_8848,N_4307,N_1871);
xor U8849 (N_8849,N_3352,N_2395);
nand U8850 (N_8850,N_2331,N_2499);
nor U8851 (N_8851,N_3286,N_866);
nor U8852 (N_8852,N_4499,N_4289);
or U8853 (N_8853,N_1033,N_3936);
or U8854 (N_8854,N_2289,N_4519);
and U8855 (N_8855,N_3501,N_636);
nor U8856 (N_8856,N_1646,N_3547);
or U8857 (N_8857,N_292,N_3473);
and U8858 (N_8858,N_1695,N_652);
nand U8859 (N_8859,N_2736,N_844);
and U8860 (N_8860,N_3739,N_2702);
and U8861 (N_8861,N_482,N_1176);
nand U8862 (N_8862,N_1630,N_2006);
or U8863 (N_8863,N_244,N_4405);
and U8864 (N_8864,N_3445,N_4814);
or U8865 (N_8865,N_275,N_4168);
nand U8866 (N_8866,N_1678,N_913);
or U8867 (N_8867,N_3705,N_1453);
and U8868 (N_8868,N_3688,N_282);
and U8869 (N_8869,N_1617,N_4126);
nand U8870 (N_8870,N_3956,N_2369);
nand U8871 (N_8871,N_2662,N_3993);
nor U8872 (N_8872,N_3891,N_4555);
nand U8873 (N_8873,N_3559,N_2514);
nand U8874 (N_8874,N_618,N_127);
or U8875 (N_8875,N_3623,N_318);
nor U8876 (N_8876,N_1025,N_1252);
nor U8877 (N_8877,N_1331,N_1518);
xor U8878 (N_8878,N_810,N_4368);
nor U8879 (N_8879,N_651,N_4796);
or U8880 (N_8880,N_4119,N_4787);
nor U8881 (N_8881,N_516,N_1162);
and U8882 (N_8882,N_0,N_1278);
and U8883 (N_8883,N_3512,N_769);
and U8884 (N_8884,N_1467,N_1326);
or U8885 (N_8885,N_1004,N_1844);
and U8886 (N_8886,N_2980,N_513);
nand U8887 (N_8887,N_1673,N_441);
nand U8888 (N_8888,N_3744,N_3609);
nor U8889 (N_8889,N_4725,N_970);
or U8890 (N_8890,N_3290,N_2633);
nand U8891 (N_8891,N_973,N_197);
nand U8892 (N_8892,N_2260,N_4303);
nand U8893 (N_8893,N_681,N_4132);
and U8894 (N_8894,N_3694,N_436);
nand U8895 (N_8895,N_3641,N_2802);
nand U8896 (N_8896,N_4457,N_2393);
nand U8897 (N_8897,N_3061,N_2553);
and U8898 (N_8898,N_2314,N_3053);
nand U8899 (N_8899,N_410,N_2669);
xor U8900 (N_8900,N_3968,N_3678);
nand U8901 (N_8901,N_3009,N_3083);
nor U8902 (N_8902,N_3094,N_4439);
nor U8903 (N_8903,N_3882,N_3385);
and U8904 (N_8904,N_1048,N_3718);
nand U8905 (N_8905,N_2235,N_3799);
nor U8906 (N_8906,N_3327,N_4385);
nand U8907 (N_8907,N_383,N_2012);
nand U8908 (N_8908,N_2069,N_2725);
or U8909 (N_8909,N_4931,N_1381);
nor U8910 (N_8910,N_1773,N_2800);
nand U8911 (N_8911,N_4982,N_2245);
nand U8912 (N_8912,N_3259,N_3734);
nor U8913 (N_8913,N_2140,N_2250);
or U8914 (N_8914,N_3839,N_4088);
or U8915 (N_8915,N_67,N_1208);
nor U8916 (N_8916,N_1115,N_2144);
or U8917 (N_8917,N_1189,N_134);
nor U8918 (N_8918,N_3849,N_3900);
and U8919 (N_8919,N_1291,N_1256);
and U8920 (N_8920,N_1341,N_3535);
nor U8921 (N_8921,N_492,N_3353);
nand U8922 (N_8922,N_4278,N_352);
and U8923 (N_8923,N_4100,N_248);
nand U8924 (N_8924,N_4831,N_1103);
and U8925 (N_8925,N_2243,N_799);
nor U8926 (N_8926,N_1011,N_206);
nor U8927 (N_8927,N_1589,N_3544);
and U8928 (N_8928,N_630,N_4002);
or U8929 (N_8929,N_4241,N_4579);
nor U8930 (N_8930,N_4946,N_2180);
nand U8931 (N_8931,N_4601,N_3433);
or U8932 (N_8932,N_2766,N_2760);
and U8933 (N_8933,N_1217,N_1102);
or U8934 (N_8934,N_4544,N_2117);
nor U8935 (N_8935,N_2026,N_2647);
or U8936 (N_8936,N_2583,N_1302);
or U8937 (N_8937,N_4980,N_3869);
nand U8938 (N_8938,N_2197,N_2973);
and U8939 (N_8939,N_3704,N_491);
or U8940 (N_8940,N_679,N_4262);
nor U8941 (N_8941,N_4047,N_2022);
nand U8942 (N_8942,N_917,N_2892);
or U8943 (N_8943,N_4248,N_1676);
nand U8944 (N_8944,N_4296,N_2669);
nand U8945 (N_8945,N_2553,N_329);
nand U8946 (N_8946,N_148,N_4210);
or U8947 (N_8947,N_979,N_203);
and U8948 (N_8948,N_4691,N_4278);
nor U8949 (N_8949,N_1837,N_3117);
nand U8950 (N_8950,N_1662,N_2253);
and U8951 (N_8951,N_4090,N_914);
nand U8952 (N_8952,N_3548,N_709);
and U8953 (N_8953,N_4031,N_2685);
nand U8954 (N_8954,N_4086,N_4581);
or U8955 (N_8955,N_4871,N_815);
and U8956 (N_8956,N_4709,N_1623);
and U8957 (N_8957,N_331,N_2709);
nand U8958 (N_8958,N_4509,N_476);
and U8959 (N_8959,N_3693,N_786);
nand U8960 (N_8960,N_3051,N_1925);
nand U8961 (N_8961,N_4788,N_1003);
or U8962 (N_8962,N_3773,N_1517);
or U8963 (N_8963,N_1105,N_427);
nor U8964 (N_8964,N_2169,N_1303);
nand U8965 (N_8965,N_2127,N_587);
or U8966 (N_8966,N_3689,N_3482);
and U8967 (N_8967,N_1935,N_3679);
or U8968 (N_8968,N_621,N_1717);
nor U8969 (N_8969,N_3756,N_998);
nor U8970 (N_8970,N_4967,N_1445);
nor U8971 (N_8971,N_4544,N_345);
and U8972 (N_8972,N_4690,N_3641);
nor U8973 (N_8973,N_4556,N_3086);
nor U8974 (N_8974,N_2808,N_3498);
nor U8975 (N_8975,N_3709,N_2533);
and U8976 (N_8976,N_3727,N_218);
nor U8977 (N_8977,N_3878,N_2251);
nand U8978 (N_8978,N_427,N_2004);
and U8979 (N_8979,N_4301,N_1800);
or U8980 (N_8980,N_1259,N_3733);
nor U8981 (N_8981,N_356,N_873);
and U8982 (N_8982,N_3632,N_888);
nor U8983 (N_8983,N_4703,N_4879);
nor U8984 (N_8984,N_626,N_1227);
nor U8985 (N_8985,N_1143,N_208);
nor U8986 (N_8986,N_3663,N_810);
or U8987 (N_8987,N_2650,N_2046);
and U8988 (N_8988,N_2400,N_2414);
nor U8989 (N_8989,N_808,N_4518);
nor U8990 (N_8990,N_4123,N_4311);
nor U8991 (N_8991,N_3495,N_2073);
and U8992 (N_8992,N_606,N_2869);
nor U8993 (N_8993,N_4068,N_329);
nor U8994 (N_8994,N_2841,N_759);
and U8995 (N_8995,N_4128,N_2810);
nand U8996 (N_8996,N_1226,N_4675);
and U8997 (N_8997,N_896,N_2795);
nor U8998 (N_8998,N_4963,N_3754);
and U8999 (N_8999,N_2485,N_343);
nand U9000 (N_9000,N_3630,N_2768);
and U9001 (N_9001,N_4293,N_1854);
and U9002 (N_9002,N_4860,N_2338);
and U9003 (N_9003,N_1534,N_1497);
nor U9004 (N_9004,N_1969,N_1509);
nor U9005 (N_9005,N_4841,N_3999);
or U9006 (N_9006,N_4851,N_890);
and U9007 (N_9007,N_651,N_1223);
or U9008 (N_9008,N_2565,N_2212);
nor U9009 (N_9009,N_4861,N_628);
and U9010 (N_9010,N_4025,N_4778);
or U9011 (N_9011,N_167,N_1704);
or U9012 (N_9012,N_3096,N_426);
nor U9013 (N_9013,N_3609,N_2832);
or U9014 (N_9014,N_2927,N_47);
nor U9015 (N_9015,N_4951,N_1261);
and U9016 (N_9016,N_3401,N_2445);
nor U9017 (N_9017,N_4002,N_2993);
nand U9018 (N_9018,N_1832,N_4308);
nor U9019 (N_9019,N_2387,N_2847);
and U9020 (N_9020,N_4968,N_1363);
and U9021 (N_9021,N_1634,N_1917);
or U9022 (N_9022,N_4045,N_3698);
nor U9023 (N_9023,N_809,N_2938);
or U9024 (N_9024,N_2669,N_830);
nand U9025 (N_9025,N_3525,N_1344);
nand U9026 (N_9026,N_2745,N_4341);
nand U9027 (N_9027,N_1425,N_1977);
nand U9028 (N_9028,N_2940,N_1597);
or U9029 (N_9029,N_652,N_1010);
nor U9030 (N_9030,N_1709,N_1472);
and U9031 (N_9031,N_305,N_4121);
nand U9032 (N_9032,N_3988,N_1019);
nand U9033 (N_9033,N_575,N_4362);
nor U9034 (N_9034,N_3439,N_3421);
and U9035 (N_9035,N_2640,N_2077);
nor U9036 (N_9036,N_1810,N_4034);
and U9037 (N_9037,N_801,N_1028);
nor U9038 (N_9038,N_2560,N_3950);
nand U9039 (N_9039,N_4926,N_1436);
nand U9040 (N_9040,N_84,N_4623);
nand U9041 (N_9041,N_1454,N_3683);
and U9042 (N_9042,N_4412,N_4023);
or U9043 (N_9043,N_4624,N_1254);
and U9044 (N_9044,N_915,N_3521);
nand U9045 (N_9045,N_829,N_4686);
nor U9046 (N_9046,N_2840,N_2325);
nand U9047 (N_9047,N_4258,N_4539);
or U9048 (N_9048,N_4613,N_804);
and U9049 (N_9049,N_927,N_1606);
nand U9050 (N_9050,N_805,N_3188);
nor U9051 (N_9051,N_4247,N_1192);
and U9052 (N_9052,N_1813,N_1126);
or U9053 (N_9053,N_167,N_914);
or U9054 (N_9054,N_1717,N_4035);
nor U9055 (N_9055,N_3210,N_732);
nand U9056 (N_9056,N_3332,N_3239);
and U9057 (N_9057,N_2883,N_3697);
nor U9058 (N_9058,N_3605,N_1017);
or U9059 (N_9059,N_3841,N_314);
nand U9060 (N_9060,N_1585,N_4878);
nand U9061 (N_9061,N_3004,N_4950);
or U9062 (N_9062,N_4435,N_418);
and U9063 (N_9063,N_2825,N_2202);
or U9064 (N_9064,N_178,N_21);
nor U9065 (N_9065,N_3668,N_2117);
and U9066 (N_9066,N_2898,N_3992);
or U9067 (N_9067,N_3364,N_3089);
nand U9068 (N_9068,N_4260,N_3306);
or U9069 (N_9069,N_388,N_1226);
or U9070 (N_9070,N_4387,N_1166);
nor U9071 (N_9071,N_4220,N_1709);
nor U9072 (N_9072,N_3424,N_3895);
and U9073 (N_9073,N_4713,N_4917);
xor U9074 (N_9074,N_4385,N_1981);
or U9075 (N_9075,N_1049,N_4830);
nor U9076 (N_9076,N_2040,N_1916);
or U9077 (N_9077,N_1955,N_233);
nor U9078 (N_9078,N_318,N_4943);
nand U9079 (N_9079,N_3158,N_768);
nor U9080 (N_9080,N_4869,N_2673);
and U9081 (N_9081,N_3903,N_97);
xnor U9082 (N_9082,N_3566,N_1287);
or U9083 (N_9083,N_491,N_289);
nor U9084 (N_9084,N_4581,N_1106);
and U9085 (N_9085,N_42,N_2800);
or U9086 (N_9086,N_3946,N_4969);
nand U9087 (N_9087,N_1485,N_1978);
nand U9088 (N_9088,N_656,N_1529);
nand U9089 (N_9089,N_3810,N_574);
or U9090 (N_9090,N_2371,N_4125);
xor U9091 (N_9091,N_168,N_4157);
or U9092 (N_9092,N_490,N_2215);
nand U9093 (N_9093,N_798,N_1584);
or U9094 (N_9094,N_4583,N_4407);
and U9095 (N_9095,N_3467,N_233);
and U9096 (N_9096,N_2853,N_233);
nor U9097 (N_9097,N_3058,N_3602);
nand U9098 (N_9098,N_1624,N_4431);
nand U9099 (N_9099,N_4059,N_1188);
nand U9100 (N_9100,N_939,N_71);
or U9101 (N_9101,N_2723,N_1198);
and U9102 (N_9102,N_4662,N_4562);
nand U9103 (N_9103,N_2397,N_3991);
and U9104 (N_9104,N_690,N_3377);
nor U9105 (N_9105,N_4485,N_2021);
and U9106 (N_9106,N_1148,N_1409);
nor U9107 (N_9107,N_4446,N_1255);
nand U9108 (N_9108,N_301,N_1174);
nor U9109 (N_9109,N_2227,N_808);
nand U9110 (N_9110,N_1135,N_4428);
nor U9111 (N_9111,N_32,N_4131);
and U9112 (N_9112,N_3101,N_2324);
and U9113 (N_9113,N_1328,N_2978);
nor U9114 (N_9114,N_3058,N_1583);
nand U9115 (N_9115,N_3869,N_867);
and U9116 (N_9116,N_3143,N_1801);
nand U9117 (N_9117,N_2299,N_556);
nand U9118 (N_9118,N_1975,N_4053);
nand U9119 (N_9119,N_2688,N_3696);
nand U9120 (N_9120,N_231,N_4369);
or U9121 (N_9121,N_3143,N_2139);
and U9122 (N_9122,N_3657,N_2938);
nand U9123 (N_9123,N_2228,N_1161);
or U9124 (N_9124,N_1211,N_2797);
and U9125 (N_9125,N_1451,N_2800);
or U9126 (N_9126,N_393,N_409);
and U9127 (N_9127,N_1770,N_156);
and U9128 (N_9128,N_146,N_1257);
and U9129 (N_9129,N_388,N_403);
nor U9130 (N_9130,N_2213,N_3184);
nand U9131 (N_9131,N_771,N_173);
or U9132 (N_9132,N_2393,N_1568);
nor U9133 (N_9133,N_4844,N_4979);
and U9134 (N_9134,N_2300,N_1615);
nor U9135 (N_9135,N_3235,N_420);
or U9136 (N_9136,N_3387,N_1010);
nor U9137 (N_9137,N_2723,N_3073);
and U9138 (N_9138,N_4412,N_4602);
and U9139 (N_9139,N_3641,N_1666);
or U9140 (N_9140,N_3845,N_1298);
or U9141 (N_9141,N_3108,N_36);
xnor U9142 (N_9142,N_1597,N_301);
nand U9143 (N_9143,N_940,N_1239);
nor U9144 (N_9144,N_4873,N_4281);
or U9145 (N_9145,N_2068,N_3689);
and U9146 (N_9146,N_3996,N_2308);
nor U9147 (N_9147,N_1237,N_4291);
nand U9148 (N_9148,N_4333,N_3412);
nand U9149 (N_9149,N_4010,N_2790);
and U9150 (N_9150,N_2304,N_4555);
nand U9151 (N_9151,N_4722,N_2980);
and U9152 (N_9152,N_3875,N_2538);
xor U9153 (N_9153,N_740,N_4628);
nand U9154 (N_9154,N_4349,N_4097);
or U9155 (N_9155,N_48,N_195);
and U9156 (N_9156,N_3413,N_1997);
nand U9157 (N_9157,N_1434,N_3068);
nor U9158 (N_9158,N_2414,N_2360);
or U9159 (N_9159,N_2167,N_3229);
or U9160 (N_9160,N_3533,N_1250);
nor U9161 (N_9161,N_1513,N_2281);
nor U9162 (N_9162,N_1980,N_4017);
nor U9163 (N_9163,N_3230,N_2196);
nand U9164 (N_9164,N_1918,N_290);
or U9165 (N_9165,N_2033,N_1455);
nor U9166 (N_9166,N_2818,N_2971);
and U9167 (N_9167,N_3301,N_2154);
nand U9168 (N_9168,N_1393,N_2070);
nand U9169 (N_9169,N_734,N_2672);
or U9170 (N_9170,N_2677,N_406);
nand U9171 (N_9171,N_3479,N_3456);
or U9172 (N_9172,N_4769,N_4156);
or U9173 (N_9173,N_1345,N_2612);
or U9174 (N_9174,N_4072,N_3521);
and U9175 (N_9175,N_4368,N_1196);
nor U9176 (N_9176,N_3772,N_3444);
xor U9177 (N_9177,N_964,N_4551);
nand U9178 (N_9178,N_2281,N_4473);
nor U9179 (N_9179,N_2799,N_36);
nor U9180 (N_9180,N_1600,N_3470);
or U9181 (N_9181,N_3932,N_138);
and U9182 (N_9182,N_4029,N_3598);
or U9183 (N_9183,N_4693,N_3562);
nand U9184 (N_9184,N_579,N_3079);
and U9185 (N_9185,N_4237,N_74);
or U9186 (N_9186,N_5,N_3029);
and U9187 (N_9187,N_1918,N_4743);
and U9188 (N_9188,N_2474,N_4833);
or U9189 (N_9189,N_662,N_3111);
or U9190 (N_9190,N_4578,N_4101);
nand U9191 (N_9191,N_3456,N_1394);
and U9192 (N_9192,N_3003,N_2340);
and U9193 (N_9193,N_3210,N_1193);
nor U9194 (N_9194,N_4767,N_895);
and U9195 (N_9195,N_3685,N_3473);
and U9196 (N_9196,N_1885,N_2697);
or U9197 (N_9197,N_2743,N_434);
and U9198 (N_9198,N_4755,N_4919);
or U9199 (N_9199,N_2495,N_2152);
or U9200 (N_9200,N_2045,N_1802);
nand U9201 (N_9201,N_2336,N_1027);
or U9202 (N_9202,N_4683,N_4451);
nand U9203 (N_9203,N_2756,N_1784);
nand U9204 (N_9204,N_587,N_4505);
nand U9205 (N_9205,N_4179,N_1191);
or U9206 (N_9206,N_2011,N_2537);
nor U9207 (N_9207,N_4375,N_2273);
nor U9208 (N_9208,N_751,N_4389);
and U9209 (N_9209,N_4441,N_4291);
nand U9210 (N_9210,N_2813,N_4411);
nor U9211 (N_9211,N_811,N_3841);
or U9212 (N_9212,N_4571,N_2029);
or U9213 (N_9213,N_1618,N_2686);
and U9214 (N_9214,N_1870,N_3678);
and U9215 (N_9215,N_3994,N_1788);
nand U9216 (N_9216,N_1507,N_1252);
nand U9217 (N_9217,N_1417,N_3749);
or U9218 (N_9218,N_1947,N_4620);
nand U9219 (N_9219,N_112,N_1687);
xnor U9220 (N_9220,N_2214,N_653);
nand U9221 (N_9221,N_3841,N_4465);
or U9222 (N_9222,N_930,N_524);
and U9223 (N_9223,N_2106,N_1362);
or U9224 (N_9224,N_231,N_4934);
and U9225 (N_9225,N_2850,N_2656);
and U9226 (N_9226,N_2460,N_1767);
or U9227 (N_9227,N_3675,N_734);
nor U9228 (N_9228,N_3958,N_3919);
nor U9229 (N_9229,N_1768,N_4501);
or U9230 (N_9230,N_1924,N_1064);
nor U9231 (N_9231,N_4807,N_352);
nand U9232 (N_9232,N_673,N_3017);
or U9233 (N_9233,N_3096,N_3773);
nand U9234 (N_9234,N_3176,N_4406);
nand U9235 (N_9235,N_2471,N_667);
and U9236 (N_9236,N_211,N_1733);
nand U9237 (N_9237,N_616,N_3405);
and U9238 (N_9238,N_4067,N_41);
nand U9239 (N_9239,N_2788,N_3997);
nor U9240 (N_9240,N_1497,N_4681);
or U9241 (N_9241,N_1648,N_3800);
nor U9242 (N_9242,N_3867,N_781);
nand U9243 (N_9243,N_2434,N_869);
or U9244 (N_9244,N_3520,N_3526);
nand U9245 (N_9245,N_3125,N_69);
or U9246 (N_9246,N_1434,N_1570);
or U9247 (N_9247,N_4950,N_1796);
nand U9248 (N_9248,N_556,N_501);
and U9249 (N_9249,N_1522,N_4997);
and U9250 (N_9250,N_3566,N_80);
nor U9251 (N_9251,N_1250,N_3813);
and U9252 (N_9252,N_4933,N_2040);
xnor U9253 (N_9253,N_243,N_879);
and U9254 (N_9254,N_4604,N_560);
nand U9255 (N_9255,N_2328,N_2890);
nand U9256 (N_9256,N_1319,N_1324);
nor U9257 (N_9257,N_3506,N_4673);
nand U9258 (N_9258,N_1387,N_950);
or U9259 (N_9259,N_3768,N_1036);
xor U9260 (N_9260,N_1390,N_4197);
nor U9261 (N_9261,N_3477,N_4554);
nand U9262 (N_9262,N_4219,N_3991);
and U9263 (N_9263,N_4060,N_643);
and U9264 (N_9264,N_2501,N_1389);
nand U9265 (N_9265,N_3320,N_572);
nand U9266 (N_9266,N_4359,N_1882);
nor U9267 (N_9267,N_3239,N_4612);
or U9268 (N_9268,N_3247,N_1162);
and U9269 (N_9269,N_1726,N_3645);
nor U9270 (N_9270,N_3065,N_2521);
xor U9271 (N_9271,N_2301,N_4628);
and U9272 (N_9272,N_2186,N_3733);
or U9273 (N_9273,N_4562,N_4286);
nand U9274 (N_9274,N_4490,N_4924);
or U9275 (N_9275,N_1436,N_1305);
nor U9276 (N_9276,N_4585,N_3228);
nor U9277 (N_9277,N_3953,N_4524);
and U9278 (N_9278,N_3112,N_143);
nor U9279 (N_9279,N_904,N_455);
or U9280 (N_9280,N_4630,N_2631);
nand U9281 (N_9281,N_4103,N_3794);
and U9282 (N_9282,N_2156,N_4366);
or U9283 (N_9283,N_4649,N_4334);
and U9284 (N_9284,N_126,N_1795);
or U9285 (N_9285,N_1694,N_2097);
nor U9286 (N_9286,N_664,N_2850);
and U9287 (N_9287,N_4780,N_4696);
or U9288 (N_9288,N_1319,N_3893);
nand U9289 (N_9289,N_1,N_191);
and U9290 (N_9290,N_2598,N_2933);
nand U9291 (N_9291,N_4052,N_2680);
or U9292 (N_9292,N_3659,N_1110);
nor U9293 (N_9293,N_2385,N_390);
or U9294 (N_9294,N_2018,N_577);
nor U9295 (N_9295,N_3437,N_1902);
and U9296 (N_9296,N_3468,N_4017);
nand U9297 (N_9297,N_4332,N_3177);
or U9298 (N_9298,N_3261,N_3046);
and U9299 (N_9299,N_498,N_599);
or U9300 (N_9300,N_3813,N_1217);
or U9301 (N_9301,N_4293,N_2010);
nor U9302 (N_9302,N_884,N_1576);
and U9303 (N_9303,N_2164,N_1740);
nand U9304 (N_9304,N_4874,N_695);
and U9305 (N_9305,N_2359,N_2311);
and U9306 (N_9306,N_4662,N_2302);
nor U9307 (N_9307,N_2817,N_3371);
or U9308 (N_9308,N_4936,N_291);
nand U9309 (N_9309,N_3637,N_4885);
and U9310 (N_9310,N_35,N_3086);
nand U9311 (N_9311,N_4235,N_3994);
nor U9312 (N_9312,N_350,N_3047);
or U9313 (N_9313,N_883,N_4142);
nor U9314 (N_9314,N_4763,N_3068);
or U9315 (N_9315,N_2903,N_2101);
and U9316 (N_9316,N_46,N_2902);
or U9317 (N_9317,N_1048,N_1510);
or U9318 (N_9318,N_806,N_1532);
and U9319 (N_9319,N_2453,N_124);
and U9320 (N_9320,N_4656,N_4151);
and U9321 (N_9321,N_1698,N_3635);
nand U9322 (N_9322,N_2097,N_3351);
nor U9323 (N_9323,N_2155,N_4032);
and U9324 (N_9324,N_3928,N_1953);
nor U9325 (N_9325,N_1980,N_1460);
or U9326 (N_9326,N_3305,N_3468);
nor U9327 (N_9327,N_4837,N_3034);
nand U9328 (N_9328,N_2996,N_2601);
and U9329 (N_9329,N_3743,N_1659);
or U9330 (N_9330,N_4070,N_1310);
and U9331 (N_9331,N_3698,N_4648);
nor U9332 (N_9332,N_2389,N_1620);
and U9333 (N_9333,N_4763,N_193);
and U9334 (N_9334,N_1156,N_4349);
nand U9335 (N_9335,N_4715,N_1123);
and U9336 (N_9336,N_2622,N_1947);
and U9337 (N_9337,N_3295,N_2190);
nor U9338 (N_9338,N_4079,N_3359);
nand U9339 (N_9339,N_517,N_4845);
or U9340 (N_9340,N_4756,N_3951);
nor U9341 (N_9341,N_3346,N_1788);
and U9342 (N_9342,N_4332,N_2119);
or U9343 (N_9343,N_1993,N_4473);
nand U9344 (N_9344,N_2565,N_1950);
or U9345 (N_9345,N_2755,N_4709);
or U9346 (N_9346,N_3880,N_4833);
nor U9347 (N_9347,N_4245,N_22);
and U9348 (N_9348,N_2260,N_4593);
nor U9349 (N_9349,N_190,N_3514);
nor U9350 (N_9350,N_3383,N_1557);
and U9351 (N_9351,N_3324,N_4448);
and U9352 (N_9352,N_1491,N_2653);
nand U9353 (N_9353,N_4820,N_1586);
or U9354 (N_9354,N_1099,N_3188);
or U9355 (N_9355,N_3639,N_2746);
nand U9356 (N_9356,N_2067,N_1075);
nand U9357 (N_9357,N_2237,N_4887);
nor U9358 (N_9358,N_4619,N_1154);
nor U9359 (N_9359,N_631,N_1914);
nor U9360 (N_9360,N_4939,N_975);
nand U9361 (N_9361,N_4855,N_2864);
or U9362 (N_9362,N_507,N_3986);
and U9363 (N_9363,N_4353,N_4372);
nand U9364 (N_9364,N_4655,N_686);
xnor U9365 (N_9365,N_102,N_4407);
nor U9366 (N_9366,N_2731,N_239);
nor U9367 (N_9367,N_459,N_3823);
nor U9368 (N_9368,N_4907,N_3391);
or U9369 (N_9369,N_3006,N_4117);
nor U9370 (N_9370,N_4593,N_1063);
or U9371 (N_9371,N_2904,N_892);
nor U9372 (N_9372,N_2211,N_975);
nor U9373 (N_9373,N_4414,N_1277);
and U9374 (N_9374,N_2869,N_4340);
and U9375 (N_9375,N_1192,N_2545);
and U9376 (N_9376,N_2000,N_2485);
and U9377 (N_9377,N_4946,N_4196);
nand U9378 (N_9378,N_4448,N_1962);
or U9379 (N_9379,N_1966,N_3274);
and U9380 (N_9380,N_2721,N_3645);
nor U9381 (N_9381,N_2341,N_1534);
and U9382 (N_9382,N_4160,N_159);
and U9383 (N_9383,N_2617,N_3090);
or U9384 (N_9384,N_1104,N_4870);
and U9385 (N_9385,N_4987,N_4943);
or U9386 (N_9386,N_976,N_1682);
and U9387 (N_9387,N_4716,N_4218);
or U9388 (N_9388,N_4800,N_1042);
or U9389 (N_9389,N_396,N_1169);
nor U9390 (N_9390,N_350,N_1139);
nor U9391 (N_9391,N_4203,N_4006);
nor U9392 (N_9392,N_1732,N_4018);
and U9393 (N_9393,N_3572,N_4424);
nand U9394 (N_9394,N_1531,N_4844);
nand U9395 (N_9395,N_988,N_3860);
nand U9396 (N_9396,N_3180,N_810);
nand U9397 (N_9397,N_1739,N_319);
nand U9398 (N_9398,N_312,N_4430);
and U9399 (N_9399,N_4029,N_3134);
nand U9400 (N_9400,N_3834,N_665);
and U9401 (N_9401,N_680,N_1395);
nand U9402 (N_9402,N_4113,N_2769);
and U9403 (N_9403,N_3877,N_3661);
and U9404 (N_9404,N_2981,N_1345);
nand U9405 (N_9405,N_841,N_3184);
nor U9406 (N_9406,N_657,N_4607);
nor U9407 (N_9407,N_2551,N_2943);
and U9408 (N_9408,N_2306,N_3038);
nand U9409 (N_9409,N_4285,N_3185);
and U9410 (N_9410,N_1620,N_383);
or U9411 (N_9411,N_4716,N_1119);
and U9412 (N_9412,N_3567,N_2696);
nor U9413 (N_9413,N_3532,N_3398);
and U9414 (N_9414,N_4733,N_4177);
nor U9415 (N_9415,N_1714,N_1622);
nor U9416 (N_9416,N_3577,N_3027);
nor U9417 (N_9417,N_1286,N_1172);
nand U9418 (N_9418,N_2302,N_2463);
and U9419 (N_9419,N_2257,N_1430);
or U9420 (N_9420,N_3190,N_2137);
nand U9421 (N_9421,N_919,N_1077);
and U9422 (N_9422,N_1149,N_4094);
nand U9423 (N_9423,N_503,N_609);
and U9424 (N_9424,N_2169,N_2179);
or U9425 (N_9425,N_1967,N_2539);
nor U9426 (N_9426,N_1419,N_3530);
and U9427 (N_9427,N_2315,N_2221);
or U9428 (N_9428,N_1245,N_2674);
nand U9429 (N_9429,N_1299,N_724);
nand U9430 (N_9430,N_1611,N_965);
and U9431 (N_9431,N_1913,N_215);
nand U9432 (N_9432,N_3501,N_1509);
and U9433 (N_9433,N_219,N_2075);
nor U9434 (N_9434,N_2781,N_795);
and U9435 (N_9435,N_1447,N_4478);
or U9436 (N_9436,N_1745,N_2985);
nor U9437 (N_9437,N_3056,N_737);
xor U9438 (N_9438,N_810,N_494);
nor U9439 (N_9439,N_3379,N_2832);
nand U9440 (N_9440,N_2979,N_3747);
nor U9441 (N_9441,N_1478,N_4913);
nor U9442 (N_9442,N_152,N_2091);
or U9443 (N_9443,N_1684,N_2585);
nor U9444 (N_9444,N_2213,N_3073);
and U9445 (N_9445,N_3914,N_4261);
or U9446 (N_9446,N_618,N_4189);
and U9447 (N_9447,N_3328,N_3723);
nor U9448 (N_9448,N_2615,N_2312);
nor U9449 (N_9449,N_1974,N_4198);
or U9450 (N_9450,N_4790,N_3212);
and U9451 (N_9451,N_4062,N_496);
nor U9452 (N_9452,N_1426,N_2979);
or U9453 (N_9453,N_4134,N_103);
nor U9454 (N_9454,N_4238,N_2189);
and U9455 (N_9455,N_172,N_2311);
nand U9456 (N_9456,N_3175,N_4717);
or U9457 (N_9457,N_1276,N_2858);
and U9458 (N_9458,N_3987,N_2253);
and U9459 (N_9459,N_1671,N_4487);
and U9460 (N_9460,N_851,N_3579);
nor U9461 (N_9461,N_4354,N_338);
or U9462 (N_9462,N_3254,N_2825);
nand U9463 (N_9463,N_1131,N_1171);
nand U9464 (N_9464,N_4633,N_4425);
nor U9465 (N_9465,N_3299,N_2765);
or U9466 (N_9466,N_3079,N_866);
and U9467 (N_9467,N_3152,N_2460);
or U9468 (N_9468,N_25,N_4522);
nor U9469 (N_9469,N_3010,N_2490);
or U9470 (N_9470,N_862,N_1706);
or U9471 (N_9471,N_1848,N_487);
or U9472 (N_9472,N_1890,N_4525);
or U9473 (N_9473,N_4766,N_1804);
and U9474 (N_9474,N_3802,N_791);
or U9475 (N_9475,N_3774,N_4376);
nand U9476 (N_9476,N_2866,N_1360);
and U9477 (N_9477,N_2857,N_4517);
nor U9478 (N_9478,N_4722,N_419);
nor U9479 (N_9479,N_2971,N_3363);
nand U9480 (N_9480,N_3240,N_1792);
or U9481 (N_9481,N_1667,N_1916);
nor U9482 (N_9482,N_1300,N_4653);
nand U9483 (N_9483,N_4594,N_3000);
nor U9484 (N_9484,N_4352,N_845);
nand U9485 (N_9485,N_592,N_2328);
or U9486 (N_9486,N_1210,N_3526);
and U9487 (N_9487,N_3940,N_4000);
or U9488 (N_9488,N_3935,N_4952);
nor U9489 (N_9489,N_2583,N_14);
and U9490 (N_9490,N_852,N_4605);
nand U9491 (N_9491,N_1613,N_2743);
nand U9492 (N_9492,N_938,N_1628);
nor U9493 (N_9493,N_4640,N_1874);
nand U9494 (N_9494,N_2613,N_2570);
or U9495 (N_9495,N_999,N_1902);
or U9496 (N_9496,N_3136,N_495);
nor U9497 (N_9497,N_4764,N_145);
and U9498 (N_9498,N_1752,N_4290);
or U9499 (N_9499,N_2908,N_579);
nor U9500 (N_9500,N_4667,N_1192);
or U9501 (N_9501,N_4336,N_1320);
nand U9502 (N_9502,N_238,N_2297);
nor U9503 (N_9503,N_1686,N_4005);
or U9504 (N_9504,N_3539,N_1316);
nand U9505 (N_9505,N_1744,N_2064);
nor U9506 (N_9506,N_629,N_4636);
nand U9507 (N_9507,N_3694,N_3750);
nand U9508 (N_9508,N_4198,N_4661);
nor U9509 (N_9509,N_1613,N_2496);
nor U9510 (N_9510,N_544,N_3673);
nor U9511 (N_9511,N_1850,N_1583);
nor U9512 (N_9512,N_4789,N_1426);
nand U9513 (N_9513,N_1631,N_1274);
nor U9514 (N_9514,N_1187,N_2141);
or U9515 (N_9515,N_523,N_3321);
and U9516 (N_9516,N_4712,N_989);
and U9517 (N_9517,N_1008,N_1269);
or U9518 (N_9518,N_2593,N_651);
nand U9519 (N_9519,N_2562,N_295);
nor U9520 (N_9520,N_4579,N_294);
nand U9521 (N_9521,N_921,N_695);
or U9522 (N_9522,N_579,N_666);
and U9523 (N_9523,N_4745,N_3341);
nand U9524 (N_9524,N_2373,N_1337);
nand U9525 (N_9525,N_1076,N_1910);
or U9526 (N_9526,N_1208,N_1960);
nand U9527 (N_9527,N_247,N_1470);
and U9528 (N_9528,N_2086,N_785);
and U9529 (N_9529,N_4093,N_944);
or U9530 (N_9530,N_3792,N_3519);
and U9531 (N_9531,N_4604,N_4239);
and U9532 (N_9532,N_432,N_3726);
nand U9533 (N_9533,N_4764,N_120);
nor U9534 (N_9534,N_1579,N_4351);
or U9535 (N_9535,N_3536,N_4810);
nor U9536 (N_9536,N_4724,N_2265);
nand U9537 (N_9537,N_3853,N_2395);
nand U9538 (N_9538,N_3967,N_3756);
xor U9539 (N_9539,N_1216,N_1689);
and U9540 (N_9540,N_3156,N_2639);
and U9541 (N_9541,N_1655,N_2609);
and U9542 (N_9542,N_4769,N_1598);
nand U9543 (N_9543,N_2490,N_4796);
nor U9544 (N_9544,N_22,N_4641);
nor U9545 (N_9545,N_98,N_3110);
nor U9546 (N_9546,N_3954,N_1347);
and U9547 (N_9547,N_2923,N_4394);
and U9548 (N_9548,N_34,N_2780);
nand U9549 (N_9549,N_3356,N_2098);
or U9550 (N_9550,N_3797,N_518);
and U9551 (N_9551,N_4271,N_2421);
or U9552 (N_9552,N_4806,N_2653);
nand U9553 (N_9553,N_4659,N_1275);
or U9554 (N_9554,N_2234,N_4588);
nor U9555 (N_9555,N_4890,N_2434);
nor U9556 (N_9556,N_3500,N_750);
nor U9557 (N_9557,N_2811,N_181);
nand U9558 (N_9558,N_1153,N_1781);
nand U9559 (N_9559,N_4760,N_4391);
or U9560 (N_9560,N_4800,N_2717);
nor U9561 (N_9561,N_3383,N_914);
nor U9562 (N_9562,N_3348,N_1281);
and U9563 (N_9563,N_1745,N_3943);
and U9564 (N_9564,N_3865,N_3569);
nor U9565 (N_9565,N_1832,N_2989);
or U9566 (N_9566,N_1260,N_3997);
or U9567 (N_9567,N_4385,N_2735);
nor U9568 (N_9568,N_1550,N_4658);
nor U9569 (N_9569,N_4798,N_131);
and U9570 (N_9570,N_484,N_358);
and U9571 (N_9571,N_1675,N_397);
nor U9572 (N_9572,N_324,N_730);
and U9573 (N_9573,N_766,N_3326);
nand U9574 (N_9574,N_154,N_1401);
or U9575 (N_9575,N_266,N_3426);
nor U9576 (N_9576,N_4423,N_4838);
nand U9577 (N_9577,N_5,N_3553);
nand U9578 (N_9578,N_2127,N_3673);
and U9579 (N_9579,N_1551,N_1263);
and U9580 (N_9580,N_2705,N_1712);
nand U9581 (N_9581,N_1627,N_4567);
or U9582 (N_9582,N_1938,N_531);
nor U9583 (N_9583,N_4970,N_3114);
or U9584 (N_9584,N_537,N_4003);
nor U9585 (N_9585,N_3661,N_130);
nor U9586 (N_9586,N_4180,N_1223);
or U9587 (N_9587,N_4530,N_4586);
nor U9588 (N_9588,N_1126,N_438);
nor U9589 (N_9589,N_4614,N_475);
or U9590 (N_9590,N_413,N_2288);
and U9591 (N_9591,N_4885,N_1514);
nor U9592 (N_9592,N_643,N_4203);
nor U9593 (N_9593,N_1246,N_1022);
nor U9594 (N_9594,N_1703,N_4398);
or U9595 (N_9595,N_216,N_3638);
nor U9596 (N_9596,N_2239,N_2136);
nor U9597 (N_9597,N_4122,N_2473);
or U9598 (N_9598,N_3012,N_2612);
and U9599 (N_9599,N_1938,N_1801);
and U9600 (N_9600,N_4746,N_3150);
or U9601 (N_9601,N_4357,N_1477);
and U9602 (N_9602,N_1412,N_3860);
nand U9603 (N_9603,N_4157,N_568);
and U9604 (N_9604,N_4965,N_3998);
nor U9605 (N_9605,N_4380,N_2311);
and U9606 (N_9606,N_1203,N_164);
nand U9607 (N_9607,N_3675,N_3788);
and U9608 (N_9608,N_1430,N_4059);
nor U9609 (N_9609,N_4904,N_4577);
or U9610 (N_9610,N_4341,N_4541);
or U9611 (N_9611,N_678,N_1631);
xnor U9612 (N_9612,N_590,N_2432);
or U9613 (N_9613,N_2406,N_540);
and U9614 (N_9614,N_842,N_1062);
xnor U9615 (N_9615,N_3178,N_1174);
nand U9616 (N_9616,N_1332,N_854);
and U9617 (N_9617,N_3273,N_4613);
and U9618 (N_9618,N_1688,N_3698);
nand U9619 (N_9619,N_173,N_3437);
or U9620 (N_9620,N_3768,N_514);
nor U9621 (N_9621,N_3084,N_1467);
nand U9622 (N_9622,N_2084,N_2864);
and U9623 (N_9623,N_4677,N_3823);
nand U9624 (N_9624,N_2050,N_2264);
and U9625 (N_9625,N_2180,N_189);
nand U9626 (N_9626,N_4971,N_504);
or U9627 (N_9627,N_889,N_1960);
or U9628 (N_9628,N_2669,N_4266);
nor U9629 (N_9629,N_2371,N_4224);
nand U9630 (N_9630,N_3414,N_2799);
nor U9631 (N_9631,N_4780,N_741);
nor U9632 (N_9632,N_4007,N_2361);
nor U9633 (N_9633,N_1944,N_3039);
and U9634 (N_9634,N_4323,N_3547);
or U9635 (N_9635,N_206,N_4215);
nor U9636 (N_9636,N_439,N_3419);
or U9637 (N_9637,N_3952,N_2354);
nor U9638 (N_9638,N_2756,N_3560);
and U9639 (N_9639,N_2641,N_2708);
nand U9640 (N_9640,N_4857,N_2313);
nand U9641 (N_9641,N_2378,N_990);
or U9642 (N_9642,N_1355,N_487);
and U9643 (N_9643,N_1790,N_426);
nor U9644 (N_9644,N_1008,N_2997);
and U9645 (N_9645,N_8,N_3423);
nand U9646 (N_9646,N_909,N_2842);
and U9647 (N_9647,N_712,N_2109);
nand U9648 (N_9648,N_2393,N_1775);
and U9649 (N_9649,N_3306,N_4259);
nand U9650 (N_9650,N_115,N_1803);
nor U9651 (N_9651,N_4644,N_300);
nor U9652 (N_9652,N_3468,N_3530);
or U9653 (N_9653,N_2185,N_480);
and U9654 (N_9654,N_3193,N_920);
nor U9655 (N_9655,N_760,N_703);
and U9656 (N_9656,N_2114,N_4208);
and U9657 (N_9657,N_1222,N_3962);
or U9658 (N_9658,N_207,N_1472);
xnor U9659 (N_9659,N_3204,N_424);
and U9660 (N_9660,N_328,N_1538);
or U9661 (N_9661,N_168,N_4913);
nand U9662 (N_9662,N_1772,N_1227);
and U9663 (N_9663,N_634,N_1998);
or U9664 (N_9664,N_3474,N_3286);
nand U9665 (N_9665,N_701,N_3440);
and U9666 (N_9666,N_1459,N_1857);
nand U9667 (N_9667,N_4477,N_4029);
nor U9668 (N_9668,N_4160,N_2842);
and U9669 (N_9669,N_4485,N_2487);
or U9670 (N_9670,N_2913,N_1137);
nand U9671 (N_9671,N_789,N_2089);
and U9672 (N_9672,N_3251,N_3787);
nand U9673 (N_9673,N_3825,N_4456);
and U9674 (N_9674,N_2301,N_1241);
or U9675 (N_9675,N_856,N_3293);
nor U9676 (N_9676,N_3792,N_4849);
nand U9677 (N_9677,N_936,N_3092);
or U9678 (N_9678,N_4847,N_1835);
or U9679 (N_9679,N_819,N_401);
and U9680 (N_9680,N_1242,N_3063);
nand U9681 (N_9681,N_342,N_2302);
nand U9682 (N_9682,N_1606,N_285);
nor U9683 (N_9683,N_4698,N_2652);
and U9684 (N_9684,N_1527,N_3766);
and U9685 (N_9685,N_2166,N_4942);
nand U9686 (N_9686,N_1323,N_4884);
or U9687 (N_9687,N_4109,N_4207);
nand U9688 (N_9688,N_1280,N_3479);
nor U9689 (N_9689,N_13,N_1619);
xor U9690 (N_9690,N_4825,N_4495);
nor U9691 (N_9691,N_3778,N_3223);
nand U9692 (N_9692,N_349,N_1262);
nand U9693 (N_9693,N_3506,N_2010);
nor U9694 (N_9694,N_4451,N_1115);
and U9695 (N_9695,N_4382,N_1258);
nand U9696 (N_9696,N_1605,N_2958);
nand U9697 (N_9697,N_2560,N_2963);
nor U9698 (N_9698,N_3497,N_232);
nor U9699 (N_9699,N_4162,N_436);
nor U9700 (N_9700,N_4283,N_2239);
or U9701 (N_9701,N_3743,N_56);
nor U9702 (N_9702,N_3867,N_4581);
or U9703 (N_9703,N_4569,N_209);
and U9704 (N_9704,N_4192,N_1231);
nor U9705 (N_9705,N_177,N_247);
or U9706 (N_9706,N_3641,N_3728);
and U9707 (N_9707,N_1090,N_4369);
nor U9708 (N_9708,N_4342,N_747);
and U9709 (N_9709,N_3348,N_681);
nor U9710 (N_9710,N_4203,N_2076);
and U9711 (N_9711,N_3797,N_4968);
nand U9712 (N_9712,N_2662,N_4747);
nand U9713 (N_9713,N_4606,N_4957);
or U9714 (N_9714,N_3804,N_4645);
nand U9715 (N_9715,N_3177,N_662);
nor U9716 (N_9716,N_4584,N_1849);
or U9717 (N_9717,N_67,N_3229);
nor U9718 (N_9718,N_908,N_3576);
or U9719 (N_9719,N_3286,N_4074);
nor U9720 (N_9720,N_3533,N_4134);
nand U9721 (N_9721,N_926,N_2756);
nand U9722 (N_9722,N_3434,N_454);
and U9723 (N_9723,N_4745,N_2822);
and U9724 (N_9724,N_2263,N_5);
nand U9725 (N_9725,N_525,N_4181);
and U9726 (N_9726,N_323,N_3746);
and U9727 (N_9727,N_3143,N_4666);
nor U9728 (N_9728,N_1923,N_3771);
or U9729 (N_9729,N_4400,N_2961);
nor U9730 (N_9730,N_1635,N_258);
and U9731 (N_9731,N_4982,N_1542);
and U9732 (N_9732,N_4489,N_2658);
or U9733 (N_9733,N_707,N_3395);
nand U9734 (N_9734,N_2305,N_1836);
and U9735 (N_9735,N_2059,N_1278);
or U9736 (N_9736,N_4336,N_196);
or U9737 (N_9737,N_4371,N_70);
or U9738 (N_9738,N_534,N_2811);
nand U9739 (N_9739,N_362,N_3457);
nor U9740 (N_9740,N_2043,N_300);
or U9741 (N_9741,N_1612,N_3430);
nand U9742 (N_9742,N_2198,N_1643);
or U9743 (N_9743,N_1279,N_3025);
and U9744 (N_9744,N_3210,N_478);
or U9745 (N_9745,N_1963,N_4541);
nand U9746 (N_9746,N_4921,N_4180);
or U9747 (N_9747,N_2989,N_3417);
nand U9748 (N_9748,N_144,N_1279);
nor U9749 (N_9749,N_4620,N_2690);
and U9750 (N_9750,N_1244,N_457);
nor U9751 (N_9751,N_4138,N_2663);
nand U9752 (N_9752,N_2829,N_4869);
or U9753 (N_9753,N_4355,N_492);
or U9754 (N_9754,N_728,N_3192);
and U9755 (N_9755,N_3974,N_646);
nor U9756 (N_9756,N_3099,N_2246);
nor U9757 (N_9757,N_2451,N_3449);
nand U9758 (N_9758,N_4808,N_1553);
or U9759 (N_9759,N_1618,N_2022);
and U9760 (N_9760,N_4870,N_3292);
or U9761 (N_9761,N_2626,N_562);
nor U9762 (N_9762,N_2546,N_4033);
nand U9763 (N_9763,N_3622,N_4622);
nor U9764 (N_9764,N_2646,N_49);
or U9765 (N_9765,N_4607,N_418);
nor U9766 (N_9766,N_1719,N_1218);
nor U9767 (N_9767,N_3792,N_1914);
nor U9768 (N_9768,N_738,N_351);
and U9769 (N_9769,N_2857,N_4899);
nand U9770 (N_9770,N_1539,N_3487);
nand U9771 (N_9771,N_3035,N_1762);
nor U9772 (N_9772,N_2632,N_1450);
or U9773 (N_9773,N_3176,N_1830);
nand U9774 (N_9774,N_1313,N_2405);
or U9775 (N_9775,N_445,N_3442);
nand U9776 (N_9776,N_234,N_1335);
nand U9777 (N_9777,N_4975,N_2943);
or U9778 (N_9778,N_4108,N_4241);
xnor U9779 (N_9779,N_3074,N_1704);
and U9780 (N_9780,N_379,N_4882);
nand U9781 (N_9781,N_2131,N_2366);
nand U9782 (N_9782,N_1813,N_4773);
and U9783 (N_9783,N_2184,N_3432);
nor U9784 (N_9784,N_2720,N_714);
nand U9785 (N_9785,N_270,N_469);
and U9786 (N_9786,N_4990,N_3301);
nor U9787 (N_9787,N_186,N_275);
and U9788 (N_9788,N_4237,N_1393);
and U9789 (N_9789,N_4377,N_4304);
nor U9790 (N_9790,N_3182,N_594);
and U9791 (N_9791,N_3531,N_3042);
nor U9792 (N_9792,N_1663,N_3796);
or U9793 (N_9793,N_394,N_1892);
and U9794 (N_9794,N_4341,N_358);
or U9795 (N_9795,N_2120,N_4960);
nor U9796 (N_9796,N_4851,N_2292);
or U9797 (N_9797,N_1109,N_19);
nor U9798 (N_9798,N_1098,N_990);
and U9799 (N_9799,N_2883,N_538);
nand U9800 (N_9800,N_3261,N_837);
and U9801 (N_9801,N_3205,N_2004);
and U9802 (N_9802,N_2284,N_3136);
or U9803 (N_9803,N_2863,N_4334);
and U9804 (N_9804,N_1908,N_1491);
or U9805 (N_9805,N_3674,N_4983);
and U9806 (N_9806,N_1113,N_866);
and U9807 (N_9807,N_1084,N_2601);
and U9808 (N_9808,N_2053,N_4668);
nor U9809 (N_9809,N_340,N_4572);
and U9810 (N_9810,N_1603,N_555);
and U9811 (N_9811,N_1000,N_1307);
and U9812 (N_9812,N_4239,N_567);
or U9813 (N_9813,N_1251,N_27);
and U9814 (N_9814,N_4108,N_2397);
nor U9815 (N_9815,N_4112,N_971);
or U9816 (N_9816,N_272,N_3772);
and U9817 (N_9817,N_926,N_4327);
nor U9818 (N_9818,N_1098,N_1254);
and U9819 (N_9819,N_4115,N_597);
or U9820 (N_9820,N_1875,N_1617);
nand U9821 (N_9821,N_3641,N_1872);
nor U9822 (N_9822,N_4893,N_3151);
nand U9823 (N_9823,N_4082,N_1915);
nand U9824 (N_9824,N_4410,N_275);
or U9825 (N_9825,N_2469,N_3057);
and U9826 (N_9826,N_1525,N_776);
or U9827 (N_9827,N_2669,N_1537);
nand U9828 (N_9828,N_2935,N_4634);
nor U9829 (N_9829,N_1453,N_2265);
and U9830 (N_9830,N_732,N_1772);
nand U9831 (N_9831,N_1824,N_3085);
nand U9832 (N_9832,N_3183,N_3942);
nor U9833 (N_9833,N_2910,N_562);
nor U9834 (N_9834,N_4616,N_1578);
or U9835 (N_9835,N_444,N_1731);
or U9836 (N_9836,N_2174,N_3649);
nor U9837 (N_9837,N_882,N_1350);
nor U9838 (N_9838,N_1766,N_3015);
and U9839 (N_9839,N_4612,N_475);
nor U9840 (N_9840,N_2457,N_1293);
or U9841 (N_9841,N_4889,N_2913);
nand U9842 (N_9842,N_3763,N_1782);
nor U9843 (N_9843,N_4133,N_738);
and U9844 (N_9844,N_3268,N_3553);
nor U9845 (N_9845,N_1605,N_1811);
or U9846 (N_9846,N_2384,N_824);
and U9847 (N_9847,N_1061,N_510);
nand U9848 (N_9848,N_3755,N_129);
or U9849 (N_9849,N_1183,N_911);
and U9850 (N_9850,N_1496,N_1235);
nand U9851 (N_9851,N_1399,N_3398);
or U9852 (N_9852,N_4855,N_2378);
nand U9853 (N_9853,N_263,N_702);
xnor U9854 (N_9854,N_2461,N_3992);
nor U9855 (N_9855,N_1904,N_2690);
and U9856 (N_9856,N_2567,N_4048);
and U9857 (N_9857,N_2197,N_378);
nor U9858 (N_9858,N_1572,N_2707);
nor U9859 (N_9859,N_2622,N_4512);
or U9860 (N_9860,N_2932,N_1903);
or U9861 (N_9861,N_4971,N_2799);
and U9862 (N_9862,N_2260,N_270);
nor U9863 (N_9863,N_1138,N_4026);
or U9864 (N_9864,N_3561,N_3907);
nand U9865 (N_9865,N_3235,N_1425);
and U9866 (N_9866,N_63,N_854);
nor U9867 (N_9867,N_424,N_1022);
or U9868 (N_9868,N_2331,N_3909);
and U9869 (N_9869,N_1964,N_3905);
nand U9870 (N_9870,N_1038,N_3171);
nor U9871 (N_9871,N_2649,N_2301);
nor U9872 (N_9872,N_239,N_2548);
nand U9873 (N_9873,N_4209,N_2649);
nand U9874 (N_9874,N_488,N_142);
nor U9875 (N_9875,N_1192,N_2035);
and U9876 (N_9876,N_1663,N_152);
or U9877 (N_9877,N_4205,N_377);
nand U9878 (N_9878,N_4278,N_1503);
or U9879 (N_9879,N_1301,N_2149);
or U9880 (N_9880,N_1117,N_885);
nor U9881 (N_9881,N_2236,N_105);
and U9882 (N_9882,N_1192,N_2484);
nand U9883 (N_9883,N_927,N_1255);
or U9884 (N_9884,N_1157,N_1774);
nand U9885 (N_9885,N_2822,N_1396);
nand U9886 (N_9886,N_2314,N_2484);
and U9887 (N_9887,N_1513,N_248);
nand U9888 (N_9888,N_289,N_1532);
or U9889 (N_9889,N_3520,N_4047);
or U9890 (N_9890,N_4090,N_4700);
or U9891 (N_9891,N_1311,N_44);
or U9892 (N_9892,N_3156,N_3271);
and U9893 (N_9893,N_3830,N_2463);
nor U9894 (N_9894,N_3643,N_4949);
or U9895 (N_9895,N_1509,N_231);
and U9896 (N_9896,N_2045,N_1049);
and U9897 (N_9897,N_2109,N_4238);
nand U9898 (N_9898,N_2069,N_2061);
nand U9899 (N_9899,N_3019,N_3865);
or U9900 (N_9900,N_3023,N_206);
nand U9901 (N_9901,N_4290,N_3554);
nand U9902 (N_9902,N_4768,N_3660);
and U9903 (N_9903,N_4389,N_2743);
and U9904 (N_9904,N_4367,N_1488);
and U9905 (N_9905,N_3632,N_4889);
nand U9906 (N_9906,N_2574,N_3668);
and U9907 (N_9907,N_446,N_868);
or U9908 (N_9908,N_4095,N_632);
and U9909 (N_9909,N_1812,N_3694);
and U9910 (N_9910,N_3910,N_2927);
and U9911 (N_9911,N_2393,N_4408);
and U9912 (N_9912,N_4889,N_4602);
nor U9913 (N_9913,N_1223,N_4069);
nand U9914 (N_9914,N_682,N_3335);
and U9915 (N_9915,N_3073,N_228);
and U9916 (N_9916,N_2860,N_878);
or U9917 (N_9917,N_4416,N_4440);
nand U9918 (N_9918,N_2696,N_1005);
nor U9919 (N_9919,N_2813,N_470);
and U9920 (N_9920,N_3090,N_799);
and U9921 (N_9921,N_1481,N_1400);
nor U9922 (N_9922,N_4129,N_1720);
nor U9923 (N_9923,N_980,N_1866);
or U9924 (N_9924,N_4648,N_3070);
or U9925 (N_9925,N_1528,N_658);
and U9926 (N_9926,N_1587,N_3678);
nand U9927 (N_9927,N_365,N_2843);
nor U9928 (N_9928,N_865,N_3522);
nor U9929 (N_9929,N_3467,N_3044);
nor U9930 (N_9930,N_1940,N_1087);
nand U9931 (N_9931,N_4271,N_1694);
and U9932 (N_9932,N_2929,N_1991);
nor U9933 (N_9933,N_1169,N_1020);
and U9934 (N_9934,N_4644,N_4996);
nand U9935 (N_9935,N_4512,N_3004);
nand U9936 (N_9936,N_3204,N_4086);
nand U9937 (N_9937,N_3508,N_3775);
nand U9938 (N_9938,N_1158,N_1911);
and U9939 (N_9939,N_1171,N_1082);
nand U9940 (N_9940,N_2460,N_4566);
nand U9941 (N_9941,N_875,N_1859);
nor U9942 (N_9942,N_1182,N_4489);
nand U9943 (N_9943,N_3168,N_924);
nand U9944 (N_9944,N_2005,N_2059);
nor U9945 (N_9945,N_3819,N_3816);
xor U9946 (N_9946,N_3967,N_952);
nor U9947 (N_9947,N_988,N_2756);
or U9948 (N_9948,N_470,N_3663);
nor U9949 (N_9949,N_1432,N_4700);
or U9950 (N_9950,N_2853,N_1337);
or U9951 (N_9951,N_1265,N_1190);
nand U9952 (N_9952,N_817,N_645);
nand U9953 (N_9953,N_2495,N_468);
nand U9954 (N_9954,N_377,N_2625);
or U9955 (N_9955,N_2128,N_193);
nor U9956 (N_9956,N_4213,N_4303);
and U9957 (N_9957,N_2350,N_507);
and U9958 (N_9958,N_1981,N_4334);
nor U9959 (N_9959,N_2433,N_414);
nor U9960 (N_9960,N_2503,N_1828);
and U9961 (N_9961,N_1179,N_3737);
or U9962 (N_9962,N_4270,N_3702);
or U9963 (N_9963,N_1344,N_1817);
and U9964 (N_9964,N_3491,N_1580);
nor U9965 (N_9965,N_3670,N_4622);
nor U9966 (N_9966,N_3661,N_1623);
nand U9967 (N_9967,N_76,N_3356);
and U9968 (N_9968,N_2045,N_4556);
nor U9969 (N_9969,N_965,N_977);
nand U9970 (N_9970,N_3748,N_3073);
nor U9971 (N_9971,N_4298,N_3143);
xor U9972 (N_9972,N_1700,N_2147);
nand U9973 (N_9973,N_3446,N_1075);
nor U9974 (N_9974,N_4306,N_4545);
nand U9975 (N_9975,N_3197,N_4722);
nand U9976 (N_9976,N_251,N_1988);
nand U9977 (N_9977,N_2261,N_365);
and U9978 (N_9978,N_1116,N_1455);
nor U9979 (N_9979,N_1224,N_1257);
or U9980 (N_9980,N_3582,N_2512);
or U9981 (N_9981,N_4000,N_607);
or U9982 (N_9982,N_2362,N_4552);
and U9983 (N_9983,N_1936,N_1921);
nand U9984 (N_9984,N_1464,N_2484);
nand U9985 (N_9985,N_1210,N_1028);
nand U9986 (N_9986,N_4600,N_2780);
nor U9987 (N_9987,N_1371,N_4306);
and U9988 (N_9988,N_1137,N_2036);
or U9989 (N_9989,N_1639,N_4880);
nor U9990 (N_9990,N_2822,N_3815);
nand U9991 (N_9991,N_4235,N_2939);
nor U9992 (N_9992,N_3899,N_1088);
nand U9993 (N_9993,N_417,N_134);
nand U9994 (N_9994,N_3223,N_3606);
nand U9995 (N_9995,N_898,N_484);
nor U9996 (N_9996,N_3006,N_4525);
or U9997 (N_9997,N_760,N_1637);
or U9998 (N_9998,N_3526,N_4399);
nand U9999 (N_9999,N_45,N_982);
nor UO_0 (O_0,N_9686,N_9403);
nor UO_1 (O_1,N_5684,N_7062);
nand UO_2 (O_2,N_9025,N_7969);
nand UO_3 (O_3,N_8971,N_7994);
nand UO_4 (O_4,N_7185,N_5850);
nand UO_5 (O_5,N_7478,N_5802);
nor UO_6 (O_6,N_5726,N_6708);
nor UO_7 (O_7,N_6286,N_9252);
nor UO_8 (O_8,N_6086,N_9189);
nand UO_9 (O_9,N_9317,N_9114);
nor UO_10 (O_10,N_5887,N_6328);
and UO_11 (O_11,N_7581,N_5768);
or UO_12 (O_12,N_5190,N_6726);
nand UO_13 (O_13,N_5324,N_5013);
nor UO_14 (O_14,N_9571,N_5408);
nor UO_15 (O_15,N_5737,N_6850);
and UO_16 (O_16,N_6514,N_6002);
nand UO_17 (O_17,N_7670,N_6497);
and UO_18 (O_18,N_8234,N_5291);
or UO_19 (O_19,N_7584,N_9090);
or UO_20 (O_20,N_8317,N_6021);
nor UO_21 (O_21,N_9168,N_5168);
and UO_22 (O_22,N_9338,N_7724);
and UO_23 (O_23,N_7431,N_7597);
or UO_24 (O_24,N_9225,N_6238);
or UO_25 (O_25,N_6954,N_8526);
nand UO_26 (O_26,N_9823,N_9272);
or UO_27 (O_27,N_8373,N_8909);
and UO_28 (O_28,N_8865,N_6487);
and UO_29 (O_29,N_9246,N_6431);
nand UO_30 (O_30,N_6541,N_9832);
or UO_31 (O_31,N_9986,N_6999);
nor UO_32 (O_32,N_9611,N_8030);
nand UO_33 (O_33,N_6396,N_9532);
nor UO_34 (O_34,N_6660,N_9794);
and UO_35 (O_35,N_7685,N_6244);
and UO_36 (O_36,N_9348,N_9300);
nor UO_37 (O_37,N_7818,N_8149);
or UO_38 (O_38,N_9274,N_6160);
nor UO_39 (O_39,N_6118,N_8981);
and UO_40 (O_40,N_5963,N_8578);
nor UO_41 (O_41,N_8276,N_8318);
nor UO_42 (O_42,N_8780,N_9449);
or UO_43 (O_43,N_8035,N_7980);
nand UO_44 (O_44,N_8342,N_5480);
or UO_45 (O_45,N_6947,N_8880);
and UO_46 (O_46,N_6608,N_8139);
nand UO_47 (O_47,N_8518,N_8481);
nor UO_48 (O_48,N_7860,N_9562);
nand UO_49 (O_49,N_8912,N_9737);
nor UO_50 (O_50,N_8290,N_8701);
or UO_51 (O_51,N_5331,N_8224);
and UO_52 (O_52,N_5389,N_8019);
nor UO_53 (O_53,N_7651,N_9254);
or UO_54 (O_54,N_9067,N_6776);
nor UO_55 (O_55,N_6820,N_5241);
nor UO_56 (O_56,N_6449,N_9164);
and UO_57 (O_57,N_7666,N_7618);
nor UO_58 (O_58,N_8455,N_9423);
or UO_59 (O_59,N_6178,N_8013);
nand UO_60 (O_60,N_6437,N_8037);
or UO_61 (O_61,N_5580,N_5263);
and UO_62 (O_62,N_6798,N_8836);
nand UO_63 (O_63,N_8848,N_6029);
nand UO_64 (O_64,N_6050,N_9869);
nand UO_65 (O_65,N_5335,N_5565);
nor UO_66 (O_66,N_6283,N_9646);
or UO_67 (O_67,N_9668,N_7540);
and UO_68 (O_68,N_9316,N_5567);
or UO_69 (O_69,N_5847,N_6680);
nor UO_70 (O_70,N_5513,N_8334);
and UO_71 (O_71,N_8169,N_6827);
or UO_72 (O_72,N_9065,N_5119);
or UO_73 (O_73,N_9356,N_6556);
nand UO_74 (O_74,N_9007,N_6241);
nor UO_75 (O_75,N_7078,N_9868);
and UO_76 (O_76,N_7226,N_5627);
nand UO_77 (O_77,N_6205,N_5999);
or UO_78 (O_78,N_9401,N_6710);
nand UO_79 (O_79,N_9191,N_6550);
nor UO_80 (O_80,N_9992,N_7481);
or UO_81 (O_81,N_5148,N_9564);
or UO_82 (O_82,N_7641,N_6394);
or UO_83 (O_83,N_5778,N_7875);
nor UO_84 (O_84,N_5258,N_9216);
and UO_85 (O_85,N_8284,N_8304);
and UO_86 (O_86,N_7331,N_6853);
or UO_87 (O_87,N_5920,N_5493);
and UO_88 (O_88,N_8840,N_9364);
or UO_89 (O_89,N_8313,N_6572);
and UO_90 (O_90,N_5419,N_6662);
nand UO_91 (O_91,N_6285,N_7706);
nand UO_92 (O_92,N_8468,N_6518);
nor UO_93 (O_93,N_9163,N_6398);
or UO_94 (O_94,N_5036,N_5162);
and UO_95 (O_95,N_8914,N_6653);
nor UO_96 (O_96,N_6494,N_7775);
or UO_97 (O_97,N_6949,N_6875);
and UO_98 (O_98,N_6735,N_8948);
and UO_99 (O_99,N_7887,N_9087);
nand UO_100 (O_100,N_7275,N_9277);
and UO_101 (O_101,N_6416,N_8670);
and UO_102 (O_102,N_7323,N_8888);
nor UO_103 (O_103,N_8967,N_5800);
or UO_104 (O_104,N_5523,N_6800);
or UO_105 (O_105,N_5197,N_6466);
nand UO_106 (O_106,N_7156,N_8921);
or UO_107 (O_107,N_6485,N_6970);
or UO_108 (O_108,N_5556,N_7788);
and UO_109 (O_109,N_8849,N_8055);
or UO_110 (O_110,N_6352,N_8655);
and UO_111 (O_111,N_7038,N_8159);
nand UO_112 (O_112,N_8011,N_6834);
nand UO_113 (O_113,N_6807,N_6441);
nand UO_114 (O_114,N_7375,N_9526);
nor UO_115 (O_115,N_7059,N_7332);
nand UO_116 (O_116,N_5485,N_5441);
or UO_117 (O_117,N_9559,N_5630);
nor UO_118 (O_118,N_5128,N_6468);
nor UO_119 (O_119,N_9700,N_7872);
nor UO_120 (O_120,N_9514,N_7088);
and UO_121 (O_121,N_9952,N_6705);
or UO_122 (O_122,N_8475,N_5172);
nor UO_123 (O_123,N_6706,N_5863);
nor UO_124 (O_124,N_7210,N_5189);
nand UO_125 (O_125,N_7535,N_7491);
nand UO_126 (O_126,N_7648,N_6276);
or UO_127 (O_127,N_9783,N_8144);
nor UO_128 (O_128,N_7679,N_9578);
and UO_129 (O_129,N_5075,N_8765);
nand UO_130 (O_130,N_7640,N_7264);
or UO_131 (O_131,N_7205,N_6020);
nor UO_132 (O_132,N_7054,N_8513);
nor UO_133 (O_133,N_6410,N_8077);
or UO_134 (O_134,N_9570,N_8557);
nor UO_135 (O_135,N_5175,N_5058);
and UO_136 (O_136,N_5600,N_5210);
nand UO_137 (O_137,N_5846,N_8316);
nand UO_138 (O_138,N_7838,N_7855);
or UO_139 (O_139,N_9260,N_9921);
or UO_140 (O_140,N_7978,N_8874);
nand UO_141 (O_141,N_7711,N_9071);
and UO_142 (O_142,N_7113,N_5555);
or UO_143 (O_143,N_9502,N_9419);
nand UO_144 (O_144,N_9402,N_5099);
and UO_145 (O_145,N_9619,N_5299);
nor UO_146 (O_146,N_6240,N_5327);
or UO_147 (O_147,N_5173,N_7765);
nor UO_148 (O_148,N_7119,N_9516);
nand UO_149 (O_149,N_7506,N_9670);
xnor UO_150 (O_150,N_7453,N_5717);
nor UO_151 (O_151,N_9733,N_8173);
nor UO_152 (O_152,N_7793,N_8106);
nor UO_153 (O_153,N_8076,N_7663);
and UO_154 (O_154,N_9698,N_6440);
nor UO_155 (O_155,N_6887,N_8141);
or UO_156 (O_156,N_9209,N_9266);
nor UO_157 (O_157,N_6661,N_6009);
nand UO_158 (O_158,N_5363,N_6505);
or UO_159 (O_159,N_6771,N_9273);
nand UO_160 (O_160,N_7722,N_7090);
nor UO_161 (O_161,N_9996,N_9424);
nand UO_162 (O_162,N_5370,N_9186);
xnor UO_163 (O_163,N_8209,N_7399);
and UO_164 (O_164,N_6072,N_5704);
or UO_165 (O_165,N_5640,N_5552);
and UO_166 (O_166,N_7668,N_7988);
and UO_167 (O_167,N_5096,N_7507);
nand UO_168 (O_168,N_5361,N_6052);
nand UO_169 (O_169,N_6811,N_5870);
or UO_170 (O_170,N_9490,N_9411);
nor UO_171 (O_171,N_9194,N_5215);
and UO_172 (O_172,N_6749,N_7058);
nor UO_173 (O_173,N_6469,N_5071);
and UO_174 (O_174,N_5614,N_6473);
and UO_175 (O_175,N_8222,N_7509);
nand UO_176 (O_176,N_8353,N_7099);
and UO_177 (O_177,N_6450,N_6134);
or UO_178 (O_178,N_6108,N_9732);
nand UO_179 (O_179,N_8932,N_9534);
and UO_180 (O_180,N_9658,N_8550);
or UO_181 (O_181,N_8768,N_9543);
nand UO_182 (O_182,N_5406,N_6625);
nand UO_183 (O_183,N_9941,N_7510);
or UO_184 (O_184,N_9734,N_5725);
nor UO_185 (O_185,N_8985,N_9031);
nand UO_186 (O_186,N_9097,N_6979);
and UO_187 (O_187,N_5385,N_6388);
nand UO_188 (O_188,N_9776,N_9000);
nand UO_189 (O_189,N_5558,N_9192);
nand UO_190 (O_190,N_6075,N_6775);
or UO_191 (O_191,N_5392,N_8669);
and UO_192 (O_192,N_6768,N_5752);
nand UO_193 (O_193,N_9682,N_5618);
nand UO_194 (O_194,N_8328,N_9594);
nand UO_195 (O_195,N_9426,N_9236);
and UO_196 (O_196,N_9760,N_5824);
nand UO_197 (O_197,N_5223,N_8123);
nand UO_198 (O_198,N_7891,N_6913);
or UO_199 (O_199,N_7699,N_9220);
nand UO_200 (O_200,N_5158,N_7394);
nand UO_201 (O_201,N_9711,N_6833);
or UO_202 (O_202,N_6089,N_8769);
nor UO_203 (O_203,N_9204,N_5702);
and UO_204 (O_204,N_5689,N_6770);
and UO_205 (O_205,N_5193,N_5268);
or UO_206 (O_206,N_5753,N_8799);
and UO_207 (O_207,N_8908,N_8790);
or UO_208 (O_208,N_7594,N_5089);
nand UO_209 (O_209,N_8125,N_7716);
or UO_210 (O_210,N_8938,N_7476);
nand UO_211 (O_211,N_8961,N_7463);
or UO_212 (O_212,N_5893,N_5652);
nand UO_213 (O_213,N_9590,N_7999);
or UO_214 (O_214,N_5891,N_5792);
nor UO_215 (O_215,N_6890,N_5364);
or UO_216 (O_216,N_7528,N_9595);
nand UO_217 (O_217,N_7292,N_6841);
and UO_218 (O_218,N_5211,N_8675);
nand UO_219 (O_219,N_6418,N_8315);
and UO_220 (O_220,N_5034,N_8476);
nand UO_221 (O_221,N_9215,N_6208);
nor UO_222 (O_222,N_5352,N_8746);
nor UO_223 (O_223,N_6737,N_7060);
nor UO_224 (O_224,N_7228,N_6733);
nand UO_225 (O_225,N_9556,N_8762);
or UO_226 (O_226,N_9971,N_8409);
or UO_227 (O_227,N_7846,N_8435);
and UO_228 (O_228,N_5719,N_8531);
and UO_229 (O_229,N_9550,N_6934);
and UO_230 (O_230,N_6526,N_5581);
or UO_231 (O_231,N_9349,N_5796);
nor UO_232 (O_232,N_8464,N_7754);
or UO_233 (O_233,N_8289,N_7080);
nand UO_234 (O_234,N_7250,N_9145);
nor UO_235 (O_235,N_7779,N_7384);
or UO_236 (O_236,N_9985,N_6647);
and UO_237 (O_237,N_5654,N_6976);
nor UO_238 (O_238,N_6822,N_5995);
nand UO_239 (O_239,N_9951,N_7773);
or UO_240 (O_240,N_8543,N_8177);
nand UO_241 (O_241,N_8639,N_5766);
nor UO_242 (O_242,N_7676,N_9098);
or UO_243 (O_243,N_5339,N_7559);
nand UO_244 (O_244,N_6364,N_7044);
and UO_245 (O_245,N_9774,N_7627);
and UO_246 (O_246,N_9903,N_6849);
nor UO_247 (O_247,N_5199,N_8621);
nor UO_248 (O_248,N_6783,N_7385);
or UO_249 (O_249,N_7746,N_9415);
nand UO_250 (O_250,N_9956,N_9575);
nand UO_251 (O_251,N_8431,N_6985);
nor UO_252 (O_252,N_5804,N_7885);
nand UO_253 (O_253,N_9435,N_9409);
or UO_254 (O_254,N_6991,N_5718);
nor UO_255 (O_255,N_5117,N_7012);
and UO_256 (O_256,N_7452,N_5218);
and UO_257 (O_257,N_7374,N_8015);
nand UO_258 (O_258,N_6324,N_7516);
or UO_259 (O_259,N_9916,N_8158);
nor UO_260 (O_260,N_6829,N_8422);
nor UO_261 (O_261,N_5711,N_7284);
or UO_262 (O_262,N_5468,N_6353);
nor UO_263 (O_263,N_8324,N_7810);
nand UO_264 (O_264,N_7175,N_9059);
and UO_265 (O_265,N_9885,N_8038);
or UO_266 (O_266,N_9281,N_7958);
or UO_267 (O_267,N_5458,N_8761);
or UO_268 (O_268,N_6476,N_9879);
or UO_269 (O_269,N_6200,N_9487);
nand UO_270 (O_270,N_7592,N_8403);
nand UO_271 (O_271,N_7564,N_8446);
or UO_272 (O_272,N_7282,N_8868);
nand UO_273 (O_273,N_6078,N_6684);
nor UO_274 (O_274,N_5966,N_8171);
and UO_275 (O_275,N_8206,N_8372);
nor UO_276 (O_276,N_8052,N_9875);
nand UO_277 (O_277,N_8617,N_7072);
and UO_278 (O_278,N_6683,N_6033);
nor UO_279 (O_279,N_8584,N_9328);
or UO_280 (O_280,N_6851,N_7360);
nor UO_281 (O_281,N_9808,N_9144);
and UO_282 (O_282,N_9631,N_9661);
or UO_283 (O_283,N_8295,N_6498);
nor UO_284 (O_284,N_6763,N_6609);
nor UO_285 (O_285,N_8140,N_9036);
and UO_286 (O_286,N_9926,N_5350);
and UO_287 (O_287,N_6370,N_7993);
nor UO_288 (O_288,N_8825,N_9881);
or UO_289 (O_289,N_9029,N_6342);
nand UO_290 (O_290,N_9662,N_6983);
or UO_291 (O_291,N_9560,N_9171);
nor UO_292 (O_292,N_6098,N_7112);
and UO_293 (O_293,N_6998,N_9458);
or UO_294 (O_294,N_7790,N_9890);
nand UO_295 (O_295,N_6793,N_7174);
nor UO_296 (O_296,N_9958,N_9462);
nand UO_297 (O_297,N_6835,N_5703);
nand UO_298 (O_298,N_6138,N_6993);
nor UO_299 (O_299,N_6452,N_5054);
nor UO_300 (O_300,N_9864,N_6839);
nand UO_301 (O_301,N_5252,N_8470);
nand UO_302 (O_302,N_9810,N_5878);
and UO_303 (O_303,N_5225,N_8837);
and UO_304 (O_304,N_6090,N_7221);
or UO_305 (O_305,N_5839,N_7525);
and UO_306 (O_306,N_8649,N_5420);
nor UO_307 (O_307,N_9858,N_5247);
and UO_308 (O_308,N_5639,N_9505);
nand UO_309 (O_309,N_5732,N_9841);
or UO_310 (O_310,N_8340,N_8124);
or UO_311 (O_311,N_5574,N_9327);
and UO_312 (O_312,N_6799,N_9637);
or UO_313 (O_313,N_7290,N_5476);
or UO_314 (O_314,N_9857,N_5355);
and UO_315 (O_315,N_5811,N_9363);
nor UO_316 (O_316,N_6067,N_6109);
xnor UO_317 (O_317,N_9758,N_5019);
and UO_318 (O_318,N_9250,N_6198);
nand UO_319 (O_319,N_7857,N_9080);
and UO_320 (O_320,N_8569,N_7364);
nand UO_321 (O_321,N_6920,N_7029);
nor UO_322 (O_322,N_7419,N_8867);
nand UO_323 (O_323,N_5705,N_7124);
and UO_324 (O_324,N_9888,N_6825);
and UO_325 (O_325,N_5470,N_8823);
and UO_326 (O_326,N_6711,N_5050);
nor UO_327 (O_327,N_7459,N_5923);
nand UO_328 (O_328,N_8116,N_9513);
nor UO_329 (O_329,N_9337,N_8219);
and UO_330 (O_330,N_7222,N_8764);
or UO_331 (O_331,N_6966,N_6459);
nand UO_332 (O_332,N_9877,N_7574);
or UO_333 (O_333,N_9443,N_5216);
and UO_334 (O_334,N_5312,N_6821);
and UO_335 (O_335,N_8410,N_5068);
nor UO_336 (O_336,N_6562,N_8078);
and UO_337 (O_337,N_6577,N_5032);
or UO_338 (O_338,N_6219,N_5965);
nand UO_339 (O_339,N_9024,N_6615);
nor UO_340 (O_340,N_6560,N_5947);
nor UO_341 (O_341,N_9805,N_9261);
nor UO_342 (O_342,N_8103,N_8433);
nand UO_343 (O_343,N_8311,N_8873);
nand UO_344 (O_344,N_5576,N_8390);
nand UO_345 (O_345,N_5914,N_5592);
nand UO_346 (O_346,N_8969,N_8785);
nor UO_347 (O_347,N_7515,N_7424);
nand UO_348 (O_348,N_7457,N_8508);
nand UO_349 (O_349,N_7954,N_7024);
nand UO_350 (O_350,N_5516,N_8120);
nand UO_351 (O_351,N_7938,N_8230);
and UO_352 (O_352,N_9016,N_7154);
nand UO_353 (O_353,N_7998,N_5590);
nand UO_354 (O_354,N_7986,N_8916);
and UO_355 (O_355,N_5960,N_8192);
and UO_356 (O_356,N_6153,N_6216);
nand UO_357 (O_357,N_7203,N_8889);
or UO_358 (O_358,N_5400,N_6766);
nor UO_359 (O_359,N_6412,N_6861);
xnor UO_360 (O_360,N_5213,N_9492);
and UO_361 (O_361,N_8412,N_8747);
or UO_362 (O_362,N_5646,N_9035);
and UO_363 (O_363,N_9908,N_5272);
nand UO_364 (O_364,N_7046,N_6015);
and UO_365 (O_365,N_5394,N_7695);
and UO_366 (O_366,N_9285,N_5981);
or UO_367 (O_367,N_5530,N_5706);
or UO_368 (O_368,N_6338,N_6912);
nand UO_369 (O_369,N_7319,N_8101);
or UO_370 (O_370,N_8516,N_6652);
nand UO_371 (O_371,N_9838,N_9353);
nand UO_372 (O_372,N_7182,N_7805);
and UO_373 (O_373,N_6266,N_7079);
nand UO_374 (O_374,N_8520,N_8216);
nor UO_375 (O_375,N_5212,N_6040);
and UO_376 (O_376,N_5860,N_7251);
nor UO_377 (O_377,N_6553,N_8269);
or UO_378 (O_378,N_5345,N_6159);
nor UO_379 (O_379,N_9600,N_9053);
nor UO_380 (O_380,N_9673,N_5055);
or UO_381 (O_381,N_8203,N_9507);
or UO_382 (O_382,N_8138,N_7101);
and UO_383 (O_383,N_5510,N_5267);
nand UO_384 (O_384,N_6986,N_7216);
nand UO_385 (O_385,N_6061,N_8729);
nand UO_386 (O_386,N_8211,N_8479);
nor UO_387 (O_387,N_7977,N_9775);
or UO_388 (O_388,N_5396,N_9048);
and UO_389 (O_389,N_5713,N_5518);
nor UO_390 (O_390,N_7190,N_5319);
nand UO_391 (O_391,N_8707,N_7092);
nand UO_392 (O_392,N_7145,N_9837);
and UO_393 (O_393,N_7026,N_5201);
or UO_394 (O_394,N_6211,N_5155);
or UO_395 (O_395,N_9953,N_5823);
or UO_396 (O_396,N_7278,N_8565);
nand UO_397 (O_397,N_8990,N_7837);
and UO_398 (O_398,N_5791,N_9150);
nand UO_399 (O_399,N_7249,N_8355);
xnor UO_400 (O_400,N_6975,N_9685);
nand UO_401 (O_401,N_8056,N_8453);
nand UO_402 (O_402,N_5484,N_5275);
nand UO_403 (O_403,N_7981,N_7701);
and UO_404 (O_404,N_7265,N_6689);
and UO_405 (O_405,N_6929,N_5340);
or UO_406 (O_406,N_8757,N_9862);
nand UO_407 (O_407,N_9621,N_9970);
and UO_408 (O_408,N_6023,N_6651);
nand UO_409 (O_409,N_6731,N_5970);
nor UO_410 (O_410,N_5783,N_8751);
or UO_411 (O_411,N_7253,N_7611);
or UO_412 (O_412,N_9296,N_6965);
nand UO_413 (O_413,N_7570,N_9179);
nand UO_414 (O_414,N_6959,N_5820);
nor UO_415 (O_415,N_9015,N_6532);
or UO_416 (O_416,N_9520,N_7612);
nor UO_417 (O_417,N_8310,N_8620);
or UO_418 (O_418,N_5294,N_7379);
nand UO_419 (O_419,N_5296,N_7814);
nor UO_420 (O_420,N_7106,N_6495);
nand UO_421 (O_421,N_5375,N_7839);
and UO_422 (O_422,N_7373,N_8093);
nor UO_423 (O_423,N_7126,N_8946);
nor UO_424 (O_424,N_7461,N_9452);
and UO_425 (O_425,N_9284,N_6464);
or UO_426 (O_426,N_9131,N_9213);
or UO_427 (O_427,N_6826,N_6719);
nand UO_428 (O_428,N_9535,N_7952);
nand UO_429 (O_429,N_9023,N_6808);
and UO_430 (O_430,N_7285,N_6903);
or UO_431 (O_431,N_6539,N_6107);
and UO_432 (O_432,N_6003,N_5332);
nor UO_433 (O_433,N_6483,N_8406);
and UO_434 (O_434,N_8187,N_9551);
and UO_435 (O_435,N_9628,N_8536);
and UO_436 (O_436,N_7252,N_8388);
or UO_437 (O_437,N_6784,N_9795);
nor UO_438 (O_438,N_5833,N_9644);
nor UO_439 (O_439,N_9269,N_7191);
and UO_440 (O_440,N_8156,N_5787);
or UO_441 (O_441,N_6641,N_8198);
or UO_442 (O_442,N_5368,N_6239);
and UO_443 (O_443,N_5100,N_9601);
nor UO_444 (O_444,N_7966,N_8775);
and UO_445 (O_445,N_8819,N_5975);
and UO_446 (O_446,N_5894,N_8245);
and UO_447 (O_447,N_7542,N_6404);
nor UO_448 (O_448,N_5908,N_5478);
nand UO_449 (O_449,N_9822,N_6128);
nor UO_450 (O_450,N_6312,N_9480);
and UO_451 (O_451,N_7806,N_7883);
and UO_452 (O_452,N_6848,N_9368);
nor UO_453 (O_453,N_8534,N_5414);
nor UO_454 (O_454,N_7325,N_9472);
or UO_455 (O_455,N_7223,N_6669);
nor UO_456 (O_456,N_9581,N_5683);
or UO_457 (O_457,N_5451,N_6036);
or UO_458 (O_458,N_5380,N_5972);
nor UO_459 (O_459,N_6831,N_9641);
or UO_460 (O_460,N_9624,N_7889);
nor UO_461 (O_461,N_5911,N_5864);
nand UO_462 (O_462,N_7454,N_5221);
nor UO_463 (O_463,N_8693,N_9371);
nor UO_464 (O_464,N_6872,N_7635);
and UO_465 (O_465,N_6792,N_8277);
nand UO_466 (O_466,N_8885,N_5519);
or UO_467 (O_467,N_8692,N_6399);
and UO_468 (O_468,N_9287,N_9955);
or UO_469 (O_469,N_6112,N_8977);
nor UO_470 (O_470,N_5943,N_7517);
or UO_471 (O_471,N_5935,N_6585);
nor UO_472 (O_472,N_5644,N_6369);
and UO_473 (O_473,N_9583,N_8312);
nand UO_474 (O_474,N_6011,N_7582);
nor UO_475 (O_475,N_6335,N_5379);
and UO_476 (O_476,N_7601,N_8890);
and UO_477 (O_477,N_7927,N_8448);
and UO_478 (O_478,N_5632,N_9859);
or UO_479 (O_479,N_9033,N_6039);
or UO_480 (O_480,N_5235,N_5903);
or UO_481 (O_481,N_5940,N_5301);
nand UO_482 (O_482,N_9085,N_9651);
or UO_483 (O_483,N_5035,N_8439);
nand UO_484 (O_484,N_5060,N_7403);
and UO_485 (O_485,N_7393,N_8163);
or UO_486 (O_486,N_9099,N_8993);
nor UO_487 (O_487,N_7686,N_8529);
and UO_488 (O_488,N_6629,N_9940);
nor UO_489 (O_489,N_5390,N_7937);
and UO_490 (O_490,N_5877,N_5769);
or UO_491 (O_491,N_6867,N_7577);
or UO_492 (O_492,N_6589,N_6860);
and UO_493 (O_493,N_8727,N_8734);
nor UO_494 (O_494,N_5727,N_7492);
and UO_495 (O_495,N_9456,N_6115);
nor UO_496 (O_496,N_5374,N_5821);
nand UO_497 (O_497,N_9539,N_5421);
or UO_498 (O_498,N_8387,N_8766);
nand UO_499 (O_499,N_5907,N_7743);
nor UO_500 (O_500,N_8660,N_7484);
or UO_501 (O_501,N_8283,N_5164);
and UO_502 (O_502,N_8533,N_7503);
nor UO_503 (O_503,N_5261,N_7742);
nor UO_504 (O_504,N_5397,N_6794);
nand UO_505 (O_505,N_6150,N_9796);
and UO_506 (O_506,N_5171,N_9814);
and UO_507 (O_507,N_7925,N_7854);
nor UO_508 (O_508,N_7858,N_7085);
and UO_509 (O_509,N_9965,N_5777);
or UO_510 (O_510,N_7940,N_5569);
or UO_511 (O_511,N_6681,N_8263);
or UO_512 (O_512,N_5641,N_5563);
nand UO_513 (O_513,N_8683,N_7115);
or UO_514 (O_514,N_9899,N_5404);
and UO_515 (O_515,N_9634,N_6308);
and UO_516 (O_516,N_6673,N_7614);
xnor UO_517 (O_517,N_7412,N_5952);
and UO_518 (O_518,N_5187,N_9185);
or UO_519 (O_519,N_9103,N_9753);
nand UO_520 (O_520,N_7951,N_6503);
or UO_521 (O_521,N_9135,N_5738);
nand UO_522 (O_522,N_5194,N_6712);
or UO_523 (O_523,N_6041,N_8121);
and UO_524 (O_524,N_8255,N_7644);
and UO_525 (O_525,N_5300,N_5798);
nand UO_526 (O_526,N_8074,N_7368);
nand UO_527 (O_527,N_6278,N_9196);
and UO_528 (O_528,N_8393,N_9647);
nand UO_529 (O_529,N_8204,N_5501);
or UO_530 (O_530,N_7802,N_8635);
nand UO_531 (O_531,N_9430,N_8861);
nand UO_532 (O_532,N_6902,N_9994);
or UO_533 (O_533,N_9101,N_8039);
and UO_534 (O_534,N_8329,N_6343);
and UO_535 (O_535,N_5764,N_8205);
or UO_536 (O_536,N_9576,N_8275);
and UO_537 (O_537,N_6642,N_7086);
nand UO_538 (O_538,N_7930,N_9467);
or UO_539 (O_539,N_9598,N_7254);
or UO_540 (O_540,N_7776,N_7888);
or UO_541 (O_541,N_7474,N_9398);
nor UO_542 (O_542,N_8178,N_8895);
nand UO_543 (O_543,N_5898,N_5544);
nor UO_544 (O_544,N_6666,N_6502);
nand UO_545 (O_545,N_7367,N_5526);
or UO_546 (O_546,N_6846,N_7941);
and UO_547 (O_547,N_8677,N_8365);
or UO_548 (O_548,N_7483,N_5239);
nor UO_549 (O_549,N_9613,N_5188);
or UO_550 (O_550,N_9835,N_9716);
and UO_551 (O_551,N_8148,N_7070);
nand UO_552 (O_552,N_7041,N_7893);
and UO_553 (O_553,N_6730,N_6062);
nor UO_554 (O_554,N_8114,N_5465);
or UO_555 (O_555,N_5376,N_7907);
or UO_556 (O_556,N_7926,N_5697);
or UO_557 (O_557,N_6535,N_9482);
or UO_558 (O_558,N_6525,N_7964);
nor UO_559 (O_559,N_8595,N_9844);
nor UO_560 (O_560,N_5655,N_6031);
or UO_561 (O_561,N_5104,N_7973);
nor UO_562 (O_562,N_5341,N_7000);
xnor UO_563 (O_563,N_7645,N_9175);
and UO_564 (O_564,N_7413,N_9126);
and UO_565 (O_565,N_5346,N_6878);
nand UO_566 (O_566,N_7864,N_8519);
nand UO_567 (O_567,N_7780,N_7168);
nand UO_568 (O_568,N_5152,N_7939);
nor UO_569 (O_569,N_9184,N_9157);
and UO_570 (O_570,N_6511,N_5295);
nand UO_571 (O_571,N_7524,N_5457);
nand UO_572 (O_572,N_5342,N_8678);
or UO_573 (O_573,N_6894,N_7017);
or UO_574 (O_574,N_7300,N_8725);
nand UO_575 (O_575,N_8637,N_8326);
or UO_576 (O_576,N_9904,N_9506);
and UO_577 (O_577,N_5742,N_9257);
or UO_578 (O_578,N_8032,N_6197);
and UO_579 (O_579,N_5979,N_7144);
nor UO_580 (O_580,N_8413,N_8842);
nor UO_581 (O_581,N_8847,N_6417);
nor UO_582 (O_582,N_8258,N_5454);
and UO_583 (O_583,N_7084,N_9652);
or UO_584 (O_584,N_6147,N_6687);
xor UO_585 (O_585,N_7322,N_5866);
or UO_586 (O_586,N_8063,N_8742);
nor UO_587 (O_587,N_6135,N_7703);
and UO_588 (O_588,N_5249,N_6524);
and UO_589 (O_589,N_8651,N_8073);
or UO_590 (O_590,N_7007,N_5997);
and UO_591 (O_591,N_5694,N_7397);
and UO_592 (O_592,N_7055,N_8415);
or UO_593 (O_593,N_6529,N_6720);
or UO_594 (O_594,N_5321,N_9809);
and UO_595 (O_595,N_7442,N_9178);
and UO_596 (O_596,N_9684,N_6893);
nand UO_597 (O_597,N_8152,N_7333);
and UO_598 (O_598,N_9224,N_8408);
nand UO_599 (O_599,N_8157,N_5656);
and UO_600 (O_600,N_8506,N_8924);
or UO_601 (O_601,N_5251,N_6260);
or UO_602 (O_602,N_7047,N_8385);
and UO_603 (O_603,N_5153,N_9587);
and UO_604 (O_604,N_8883,N_6773);
or UO_605 (O_605,N_8236,N_7266);
nand UO_606 (O_606,N_8092,N_5784);
nor UO_607 (O_607,N_8306,N_5896);
nor UO_608 (O_608,N_9508,N_5770);
nand UO_609 (O_609,N_5710,N_8054);
or UO_610 (O_610,N_9201,N_5464);
or UO_611 (O_611,N_6385,N_9812);
nor UO_612 (O_612,N_6513,N_8958);
and UO_613 (O_613,N_9945,N_5418);
or UO_614 (O_614,N_9064,N_7783);
or UO_615 (O_615,N_6183,N_5088);
or UO_616 (O_616,N_8859,N_9248);
and UO_617 (O_617,N_8665,N_9763);
nor UO_618 (O_618,N_8572,N_6114);
nand UO_619 (O_619,N_6695,N_8714);
and UO_620 (O_620,N_6310,N_9558);
and UO_621 (O_621,N_8086,N_7415);
or UO_622 (O_622,N_7896,N_9293);
nor UO_623 (O_623,N_7147,N_8911);
nand UO_624 (O_624,N_8695,N_7445);
and UO_625 (O_625,N_8694,N_6207);
and UO_626 (O_626,N_5140,N_5721);
and UO_627 (O_627,N_5874,N_5041);
nand UO_628 (O_628,N_6005,N_8427);
xor UO_629 (O_629,N_7016,N_8976);
nand UO_630 (O_630,N_6777,N_9709);
nand UO_631 (O_631,N_9385,N_9491);
or UO_632 (O_632,N_7406,N_6565);
nor UO_633 (O_633,N_7830,N_5775);
nor UO_634 (O_634,N_5714,N_7365);
nand UO_635 (O_635,N_5284,N_5483);
and UO_636 (O_636,N_9524,N_6739);
nor UO_637 (O_637,N_8134,N_9127);
or UO_638 (O_638,N_6877,N_7778);
nor UO_639 (O_639,N_8537,N_6928);
xnor UO_640 (O_640,N_6664,N_8089);
and UO_641 (O_641,N_9518,N_9470);
nand UO_642 (O_642,N_5449,N_8094);
nor UO_643 (O_643,N_6329,N_9517);
or UO_644 (O_644,N_9762,N_9463);
nor UO_645 (O_645,N_5635,N_5762);
nand UO_646 (O_646,N_5230,N_7104);
nor UO_647 (O_647,N_9149,N_5901);
nand UO_648 (O_648,N_7338,N_7572);
nor UO_649 (O_649,N_5698,N_8142);
and UO_650 (O_650,N_5888,N_9251);
or UO_651 (O_651,N_6180,N_9012);
nand UO_652 (O_652,N_9304,N_7541);
or UO_653 (O_653,N_8596,N_8830);
nand UO_654 (O_654,N_5942,N_6306);
and UO_655 (O_655,N_5442,N_5744);
or UO_656 (O_656,N_9278,N_8705);
and UO_657 (O_657,N_7303,N_9937);
nor UO_658 (O_658,N_6351,N_9866);
xor UO_659 (O_659,N_6463,N_9437);
nand UO_660 (O_660,N_5531,N_6038);
nor UO_661 (O_661,N_9542,N_9607);
nand UO_662 (O_662,N_8248,N_7318);
or UO_663 (O_663,N_5837,N_7848);
nand UO_664 (O_664,N_5146,N_7752);
nor UO_665 (O_665,N_6406,N_8900);
nor UO_666 (O_666,N_5809,N_5918);
nor UO_667 (O_667,N_5924,N_5078);
or UO_668 (O_668,N_5938,N_6806);
and UO_669 (O_669,N_5471,N_8443);
and UO_670 (O_670,N_5575,N_8379);
or UO_671 (O_671,N_7967,N_5948);
nor UO_672 (O_672,N_6374,N_7677);
nand UO_673 (O_673,N_5432,N_7179);
nor UO_674 (O_674,N_5735,N_7390);
or UO_675 (O_675,N_8502,N_7139);
nor UO_676 (O_676,N_8835,N_6533);
and UO_677 (O_677,N_6745,N_7330);
and UO_678 (O_678,N_5014,N_6217);
and UO_679 (O_679,N_7159,N_8510);
or UO_680 (O_680,N_7131,N_8023);
and UO_681 (O_681,N_6918,N_5667);
or UO_682 (O_682,N_5425,N_9856);
and UO_683 (O_683,N_9865,N_8349);
and UO_684 (O_684,N_5801,N_9643);
nand UO_685 (O_685,N_5381,N_5462);
nor UO_686 (O_686,N_6077,N_8528);
or UO_687 (O_687,N_6512,N_8221);
xor UO_688 (O_688,N_6282,N_8696);
nand UO_689 (O_689,N_8844,N_8656);
nor UO_690 (O_690,N_9793,N_9198);
and UO_691 (O_691,N_8362,N_9418);
nand UO_692 (O_692,N_5349,N_6423);
or UO_693 (O_693,N_5037,N_6597);
or UO_694 (O_694,N_7436,N_8604);
nor UO_695 (O_695,N_8759,N_5829);
nand UO_696 (O_696,N_8979,N_6769);
or UO_697 (O_697,N_6544,N_9440);
nand UO_698 (O_698,N_9820,N_5844);
and UO_699 (O_699,N_5927,N_5554);
nand UO_700 (O_700,N_6698,N_7215);
nand UO_701 (O_701,N_6069,N_8616);
and UO_702 (O_702,N_7551,N_9239);
nor UO_703 (O_703,N_9030,N_6475);
nor UO_704 (O_704,N_5749,N_6419);
and UO_705 (O_705,N_6791,N_7232);
and UO_706 (O_706,N_5372,N_8416);
or UO_707 (O_707,N_5817,N_7709);
nor UO_708 (O_708,N_9749,N_5665);
and UO_709 (O_709,N_7843,N_8264);
nor UO_710 (O_710,N_6000,N_6815);
nand UO_711 (O_711,N_9347,N_6696);
or UO_712 (O_712,N_5666,N_5548);
and UO_713 (O_713,N_7869,N_6637);
or UO_714 (O_714,N_8640,N_6355);
or UO_715 (O_715,N_6830,N_8208);
and UO_716 (O_716,N_8797,N_7089);
or UO_717 (O_717,N_5313,N_5834);
and UO_718 (O_718,N_5098,N_8629);
nor UO_719 (O_719,N_5459,N_5315);
nor UO_720 (O_720,N_5154,N_5603);
nand UO_721 (O_721,N_6043,N_6327);
nand UO_722 (O_722,N_9336,N_6523);
nand UO_723 (O_723,N_5551,N_8681);
nor UO_724 (O_724,N_5437,N_8605);
or UO_725 (O_725,N_5463,N_7421);
nand UO_726 (O_726,N_8779,N_8891);
or UO_727 (O_727,N_8625,N_6121);
or UO_728 (O_728,N_5048,N_7354);
or UO_729 (O_729,N_8688,N_9612);
nor UO_730 (O_730,N_9340,N_6156);
or UO_731 (O_731,N_8614,N_6409);
or UO_732 (O_732,N_9664,N_8802);
nand UO_733 (O_733,N_8252,N_5005);
nand UO_734 (O_734,N_7438,N_7262);
or UO_735 (O_735,N_6531,N_8395);
and UO_736 (O_736,N_7212,N_9155);
nor UO_737 (O_737,N_8361,N_6218);
or UO_738 (O_738,N_9061,N_7378);
nand UO_739 (O_739,N_9410,N_9330);
nand UO_740 (O_740,N_8813,N_8309);
and UO_741 (O_741,N_9109,N_9565);
nand UO_742 (O_742,N_7409,N_8057);
nand UO_743 (O_743,N_6246,N_6570);
nor UO_744 (O_744,N_6522,N_5750);
and UO_745 (O_745,N_6575,N_6623);
and UO_746 (O_746,N_7277,N_5309);
nand UO_747 (O_747,N_7849,N_8532);
or UO_748 (O_748,N_9152,N_5027);
or UO_749 (O_749,N_6717,N_7298);
and UO_750 (O_750,N_8700,N_8673);
nand UO_751 (O_751,N_9813,N_8723);
nand UO_752 (O_752,N_5450,N_5693);
nor UO_753 (O_753,N_6667,N_7991);
nor UO_754 (O_754,N_8796,N_7472);
nor UO_755 (O_755,N_8767,N_6175);
or UO_756 (O_756,N_8332,N_8787);
nand UO_757 (O_757,N_9406,N_9052);
and UO_758 (O_758,N_6931,N_5584);
nor UO_759 (O_759,N_7342,N_7289);
and UO_760 (O_760,N_9331,N_5120);
and UO_761 (O_761,N_5939,N_6648);
or UO_762 (O_762,N_6026,N_9222);
nand UO_763 (O_763,N_6559,N_5734);
and UO_764 (O_764,N_7659,N_6162);
nand UO_765 (O_765,N_9761,N_6271);
nor UO_766 (O_766,N_7610,N_5070);
nand UO_767 (O_767,N_7556,N_9792);
and UO_768 (O_768,N_5047,N_9380);
and UO_769 (O_769,N_6213,N_7575);
nand UO_770 (O_770,N_7717,N_9313);
and UO_771 (O_771,N_8085,N_5897);
nor UO_772 (O_772,N_8994,N_7508);
nand UO_773 (O_773,N_8703,N_9750);
or UO_774 (O_774,N_9392,N_9457);
or UO_775 (O_775,N_7263,N_5912);
nand UO_776 (O_776,N_9132,N_6674);
nor UO_777 (O_777,N_6095,N_5508);
and UO_778 (O_778,N_6756,N_9124);
nor UO_779 (O_779,N_5988,N_9689);
or UO_780 (O_780,N_6616,N_6964);
and UO_781 (O_781,N_9927,N_8348);
and UO_782 (O_782,N_7009,N_9383);
and UO_783 (O_783,N_5849,N_5546);
or UO_784 (O_784,N_8368,N_5009);
nand UO_785 (O_785,N_6300,N_7548);
and UO_786 (O_786,N_8319,N_9574);
nor UO_787 (O_787,N_8926,N_7048);
nor UO_788 (O_788,N_9976,N_9690);
nand UO_789 (O_789,N_8983,N_8065);
nor UO_790 (O_790,N_5277,N_6184);
nor UO_791 (O_791,N_9276,N_7151);
and UO_792 (O_792,N_9240,N_5862);
or UO_793 (O_793,N_8378,N_9917);
nor UO_794 (O_794,N_9143,N_9221);
nand UO_795 (O_795,N_7530,N_7656);
nand UO_796 (O_796,N_5305,N_7395);
nor UO_797 (O_797,N_9388,N_5517);
nand UO_798 (O_798,N_9102,N_8542);
and UO_799 (O_799,N_6738,N_9799);
nor UO_800 (O_800,N_6102,N_9084);
and UO_801 (O_801,N_6746,N_8343);
nor UO_802 (O_802,N_5871,N_8804);
nor UO_803 (O_803,N_5248,N_7123);
nand UO_804 (O_804,N_6154,N_5330);
nand UO_805 (O_805,N_7176,N_5557);
nand UO_806 (O_806,N_9717,N_5255);
and UO_807 (O_807,N_7555,N_6027);
and UO_808 (O_808,N_6704,N_8242);
nand UO_809 (O_809,N_5007,N_6141);
nor UO_810 (O_810,N_7235,N_5814);
nand UO_811 (O_811,N_6963,N_8008);
or UO_812 (O_812,N_6491,N_5566);
nor UO_813 (O_813,N_8210,N_8190);
nand UO_814 (O_814,N_8366,N_5080);
or UO_815 (O_815,N_5612,N_7696);
nand UO_816 (O_816,N_8225,N_6194);
or UO_817 (O_817,N_8499,N_5122);
and UO_818 (O_818,N_9270,N_6155);
and UO_819 (O_819,N_7359,N_6059);
nand UO_820 (O_820,N_9227,N_5074);
or UO_821 (O_821,N_9253,N_9525);
nand UO_822 (O_822,N_7613,N_7021);
nand UO_823 (O_823,N_6499,N_5522);
nor UO_824 (O_824,N_5334,N_7425);
nand UO_825 (O_825,N_8611,N_8603);
nor UO_826 (O_826,N_8690,N_5739);
xnor UO_827 (O_827,N_8246,N_9582);
nand UO_828 (O_828,N_5053,N_9489);
and UO_829 (O_829,N_6305,N_7796);
or UO_830 (O_830,N_5889,N_7957);
or UO_831 (O_831,N_7985,N_9924);
or UO_832 (O_832,N_6408,N_5647);
nor UO_833 (O_833,N_8112,N_9471);
nand UO_834 (O_834,N_7526,N_8394);
nand UO_835 (O_835,N_9798,N_5536);
nand UO_836 (O_836,N_7913,N_5695);
nor UO_837 (O_837,N_7918,N_5827);
or UO_838 (O_838,N_9998,N_7987);
nor UO_839 (O_839,N_8397,N_9663);
nor UO_840 (O_840,N_6935,N_8027);
nor UO_841 (O_841,N_7650,N_9553);
nand UO_842 (O_842,N_5090,N_6130);
and UO_843 (O_843,N_7240,N_6568);
nand UO_844 (O_844,N_8894,N_8195);
and UO_845 (O_845,N_6170,N_6953);
nand UO_846 (O_846,N_7170,N_7141);
nor UO_847 (O_847,N_7673,N_6037);
nand UO_848 (O_848,N_6933,N_8601);
and UO_849 (O_849,N_6018,N_5343);
or UO_850 (O_850,N_9190,N_5144);
nor UO_851 (O_851,N_9993,N_7646);
nor UO_852 (O_852,N_8568,N_6895);
nand UO_853 (O_853,N_9618,N_9360);
or UO_854 (O_854,N_5422,N_7593);
nor UO_855 (O_855,N_7349,N_7272);
nand UO_856 (O_856,N_7904,N_9804);
or UO_857 (O_857,N_7726,N_6250);
or UO_858 (O_858,N_9989,N_7653);
and UO_859 (O_859,N_5609,N_8180);
nand UO_860 (O_860,N_7989,N_7750);
nand UO_861 (O_861,N_7836,N_5622);
nor UO_862 (O_862,N_6486,N_9544);
or UO_863 (O_863,N_8915,N_5280);
nand UO_864 (O_864,N_5680,N_6507);
or UO_865 (O_865,N_6870,N_9256);
nand UO_866 (O_866,N_6937,N_5244);
nor UO_867 (O_867,N_7288,N_6085);
or UO_868 (O_868,N_5984,N_9112);
and UO_869 (O_869,N_8942,N_6678);
and UO_870 (O_870,N_5026,N_8197);
or UO_871 (O_871,N_6166,N_7688);
nand UO_872 (O_872,N_5006,N_7475);
and UO_873 (O_873,N_7369,N_6663);
or UO_874 (O_874,N_8273,N_5540);
and UO_875 (O_875,N_8104,N_6789);
nand UO_876 (O_876,N_9603,N_5916);
and UO_877 (O_877,N_7680,N_9830);
or UO_878 (O_878,N_9821,N_9747);
and UO_879 (O_879,N_6823,N_9609);
and UO_880 (O_880,N_5754,N_6601);
nand UO_881 (O_881,N_8053,N_9977);
nand UO_882 (O_882,N_8964,N_8706);
or UO_883 (O_883,N_6671,N_6907);
xor UO_884 (O_884,N_9961,N_6137);
nand UO_885 (O_885,N_9354,N_5743);
or UO_886 (O_886,N_6876,N_9297);
and UO_887 (O_887,N_8087,N_7560);
nor UO_888 (O_888,N_9288,N_8709);
nor UO_889 (O_889,N_7337,N_7053);
and UO_890 (O_890,N_5362,N_8839);
and UO_891 (O_891,N_6581,N_5539);
and UO_892 (O_892,N_7494,N_9791);
and UO_893 (O_893,N_9073,N_9846);
or UO_894 (O_894,N_9267,N_6291);
or UO_895 (O_895,N_5507,N_6167);
nand UO_896 (O_896,N_7608,N_7826);
and UO_897 (O_897,N_5167,N_7518);
and UO_898 (O_898,N_8573,N_9436);
and UO_899 (O_899,N_6196,N_8710);
nor UO_900 (O_900,N_8305,N_7691);
nor UO_901 (O_901,N_5991,N_5904);
nand UO_902 (O_902,N_7427,N_5786);
nor UO_903 (O_903,N_9767,N_5857);
xor UO_904 (O_904,N_9229,N_5398);
or UO_905 (O_905,N_8862,N_5079);
or UO_906 (O_906,N_7799,N_5109);
and UO_907 (O_907,N_9897,N_6277);
nor UO_908 (O_908,N_8992,N_5033);
or UO_909 (O_909,N_8791,N_7051);
nor UO_910 (O_910,N_5906,N_5797);
nand UO_911 (O_911,N_9358,N_9649);
nand UO_912 (O_912,N_7878,N_5439);
nand UO_913 (O_913,N_8959,N_6330);
nor UO_914 (O_914,N_8051,N_9773);
nor UO_915 (O_915,N_6774,N_5949);
nand UO_916 (O_916,N_9784,N_7723);
or UO_917 (O_917,N_9465,N_5594);
or UO_918 (O_918,N_8428,N_5040);
or UO_919 (O_919,N_6255,N_9800);
nand UO_920 (O_920,N_9233,N_7616);
or UO_921 (O_921,N_7261,N_5722);
nand UO_922 (O_922,N_8923,N_6960);
nor UO_923 (O_923,N_9589,N_9060);
or UO_924 (O_924,N_9679,N_5971);
and UO_925 (O_925,N_7654,N_5452);
nand UO_926 (O_926,N_8452,N_6326);
or UO_927 (O_927,N_9247,N_8636);
or UO_928 (O_928,N_5985,N_7352);
and UO_929 (O_929,N_6626,N_8750);
nand UO_930 (O_930,N_5686,N_8552);
nor UO_931 (O_931,N_7628,N_9433);
and UO_932 (O_932,N_8215,N_6345);
nand UO_933 (O_933,N_7901,N_5578);
and UO_934 (O_934,N_8641,N_6272);
and UO_935 (O_935,N_9208,N_8521);
and UO_936 (O_936,N_5150,N_9742);
and UO_937 (O_937,N_8367,N_6816);
and UO_938 (O_938,N_5412,N_8735);
xnor UO_939 (O_939,N_6923,N_7040);
or UO_940 (O_940,N_6961,N_9692);
or UO_941 (O_941,N_6640,N_7181);
or UO_942 (O_942,N_7662,N_5403);
nand UO_943 (O_943,N_6668,N_6331);
or UO_944 (O_944,N_5232,N_9983);
or UO_945 (O_945,N_7811,N_6356);
and UO_946 (O_946,N_9653,N_7357);
nand UO_947 (O_947,N_6436,N_9497);
nor UO_948 (O_948,N_8931,N_6534);
nand UO_949 (O_949,N_5895,N_7975);
and UO_950 (O_950,N_7372,N_8876);
and UO_951 (O_951,N_6132,N_8251);
and UO_952 (O_952,N_7558,N_5012);
nor UO_953 (O_953,N_8467,N_5137);
nand UO_954 (O_954,N_6397,N_7737);
and UO_955 (O_955,N_5599,N_9944);
or UO_956 (O_956,N_8147,N_7992);
and UO_957 (O_957,N_6104,N_8571);
or UO_958 (O_958,N_7153,N_9703);
and UO_959 (O_959,N_5226,N_9001);
nand UO_960 (O_960,N_9840,N_5954);
and UO_961 (O_961,N_7392,N_6573);
or UO_962 (O_962,N_7127,N_7538);
or UO_963 (O_963,N_7871,N_7304);
or UO_964 (O_964,N_6549,N_8029);
nand UO_965 (O_965,N_9626,N_7625);
and UO_966 (O_966,N_5840,N_7033);
nor UO_967 (O_967,N_6930,N_5613);
or UO_968 (O_968,N_8642,N_6247);
and UO_969 (O_969,N_8383,N_9640);
nor UO_970 (O_970,N_8980,N_6941);
nand UO_971 (O_971,N_5147,N_6509);
and UO_972 (O_972,N_7800,N_5953);
nand UO_973 (O_973,N_8447,N_6325);
nor UO_974 (O_974,N_5992,N_8228);
nand UO_975 (O_975,N_5491,N_6677);
nor UO_976 (O_976,N_8730,N_8821);
or UO_977 (O_977,N_9294,N_5498);
nor UO_978 (O_978,N_8043,N_8586);
or UO_979 (O_979,N_8024,N_9632);
and UO_980 (O_980,N_6432,N_6995);
and UO_981 (O_981,N_8067,N_8151);
nand UO_982 (O_982,N_8917,N_7536);
nor UO_983 (O_983,N_5772,N_5779);
and UO_984 (O_984,N_5662,N_9566);
nand UO_985 (O_985,N_7308,N_6478);
nand UO_986 (O_986,N_5649,N_7720);
nand UO_987 (O_987,N_9301,N_7137);
nand UO_988 (O_988,N_7816,N_8719);
nand UO_989 (O_989,N_6365,N_8243);
and UO_990 (O_990,N_7529,N_8323);
and UO_991 (O_991,N_7243,N_8130);
nor UO_992 (O_992,N_5685,N_6164);
nor UO_993 (O_993,N_6856,N_6915);
or UO_994 (O_994,N_9153,N_6461);
and UO_995 (O_995,N_5469,N_5668);
or UO_996 (O_996,N_5039,N_8815);
or UO_997 (O_997,N_7774,N_5304);
and UO_998 (O_998,N_8136,N_6740);
nor UO_999 (O_999,N_5657,N_8530);
nand UO_1000 (O_1000,N_6280,N_9483);
and UO_1001 (O_1001,N_7432,N_9764);
nand UO_1002 (O_1002,N_6620,N_8607);
and UO_1003 (O_1003,N_8512,N_6676);
nand UO_1004 (O_1004,N_7815,N_9770);
or UO_1005 (O_1005,N_7224,N_8012);
nand UO_1006 (O_1006,N_5347,N_9323);
or UO_1007 (O_1007,N_8771,N_7197);
nand UO_1008 (O_1008,N_7820,N_7239);
nor UO_1009 (O_1009,N_8794,N_9453);
nor UO_1010 (O_1010,N_5095,N_9228);
nand UO_1011 (O_1011,N_5281,N_9004);
nor UO_1012 (O_1012,N_5589,N_5443);
or UO_1013 (O_1013,N_9034,N_7404);
or UO_1014 (O_1014,N_5532,N_7171);
nor UO_1015 (O_1015,N_8991,N_6932);
or UO_1016 (O_1016,N_6457,N_6840);
or UO_1017 (O_1017,N_7270,N_8489);
and UO_1018 (O_1018,N_8698,N_8424);
nand UO_1019 (O_1019,N_6455,N_6496);
nor UO_1020 (O_1020,N_7908,N_8418);
and UO_1021 (O_1021,N_7091,N_9833);
nor UO_1022 (O_1022,N_7866,N_5785);
and UO_1023 (O_1023,N_7850,N_8025);
or UO_1024 (O_1024,N_9302,N_7734);
or UO_1025 (O_1025,N_5115,N_6008);
nand UO_1026 (O_1026,N_9375,N_6339);
and UO_1027 (O_1027,N_5348,N_8901);
or UO_1028 (O_1028,N_5634,N_7578);
and UO_1029 (O_1029,N_9242,N_7997);
nor UO_1030 (O_1030,N_8661,N_7493);
nand UO_1031 (O_1031,N_6014,N_7652);
or UO_1032 (O_1032,N_7448,N_7075);
nor UO_1033 (O_1033,N_6936,N_5205);
and UO_1034 (O_1034,N_6658,N_8061);
and UO_1035 (O_1035,N_6017,N_6103);
or UO_1036 (O_1036,N_7401,N_5848);
and UO_1037 (O_1037,N_6692,N_7702);
and UO_1038 (O_1038,N_9362,N_8776);
nand UO_1039 (O_1039,N_5959,N_6790);
and UO_1040 (O_1040,N_8685,N_6593);
nor UO_1041 (O_1041,N_8262,N_5527);
or UO_1042 (O_1042,N_9498,N_5990);
or UO_1043 (O_1043,N_8350,N_8986);
and UO_1044 (O_1044,N_8740,N_7567);
or UO_1045 (O_1045,N_5645,N_9669);
and UO_1046 (O_1046,N_7861,N_5413);
or UO_1047 (O_1047,N_5428,N_6110);
and UO_1048 (O_1048,N_9757,N_6688);
and UO_1049 (O_1049,N_9095,N_9326);
nor UO_1050 (O_1050,N_9915,N_7600);
and UO_1051 (O_1051,N_9959,N_7184);
nand UO_1052 (O_1052,N_8950,N_6536);
and UO_1053 (O_1053,N_6287,N_7735);
nor UO_1054 (O_1054,N_5395,N_9104);
and UO_1055 (O_1055,N_7327,N_5402);
or UO_1056 (O_1056,N_7713,N_7417);
or UO_1057 (O_1057,N_7835,N_6992);
nand UO_1058 (O_1058,N_9567,N_5200);
or UO_1059 (O_1059,N_9949,N_7473);
and UO_1060 (O_1060,N_5573,N_9914);
and UO_1061 (O_1061,N_6813,N_7697);
or UO_1062 (O_1062,N_6322,N_8360);
nand UO_1063 (O_1063,N_7751,N_5298);
nand UO_1064 (O_1064,N_5302,N_8425);
nor UO_1065 (O_1065,N_9622,N_6395);
nand UO_1066 (O_1066,N_7531,N_6882);
nor UO_1067 (O_1067,N_6165,N_5842);
and UO_1068 (O_1068,N_7295,N_6251);
nor UO_1069 (O_1069,N_9706,N_7719);
nand UO_1070 (O_1070,N_8680,N_7533);
nand UO_1071 (O_1071,N_9878,N_7164);
nand UO_1072 (O_1072,N_7970,N_8145);
nor UO_1073 (O_1073,N_5359,N_7336);
or UO_1074 (O_1074,N_7758,N_8589);
nand UO_1075 (O_1075,N_5445,N_8676);
nand UO_1076 (O_1076,N_7209,N_9712);
or UO_1077 (O_1077,N_5905,N_7037);
nand UO_1078 (O_1078,N_7785,N_5250);
or UO_1079 (O_1079,N_7370,N_6617);
and UO_1080 (O_1080,N_6548,N_9212);
and UO_1081 (O_1081,N_5926,N_7187);
or UO_1082 (O_1082,N_8150,N_9563);
nand UO_1083 (O_1083,N_9635,N_7817);
and UO_1084 (O_1084,N_5925,N_5998);
nor UO_1085 (O_1085,N_7801,N_6996);
nor UO_1086 (O_1086,N_6092,N_6401);
nand UO_1087 (O_1087,N_9636,N_7690);
and UO_1088 (O_1088,N_7152,N_9756);
nor UO_1089 (O_1089,N_6222,N_9625);
nand UO_1090 (O_1090,N_6656,N_5360);
or UO_1091 (O_1091,N_8160,N_9039);
xor UO_1092 (O_1092,N_8738,N_8800);
or UO_1093 (O_1093,N_8574,N_8174);
nand UO_1094 (O_1094,N_5790,N_7416);
or UO_1095 (O_1095,N_6724,N_9979);
and UO_1096 (O_1096,N_7246,N_8704);
nand UO_1097 (O_1097,N_6643,N_5056);
or UO_1098 (O_1098,N_6659,N_8040);
and UO_1099 (O_1099,N_8166,N_9911);
nand UO_1100 (O_1100,N_8763,N_8907);
or UO_1101 (O_1101,N_9966,N_8082);
nand UO_1102 (O_1102,N_5336,N_8793);
nand UO_1103 (O_1103,N_9038,N_8084);
or UO_1104 (O_1104,N_8107,N_9588);
nor UO_1105 (O_1105,N_5073,N_7505);
or UO_1106 (O_1106,N_9766,N_5951);
nand UO_1107 (O_1107,N_5561,N_9298);
or UO_1108 (O_1108,N_7622,N_7260);
and UO_1109 (O_1109,N_5286,N_6311);
nand UO_1110 (O_1110,N_8674,N_9967);
or UO_1111 (O_1111,N_6318,N_9245);
and UO_1112 (O_1112,N_7297,N_7103);
nor UO_1113 (O_1113,N_8375,N_8905);
and UO_1114 (O_1114,N_8754,N_9675);
or UO_1115 (O_1115,N_7725,N_6500);
and UO_1116 (O_1116,N_9068,N_9329);
nand UO_1117 (O_1117,N_5290,N_5521);
and UO_1118 (O_1118,N_6588,N_6898);
and UO_1119 (O_1119,N_7915,N_7408);
nor UO_1120 (O_1120,N_5628,N_6751);
nand UO_1121 (O_1121,N_9736,N_9584);
and UO_1122 (O_1122,N_9740,N_6293);
nand UO_1123 (O_1123,N_8581,N_7162);
nand UO_1124 (O_1124,N_6133,N_9831);
and UO_1125 (O_1125,N_5165,N_7658);
or UO_1126 (O_1126,N_9765,N_6243);
or UO_1127 (O_1127,N_5333,N_6874);
nor UO_1128 (O_1128,N_8369,N_8256);
nor UO_1129 (O_1129,N_6257,N_5203);
and UO_1130 (O_1130,N_6101,N_6234);
or UO_1131 (O_1131,N_9882,N_5808);
xnor UO_1132 (O_1132,N_7804,N_6317);
nor UO_1133 (O_1133,N_6906,N_7867);
nand UO_1134 (O_1134,N_8135,N_6649);
and UO_1135 (O_1135,N_8001,N_7320);
nand UO_1136 (O_1136,N_7433,N_9980);
nand UO_1137 (O_1137,N_6245,N_9802);
nand UO_1138 (O_1138,N_8034,N_8608);
or UO_1139 (O_1139,N_9901,N_7479);
nor UO_1140 (O_1140,N_9960,N_8963);
nor UO_1141 (O_1141,N_8088,N_7803);
and UO_1142 (O_1142,N_7098,N_8858);
nor UO_1143 (O_1143,N_5983,N_6136);
nand UO_1144 (O_1144,N_6193,N_5496);
nor UO_1145 (O_1145,N_6189,N_5803);
and UO_1146 (O_1146,N_9172,N_8920);
or UO_1147 (O_1147,N_5729,N_6139);
nor UO_1148 (O_1148,N_9528,N_5159);
or UO_1149 (O_1149,N_5664,N_5794);
nand UO_1150 (O_1150,N_8687,N_8492);
and UO_1151 (O_1151,N_7870,N_7514);
nor UO_1152 (O_1152,N_5227,N_6990);
nand UO_1153 (O_1153,N_6901,N_9350);
or UO_1154 (O_1154,N_5899,N_8547);
nand UO_1155 (O_1155,N_5720,N_8396);
xnor UO_1156 (O_1156,N_6614,N_8551);
and UO_1157 (O_1157,N_8783,N_7117);
nand UO_1158 (O_1158,N_7710,N_9399);
and UO_1159 (O_1159,N_5852,N_7281);
nor UO_1160 (O_1160,N_7165,N_7296);
or UO_1161 (O_1161,N_5696,N_6346);
nor UO_1162 (O_1162,N_9851,N_6263);
nor UO_1163 (O_1163,N_6703,N_6366);
and UO_1164 (O_1164,N_9615,N_8570);
or UO_1165 (O_1165,N_6686,N_7971);
nor UO_1166 (O_1166,N_6752,N_6056);
nand UO_1167 (O_1167,N_9779,N_7906);
nand UO_1168 (O_1168,N_6261,N_9863);
nor UO_1169 (O_1169,N_9473,N_8325);
or UO_1170 (O_1170,N_5106,N_8856);
and UO_1171 (O_1171,N_8855,N_8567);
and UO_1172 (O_1172,N_6489,N_5587);
nand UO_1173 (O_1173,N_7795,N_9782);
nor UO_1174 (O_1174,N_8753,N_6718);
and UO_1175 (O_1175,N_6225,N_6357);
nor UO_1176 (O_1176,N_7120,N_9531);
and UO_1177 (O_1177,N_8812,N_8507);
nand UO_1178 (O_1178,N_5913,N_5658);
and UO_1179 (O_1179,N_7096,N_9116);
nor UO_1180 (O_1180,N_8896,N_9051);
or UO_1181 (O_1181,N_5869,N_6199);
and UO_1182 (O_1182,N_9387,N_9359);
and UO_1183 (O_1183,N_9203,N_7353);
and UO_1184 (O_1184,N_6454,N_6540);
or UO_1185 (O_1185,N_5209,N_5179);
or UO_1186 (O_1186,N_9444,N_7643);
and UO_1187 (O_1187,N_6778,N_5472);
and UO_1188 (O_1188,N_8496,N_6916);
and UO_1189 (O_1189,N_8308,N_7102);
nor UO_1190 (O_1190,N_8420,N_7042);
and UO_1191 (O_1191,N_5859,N_6638);
and UO_1192 (O_1192,N_8882,N_9968);
nand UO_1193 (O_1193,N_7898,N_8989);
and UO_1194 (O_1194,N_8906,N_9629);
and UO_1195 (O_1195,N_6381,N_8798);
or UO_1196 (O_1196,N_6604,N_6569);
nor UO_1197 (O_1197,N_7143,N_8469);
nand UO_1198 (O_1198,N_5160,N_5310);
and UO_1199 (O_1199,N_7482,N_9137);
or UO_1200 (O_1200,N_6868,N_7631);
nor UO_1201 (O_1201,N_7455,N_7087);
nor UO_1202 (O_1202,N_6185,N_9047);
nor UO_1203 (O_1203,N_5314,N_6635);
nor UO_1204 (O_1204,N_5001,N_9728);
nor UO_1205 (O_1205,N_6788,N_7890);
and UO_1206 (O_1206,N_6191,N_9723);
or UO_1207 (O_1207,N_7128,N_6083);
nor UO_1208 (O_1208,N_6145,N_9704);
nor UO_1209 (O_1209,N_8113,N_9089);
nand UO_1210 (O_1210,N_7355,N_5543);
nand UO_1211 (O_1211,N_5191,N_9306);
or UO_1212 (O_1212,N_9429,N_8293);
or UO_1213 (O_1213,N_5011,N_7892);
nor UO_1214 (O_1214,N_8702,N_5134);
nand UO_1215 (O_1215,N_8566,N_8638);
and UO_1216 (O_1216,N_7105,N_9026);
or UO_1217 (O_1217,N_7770,N_9939);
or UO_1218 (O_1218,N_8079,N_8331);
nand UO_1219 (O_1219,N_6863,N_9231);
nand UO_1220 (O_1220,N_5885,N_6425);
nand UO_1221 (O_1221,N_8587,N_6163);
nand UO_1222 (O_1222,N_8132,N_9922);
or UO_1223 (O_1223,N_9702,N_9933);
or UO_1224 (O_1224,N_6474,N_7248);
nand UO_1225 (O_1225,N_5621,N_6612);
nor UO_1226 (O_1226,N_6400,N_6555);
or UO_1227 (O_1227,N_7447,N_9909);
nand UO_1228 (O_1228,N_6051,N_8445);
nor UO_1229 (O_1229,N_5969,N_9982);
and UO_1230 (O_1230,N_5337,N_7464);
or UO_1231 (O_1231,N_5004,N_9701);
or UO_1232 (O_1232,N_8869,N_9828);
and UO_1233 (O_1233,N_7678,N_5477);
nand UO_1234 (O_1234,N_8069,N_9746);
or UO_1235 (O_1235,N_9003,N_9568);
or UO_1236 (O_1236,N_7458,N_9232);
or UO_1237 (O_1237,N_5506,N_6129);
or UO_1238 (O_1238,N_5650,N_5101);
or UO_1239 (O_1239,N_7629,N_9050);
or UO_1240 (O_1240,N_8235,N_6362);
or UO_1241 (O_1241,N_6088,N_7132);
or UO_1242 (O_1242,N_9900,N_6583);
nor UO_1243 (O_1243,N_9741,N_6697);
nand UO_1244 (O_1244,N_7324,N_8689);
xnor UO_1245 (O_1245,N_6148,N_8720);
nor UO_1246 (O_1246,N_7856,N_6782);
nor UO_1247 (O_1247,N_6186,N_5018);
or UO_1248 (O_1248,N_9533,N_5393);
nor UO_1249 (O_1249,N_5228,N_8831);
nand UO_1250 (O_1250,N_8080,N_9076);
or UO_1251 (O_1251,N_9441,N_6580);
and UO_1252 (O_1252,N_9091,N_7667);
and UO_1253 (O_1253,N_5928,N_9319);
nor UO_1254 (O_1254,N_5111,N_9129);
nand UO_1255 (O_1255,N_7142,N_7396);
and UO_1256 (O_1256,N_5130,N_5986);
nor UO_1257 (O_1257,N_6741,N_9602);
nor UO_1258 (O_1258,N_8667,N_5919);
nor UO_1259 (O_1259,N_7764,N_7376);
nand UO_1260 (O_1260,N_5426,N_7314);
and UO_1261 (O_1261,N_6968,N_8505);
nor UO_1262 (O_1262,N_5810,N_6542);
nor UO_1263 (O_1263,N_5367,N_9439);
nor UO_1264 (O_1264,N_9873,N_6227);
nor UO_1265 (O_1265,N_6582,N_9181);
or UO_1266 (O_1266,N_6956,N_5690);
or UO_1267 (O_1267,N_9943,N_6016);
nand UO_1268 (O_1268,N_7621,N_5883);
nor UO_1269 (O_1269,N_9262,N_8739);
and UO_1270 (O_1270,N_8320,N_5880);
or UO_1271 (O_1271,N_7097,N_8058);
nand UO_1272 (O_1272,N_7348,N_7671);
nand UO_1273 (O_1273,N_9032,N_7259);
nand UO_1274 (O_1274,N_5867,N_5169);
nand UO_1275 (O_1275,N_6520,N_6859);
nor UO_1276 (O_1276,N_9056,N_9318);
and UO_1277 (O_1277,N_8357,N_5003);
nand UO_1278 (O_1278,N_5826,N_6682);
nor UO_1279 (O_1279,N_6354,N_8934);
nor UO_1280 (O_1280,N_6837,N_6226);
and UO_1281 (O_1281,N_5233,N_9667);
nand UO_1282 (O_1282,N_6140,N_8028);
nand UO_1283 (O_1283,N_5446,N_9860);
and UO_1284 (O_1284,N_6064,N_6624);
and UO_1285 (O_1285,N_7435,N_5958);
and UO_1286 (O_1286,N_9119,N_6421);
or UO_1287 (O_1287,N_5934,N_5423);
nor UO_1288 (O_1288,N_9719,N_6359);
or UO_1289 (O_1289,N_6796,N_6603);
nand UO_1290 (O_1290,N_9485,N_5815);
nor UO_1291 (O_1291,N_9451,N_7150);
nand UO_1292 (O_1292,N_6939,N_7580);
or UO_1293 (O_1293,N_5184,N_9642);
nand UO_1294 (O_1294,N_7587,N_5782);
nor UO_1295 (O_1295,N_6350,N_9500);
nor UO_1296 (O_1296,N_6375,N_8359);
or UO_1297 (O_1297,N_5083,N_8402);
or UO_1298 (O_1298,N_6131,N_5317);
or UO_1299 (O_1299,N_9182,N_6728);
nand UO_1300 (O_1300,N_5671,N_9735);
nand UO_1301 (O_1301,N_9265,N_9510);
or UO_1302 (O_1302,N_6810,N_5931);
or UO_1303 (O_1303,N_9870,N_9934);
or UO_1304 (O_1304,N_8845,N_8442);
and UO_1305 (O_1305,N_8167,N_9014);
or UO_1306 (O_1306,N_7728,N_5391);
or UO_1307 (O_1307,N_6224,N_8196);
nor UO_1308 (O_1308,N_5873,N_7852);
or UO_1309 (O_1309,N_8870,N_5812);
or UO_1310 (O_1310,N_8282,N_9133);
or UO_1311 (O_1311,N_7609,N_9699);
and UO_1312 (O_1312,N_7596,N_5289);
nor UO_1313 (O_1313,N_8615,N_9730);
or UO_1314 (O_1314,N_8630,N_8154);
and UO_1315 (O_1315,N_7293,N_8664);
and UO_1316 (O_1316,N_9351,N_8189);
nand UO_1317 (O_1317,N_8833,N_8354);
nand UO_1318 (O_1318,N_8807,N_7134);
nand UO_1319 (O_1319,N_9479,N_5297);
and UO_1320 (O_1320,N_9320,N_9495);
or UO_1321 (O_1321,N_6221,N_6817);
and UO_1322 (O_1322,N_6415,N_5608);
and UO_1323 (O_1323,N_5605,N_5022);
or UO_1324 (O_1324,N_9384,N_5973);
and UO_1325 (O_1325,N_8257,N_8184);
nand UO_1326 (O_1326,N_6347,N_5733);
or UO_1327 (O_1327,N_8314,N_9341);
and UO_1328 (O_1328,N_8755,N_8576);
nor UO_1329 (O_1329,N_6274,N_6279);
or UO_1330 (O_1330,N_7744,N_8650);
and UO_1331 (O_1331,N_7730,N_6254);
nand UO_1332 (O_1332,N_8951,N_8503);
and UO_1333 (O_1333,N_8622,N_9787);
and UO_1334 (O_1334,N_8066,N_9677);
and UO_1335 (O_1335,N_5541,N_5789);
nand UO_1336 (O_1336,N_8748,N_6590);
nor UO_1337 (O_1337,N_6675,N_8987);
or UO_1338 (O_1338,N_5087,N_6363);
nor UO_1339 (O_1339,N_7446,N_8398);
or UO_1340 (O_1340,N_9235,N_7023);
nor UO_1341 (O_1341,N_6493,N_9537);
nor UO_1342 (O_1342,N_6127,N_8285);
or UO_1343 (O_1343,N_9826,N_9027);
nor UO_1344 (O_1344,N_9391,N_9206);
and UO_1345 (O_1345,N_9086,N_9017);
nor UO_1346 (O_1346,N_6173,N_7763);
or UO_1347 (O_1347,N_6125,N_9369);
or UO_1348 (O_1348,N_7340,N_8250);
or UO_1349 (O_1349,N_6567,N_5094);
nand UO_1350 (O_1350,N_6732,N_8480);
and UO_1351 (O_1351,N_8483,N_9991);
nor UO_1352 (O_1352,N_6249,N_5174);
nand UO_1353 (O_1353,N_8697,N_5436);
or UO_1354 (O_1354,N_5611,N_6367);
nor UO_1355 (O_1355,N_9964,N_8018);
nor UO_1356 (O_1356,N_6905,N_9501);
or UO_1357 (O_1357,N_8466,N_9159);
and UO_1358 (O_1358,N_9420,N_6994);
and UO_1359 (O_1359,N_8436,N_7429);
nand UO_1360 (O_1360,N_5955,N_6079);
nor UO_1361 (O_1361,N_6952,N_9777);
nor UO_1362 (O_1362,N_7620,N_5021);
or UO_1363 (O_1363,N_7108,N_9373);
nor UO_1364 (O_1364,N_5765,N_7217);
nor UO_1365 (O_1365,N_8853,N_6304);
and UO_1366 (O_1366,N_6734,N_9455);
and UO_1367 (O_1367,N_8168,N_8965);
or UO_1368 (O_1368,N_8185,N_6699);
nand UO_1369 (O_1369,N_7694,N_6843);
nand UO_1370 (O_1370,N_8956,N_7206);
nor UO_1371 (O_1371,N_7557,N_9751);
and UO_1372 (O_1372,N_7905,N_9827);
nor UO_1373 (O_1373,N_9883,N_5856);
or UO_1374 (O_1374,N_8699,N_7020);
or UO_1375 (O_1375,N_7976,N_6093);
or UO_1376 (O_1376,N_6203,N_8606);
or UO_1377 (O_1377,N_8511,N_5141);
nand UO_1378 (O_1378,N_8624,N_9448);
or UO_1379 (O_1379,N_9803,N_9855);
or UO_1380 (O_1380,N_8042,N_8792);
nand UO_1381 (O_1381,N_6373,N_6594);
or UO_1382 (O_1382,N_8737,N_6938);
or UO_1383 (O_1383,N_7003,N_6892);
nand UO_1384 (O_1384,N_5043,N_7496);
or UO_1385 (O_1385,N_9136,N_5077);
nor UO_1386 (O_1386,N_6377,N_5623);
or UO_1387 (O_1387,N_5625,N_9395);
and UO_1388 (O_1388,N_8478,N_9780);
or UO_1389 (O_1389,N_5279,N_8400);
or UO_1390 (O_1390,N_7410,N_5093);
or UO_1391 (O_1391,N_8884,N_9633);
nor UO_1392 (O_1392,N_5677,N_6004);
or UO_1393 (O_1393,N_8663,N_6508);
and UO_1394 (O_1394,N_7853,N_6228);
or UO_1395 (O_1395,N_7095,N_7005);
and UO_1396 (O_1396,N_7974,N_7740);
and UO_1397 (O_1397,N_9425,N_7712);
and UO_1398 (O_1398,N_7172,N_7924);
nor UO_1399 (O_1399,N_9404,N_6099);
nor UO_1400 (O_1400,N_6528,N_7942);
nand UO_1401 (O_1401,N_8525,N_8341);
or UO_1402 (O_1402,N_9616,N_8949);
nor UO_1403 (O_1403,N_7502,N_6252);
nand UO_1404 (O_1404,N_9938,N_7356);
and UO_1405 (O_1405,N_8004,N_6873);
and UO_1406 (O_1406,N_5287,N_6611);
nand UO_1407 (O_1407,N_5494,N_5805);
xor UO_1408 (O_1408,N_8984,N_8995);
and UO_1409 (O_1409,N_8887,N_6899);
and UO_1410 (O_1410,N_6034,N_7423);
nand UO_1411 (O_1411,N_5700,N_8564);
nand UO_1412 (O_1412,N_5069,N_7922);
nor UO_1413 (O_1413,N_6177,N_7358);
or UO_1414 (O_1414,N_8899,N_6818);
nand UO_1415 (O_1415,N_7965,N_7638);
nor UO_1416 (O_1416,N_9907,N_5344);
nand UO_1417 (O_1417,N_5868,N_5881);
nand UO_1418 (O_1418,N_8562,N_7140);
nor UO_1419 (O_1419,N_8351,N_5669);
nand UO_1420 (O_1420,N_9396,N_9315);
nand UO_1421 (O_1421,N_6146,N_8172);
or UO_1422 (O_1422,N_9829,N_7753);
or UO_1423 (O_1423,N_8347,N_6382);
nand UO_1424 (O_1424,N_6270,N_9291);
nand UO_1425 (O_1425,N_6275,N_7797);
or UO_1426 (O_1426,N_7380,N_7014);
or UO_1427 (O_1427,N_7589,N_8218);
and UO_1428 (O_1428,N_7851,N_7920);
and UO_1429 (O_1429,N_6470,N_7309);
nand UO_1430 (O_1430,N_6701,N_6169);
nand UO_1431 (O_1431,N_7312,N_5761);
or UO_1432 (O_1432,N_6262,N_7255);
or UO_1433 (O_1433,N_8449,N_9110);
or UO_1434 (O_1434,N_5417,N_8137);
or UO_1435 (O_1435,N_9623,N_6429);
nand UO_1436 (O_1436,N_9973,N_8777);
or UO_1437 (O_1437,N_7718,N_6962);
and UO_1438 (O_1438,N_7834,N_5930);
and UO_1439 (O_1439,N_9557,N_6797);
nor UO_1440 (O_1440,N_8091,N_7129);
and UO_1441 (O_1441,N_7874,N_5909);
or UO_1442 (O_1442,N_6772,N_9413);
nor UO_1443 (O_1443,N_9850,N_7894);
and UO_1444 (O_1444,N_5741,N_7213);
nor UO_1445 (O_1445,N_9853,N_8463);
or UO_1446 (O_1446,N_9160,N_7946);
and UO_1447 (O_1447,N_7242,N_8732);
or UO_1448 (O_1448,N_9045,N_8128);
and UO_1449 (O_1449,N_9037,N_8877);
nand UO_1450 (O_1450,N_9727,N_5386);
xnor UO_1451 (O_1451,N_8487,N_6057);
and UO_1452 (O_1452,N_7160,N_9195);
nand UO_1453 (O_1453,N_9910,N_8940);
nor UO_1454 (O_1454,N_9438,N_5756);
nor UO_1455 (O_1455,N_6897,N_8816);
nand UO_1456 (O_1456,N_6070,N_8749);
nor UO_1457 (O_1457,N_9170,N_7798);
nand UO_1458 (O_1458,N_7027,N_5243);
nand UO_1459 (O_1459,N_6268,N_9268);
nand UO_1460 (O_1460,N_8633,N_5682);
nand UO_1461 (O_1461,N_7487,N_8045);
or UO_1462 (O_1462,N_7485,N_9346);
nand UO_1463 (O_1463,N_7081,N_6982);
and UO_1464 (O_1464,N_6212,N_6586);
or UO_1465 (O_1465,N_7028,N_7237);
and UO_1466 (O_1466,N_9094,N_7443);
or UO_1467 (O_1467,N_7873,N_9954);
nor UO_1468 (O_1468,N_9592,N_8426);
or UO_1469 (O_1469,N_5776,N_6340);
or UO_1470 (O_1470,N_5325,N_6879);
and UO_1471 (O_1471,N_5139,N_6119);
and UO_1472 (O_1472,N_8954,N_8401);
nor UO_1473 (O_1473,N_7689,N_6320);
or UO_1474 (O_1474,N_5701,N_7280);
and UO_1475 (O_1475,N_6691,N_5416);
or UO_1476 (O_1476,N_8430,N_5858);
and UO_1477 (O_1477,N_7660,N_9790);
nand UO_1478 (O_1478,N_5023,N_7450);
nand UO_1479 (O_1479,N_9681,N_6958);
nor UO_1480 (O_1480,N_8484,N_7236);
or UO_1481 (O_1481,N_6049,N_7809);
nor UO_1482 (O_1482,N_7636,N_5767);
or UO_1483 (O_1483,N_8081,N_5499);
nor UO_1484 (O_1484,N_7166,N_5831);
and UO_1485 (O_1485,N_7822,N_7056);
or UO_1486 (O_1486,N_9147,N_7049);
nor UO_1487 (O_1487,N_9107,N_7842);
or UO_1488 (O_1488,N_6753,N_7903);
or UO_1489 (O_1489,N_9305,N_7500);
or UO_1490 (O_1490,N_6444,N_9058);
nand UO_1491 (O_1491,N_8272,N_8580);
nand UO_1492 (O_1492,N_9946,N_6700);
nand UO_1493 (O_1493,N_8758,N_9529);
nand UO_1494 (O_1494,N_7441,N_9599);
nor UO_1495 (O_1495,N_9207,N_7067);
and UO_1496 (O_1496,N_9093,N_8646);
or UO_1497 (O_1497,N_9739,N_9894);
nor UO_1498 (O_1498,N_6188,N_6204);
nand UO_1499 (O_1499,N_8017,N_9889);
endmodule