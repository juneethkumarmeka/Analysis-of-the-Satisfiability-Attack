module basic_1500_15000_2000_120_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_689,In_1426);
xnor U1 (N_1,In_475,In_41);
nor U2 (N_2,In_1428,In_1137);
nand U3 (N_3,In_1100,In_1129);
nand U4 (N_4,In_488,In_1212);
nand U5 (N_5,In_214,In_1051);
nand U6 (N_6,In_1374,In_880);
or U7 (N_7,In_96,In_1024);
and U8 (N_8,In_504,In_1148);
or U9 (N_9,In_857,In_805);
or U10 (N_10,In_1081,In_1273);
xnor U11 (N_11,In_236,In_453);
or U12 (N_12,In_86,In_381);
xnor U13 (N_13,In_1074,In_1206);
and U14 (N_14,In_121,In_279);
and U15 (N_15,In_1142,In_94);
and U16 (N_16,In_1236,In_319);
or U17 (N_17,In_1485,In_1494);
or U18 (N_18,In_545,In_202);
nor U19 (N_19,In_1497,In_476);
nand U20 (N_20,In_1203,In_1420);
xor U21 (N_21,In_1272,In_392);
nand U22 (N_22,In_996,In_1076);
nor U23 (N_23,In_553,In_1477);
and U24 (N_24,In_410,In_1361);
and U25 (N_25,In_985,In_704);
or U26 (N_26,In_1136,In_181);
xor U27 (N_27,In_1063,In_558);
nand U28 (N_28,In_934,In_728);
or U29 (N_29,In_444,In_1390);
or U30 (N_30,In_574,In_598);
nand U31 (N_31,In_217,In_235);
nand U32 (N_32,In_1198,In_14);
xor U33 (N_33,In_867,In_419);
or U34 (N_34,In_1437,In_1407);
and U35 (N_35,In_1289,In_834);
xor U36 (N_36,In_532,In_820);
or U37 (N_37,In_683,In_1143);
nor U38 (N_38,In_599,In_995);
nand U39 (N_39,In_1095,In_53);
and U40 (N_40,In_1466,In_988);
xor U41 (N_41,In_597,In_215);
xnor U42 (N_42,In_112,In_1128);
nand U43 (N_43,In_1171,In_42);
and U44 (N_44,In_485,In_740);
nor U45 (N_45,In_354,In_6);
nand U46 (N_46,In_974,In_631);
xor U47 (N_47,In_288,In_840);
nand U48 (N_48,In_695,In_729);
nor U49 (N_49,In_682,In_1144);
and U50 (N_50,In_941,In_625);
nand U51 (N_51,In_477,In_958);
and U52 (N_52,In_1090,In_1164);
or U53 (N_53,In_1228,In_1082);
nor U54 (N_54,In_464,In_1282);
and U55 (N_55,In_752,In_1257);
nand U56 (N_56,In_1232,In_1154);
or U57 (N_57,In_1334,In_1472);
and U58 (N_58,In_69,In_253);
xnor U59 (N_59,In_1481,In_844);
and U60 (N_60,In_736,In_314);
and U61 (N_61,In_1209,In_637);
or U62 (N_62,In_1172,In_1107);
nand U63 (N_63,In_1329,In_302);
or U64 (N_64,In_82,In_753);
nor U65 (N_65,In_808,In_676);
and U66 (N_66,In_339,In_956);
nor U67 (N_67,In_1155,In_1127);
or U68 (N_68,In_299,In_940);
nor U69 (N_69,In_539,In_493);
or U70 (N_70,In_1303,In_427);
and U71 (N_71,In_648,In_911);
xnor U72 (N_72,In_118,In_228);
or U73 (N_73,In_107,In_706);
xnor U74 (N_74,In_807,In_409);
nor U75 (N_75,In_1071,In_1386);
or U76 (N_76,In_1445,In_333);
nor U77 (N_77,In_126,In_1185);
xnor U78 (N_78,In_977,In_1021);
nand U79 (N_79,In_458,In_639);
and U80 (N_80,In_700,In_904);
or U81 (N_81,In_611,In_165);
or U82 (N_82,In_1369,In_201);
and U83 (N_83,In_1193,In_1299);
and U84 (N_84,In_106,In_1371);
nand U85 (N_85,In_984,In_1068);
and U86 (N_86,In_883,In_2);
nor U87 (N_87,In_735,In_848);
nor U88 (N_88,In_937,In_1380);
nand U89 (N_89,In_803,In_30);
and U90 (N_90,In_1139,In_167);
nand U91 (N_91,In_876,In_242);
nand U92 (N_92,In_1367,In_932);
xnor U93 (N_93,In_953,In_1269);
and U94 (N_94,In_1318,In_500);
nand U95 (N_95,In_12,In_635);
and U96 (N_96,In_100,In_1383);
nor U97 (N_97,In_566,In_11);
nand U98 (N_98,In_318,In_46);
or U99 (N_99,In_76,In_793);
nor U100 (N_100,In_962,In_744);
and U101 (N_101,In_1032,In_713);
xor U102 (N_102,In_408,In_200);
or U103 (N_103,In_285,In_1001);
nor U104 (N_104,In_1457,In_1266);
xnor U105 (N_105,In_1216,In_21);
or U106 (N_106,In_542,In_709);
nor U107 (N_107,In_74,In_1311);
or U108 (N_108,In_62,In_415);
xor U109 (N_109,In_1247,In_1087);
xor U110 (N_110,In_1031,In_523);
or U111 (N_111,In_32,In_733);
nand U112 (N_112,In_468,In_534);
nand U113 (N_113,In_1058,In_417);
nor U114 (N_114,In_677,In_1158);
and U115 (N_115,In_134,In_1274);
nand U116 (N_116,In_60,In_1204);
or U117 (N_117,In_222,In_473);
and U118 (N_118,In_1341,In_927);
or U119 (N_119,In_268,In_612);
or U120 (N_120,In_124,In_555);
nor U121 (N_121,In_1450,In_1438);
nand U122 (N_122,In_496,In_1121);
or U123 (N_123,In_638,In_1306);
nor U124 (N_124,In_860,In_331);
and U125 (N_125,In_1381,In_745);
nor U126 (N_126,N_55,In_686);
nor U127 (N_127,In_84,In_697);
or U128 (N_128,In_194,In_1478);
and U129 (N_129,In_1053,In_852);
nand U130 (N_130,In_673,In_864);
nor U131 (N_131,In_1243,In_1059);
xor U132 (N_132,In_636,In_190);
xnor U133 (N_133,In_1008,In_168);
xor U134 (N_134,In_845,In_366);
or U135 (N_135,In_916,In_1217);
nand U136 (N_136,N_107,In_1084);
or U137 (N_137,In_522,In_157);
or U138 (N_138,In_981,In_872);
xnor U139 (N_139,In_284,In_721);
and U140 (N_140,In_499,In_1416);
or U141 (N_141,In_92,In_795);
nand U142 (N_142,In_655,In_554);
nand U143 (N_143,In_884,In_544);
nand U144 (N_144,In_921,In_1234);
nand U145 (N_145,In_494,In_1349);
nand U146 (N_146,In_247,In_1332);
or U147 (N_147,In_780,In_505);
xnor U148 (N_148,In_293,In_972);
xnor U149 (N_149,In_128,In_1249);
nand U150 (N_150,In_1330,In_584);
nor U151 (N_151,In_1186,In_1250);
xnor U152 (N_152,N_30,In_212);
nand U153 (N_153,In_698,In_186);
and U154 (N_154,In_1006,In_1468);
nand U155 (N_155,In_1321,In_231);
and U156 (N_156,In_1169,In_358);
xor U157 (N_157,In_258,In_547);
nand U158 (N_158,In_125,In_731);
or U159 (N_159,In_1030,In_1037);
and U160 (N_160,In_540,In_188);
or U161 (N_161,In_561,In_1434);
xnor U162 (N_162,In_798,In_1218);
and U163 (N_163,In_1175,N_67);
nor U164 (N_164,In_1072,In_371);
or U165 (N_165,In_317,In_789);
nand U166 (N_166,In_1098,In_315);
xor U167 (N_167,In_609,N_97);
xnor U168 (N_168,In_394,In_758);
nor U169 (N_169,In_466,N_75);
xor U170 (N_170,In_295,N_99);
nand U171 (N_171,In_831,In_1079);
or U172 (N_172,N_4,In_537);
or U173 (N_173,N_21,In_1356);
nor U174 (N_174,In_647,In_311);
and U175 (N_175,In_1404,In_640);
nor U176 (N_176,N_53,In_777);
nor U177 (N_177,In_1056,In_913);
nand U178 (N_178,In_31,In_1373);
or U179 (N_179,In_684,In_862);
xnor U180 (N_180,In_632,In_237);
xor U181 (N_181,N_84,In_122);
nand U182 (N_182,In_260,In_1446);
and U183 (N_183,In_306,In_1038);
nand U184 (N_184,In_206,In_634);
or U185 (N_185,In_440,In_197);
and U186 (N_186,In_1042,In_738);
nand U187 (N_187,In_869,In_300);
or U188 (N_188,In_1255,In_1132);
or U189 (N_189,N_69,In_910);
or U190 (N_190,In_57,In_658);
xor U191 (N_191,In_1043,N_6);
and U192 (N_192,In_665,In_1421);
xnor U193 (N_193,In_1425,In_716);
xnor U194 (N_194,In_406,In_450);
nand U195 (N_195,In_359,In_671);
or U196 (N_196,In_379,In_172);
and U197 (N_197,In_340,In_887);
and U198 (N_198,In_601,In_866);
nor U199 (N_199,In_560,In_1474);
or U200 (N_200,In_816,In_1115);
nor U201 (N_201,In_322,In_383);
nor U202 (N_202,In_743,In_363);
nand U203 (N_203,In_1458,In_707);
and U204 (N_204,N_113,In_297);
xnor U205 (N_205,In_1123,In_1368);
nor U206 (N_206,In_570,In_589);
or U207 (N_207,In_1133,In_770);
nand U208 (N_208,In_449,In_567);
and U209 (N_209,In_1202,In_1167);
nor U210 (N_210,In_309,In_492);
or U211 (N_211,N_124,N_14);
and U212 (N_212,In_1331,In_273);
or U213 (N_213,In_180,In_606);
nand U214 (N_214,In_1151,In_275);
nand U215 (N_215,In_259,In_936);
and U216 (N_216,In_813,In_1233);
xor U217 (N_217,In_859,In_33);
nand U218 (N_218,In_1376,In_1360);
nor U219 (N_219,N_43,In_502);
or U220 (N_220,In_70,In_990);
nor U221 (N_221,In_833,In_442);
xnor U222 (N_222,In_143,In_952);
xor U223 (N_223,In_694,In_1414);
or U224 (N_224,In_1138,In_1382);
or U225 (N_225,In_797,In_216);
or U226 (N_226,In_1280,In_755);
nand U227 (N_227,In_1141,In_1353);
nand U228 (N_228,In_454,In_1323);
and U229 (N_229,In_471,In_1065);
or U230 (N_230,In_1105,In_1170);
or U231 (N_231,In_189,In_1027);
nor U232 (N_232,In_1075,In_252);
xnor U233 (N_233,In_65,In_68);
xor U234 (N_234,In_16,In_1213);
or U235 (N_235,In_696,In_865);
or U236 (N_236,In_938,In_0);
or U237 (N_237,In_199,In_1372);
xnor U238 (N_238,In_1184,N_52);
xnor U239 (N_239,In_1176,In_316);
nor U240 (N_240,In_681,In_593);
and U241 (N_241,In_210,In_142);
or U242 (N_242,In_262,In_432);
or U243 (N_243,In_1099,In_619);
and U244 (N_244,In_835,In_338);
or U245 (N_245,In_823,N_102);
nor U246 (N_246,In_341,In_480);
nand U247 (N_247,In_1224,In_902);
and U248 (N_248,In_1417,In_991);
xor U249 (N_249,In_583,In_747);
nand U250 (N_250,In_588,In_1482);
nor U251 (N_251,In_343,N_195);
nor U252 (N_252,In_263,In_151);
and U253 (N_253,In_1124,In_919);
xnor U254 (N_254,In_668,N_90);
nor U255 (N_255,In_360,In_1480);
nand U256 (N_256,In_970,In_899);
and U257 (N_257,N_188,In_512);
xnor U258 (N_258,In_535,In_39);
xor U259 (N_259,In_832,In_158);
nand U260 (N_260,In_1431,In_49);
nor U261 (N_261,In_827,In_355);
or U262 (N_262,N_37,In_772);
nand U263 (N_263,In_1254,In_1487);
nor U264 (N_264,N_219,In_95);
xnor U265 (N_265,N_20,N_33);
xor U266 (N_266,In_771,N_111);
nand U267 (N_267,In_1118,In_248);
nor U268 (N_268,N_222,In_400);
and U269 (N_269,In_531,In_621);
nand U270 (N_270,In_1069,In_594);
xor U271 (N_271,In_907,In_871);
and U272 (N_272,In_1149,In_1239);
nor U273 (N_273,In_855,In_490);
nor U274 (N_274,In_817,In_1322);
and U275 (N_275,In_1454,In_939);
and U276 (N_276,In_822,In_1028);
nor U277 (N_277,In_895,In_244);
or U278 (N_278,In_1263,In_660);
and U279 (N_279,N_128,In_727);
nor U280 (N_280,In_949,In_1180);
xor U281 (N_281,In_965,In_1242);
and U282 (N_282,In_659,In_1489);
and U283 (N_283,In_378,N_198);
xor U284 (N_284,In_1086,N_39);
and U285 (N_285,N_205,In_1003);
or U286 (N_286,In_397,In_85);
nor U287 (N_287,In_83,In_1000);
nand U288 (N_288,N_155,In_418);
or U289 (N_289,N_105,N_239);
nand U290 (N_290,In_28,N_25);
and U291 (N_291,In_1357,N_62);
or U292 (N_292,N_59,In_218);
and U293 (N_293,In_420,In_508);
nand U294 (N_294,In_1117,In_1040);
xor U295 (N_295,N_112,N_127);
nand U296 (N_296,In_428,In_596);
and U297 (N_297,N_44,In_1347);
and U298 (N_298,In_873,In_1490);
nor U299 (N_299,In_352,In_875);
xnor U300 (N_300,In_749,In_918);
and U301 (N_301,N_158,In_801);
xor U302 (N_302,In_88,In_1456);
or U303 (N_303,In_1275,In_344);
or U304 (N_304,In_1286,In_1297);
nand U305 (N_305,In_127,In_511);
nand U306 (N_306,In_162,In_87);
or U307 (N_307,In_1302,N_88);
nor U308 (N_308,In_1486,In_1049);
xor U309 (N_309,In_585,In_1348);
nand U310 (N_310,In_811,In_931);
nor U311 (N_311,In_791,N_165);
nand U312 (N_312,In_482,In_1078);
or U313 (N_313,N_51,N_79);
nand U314 (N_314,In_230,In_830);
nor U315 (N_315,In_888,N_130);
or U316 (N_316,In_396,In_1295);
nor U317 (N_317,In_467,In_896);
nand U318 (N_318,In_43,N_78);
nand U319 (N_319,In_1358,In_1150);
nand U320 (N_320,N_96,In_135);
nor U321 (N_321,In_232,In_56);
nor U322 (N_322,In_221,In_1448);
and U323 (N_323,N_206,In_1062);
or U324 (N_324,In_211,In_399);
or U325 (N_325,In_781,In_481);
or U326 (N_326,In_99,In_348);
xnor U327 (N_327,In_462,In_101);
and U328 (N_328,In_524,In_507);
xnor U329 (N_329,In_1182,In_1061);
and U330 (N_330,In_486,N_180);
and U331 (N_331,In_117,In_1012);
or U332 (N_332,In_1325,In_298);
nand U333 (N_333,N_136,In_997);
xor U334 (N_334,In_224,In_174);
nor U335 (N_335,In_975,In_78);
xor U336 (N_336,In_863,In_576);
xor U337 (N_337,In_75,N_215);
and U338 (N_338,N_81,In_964);
and U339 (N_339,N_230,In_1377);
nor U340 (N_340,In_384,In_769);
and U341 (N_341,In_900,In_54);
nor U342 (N_342,In_679,N_213);
or U343 (N_343,In_1315,N_82);
nor U344 (N_344,In_569,In_1310);
or U345 (N_345,N_154,In_739);
and U346 (N_346,In_963,In_821);
xnor U347 (N_347,In_802,N_31);
nand U348 (N_348,In_1187,In_768);
or U349 (N_349,In_1467,N_172);
nor U350 (N_350,N_173,In_715);
and U351 (N_351,In_579,In_1134);
and U352 (N_352,In_592,N_70);
and U353 (N_353,In_691,N_116);
nand U354 (N_354,N_243,In_336);
nor U355 (N_355,In_1146,In_944);
nor U356 (N_356,In_103,In_116);
and U357 (N_357,In_20,In_7);
or U358 (N_358,In_765,In_1298);
xnor U359 (N_359,In_1409,In_66);
or U360 (N_360,N_248,In_690);
or U361 (N_361,In_1,In_732);
nand U362 (N_362,In_550,In_565);
and U363 (N_363,N_183,In_1166);
nor U364 (N_364,In_1014,In_849);
or U365 (N_365,In_1344,In_675);
nand U366 (N_366,In_431,In_1461);
xor U367 (N_367,N_196,N_22);
nor U368 (N_368,In_1122,N_151);
nor U369 (N_369,In_1433,In_784);
nor U370 (N_370,In_47,N_143);
xor U371 (N_371,In_1160,In_1097);
nor U372 (N_372,In_1392,In_650);
or U373 (N_373,In_767,In_1109);
xor U374 (N_374,In_1196,In_404);
nor U375 (N_375,In_1080,N_123);
and U376 (N_376,In_856,N_171);
nand U377 (N_377,In_717,N_18);
or U378 (N_378,N_131,In_72);
xor U379 (N_379,In_685,In_1221);
and U380 (N_380,In_1294,In_234);
xor U381 (N_381,In_495,In_1214);
or U382 (N_382,In_163,N_161);
and U383 (N_383,In_653,In_711);
xnor U384 (N_384,In_1002,In_474);
or U385 (N_385,In_332,N_74);
xnor U386 (N_386,In_133,N_0);
nor U387 (N_387,N_114,In_552);
xor U388 (N_388,In_153,In_1034);
nand U389 (N_389,N_344,N_323);
and U390 (N_390,N_32,In_1220);
nand U391 (N_391,In_367,In_421);
or U392 (N_392,In_350,In_1211);
nor U393 (N_393,In_1248,N_200);
and U394 (N_394,N_264,In_90);
xnor U395 (N_395,N_324,N_42);
nand U396 (N_396,In_829,In_385);
or U397 (N_397,In_825,In_645);
nand U398 (N_398,N_119,In_933);
and U399 (N_399,In_388,In_750);
nor U400 (N_400,In_1492,In_714);
xnor U401 (N_401,N_108,In_1244);
nand U402 (N_402,In_1406,N_246);
or U403 (N_403,In_577,In_882);
nand U404 (N_404,In_254,N_89);
nand U405 (N_405,In_980,In_10);
or U406 (N_406,N_301,N_289);
nor U407 (N_407,In_447,In_943);
xor U408 (N_408,In_761,In_155);
and U409 (N_409,In_23,In_722);
nand U410 (N_410,In_559,In_386);
nand U411 (N_411,In_1119,In_169);
nor U412 (N_412,N_327,N_259);
or U413 (N_413,In_948,In_1443);
nand U414 (N_414,In_469,In_1333);
nor U415 (N_415,In_131,In_548);
nor U416 (N_416,In_950,N_201);
and U417 (N_417,In_171,N_365);
and U418 (N_418,N_252,In_868);
nand U419 (N_419,In_1283,N_247);
xnor U420 (N_420,N_340,In_204);
or U421 (N_421,In_1055,In_81);
and U422 (N_422,N_322,In_1422);
nor U423 (N_423,N_266,In_1064);
and U424 (N_424,In_776,In_573);
nor U425 (N_425,In_1066,In_144);
or U426 (N_426,In_1432,N_285);
or U427 (N_427,In_986,N_193);
and U428 (N_428,In_838,In_656);
or U429 (N_429,In_170,In_307);
nor U430 (N_430,N_314,In_207);
or U431 (N_431,In_925,In_347);
or U432 (N_432,In_277,N_15);
and U433 (N_433,In_265,In_1285);
and U434 (N_434,In_1041,N_313);
and U435 (N_435,In_756,N_118);
or U436 (N_436,N_85,In_898);
or U437 (N_437,In_966,In_819);
nand U438 (N_438,In_430,In_957);
and U439 (N_439,In_413,In_1340);
or U440 (N_440,In_61,In_372);
and U441 (N_441,N_91,N_374);
nor U442 (N_442,In_1178,N_342);
and U443 (N_443,In_152,In_292);
and U444 (N_444,In_1145,In_98);
nor U445 (N_445,N_140,N_287);
nor U446 (N_446,N_16,N_66);
nor U447 (N_447,In_543,In_794);
nor U448 (N_448,In_1324,In_894);
nand U449 (N_449,In_917,In_853);
nor U450 (N_450,In_267,In_556);
nor U451 (N_451,In_536,N_227);
or U452 (N_452,In_666,In_1108);
nand U453 (N_453,In_983,In_533);
and U454 (N_454,In_368,In_498);
and U455 (N_455,N_186,N_117);
xnor U456 (N_456,In_1256,N_260);
and U457 (N_457,In_281,In_1036);
xor U458 (N_458,N_192,N_346);
xnor U459 (N_459,In_692,N_7);
or U460 (N_460,In_1309,In_55);
or U461 (N_461,In_402,N_178);
and U462 (N_462,N_351,N_255);
or U463 (N_463,N_129,In_818);
nand U464 (N_464,In_1215,In_375);
nand U465 (N_465,In_562,In_1190);
nor U466 (N_466,N_292,In_479);
nand U467 (N_467,N_241,In_1103);
xor U468 (N_468,In_568,In_1316);
nor U469 (N_469,N_363,In_602);
nand U470 (N_470,In_1473,In_433);
nor U471 (N_471,In_1252,In_1307);
xnor U472 (N_472,In_538,In_403);
nand U473 (N_473,In_1230,N_373);
xor U474 (N_474,In_414,In_1201);
and U475 (N_475,In_1265,N_214);
nor U476 (N_476,N_278,In_1395);
or U477 (N_477,N_1,N_325);
or U478 (N_478,In_423,N_304);
xor U479 (N_479,N_13,In_195);
nor U480 (N_480,In_1157,N_353);
nor U481 (N_481,In_179,In_874);
nand U482 (N_482,In_487,N_208);
nand U483 (N_483,N_203,N_318);
and U484 (N_484,In_654,In_519);
or U485 (N_485,In_901,In_1131);
or U486 (N_486,N_156,N_83);
and U487 (N_487,N_279,In_580);
nor U488 (N_488,In_264,In_1054);
or U489 (N_489,In_335,In_1436);
nor U490 (N_490,In_97,In_775);
and U491 (N_491,In_398,In_241);
or U492 (N_492,In_115,In_1181);
or U493 (N_493,In_506,N_212);
or U494 (N_494,N_5,In_59);
xnor U495 (N_495,In_1270,In_1271);
nand U496 (N_496,In_1379,In_858);
nor U497 (N_497,In_699,In_1005);
or U498 (N_498,In_994,In_1092);
nor U499 (N_499,N_293,In_930);
xnor U500 (N_500,N_399,In_667);
nand U501 (N_501,In_227,N_277);
or U502 (N_502,N_375,N_435);
nand U503 (N_503,N_209,In_642);
and U504 (N_504,In_976,N_362);
nand U505 (N_505,N_453,N_468);
or U506 (N_506,In_1083,In_971);
nor U507 (N_507,N_450,In_63);
or U508 (N_508,In_1385,In_52);
nand U509 (N_509,In_1339,In_193);
and U510 (N_510,In_164,In_1396);
xnor U511 (N_511,N_480,In_1007);
xor U512 (N_512,In_233,N_150);
nor U513 (N_513,N_276,N_334);
or U514 (N_514,N_149,In_551);
and U515 (N_515,In_670,N_290);
xor U516 (N_516,In_708,N_372);
nor U517 (N_517,In_296,In_847);
nand U518 (N_518,In_942,N_109);
nand U519 (N_519,In_510,In_730);
nand U520 (N_520,In_1449,In_278);
xor U521 (N_521,N_319,In_877);
or U522 (N_522,In_1281,In_1479);
nand U523 (N_523,N_234,In_286);
or U524 (N_524,In_71,In_51);
or U525 (N_525,In_979,In_356);
nor U526 (N_526,N_226,In_1192);
nor U527 (N_527,In_80,N_386);
nor U528 (N_528,N_103,N_9);
xor U529 (N_529,In_622,N_412);
nor U530 (N_530,In_1238,In_973);
nor U531 (N_531,N_302,N_282);
nor U532 (N_532,In_34,N_47);
nand U533 (N_533,N_497,N_121);
nor U534 (N_534,In_1018,In_1469);
nand U535 (N_535,N_288,In_615);
or U536 (N_536,N_384,In_1498);
nand U537 (N_537,N_433,In_77);
and U538 (N_538,In_790,In_1067);
and U539 (N_539,N_432,In_489);
nand U540 (N_540,N_8,In_703);
and U541 (N_541,N_484,N_461);
or U542 (N_542,N_58,N_482);
nor U543 (N_543,In_513,In_1114);
xor U544 (N_544,N_441,N_400);
nor U545 (N_545,N_354,In_1011);
xnor U546 (N_546,N_194,N_50);
or U547 (N_547,In_1262,In_678);
nand U548 (N_548,In_851,In_617);
or U549 (N_549,N_225,N_191);
or U550 (N_550,N_499,In_1231);
and U551 (N_551,In_35,In_712);
nand U552 (N_552,N_257,N_309);
nor U553 (N_553,In_662,In_1241);
or U554 (N_554,N_444,In_203);
nand U555 (N_555,N_472,In_1288);
xor U556 (N_556,In_718,In_438);
xor U557 (N_557,In_792,In_3);
or U558 (N_558,N_368,N_364);
nand U559 (N_559,In_395,N_125);
and U560 (N_560,N_162,In_719);
nor U561 (N_561,N_216,N_406);
xnor U562 (N_562,In_1089,N_232);
xnor U563 (N_563,N_197,In_187);
xnor U564 (N_564,In_903,In_196);
nand U565 (N_565,N_281,In_842);
and U566 (N_566,In_701,N_133);
and U567 (N_567,In_503,In_357);
and U568 (N_568,N_139,In_1130);
nor U569 (N_569,N_95,In_437);
nor U570 (N_570,N_296,N_249);
or U571 (N_571,In_251,In_626);
and U572 (N_572,In_720,N_455);
xnor U573 (N_573,In_680,In_1268);
and U574 (N_574,In_1491,In_1337);
xnor U575 (N_575,In_628,In_779);
nand U576 (N_576,In_608,N_12);
or U577 (N_577,In_274,In_1447);
nor U578 (N_578,In_1405,In_881);
and U579 (N_579,In_1441,In_1227);
or U580 (N_580,In_1401,N_28);
or U581 (N_581,In_1493,N_258);
nand U582 (N_582,In_1398,In_614);
or U583 (N_583,In_15,In_890);
xnor U584 (N_584,In_1033,N_310);
nand U585 (N_585,In_44,N_475);
xor U586 (N_586,In_294,In_644);
and U587 (N_587,In_337,N_380);
xnor U588 (N_588,In_726,N_54);
xnor U589 (N_589,N_462,In_603);
or U590 (N_590,In_405,In_1484);
or U591 (N_591,In_1363,In_604);
xnor U592 (N_592,In_213,In_1319);
nor U593 (N_593,In_530,N_348);
and U594 (N_594,In_1174,In_1152);
nand U595 (N_595,In_452,In_1125);
nor U596 (N_596,N_371,In_361);
nand U597 (N_597,In_497,N_253);
or U598 (N_598,In_26,N_40);
and U599 (N_599,N_27,In_37);
nand U600 (N_600,In_796,N_355);
nor U601 (N_601,In_17,In_150);
nand U602 (N_602,In_786,N_80);
nor U603 (N_603,In_351,N_77);
nor U604 (N_604,N_35,N_397);
nor U605 (N_605,In_891,In_19);
or U606 (N_606,N_361,In_1260);
xor U607 (N_607,In_435,In_1016);
or U608 (N_608,In_1229,In_1430);
and U609 (N_609,N_312,In_191);
or U610 (N_610,N_166,In_549);
xnor U611 (N_611,In_514,In_1153);
nand U612 (N_612,N_284,In_1060);
nor U613 (N_613,N_379,In_657);
or U614 (N_614,N_187,In_1293);
or U615 (N_615,In_841,In_861);
nor U616 (N_616,In_893,In_369);
nor U617 (N_617,N_470,In_1342);
and U618 (N_618,N_298,In_1384);
nand U619 (N_619,In_380,In_48);
xnor U620 (N_620,In_1223,In_303);
nand U621 (N_621,In_401,N_48);
or U622 (N_622,In_947,N_147);
or U623 (N_623,In_240,N_291);
nor U624 (N_624,In_605,N_465);
xor U625 (N_625,In_1345,In_1397);
nor U626 (N_626,In_426,N_500);
or U627 (N_627,N_541,N_545);
nand U628 (N_628,In_1017,N_396);
xor U629 (N_629,N_256,In_773);
or U630 (N_630,N_377,In_1442);
and U631 (N_631,N_538,In_1427);
nand U632 (N_632,In_136,In_1471);
nor U633 (N_633,In_998,In_664);
nor U634 (N_634,N_330,N_320);
and U635 (N_635,In_929,In_581);
nor U636 (N_636,In_50,N_87);
nand U637 (N_637,N_544,In_478);
xnor U638 (N_638,In_1101,In_1410);
nand U639 (N_639,N_570,N_185);
xnor U640 (N_640,N_563,In_205);
nand U641 (N_641,N_617,In_1177);
xnor U642 (N_642,N_576,In_1423);
nor U643 (N_643,N_469,N_182);
or U644 (N_644,In_897,N_168);
nand U645 (N_645,N_588,In_516);
and U646 (N_646,In_219,N_495);
and U647 (N_647,In_463,N_283);
nand U648 (N_648,In_220,In_460);
or U649 (N_649,N_542,N_466);
xnor U650 (N_650,N_555,In_374);
nand U651 (N_651,N_426,In_208);
nand U652 (N_652,In_1465,N_3);
and U653 (N_653,N_512,N_271);
xor U654 (N_654,In_1045,N_427);
nand U655 (N_655,In_1207,N_618);
or U656 (N_656,In_443,In_892);
and U657 (N_657,In_1147,N_306);
and U658 (N_658,In_1267,In_353);
or U659 (N_659,In_1120,N_235);
nor U660 (N_660,In_1191,In_613);
xor U661 (N_661,In_541,In_1025);
nor U662 (N_662,In_595,In_1259);
nor U663 (N_663,In_1343,In_922);
and U664 (N_664,In_623,In_607);
nor U665 (N_665,In_484,N_240);
or U666 (N_666,In_1199,In_646);
nor U667 (N_667,In_91,N_303);
and U668 (N_668,In_305,In_627);
nand U669 (N_669,N_596,In_1116);
xnor U670 (N_670,In_1222,In_912);
nor U671 (N_671,In_906,N_622);
or U672 (N_672,In_257,In_1050);
xnor U673 (N_673,In_1400,N_430);
nor U674 (N_674,In_1455,N_423);
or U675 (N_675,In_1179,In_1140);
or U676 (N_676,In_1408,N_530);
nand U677 (N_677,In_161,In_1022);
and U678 (N_678,N_145,N_152);
and U679 (N_679,N_572,In_1135);
nor U680 (N_680,In_501,N_456);
nand U681 (N_681,N_229,N_142);
and U682 (N_682,N_174,N_516);
or U683 (N_683,N_611,In_451);
nor U684 (N_684,In_1475,N_428);
and U685 (N_685,In_160,In_1091);
and U686 (N_686,In_1362,In_546);
and U687 (N_687,N_534,In_809);
nand U688 (N_688,N_549,In_123);
or U689 (N_689,In_1035,N_49);
and U690 (N_690,In_1276,N_101);
xor U691 (N_691,N_343,In_198);
xnor U692 (N_692,In_725,In_40);
xor U693 (N_693,In_1300,N_394);
or U694 (N_694,In_1327,In_1488);
xor U695 (N_695,N_418,N_137);
nor U696 (N_696,In_968,N_308);
or U697 (N_697,In_79,In_36);
nor U698 (N_698,N_419,In_1403);
and U699 (N_699,In_517,N_228);
nor U700 (N_700,In_1470,N_491);
and U701 (N_701,N_610,In_119);
xnor U702 (N_702,In_624,In_1391);
nand U703 (N_703,N_594,In_1226);
and U704 (N_704,In_961,In_978);
nor U705 (N_705,In_787,In_1264);
and U706 (N_706,In_269,N_175);
xnor U707 (N_707,N_415,N_473);
nand U708 (N_708,In_741,In_1278);
nand U709 (N_709,N_440,In_836);
or U710 (N_710,N_561,N_589);
or U711 (N_711,In_183,In_1046);
nand U712 (N_712,In_663,In_114);
nand U713 (N_713,N_540,N_416);
nor U714 (N_714,N_376,In_563);
nor U715 (N_715,In_688,N_537);
and U716 (N_716,In_1245,In_641);
xnor U717 (N_717,In_1354,N_606);
nand U718 (N_718,N_571,In_1162);
or U719 (N_719,N_585,In_905);
and U720 (N_720,In_362,In_483);
nand U721 (N_721,N_436,In_329);
xor U722 (N_722,In_229,N_522);
nand U723 (N_723,N_607,N_535);
nor U724 (N_724,In_301,N_547);
nand U725 (N_725,N_120,In_328);
and U726 (N_726,N_265,In_782);
nand U727 (N_727,In_669,N_387);
nand U728 (N_728,In_526,N_529);
or U729 (N_729,In_280,N_525);
and U730 (N_730,N_92,In_1251);
or U731 (N_731,N_63,In_289);
nand U732 (N_732,In_529,In_521);
and U733 (N_733,N_176,In_1237);
nand U734 (N_734,In_1106,N_590);
or U735 (N_735,N_122,N_169);
nor U736 (N_736,N_494,N_238);
or U737 (N_737,In_1102,N_493);
nor U738 (N_738,In_1225,N_598);
or U739 (N_739,N_254,N_381);
and U740 (N_740,N_19,N_100);
xnor U741 (N_741,In_446,N_492);
nand U742 (N_742,N_210,In_1194);
nor U743 (N_743,N_135,N_414);
nor U744 (N_744,In_1326,In_102);
xor U745 (N_745,N_425,In_1499);
nor U746 (N_746,N_38,N_434);
nand U747 (N_747,N_189,N_533);
and U748 (N_748,In_1452,In_1394);
and U749 (N_749,In_1320,N_370);
nand U750 (N_750,N_578,In_445);
nor U751 (N_751,N_505,N_98);
xnor U752 (N_752,N_627,N_595);
nor U753 (N_753,N_170,In_1365);
nand U754 (N_754,In_1015,N_245);
xor U755 (N_755,In_1258,In_422);
xor U756 (N_756,In_629,In_441);
and U757 (N_757,N_223,In_141);
nor U758 (N_758,N_514,N_543);
xor U759 (N_759,N_565,N_556);
and U760 (N_760,N_496,N_697);
or U761 (N_761,In_320,N_661);
or U762 (N_762,In_1235,N_467);
and U763 (N_763,N_729,N_630);
or U764 (N_764,N_204,In_184);
nand U765 (N_765,In_1013,N_601);
xnor U766 (N_766,In_182,N_734);
and U767 (N_767,N_519,N_737);
nor U768 (N_768,N_231,N_652);
or U769 (N_769,N_609,N_407);
and U770 (N_770,N_267,In_1195);
or U771 (N_771,N_315,N_501);
nand U772 (N_772,In_387,In_313);
xor U773 (N_773,N_94,In_455);
nor U774 (N_774,N_106,N_503);
nor U775 (N_775,N_658,In_9);
xnor U776 (N_776,In_1476,N_721);
or U777 (N_777,N_517,In_434);
or U778 (N_778,In_760,N_586);
and U779 (N_779,N_605,In_370);
xor U780 (N_780,N_671,N_748);
and U781 (N_781,In_1010,In_815);
and U782 (N_782,N_359,In_1464);
or U783 (N_783,In_1387,N_487);
nand U784 (N_784,In_1429,N_648);
xnor U785 (N_785,N_573,N_36);
nor U786 (N_786,N_305,N_667);
and U787 (N_787,In_105,N_483);
xnor U788 (N_788,N_620,N_506);
or U789 (N_789,In_571,In_110);
xor U790 (N_790,N_45,N_481);
xnor U791 (N_791,N_743,In_1411);
nor U792 (N_792,N_682,N_651);
nand U793 (N_793,In_1291,N_68);
xnor U794 (N_794,In_1188,In_1287);
nand U795 (N_795,In_412,N_382);
or U796 (N_796,N_300,N_735);
xor U797 (N_797,N_568,In_525);
or U798 (N_798,N_502,N_732);
xnor U799 (N_799,N_138,In_1094);
nand U800 (N_800,In_18,N_263);
and U801 (N_801,In_1460,N_647);
and U802 (N_802,N_339,N_747);
or U803 (N_803,N_696,In_349);
or U804 (N_804,In_610,N_713);
xnor U805 (N_805,In_245,N_356);
nand U806 (N_806,In_737,N_218);
nand U807 (N_807,In_1336,N_146);
and U808 (N_808,N_657,N_631);
and U809 (N_809,N_489,In_393);
and U810 (N_810,N_659,In_345);
or U811 (N_811,In_425,In_575);
xor U812 (N_812,N_86,In_746);
and U813 (N_813,N_393,N_11);
xnor U814 (N_814,N_679,N_562);
or U815 (N_815,In_1351,In_376);
nor U816 (N_816,In_1126,In_178);
or U817 (N_817,N_338,N_681);
or U818 (N_818,In_1389,N_708);
xnor U819 (N_819,In_812,N_477);
or U820 (N_820,N_727,N_413);
or U821 (N_821,In_837,N_439);
and U822 (N_822,N_642,N_237);
or U823 (N_823,N_504,In_239);
or U824 (N_824,N_389,In_702);
and U825 (N_825,N_509,N_566);
nor U826 (N_826,N_689,In_1350);
and U827 (N_827,In_1189,N_688);
xnor U828 (N_828,N_390,In_149);
xor U829 (N_829,N_294,In_889);
nand U830 (N_830,In_1277,N_395);
or U831 (N_831,N_72,N_518);
nand U832 (N_832,In_557,In_1070);
and U833 (N_833,In_209,N_645);
nand U834 (N_834,In_586,N_731);
nand U835 (N_835,In_967,In_342);
nor U836 (N_836,In_518,In_1110);
and U837 (N_837,N_337,In_334);
or U838 (N_838,N_587,N_699);
nor U839 (N_839,N_275,In_146);
xnor U840 (N_840,In_1424,In_693);
nand U841 (N_841,N_357,In_1210);
or U842 (N_842,In_935,N_217);
xnor U843 (N_843,In_310,N_615);
nand U844 (N_844,In_389,N_546);
and U845 (N_845,In_109,In_192);
and U846 (N_846,N_558,N_474);
and U847 (N_847,In_908,In_1104);
xnor U848 (N_848,N_349,In_365);
nand U849 (N_849,In_166,N_366);
and U850 (N_850,In_1208,In_145);
and U851 (N_851,In_987,N_369);
nand U852 (N_852,In_1328,N_476);
nor U853 (N_853,N_684,N_741);
or U854 (N_854,In_946,N_709);
or U855 (N_855,In_104,N_104);
nand U856 (N_856,N_531,N_56);
xnor U857 (N_857,N_655,In_330);
xnor U858 (N_858,N_2,N_507);
and U859 (N_859,N_629,N_46);
nand U860 (N_860,N_669,N_628);
xnor U861 (N_861,N_580,In_926);
xnor U862 (N_862,In_1305,In_1296);
or U863 (N_863,In_945,In_687);
xnor U864 (N_864,N_60,In_826);
nand U865 (N_865,N_417,In_1023);
or U866 (N_866,In_93,In_814);
or U867 (N_867,In_1048,In_1057);
or U868 (N_868,In_147,N_26);
nand U869 (N_869,N_479,In_108);
or U870 (N_870,In_1279,In_1219);
nor U871 (N_871,In_1029,In_705);
and U872 (N_872,N_405,In_45);
nor U873 (N_873,N_41,N_574);
nand U874 (N_874,In_1495,In_137);
or U875 (N_875,In_1388,N_569);
or U876 (N_876,N_331,In_58);
or U877 (N_877,In_672,N_299);
xor U878 (N_878,In_1200,N_872);
nor U879 (N_879,N_662,N_392);
nand U880 (N_880,In_759,N_848);
nor U881 (N_881,In_1370,N_795);
or U882 (N_882,N_745,In_778);
nor U883 (N_883,In_459,N_179);
nor U884 (N_884,N_126,In_969);
nor U885 (N_885,N_739,In_754);
nor U886 (N_886,N_181,In_1335);
xor U887 (N_887,N_592,N_836);
or U888 (N_888,In_139,In_528);
nor U889 (N_889,N_720,N_711);
nand U890 (N_890,In_630,N_608);
or U891 (N_891,In_1113,N_860);
nand U892 (N_892,N_297,N_673);
nor U893 (N_893,N_789,N_827);
nor U894 (N_894,N_488,N_722);
nor U895 (N_895,N_341,N_775);
or U896 (N_896,N_830,N_753);
nor U897 (N_897,N_311,N_839);
xnor U898 (N_898,N_670,N_478);
xnor U899 (N_899,N_700,N_420);
and U900 (N_900,N_445,N_251);
or U901 (N_901,N_490,N_485);
or U902 (N_902,N_640,N_873);
and U903 (N_903,In_321,N_464);
xnor U904 (N_904,N_268,N_763);
xor U905 (N_905,N_866,In_1301);
nor U906 (N_906,N_824,In_1163);
xor U907 (N_907,In_846,N_646);
and U908 (N_908,N_704,N_768);
nor U909 (N_909,In_955,N_665);
nor U910 (N_910,N_653,In_373);
and U911 (N_911,N_458,N_835);
xor U912 (N_912,N_779,In_1039);
and U913 (N_913,N_57,N_851);
nand U914 (N_914,N_761,N_442);
nor U915 (N_915,N_61,In_290);
or U916 (N_916,N_134,N_644);
xor U917 (N_917,N_874,In_1402);
or U918 (N_918,In_1359,In_600);
xor U919 (N_919,In_810,N_832);
nand U920 (N_920,N_660,N_842);
nand U921 (N_921,N_649,In_439);
and U922 (N_922,In_38,N_809);
nand U923 (N_923,In_766,In_1304);
or U924 (N_924,In_1168,N_817);
nand U925 (N_925,In_250,In_5);
xnor U926 (N_926,In_8,In_785);
xnor U927 (N_927,N_846,N_676);
nor U928 (N_928,N_144,N_508);
nand U929 (N_929,N_870,N_164);
and U930 (N_930,N_702,N_575);
nor U931 (N_931,In_223,N_829);
or U932 (N_932,N_632,In_67);
xnor U933 (N_933,N_742,In_643);
or U934 (N_934,In_828,N_840);
and U935 (N_935,N_272,N_329);
and U936 (N_936,In_327,In_1453);
or U937 (N_937,In_456,N_808);
or U938 (N_938,N_707,N_855);
nor U939 (N_939,N_856,N_64);
and U940 (N_940,In_424,In_710);
nor U941 (N_941,In_225,N_332);
and U942 (N_942,N_564,In_804);
nor U943 (N_943,N_773,N_668);
nor U944 (N_944,In_243,N_110);
nand U945 (N_945,In_734,N_616);
and U946 (N_946,In_291,In_256);
nor U947 (N_947,N_718,N_755);
xnor U948 (N_948,N_796,N_409);
and U949 (N_949,In_924,N_758);
nor U950 (N_950,In_839,N_710);
xor U951 (N_951,In_1292,N_831);
nand U952 (N_952,In_1355,N_811);
or U953 (N_953,N_771,N_378);
or U954 (N_954,In_1019,N_862);
xor U955 (N_955,In_1415,N_638);
nor U956 (N_956,In_633,In_649);
xor U957 (N_957,In_13,N_834);
xnor U958 (N_958,In_1346,In_520);
nor U959 (N_959,In_238,N_551);
nor U960 (N_960,N_621,In_999);
nand U961 (N_961,N_280,N_800);
and U962 (N_962,N_650,N_261);
xnor U963 (N_963,In_724,N_792);
nand U964 (N_964,In_1009,N_814);
xor U965 (N_965,N_557,N_806);
xor U966 (N_966,In_774,In_1246);
xor U967 (N_967,In_1312,N_782);
or U968 (N_968,In_1393,In_271);
nor U969 (N_969,N_602,N_24);
nand U970 (N_970,N_635,N_849);
and U971 (N_971,N_326,N_784);
or U972 (N_972,N_457,In_763);
nand U973 (N_973,N_220,N_597);
and U974 (N_974,In_1366,N_633);
nor U975 (N_975,N_115,In_491);
nor U976 (N_976,In_185,N_683);
or U977 (N_977,In_29,N_705);
or U978 (N_978,N_583,In_1165);
nor U979 (N_979,N_812,N_65);
and U980 (N_980,In_591,In_748);
xor U981 (N_981,N_858,N_190);
nand U982 (N_982,N_803,N_548);
nor U983 (N_983,N_577,In_382);
nor U984 (N_984,N_498,N_841);
and U985 (N_985,In_1435,N_76);
xor U986 (N_986,N_132,In_572);
xnor U987 (N_987,N_869,N_446);
or U988 (N_988,N_786,N_850);
xor U989 (N_989,N_333,N_599);
and U990 (N_990,In_783,In_850);
nor U991 (N_991,In_909,N_719);
xor U992 (N_992,In_960,N_528);
xor U993 (N_993,In_64,In_923);
or U994 (N_994,N_810,N_459);
nand U995 (N_995,In_113,In_390);
xnor U996 (N_996,In_130,N_863);
or U997 (N_997,N_675,N_733);
nor U998 (N_998,In_914,In_266);
and U999 (N_999,In_177,N_744);
xnor U1000 (N_1000,N_581,N_422);
nor U1001 (N_1001,In_870,N_805);
and U1002 (N_1002,N_956,N_716);
xor U1003 (N_1003,N_906,N_17);
nor U1004 (N_1004,N_911,N_791);
nand U1005 (N_1005,N_160,N_968);
nor U1006 (N_1006,N_785,In_879);
nand U1007 (N_1007,N_636,N_471);
xor U1008 (N_1008,N_286,In_377);
nand U1009 (N_1009,N_988,N_818);
or U1010 (N_1010,In_1451,N_411);
xnor U1011 (N_1011,N_604,N_790);
nand U1012 (N_1012,In_324,N_859);
xor U1013 (N_1013,N_801,N_754);
xnor U1014 (N_1014,N_207,N_29);
or U1015 (N_1015,In_616,N_912);
and U1016 (N_1016,In_436,In_159);
nand U1017 (N_1017,In_1338,N_527);
nand U1018 (N_1018,In_27,N_781);
or U1019 (N_1019,In_1173,In_173);
or U1020 (N_1020,N_686,N_270);
nor U1021 (N_1021,N_854,N_674);
nand U1022 (N_1022,N_989,In_652);
nand U1023 (N_1023,In_249,N_706);
or U1024 (N_1024,In_22,N_940);
or U1025 (N_1025,N_955,N_295);
or U1026 (N_1026,N_915,In_154);
xor U1027 (N_1027,N_961,N_979);
nand U1028 (N_1028,N_930,N_553);
or U1029 (N_1029,In_261,N_944);
or U1030 (N_1030,In_993,N_398);
or U1031 (N_1031,N_804,In_226);
nor U1032 (N_1032,In_1496,In_457);
nor U1033 (N_1033,N_904,N_678);
xor U1034 (N_1034,In_1044,N_693);
or U1035 (N_1035,N_157,N_838);
xnor U1036 (N_1036,N_695,N_780);
or U1037 (N_1037,N_746,N_750);
and U1038 (N_1038,In_1205,N_821);
nor U1039 (N_1039,N_579,In_1093);
and U1040 (N_1040,N_402,N_901);
xnor U1041 (N_1041,N_766,N_909);
nor U1042 (N_1042,N_756,In_120);
nand U1043 (N_1043,N_148,N_973);
nand U1044 (N_1044,N_895,N_199);
xor U1045 (N_1045,N_725,N_816);
nand U1046 (N_1046,In_1439,N_905);
nor U1047 (N_1047,N_626,N_424);
nand U1048 (N_1048,N_524,N_890);
nor U1049 (N_1049,N_996,N_900);
or U1050 (N_1050,N_883,N_910);
nand U1051 (N_1051,In_472,N_656);
or U1052 (N_1052,N_593,N_880);
and U1053 (N_1053,N_991,N_749);
nand U1054 (N_1054,In_885,N_429);
and U1055 (N_1055,In_742,N_521);
xnor U1056 (N_1056,N_828,N_762);
xor U1057 (N_1057,N_926,N_985);
xor U1058 (N_1058,N_952,N_560);
and U1059 (N_1059,N_760,In_920);
xor U1060 (N_1060,In_751,In_1314);
nor U1061 (N_1061,N_764,N_939);
nor U1062 (N_1062,N_797,In_1112);
nor U1063 (N_1063,In_73,N_403);
nand U1064 (N_1064,N_34,N_776);
xnor U1065 (N_1065,N_844,N_923);
xor U1066 (N_1066,N_868,In_1483);
or U1067 (N_1067,N_307,In_992);
nand U1068 (N_1068,N_236,In_618);
nand U1069 (N_1069,N_947,N_677);
nand U1070 (N_1070,N_953,N_273);
nor U1071 (N_1071,In_282,N_486);
nor U1072 (N_1072,N_347,N_787);
nand U1073 (N_1073,N_957,N_603);
or U1074 (N_1074,In_1253,N_871);
nand U1075 (N_1075,N_891,N_922);
xor U1076 (N_1076,In_878,N_799);
xnor U1077 (N_1077,N_853,N_970);
xor U1078 (N_1078,N_962,N_454);
nor U1079 (N_1079,N_950,N_447);
nor U1080 (N_1080,In_620,N_938);
or U1081 (N_1081,N_933,N_539);
and U1082 (N_1082,N_698,N_717);
nor U1083 (N_1083,N_685,N_975);
nor U1084 (N_1084,In_1004,In_246);
nor U1085 (N_1085,In_854,In_1073);
xnor U1086 (N_1086,N_703,In_590);
or U1087 (N_1087,In_140,N_619);
nand U1088 (N_1088,N_443,N_896);
xnor U1089 (N_1089,N_943,N_982);
nand U1090 (N_1090,N_680,In_1183);
nor U1091 (N_1091,In_757,N_317);
and U1092 (N_1092,N_345,N_451);
nor U1093 (N_1093,N_23,N_410);
nor U1094 (N_1094,In_1156,N_807);
xor U1095 (N_1095,In_270,In_325);
nand U1096 (N_1096,N_93,N_233);
xor U1097 (N_1097,N_141,N_783);
nor U1098 (N_1098,In_1088,N_10);
xor U1099 (N_1099,N_591,N_949);
nand U1100 (N_1100,N_520,N_845);
xnor U1101 (N_1101,N_879,N_692);
and U1102 (N_1102,In_1459,N_751);
or U1103 (N_1103,In_564,N_994);
nand U1104 (N_1104,N_981,N_437);
or U1105 (N_1105,N_715,N_274);
nand U1106 (N_1106,In_4,In_1197);
nand U1107 (N_1107,N_163,N_159);
or U1108 (N_1108,In_1419,N_825);
or U1109 (N_1109,N_886,N_360);
or U1110 (N_1110,N_899,N_865);
or U1111 (N_1111,N_788,N_945);
or U1112 (N_1112,N_153,N_770);
xnor U1113 (N_1113,In_509,N_769);
xnor U1114 (N_1114,In_799,N_963);
nand U1115 (N_1115,In_272,N_937);
nand U1116 (N_1116,In_364,N_663);
nor U1117 (N_1117,N_964,N_974);
or U1118 (N_1118,N_765,N_614);
nor U1119 (N_1119,In_470,N_972);
and U1120 (N_1120,N_738,N_954);
nand U1121 (N_1121,N_358,N_536);
xnor U1122 (N_1122,In_323,In_928);
nand U1123 (N_1123,In_312,N_864);
or U1124 (N_1124,N_847,In_954);
and U1125 (N_1125,N_262,N_1045);
and U1126 (N_1126,N_559,N_1069);
nor U1127 (N_1127,N_511,In_1375);
nand U1128 (N_1128,N_532,In_176);
and U1129 (N_1129,In_1399,In_1111);
nand U1130 (N_1130,N_1009,N_1104);
nand U1131 (N_1131,N_167,In_1364);
xor U1132 (N_1132,N_1062,In_346);
xor U1133 (N_1133,N_1066,N_774);
nand U1134 (N_1134,In_308,N_1103);
nand U1135 (N_1135,N_935,N_876);
or U1136 (N_1136,N_1067,N_1053);
and U1137 (N_1137,N_1010,N_730);
nand U1138 (N_1138,In_1412,N_1043);
xor U1139 (N_1139,N_1026,N_1097);
nand U1140 (N_1140,N_1122,In_24);
or U1141 (N_1141,N_1090,N_1056);
nand U1142 (N_1142,N_852,N_843);
or U1143 (N_1143,N_798,N_1063);
nor U1144 (N_1144,N_1044,N_1041);
xnor U1145 (N_1145,N_977,N_857);
nand U1146 (N_1146,N_819,N_861);
xor U1147 (N_1147,N_998,N_1018);
and U1148 (N_1148,N_712,N_1019);
or U1149 (N_1149,In_1378,N_449);
and U1150 (N_1150,In_1096,N_177);
xor U1151 (N_1151,N_826,N_1068);
xor U1152 (N_1152,In_762,N_211);
nand U1153 (N_1153,In_1313,In_304);
nand U1154 (N_1154,N_951,N_1077);
and U1155 (N_1155,In_89,N_1102);
or U1156 (N_1156,N_1059,N_1030);
nor U1157 (N_1157,In_788,N_664);
and U1158 (N_1158,N_1029,In_1284);
or U1159 (N_1159,N_438,N_987);
xor U1160 (N_1160,N_1092,N_515);
xor U1161 (N_1161,N_1031,N_759);
nor U1162 (N_1162,N_1115,N_624);
nor U1163 (N_1163,N_1040,N_639);
or U1164 (N_1164,In_959,N_1037);
nand U1165 (N_1165,N_924,N_884);
xnor U1166 (N_1166,N_918,N_1058);
nor U1167 (N_1167,N_567,N_936);
or U1168 (N_1168,N_778,In_407);
nor U1169 (N_1169,N_740,N_929);
xor U1170 (N_1170,N_813,In_156);
and U1171 (N_1171,N_931,In_411);
and U1172 (N_1172,N_1098,N_691);
or U1173 (N_1173,N_978,N_1083);
and U1174 (N_1174,N_1070,N_984);
nor U1175 (N_1175,N_383,N_1027);
or U1176 (N_1176,N_980,N_1012);
nand U1177 (N_1177,N_1046,N_1007);
or U1178 (N_1178,N_903,In_1352);
or U1179 (N_1179,N_1080,In_674);
nor U1180 (N_1180,N_960,N_902);
or U1181 (N_1181,N_1000,In_416);
or U1182 (N_1182,N_224,In_391);
nor U1183 (N_1183,N_1108,N_613);
or U1184 (N_1184,N_882,N_875);
and U1185 (N_1185,N_995,In_465);
nor U1186 (N_1186,N_920,N_921);
or U1187 (N_1187,In_764,N_687);
nand U1188 (N_1188,N_877,N_1106);
nand U1189 (N_1189,In_1418,N_1072);
xor U1190 (N_1190,N_913,In_138);
nor U1191 (N_1191,In_582,In_806);
nor U1192 (N_1192,In_886,N_641);
nand U1193 (N_1193,N_1065,N_767);
xor U1194 (N_1194,N_867,N_969);
nor U1195 (N_1195,N_1099,In_1413);
nand U1196 (N_1196,N_772,In_527);
nor U1197 (N_1197,N_350,N_582);
xnor U1198 (N_1198,In_111,In_448);
xnor U1199 (N_1199,N_1111,N_1096);
nand U1200 (N_1200,N_321,N_997);
nand U1201 (N_1201,N_934,N_1101);
nand U1202 (N_1202,N_335,N_510);
nor U1203 (N_1203,N_1034,N_1047);
nor U1204 (N_1204,In_578,N_837);
xor U1205 (N_1205,N_986,N_1089);
xnor U1206 (N_1206,N_1087,In_1020);
and U1207 (N_1207,In_723,N_1076);
nand U1208 (N_1208,N_1023,In_1052);
and U1209 (N_1209,N_1038,N_726);
or U1210 (N_1210,In_255,N_946);
xor U1211 (N_1211,N_958,N_184);
or U1212 (N_1212,N_584,N_1015);
and U1213 (N_1213,N_250,N_526);
or U1214 (N_1214,In_1085,In_148);
and U1215 (N_1215,N_967,In_1047);
and U1216 (N_1216,N_1024,N_736);
xor U1217 (N_1217,N_752,N_728);
and U1218 (N_1218,N_959,N_623);
nand U1219 (N_1219,N_965,N_1036);
and U1220 (N_1220,N_1085,In_800);
xor U1221 (N_1221,N_1006,N_1035);
and U1222 (N_1222,N_1119,In_1463);
xor U1223 (N_1223,N_898,N_714);
or U1224 (N_1224,N_637,In_915);
or U1225 (N_1225,N_242,N_892);
xnor U1226 (N_1226,N_1112,N_385);
nor U1227 (N_1227,N_202,N_1055);
nand U1228 (N_1228,N_694,N_1084);
and U1229 (N_1229,N_523,In_1240);
nor U1230 (N_1230,N_1093,N_1114);
or U1231 (N_1231,In_276,N_1105);
and U1232 (N_1232,N_71,N_1075);
xnor U1233 (N_1233,N_391,In_132);
and U1234 (N_1234,N_1005,In_175);
or U1235 (N_1235,N_897,N_893);
and U1236 (N_1236,N_421,N_1086);
nor U1237 (N_1237,N_1071,In_287);
or U1238 (N_1238,N_73,N_1107);
or U1239 (N_1239,N_634,N_1081);
nand U1240 (N_1240,N_1048,In_843);
and U1241 (N_1241,In_587,N_600);
or U1242 (N_1242,N_463,N_1117);
or U1243 (N_1243,In_1077,N_1021);
and U1244 (N_1244,N_1118,N_1094);
nor U1245 (N_1245,In_283,N_916);
xor U1246 (N_1246,In_989,N_328);
xnor U1247 (N_1247,N_452,N_1028);
or U1248 (N_1248,N_802,N_552);
nand U1249 (N_1249,In_515,N_1110);
and U1250 (N_1250,N_1144,N_1187);
nand U1251 (N_1251,N_793,N_1134);
xor U1252 (N_1252,N_625,N_1051);
and U1253 (N_1253,N_1211,N_1082);
and U1254 (N_1254,N_1238,N_1174);
or U1255 (N_1255,N_1128,N_1145);
nand U1256 (N_1256,N_1204,N_1179);
and U1257 (N_1257,N_889,N_1192);
and U1258 (N_1258,N_1175,N_1033);
or U1259 (N_1259,In_25,N_1241);
nor U1260 (N_1260,N_1199,N_1232);
and U1261 (N_1261,N_513,N_887);
xor U1262 (N_1262,N_1191,N_1124);
and U1263 (N_1263,N_448,N_1088);
or U1264 (N_1264,N_1149,N_1132);
and U1265 (N_1265,N_1140,N_1141);
and U1266 (N_1266,N_1060,N_823);
nand U1267 (N_1267,N_1061,N_1156);
and U1268 (N_1268,N_1209,N_1020);
or U1269 (N_1269,N_1248,In_429);
nor U1270 (N_1270,N_888,N_1198);
nand U1271 (N_1271,N_1226,In_1159);
nand U1272 (N_1272,N_1074,N_1123);
nor U1273 (N_1273,N_460,N_1220);
or U1274 (N_1274,N_1231,N_431);
nand U1275 (N_1275,N_1042,N_690);
xnor U1276 (N_1276,N_1216,N_1109);
xor U1277 (N_1277,N_1146,N_976);
and U1278 (N_1278,N_1221,N_1172);
or U1279 (N_1279,N_894,N_1166);
xor U1280 (N_1280,N_1161,N_221);
and U1281 (N_1281,N_1197,In_326);
nor U1282 (N_1282,N_1185,N_612);
or U1283 (N_1283,N_1017,N_1163);
or U1284 (N_1284,N_550,N_1233);
nor U1285 (N_1285,N_269,N_1126);
or U1286 (N_1286,N_1178,N_1165);
and U1287 (N_1287,N_1078,N_1223);
nor U1288 (N_1288,N_666,In_1462);
and U1289 (N_1289,In_1261,N_1168);
and U1290 (N_1290,N_1002,N_1171);
nand U1291 (N_1291,N_1193,N_1153);
nand U1292 (N_1292,N_1025,N_932);
nor U1293 (N_1293,N_1222,N_1224);
or U1294 (N_1294,In_1440,N_820);
nand U1295 (N_1295,N_919,N_1249);
or U1296 (N_1296,N_1236,In_661);
or U1297 (N_1297,N_1169,N_408);
or U1298 (N_1298,In_1317,N_966);
and U1299 (N_1299,N_1235,In_1444);
or U1300 (N_1300,N_1239,N_1189);
and U1301 (N_1301,In_1308,N_1160);
nand U1302 (N_1302,N_1057,N_244);
nor U1303 (N_1303,N_1001,N_1181);
and U1304 (N_1304,N_1150,N_1162);
or U1305 (N_1305,N_1210,N_1022);
nand U1306 (N_1306,N_367,N_1214);
or U1307 (N_1307,N_1202,N_881);
and U1308 (N_1308,N_1073,N_1054);
and U1309 (N_1309,N_1159,In_129);
xnor U1310 (N_1310,N_352,N_1167);
and U1311 (N_1311,N_1052,N_1016);
nor U1312 (N_1312,N_1182,N_927);
nand U1313 (N_1313,N_1184,N_942);
xnor U1314 (N_1314,N_990,N_1203);
or U1315 (N_1315,N_316,N_1032);
xnor U1316 (N_1316,N_1135,N_777);
or U1317 (N_1317,N_554,N_1240);
and U1318 (N_1318,N_723,N_971);
or U1319 (N_1319,N_1116,N_1194);
nor U1320 (N_1320,N_404,N_1151);
xnor U1321 (N_1321,N_1180,N_1206);
or U1322 (N_1322,N_336,N_1129);
and U1323 (N_1323,N_1188,N_654);
nand U1324 (N_1324,N_1143,N_1147);
nor U1325 (N_1325,N_878,N_1200);
nand U1326 (N_1326,N_1120,N_1217);
and U1327 (N_1327,N_1142,N_1130);
nand U1328 (N_1328,N_1139,In_1161);
nor U1329 (N_1329,N_1121,N_1131);
and U1330 (N_1330,N_1246,N_701);
and U1331 (N_1331,In_651,N_1113);
or U1332 (N_1332,N_724,N_1183);
and U1333 (N_1333,N_1164,N_1219);
nor U1334 (N_1334,In_1290,N_1176);
and U1335 (N_1335,N_1190,N_1157);
or U1336 (N_1336,N_1158,N_925);
xnor U1337 (N_1337,N_1049,N_1154);
nor U1338 (N_1338,N_1136,N_1138);
xor U1339 (N_1339,N_672,N_1215);
nor U1340 (N_1340,N_1064,N_907);
nor U1341 (N_1341,N_1229,N_999);
nor U1342 (N_1342,N_1014,N_992);
nor U1343 (N_1343,N_1225,N_1208);
xnor U1344 (N_1344,In_461,N_1245);
or U1345 (N_1345,N_401,N_1095);
or U1346 (N_1346,N_1212,N_1230);
nor U1347 (N_1347,N_1079,N_822);
xor U1348 (N_1348,N_757,N_1148);
nor U1349 (N_1349,N_1201,N_1186);
xor U1350 (N_1350,N_1133,N_1008);
nor U1351 (N_1351,In_951,N_1234);
or U1352 (N_1352,In_1026,N_1195);
nor U1353 (N_1353,N_928,N_1213);
and U1354 (N_1354,In_824,N_1127);
nand U1355 (N_1355,N_983,N_1207);
nand U1356 (N_1356,N_993,N_1228);
nor U1357 (N_1357,N_815,N_643);
nand U1358 (N_1358,N_1177,N_1011);
xnor U1359 (N_1359,N_885,N_1003);
and U1360 (N_1360,N_1050,N_1173);
nor U1361 (N_1361,N_1125,N_1004);
nand U1362 (N_1362,N_1218,N_941);
and U1363 (N_1363,N_948,In_982);
nand U1364 (N_1364,N_1170,N_794);
nor U1365 (N_1365,N_1100,N_833);
and U1366 (N_1366,N_917,N_1243);
xnor U1367 (N_1367,N_1205,N_1244);
nor U1368 (N_1368,N_1137,N_914);
xnor U1369 (N_1369,N_908,N_1237);
and U1370 (N_1370,N_1227,N_1152);
xor U1371 (N_1371,N_1242,N_388);
or U1372 (N_1372,N_1247,N_1091);
nor U1373 (N_1373,N_1013,N_1196);
xnor U1374 (N_1374,N_1155,N_1039);
nand U1375 (N_1375,N_1363,N_1262);
xor U1376 (N_1376,N_1346,N_1275);
or U1377 (N_1377,N_1310,N_1261);
xor U1378 (N_1378,N_1250,N_1355);
and U1379 (N_1379,N_1307,N_1285);
xor U1380 (N_1380,N_1282,N_1364);
nand U1381 (N_1381,N_1277,N_1337);
xor U1382 (N_1382,N_1256,N_1362);
nand U1383 (N_1383,N_1257,N_1328);
nand U1384 (N_1384,N_1353,N_1318);
xor U1385 (N_1385,N_1343,N_1359);
or U1386 (N_1386,N_1293,N_1267);
nor U1387 (N_1387,N_1370,N_1356);
or U1388 (N_1388,N_1340,N_1268);
nand U1389 (N_1389,N_1294,N_1271);
xnor U1390 (N_1390,N_1305,N_1350);
nand U1391 (N_1391,N_1361,N_1254);
and U1392 (N_1392,N_1352,N_1351);
or U1393 (N_1393,N_1321,N_1258);
nor U1394 (N_1394,N_1300,N_1276);
nor U1395 (N_1395,N_1279,N_1368);
or U1396 (N_1396,N_1316,N_1345);
and U1397 (N_1397,N_1309,N_1304);
nand U1398 (N_1398,N_1292,N_1325);
nand U1399 (N_1399,N_1374,N_1303);
xnor U1400 (N_1400,N_1357,N_1334);
nor U1401 (N_1401,N_1358,N_1255);
and U1402 (N_1402,N_1348,N_1284);
xnor U1403 (N_1403,N_1270,N_1280);
nand U1404 (N_1404,N_1299,N_1313);
nand U1405 (N_1405,N_1320,N_1286);
or U1406 (N_1406,N_1291,N_1281);
nand U1407 (N_1407,N_1327,N_1323);
nand U1408 (N_1408,N_1312,N_1333);
nand U1409 (N_1409,N_1287,N_1344);
nor U1410 (N_1410,N_1265,N_1349);
nand U1411 (N_1411,N_1260,N_1331);
xnor U1412 (N_1412,N_1295,N_1302);
nand U1413 (N_1413,N_1336,N_1366);
nand U1414 (N_1414,N_1332,N_1324);
or U1415 (N_1415,N_1308,N_1272);
or U1416 (N_1416,N_1252,N_1369);
xnor U1417 (N_1417,N_1354,N_1371);
nand U1418 (N_1418,N_1311,N_1347);
xnor U1419 (N_1419,N_1259,N_1365);
nor U1420 (N_1420,N_1372,N_1330);
xnor U1421 (N_1421,N_1301,N_1296);
xnor U1422 (N_1422,N_1341,N_1273);
nand U1423 (N_1423,N_1297,N_1306);
or U1424 (N_1424,N_1335,N_1269);
nand U1425 (N_1425,N_1278,N_1319);
nand U1426 (N_1426,N_1263,N_1367);
nand U1427 (N_1427,N_1298,N_1329);
and U1428 (N_1428,N_1290,N_1283);
nor U1429 (N_1429,N_1264,N_1253);
nor U1430 (N_1430,N_1266,N_1338);
and U1431 (N_1431,N_1339,N_1315);
and U1432 (N_1432,N_1289,N_1326);
xor U1433 (N_1433,N_1317,N_1274);
xnor U1434 (N_1434,N_1314,N_1251);
and U1435 (N_1435,N_1360,N_1373);
nor U1436 (N_1436,N_1288,N_1322);
and U1437 (N_1437,N_1342,N_1337);
nand U1438 (N_1438,N_1253,N_1309);
or U1439 (N_1439,N_1258,N_1294);
and U1440 (N_1440,N_1329,N_1292);
and U1441 (N_1441,N_1363,N_1341);
or U1442 (N_1442,N_1268,N_1262);
xnor U1443 (N_1443,N_1342,N_1355);
nor U1444 (N_1444,N_1287,N_1253);
or U1445 (N_1445,N_1333,N_1281);
nor U1446 (N_1446,N_1282,N_1298);
xnor U1447 (N_1447,N_1296,N_1344);
or U1448 (N_1448,N_1373,N_1273);
nand U1449 (N_1449,N_1314,N_1270);
nor U1450 (N_1450,N_1372,N_1314);
and U1451 (N_1451,N_1310,N_1309);
nand U1452 (N_1452,N_1356,N_1324);
xnor U1453 (N_1453,N_1299,N_1349);
nand U1454 (N_1454,N_1369,N_1302);
nand U1455 (N_1455,N_1311,N_1263);
nand U1456 (N_1456,N_1315,N_1367);
xnor U1457 (N_1457,N_1321,N_1306);
nor U1458 (N_1458,N_1250,N_1321);
xor U1459 (N_1459,N_1263,N_1351);
xor U1460 (N_1460,N_1307,N_1370);
or U1461 (N_1461,N_1346,N_1316);
nor U1462 (N_1462,N_1292,N_1341);
nand U1463 (N_1463,N_1296,N_1347);
nor U1464 (N_1464,N_1349,N_1365);
nor U1465 (N_1465,N_1250,N_1366);
nor U1466 (N_1466,N_1270,N_1272);
xnor U1467 (N_1467,N_1327,N_1304);
xnor U1468 (N_1468,N_1333,N_1252);
or U1469 (N_1469,N_1323,N_1328);
nand U1470 (N_1470,N_1261,N_1300);
nor U1471 (N_1471,N_1263,N_1286);
xnor U1472 (N_1472,N_1333,N_1282);
nand U1473 (N_1473,N_1374,N_1352);
nor U1474 (N_1474,N_1282,N_1268);
xor U1475 (N_1475,N_1294,N_1286);
and U1476 (N_1476,N_1250,N_1343);
xor U1477 (N_1477,N_1269,N_1330);
and U1478 (N_1478,N_1290,N_1361);
nor U1479 (N_1479,N_1275,N_1259);
nand U1480 (N_1480,N_1255,N_1267);
nand U1481 (N_1481,N_1282,N_1270);
nor U1482 (N_1482,N_1340,N_1266);
xnor U1483 (N_1483,N_1262,N_1305);
or U1484 (N_1484,N_1321,N_1315);
nor U1485 (N_1485,N_1369,N_1364);
nand U1486 (N_1486,N_1283,N_1286);
nor U1487 (N_1487,N_1348,N_1345);
nor U1488 (N_1488,N_1339,N_1299);
and U1489 (N_1489,N_1351,N_1354);
xor U1490 (N_1490,N_1348,N_1351);
and U1491 (N_1491,N_1284,N_1326);
xor U1492 (N_1492,N_1331,N_1250);
or U1493 (N_1493,N_1284,N_1305);
nand U1494 (N_1494,N_1320,N_1258);
and U1495 (N_1495,N_1374,N_1270);
nand U1496 (N_1496,N_1348,N_1333);
nand U1497 (N_1497,N_1287,N_1350);
or U1498 (N_1498,N_1296,N_1286);
nand U1499 (N_1499,N_1344,N_1257);
nor U1500 (N_1500,N_1474,N_1493);
or U1501 (N_1501,N_1378,N_1415);
and U1502 (N_1502,N_1422,N_1487);
and U1503 (N_1503,N_1477,N_1483);
and U1504 (N_1504,N_1490,N_1453);
xor U1505 (N_1505,N_1495,N_1430);
nand U1506 (N_1506,N_1395,N_1438);
nor U1507 (N_1507,N_1407,N_1467);
nand U1508 (N_1508,N_1377,N_1496);
xor U1509 (N_1509,N_1416,N_1442);
xnor U1510 (N_1510,N_1476,N_1478);
or U1511 (N_1511,N_1439,N_1441);
nor U1512 (N_1512,N_1394,N_1457);
xnor U1513 (N_1513,N_1402,N_1473);
or U1514 (N_1514,N_1421,N_1385);
and U1515 (N_1515,N_1425,N_1452);
and U1516 (N_1516,N_1494,N_1498);
xnor U1517 (N_1517,N_1440,N_1449);
or U1518 (N_1518,N_1383,N_1489);
nor U1519 (N_1519,N_1399,N_1437);
xnor U1520 (N_1520,N_1409,N_1451);
xnor U1521 (N_1521,N_1488,N_1432);
nand U1522 (N_1522,N_1387,N_1391);
or U1523 (N_1523,N_1403,N_1389);
xor U1524 (N_1524,N_1390,N_1386);
xnor U1525 (N_1525,N_1384,N_1435);
xnor U1526 (N_1526,N_1427,N_1454);
xnor U1527 (N_1527,N_1461,N_1418);
xnor U1528 (N_1528,N_1396,N_1382);
xor U1529 (N_1529,N_1443,N_1456);
or U1530 (N_1530,N_1376,N_1499);
xor U1531 (N_1531,N_1468,N_1419);
nand U1532 (N_1532,N_1471,N_1408);
and U1533 (N_1533,N_1431,N_1466);
nor U1534 (N_1534,N_1460,N_1463);
and U1535 (N_1535,N_1459,N_1446);
xnor U1536 (N_1536,N_1401,N_1469);
and U1537 (N_1537,N_1436,N_1413);
nor U1538 (N_1538,N_1375,N_1428);
xnor U1539 (N_1539,N_1414,N_1405);
nand U1540 (N_1540,N_1429,N_1479);
and U1541 (N_1541,N_1423,N_1491);
nor U1542 (N_1542,N_1388,N_1481);
or U1543 (N_1543,N_1404,N_1412);
nor U1544 (N_1544,N_1444,N_1424);
nor U1545 (N_1545,N_1411,N_1485);
nand U1546 (N_1546,N_1381,N_1450);
nor U1547 (N_1547,N_1400,N_1410);
xnor U1548 (N_1548,N_1380,N_1480);
xor U1549 (N_1549,N_1475,N_1379);
xnor U1550 (N_1550,N_1497,N_1434);
xor U1551 (N_1551,N_1472,N_1426);
nand U1552 (N_1552,N_1448,N_1455);
and U1553 (N_1553,N_1484,N_1492);
or U1554 (N_1554,N_1406,N_1398);
nor U1555 (N_1555,N_1447,N_1465);
nand U1556 (N_1556,N_1462,N_1393);
nand U1557 (N_1557,N_1464,N_1417);
and U1558 (N_1558,N_1397,N_1486);
xor U1559 (N_1559,N_1458,N_1445);
nand U1560 (N_1560,N_1433,N_1470);
or U1561 (N_1561,N_1392,N_1420);
and U1562 (N_1562,N_1482,N_1498);
xnor U1563 (N_1563,N_1417,N_1406);
nor U1564 (N_1564,N_1389,N_1376);
nand U1565 (N_1565,N_1485,N_1482);
nor U1566 (N_1566,N_1427,N_1408);
nor U1567 (N_1567,N_1452,N_1408);
and U1568 (N_1568,N_1422,N_1396);
xnor U1569 (N_1569,N_1464,N_1416);
and U1570 (N_1570,N_1493,N_1443);
or U1571 (N_1571,N_1445,N_1470);
nand U1572 (N_1572,N_1492,N_1421);
nand U1573 (N_1573,N_1462,N_1380);
or U1574 (N_1574,N_1392,N_1490);
nand U1575 (N_1575,N_1377,N_1479);
or U1576 (N_1576,N_1386,N_1398);
xnor U1577 (N_1577,N_1483,N_1452);
xnor U1578 (N_1578,N_1436,N_1455);
nor U1579 (N_1579,N_1379,N_1418);
nor U1580 (N_1580,N_1385,N_1461);
nor U1581 (N_1581,N_1426,N_1390);
nor U1582 (N_1582,N_1407,N_1392);
nor U1583 (N_1583,N_1455,N_1385);
xnor U1584 (N_1584,N_1440,N_1375);
or U1585 (N_1585,N_1384,N_1377);
nand U1586 (N_1586,N_1473,N_1434);
xnor U1587 (N_1587,N_1495,N_1379);
and U1588 (N_1588,N_1409,N_1491);
and U1589 (N_1589,N_1499,N_1457);
or U1590 (N_1590,N_1395,N_1425);
nand U1591 (N_1591,N_1421,N_1496);
nor U1592 (N_1592,N_1397,N_1385);
and U1593 (N_1593,N_1438,N_1473);
xor U1594 (N_1594,N_1408,N_1389);
nand U1595 (N_1595,N_1478,N_1400);
nand U1596 (N_1596,N_1382,N_1438);
xnor U1597 (N_1597,N_1465,N_1467);
nand U1598 (N_1598,N_1383,N_1472);
xnor U1599 (N_1599,N_1423,N_1463);
nand U1600 (N_1600,N_1426,N_1379);
nor U1601 (N_1601,N_1451,N_1447);
nor U1602 (N_1602,N_1478,N_1437);
nor U1603 (N_1603,N_1428,N_1483);
nand U1604 (N_1604,N_1439,N_1487);
and U1605 (N_1605,N_1488,N_1485);
nand U1606 (N_1606,N_1413,N_1461);
nand U1607 (N_1607,N_1378,N_1482);
nand U1608 (N_1608,N_1389,N_1480);
or U1609 (N_1609,N_1380,N_1445);
or U1610 (N_1610,N_1399,N_1431);
nand U1611 (N_1611,N_1479,N_1396);
or U1612 (N_1612,N_1488,N_1492);
nand U1613 (N_1613,N_1471,N_1393);
xor U1614 (N_1614,N_1434,N_1466);
nand U1615 (N_1615,N_1469,N_1406);
or U1616 (N_1616,N_1479,N_1417);
nor U1617 (N_1617,N_1495,N_1414);
and U1618 (N_1618,N_1436,N_1390);
nand U1619 (N_1619,N_1381,N_1467);
or U1620 (N_1620,N_1433,N_1465);
nor U1621 (N_1621,N_1483,N_1473);
nor U1622 (N_1622,N_1472,N_1410);
nor U1623 (N_1623,N_1426,N_1444);
nor U1624 (N_1624,N_1479,N_1424);
nand U1625 (N_1625,N_1548,N_1516);
nand U1626 (N_1626,N_1617,N_1541);
xnor U1627 (N_1627,N_1534,N_1568);
and U1628 (N_1628,N_1526,N_1549);
nand U1629 (N_1629,N_1545,N_1509);
nand U1630 (N_1630,N_1607,N_1585);
xor U1631 (N_1631,N_1610,N_1606);
and U1632 (N_1632,N_1561,N_1618);
nand U1633 (N_1633,N_1578,N_1592);
or U1634 (N_1634,N_1587,N_1544);
nor U1635 (N_1635,N_1570,N_1555);
and U1636 (N_1636,N_1563,N_1581);
nor U1637 (N_1637,N_1623,N_1537);
nor U1638 (N_1638,N_1591,N_1566);
xor U1639 (N_1639,N_1624,N_1553);
or U1640 (N_1640,N_1574,N_1572);
xnor U1641 (N_1641,N_1595,N_1609);
xor U1642 (N_1642,N_1546,N_1521);
and U1643 (N_1643,N_1525,N_1613);
xnor U1644 (N_1644,N_1508,N_1515);
nor U1645 (N_1645,N_1535,N_1589);
nand U1646 (N_1646,N_1611,N_1512);
nand U1647 (N_1647,N_1506,N_1522);
nand U1648 (N_1648,N_1567,N_1518);
nor U1649 (N_1649,N_1619,N_1604);
nor U1650 (N_1650,N_1565,N_1536);
xor U1651 (N_1651,N_1519,N_1575);
xor U1652 (N_1652,N_1556,N_1596);
or U1653 (N_1653,N_1579,N_1603);
xor U1654 (N_1654,N_1576,N_1500);
nor U1655 (N_1655,N_1540,N_1505);
and U1656 (N_1656,N_1622,N_1530);
nor U1657 (N_1657,N_1547,N_1582);
xnor U1658 (N_1658,N_1513,N_1539);
or U1659 (N_1659,N_1614,N_1550);
and U1660 (N_1660,N_1538,N_1503);
xnor U1661 (N_1661,N_1501,N_1529);
or U1662 (N_1662,N_1524,N_1562);
and U1663 (N_1663,N_1520,N_1510);
xor U1664 (N_1664,N_1573,N_1514);
or U1665 (N_1665,N_1569,N_1559);
and U1666 (N_1666,N_1588,N_1533);
nand U1667 (N_1667,N_1615,N_1532);
xnor U1668 (N_1668,N_1551,N_1598);
nor U1669 (N_1669,N_1571,N_1602);
and U1670 (N_1670,N_1552,N_1517);
nor U1671 (N_1671,N_1511,N_1554);
and U1672 (N_1672,N_1583,N_1590);
nor U1673 (N_1673,N_1564,N_1577);
or U1674 (N_1674,N_1594,N_1612);
nor U1675 (N_1675,N_1601,N_1543);
nand U1676 (N_1676,N_1527,N_1605);
nor U1677 (N_1677,N_1558,N_1507);
and U1678 (N_1678,N_1600,N_1608);
or U1679 (N_1679,N_1616,N_1528);
xor U1680 (N_1680,N_1557,N_1584);
or U1681 (N_1681,N_1531,N_1597);
and U1682 (N_1682,N_1523,N_1542);
nand U1683 (N_1683,N_1593,N_1586);
and U1684 (N_1684,N_1599,N_1580);
xor U1685 (N_1685,N_1560,N_1620);
nand U1686 (N_1686,N_1621,N_1502);
and U1687 (N_1687,N_1504,N_1613);
nor U1688 (N_1688,N_1606,N_1622);
xor U1689 (N_1689,N_1603,N_1508);
or U1690 (N_1690,N_1555,N_1577);
nand U1691 (N_1691,N_1579,N_1546);
nor U1692 (N_1692,N_1525,N_1524);
xor U1693 (N_1693,N_1554,N_1588);
nor U1694 (N_1694,N_1517,N_1590);
xnor U1695 (N_1695,N_1618,N_1597);
nor U1696 (N_1696,N_1501,N_1624);
nor U1697 (N_1697,N_1531,N_1506);
or U1698 (N_1698,N_1551,N_1512);
nand U1699 (N_1699,N_1621,N_1520);
nand U1700 (N_1700,N_1607,N_1538);
nand U1701 (N_1701,N_1542,N_1598);
xnor U1702 (N_1702,N_1517,N_1601);
nor U1703 (N_1703,N_1621,N_1531);
xnor U1704 (N_1704,N_1504,N_1553);
nor U1705 (N_1705,N_1546,N_1512);
and U1706 (N_1706,N_1619,N_1567);
and U1707 (N_1707,N_1509,N_1576);
nor U1708 (N_1708,N_1592,N_1554);
nand U1709 (N_1709,N_1521,N_1504);
nand U1710 (N_1710,N_1621,N_1562);
and U1711 (N_1711,N_1576,N_1518);
nor U1712 (N_1712,N_1518,N_1623);
and U1713 (N_1713,N_1604,N_1623);
xnor U1714 (N_1714,N_1596,N_1573);
and U1715 (N_1715,N_1552,N_1512);
nand U1716 (N_1716,N_1536,N_1613);
and U1717 (N_1717,N_1622,N_1560);
nand U1718 (N_1718,N_1614,N_1547);
or U1719 (N_1719,N_1621,N_1605);
or U1720 (N_1720,N_1504,N_1538);
nand U1721 (N_1721,N_1564,N_1513);
nor U1722 (N_1722,N_1568,N_1564);
and U1723 (N_1723,N_1618,N_1607);
nand U1724 (N_1724,N_1587,N_1574);
nor U1725 (N_1725,N_1594,N_1561);
nand U1726 (N_1726,N_1621,N_1510);
nand U1727 (N_1727,N_1505,N_1500);
nor U1728 (N_1728,N_1524,N_1610);
nand U1729 (N_1729,N_1613,N_1526);
nand U1730 (N_1730,N_1549,N_1511);
nand U1731 (N_1731,N_1581,N_1592);
and U1732 (N_1732,N_1618,N_1624);
nand U1733 (N_1733,N_1569,N_1536);
nand U1734 (N_1734,N_1525,N_1581);
or U1735 (N_1735,N_1571,N_1508);
or U1736 (N_1736,N_1596,N_1503);
nand U1737 (N_1737,N_1617,N_1561);
and U1738 (N_1738,N_1614,N_1565);
nor U1739 (N_1739,N_1510,N_1599);
and U1740 (N_1740,N_1515,N_1575);
nand U1741 (N_1741,N_1606,N_1619);
or U1742 (N_1742,N_1556,N_1582);
nand U1743 (N_1743,N_1571,N_1544);
and U1744 (N_1744,N_1562,N_1567);
nor U1745 (N_1745,N_1518,N_1608);
nor U1746 (N_1746,N_1521,N_1542);
and U1747 (N_1747,N_1547,N_1550);
or U1748 (N_1748,N_1608,N_1529);
xnor U1749 (N_1749,N_1603,N_1546);
xor U1750 (N_1750,N_1727,N_1712);
or U1751 (N_1751,N_1625,N_1680);
or U1752 (N_1752,N_1636,N_1742);
xnor U1753 (N_1753,N_1658,N_1737);
xnor U1754 (N_1754,N_1630,N_1648);
and U1755 (N_1755,N_1717,N_1748);
nand U1756 (N_1756,N_1720,N_1741);
nand U1757 (N_1757,N_1651,N_1744);
nand U1758 (N_1758,N_1738,N_1694);
nand U1759 (N_1759,N_1735,N_1687);
nor U1760 (N_1760,N_1743,N_1685);
and U1761 (N_1761,N_1718,N_1682);
or U1762 (N_1762,N_1660,N_1674);
or U1763 (N_1763,N_1635,N_1628);
xor U1764 (N_1764,N_1663,N_1659);
nor U1765 (N_1765,N_1733,N_1715);
xnor U1766 (N_1766,N_1672,N_1647);
xnor U1767 (N_1767,N_1649,N_1678);
nand U1768 (N_1768,N_1637,N_1686);
and U1769 (N_1769,N_1699,N_1706);
nor U1770 (N_1770,N_1708,N_1657);
or U1771 (N_1771,N_1676,N_1656);
or U1772 (N_1772,N_1688,N_1642);
or U1773 (N_1773,N_1713,N_1725);
nand U1774 (N_1774,N_1731,N_1716);
or U1775 (N_1775,N_1721,N_1696);
nor U1776 (N_1776,N_1677,N_1700);
or U1777 (N_1777,N_1690,N_1675);
or U1778 (N_1778,N_1684,N_1638);
and U1779 (N_1779,N_1711,N_1640);
xor U1780 (N_1780,N_1736,N_1646);
nor U1781 (N_1781,N_1732,N_1655);
nand U1782 (N_1782,N_1705,N_1681);
and U1783 (N_1783,N_1726,N_1719);
nor U1784 (N_1784,N_1693,N_1661);
xnor U1785 (N_1785,N_1689,N_1734);
and U1786 (N_1786,N_1740,N_1679);
nor U1787 (N_1787,N_1667,N_1669);
nor U1788 (N_1788,N_1668,N_1643);
or U1789 (N_1789,N_1692,N_1670);
nand U1790 (N_1790,N_1666,N_1697);
and U1791 (N_1791,N_1746,N_1709);
or U1792 (N_1792,N_1641,N_1633);
nor U1793 (N_1793,N_1631,N_1654);
nor U1794 (N_1794,N_1665,N_1691);
or U1795 (N_1795,N_1745,N_1729);
or U1796 (N_1796,N_1714,N_1632);
nor U1797 (N_1797,N_1702,N_1701);
nor U1798 (N_1798,N_1722,N_1664);
nand U1799 (N_1799,N_1627,N_1629);
xnor U1800 (N_1800,N_1644,N_1626);
xor U1801 (N_1801,N_1673,N_1728);
xnor U1802 (N_1802,N_1724,N_1634);
and U1803 (N_1803,N_1723,N_1683);
and U1804 (N_1804,N_1698,N_1747);
nor U1805 (N_1805,N_1662,N_1707);
nor U1806 (N_1806,N_1639,N_1650);
or U1807 (N_1807,N_1695,N_1710);
nor U1808 (N_1808,N_1739,N_1730);
and U1809 (N_1809,N_1653,N_1645);
xnor U1810 (N_1810,N_1652,N_1704);
nand U1811 (N_1811,N_1703,N_1749);
nor U1812 (N_1812,N_1671,N_1672);
or U1813 (N_1813,N_1746,N_1748);
and U1814 (N_1814,N_1724,N_1704);
nor U1815 (N_1815,N_1744,N_1666);
and U1816 (N_1816,N_1685,N_1666);
nand U1817 (N_1817,N_1631,N_1638);
and U1818 (N_1818,N_1710,N_1705);
nand U1819 (N_1819,N_1745,N_1697);
or U1820 (N_1820,N_1719,N_1653);
and U1821 (N_1821,N_1748,N_1742);
xnor U1822 (N_1822,N_1673,N_1699);
nor U1823 (N_1823,N_1736,N_1639);
xor U1824 (N_1824,N_1693,N_1710);
or U1825 (N_1825,N_1673,N_1708);
and U1826 (N_1826,N_1706,N_1720);
nor U1827 (N_1827,N_1707,N_1697);
xor U1828 (N_1828,N_1658,N_1653);
or U1829 (N_1829,N_1716,N_1742);
and U1830 (N_1830,N_1745,N_1653);
xor U1831 (N_1831,N_1712,N_1662);
nand U1832 (N_1832,N_1680,N_1712);
nor U1833 (N_1833,N_1629,N_1733);
and U1834 (N_1834,N_1686,N_1733);
nand U1835 (N_1835,N_1637,N_1638);
nor U1836 (N_1836,N_1650,N_1660);
and U1837 (N_1837,N_1737,N_1677);
xor U1838 (N_1838,N_1667,N_1719);
and U1839 (N_1839,N_1706,N_1743);
xnor U1840 (N_1840,N_1691,N_1698);
and U1841 (N_1841,N_1728,N_1704);
or U1842 (N_1842,N_1647,N_1660);
xnor U1843 (N_1843,N_1679,N_1634);
nor U1844 (N_1844,N_1735,N_1695);
and U1845 (N_1845,N_1706,N_1649);
or U1846 (N_1846,N_1639,N_1742);
xor U1847 (N_1847,N_1714,N_1628);
and U1848 (N_1848,N_1731,N_1715);
xor U1849 (N_1849,N_1714,N_1710);
or U1850 (N_1850,N_1669,N_1657);
or U1851 (N_1851,N_1683,N_1686);
nand U1852 (N_1852,N_1641,N_1737);
nand U1853 (N_1853,N_1711,N_1684);
or U1854 (N_1854,N_1728,N_1701);
nand U1855 (N_1855,N_1650,N_1645);
nor U1856 (N_1856,N_1649,N_1675);
and U1857 (N_1857,N_1642,N_1742);
and U1858 (N_1858,N_1670,N_1747);
or U1859 (N_1859,N_1670,N_1712);
and U1860 (N_1860,N_1682,N_1698);
or U1861 (N_1861,N_1640,N_1745);
or U1862 (N_1862,N_1628,N_1625);
nand U1863 (N_1863,N_1664,N_1630);
nor U1864 (N_1864,N_1672,N_1727);
nor U1865 (N_1865,N_1738,N_1649);
and U1866 (N_1866,N_1686,N_1706);
and U1867 (N_1867,N_1641,N_1711);
nor U1868 (N_1868,N_1634,N_1747);
nor U1869 (N_1869,N_1694,N_1748);
or U1870 (N_1870,N_1696,N_1672);
xnor U1871 (N_1871,N_1702,N_1640);
nor U1872 (N_1872,N_1643,N_1706);
nand U1873 (N_1873,N_1630,N_1677);
xnor U1874 (N_1874,N_1659,N_1642);
xnor U1875 (N_1875,N_1807,N_1834);
xnor U1876 (N_1876,N_1797,N_1817);
and U1877 (N_1877,N_1811,N_1809);
and U1878 (N_1878,N_1847,N_1787);
nand U1879 (N_1879,N_1767,N_1829);
xor U1880 (N_1880,N_1815,N_1868);
nor U1881 (N_1881,N_1757,N_1803);
and U1882 (N_1882,N_1837,N_1827);
xor U1883 (N_1883,N_1862,N_1864);
and U1884 (N_1884,N_1866,N_1821);
nor U1885 (N_1885,N_1760,N_1773);
xnor U1886 (N_1886,N_1792,N_1819);
or U1887 (N_1887,N_1765,N_1857);
xnor U1888 (N_1888,N_1838,N_1808);
nand U1889 (N_1889,N_1830,N_1863);
or U1890 (N_1890,N_1799,N_1752);
xor U1891 (N_1891,N_1826,N_1790);
and U1892 (N_1892,N_1822,N_1779);
and U1893 (N_1893,N_1853,N_1854);
xnor U1894 (N_1894,N_1831,N_1820);
or U1895 (N_1895,N_1791,N_1769);
xnor U1896 (N_1896,N_1836,N_1867);
nor U1897 (N_1897,N_1781,N_1756);
nand U1898 (N_1898,N_1771,N_1849);
xor U1899 (N_1899,N_1798,N_1825);
or U1900 (N_1900,N_1845,N_1818);
nor U1901 (N_1901,N_1776,N_1758);
nand U1902 (N_1902,N_1751,N_1750);
nor U1903 (N_1903,N_1874,N_1828);
xnor U1904 (N_1904,N_1763,N_1842);
nand U1905 (N_1905,N_1786,N_1780);
nor U1906 (N_1906,N_1851,N_1761);
nand U1907 (N_1907,N_1840,N_1861);
or U1908 (N_1908,N_1843,N_1783);
xor U1909 (N_1909,N_1775,N_1806);
and U1910 (N_1910,N_1764,N_1754);
nand U1911 (N_1911,N_1832,N_1802);
nor U1912 (N_1912,N_1839,N_1841);
or U1913 (N_1913,N_1789,N_1870);
nand U1914 (N_1914,N_1782,N_1755);
xnor U1915 (N_1915,N_1848,N_1856);
nor U1916 (N_1916,N_1855,N_1778);
and U1917 (N_1917,N_1873,N_1846);
nand U1918 (N_1918,N_1860,N_1804);
xnor U1919 (N_1919,N_1872,N_1753);
and U1920 (N_1920,N_1785,N_1865);
xnor U1921 (N_1921,N_1772,N_1777);
nor U1922 (N_1922,N_1801,N_1869);
or U1923 (N_1923,N_1768,N_1796);
nand U1924 (N_1924,N_1770,N_1816);
xor U1925 (N_1925,N_1805,N_1823);
and U1926 (N_1926,N_1784,N_1759);
nand U1927 (N_1927,N_1774,N_1850);
or U1928 (N_1928,N_1835,N_1794);
and U1929 (N_1929,N_1814,N_1762);
or U1930 (N_1930,N_1871,N_1858);
or U1931 (N_1931,N_1844,N_1813);
nor U1932 (N_1932,N_1793,N_1795);
xnor U1933 (N_1933,N_1810,N_1766);
or U1934 (N_1934,N_1812,N_1800);
nor U1935 (N_1935,N_1833,N_1852);
xnor U1936 (N_1936,N_1788,N_1859);
nor U1937 (N_1937,N_1824,N_1838);
nand U1938 (N_1938,N_1823,N_1758);
nor U1939 (N_1939,N_1852,N_1815);
and U1940 (N_1940,N_1779,N_1841);
xor U1941 (N_1941,N_1753,N_1768);
or U1942 (N_1942,N_1821,N_1759);
or U1943 (N_1943,N_1871,N_1874);
and U1944 (N_1944,N_1776,N_1800);
or U1945 (N_1945,N_1816,N_1871);
nor U1946 (N_1946,N_1817,N_1755);
nor U1947 (N_1947,N_1834,N_1771);
xnor U1948 (N_1948,N_1754,N_1805);
xor U1949 (N_1949,N_1802,N_1788);
xor U1950 (N_1950,N_1792,N_1812);
and U1951 (N_1951,N_1840,N_1758);
xnor U1952 (N_1952,N_1779,N_1837);
xnor U1953 (N_1953,N_1750,N_1867);
or U1954 (N_1954,N_1768,N_1813);
or U1955 (N_1955,N_1758,N_1834);
and U1956 (N_1956,N_1860,N_1871);
nand U1957 (N_1957,N_1788,N_1838);
nor U1958 (N_1958,N_1813,N_1818);
nand U1959 (N_1959,N_1803,N_1767);
nor U1960 (N_1960,N_1807,N_1858);
xnor U1961 (N_1961,N_1778,N_1851);
nand U1962 (N_1962,N_1805,N_1853);
nor U1963 (N_1963,N_1753,N_1841);
nor U1964 (N_1964,N_1769,N_1807);
xor U1965 (N_1965,N_1768,N_1772);
xnor U1966 (N_1966,N_1845,N_1850);
or U1967 (N_1967,N_1769,N_1855);
and U1968 (N_1968,N_1807,N_1770);
xnor U1969 (N_1969,N_1806,N_1842);
xnor U1970 (N_1970,N_1765,N_1784);
nor U1971 (N_1971,N_1848,N_1762);
xnor U1972 (N_1972,N_1783,N_1800);
and U1973 (N_1973,N_1758,N_1772);
nand U1974 (N_1974,N_1784,N_1773);
xor U1975 (N_1975,N_1843,N_1767);
nand U1976 (N_1976,N_1872,N_1866);
nor U1977 (N_1977,N_1845,N_1825);
xor U1978 (N_1978,N_1823,N_1799);
xnor U1979 (N_1979,N_1869,N_1813);
nor U1980 (N_1980,N_1843,N_1785);
xnor U1981 (N_1981,N_1832,N_1853);
nand U1982 (N_1982,N_1779,N_1847);
and U1983 (N_1983,N_1765,N_1868);
xnor U1984 (N_1984,N_1834,N_1863);
and U1985 (N_1985,N_1768,N_1851);
or U1986 (N_1986,N_1763,N_1813);
xor U1987 (N_1987,N_1801,N_1775);
nor U1988 (N_1988,N_1812,N_1765);
nand U1989 (N_1989,N_1783,N_1851);
and U1990 (N_1990,N_1812,N_1798);
and U1991 (N_1991,N_1806,N_1760);
and U1992 (N_1992,N_1763,N_1799);
nor U1993 (N_1993,N_1857,N_1798);
nand U1994 (N_1994,N_1760,N_1869);
nor U1995 (N_1995,N_1831,N_1805);
and U1996 (N_1996,N_1785,N_1778);
xnor U1997 (N_1997,N_1761,N_1778);
nand U1998 (N_1998,N_1762,N_1768);
xnor U1999 (N_1999,N_1807,N_1813);
nand U2000 (N_2000,N_1965,N_1904);
and U2001 (N_2001,N_1994,N_1893);
or U2002 (N_2002,N_1946,N_1888);
nor U2003 (N_2003,N_1892,N_1922);
or U2004 (N_2004,N_1934,N_1891);
xnor U2005 (N_2005,N_1945,N_1930);
nand U2006 (N_2006,N_1913,N_1876);
nor U2007 (N_2007,N_1983,N_1931);
or U2008 (N_2008,N_1972,N_1917);
or U2009 (N_2009,N_1991,N_1995);
nor U2010 (N_2010,N_1920,N_1981);
and U2011 (N_2011,N_1921,N_1890);
xnor U2012 (N_2012,N_1967,N_1954);
or U2013 (N_2013,N_1900,N_1955);
xnor U2014 (N_2014,N_1974,N_1939);
or U2015 (N_2015,N_1950,N_1977);
nor U2016 (N_2016,N_1948,N_1951);
or U2017 (N_2017,N_1886,N_1881);
nor U2018 (N_2018,N_1949,N_1971);
and U2019 (N_2019,N_1924,N_1907);
or U2020 (N_2020,N_1889,N_1928);
xor U2021 (N_2021,N_1998,N_1993);
nand U2022 (N_2022,N_1875,N_1968);
nand U2023 (N_2023,N_1986,N_1941);
and U2024 (N_2024,N_1887,N_1897);
and U2025 (N_2025,N_1959,N_1878);
xnor U2026 (N_2026,N_1999,N_1915);
and U2027 (N_2027,N_1926,N_1990);
and U2028 (N_2028,N_1992,N_1879);
or U2029 (N_2029,N_1942,N_1957);
or U2030 (N_2030,N_1936,N_1979);
xnor U2031 (N_2031,N_1883,N_1884);
or U2032 (N_2032,N_1958,N_1982);
nand U2033 (N_2033,N_1899,N_1947);
and U2034 (N_2034,N_1961,N_1927);
nor U2035 (N_2035,N_1937,N_1970);
and U2036 (N_2036,N_1952,N_1910);
nor U2037 (N_2037,N_1901,N_1989);
nor U2038 (N_2038,N_1978,N_1969);
xnor U2039 (N_2039,N_1903,N_1996);
xor U2040 (N_2040,N_1962,N_1929);
and U2041 (N_2041,N_1964,N_1975);
and U2042 (N_2042,N_1997,N_1987);
xor U2043 (N_2043,N_1988,N_1956);
or U2044 (N_2044,N_1912,N_1919);
nor U2045 (N_2045,N_1960,N_1896);
nand U2046 (N_2046,N_1908,N_1985);
and U2047 (N_2047,N_1932,N_1895);
nand U2048 (N_2048,N_1885,N_1966);
nor U2049 (N_2049,N_1925,N_1914);
and U2050 (N_2050,N_1973,N_1944);
nor U2051 (N_2051,N_1911,N_1984);
nand U2052 (N_2052,N_1953,N_1963);
and U2053 (N_2053,N_1877,N_1935);
xor U2054 (N_2054,N_1916,N_1940);
nor U2055 (N_2055,N_1906,N_1933);
xor U2056 (N_2056,N_1905,N_1923);
xnor U2057 (N_2057,N_1909,N_1902);
xnor U2058 (N_2058,N_1880,N_1976);
or U2059 (N_2059,N_1938,N_1898);
nand U2060 (N_2060,N_1918,N_1980);
nor U2061 (N_2061,N_1894,N_1882);
nand U2062 (N_2062,N_1943,N_1885);
nor U2063 (N_2063,N_1886,N_1949);
nor U2064 (N_2064,N_1939,N_1946);
and U2065 (N_2065,N_1981,N_1910);
nand U2066 (N_2066,N_1920,N_1926);
xor U2067 (N_2067,N_1911,N_1976);
and U2068 (N_2068,N_1925,N_1904);
xnor U2069 (N_2069,N_1920,N_1880);
and U2070 (N_2070,N_1882,N_1907);
nor U2071 (N_2071,N_1998,N_1986);
and U2072 (N_2072,N_1990,N_1921);
nor U2073 (N_2073,N_1893,N_1997);
nor U2074 (N_2074,N_1915,N_1975);
nor U2075 (N_2075,N_1986,N_1917);
nor U2076 (N_2076,N_1906,N_1969);
and U2077 (N_2077,N_1895,N_1884);
or U2078 (N_2078,N_1968,N_1969);
or U2079 (N_2079,N_1955,N_1919);
nor U2080 (N_2080,N_1993,N_1926);
and U2081 (N_2081,N_1881,N_1986);
nor U2082 (N_2082,N_1899,N_1973);
xnor U2083 (N_2083,N_1906,N_1907);
xor U2084 (N_2084,N_1875,N_1995);
or U2085 (N_2085,N_1947,N_1969);
and U2086 (N_2086,N_1906,N_1903);
xor U2087 (N_2087,N_1952,N_1959);
nand U2088 (N_2088,N_1909,N_1899);
and U2089 (N_2089,N_1947,N_1987);
xnor U2090 (N_2090,N_1931,N_1876);
nor U2091 (N_2091,N_1989,N_1921);
nor U2092 (N_2092,N_1983,N_1981);
and U2093 (N_2093,N_1980,N_1916);
and U2094 (N_2094,N_1947,N_1910);
nor U2095 (N_2095,N_1929,N_1923);
and U2096 (N_2096,N_1970,N_1993);
nor U2097 (N_2097,N_1936,N_1912);
or U2098 (N_2098,N_1884,N_1966);
nand U2099 (N_2099,N_1897,N_1900);
nor U2100 (N_2100,N_1878,N_1984);
nand U2101 (N_2101,N_1943,N_1977);
and U2102 (N_2102,N_1928,N_1900);
or U2103 (N_2103,N_1934,N_1935);
and U2104 (N_2104,N_1980,N_1930);
nor U2105 (N_2105,N_1944,N_1882);
or U2106 (N_2106,N_1883,N_1973);
and U2107 (N_2107,N_1985,N_1921);
and U2108 (N_2108,N_1949,N_1957);
xnor U2109 (N_2109,N_1965,N_1893);
xor U2110 (N_2110,N_1943,N_1945);
nor U2111 (N_2111,N_1889,N_1954);
or U2112 (N_2112,N_1934,N_1877);
and U2113 (N_2113,N_1932,N_1901);
nand U2114 (N_2114,N_1926,N_1942);
or U2115 (N_2115,N_1895,N_1982);
and U2116 (N_2116,N_1920,N_1911);
or U2117 (N_2117,N_1916,N_1883);
or U2118 (N_2118,N_1981,N_1935);
nor U2119 (N_2119,N_1990,N_1976);
and U2120 (N_2120,N_1893,N_1945);
or U2121 (N_2121,N_1961,N_1911);
and U2122 (N_2122,N_1919,N_1961);
nor U2123 (N_2123,N_1921,N_1919);
or U2124 (N_2124,N_1980,N_1968);
nor U2125 (N_2125,N_2091,N_2108);
nand U2126 (N_2126,N_2047,N_2070);
xnor U2127 (N_2127,N_2037,N_2004);
or U2128 (N_2128,N_2112,N_2102);
xnor U2129 (N_2129,N_2022,N_2040);
and U2130 (N_2130,N_2012,N_2113);
nand U2131 (N_2131,N_2018,N_2034);
nor U2132 (N_2132,N_2065,N_2080);
and U2133 (N_2133,N_2021,N_2031);
or U2134 (N_2134,N_2086,N_2024);
xor U2135 (N_2135,N_2089,N_2050);
nand U2136 (N_2136,N_2038,N_2001);
and U2137 (N_2137,N_2105,N_2119);
nor U2138 (N_2138,N_2107,N_2093);
xor U2139 (N_2139,N_2058,N_2109);
or U2140 (N_2140,N_2114,N_2039);
and U2141 (N_2141,N_2095,N_2059);
nand U2142 (N_2142,N_2096,N_2009);
and U2143 (N_2143,N_2100,N_2072);
and U2144 (N_2144,N_2000,N_2120);
and U2145 (N_2145,N_2116,N_2055);
nor U2146 (N_2146,N_2013,N_2076);
or U2147 (N_2147,N_2068,N_2062);
nand U2148 (N_2148,N_2085,N_2002);
nand U2149 (N_2149,N_2008,N_2081);
and U2150 (N_2150,N_2075,N_2073);
nor U2151 (N_2151,N_2099,N_2051);
and U2152 (N_2152,N_2019,N_2123);
and U2153 (N_2153,N_2117,N_2029);
nor U2154 (N_2154,N_2005,N_2124);
and U2155 (N_2155,N_2097,N_2111);
or U2156 (N_2156,N_2044,N_2011);
xnor U2157 (N_2157,N_2049,N_2042);
or U2158 (N_2158,N_2084,N_2071);
nor U2159 (N_2159,N_2007,N_2006);
and U2160 (N_2160,N_2069,N_2079);
nand U2161 (N_2161,N_2027,N_2017);
and U2162 (N_2162,N_2028,N_2048);
or U2163 (N_2163,N_2035,N_2064);
and U2164 (N_2164,N_2063,N_2030);
xnor U2165 (N_2165,N_2121,N_2110);
nand U2166 (N_2166,N_2098,N_2032);
xor U2167 (N_2167,N_2052,N_2061);
or U2168 (N_2168,N_2067,N_2016);
and U2169 (N_2169,N_2033,N_2056);
or U2170 (N_2170,N_2045,N_2041);
xnor U2171 (N_2171,N_2043,N_2103);
or U2172 (N_2172,N_2106,N_2092);
and U2173 (N_2173,N_2101,N_2122);
and U2174 (N_2174,N_2083,N_2088);
and U2175 (N_2175,N_2003,N_2025);
nor U2176 (N_2176,N_2087,N_2115);
and U2177 (N_2177,N_2066,N_2026);
nand U2178 (N_2178,N_2015,N_2060);
and U2179 (N_2179,N_2094,N_2054);
nor U2180 (N_2180,N_2036,N_2074);
nand U2181 (N_2181,N_2077,N_2082);
nor U2182 (N_2182,N_2078,N_2020);
or U2183 (N_2183,N_2057,N_2010);
or U2184 (N_2184,N_2046,N_2014);
nand U2185 (N_2185,N_2104,N_2053);
and U2186 (N_2186,N_2118,N_2023);
nor U2187 (N_2187,N_2090,N_2023);
nor U2188 (N_2188,N_2109,N_2008);
nor U2189 (N_2189,N_2108,N_2048);
nand U2190 (N_2190,N_2120,N_2075);
or U2191 (N_2191,N_2010,N_2077);
xor U2192 (N_2192,N_2080,N_2021);
xnor U2193 (N_2193,N_2014,N_2055);
or U2194 (N_2194,N_2042,N_2079);
nor U2195 (N_2195,N_2059,N_2070);
and U2196 (N_2196,N_2017,N_2033);
nand U2197 (N_2197,N_2013,N_2001);
nor U2198 (N_2198,N_2074,N_2035);
or U2199 (N_2199,N_2102,N_2010);
xor U2200 (N_2200,N_2039,N_2122);
nand U2201 (N_2201,N_2033,N_2026);
nand U2202 (N_2202,N_2069,N_2102);
and U2203 (N_2203,N_2038,N_2035);
xor U2204 (N_2204,N_2051,N_2066);
xnor U2205 (N_2205,N_2103,N_2030);
nand U2206 (N_2206,N_2062,N_2076);
or U2207 (N_2207,N_2109,N_2068);
nor U2208 (N_2208,N_2025,N_2000);
xnor U2209 (N_2209,N_2083,N_2073);
or U2210 (N_2210,N_2064,N_2092);
and U2211 (N_2211,N_2097,N_2078);
and U2212 (N_2212,N_2108,N_2025);
xnor U2213 (N_2213,N_2055,N_2074);
or U2214 (N_2214,N_2089,N_2059);
or U2215 (N_2215,N_2070,N_2121);
nand U2216 (N_2216,N_2084,N_2070);
or U2217 (N_2217,N_2004,N_2062);
or U2218 (N_2218,N_2048,N_2003);
xor U2219 (N_2219,N_2012,N_2017);
xnor U2220 (N_2220,N_2034,N_2095);
or U2221 (N_2221,N_2116,N_2121);
nand U2222 (N_2222,N_2013,N_2101);
nand U2223 (N_2223,N_2038,N_2112);
and U2224 (N_2224,N_2083,N_2001);
or U2225 (N_2225,N_2083,N_2042);
and U2226 (N_2226,N_2094,N_2111);
nor U2227 (N_2227,N_2045,N_2100);
and U2228 (N_2228,N_2063,N_2073);
nor U2229 (N_2229,N_2121,N_2065);
nor U2230 (N_2230,N_2120,N_2089);
nand U2231 (N_2231,N_2059,N_2103);
nor U2232 (N_2232,N_2090,N_2054);
or U2233 (N_2233,N_2003,N_2109);
or U2234 (N_2234,N_2091,N_2058);
nand U2235 (N_2235,N_2070,N_2045);
nand U2236 (N_2236,N_2057,N_2051);
xor U2237 (N_2237,N_2007,N_2065);
or U2238 (N_2238,N_2078,N_2061);
or U2239 (N_2239,N_2040,N_2054);
or U2240 (N_2240,N_2086,N_2062);
and U2241 (N_2241,N_2123,N_2028);
or U2242 (N_2242,N_2000,N_2057);
or U2243 (N_2243,N_2067,N_2063);
and U2244 (N_2244,N_2090,N_2056);
xnor U2245 (N_2245,N_2041,N_2090);
and U2246 (N_2246,N_2037,N_2117);
xnor U2247 (N_2247,N_2116,N_2063);
xnor U2248 (N_2248,N_2026,N_2058);
nor U2249 (N_2249,N_2080,N_2110);
xnor U2250 (N_2250,N_2219,N_2167);
nand U2251 (N_2251,N_2143,N_2214);
and U2252 (N_2252,N_2128,N_2220);
nand U2253 (N_2253,N_2247,N_2157);
or U2254 (N_2254,N_2237,N_2190);
xor U2255 (N_2255,N_2147,N_2195);
nand U2256 (N_2256,N_2154,N_2192);
and U2257 (N_2257,N_2194,N_2131);
xnor U2258 (N_2258,N_2229,N_2235);
and U2259 (N_2259,N_2156,N_2199);
or U2260 (N_2260,N_2197,N_2221);
and U2261 (N_2261,N_2243,N_2232);
xor U2262 (N_2262,N_2240,N_2225);
xor U2263 (N_2263,N_2149,N_2127);
and U2264 (N_2264,N_2152,N_2168);
or U2265 (N_2265,N_2171,N_2129);
xor U2266 (N_2266,N_2153,N_2148);
and U2267 (N_2267,N_2215,N_2165);
xor U2268 (N_2268,N_2205,N_2233);
nand U2269 (N_2269,N_2142,N_2151);
xor U2270 (N_2270,N_2198,N_2177);
xor U2271 (N_2271,N_2180,N_2238);
or U2272 (N_2272,N_2242,N_2174);
xnor U2273 (N_2273,N_2136,N_2126);
nand U2274 (N_2274,N_2163,N_2227);
and U2275 (N_2275,N_2223,N_2150);
nor U2276 (N_2276,N_2155,N_2201);
xor U2277 (N_2277,N_2135,N_2211);
or U2278 (N_2278,N_2169,N_2133);
nand U2279 (N_2279,N_2207,N_2204);
or U2280 (N_2280,N_2183,N_2184);
and U2281 (N_2281,N_2212,N_2141);
nor U2282 (N_2282,N_2179,N_2213);
and U2283 (N_2283,N_2160,N_2226);
or U2284 (N_2284,N_2228,N_2134);
xnor U2285 (N_2285,N_2178,N_2132);
nor U2286 (N_2286,N_2188,N_2216);
nand U2287 (N_2287,N_2203,N_2248);
nand U2288 (N_2288,N_2245,N_2170);
or U2289 (N_2289,N_2196,N_2217);
xor U2290 (N_2290,N_2159,N_2172);
or U2291 (N_2291,N_2202,N_2182);
nand U2292 (N_2292,N_2208,N_2185);
or U2293 (N_2293,N_2166,N_2145);
and U2294 (N_2294,N_2246,N_2137);
or U2295 (N_2295,N_2210,N_2146);
xnor U2296 (N_2296,N_2144,N_2230);
nor U2297 (N_2297,N_2191,N_2222);
and U2298 (N_2298,N_2181,N_2234);
nand U2299 (N_2299,N_2173,N_2206);
and U2300 (N_2300,N_2231,N_2161);
or U2301 (N_2301,N_2186,N_2158);
xnor U2302 (N_2302,N_2218,N_2164);
nand U2303 (N_2303,N_2139,N_2239);
and U2304 (N_2304,N_2189,N_2162);
nand U2305 (N_2305,N_2187,N_2130);
nand U2306 (N_2306,N_2236,N_2200);
nand U2307 (N_2307,N_2138,N_2241);
nand U2308 (N_2308,N_2209,N_2224);
xor U2309 (N_2309,N_2140,N_2176);
and U2310 (N_2310,N_2175,N_2125);
and U2311 (N_2311,N_2193,N_2249);
nand U2312 (N_2312,N_2244,N_2137);
nand U2313 (N_2313,N_2228,N_2227);
nor U2314 (N_2314,N_2226,N_2140);
and U2315 (N_2315,N_2230,N_2182);
and U2316 (N_2316,N_2185,N_2218);
nor U2317 (N_2317,N_2228,N_2197);
or U2318 (N_2318,N_2195,N_2155);
nor U2319 (N_2319,N_2156,N_2169);
nor U2320 (N_2320,N_2226,N_2188);
nand U2321 (N_2321,N_2211,N_2126);
and U2322 (N_2322,N_2206,N_2189);
xnor U2323 (N_2323,N_2226,N_2206);
xor U2324 (N_2324,N_2151,N_2236);
or U2325 (N_2325,N_2186,N_2189);
nand U2326 (N_2326,N_2144,N_2199);
nor U2327 (N_2327,N_2180,N_2127);
nand U2328 (N_2328,N_2215,N_2232);
or U2329 (N_2329,N_2162,N_2180);
nor U2330 (N_2330,N_2219,N_2243);
or U2331 (N_2331,N_2234,N_2224);
nor U2332 (N_2332,N_2127,N_2179);
nor U2333 (N_2333,N_2136,N_2196);
and U2334 (N_2334,N_2136,N_2207);
or U2335 (N_2335,N_2126,N_2132);
xnor U2336 (N_2336,N_2146,N_2204);
xnor U2337 (N_2337,N_2155,N_2213);
and U2338 (N_2338,N_2128,N_2169);
and U2339 (N_2339,N_2156,N_2211);
xor U2340 (N_2340,N_2127,N_2198);
and U2341 (N_2341,N_2239,N_2198);
or U2342 (N_2342,N_2181,N_2247);
xor U2343 (N_2343,N_2151,N_2210);
or U2344 (N_2344,N_2224,N_2125);
or U2345 (N_2345,N_2246,N_2133);
nand U2346 (N_2346,N_2167,N_2214);
or U2347 (N_2347,N_2232,N_2248);
xnor U2348 (N_2348,N_2247,N_2135);
xor U2349 (N_2349,N_2246,N_2197);
or U2350 (N_2350,N_2237,N_2134);
xnor U2351 (N_2351,N_2153,N_2217);
nand U2352 (N_2352,N_2145,N_2244);
nor U2353 (N_2353,N_2231,N_2202);
or U2354 (N_2354,N_2132,N_2247);
nand U2355 (N_2355,N_2215,N_2133);
or U2356 (N_2356,N_2162,N_2210);
xnor U2357 (N_2357,N_2199,N_2146);
or U2358 (N_2358,N_2209,N_2180);
nor U2359 (N_2359,N_2210,N_2240);
nor U2360 (N_2360,N_2164,N_2157);
nor U2361 (N_2361,N_2236,N_2246);
or U2362 (N_2362,N_2162,N_2152);
xor U2363 (N_2363,N_2204,N_2191);
nand U2364 (N_2364,N_2241,N_2202);
nand U2365 (N_2365,N_2148,N_2181);
nand U2366 (N_2366,N_2236,N_2180);
nor U2367 (N_2367,N_2135,N_2219);
nor U2368 (N_2368,N_2200,N_2241);
or U2369 (N_2369,N_2136,N_2202);
nand U2370 (N_2370,N_2135,N_2217);
xor U2371 (N_2371,N_2214,N_2127);
and U2372 (N_2372,N_2216,N_2137);
or U2373 (N_2373,N_2126,N_2146);
or U2374 (N_2374,N_2189,N_2191);
or U2375 (N_2375,N_2371,N_2347);
or U2376 (N_2376,N_2292,N_2304);
nand U2377 (N_2377,N_2287,N_2300);
xnor U2378 (N_2378,N_2291,N_2261);
xor U2379 (N_2379,N_2281,N_2363);
and U2380 (N_2380,N_2301,N_2266);
nor U2381 (N_2381,N_2359,N_2367);
xor U2382 (N_2382,N_2361,N_2267);
nor U2383 (N_2383,N_2336,N_2271);
and U2384 (N_2384,N_2268,N_2330);
xor U2385 (N_2385,N_2370,N_2295);
nor U2386 (N_2386,N_2286,N_2358);
nand U2387 (N_2387,N_2319,N_2323);
nor U2388 (N_2388,N_2256,N_2345);
nand U2389 (N_2389,N_2298,N_2368);
nor U2390 (N_2390,N_2307,N_2269);
and U2391 (N_2391,N_2275,N_2333);
xor U2392 (N_2392,N_2284,N_2348);
nand U2393 (N_2393,N_2343,N_2313);
nand U2394 (N_2394,N_2369,N_2290);
nor U2395 (N_2395,N_2356,N_2342);
xnor U2396 (N_2396,N_2278,N_2344);
or U2397 (N_2397,N_2276,N_2351);
nor U2398 (N_2398,N_2337,N_2353);
nand U2399 (N_2399,N_2263,N_2255);
or U2400 (N_2400,N_2360,N_2331);
nor U2401 (N_2401,N_2254,N_2325);
nor U2402 (N_2402,N_2277,N_2280);
nor U2403 (N_2403,N_2322,N_2314);
and U2404 (N_2404,N_2315,N_2366);
xor U2405 (N_2405,N_2309,N_2365);
nor U2406 (N_2406,N_2334,N_2299);
nor U2407 (N_2407,N_2262,N_2357);
xnor U2408 (N_2408,N_2346,N_2354);
nor U2409 (N_2409,N_2318,N_2253);
xnor U2410 (N_2410,N_2339,N_2282);
or U2411 (N_2411,N_2311,N_2296);
and U2412 (N_2412,N_2335,N_2329);
xor U2413 (N_2413,N_2285,N_2312);
nor U2414 (N_2414,N_2373,N_2279);
xnor U2415 (N_2415,N_2372,N_2274);
nand U2416 (N_2416,N_2364,N_2257);
and U2417 (N_2417,N_2324,N_2264);
nand U2418 (N_2418,N_2260,N_2306);
and U2419 (N_2419,N_2328,N_2250);
nand U2420 (N_2420,N_2316,N_2270);
nand U2421 (N_2421,N_2349,N_2352);
nor U2422 (N_2422,N_2251,N_2303);
and U2423 (N_2423,N_2327,N_2338);
nor U2424 (N_2424,N_2374,N_2362);
or U2425 (N_2425,N_2294,N_2321);
or U2426 (N_2426,N_2310,N_2297);
or U2427 (N_2427,N_2320,N_2305);
and U2428 (N_2428,N_2332,N_2341);
nor U2429 (N_2429,N_2265,N_2258);
or U2430 (N_2430,N_2302,N_2293);
or U2431 (N_2431,N_2355,N_2252);
nand U2432 (N_2432,N_2283,N_2340);
nand U2433 (N_2433,N_2308,N_2289);
xor U2434 (N_2434,N_2273,N_2317);
nor U2435 (N_2435,N_2272,N_2259);
nor U2436 (N_2436,N_2326,N_2350);
nor U2437 (N_2437,N_2288,N_2301);
and U2438 (N_2438,N_2311,N_2279);
nand U2439 (N_2439,N_2326,N_2324);
xnor U2440 (N_2440,N_2288,N_2354);
or U2441 (N_2441,N_2254,N_2292);
nand U2442 (N_2442,N_2365,N_2284);
xnor U2443 (N_2443,N_2292,N_2349);
and U2444 (N_2444,N_2254,N_2253);
and U2445 (N_2445,N_2295,N_2302);
nor U2446 (N_2446,N_2327,N_2326);
or U2447 (N_2447,N_2358,N_2370);
and U2448 (N_2448,N_2362,N_2289);
and U2449 (N_2449,N_2308,N_2288);
or U2450 (N_2450,N_2329,N_2306);
nor U2451 (N_2451,N_2332,N_2314);
nor U2452 (N_2452,N_2277,N_2274);
and U2453 (N_2453,N_2322,N_2323);
nor U2454 (N_2454,N_2364,N_2277);
nor U2455 (N_2455,N_2335,N_2359);
xnor U2456 (N_2456,N_2360,N_2307);
nand U2457 (N_2457,N_2276,N_2364);
xor U2458 (N_2458,N_2297,N_2352);
and U2459 (N_2459,N_2262,N_2295);
and U2460 (N_2460,N_2339,N_2290);
nand U2461 (N_2461,N_2345,N_2332);
or U2462 (N_2462,N_2302,N_2281);
and U2463 (N_2463,N_2329,N_2289);
xor U2464 (N_2464,N_2294,N_2267);
xnor U2465 (N_2465,N_2351,N_2250);
nor U2466 (N_2466,N_2284,N_2335);
nor U2467 (N_2467,N_2372,N_2371);
or U2468 (N_2468,N_2364,N_2335);
xor U2469 (N_2469,N_2359,N_2290);
xor U2470 (N_2470,N_2277,N_2256);
or U2471 (N_2471,N_2316,N_2325);
xnor U2472 (N_2472,N_2295,N_2312);
nand U2473 (N_2473,N_2251,N_2370);
nand U2474 (N_2474,N_2344,N_2279);
nor U2475 (N_2475,N_2279,N_2267);
xor U2476 (N_2476,N_2288,N_2318);
nand U2477 (N_2477,N_2351,N_2315);
and U2478 (N_2478,N_2291,N_2290);
and U2479 (N_2479,N_2269,N_2323);
nand U2480 (N_2480,N_2316,N_2342);
nor U2481 (N_2481,N_2276,N_2352);
nand U2482 (N_2482,N_2350,N_2305);
nor U2483 (N_2483,N_2351,N_2272);
or U2484 (N_2484,N_2255,N_2365);
or U2485 (N_2485,N_2307,N_2304);
xnor U2486 (N_2486,N_2314,N_2321);
or U2487 (N_2487,N_2303,N_2324);
or U2488 (N_2488,N_2309,N_2290);
and U2489 (N_2489,N_2323,N_2252);
xnor U2490 (N_2490,N_2279,N_2367);
nand U2491 (N_2491,N_2350,N_2320);
nor U2492 (N_2492,N_2250,N_2359);
xor U2493 (N_2493,N_2347,N_2271);
nand U2494 (N_2494,N_2313,N_2315);
nand U2495 (N_2495,N_2304,N_2270);
or U2496 (N_2496,N_2336,N_2315);
and U2497 (N_2497,N_2257,N_2359);
and U2498 (N_2498,N_2311,N_2330);
and U2499 (N_2499,N_2317,N_2334);
xor U2500 (N_2500,N_2461,N_2425);
xnor U2501 (N_2501,N_2402,N_2454);
nand U2502 (N_2502,N_2403,N_2422);
nand U2503 (N_2503,N_2457,N_2383);
xnor U2504 (N_2504,N_2441,N_2445);
nor U2505 (N_2505,N_2410,N_2452);
and U2506 (N_2506,N_2380,N_2492);
nand U2507 (N_2507,N_2427,N_2473);
xnor U2508 (N_2508,N_2419,N_2417);
or U2509 (N_2509,N_2499,N_2399);
or U2510 (N_2510,N_2389,N_2375);
and U2511 (N_2511,N_2409,N_2448);
xor U2512 (N_2512,N_2485,N_2450);
nor U2513 (N_2513,N_2401,N_2381);
or U2514 (N_2514,N_2479,N_2416);
nand U2515 (N_2515,N_2376,N_2426);
xor U2516 (N_2516,N_2434,N_2446);
xor U2517 (N_2517,N_2379,N_2435);
and U2518 (N_2518,N_2405,N_2394);
and U2519 (N_2519,N_2391,N_2397);
nand U2520 (N_2520,N_2487,N_2476);
and U2521 (N_2521,N_2398,N_2486);
xnor U2522 (N_2522,N_2498,N_2431);
nand U2523 (N_2523,N_2449,N_2474);
and U2524 (N_2524,N_2411,N_2404);
nor U2525 (N_2525,N_2463,N_2413);
or U2526 (N_2526,N_2493,N_2482);
or U2527 (N_2527,N_2384,N_2386);
nand U2528 (N_2528,N_2407,N_2400);
nor U2529 (N_2529,N_2390,N_2388);
and U2530 (N_2530,N_2443,N_2478);
nand U2531 (N_2531,N_2387,N_2393);
or U2532 (N_2532,N_2494,N_2464);
nor U2533 (N_2533,N_2423,N_2440);
xnor U2534 (N_2534,N_2472,N_2438);
nand U2535 (N_2535,N_2469,N_2475);
xnor U2536 (N_2536,N_2483,N_2458);
nand U2537 (N_2537,N_2421,N_2432);
nor U2538 (N_2538,N_2451,N_2471);
nor U2539 (N_2539,N_2382,N_2496);
and U2540 (N_2540,N_2395,N_2385);
nand U2541 (N_2541,N_2453,N_2490);
or U2542 (N_2542,N_2488,N_2459);
nor U2543 (N_2543,N_2424,N_2439);
and U2544 (N_2544,N_2442,N_2433);
nor U2545 (N_2545,N_2430,N_2481);
xnor U2546 (N_2546,N_2489,N_2462);
nor U2547 (N_2547,N_2447,N_2480);
nand U2548 (N_2548,N_2396,N_2418);
xnor U2549 (N_2549,N_2436,N_2412);
xor U2550 (N_2550,N_2466,N_2495);
or U2551 (N_2551,N_2414,N_2444);
nor U2552 (N_2552,N_2491,N_2484);
and U2553 (N_2553,N_2468,N_2455);
xor U2554 (N_2554,N_2429,N_2470);
nor U2555 (N_2555,N_2408,N_2420);
xor U2556 (N_2556,N_2477,N_2460);
and U2557 (N_2557,N_2415,N_2428);
and U2558 (N_2558,N_2377,N_2406);
or U2559 (N_2559,N_2392,N_2465);
and U2560 (N_2560,N_2497,N_2456);
and U2561 (N_2561,N_2437,N_2467);
nor U2562 (N_2562,N_2378,N_2467);
and U2563 (N_2563,N_2392,N_2481);
nand U2564 (N_2564,N_2459,N_2402);
nor U2565 (N_2565,N_2443,N_2453);
and U2566 (N_2566,N_2475,N_2391);
xnor U2567 (N_2567,N_2486,N_2411);
and U2568 (N_2568,N_2383,N_2498);
nand U2569 (N_2569,N_2490,N_2471);
or U2570 (N_2570,N_2434,N_2410);
xor U2571 (N_2571,N_2462,N_2434);
or U2572 (N_2572,N_2409,N_2457);
xor U2573 (N_2573,N_2417,N_2404);
nor U2574 (N_2574,N_2396,N_2460);
nand U2575 (N_2575,N_2418,N_2481);
xor U2576 (N_2576,N_2454,N_2417);
nor U2577 (N_2577,N_2466,N_2470);
nand U2578 (N_2578,N_2468,N_2425);
and U2579 (N_2579,N_2394,N_2420);
xor U2580 (N_2580,N_2461,N_2411);
nand U2581 (N_2581,N_2461,N_2426);
or U2582 (N_2582,N_2378,N_2458);
nand U2583 (N_2583,N_2379,N_2426);
and U2584 (N_2584,N_2402,N_2378);
nand U2585 (N_2585,N_2496,N_2458);
nand U2586 (N_2586,N_2399,N_2418);
xnor U2587 (N_2587,N_2413,N_2390);
nand U2588 (N_2588,N_2450,N_2427);
nor U2589 (N_2589,N_2426,N_2405);
and U2590 (N_2590,N_2438,N_2452);
nand U2591 (N_2591,N_2436,N_2423);
or U2592 (N_2592,N_2460,N_2445);
or U2593 (N_2593,N_2453,N_2482);
and U2594 (N_2594,N_2401,N_2426);
nor U2595 (N_2595,N_2458,N_2434);
and U2596 (N_2596,N_2417,N_2486);
or U2597 (N_2597,N_2377,N_2402);
nor U2598 (N_2598,N_2386,N_2405);
xnor U2599 (N_2599,N_2432,N_2446);
and U2600 (N_2600,N_2432,N_2403);
nand U2601 (N_2601,N_2398,N_2455);
nor U2602 (N_2602,N_2375,N_2478);
or U2603 (N_2603,N_2483,N_2409);
nand U2604 (N_2604,N_2405,N_2423);
or U2605 (N_2605,N_2481,N_2484);
xor U2606 (N_2606,N_2490,N_2498);
xor U2607 (N_2607,N_2448,N_2467);
nor U2608 (N_2608,N_2403,N_2451);
or U2609 (N_2609,N_2484,N_2465);
and U2610 (N_2610,N_2466,N_2404);
xor U2611 (N_2611,N_2383,N_2424);
xor U2612 (N_2612,N_2461,N_2387);
or U2613 (N_2613,N_2450,N_2489);
nand U2614 (N_2614,N_2400,N_2406);
or U2615 (N_2615,N_2457,N_2377);
and U2616 (N_2616,N_2450,N_2429);
nand U2617 (N_2617,N_2455,N_2473);
nand U2618 (N_2618,N_2455,N_2447);
xnor U2619 (N_2619,N_2380,N_2391);
xor U2620 (N_2620,N_2477,N_2430);
nand U2621 (N_2621,N_2397,N_2498);
and U2622 (N_2622,N_2491,N_2420);
and U2623 (N_2623,N_2436,N_2497);
nand U2624 (N_2624,N_2456,N_2384);
nand U2625 (N_2625,N_2575,N_2550);
nor U2626 (N_2626,N_2614,N_2606);
nor U2627 (N_2627,N_2610,N_2539);
nor U2628 (N_2628,N_2583,N_2594);
xor U2629 (N_2629,N_2566,N_2522);
nand U2630 (N_2630,N_2555,N_2615);
nand U2631 (N_2631,N_2565,N_2556);
nand U2632 (N_2632,N_2502,N_2611);
xnor U2633 (N_2633,N_2616,N_2609);
nor U2634 (N_2634,N_2524,N_2536);
nor U2635 (N_2635,N_2603,N_2588);
nor U2636 (N_2636,N_2505,N_2532);
nand U2637 (N_2637,N_2595,N_2604);
xor U2638 (N_2638,N_2562,N_2618);
or U2639 (N_2639,N_2589,N_2548);
nand U2640 (N_2640,N_2518,N_2520);
nor U2641 (N_2641,N_2587,N_2612);
and U2642 (N_2642,N_2602,N_2582);
xor U2643 (N_2643,N_2507,N_2531);
xnor U2644 (N_2644,N_2503,N_2601);
nand U2645 (N_2645,N_2546,N_2534);
and U2646 (N_2646,N_2519,N_2596);
xnor U2647 (N_2647,N_2513,N_2511);
nand U2648 (N_2648,N_2574,N_2598);
and U2649 (N_2649,N_2576,N_2500);
nand U2650 (N_2650,N_2591,N_2553);
nand U2651 (N_2651,N_2542,N_2581);
nand U2652 (N_2652,N_2559,N_2577);
or U2653 (N_2653,N_2563,N_2558);
or U2654 (N_2654,N_2564,N_2620);
and U2655 (N_2655,N_2549,N_2585);
xor U2656 (N_2656,N_2557,N_2607);
and U2657 (N_2657,N_2540,N_2521);
and U2658 (N_2658,N_2597,N_2608);
and U2659 (N_2659,N_2569,N_2623);
nand U2660 (N_2660,N_2568,N_2537);
nand U2661 (N_2661,N_2624,N_2501);
nand U2662 (N_2662,N_2529,N_2523);
and U2663 (N_2663,N_2516,N_2592);
xor U2664 (N_2664,N_2619,N_2605);
and U2665 (N_2665,N_2528,N_2573);
nor U2666 (N_2666,N_2506,N_2580);
nor U2667 (N_2667,N_2533,N_2541);
xnor U2668 (N_2668,N_2552,N_2547);
and U2669 (N_2669,N_2526,N_2525);
and U2670 (N_2670,N_2504,N_2545);
or U2671 (N_2671,N_2515,N_2570);
and U2672 (N_2672,N_2512,N_2593);
and U2673 (N_2673,N_2578,N_2561);
and U2674 (N_2674,N_2599,N_2567);
nor U2675 (N_2675,N_2560,N_2514);
nand U2676 (N_2676,N_2510,N_2584);
and U2677 (N_2677,N_2543,N_2551);
or U2678 (N_2678,N_2535,N_2613);
or U2679 (N_2679,N_2572,N_2544);
and U2680 (N_2680,N_2517,N_2508);
nor U2681 (N_2681,N_2600,N_2571);
xor U2682 (N_2682,N_2586,N_2509);
xnor U2683 (N_2683,N_2538,N_2621);
nand U2684 (N_2684,N_2579,N_2590);
nor U2685 (N_2685,N_2617,N_2530);
or U2686 (N_2686,N_2527,N_2554);
nor U2687 (N_2687,N_2622,N_2593);
nor U2688 (N_2688,N_2530,N_2513);
or U2689 (N_2689,N_2596,N_2593);
or U2690 (N_2690,N_2528,N_2544);
nor U2691 (N_2691,N_2620,N_2558);
and U2692 (N_2692,N_2530,N_2608);
nor U2693 (N_2693,N_2530,N_2603);
or U2694 (N_2694,N_2566,N_2592);
and U2695 (N_2695,N_2602,N_2511);
xor U2696 (N_2696,N_2592,N_2601);
nand U2697 (N_2697,N_2618,N_2616);
xor U2698 (N_2698,N_2535,N_2568);
nor U2699 (N_2699,N_2582,N_2585);
xnor U2700 (N_2700,N_2527,N_2558);
nor U2701 (N_2701,N_2544,N_2619);
xnor U2702 (N_2702,N_2546,N_2619);
nand U2703 (N_2703,N_2574,N_2540);
and U2704 (N_2704,N_2562,N_2500);
xor U2705 (N_2705,N_2589,N_2518);
or U2706 (N_2706,N_2554,N_2617);
nor U2707 (N_2707,N_2559,N_2566);
and U2708 (N_2708,N_2559,N_2512);
or U2709 (N_2709,N_2623,N_2548);
nand U2710 (N_2710,N_2537,N_2538);
xnor U2711 (N_2711,N_2573,N_2523);
nand U2712 (N_2712,N_2507,N_2585);
or U2713 (N_2713,N_2620,N_2595);
xor U2714 (N_2714,N_2591,N_2584);
xnor U2715 (N_2715,N_2526,N_2619);
xnor U2716 (N_2716,N_2601,N_2506);
xor U2717 (N_2717,N_2594,N_2501);
nor U2718 (N_2718,N_2563,N_2578);
and U2719 (N_2719,N_2535,N_2536);
and U2720 (N_2720,N_2530,N_2575);
xnor U2721 (N_2721,N_2526,N_2559);
nor U2722 (N_2722,N_2569,N_2592);
xnor U2723 (N_2723,N_2576,N_2586);
xnor U2724 (N_2724,N_2514,N_2523);
nor U2725 (N_2725,N_2567,N_2501);
xor U2726 (N_2726,N_2549,N_2603);
xnor U2727 (N_2727,N_2579,N_2538);
nand U2728 (N_2728,N_2586,N_2580);
or U2729 (N_2729,N_2557,N_2554);
nor U2730 (N_2730,N_2507,N_2542);
nor U2731 (N_2731,N_2611,N_2528);
nand U2732 (N_2732,N_2595,N_2547);
nand U2733 (N_2733,N_2620,N_2530);
nor U2734 (N_2734,N_2562,N_2593);
nor U2735 (N_2735,N_2615,N_2589);
xnor U2736 (N_2736,N_2598,N_2579);
or U2737 (N_2737,N_2608,N_2614);
or U2738 (N_2738,N_2560,N_2591);
nor U2739 (N_2739,N_2525,N_2501);
or U2740 (N_2740,N_2509,N_2545);
nand U2741 (N_2741,N_2581,N_2525);
nand U2742 (N_2742,N_2510,N_2567);
nor U2743 (N_2743,N_2622,N_2568);
or U2744 (N_2744,N_2602,N_2567);
nand U2745 (N_2745,N_2584,N_2610);
nand U2746 (N_2746,N_2513,N_2598);
and U2747 (N_2747,N_2519,N_2618);
nand U2748 (N_2748,N_2528,N_2505);
nand U2749 (N_2749,N_2598,N_2565);
and U2750 (N_2750,N_2727,N_2681);
or U2751 (N_2751,N_2662,N_2649);
or U2752 (N_2752,N_2725,N_2708);
nor U2753 (N_2753,N_2728,N_2719);
and U2754 (N_2754,N_2690,N_2736);
or U2755 (N_2755,N_2655,N_2671);
nand U2756 (N_2756,N_2700,N_2633);
xnor U2757 (N_2757,N_2718,N_2626);
and U2758 (N_2758,N_2643,N_2711);
nand U2759 (N_2759,N_2737,N_2667);
or U2760 (N_2760,N_2706,N_2721);
and U2761 (N_2761,N_2640,N_2741);
and U2762 (N_2762,N_2664,N_2692);
xnor U2763 (N_2763,N_2694,N_2720);
and U2764 (N_2764,N_2687,N_2650);
or U2765 (N_2765,N_2749,N_2723);
nand U2766 (N_2766,N_2709,N_2638);
nand U2767 (N_2767,N_2689,N_2651);
or U2768 (N_2768,N_2666,N_2740);
and U2769 (N_2769,N_2631,N_2629);
nor U2770 (N_2770,N_2663,N_2634);
nor U2771 (N_2771,N_2665,N_2743);
nand U2772 (N_2772,N_2734,N_2748);
nand U2773 (N_2773,N_2672,N_2714);
xnor U2774 (N_2774,N_2744,N_2716);
or U2775 (N_2775,N_2722,N_2659);
nand U2776 (N_2776,N_2644,N_2642);
nor U2777 (N_2777,N_2701,N_2698);
nor U2778 (N_2778,N_2691,N_2747);
and U2779 (N_2779,N_2679,N_2695);
nand U2780 (N_2780,N_2646,N_2738);
and U2781 (N_2781,N_2712,N_2731);
nor U2782 (N_2782,N_2680,N_2677);
xnor U2783 (N_2783,N_2697,N_2715);
xor U2784 (N_2784,N_2636,N_2746);
nand U2785 (N_2785,N_2630,N_2641);
and U2786 (N_2786,N_2683,N_2688);
nor U2787 (N_2787,N_2703,N_2678);
and U2788 (N_2788,N_2658,N_2656);
xnor U2789 (N_2789,N_2628,N_2745);
or U2790 (N_2790,N_2674,N_2735);
xnor U2791 (N_2791,N_2730,N_2635);
nand U2792 (N_2792,N_2686,N_2668);
xnor U2793 (N_2793,N_2732,N_2627);
nand U2794 (N_2794,N_2705,N_2637);
nor U2795 (N_2795,N_2675,N_2682);
nand U2796 (N_2796,N_2657,N_2661);
xnor U2797 (N_2797,N_2710,N_2713);
xor U2798 (N_2798,N_2625,N_2652);
nand U2799 (N_2799,N_2647,N_2676);
and U2800 (N_2800,N_2704,N_2685);
xor U2801 (N_2801,N_2742,N_2660);
and U2802 (N_2802,N_2645,N_2729);
and U2803 (N_2803,N_2653,N_2648);
xnor U2804 (N_2804,N_2673,N_2726);
nor U2805 (N_2805,N_2670,N_2724);
xor U2806 (N_2806,N_2707,N_2632);
and U2807 (N_2807,N_2669,N_2702);
nor U2808 (N_2808,N_2699,N_2696);
nand U2809 (N_2809,N_2684,N_2639);
xor U2810 (N_2810,N_2717,N_2739);
nor U2811 (N_2811,N_2654,N_2693);
or U2812 (N_2812,N_2733,N_2732);
nand U2813 (N_2813,N_2660,N_2642);
and U2814 (N_2814,N_2675,N_2724);
and U2815 (N_2815,N_2679,N_2632);
nor U2816 (N_2816,N_2655,N_2714);
xnor U2817 (N_2817,N_2660,N_2675);
and U2818 (N_2818,N_2682,N_2657);
nor U2819 (N_2819,N_2725,N_2662);
and U2820 (N_2820,N_2637,N_2718);
xnor U2821 (N_2821,N_2716,N_2635);
xor U2822 (N_2822,N_2743,N_2663);
or U2823 (N_2823,N_2692,N_2738);
nand U2824 (N_2824,N_2635,N_2727);
xnor U2825 (N_2825,N_2698,N_2650);
and U2826 (N_2826,N_2661,N_2636);
and U2827 (N_2827,N_2660,N_2666);
nand U2828 (N_2828,N_2640,N_2658);
and U2829 (N_2829,N_2721,N_2723);
nand U2830 (N_2830,N_2637,N_2738);
nor U2831 (N_2831,N_2714,N_2642);
xnor U2832 (N_2832,N_2632,N_2669);
and U2833 (N_2833,N_2727,N_2634);
or U2834 (N_2834,N_2691,N_2657);
and U2835 (N_2835,N_2678,N_2741);
nand U2836 (N_2836,N_2666,N_2749);
and U2837 (N_2837,N_2708,N_2743);
nor U2838 (N_2838,N_2701,N_2644);
xor U2839 (N_2839,N_2703,N_2719);
nor U2840 (N_2840,N_2709,N_2728);
and U2841 (N_2841,N_2628,N_2636);
xnor U2842 (N_2842,N_2723,N_2729);
xor U2843 (N_2843,N_2640,N_2649);
nor U2844 (N_2844,N_2683,N_2741);
and U2845 (N_2845,N_2705,N_2648);
nor U2846 (N_2846,N_2652,N_2720);
xnor U2847 (N_2847,N_2691,N_2638);
or U2848 (N_2848,N_2653,N_2636);
nand U2849 (N_2849,N_2653,N_2643);
xor U2850 (N_2850,N_2717,N_2709);
nor U2851 (N_2851,N_2698,N_2662);
and U2852 (N_2852,N_2718,N_2660);
nand U2853 (N_2853,N_2625,N_2736);
nor U2854 (N_2854,N_2707,N_2676);
or U2855 (N_2855,N_2649,N_2725);
xnor U2856 (N_2856,N_2686,N_2629);
nor U2857 (N_2857,N_2676,N_2639);
and U2858 (N_2858,N_2726,N_2692);
and U2859 (N_2859,N_2700,N_2749);
nor U2860 (N_2860,N_2660,N_2705);
nor U2861 (N_2861,N_2697,N_2744);
and U2862 (N_2862,N_2685,N_2662);
nor U2863 (N_2863,N_2740,N_2706);
nand U2864 (N_2864,N_2725,N_2683);
and U2865 (N_2865,N_2695,N_2643);
and U2866 (N_2866,N_2741,N_2718);
xor U2867 (N_2867,N_2708,N_2651);
and U2868 (N_2868,N_2654,N_2742);
nand U2869 (N_2869,N_2694,N_2707);
xor U2870 (N_2870,N_2742,N_2712);
nand U2871 (N_2871,N_2699,N_2636);
or U2872 (N_2872,N_2719,N_2688);
nand U2873 (N_2873,N_2651,N_2735);
xor U2874 (N_2874,N_2708,N_2726);
and U2875 (N_2875,N_2810,N_2834);
or U2876 (N_2876,N_2750,N_2829);
and U2877 (N_2877,N_2809,N_2846);
and U2878 (N_2878,N_2822,N_2804);
nand U2879 (N_2879,N_2780,N_2856);
xor U2880 (N_2880,N_2815,N_2869);
nand U2881 (N_2881,N_2801,N_2765);
and U2882 (N_2882,N_2831,N_2862);
or U2883 (N_2883,N_2770,N_2867);
or U2884 (N_2884,N_2850,N_2786);
or U2885 (N_2885,N_2769,N_2845);
and U2886 (N_2886,N_2772,N_2787);
nand U2887 (N_2887,N_2841,N_2835);
nor U2888 (N_2888,N_2774,N_2762);
nand U2889 (N_2889,N_2756,N_2795);
nand U2890 (N_2890,N_2778,N_2861);
xor U2891 (N_2891,N_2783,N_2782);
nor U2892 (N_2892,N_2812,N_2788);
nand U2893 (N_2893,N_2807,N_2757);
and U2894 (N_2894,N_2870,N_2853);
nand U2895 (N_2895,N_2858,N_2817);
nand U2896 (N_2896,N_2784,N_2775);
xnor U2897 (N_2897,N_2854,N_2839);
and U2898 (N_2898,N_2803,N_2816);
xor U2899 (N_2899,N_2806,N_2802);
xnor U2900 (N_2900,N_2796,N_2830);
or U2901 (N_2901,N_2833,N_2821);
and U2902 (N_2902,N_2863,N_2755);
or U2903 (N_2903,N_2826,N_2820);
nor U2904 (N_2904,N_2813,N_2793);
and U2905 (N_2905,N_2790,N_2859);
nor U2906 (N_2906,N_2865,N_2851);
or U2907 (N_2907,N_2842,N_2792);
nand U2908 (N_2908,N_2773,N_2832);
and U2909 (N_2909,N_2799,N_2798);
nor U2910 (N_2910,N_2855,N_2843);
nor U2911 (N_2911,N_2819,N_2873);
xor U2912 (N_2912,N_2860,N_2866);
xor U2913 (N_2913,N_2753,N_2847);
or U2914 (N_2914,N_2825,N_2752);
and U2915 (N_2915,N_2823,N_2771);
nor U2916 (N_2916,N_2781,N_2764);
and U2917 (N_2917,N_2837,N_2768);
nor U2918 (N_2918,N_2838,N_2868);
nand U2919 (N_2919,N_2766,N_2763);
xor U2920 (N_2920,N_2800,N_2751);
and U2921 (N_2921,N_2871,N_2754);
xor U2922 (N_2922,N_2789,N_2791);
nor U2923 (N_2923,N_2797,N_2776);
or U2924 (N_2924,N_2760,N_2779);
xor U2925 (N_2925,N_2761,N_2857);
or U2926 (N_2926,N_2840,N_2828);
nor U2927 (N_2927,N_2852,N_2836);
or U2928 (N_2928,N_2818,N_2785);
and U2929 (N_2929,N_2849,N_2808);
or U2930 (N_2930,N_2824,N_2811);
xnor U2931 (N_2931,N_2759,N_2844);
nand U2932 (N_2932,N_2874,N_2864);
or U2933 (N_2933,N_2827,N_2805);
and U2934 (N_2934,N_2872,N_2777);
nand U2935 (N_2935,N_2848,N_2758);
nand U2936 (N_2936,N_2767,N_2794);
or U2937 (N_2937,N_2814,N_2765);
and U2938 (N_2938,N_2807,N_2831);
nand U2939 (N_2939,N_2813,N_2762);
or U2940 (N_2940,N_2862,N_2849);
or U2941 (N_2941,N_2751,N_2804);
and U2942 (N_2942,N_2761,N_2873);
xor U2943 (N_2943,N_2817,N_2796);
xnor U2944 (N_2944,N_2832,N_2836);
and U2945 (N_2945,N_2828,N_2819);
nor U2946 (N_2946,N_2810,N_2865);
or U2947 (N_2947,N_2758,N_2802);
and U2948 (N_2948,N_2758,N_2786);
xnor U2949 (N_2949,N_2823,N_2838);
and U2950 (N_2950,N_2846,N_2783);
and U2951 (N_2951,N_2791,N_2823);
nor U2952 (N_2952,N_2835,N_2866);
xnor U2953 (N_2953,N_2798,N_2793);
and U2954 (N_2954,N_2825,N_2866);
nand U2955 (N_2955,N_2855,N_2775);
nor U2956 (N_2956,N_2778,N_2797);
nand U2957 (N_2957,N_2755,N_2753);
nand U2958 (N_2958,N_2849,N_2763);
and U2959 (N_2959,N_2762,N_2816);
nand U2960 (N_2960,N_2853,N_2817);
xnor U2961 (N_2961,N_2752,N_2826);
and U2962 (N_2962,N_2764,N_2765);
or U2963 (N_2963,N_2776,N_2848);
nor U2964 (N_2964,N_2774,N_2780);
or U2965 (N_2965,N_2825,N_2793);
or U2966 (N_2966,N_2837,N_2839);
nand U2967 (N_2967,N_2805,N_2775);
or U2968 (N_2968,N_2820,N_2862);
and U2969 (N_2969,N_2867,N_2858);
nor U2970 (N_2970,N_2812,N_2830);
nand U2971 (N_2971,N_2810,N_2781);
xor U2972 (N_2972,N_2841,N_2780);
nand U2973 (N_2973,N_2786,N_2804);
nor U2974 (N_2974,N_2866,N_2777);
and U2975 (N_2975,N_2861,N_2822);
xor U2976 (N_2976,N_2792,N_2860);
and U2977 (N_2977,N_2762,N_2866);
nor U2978 (N_2978,N_2763,N_2788);
nand U2979 (N_2979,N_2820,N_2870);
xnor U2980 (N_2980,N_2767,N_2832);
or U2981 (N_2981,N_2766,N_2780);
or U2982 (N_2982,N_2808,N_2857);
nor U2983 (N_2983,N_2815,N_2871);
nor U2984 (N_2984,N_2852,N_2857);
nand U2985 (N_2985,N_2849,N_2779);
nor U2986 (N_2986,N_2855,N_2796);
or U2987 (N_2987,N_2874,N_2866);
nand U2988 (N_2988,N_2766,N_2871);
or U2989 (N_2989,N_2828,N_2810);
nand U2990 (N_2990,N_2858,N_2800);
xor U2991 (N_2991,N_2799,N_2785);
nor U2992 (N_2992,N_2871,N_2843);
xor U2993 (N_2993,N_2829,N_2855);
and U2994 (N_2994,N_2766,N_2844);
xor U2995 (N_2995,N_2759,N_2839);
and U2996 (N_2996,N_2859,N_2805);
xnor U2997 (N_2997,N_2787,N_2866);
nor U2998 (N_2998,N_2786,N_2795);
nand U2999 (N_2999,N_2815,N_2826);
nand U3000 (N_3000,N_2990,N_2917);
nand U3001 (N_3001,N_2896,N_2890);
nand U3002 (N_3002,N_2983,N_2883);
nor U3003 (N_3003,N_2976,N_2986);
xor U3004 (N_3004,N_2880,N_2909);
xnor U3005 (N_3005,N_2975,N_2964);
nor U3006 (N_3006,N_2980,N_2997);
nor U3007 (N_3007,N_2891,N_2942);
xor U3008 (N_3008,N_2932,N_2879);
nand U3009 (N_3009,N_2974,N_2957);
xnor U3010 (N_3010,N_2882,N_2999);
and U3011 (N_3011,N_2969,N_2938);
or U3012 (N_3012,N_2902,N_2918);
nand U3013 (N_3013,N_2914,N_2978);
nand U3014 (N_3014,N_2885,N_2961);
nor U3015 (N_3015,N_2971,N_2888);
nor U3016 (N_3016,N_2900,N_2970);
nor U3017 (N_3017,N_2993,N_2939);
nor U3018 (N_3018,N_2931,N_2958);
nand U3019 (N_3019,N_2952,N_2965);
nor U3020 (N_3020,N_2928,N_2989);
or U3021 (N_3021,N_2940,N_2948);
nor U3022 (N_3022,N_2887,N_2906);
and U3023 (N_3023,N_2915,N_2925);
or U3024 (N_3024,N_2959,N_2954);
nand U3025 (N_3025,N_2972,N_2953);
nand U3026 (N_3026,N_2889,N_2996);
and U3027 (N_3027,N_2984,N_2876);
nor U3028 (N_3028,N_2988,N_2956);
and U3029 (N_3029,N_2893,N_2911);
xor U3030 (N_3030,N_2935,N_2897);
xor U3031 (N_3031,N_2947,N_2994);
or U3032 (N_3032,N_2944,N_2927);
and U3033 (N_3033,N_2910,N_2987);
nand U3034 (N_3034,N_2923,N_2963);
nor U3035 (N_3035,N_2875,N_2901);
or U3036 (N_3036,N_2941,N_2877);
xor U3037 (N_3037,N_2907,N_2929);
nand U3038 (N_3038,N_2933,N_2898);
xor U3039 (N_3039,N_2979,N_2905);
nand U3040 (N_3040,N_2960,N_2919);
or U3041 (N_3041,N_2945,N_2950);
nor U3042 (N_3042,N_2894,N_2922);
nand U3043 (N_3043,N_2995,N_2921);
xor U3044 (N_3044,N_2943,N_2924);
and U3045 (N_3045,N_2892,N_2930);
or U3046 (N_3046,N_2916,N_2985);
xor U3047 (N_3047,N_2903,N_2908);
nor U3048 (N_3048,N_2991,N_2955);
and U3049 (N_3049,N_2884,N_2951);
nor U3050 (N_3050,N_2936,N_2998);
or U3051 (N_3051,N_2968,N_2977);
nand U3052 (N_3052,N_2881,N_2926);
and U3053 (N_3053,N_2920,N_2912);
nand U3054 (N_3054,N_2899,N_2895);
or U3055 (N_3055,N_2934,N_2966);
nand U3056 (N_3056,N_2913,N_2946);
nand U3057 (N_3057,N_2973,N_2878);
or U3058 (N_3058,N_2962,N_2886);
and U3059 (N_3059,N_2937,N_2949);
or U3060 (N_3060,N_2981,N_2982);
and U3061 (N_3061,N_2904,N_2967);
nand U3062 (N_3062,N_2992,N_2916);
and U3063 (N_3063,N_2990,N_2899);
nor U3064 (N_3064,N_2910,N_2940);
nand U3065 (N_3065,N_2950,N_2877);
nor U3066 (N_3066,N_2917,N_2900);
or U3067 (N_3067,N_2999,N_2994);
nand U3068 (N_3068,N_2939,N_2886);
nand U3069 (N_3069,N_2992,N_2907);
or U3070 (N_3070,N_2967,N_2896);
or U3071 (N_3071,N_2981,N_2930);
nor U3072 (N_3072,N_2999,N_2968);
or U3073 (N_3073,N_2937,N_2969);
xor U3074 (N_3074,N_2985,N_2993);
and U3075 (N_3075,N_2999,N_2923);
xnor U3076 (N_3076,N_2933,N_2920);
xor U3077 (N_3077,N_2899,N_2894);
or U3078 (N_3078,N_2930,N_2989);
nand U3079 (N_3079,N_2909,N_2888);
nor U3080 (N_3080,N_2995,N_2883);
nor U3081 (N_3081,N_2984,N_2978);
and U3082 (N_3082,N_2995,N_2955);
nor U3083 (N_3083,N_2997,N_2883);
nor U3084 (N_3084,N_2984,N_2896);
nand U3085 (N_3085,N_2875,N_2932);
and U3086 (N_3086,N_2909,N_2946);
nand U3087 (N_3087,N_2951,N_2915);
nor U3088 (N_3088,N_2999,N_2990);
nand U3089 (N_3089,N_2985,N_2960);
nor U3090 (N_3090,N_2939,N_2957);
or U3091 (N_3091,N_2990,N_2989);
nor U3092 (N_3092,N_2937,N_2885);
nand U3093 (N_3093,N_2888,N_2992);
and U3094 (N_3094,N_2993,N_2887);
or U3095 (N_3095,N_2942,N_2879);
or U3096 (N_3096,N_2902,N_2909);
or U3097 (N_3097,N_2958,N_2875);
and U3098 (N_3098,N_2990,N_2883);
nand U3099 (N_3099,N_2893,N_2991);
and U3100 (N_3100,N_2948,N_2972);
xnor U3101 (N_3101,N_2940,N_2924);
or U3102 (N_3102,N_2914,N_2910);
and U3103 (N_3103,N_2949,N_2910);
nor U3104 (N_3104,N_2945,N_2930);
nand U3105 (N_3105,N_2900,N_2908);
nand U3106 (N_3106,N_2883,N_2968);
or U3107 (N_3107,N_2891,N_2985);
xor U3108 (N_3108,N_2963,N_2964);
xnor U3109 (N_3109,N_2950,N_2892);
or U3110 (N_3110,N_2995,N_2944);
nor U3111 (N_3111,N_2929,N_2999);
or U3112 (N_3112,N_2923,N_2925);
nor U3113 (N_3113,N_2955,N_2917);
and U3114 (N_3114,N_2984,N_2927);
nor U3115 (N_3115,N_2986,N_2894);
and U3116 (N_3116,N_2929,N_2982);
xor U3117 (N_3117,N_2939,N_2928);
xor U3118 (N_3118,N_2902,N_2964);
nand U3119 (N_3119,N_2883,N_2944);
and U3120 (N_3120,N_2909,N_2910);
or U3121 (N_3121,N_2950,N_2991);
and U3122 (N_3122,N_2899,N_2997);
nor U3123 (N_3123,N_2878,N_2949);
and U3124 (N_3124,N_2914,N_2952);
or U3125 (N_3125,N_3122,N_3019);
xor U3126 (N_3126,N_3023,N_3043);
nor U3127 (N_3127,N_3024,N_3124);
nor U3128 (N_3128,N_3080,N_3018);
and U3129 (N_3129,N_3062,N_3020);
nor U3130 (N_3130,N_3025,N_3034);
nor U3131 (N_3131,N_3075,N_3057);
nand U3132 (N_3132,N_3108,N_3009);
xor U3133 (N_3133,N_3071,N_3100);
xor U3134 (N_3134,N_3051,N_3015);
nor U3135 (N_3135,N_3065,N_3005);
nand U3136 (N_3136,N_3028,N_3040);
or U3137 (N_3137,N_3004,N_3095);
and U3138 (N_3138,N_3089,N_3116);
nand U3139 (N_3139,N_3086,N_3117);
xor U3140 (N_3140,N_3031,N_3111);
nand U3141 (N_3141,N_3002,N_3037);
and U3142 (N_3142,N_3060,N_3112);
nor U3143 (N_3143,N_3114,N_3022);
and U3144 (N_3144,N_3121,N_3068);
nor U3145 (N_3145,N_3093,N_3054);
or U3146 (N_3146,N_3044,N_3090);
nand U3147 (N_3147,N_3021,N_3096);
nand U3148 (N_3148,N_3066,N_3047);
or U3149 (N_3149,N_3049,N_3016);
nand U3150 (N_3150,N_3106,N_3052);
and U3151 (N_3151,N_3045,N_3099);
nand U3152 (N_3152,N_3115,N_3102);
xnor U3153 (N_3153,N_3030,N_3072);
or U3154 (N_3154,N_3070,N_3073);
nor U3155 (N_3155,N_3081,N_3110);
xor U3156 (N_3156,N_3076,N_3123);
or U3157 (N_3157,N_3027,N_3064);
and U3158 (N_3158,N_3101,N_3056);
and U3159 (N_3159,N_3105,N_3039);
or U3160 (N_3160,N_3085,N_3006);
xnor U3161 (N_3161,N_3011,N_3084);
nand U3162 (N_3162,N_3038,N_3067);
and U3163 (N_3163,N_3074,N_3107);
nand U3164 (N_3164,N_3098,N_3035);
and U3165 (N_3165,N_3104,N_3091);
xor U3166 (N_3166,N_3048,N_3082);
and U3167 (N_3167,N_3046,N_3120);
or U3168 (N_3168,N_3077,N_3000);
and U3169 (N_3169,N_3069,N_3103);
nand U3170 (N_3170,N_3059,N_3017);
nand U3171 (N_3171,N_3001,N_3061);
and U3172 (N_3172,N_3029,N_3113);
nand U3173 (N_3173,N_3079,N_3092);
xor U3174 (N_3174,N_3050,N_3078);
and U3175 (N_3175,N_3109,N_3026);
xor U3176 (N_3176,N_3058,N_3042);
xor U3177 (N_3177,N_3087,N_3094);
nor U3178 (N_3178,N_3119,N_3088);
or U3179 (N_3179,N_3013,N_3118);
or U3180 (N_3180,N_3014,N_3033);
or U3181 (N_3181,N_3008,N_3053);
or U3182 (N_3182,N_3063,N_3036);
and U3183 (N_3183,N_3003,N_3010);
or U3184 (N_3184,N_3012,N_3032);
xnor U3185 (N_3185,N_3007,N_3083);
nand U3186 (N_3186,N_3055,N_3097);
nor U3187 (N_3187,N_3041,N_3056);
nand U3188 (N_3188,N_3021,N_3080);
xnor U3189 (N_3189,N_3032,N_3096);
nor U3190 (N_3190,N_3002,N_3066);
xnor U3191 (N_3191,N_3026,N_3008);
nor U3192 (N_3192,N_3067,N_3081);
and U3193 (N_3193,N_3094,N_3092);
xor U3194 (N_3194,N_3099,N_3023);
nand U3195 (N_3195,N_3040,N_3026);
and U3196 (N_3196,N_3110,N_3055);
xnor U3197 (N_3197,N_3055,N_3060);
nand U3198 (N_3198,N_3013,N_3091);
and U3199 (N_3199,N_3100,N_3069);
or U3200 (N_3200,N_3032,N_3075);
xor U3201 (N_3201,N_3112,N_3011);
or U3202 (N_3202,N_3071,N_3056);
and U3203 (N_3203,N_3042,N_3060);
or U3204 (N_3204,N_3023,N_3039);
or U3205 (N_3205,N_3073,N_3050);
or U3206 (N_3206,N_3045,N_3010);
nor U3207 (N_3207,N_3112,N_3107);
and U3208 (N_3208,N_3097,N_3009);
nor U3209 (N_3209,N_3074,N_3106);
nand U3210 (N_3210,N_3089,N_3018);
nand U3211 (N_3211,N_3013,N_3060);
or U3212 (N_3212,N_3107,N_3100);
and U3213 (N_3213,N_3031,N_3010);
xor U3214 (N_3214,N_3051,N_3008);
nor U3215 (N_3215,N_3018,N_3034);
nand U3216 (N_3216,N_3101,N_3035);
or U3217 (N_3217,N_3066,N_3007);
nor U3218 (N_3218,N_3029,N_3100);
or U3219 (N_3219,N_3053,N_3013);
nand U3220 (N_3220,N_3084,N_3093);
or U3221 (N_3221,N_3069,N_3093);
nor U3222 (N_3222,N_3038,N_3090);
xor U3223 (N_3223,N_3110,N_3122);
or U3224 (N_3224,N_3047,N_3058);
or U3225 (N_3225,N_3041,N_3115);
or U3226 (N_3226,N_3076,N_3008);
and U3227 (N_3227,N_3001,N_3007);
nor U3228 (N_3228,N_3096,N_3030);
or U3229 (N_3229,N_3114,N_3025);
nand U3230 (N_3230,N_3001,N_3096);
nand U3231 (N_3231,N_3011,N_3076);
or U3232 (N_3232,N_3119,N_3019);
and U3233 (N_3233,N_3032,N_3016);
nand U3234 (N_3234,N_3029,N_3043);
xor U3235 (N_3235,N_3085,N_3092);
xor U3236 (N_3236,N_3094,N_3001);
nand U3237 (N_3237,N_3122,N_3052);
nand U3238 (N_3238,N_3113,N_3080);
nand U3239 (N_3239,N_3027,N_3007);
or U3240 (N_3240,N_3026,N_3058);
and U3241 (N_3241,N_3064,N_3079);
nand U3242 (N_3242,N_3099,N_3074);
xor U3243 (N_3243,N_3121,N_3053);
and U3244 (N_3244,N_3082,N_3072);
nand U3245 (N_3245,N_3011,N_3069);
nand U3246 (N_3246,N_3016,N_3024);
and U3247 (N_3247,N_3101,N_3055);
nand U3248 (N_3248,N_3031,N_3062);
nor U3249 (N_3249,N_3082,N_3094);
or U3250 (N_3250,N_3220,N_3216);
and U3251 (N_3251,N_3130,N_3162);
nand U3252 (N_3252,N_3153,N_3214);
and U3253 (N_3253,N_3157,N_3163);
and U3254 (N_3254,N_3226,N_3143);
xor U3255 (N_3255,N_3239,N_3243);
nand U3256 (N_3256,N_3234,N_3139);
and U3257 (N_3257,N_3183,N_3167);
nor U3258 (N_3258,N_3230,N_3225);
and U3259 (N_3259,N_3184,N_3246);
nor U3260 (N_3260,N_3231,N_3198);
nand U3261 (N_3261,N_3148,N_3127);
nand U3262 (N_3262,N_3140,N_3233);
xnor U3263 (N_3263,N_3138,N_3196);
xnor U3264 (N_3264,N_3161,N_3219);
or U3265 (N_3265,N_3141,N_3170);
or U3266 (N_3266,N_3188,N_3155);
xor U3267 (N_3267,N_3145,N_3205);
nor U3268 (N_3268,N_3142,N_3175);
and U3269 (N_3269,N_3242,N_3192);
xor U3270 (N_3270,N_3241,N_3174);
nor U3271 (N_3271,N_3187,N_3248);
nand U3272 (N_3272,N_3168,N_3222);
or U3273 (N_3273,N_3211,N_3228);
nor U3274 (N_3274,N_3247,N_3149);
nor U3275 (N_3275,N_3134,N_3165);
nor U3276 (N_3276,N_3209,N_3191);
nor U3277 (N_3277,N_3150,N_3223);
or U3278 (N_3278,N_3218,N_3186);
nor U3279 (N_3279,N_3144,N_3128);
or U3280 (N_3280,N_3129,N_3229);
nor U3281 (N_3281,N_3125,N_3210);
nor U3282 (N_3282,N_3212,N_3172);
and U3283 (N_3283,N_3202,N_3194);
or U3284 (N_3284,N_3156,N_3203);
nor U3285 (N_3285,N_3185,N_3224);
nand U3286 (N_3286,N_3206,N_3200);
or U3287 (N_3287,N_3126,N_3208);
xor U3288 (N_3288,N_3189,N_3158);
nor U3289 (N_3289,N_3180,N_3232);
xnor U3290 (N_3290,N_3204,N_3181);
xnor U3291 (N_3291,N_3227,N_3132);
or U3292 (N_3292,N_3213,N_3137);
or U3293 (N_3293,N_3146,N_3217);
nor U3294 (N_3294,N_3131,N_3182);
nand U3295 (N_3295,N_3136,N_3169);
xor U3296 (N_3296,N_3152,N_3135);
nand U3297 (N_3297,N_3173,N_3179);
or U3298 (N_3298,N_3215,N_3160);
xor U3299 (N_3299,N_3164,N_3171);
or U3300 (N_3300,N_3193,N_3190);
nand U3301 (N_3301,N_3238,N_3147);
or U3302 (N_3302,N_3195,N_3221);
xnor U3303 (N_3303,N_3236,N_3245);
or U3304 (N_3304,N_3237,N_3151);
xnor U3305 (N_3305,N_3240,N_3199);
or U3306 (N_3306,N_3176,N_3159);
xnor U3307 (N_3307,N_3249,N_3178);
and U3308 (N_3308,N_3197,N_3201);
nand U3309 (N_3309,N_3235,N_3177);
or U3310 (N_3310,N_3154,N_3207);
nor U3311 (N_3311,N_3166,N_3244);
nor U3312 (N_3312,N_3133,N_3130);
xor U3313 (N_3313,N_3226,N_3173);
or U3314 (N_3314,N_3179,N_3239);
nor U3315 (N_3315,N_3177,N_3244);
or U3316 (N_3316,N_3230,N_3166);
and U3317 (N_3317,N_3189,N_3129);
nand U3318 (N_3318,N_3136,N_3170);
nor U3319 (N_3319,N_3202,N_3211);
nor U3320 (N_3320,N_3140,N_3142);
nor U3321 (N_3321,N_3188,N_3136);
or U3322 (N_3322,N_3198,N_3189);
nand U3323 (N_3323,N_3144,N_3193);
nand U3324 (N_3324,N_3144,N_3125);
or U3325 (N_3325,N_3139,N_3236);
and U3326 (N_3326,N_3154,N_3221);
nor U3327 (N_3327,N_3143,N_3231);
nor U3328 (N_3328,N_3163,N_3165);
and U3329 (N_3329,N_3126,N_3240);
and U3330 (N_3330,N_3177,N_3154);
and U3331 (N_3331,N_3224,N_3210);
xnor U3332 (N_3332,N_3240,N_3228);
and U3333 (N_3333,N_3248,N_3148);
and U3334 (N_3334,N_3159,N_3160);
xor U3335 (N_3335,N_3175,N_3183);
nand U3336 (N_3336,N_3193,N_3236);
nand U3337 (N_3337,N_3162,N_3218);
nor U3338 (N_3338,N_3149,N_3248);
or U3339 (N_3339,N_3179,N_3185);
nand U3340 (N_3340,N_3177,N_3144);
nand U3341 (N_3341,N_3220,N_3148);
xnor U3342 (N_3342,N_3212,N_3183);
or U3343 (N_3343,N_3214,N_3234);
nand U3344 (N_3344,N_3146,N_3132);
or U3345 (N_3345,N_3133,N_3153);
nand U3346 (N_3346,N_3142,N_3176);
nand U3347 (N_3347,N_3168,N_3214);
nand U3348 (N_3348,N_3161,N_3230);
nand U3349 (N_3349,N_3228,N_3163);
or U3350 (N_3350,N_3198,N_3135);
or U3351 (N_3351,N_3145,N_3187);
nor U3352 (N_3352,N_3202,N_3234);
and U3353 (N_3353,N_3158,N_3149);
or U3354 (N_3354,N_3131,N_3167);
xnor U3355 (N_3355,N_3133,N_3211);
nor U3356 (N_3356,N_3172,N_3216);
xor U3357 (N_3357,N_3205,N_3195);
nor U3358 (N_3358,N_3225,N_3151);
or U3359 (N_3359,N_3230,N_3146);
or U3360 (N_3360,N_3164,N_3219);
or U3361 (N_3361,N_3147,N_3216);
and U3362 (N_3362,N_3225,N_3188);
xnor U3363 (N_3363,N_3231,N_3200);
or U3364 (N_3364,N_3173,N_3133);
xor U3365 (N_3365,N_3142,N_3249);
and U3366 (N_3366,N_3223,N_3160);
and U3367 (N_3367,N_3136,N_3171);
nor U3368 (N_3368,N_3130,N_3247);
nor U3369 (N_3369,N_3232,N_3135);
xor U3370 (N_3370,N_3148,N_3181);
nand U3371 (N_3371,N_3239,N_3229);
nand U3372 (N_3372,N_3236,N_3234);
and U3373 (N_3373,N_3179,N_3139);
xor U3374 (N_3374,N_3131,N_3202);
or U3375 (N_3375,N_3339,N_3290);
nor U3376 (N_3376,N_3278,N_3253);
nor U3377 (N_3377,N_3335,N_3294);
nor U3378 (N_3378,N_3336,N_3281);
nand U3379 (N_3379,N_3362,N_3292);
and U3380 (N_3380,N_3293,N_3325);
or U3381 (N_3381,N_3318,N_3264);
or U3382 (N_3382,N_3354,N_3273);
nor U3383 (N_3383,N_3313,N_3357);
xor U3384 (N_3384,N_3321,N_3355);
and U3385 (N_3385,N_3307,N_3266);
and U3386 (N_3386,N_3340,N_3261);
nand U3387 (N_3387,N_3279,N_3306);
or U3388 (N_3388,N_3271,N_3364);
nor U3389 (N_3389,N_3343,N_3342);
and U3390 (N_3390,N_3268,N_3324);
or U3391 (N_3391,N_3320,N_3298);
nand U3392 (N_3392,N_3297,N_3367);
nor U3393 (N_3393,N_3286,N_3374);
and U3394 (N_3394,N_3347,N_3295);
xnor U3395 (N_3395,N_3267,N_3304);
nor U3396 (N_3396,N_3371,N_3262);
nand U3397 (N_3397,N_3317,N_3350);
and U3398 (N_3398,N_3299,N_3257);
nand U3399 (N_3399,N_3260,N_3258);
nand U3400 (N_3400,N_3356,N_3338);
nand U3401 (N_3401,N_3323,N_3361);
xnor U3402 (N_3402,N_3359,N_3309);
xor U3403 (N_3403,N_3291,N_3308);
or U3404 (N_3404,N_3250,N_3300);
nor U3405 (N_3405,N_3327,N_3372);
nand U3406 (N_3406,N_3259,N_3277);
and U3407 (N_3407,N_3322,N_3288);
or U3408 (N_3408,N_3256,N_3283);
nand U3409 (N_3409,N_3331,N_3346);
nand U3410 (N_3410,N_3251,N_3312);
and U3411 (N_3411,N_3363,N_3255);
or U3412 (N_3412,N_3353,N_3269);
nand U3413 (N_3413,N_3272,N_3314);
nand U3414 (N_3414,N_3285,N_3280);
and U3415 (N_3415,N_3305,N_3348);
nor U3416 (N_3416,N_3275,N_3329);
nand U3417 (N_3417,N_3341,N_3284);
and U3418 (N_3418,N_3349,N_3330);
or U3419 (N_3419,N_3303,N_3287);
nor U3420 (N_3420,N_3337,N_3365);
nand U3421 (N_3421,N_3369,N_3368);
or U3422 (N_3422,N_3310,N_3352);
or U3423 (N_3423,N_3296,N_3351);
nor U3424 (N_3424,N_3282,N_3358);
and U3425 (N_3425,N_3315,N_3360);
or U3426 (N_3426,N_3319,N_3265);
nor U3427 (N_3427,N_3326,N_3302);
nor U3428 (N_3428,N_3289,N_3276);
xor U3429 (N_3429,N_3333,N_3366);
or U3430 (N_3430,N_3301,N_3332);
nand U3431 (N_3431,N_3270,N_3334);
or U3432 (N_3432,N_3252,N_3311);
and U3433 (N_3433,N_3344,N_3370);
xor U3434 (N_3434,N_3316,N_3345);
and U3435 (N_3435,N_3263,N_3328);
xor U3436 (N_3436,N_3274,N_3373);
or U3437 (N_3437,N_3254,N_3321);
and U3438 (N_3438,N_3263,N_3299);
nor U3439 (N_3439,N_3262,N_3324);
and U3440 (N_3440,N_3373,N_3310);
and U3441 (N_3441,N_3322,N_3251);
xor U3442 (N_3442,N_3366,N_3295);
and U3443 (N_3443,N_3347,N_3352);
nor U3444 (N_3444,N_3318,N_3372);
and U3445 (N_3445,N_3320,N_3274);
or U3446 (N_3446,N_3310,N_3313);
nor U3447 (N_3447,N_3258,N_3282);
xnor U3448 (N_3448,N_3271,N_3326);
and U3449 (N_3449,N_3298,N_3252);
nor U3450 (N_3450,N_3361,N_3295);
and U3451 (N_3451,N_3348,N_3337);
xnor U3452 (N_3452,N_3333,N_3257);
nand U3453 (N_3453,N_3251,N_3357);
or U3454 (N_3454,N_3311,N_3261);
or U3455 (N_3455,N_3373,N_3354);
xor U3456 (N_3456,N_3293,N_3297);
and U3457 (N_3457,N_3308,N_3314);
nand U3458 (N_3458,N_3291,N_3338);
or U3459 (N_3459,N_3288,N_3264);
and U3460 (N_3460,N_3299,N_3266);
or U3461 (N_3461,N_3363,N_3314);
xnor U3462 (N_3462,N_3331,N_3358);
or U3463 (N_3463,N_3319,N_3262);
nor U3464 (N_3464,N_3347,N_3278);
or U3465 (N_3465,N_3352,N_3290);
xnor U3466 (N_3466,N_3325,N_3261);
nor U3467 (N_3467,N_3334,N_3364);
or U3468 (N_3468,N_3303,N_3323);
or U3469 (N_3469,N_3365,N_3306);
xnor U3470 (N_3470,N_3335,N_3313);
or U3471 (N_3471,N_3267,N_3277);
nor U3472 (N_3472,N_3271,N_3358);
and U3473 (N_3473,N_3298,N_3294);
xor U3474 (N_3474,N_3335,N_3355);
or U3475 (N_3475,N_3289,N_3304);
or U3476 (N_3476,N_3339,N_3285);
xor U3477 (N_3477,N_3346,N_3368);
xnor U3478 (N_3478,N_3324,N_3306);
xnor U3479 (N_3479,N_3340,N_3329);
or U3480 (N_3480,N_3298,N_3323);
nand U3481 (N_3481,N_3319,N_3359);
nor U3482 (N_3482,N_3261,N_3289);
xor U3483 (N_3483,N_3288,N_3332);
nor U3484 (N_3484,N_3278,N_3263);
xnor U3485 (N_3485,N_3314,N_3351);
nand U3486 (N_3486,N_3349,N_3334);
xor U3487 (N_3487,N_3341,N_3266);
nand U3488 (N_3488,N_3341,N_3310);
nor U3489 (N_3489,N_3272,N_3334);
nand U3490 (N_3490,N_3335,N_3339);
and U3491 (N_3491,N_3270,N_3272);
nor U3492 (N_3492,N_3280,N_3345);
and U3493 (N_3493,N_3279,N_3320);
and U3494 (N_3494,N_3287,N_3282);
nor U3495 (N_3495,N_3282,N_3265);
and U3496 (N_3496,N_3275,N_3339);
xnor U3497 (N_3497,N_3297,N_3281);
nand U3498 (N_3498,N_3259,N_3296);
or U3499 (N_3499,N_3366,N_3305);
xnor U3500 (N_3500,N_3419,N_3436);
and U3501 (N_3501,N_3412,N_3494);
xor U3502 (N_3502,N_3440,N_3395);
and U3503 (N_3503,N_3423,N_3463);
nor U3504 (N_3504,N_3434,N_3397);
and U3505 (N_3505,N_3450,N_3420);
and U3506 (N_3506,N_3379,N_3484);
and U3507 (N_3507,N_3393,N_3443);
or U3508 (N_3508,N_3491,N_3413);
nor U3509 (N_3509,N_3407,N_3394);
or U3510 (N_3510,N_3460,N_3468);
or U3511 (N_3511,N_3469,N_3400);
nor U3512 (N_3512,N_3432,N_3483);
and U3513 (N_3513,N_3453,N_3449);
xor U3514 (N_3514,N_3384,N_3462);
and U3515 (N_3515,N_3442,N_3386);
and U3516 (N_3516,N_3459,N_3495);
nor U3517 (N_3517,N_3376,N_3416);
and U3518 (N_3518,N_3418,N_3425);
xor U3519 (N_3519,N_3485,N_3441);
and U3520 (N_3520,N_3480,N_3385);
or U3521 (N_3521,N_3435,N_3389);
and U3522 (N_3522,N_3392,N_3490);
nand U3523 (N_3523,N_3437,N_3448);
nand U3524 (N_3524,N_3438,N_3405);
nor U3525 (N_3525,N_3429,N_3482);
nor U3526 (N_3526,N_3487,N_3422);
nand U3527 (N_3527,N_3375,N_3382);
nand U3528 (N_3528,N_3421,N_3415);
or U3529 (N_3529,N_3488,N_3424);
and U3530 (N_3530,N_3479,N_3388);
xor U3531 (N_3531,N_3497,N_3433);
or U3532 (N_3532,N_3454,N_3473);
and U3533 (N_3533,N_3451,N_3409);
xnor U3534 (N_3534,N_3474,N_3410);
xnor U3535 (N_3535,N_3390,N_3466);
nor U3536 (N_3536,N_3456,N_3430);
xnor U3537 (N_3537,N_3439,N_3414);
or U3538 (N_3538,N_3486,N_3381);
and U3539 (N_3539,N_3403,N_3444);
nor U3540 (N_3540,N_3402,N_3481);
nor U3541 (N_3541,N_3489,N_3399);
and U3542 (N_3542,N_3408,N_3492);
or U3543 (N_3543,N_3417,N_3470);
nor U3544 (N_3544,N_3493,N_3461);
xor U3545 (N_3545,N_3471,N_3472);
xnor U3546 (N_3546,N_3447,N_3475);
nor U3547 (N_3547,N_3404,N_3401);
or U3548 (N_3548,N_3391,N_3455);
and U3549 (N_3549,N_3478,N_3396);
xor U3550 (N_3550,N_3427,N_3465);
xnor U3551 (N_3551,N_3498,N_3411);
nor U3552 (N_3552,N_3426,N_3445);
xnor U3553 (N_3553,N_3446,N_3452);
nand U3554 (N_3554,N_3377,N_3457);
nand U3555 (N_3555,N_3464,N_3428);
and U3556 (N_3556,N_3406,N_3499);
xnor U3557 (N_3557,N_3398,N_3387);
nor U3558 (N_3558,N_3378,N_3380);
and U3559 (N_3559,N_3383,N_3431);
nand U3560 (N_3560,N_3458,N_3496);
nor U3561 (N_3561,N_3467,N_3476);
nor U3562 (N_3562,N_3477,N_3388);
nor U3563 (N_3563,N_3466,N_3484);
and U3564 (N_3564,N_3418,N_3491);
xor U3565 (N_3565,N_3496,N_3459);
or U3566 (N_3566,N_3487,N_3389);
xnor U3567 (N_3567,N_3424,N_3400);
nor U3568 (N_3568,N_3396,N_3470);
nor U3569 (N_3569,N_3426,N_3443);
and U3570 (N_3570,N_3385,N_3437);
nor U3571 (N_3571,N_3424,N_3490);
and U3572 (N_3572,N_3395,N_3497);
nand U3573 (N_3573,N_3492,N_3444);
nor U3574 (N_3574,N_3480,N_3486);
nand U3575 (N_3575,N_3445,N_3480);
nand U3576 (N_3576,N_3435,N_3499);
nand U3577 (N_3577,N_3459,N_3476);
and U3578 (N_3578,N_3454,N_3413);
xor U3579 (N_3579,N_3480,N_3377);
nor U3580 (N_3580,N_3423,N_3469);
xor U3581 (N_3581,N_3386,N_3414);
and U3582 (N_3582,N_3462,N_3392);
and U3583 (N_3583,N_3472,N_3392);
xnor U3584 (N_3584,N_3376,N_3398);
nand U3585 (N_3585,N_3401,N_3409);
and U3586 (N_3586,N_3395,N_3472);
and U3587 (N_3587,N_3388,N_3423);
nor U3588 (N_3588,N_3399,N_3498);
or U3589 (N_3589,N_3406,N_3392);
nor U3590 (N_3590,N_3403,N_3391);
xnor U3591 (N_3591,N_3450,N_3432);
or U3592 (N_3592,N_3412,N_3459);
nor U3593 (N_3593,N_3385,N_3486);
nor U3594 (N_3594,N_3408,N_3487);
nand U3595 (N_3595,N_3460,N_3488);
and U3596 (N_3596,N_3479,N_3419);
xor U3597 (N_3597,N_3425,N_3479);
and U3598 (N_3598,N_3389,N_3419);
xnor U3599 (N_3599,N_3388,N_3411);
or U3600 (N_3600,N_3396,N_3430);
and U3601 (N_3601,N_3452,N_3432);
nor U3602 (N_3602,N_3444,N_3388);
or U3603 (N_3603,N_3447,N_3433);
or U3604 (N_3604,N_3480,N_3490);
and U3605 (N_3605,N_3399,N_3434);
or U3606 (N_3606,N_3419,N_3397);
and U3607 (N_3607,N_3469,N_3382);
or U3608 (N_3608,N_3451,N_3481);
xor U3609 (N_3609,N_3498,N_3409);
nor U3610 (N_3610,N_3438,N_3463);
or U3611 (N_3611,N_3447,N_3439);
nor U3612 (N_3612,N_3458,N_3454);
xnor U3613 (N_3613,N_3379,N_3499);
nor U3614 (N_3614,N_3410,N_3459);
nor U3615 (N_3615,N_3496,N_3394);
and U3616 (N_3616,N_3390,N_3470);
or U3617 (N_3617,N_3498,N_3497);
xnor U3618 (N_3618,N_3447,N_3480);
xor U3619 (N_3619,N_3429,N_3391);
and U3620 (N_3620,N_3390,N_3469);
nor U3621 (N_3621,N_3449,N_3380);
and U3622 (N_3622,N_3401,N_3456);
and U3623 (N_3623,N_3419,N_3483);
xor U3624 (N_3624,N_3454,N_3426);
or U3625 (N_3625,N_3510,N_3553);
or U3626 (N_3626,N_3572,N_3568);
nand U3627 (N_3627,N_3575,N_3540);
and U3628 (N_3628,N_3607,N_3574);
nand U3629 (N_3629,N_3614,N_3578);
or U3630 (N_3630,N_3587,N_3550);
xnor U3631 (N_3631,N_3582,N_3502);
nand U3632 (N_3632,N_3508,N_3544);
and U3633 (N_3633,N_3564,N_3551);
or U3634 (N_3634,N_3605,N_3532);
nor U3635 (N_3635,N_3504,N_3501);
and U3636 (N_3636,N_3511,N_3590);
and U3637 (N_3637,N_3620,N_3597);
or U3638 (N_3638,N_3616,N_3610);
nand U3639 (N_3639,N_3554,N_3580);
nand U3640 (N_3640,N_3577,N_3500);
nand U3641 (N_3641,N_3612,N_3596);
or U3642 (N_3642,N_3523,N_3604);
and U3643 (N_3643,N_3589,N_3588);
nand U3644 (N_3644,N_3558,N_3545);
xnor U3645 (N_3645,N_3624,N_3561);
or U3646 (N_3646,N_3525,N_3565);
xor U3647 (N_3647,N_3585,N_3535);
nand U3648 (N_3648,N_3514,N_3517);
nand U3649 (N_3649,N_3509,N_3524);
nor U3650 (N_3650,N_3560,N_3593);
and U3651 (N_3651,N_3506,N_3623);
nand U3652 (N_3652,N_3606,N_3542);
nand U3653 (N_3653,N_3601,N_3529);
or U3654 (N_3654,N_3536,N_3521);
or U3655 (N_3655,N_3557,N_3555);
or U3656 (N_3656,N_3622,N_3533);
and U3657 (N_3657,N_3570,N_3567);
nor U3658 (N_3658,N_3552,N_3537);
and U3659 (N_3659,N_3528,N_3512);
or U3660 (N_3660,N_3617,N_3546);
xnor U3661 (N_3661,N_3571,N_3541);
nor U3662 (N_3662,N_3548,N_3563);
nor U3663 (N_3663,N_3595,N_3549);
or U3664 (N_3664,N_3566,N_3527);
or U3665 (N_3665,N_3609,N_3538);
nor U3666 (N_3666,N_3522,N_3569);
xor U3667 (N_3667,N_3507,N_3615);
and U3668 (N_3668,N_3503,N_3576);
or U3669 (N_3669,N_3530,N_3599);
nand U3670 (N_3670,N_3583,N_3586);
and U3671 (N_3671,N_3608,N_3518);
and U3672 (N_3672,N_3584,N_3543);
xnor U3673 (N_3673,N_3516,N_3531);
xnor U3674 (N_3674,N_3621,N_3526);
and U3675 (N_3675,N_3581,N_3579);
or U3676 (N_3676,N_3573,N_3603);
nand U3677 (N_3677,N_3505,N_3592);
and U3678 (N_3678,N_3618,N_3547);
or U3679 (N_3679,N_3520,N_3539);
nor U3680 (N_3680,N_3534,N_3598);
nor U3681 (N_3681,N_3515,N_3513);
xor U3682 (N_3682,N_3619,N_3600);
xnor U3683 (N_3683,N_3556,N_3613);
and U3684 (N_3684,N_3591,N_3611);
or U3685 (N_3685,N_3519,N_3602);
nand U3686 (N_3686,N_3559,N_3562);
nand U3687 (N_3687,N_3594,N_3584);
nor U3688 (N_3688,N_3516,N_3518);
or U3689 (N_3689,N_3513,N_3559);
and U3690 (N_3690,N_3583,N_3520);
nor U3691 (N_3691,N_3505,N_3533);
or U3692 (N_3692,N_3590,N_3604);
or U3693 (N_3693,N_3509,N_3592);
nand U3694 (N_3694,N_3566,N_3501);
xnor U3695 (N_3695,N_3592,N_3569);
nand U3696 (N_3696,N_3576,N_3559);
or U3697 (N_3697,N_3505,N_3607);
xnor U3698 (N_3698,N_3604,N_3578);
xor U3699 (N_3699,N_3525,N_3544);
nand U3700 (N_3700,N_3537,N_3517);
and U3701 (N_3701,N_3582,N_3593);
xor U3702 (N_3702,N_3528,N_3566);
nand U3703 (N_3703,N_3598,N_3604);
nand U3704 (N_3704,N_3524,N_3608);
nand U3705 (N_3705,N_3616,N_3617);
or U3706 (N_3706,N_3510,N_3587);
or U3707 (N_3707,N_3613,N_3547);
nand U3708 (N_3708,N_3515,N_3530);
nand U3709 (N_3709,N_3518,N_3579);
and U3710 (N_3710,N_3537,N_3576);
nor U3711 (N_3711,N_3554,N_3512);
nor U3712 (N_3712,N_3506,N_3584);
or U3713 (N_3713,N_3531,N_3556);
and U3714 (N_3714,N_3544,N_3610);
xor U3715 (N_3715,N_3546,N_3519);
or U3716 (N_3716,N_3573,N_3539);
xnor U3717 (N_3717,N_3507,N_3538);
and U3718 (N_3718,N_3517,N_3584);
nor U3719 (N_3719,N_3566,N_3561);
nand U3720 (N_3720,N_3556,N_3535);
and U3721 (N_3721,N_3594,N_3568);
nor U3722 (N_3722,N_3597,N_3507);
nand U3723 (N_3723,N_3567,N_3521);
nand U3724 (N_3724,N_3566,N_3535);
nand U3725 (N_3725,N_3594,N_3517);
xor U3726 (N_3726,N_3514,N_3572);
nor U3727 (N_3727,N_3619,N_3520);
nor U3728 (N_3728,N_3611,N_3517);
or U3729 (N_3729,N_3573,N_3612);
or U3730 (N_3730,N_3547,N_3596);
or U3731 (N_3731,N_3594,N_3527);
or U3732 (N_3732,N_3564,N_3542);
xnor U3733 (N_3733,N_3607,N_3599);
xnor U3734 (N_3734,N_3607,N_3502);
and U3735 (N_3735,N_3595,N_3539);
nor U3736 (N_3736,N_3529,N_3554);
xnor U3737 (N_3737,N_3529,N_3571);
and U3738 (N_3738,N_3544,N_3603);
and U3739 (N_3739,N_3548,N_3602);
or U3740 (N_3740,N_3525,N_3587);
nand U3741 (N_3741,N_3545,N_3522);
and U3742 (N_3742,N_3504,N_3521);
xnor U3743 (N_3743,N_3575,N_3566);
and U3744 (N_3744,N_3585,N_3525);
xor U3745 (N_3745,N_3565,N_3547);
nor U3746 (N_3746,N_3543,N_3539);
or U3747 (N_3747,N_3615,N_3554);
xor U3748 (N_3748,N_3567,N_3510);
xor U3749 (N_3749,N_3527,N_3540);
nand U3750 (N_3750,N_3640,N_3691);
or U3751 (N_3751,N_3684,N_3629);
nand U3752 (N_3752,N_3733,N_3678);
nand U3753 (N_3753,N_3682,N_3677);
and U3754 (N_3754,N_3662,N_3741);
or U3755 (N_3755,N_3713,N_3749);
xnor U3756 (N_3756,N_3699,N_3739);
nor U3757 (N_3757,N_3709,N_3645);
and U3758 (N_3758,N_3743,N_3628);
nor U3759 (N_3759,N_3666,N_3663);
or U3760 (N_3760,N_3676,N_3675);
and U3761 (N_3761,N_3703,N_3748);
and U3762 (N_3762,N_3747,N_3670);
or U3763 (N_3763,N_3639,N_3679);
or U3764 (N_3764,N_3723,N_3731);
or U3765 (N_3765,N_3742,N_3710);
or U3766 (N_3766,N_3659,N_3664);
nor U3767 (N_3767,N_3651,N_3634);
nor U3768 (N_3768,N_3665,N_3642);
nor U3769 (N_3769,N_3697,N_3727);
and U3770 (N_3770,N_3625,N_3717);
and U3771 (N_3771,N_3744,N_3673);
xor U3772 (N_3772,N_3732,N_3680);
and U3773 (N_3773,N_3657,N_3658);
xnor U3774 (N_3774,N_3722,N_3653);
and U3775 (N_3775,N_3715,N_3668);
and U3776 (N_3776,N_3729,N_3650);
nand U3777 (N_3777,N_3736,N_3745);
or U3778 (N_3778,N_3704,N_3626);
nand U3779 (N_3779,N_3708,N_3646);
and U3780 (N_3780,N_3737,N_3740);
or U3781 (N_3781,N_3735,N_3654);
nor U3782 (N_3782,N_3672,N_3647);
or U3783 (N_3783,N_3730,N_3649);
nand U3784 (N_3784,N_3716,N_3714);
xor U3785 (N_3785,N_3683,N_3655);
or U3786 (N_3786,N_3667,N_3725);
or U3787 (N_3787,N_3643,N_3701);
nand U3788 (N_3788,N_3636,N_3706);
and U3789 (N_3789,N_3702,N_3746);
xor U3790 (N_3790,N_3671,N_3630);
or U3791 (N_3791,N_3656,N_3631);
xnor U3792 (N_3792,N_3681,N_3648);
and U3793 (N_3793,N_3728,N_3738);
nand U3794 (N_3794,N_3700,N_3652);
and U3795 (N_3795,N_3638,N_3711);
nor U3796 (N_3796,N_3660,N_3692);
or U3797 (N_3797,N_3687,N_3685);
nand U3798 (N_3798,N_3635,N_3724);
or U3799 (N_3799,N_3633,N_3669);
or U3800 (N_3800,N_3695,N_3720);
nand U3801 (N_3801,N_3734,N_3688);
nand U3802 (N_3802,N_3707,N_3632);
nor U3803 (N_3803,N_3726,N_3686);
nand U3804 (N_3804,N_3637,N_3661);
and U3805 (N_3805,N_3689,N_3627);
and U3806 (N_3806,N_3694,N_3705);
xor U3807 (N_3807,N_3644,N_3690);
or U3808 (N_3808,N_3696,N_3693);
and U3809 (N_3809,N_3712,N_3674);
and U3810 (N_3810,N_3641,N_3698);
and U3811 (N_3811,N_3718,N_3719);
xor U3812 (N_3812,N_3721,N_3682);
nor U3813 (N_3813,N_3691,N_3644);
nand U3814 (N_3814,N_3709,N_3696);
and U3815 (N_3815,N_3644,N_3721);
or U3816 (N_3816,N_3668,N_3709);
and U3817 (N_3817,N_3667,N_3663);
and U3818 (N_3818,N_3636,N_3676);
or U3819 (N_3819,N_3707,N_3638);
nand U3820 (N_3820,N_3729,N_3646);
or U3821 (N_3821,N_3652,N_3628);
and U3822 (N_3822,N_3657,N_3702);
or U3823 (N_3823,N_3652,N_3737);
xor U3824 (N_3824,N_3634,N_3725);
or U3825 (N_3825,N_3642,N_3726);
nor U3826 (N_3826,N_3733,N_3720);
nor U3827 (N_3827,N_3630,N_3697);
and U3828 (N_3828,N_3681,N_3696);
nand U3829 (N_3829,N_3634,N_3653);
or U3830 (N_3830,N_3746,N_3626);
xor U3831 (N_3831,N_3681,N_3656);
or U3832 (N_3832,N_3742,N_3659);
and U3833 (N_3833,N_3687,N_3663);
nor U3834 (N_3834,N_3730,N_3656);
nor U3835 (N_3835,N_3744,N_3746);
nor U3836 (N_3836,N_3736,N_3700);
or U3837 (N_3837,N_3687,N_3633);
nor U3838 (N_3838,N_3644,N_3670);
xor U3839 (N_3839,N_3701,N_3712);
nor U3840 (N_3840,N_3711,N_3677);
or U3841 (N_3841,N_3662,N_3632);
and U3842 (N_3842,N_3668,N_3684);
xnor U3843 (N_3843,N_3634,N_3679);
or U3844 (N_3844,N_3703,N_3720);
nor U3845 (N_3845,N_3632,N_3637);
and U3846 (N_3846,N_3661,N_3694);
nand U3847 (N_3847,N_3638,N_3747);
nor U3848 (N_3848,N_3661,N_3720);
or U3849 (N_3849,N_3687,N_3701);
nor U3850 (N_3850,N_3744,N_3650);
xnor U3851 (N_3851,N_3693,N_3660);
or U3852 (N_3852,N_3682,N_3728);
and U3853 (N_3853,N_3729,N_3707);
and U3854 (N_3854,N_3703,N_3677);
xor U3855 (N_3855,N_3711,N_3669);
and U3856 (N_3856,N_3716,N_3680);
xor U3857 (N_3857,N_3701,N_3634);
or U3858 (N_3858,N_3736,N_3659);
or U3859 (N_3859,N_3742,N_3677);
nand U3860 (N_3860,N_3676,N_3742);
or U3861 (N_3861,N_3695,N_3688);
and U3862 (N_3862,N_3748,N_3667);
nor U3863 (N_3863,N_3725,N_3737);
and U3864 (N_3864,N_3702,N_3649);
and U3865 (N_3865,N_3749,N_3665);
nand U3866 (N_3866,N_3742,N_3665);
or U3867 (N_3867,N_3675,N_3717);
xnor U3868 (N_3868,N_3718,N_3676);
xnor U3869 (N_3869,N_3657,N_3663);
and U3870 (N_3870,N_3698,N_3632);
xnor U3871 (N_3871,N_3748,N_3697);
and U3872 (N_3872,N_3721,N_3648);
or U3873 (N_3873,N_3671,N_3706);
xnor U3874 (N_3874,N_3652,N_3728);
or U3875 (N_3875,N_3766,N_3833);
nor U3876 (N_3876,N_3790,N_3847);
nand U3877 (N_3877,N_3852,N_3822);
or U3878 (N_3878,N_3785,N_3853);
nor U3879 (N_3879,N_3830,N_3816);
nor U3880 (N_3880,N_3831,N_3821);
and U3881 (N_3881,N_3820,N_3796);
and U3882 (N_3882,N_3756,N_3818);
or U3883 (N_3883,N_3841,N_3800);
xor U3884 (N_3884,N_3802,N_3771);
nor U3885 (N_3885,N_3773,N_3812);
nand U3886 (N_3886,N_3823,N_3786);
nand U3887 (N_3887,N_3778,N_3836);
or U3888 (N_3888,N_3770,N_3867);
or U3889 (N_3889,N_3835,N_3845);
nor U3890 (N_3890,N_3783,N_3752);
and U3891 (N_3891,N_3848,N_3763);
or U3892 (N_3892,N_3827,N_3750);
or U3893 (N_3893,N_3779,N_3811);
or U3894 (N_3894,N_3858,N_3799);
and U3895 (N_3895,N_3832,N_3759);
nand U3896 (N_3896,N_3774,N_3804);
nand U3897 (N_3897,N_3844,N_3767);
and U3898 (N_3898,N_3859,N_3828);
or U3899 (N_3899,N_3775,N_3871);
and U3900 (N_3900,N_3757,N_3817);
nor U3901 (N_3901,N_3872,N_3815);
or U3902 (N_3902,N_3810,N_3764);
or U3903 (N_3903,N_3795,N_3793);
nand U3904 (N_3904,N_3792,N_3824);
nand U3905 (N_3905,N_3761,N_3861);
or U3906 (N_3906,N_3806,N_3753);
nand U3907 (N_3907,N_3826,N_3851);
xor U3908 (N_3908,N_3755,N_3758);
nor U3909 (N_3909,N_3814,N_3854);
nor U3910 (N_3910,N_3808,N_3784);
xor U3911 (N_3911,N_3798,N_3754);
and U3912 (N_3912,N_3838,N_3801);
or U3913 (N_3913,N_3834,N_3865);
nor U3914 (N_3914,N_3768,N_3807);
nand U3915 (N_3915,N_3856,N_3864);
or U3916 (N_3916,N_3840,N_3781);
and U3917 (N_3917,N_3839,N_3843);
or U3918 (N_3918,N_3780,N_3849);
and U3919 (N_3919,N_3829,N_3837);
or U3920 (N_3920,N_3776,N_3825);
nor U3921 (N_3921,N_3751,N_3809);
nand U3922 (N_3922,N_3862,N_3857);
xor U3923 (N_3923,N_3772,N_3791);
and U3924 (N_3924,N_3787,N_3769);
xnor U3925 (N_3925,N_3777,N_3794);
or U3926 (N_3926,N_3765,N_3805);
or U3927 (N_3927,N_3873,N_3870);
and U3928 (N_3928,N_3860,N_3855);
xor U3929 (N_3929,N_3813,N_3863);
and U3930 (N_3930,N_3866,N_3782);
nand U3931 (N_3931,N_3869,N_3788);
nand U3932 (N_3932,N_3819,N_3762);
and U3933 (N_3933,N_3868,N_3797);
nand U3934 (N_3934,N_3789,N_3846);
nand U3935 (N_3935,N_3874,N_3850);
xnor U3936 (N_3936,N_3803,N_3842);
and U3937 (N_3937,N_3760,N_3785);
or U3938 (N_3938,N_3787,N_3803);
nand U3939 (N_3939,N_3846,N_3779);
or U3940 (N_3940,N_3820,N_3753);
and U3941 (N_3941,N_3783,N_3785);
and U3942 (N_3942,N_3768,N_3865);
and U3943 (N_3943,N_3846,N_3862);
nand U3944 (N_3944,N_3797,N_3810);
nand U3945 (N_3945,N_3752,N_3753);
nand U3946 (N_3946,N_3859,N_3762);
xor U3947 (N_3947,N_3781,N_3839);
and U3948 (N_3948,N_3873,N_3858);
or U3949 (N_3949,N_3804,N_3860);
nor U3950 (N_3950,N_3829,N_3806);
or U3951 (N_3951,N_3850,N_3823);
xor U3952 (N_3952,N_3817,N_3756);
xnor U3953 (N_3953,N_3821,N_3815);
or U3954 (N_3954,N_3828,N_3785);
or U3955 (N_3955,N_3796,N_3857);
xor U3956 (N_3956,N_3826,N_3755);
nor U3957 (N_3957,N_3777,N_3855);
nor U3958 (N_3958,N_3867,N_3774);
nand U3959 (N_3959,N_3820,N_3855);
and U3960 (N_3960,N_3814,N_3873);
xnor U3961 (N_3961,N_3785,N_3862);
nand U3962 (N_3962,N_3826,N_3872);
and U3963 (N_3963,N_3833,N_3858);
or U3964 (N_3964,N_3835,N_3853);
or U3965 (N_3965,N_3838,N_3791);
nor U3966 (N_3966,N_3764,N_3851);
nand U3967 (N_3967,N_3784,N_3768);
or U3968 (N_3968,N_3856,N_3767);
xor U3969 (N_3969,N_3821,N_3809);
xnor U3970 (N_3970,N_3750,N_3850);
and U3971 (N_3971,N_3818,N_3833);
nor U3972 (N_3972,N_3867,N_3843);
and U3973 (N_3973,N_3810,N_3873);
and U3974 (N_3974,N_3772,N_3796);
and U3975 (N_3975,N_3757,N_3803);
and U3976 (N_3976,N_3771,N_3766);
nor U3977 (N_3977,N_3870,N_3781);
and U3978 (N_3978,N_3820,N_3833);
or U3979 (N_3979,N_3824,N_3849);
and U3980 (N_3980,N_3758,N_3821);
or U3981 (N_3981,N_3864,N_3840);
nand U3982 (N_3982,N_3846,N_3780);
nand U3983 (N_3983,N_3779,N_3857);
and U3984 (N_3984,N_3757,N_3849);
and U3985 (N_3985,N_3803,N_3784);
nor U3986 (N_3986,N_3854,N_3755);
and U3987 (N_3987,N_3808,N_3840);
or U3988 (N_3988,N_3791,N_3865);
nand U3989 (N_3989,N_3830,N_3800);
or U3990 (N_3990,N_3799,N_3754);
nor U3991 (N_3991,N_3870,N_3840);
nor U3992 (N_3992,N_3833,N_3872);
and U3993 (N_3993,N_3755,N_3787);
and U3994 (N_3994,N_3787,N_3824);
or U3995 (N_3995,N_3856,N_3761);
or U3996 (N_3996,N_3754,N_3806);
xor U3997 (N_3997,N_3839,N_3811);
nor U3998 (N_3998,N_3786,N_3792);
nand U3999 (N_3999,N_3856,N_3781);
xnor U4000 (N_4000,N_3876,N_3951);
or U4001 (N_4001,N_3920,N_3939);
and U4002 (N_4002,N_3993,N_3917);
nand U4003 (N_4003,N_3954,N_3934);
nor U4004 (N_4004,N_3879,N_3964);
or U4005 (N_4005,N_3947,N_3949);
xnor U4006 (N_4006,N_3878,N_3908);
nand U4007 (N_4007,N_3907,N_3972);
or U4008 (N_4008,N_3891,N_3959);
xnor U4009 (N_4009,N_3890,N_3960);
xnor U4010 (N_4010,N_3880,N_3906);
nor U4011 (N_4011,N_3902,N_3977);
and U4012 (N_4012,N_3978,N_3999);
nand U4013 (N_4013,N_3888,N_3897);
and U4014 (N_4014,N_3982,N_3950);
and U4015 (N_4015,N_3941,N_3962);
and U4016 (N_4016,N_3905,N_3930);
nand U4017 (N_4017,N_3929,N_3928);
nor U4018 (N_4018,N_3958,N_3955);
xnor U4019 (N_4019,N_3925,N_3995);
and U4020 (N_4020,N_3985,N_3961);
and U4021 (N_4021,N_3882,N_3889);
xnor U4022 (N_4022,N_3914,N_3916);
or U4023 (N_4023,N_3921,N_3927);
nor U4024 (N_4024,N_3983,N_3967);
nor U4025 (N_4025,N_3957,N_3994);
xor U4026 (N_4026,N_3909,N_3886);
xnor U4027 (N_4027,N_3988,N_3901);
nand U4028 (N_4028,N_3919,N_3979);
nor U4029 (N_4029,N_3948,N_3936);
xor U4030 (N_4030,N_3974,N_3942);
xor U4031 (N_4031,N_3912,N_3900);
xnor U4032 (N_4032,N_3932,N_3911);
nor U4033 (N_4033,N_3894,N_3981);
or U4034 (N_4034,N_3980,N_3931);
xor U4035 (N_4035,N_3943,N_3935);
xor U4036 (N_4036,N_3998,N_3991);
or U4037 (N_4037,N_3997,N_3933);
nor U4038 (N_4038,N_3968,N_3915);
and U4039 (N_4039,N_3944,N_3904);
xor U4040 (N_4040,N_3945,N_3965);
or U4041 (N_4041,N_3883,N_3913);
and U4042 (N_4042,N_3956,N_3918);
nor U4043 (N_4043,N_3973,N_3989);
xor U4044 (N_4044,N_3899,N_3953);
nand U4045 (N_4045,N_3893,N_3924);
and U4046 (N_4046,N_3963,N_3884);
xor U4047 (N_4047,N_3896,N_3992);
nand U4048 (N_4048,N_3976,N_3937);
xnor U4049 (N_4049,N_3966,N_3969);
or U4050 (N_4050,N_3898,N_3881);
and U4051 (N_4051,N_3986,N_3984);
nand U4052 (N_4052,N_3987,N_3938);
and U4053 (N_4053,N_3946,N_3975);
nor U4054 (N_4054,N_3892,N_3923);
or U4055 (N_4055,N_3877,N_3895);
nor U4056 (N_4056,N_3910,N_3996);
or U4057 (N_4057,N_3970,N_3952);
xor U4058 (N_4058,N_3971,N_3885);
nand U4059 (N_4059,N_3926,N_3990);
nand U4060 (N_4060,N_3903,N_3875);
xnor U4061 (N_4061,N_3922,N_3940);
and U4062 (N_4062,N_3887,N_3913);
xor U4063 (N_4063,N_3945,N_3975);
and U4064 (N_4064,N_3957,N_3917);
or U4065 (N_4065,N_3992,N_3975);
nand U4066 (N_4066,N_3895,N_3985);
or U4067 (N_4067,N_3950,N_3895);
or U4068 (N_4068,N_3940,N_3957);
nor U4069 (N_4069,N_3917,N_3975);
nor U4070 (N_4070,N_3888,N_3907);
nor U4071 (N_4071,N_3963,N_3924);
xnor U4072 (N_4072,N_3945,N_3910);
nand U4073 (N_4073,N_3992,N_3933);
and U4074 (N_4074,N_3934,N_3889);
xor U4075 (N_4075,N_3989,N_3923);
nand U4076 (N_4076,N_3913,N_3892);
and U4077 (N_4077,N_3999,N_3898);
nand U4078 (N_4078,N_3934,N_3877);
xor U4079 (N_4079,N_3897,N_3933);
and U4080 (N_4080,N_3988,N_3967);
and U4081 (N_4081,N_3904,N_3937);
nand U4082 (N_4082,N_3883,N_3896);
xnor U4083 (N_4083,N_3991,N_3929);
nand U4084 (N_4084,N_3880,N_3992);
nor U4085 (N_4085,N_3997,N_3919);
and U4086 (N_4086,N_3971,N_3945);
and U4087 (N_4087,N_3982,N_3956);
xor U4088 (N_4088,N_3941,N_3985);
xnor U4089 (N_4089,N_3943,N_3939);
xnor U4090 (N_4090,N_3967,N_3908);
and U4091 (N_4091,N_3942,N_3879);
nand U4092 (N_4092,N_3981,N_3943);
and U4093 (N_4093,N_3905,N_3927);
nand U4094 (N_4094,N_3881,N_3903);
nand U4095 (N_4095,N_3907,N_3984);
nand U4096 (N_4096,N_3985,N_3931);
xnor U4097 (N_4097,N_3948,N_3923);
xor U4098 (N_4098,N_3941,N_3875);
xnor U4099 (N_4099,N_3918,N_3961);
xor U4100 (N_4100,N_3998,N_3934);
and U4101 (N_4101,N_3910,N_3999);
nand U4102 (N_4102,N_3949,N_3889);
or U4103 (N_4103,N_3882,N_3930);
nor U4104 (N_4104,N_3878,N_3877);
nor U4105 (N_4105,N_3908,N_3995);
and U4106 (N_4106,N_3997,N_3907);
or U4107 (N_4107,N_3905,N_3981);
nor U4108 (N_4108,N_3913,N_3914);
nor U4109 (N_4109,N_3948,N_3911);
nor U4110 (N_4110,N_3948,N_3977);
nand U4111 (N_4111,N_3910,N_3886);
xnor U4112 (N_4112,N_3902,N_3889);
or U4113 (N_4113,N_3877,N_3976);
or U4114 (N_4114,N_3941,N_3973);
xnor U4115 (N_4115,N_3938,N_3901);
nor U4116 (N_4116,N_3931,N_3876);
or U4117 (N_4117,N_3913,N_3961);
xor U4118 (N_4118,N_3911,N_3884);
nand U4119 (N_4119,N_3891,N_3972);
xor U4120 (N_4120,N_3937,N_3920);
or U4121 (N_4121,N_3979,N_3904);
nand U4122 (N_4122,N_3889,N_3917);
and U4123 (N_4123,N_3880,N_3888);
nor U4124 (N_4124,N_3951,N_3882);
and U4125 (N_4125,N_4025,N_4071);
nor U4126 (N_4126,N_4087,N_4064);
and U4127 (N_4127,N_4031,N_4054);
nor U4128 (N_4128,N_4003,N_4102);
nor U4129 (N_4129,N_4030,N_4088);
xnor U4130 (N_4130,N_4018,N_4084);
nand U4131 (N_4131,N_4050,N_4020);
and U4132 (N_4132,N_4067,N_4058);
nor U4133 (N_4133,N_4013,N_4118);
nand U4134 (N_4134,N_4093,N_4035);
xor U4135 (N_4135,N_4110,N_4097);
nor U4136 (N_4136,N_4032,N_4076);
nand U4137 (N_4137,N_4012,N_4055);
nand U4138 (N_4138,N_4016,N_4060);
xnor U4139 (N_4139,N_4099,N_4057);
and U4140 (N_4140,N_4123,N_4052);
xnor U4141 (N_4141,N_4002,N_4072);
and U4142 (N_4142,N_4065,N_4029);
or U4143 (N_4143,N_4090,N_4021);
nor U4144 (N_4144,N_4019,N_4045);
and U4145 (N_4145,N_4038,N_4080);
nand U4146 (N_4146,N_4047,N_4112);
or U4147 (N_4147,N_4092,N_4005);
xnor U4148 (N_4148,N_4006,N_4083);
nor U4149 (N_4149,N_4028,N_4024);
nor U4150 (N_4150,N_4100,N_4078);
xnor U4151 (N_4151,N_4051,N_4027);
or U4152 (N_4152,N_4040,N_4042);
nor U4153 (N_4153,N_4091,N_4011);
nor U4154 (N_4154,N_4023,N_4056);
nor U4155 (N_4155,N_4108,N_4074);
nor U4156 (N_4156,N_4059,N_4075);
or U4157 (N_4157,N_4022,N_4119);
xnor U4158 (N_4158,N_4120,N_4086);
nor U4159 (N_4159,N_4098,N_4033);
and U4160 (N_4160,N_4026,N_4079);
nor U4161 (N_4161,N_4077,N_4053);
and U4162 (N_4162,N_4103,N_4000);
and U4163 (N_4163,N_4082,N_4007);
or U4164 (N_4164,N_4117,N_4122);
and U4165 (N_4165,N_4089,N_4116);
nor U4166 (N_4166,N_4094,N_4069);
nand U4167 (N_4167,N_4043,N_4081);
xnor U4168 (N_4168,N_4017,N_4073);
and U4169 (N_4169,N_4046,N_4044);
or U4170 (N_4170,N_4115,N_4085);
nor U4171 (N_4171,N_4124,N_4004);
xor U4172 (N_4172,N_4014,N_4104);
or U4173 (N_4173,N_4096,N_4062);
nand U4174 (N_4174,N_4070,N_4010);
or U4175 (N_4175,N_4105,N_4037);
or U4176 (N_4176,N_4063,N_4107);
nor U4177 (N_4177,N_4106,N_4111);
xor U4178 (N_4178,N_4036,N_4041);
xnor U4179 (N_4179,N_4034,N_4101);
xor U4180 (N_4180,N_4095,N_4121);
nor U4181 (N_4181,N_4049,N_4114);
and U4182 (N_4182,N_4068,N_4039);
nand U4183 (N_4183,N_4009,N_4008);
nor U4184 (N_4184,N_4048,N_4113);
nor U4185 (N_4185,N_4015,N_4109);
nand U4186 (N_4186,N_4061,N_4001);
and U4187 (N_4187,N_4066,N_4016);
or U4188 (N_4188,N_4117,N_4114);
or U4189 (N_4189,N_4030,N_4084);
xor U4190 (N_4190,N_4054,N_4085);
nand U4191 (N_4191,N_4072,N_4021);
or U4192 (N_4192,N_4110,N_4008);
or U4193 (N_4193,N_4062,N_4123);
and U4194 (N_4194,N_4058,N_4115);
nor U4195 (N_4195,N_4071,N_4054);
and U4196 (N_4196,N_4100,N_4109);
nand U4197 (N_4197,N_4058,N_4014);
nand U4198 (N_4198,N_4103,N_4121);
nor U4199 (N_4199,N_4026,N_4108);
nand U4200 (N_4200,N_4092,N_4051);
and U4201 (N_4201,N_4113,N_4087);
or U4202 (N_4202,N_4095,N_4100);
xnor U4203 (N_4203,N_4046,N_4005);
and U4204 (N_4204,N_4006,N_4004);
and U4205 (N_4205,N_4001,N_4015);
nor U4206 (N_4206,N_4041,N_4032);
and U4207 (N_4207,N_4004,N_4106);
and U4208 (N_4208,N_4025,N_4080);
and U4209 (N_4209,N_4004,N_4070);
or U4210 (N_4210,N_4099,N_4092);
xor U4211 (N_4211,N_4061,N_4120);
nand U4212 (N_4212,N_4022,N_4006);
nor U4213 (N_4213,N_4052,N_4073);
nand U4214 (N_4214,N_4029,N_4027);
and U4215 (N_4215,N_4123,N_4087);
or U4216 (N_4216,N_4104,N_4027);
xor U4217 (N_4217,N_4021,N_4010);
xor U4218 (N_4218,N_4088,N_4109);
nor U4219 (N_4219,N_4023,N_4116);
and U4220 (N_4220,N_4115,N_4012);
nor U4221 (N_4221,N_4032,N_4025);
or U4222 (N_4222,N_4044,N_4021);
xnor U4223 (N_4223,N_4096,N_4073);
nand U4224 (N_4224,N_4124,N_4036);
and U4225 (N_4225,N_4110,N_4045);
nand U4226 (N_4226,N_4035,N_4090);
or U4227 (N_4227,N_4096,N_4032);
and U4228 (N_4228,N_4066,N_4099);
nand U4229 (N_4229,N_4113,N_4114);
and U4230 (N_4230,N_4118,N_4091);
xnor U4231 (N_4231,N_4040,N_4102);
xor U4232 (N_4232,N_4041,N_4103);
nand U4233 (N_4233,N_4093,N_4006);
xnor U4234 (N_4234,N_4090,N_4031);
and U4235 (N_4235,N_4035,N_4047);
or U4236 (N_4236,N_4006,N_4088);
and U4237 (N_4237,N_4119,N_4091);
or U4238 (N_4238,N_4123,N_4023);
and U4239 (N_4239,N_4060,N_4012);
or U4240 (N_4240,N_4096,N_4020);
and U4241 (N_4241,N_4062,N_4084);
nand U4242 (N_4242,N_4069,N_4087);
nor U4243 (N_4243,N_4031,N_4113);
xnor U4244 (N_4244,N_4117,N_4060);
xnor U4245 (N_4245,N_4119,N_4007);
nand U4246 (N_4246,N_4033,N_4011);
nand U4247 (N_4247,N_4040,N_4037);
or U4248 (N_4248,N_4000,N_4098);
or U4249 (N_4249,N_4055,N_4049);
nand U4250 (N_4250,N_4175,N_4127);
nor U4251 (N_4251,N_4188,N_4199);
or U4252 (N_4252,N_4174,N_4208);
nand U4253 (N_4253,N_4240,N_4130);
or U4254 (N_4254,N_4142,N_4219);
nand U4255 (N_4255,N_4231,N_4221);
xnor U4256 (N_4256,N_4166,N_4220);
xor U4257 (N_4257,N_4152,N_4177);
nand U4258 (N_4258,N_4209,N_4211);
and U4259 (N_4259,N_4191,N_4162);
and U4260 (N_4260,N_4150,N_4195);
nor U4261 (N_4261,N_4203,N_4238);
and U4262 (N_4262,N_4168,N_4244);
nor U4263 (N_4263,N_4228,N_4146);
and U4264 (N_4264,N_4245,N_4131);
xor U4265 (N_4265,N_4249,N_4197);
and U4266 (N_4266,N_4200,N_4171);
nor U4267 (N_4267,N_4212,N_4213);
xnor U4268 (N_4268,N_4234,N_4140);
nand U4269 (N_4269,N_4141,N_4216);
nand U4270 (N_4270,N_4187,N_4242);
or U4271 (N_4271,N_4126,N_4155);
xnor U4272 (N_4272,N_4204,N_4210);
nor U4273 (N_4273,N_4205,N_4201);
nand U4274 (N_4274,N_4158,N_4239);
nand U4275 (N_4275,N_4223,N_4170);
nand U4276 (N_4276,N_4176,N_4198);
nand U4277 (N_4277,N_4129,N_4215);
nor U4278 (N_4278,N_4139,N_4151);
nand U4279 (N_4279,N_4143,N_4226);
xor U4280 (N_4280,N_4179,N_4233);
or U4281 (N_4281,N_4149,N_4181);
or U4282 (N_4282,N_4194,N_4132);
and U4283 (N_4283,N_4164,N_4207);
xnor U4284 (N_4284,N_4165,N_4243);
nor U4285 (N_4285,N_4144,N_4182);
and U4286 (N_4286,N_4167,N_4237);
and U4287 (N_4287,N_4128,N_4134);
nor U4288 (N_4288,N_4225,N_4232);
and U4289 (N_4289,N_4138,N_4180);
or U4290 (N_4290,N_4222,N_4247);
xnor U4291 (N_4291,N_4192,N_4133);
nor U4292 (N_4292,N_4246,N_4235);
nor U4293 (N_4293,N_4229,N_4227);
and U4294 (N_4294,N_4173,N_4248);
and U4295 (N_4295,N_4136,N_4178);
nand U4296 (N_4296,N_4153,N_4236);
nor U4297 (N_4297,N_4224,N_4202);
nand U4298 (N_4298,N_4169,N_4183);
nand U4299 (N_4299,N_4125,N_4190);
and U4300 (N_4300,N_4218,N_4148);
nand U4301 (N_4301,N_4206,N_4214);
and U4302 (N_4302,N_4241,N_4157);
nor U4303 (N_4303,N_4185,N_4147);
or U4304 (N_4304,N_4184,N_4160);
nand U4305 (N_4305,N_4135,N_4230);
or U4306 (N_4306,N_4172,N_4137);
nor U4307 (N_4307,N_4189,N_4163);
or U4308 (N_4308,N_4217,N_4154);
nand U4309 (N_4309,N_4159,N_4145);
xnor U4310 (N_4310,N_4196,N_4156);
nor U4311 (N_4311,N_4193,N_4161);
and U4312 (N_4312,N_4186,N_4139);
and U4313 (N_4313,N_4249,N_4159);
and U4314 (N_4314,N_4133,N_4153);
or U4315 (N_4315,N_4236,N_4219);
nand U4316 (N_4316,N_4249,N_4175);
nor U4317 (N_4317,N_4224,N_4128);
and U4318 (N_4318,N_4179,N_4224);
nand U4319 (N_4319,N_4148,N_4244);
nor U4320 (N_4320,N_4143,N_4146);
nand U4321 (N_4321,N_4154,N_4202);
nor U4322 (N_4322,N_4223,N_4166);
nor U4323 (N_4323,N_4204,N_4217);
nand U4324 (N_4324,N_4164,N_4197);
or U4325 (N_4325,N_4226,N_4242);
and U4326 (N_4326,N_4129,N_4137);
and U4327 (N_4327,N_4156,N_4206);
and U4328 (N_4328,N_4241,N_4190);
and U4329 (N_4329,N_4240,N_4150);
nor U4330 (N_4330,N_4204,N_4234);
nor U4331 (N_4331,N_4243,N_4236);
xnor U4332 (N_4332,N_4142,N_4140);
nand U4333 (N_4333,N_4209,N_4189);
nor U4334 (N_4334,N_4155,N_4145);
xor U4335 (N_4335,N_4245,N_4128);
or U4336 (N_4336,N_4239,N_4148);
nor U4337 (N_4337,N_4162,N_4227);
nand U4338 (N_4338,N_4129,N_4125);
nand U4339 (N_4339,N_4206,N_4235);
and U4340 (N_4340,N_4194,N_4171);
nand U4341 (N_4341,N_4207,N_4133);
nand U4342 (N_4342,N_4211,N_4199);
and U4343 (N_4343,N_4132,N_4225);
and U4344 (N_4344,N_4195,N_4173);
or U4345 (N_4345,N_4237,N_4193);
or U4346 (N_4346,N_4204,N_4225);
xnor U4347 (N_4347,N_4228,N_4163);
xor U4348 (N_4348,N_4182,N_4127);
xor U4349 (N_4349,N_4232,N_4219);
xor U4350 (N_4350,N_4239,N_4195);
and U4351 (N_4351,N_4227,N_4145);
and U4352 (N_4352,N_4247,N_4212);
nor U4353 (N_4353,N_4234,N_4136);
and U4354 (N_4354,N_4143,N_4163);
nor U4355 (N_4355,N_4190,N_4159);
and U4356 (N_4356,N_4168,N_4150);
xnor U4357 (N_4357,N_4219,N_4203);
nand U4358 (N_4358,N_4142,N_4172);
nand U4359 (N_4359,N_4235,N_4223);
or U4360 (N_4360,N_4187,N_4162);
and U4361 (N_4361,N_4164,N_4171);
xor U4362 (N_4362,N_4234,N_4177);
nor U4363 (N_4363,N_4162,N_4204);
or U4364 (N_4364,N_4211,N_4154);
xor U4365 (N_4365,N_4219,N_4183);
xor U4366 (N_4366,N_4202,N_4226);
nor U4367 (N_4367,N_4201,N_4160);
xnor U4368 (N_4368,N_4229,N_4153);
nand U4369 (N_4369,N_4216,N_4222);
xor U4370 (N_4370,N_4212,N_4175);
and U4371 (N_4371,N_4226,N_4205);
xor U4372 (N_4372,N_4227,N_4172);
xor U4373 (N_4373,N_4241,N_4201);
xnor U4374 (N_4374,N_4135,N_4150);
nor U4375 (N_4375,N_4294,N_4354);
xor U4376 (N_4376,N_4252,N_4337);
nor U4377 (N_4377,N_4339,N_4343);
nor U4378 (N_4378,N_4311,N_4319);
xor U4379 (N_4379,N_4361,N_4324);
and U4380 (N_4380,N_4342,N_4272);
or U4381 (N_4381,N_4291,N_4364);
nor U4382 (N_4382,N_4279,N_4312);
or U4383 (N_4383,N_4287,N_4340);
and U4384 (N_4384,N_4258,N_4273);
nand U4385 (N_4385,N_4321,N_4269);
xor U4386 (N_4386,N_4282,N_4274);
nand U4387 (N_4387,N_4322,N_4281);
and U4388 (N_4388,N_4356,N_4261);
nand U4389 (N_4389,N_4346,N_4316);
or U4390 (N_4390,N_4367,N_4357);
or U4391 (N_4391,N_4338,N_4265);
xor U4392 (N_4392,N_4309,N_4296);
or U4393 (N_4393,N_4302,N_4353);
and U4394 (N_4394,N_4355,N_4351);
nand U4395 (N_4395,N_4326,N_4292);
or U4396 (N_4396,N_4257,N_4283);
nand U4397 (N_4397,N_4251,N_4320);
nor U4398 (N_4398,N_4371,N_4373);
or U4399 (N_4399,N_4350,N_4307);
and U4400 (N_4400,N_4331,N_4332);
xnor U4401 (N_4401,N_4365,N_4275);
xor U4402 (N_4402,N_4254,N_4317);
xor U4403 (N_4403,N_4266,N_4336);
nor U4404 (N_4404,N_4306,N_4341);
nand U4405 (N_4405,N_4370,N_4334);
and U4406 (N_4406,N_4358,N_4263);
nand U4407 (N_4407,N_4288,N_4284);
or U4408 (N_4408,N_4369,N_4285);
xnor U4409 (N_4409,N_4260,N_4277);
nand U4410 (N_4410,N_4325,N_4308);
nor U4411 (N_4411,N_4295,N_4335);
nor U4412 (N_4412,N_4278,N_4368);
nor U4413 (N_4413,N_4360,N_4255);
xnor U4414 (N_4414,N_4289,N_4333);
or U4415 (N_4415,N_4256,N_4276);
and U4416 (N_4416,N_4344,N_4298);
or U4417 (N_4417,N_4327,N_4348);
and U4418 (N_4418,N_4270,N_4299);
and U4419 (N_4419,N_4349,N_4323);
xnor U4420 (N_4420,N_4318,N_4345);
nand U4421 (N_4421,N_4330,N_4259);
nor U4422 (N_4422,N_4314,N_4253);
nor U4423 (N_4423,N_4271,N_4303);
or U4424 (N_4424,N_4290,N_4286);
or U4425 (N_4425,N_4352,N_4366);
xor U4426 (N_4426,N_4359,N_4305);
and U4427 (N_4427,N_4297,N_4300);
nand U4428 (N_4428,N_4363,N_4264);
nor U4429 (N_4429,N_4293,N_4328);
xor U4430 (N_4430,N_4304,N_4362);
and U4431 (N_4431,N_4267,N_4372);
nor U4432 (N_4432,N_4315,N_4310);
or U4433 (N_4433,N_4280,N_4301);
or U4434 (N_4434,N_4374,N_4262);
nand U4435 (N_4435,N_4313,N_4329);
or U4436 (N_4436,N_4250,N_4347);
and U4437 (N_4437,N_4268,N_4314);
nor U4438 (N_4438,N_4254,N_4353);
nand U4439 (N_4439,N_4331,N_4305);
nand U4440 (N_4440,N_4340,N_4367);
xor U4441 (N_4441,N_4263,N_4260);
and U4442 (N_4442,N_4328,N_4319);
nor U4443 (N_4443,N_4331,N_4328);
xnor U4444 (N_4444,N_4332,N_4297);
and U4445 (N_4445,N_4339,N_4349);
xor U4446 (N_4446,N_4343,N_4280);
and U4447 (N_4447,N_4320,N_4282);
xor U4448 (N_4448,N_4269,N_4284);
xnor U4449 (N_4449,N_4343,N_4366);
and U4450 (N_4450,N_4280,N_4327);
xor U4451 (N_4451,N_4363,N_4316);
nor U4452 (N_4452,N_4370,N_4285);
nor U4453 (N_4453,N_4269,N_4334);
xnor U4454 (N_4454,N_4251,N_4280);
or U4455 (N_4455,N_4260,N_4358);
or U4456 (N_4456,N_4292,N_4304);
nand U4457 (N_4457,N_4276,N_4265);
nand U4458 (N_4458,N_4288,N_4345);
xnor U4459 (N_4459,N_4316,N_4320);
xnor U4460 (N_4460,N_4357,N_4312);
or U4461 (N_4461,N_4307,N_4311);
nor U4462 (N_4462,N_4318,N_4254);
nor U4463 (N_4463,N_4293,N_4299);
nand U4464 (N_4464,N_4282,N_4289);
nor U4465 (N_4465,N_4262,N_4353);
nand U4466 (N_4466,N_4330,N_4253);
nor U4467 (N_4467,N_4262,N_4326);
nand U4468 (N_4468,N_4356,N_4346);
nand U4469 (N_4469,N_4327,N_4369);
nand U4470 (N_4470,N_4345,N_4278);
xnor U4471 (N_4471,N_4350,N_4338);
nand U4472 (N_4472,N_4281,N_4335);
nand U4473 (N_4473,N_4339,N_4324);
nor U4474 (N_4474,N_4350,N_4351);
and U4475 (N_4475,N_4295,N_4263);
and U4476 (N_4476,N_4308,N_4333);
nor U4477 (N_4477,N_4373,N_4326);
nand U4478 (N_4478,N_4298,N_4337);
nor U4479 (N_4479,N_4286,N_4352);
and U4480 (N_4480,N_4334,N_4367);
or U4481 (N_4481,N_4369,N_4309);
nor U4482 (N_4482,N_4289,N_4254);
and U4483 (N_4483,N_4264,N_4260);
xor U4484 (N_4484,N_4315,N_4280);
xor U4485 (N_4485,N_4267,N_4305);
xnor U4486 (N_4486,N_4263,N_4370);
or U4487 (N_4487,N_4258,N_4371);
nand U4488 (N_4488,N_4277,N_4328);
or U4489 (N_4489,N_4329,N_4268);
nor U4490 (N_4490,N_4323,N_4354);
nand U4491 (N_4491,N_4325,N_4326);
xnor U4492 (N_4492,N_4302,N_4329);
nor U4493 (N_4493,N_4348,N_4317);
xnor U4494 (N_4494,N_4349,N_4291);
and U4495 (N_4495,N_4359,N_4264);
and U4496 (N_4496,N_4340,N_4371);
nor U4497 (N_4497,N_4333,N_4364);
nand U4498 (N_4498,N_4335,N_4304);
and U4499 (N_4499,N_4264,N_4337);
xor U4500 (N_4500,N_4478,N_4460);
nor U4501 (N_4501,N_4425,N_4442);
or U4502 (N_4502,N_4407,N_4428);
nand U4503 (N_4503,N_4411,N_4483);
or U4504 (N_4504,N_4388,N_4431);
or U4505 (N_4505,N_4440,N_4406);
xnor U4506 (N_4506,N_4485,N_4392);
and U4507 (N_4507,N_4419,N_4418);
nand U4508 (N_4508,N_4393,N_4456);
nor U4509 (N_4509,N_4424,N_4401);
or U4510 (N_4510,N_4409,N_4414);
nand U4511 (N_4511,N_4399,N_4420);
or U4512 (N_4512,N_4416,N_4462);
nand U4513 (N_4513,N_4484,N_4463);
xor U4514 (N_4514,N_4492,N_4382);
xnor U4515 (N_4515,N_4412,N_4489);
nand U4516 (N_4516,N_4390,N_4479);
nor U4517 (N_4517,N_4432,N_4387);
nand U4518 (N_4518,N_4451,N_4398);
xnor U4519 (N_4519,N_4426,N_4391);
nor U4520 (N_4520,N_4400,N_4465);
xnor U4521 (N_4521,N_4452,N_4480);
nor U4522 (N_4522,N_4464,N_4453);
xnor U4523 (N_4523,N_4455,N_4430);
and U4524 (N_4524,N_4469,N_4415);
and U4525 (N_4525,N_4448,N_4395);
nand U4526 (N_4526,N_4461,N_4405);
and U4527 (N_4527,N_4454,N_4458);
nor U4528 (N_4528,N_4404,N_4408);
xnor U4529 (N_4529,N_4386,N_4421);
or U4530 (N_4530,N_4436,N_4445);
nor U4531 (N_4531,N_4423,N_4496);
xor U4532 (N_4532,N_4437,N_4477);
and U4533 (N_4533,N_4491,N_4488);
or U4534 (N_4534,N_4394,N_4433);
nand U4535 (N_4535,N_4446,N_4466);
and U4536 (N_4536,N_4385,N_4486);
xnor U4537 (N_4537,N_4449,N_4487);
xnor U4538 (N_4538,N_4441,N_4457);
nand U4539 (N_4539,N_4402,N_4435);
xnor U4540 (N_4540,N_4381,N_4396);
nand U4541 (N_4541,N_4473,N_4493);
nor U4542 (N_4542,N_4389,N_4378);
or U4543 (N_4543,N_4471,N_4495);
and U4544 (N_4544,N_4438,N_4481);
or U4545 (N_4545,N_4380,N_4384);
and U4546 (N_4546,N_4429,N_4498);
xor U4547 (N_4547,N_4490,N_4472);
nor U4548 (N_4548,N_4439,N_4444);
or U4549 (N_4549,N_4459,N_4397);
or U4550 (N_4550,N_4375,N_4482);
nand U4551 (N_4551,N_4403,N_4379);
nor U4552 (N_4552,N_4434,N_4447);
nand U4553 (N_4553,N_4383,N_4422);
nand U4554 (N_4554,N_4497,N_4410);
and U4555 (N_4555,N_4499,N_4427);
xor U4556 (N_4556,N_4417,N_4474);
or U4557 (N_4557,N_4467,N_4494);
xor U4558 (N_4558,N_4476,N_4443);
and U4559 (N_4559,N_4413,N_4470);
and U4560 (N_4560,N_4475,N_4377);
or U4561 (N_4561,N_4468,N_4450);
or U4562 (N_4562,N_4376,N_4492);
or U4563 (N_4563,N_4407,N_4375);
and U4564 (N_4564,N_4456,N_4463);
and U4565 (N_4565,N_4475,N_4459);
nor U4566 (N_4566,N_4391,N_4398);
nand U4567 (N_4567,N_4383,N_4455);
nand U4568 (N_4568,N_4460,N_4492);
nand U4569 (N_4569,N_4480,N_4398);
nand U4570 (N_4570,N_4458,N_4479);
or U4571 (N_4571,N_4408,N_4475);
nor U4572 (N_4572,N_4446,N_4386);
and U4573 (N_4573,N_4413,N_4403);
or U4574 (N_4574,N_4419,N_4440);
xor U4575 (N_4575,N_4408,N_4477);
nand U4576 (N_4576,N_4471,N_4446);
and U4577 (N_4577,N_4393,N_4405);
xnor U4578 (N_4578,N_4386,N_4462);
and U4579 (N_4579,N_4462,N_4471);
or U4580 (N_4580,N_4461,N_4385);
or U4581 (N_4581,N_4413,N_4390);
and U4582 (N_4582,N_4433,N_4409);
nor U4583 (N_4583,N_4396,N_4456);
nand U4584 (N_4584,N_4485,N_4497);
and U4585 (N_4585,N_4485,N_4411);
or U4586 (N_4586,N_4475,N_4418);
nor U4587 (N_4587,N_4464,N_4418);
nand U4588 (N_4588,N_4444,N_4495);
nand U4589 (N_4589,N_4476,N_4461);
or U4590 (N_4590,N_4435,N_4469);
nand U4591 (N_4591,N_4489,N_4395);
nor U4592 (N_4592,N_4479,N_4401);
xnor U4593 (N_4593,N_4429,N_4446);
or U4594 (N_4594,N_4478,N_4469);
nor U4595 (N_4595,N_4448,N_4426);
nor U4596 (N_4596,N_4477,N_4482);
nand U4597 (N_4597,N_4416,N_4455);
and U4598 (N_4598,N_4480,N_4485);
or U4599 (N_4599,N_4375,N_4406);
nand U4600 (N_4600,N_4420,N_4409);
nand U4601 (N_4601,N_4422,N_4445);
nand U4602 (N_4602,N_4388,N_4446);
nand U4603 (N_4603,N_4469,N_4392);
xnor U4604 (N_4604,N_4455,N_4431);
nor U4605 (N_4605,N_4376,N_4397);
nand U4606 (N_4606,N_4411,N_4439);
or U4607 (N_4607,N_4434,N_4470);
and U4608 (N_4608,N_4453,N_4410);
xor U4609 (N_4609,N_4439,N_4412);
xnor U4610 (N_4610,N_4398,N_4393);
nor U4611 (N_4611,N_4473,N_4380);
and U4612 (N_4612,N_4487,N_4461);
and U4613 (N_4613,N_4415,N_4499);
and U4614 (N_4614,N_4401,N_4460);
xnor U4615 (N_4615,N_4383,N_4404);
xor U4616 (N_4616,N_4419,N_4391);
xor U4617 (N_4617,N_4385,N_4401);
nor U4618 (N_4618,N_4495,N_4383);
xor U4619 (N_4619,N_4399,N_4437);
and U4620 (N_4620,N_4472,N_4395);
nor U4621 (N_4621,N_4472,N_4458);
and U4622 (N_4622,N_4438,N_4429);
and U4623 (N_4623,N_4406,N_4401);
nor U4624 (N_4624,N_4455,N_4479);
and U4625 (N_4625,N_4524,N_4587);
or U4626 (N_4626,N_4592,N_4511);
or U4627 (N_4627,N_4606,N_4500);
nand U4628 (N_4628,N_4600,N_4528);
nand U4629 (N_4629,N_4540,N_4620);
nor U4630 (N_4630,N_4605,N_4516);
and U4631 (N_4631,N_4589,N_4530);
or U4632 (N_4632,N_4607,N_4536);
xor U4633 (N_4633,N_4556,N_4577);
nand U4634 (N_4634,N_4543,N_4538);
nor U4635 (N_4635,N_4507,N_4534);
xnor U4636 (N_4636,N_4501,N_4603);
xor U4637 (N_4637,N_4504,N_4551);
xnor U4638 (N_4638,N_4619,N_4555);
nor U4639 (N_4639,N_4623,N_4505);
and U4640 (N_4640,N_4513,N_4586);
nand U4641 (N_4641,N_4596,N_4562);
nand U4642 (N_4642,N_4618,N_4613);
xnor U4643 (N_4643,N_4510,N_4579);
xnor U4644 (N_4644,N_4584,N_4594);
nand U4645 (N_4645,N_4573,N_4550);
and U4646 (N_4646,N_4535,N_4576);
and U4647 (N_4647,N_4595,N_4611);
nand U4648 (N_4648,N_4546,N_4610);
nand U4649 (N_4649,N_4544,N_4598);
and U4650 (N_4650,N_4580,N_4624);
or U4651 (N_4651,N_4585,N_4614);
xnor U4652 (N_4652,N_4566,N_4557);
and U4653 (N_4653,N_4569,N_4529);
or U4654 (N_4654,N_4616,N_4515);
nand U4655 (N_4655,N_4572,N_4582);
nor U4656 (N_4656,N_4599,N_4602);
or U4657 (N_4657,N_4519,N_4593);
xnor U4658 (N_4658,N_4553,N_4574);
nor U4659 (N_4659,N_4612,N_4548);
xnor U4660 (N_4660,N_4527,N_4571);
xor U4661 (N_4661,N_4597,N_4552);
or U4662 (N_4662,N_4526,N_4564);
nor U4663 (N_4663,N_4517,N_4575);
and U4664 (N_4664,N_4502,N_4617);
and U4665 (N_4665,N_4549,N_4523);
and U4666 (N_4666,N_4525,N_4522);
or U4667 (N_4667,N_4512,N_4558);
xor U4668 (N_4668,N_4508,N_4621);
nand U4669 (N_4669,N_4531,N_4590);
or U4670 (N_4670,N_4608,N_4588);
nand U4671 (N_4671,N_4578,N_4503);
xnor U4672 (N_4672,N_4609,N_4570);
and U4673 (N_4673,N_4583,N_4622);
or U4674 (N_4674,N_4604,N_4521);
nand U4675 (N_4675,N_4518,N_4509);
nand U4676 (N_4676,N_4560,N_4532);
nand U4677 (N_4677,N_4591,N_4568);
or U4678 (N_4678,N_4601,N_4561);
or U4679 (N_4679,N_4542,N_4567);
or U4680 (N_4680,N_4537,N_4514);
nand U4681 (N_4681,N_4506,N_4547);
nand U4682 (N_4682,N_4615,N_4533);
and U4683 (N_4683,N_4520,N_4545);
nor U4684 (N_4684,N_4563,N_4554);
or U4685 (N_4685,N_4559,N_4581);
nand U4686 (N_4686,N_4541,N_4565);
nand U4687 (N_4687,N_4539,N_4575);
and U4688 (N_4688,N_4580,N_4566);
xnor U4689 (N_4689,N_4506,N_4586);
xnor U4690 (N_4690,N_4506,N_4613);
nor U4691 (N_4691,N_4563,N_4559);
and U4692 (N_4692,N_4542,N_4535);
nand U4693 (N_4693,N_4542,N_4526);
or U4694 (N_4694,N_4571,N_4532);
and U4695 (N_4695,N_4572,N_4532);
or U4696 (N_4696,N_4623,N_4502);
nand U4697 (N_4697,N_4510,N_4596);
or U4698 (N_4698,N_4513,N_4545);
xnor U4699 (N_4699,N_4560,N_4591);
nor U4700 (N_4700,N_4576,N_4578);
and U4701 (N_4701,N_4563,N_4604);
nor U4702 (N_4702,N_4563,N_4607);
nor U4703 (N_4703,N_4573,N_4583);
and U4704 (N_4704,N_4514,N_4588);
xor U4705 (N_4705,N_4577,N_4620);
nor U4706 (N_4706,N_4579,N_4541);
and U4707 (N_4707,N_4609,N_4512);
nand U4708 (N_4708,N_4609,N_4574);
xor U4709 (N_4709,N_4579,N_4531);
or U4710 (N_4710,N_4617,N_4528);
xnor U4711 (N_4711,N_4569,N_4542);
or U4712 (N_4712,N_4558,N_4510);
xnor U4713 (N_4713,N_4585,N_4526);
and U4714 (N_4714,N_4589,N_4564);
or U4715 (N_4715,N_4579,N_4524);
nor U4716 (N_4716,N_4613,N_4581);
and U4717 (N_4717,N_4528,N_4548);
xor U4718 (N_4718,N_4507,N_4585);
nand U4719 (N_4719,N_4516,N_4531);
nor U4720 (N_4720,N_4537,N_4569);
and U4721 (N_4721,N_4544,N_4600);
and U4722 (N_4722,N_4622,N_4502);
and U4723 (N_4723,N_4586,N_4609);
xor U4724 (N_4724,N_4620,N_4621);
xor U4725 (N_4725,N_4508,N_4610);
and U4726 (N_4726,N_4592,N_4555);
xor U4727 (N_4727,N_4574,N_4517);
or U4728 (N_4728,N_4568,N_4596);
xnor U4729 (N_4729,N_4611,N_4524);
nand U4730 (N_4730,N_4621,N_4539);
nand U4731 (N_4731,N_4554,N_4574);
nand U4732 (N_4732,N_4518,N_4577);
and U4733 (N_4733,N_4543,N_4623);
or U4734 (N_4734,N_4519,N_4568);
nand U4735 (N_4735,N_4572,N_4620);
xnor U4736 (N_4736,N_4587,N_4566);
or U4737 (N_4737,N_4541,N_4532);
xnor U4738 (N_4738,N_4561,N_4546);
xor U4739 (N_4739,N_4580,N_4593);
nor U4740 (N_4740,N_4516,N_4595);
nor U4741 (N_4741,N_4540,N_4506);
nand U4742 (N_4742,N_4560,N_4564);
nor U4743 (N_4743,N_4612,N_4559);
nor U4744 (N_4744,N_4589,N_4621);
nand U4745 (N_4745,N_4603,N_4560);
nand U4746 (N_4746,N_4547,N_4559);
nand U4747 (N_4747,N_4593,N_4535);
or U4748 (N_4748,N_4624,N_4575);
nand U4749 (N_4749,N_4534,N_4565);
nand U4750 (N_4750,N_4643,N_4703);
xor U4751 (N_4751,N_4656,N_4692);
or U4752 (N_4752,N_4671,N_4710);
xnor U4753 (N_4753,N_4749,N_4704);
nand U4754 (N_4754,N_4740,N_4743);
nor U4755 (N_4755,N_4636,N_4744);
nand U4756 (N_4756,N_4661,N_4732);
or U4757 (N_4757,N_4719,N_4684);
nor U4758 (N_4758,N_4697,N_4728);
or U4759 (N_4759,N_4736,N_4628);
nor U4760 (N_4760,N_4723,N_4714);
or U4761 (N_4761,N_4668,N_4646);
nand U4762 (N_4762,N_4735,N_4669);
or U4763 (N_4763,N_4725,N_4709);
xor U4764 (N_4764,N_4625,N_4693);
xor U4765 (N_4765,N_4659,N_4678);
or U4766 (N_4766,N_4712,N_4726);
and U4767 (N_4767,N_4653,N_4665);
and U4768 (N_4768,N_4708,N_4663);
nor U4769 (N_4769,N_4730,N_4650);
xnor U4770 (N_4770,N_4655,N_4674);
nor U4771 (N_4771,N_4686,N_4688);
nor U4772 (N_4772,N_4657,N_4672);
or U4773 (N_4773,N_4742,N_4664);
or U4774 (N_4774,N_4734,N_4745);
nor U4775 (N_4775,N_4699,N_4658);
or U4776 (N_4776,N_4651,N_4748);
nor U4777 (N_4777,N_4694,N_4685);
xnor U4778 (N_4778,N_4731,N_4629);
or U4779 (N_4779,N_4687,N_4702);
or U4780 (N_4780,N_4626,N_4707);
or U4781 (N_4781,N_4641,N_4737);
xnor U4782 (N_4782,N_4640,N_4683);
nand U4783 (N_4783,N_4738,N_4635);
nand U4784 (N_4784,N_4638,N_4670);
nand U4785 (N_4785,N_4724,N_4673);
xnor U4786 (N_4786,N_4729,N_4682);
nor U4787 (N_4787,N_4741,N_4713);
nor U4788 (N_4788,N_4667,N_4679);
nor U4789 (N_4789,N_4689,N_4716);
nand U4790 (N_4790,N_4700,N_4698);
or U4791 (N_4791,N_4662,N_4633);
and U4792 (N_4792,N_4715,N_4747);
or U4793 (N_4793,N_4642,N_4739);
nand U4794 (N_4794,N_4660,N_4634);
or U4795 (N_4795,N_4705,N_4675);
and U4796 (N_4796,N_4639,N_4644);
and U4797 (N_4797,N_4632,N_4637);
xor U4798 (N_4798,N_4720,N_4721);
xnor U4799 (N_4799,N_4630,N_4649);
and U4800 (N_4800,N_4722,N_4718);
or U4801 (N_4801,N_4648,N_4652);
nor U4802 (N_4802,N_4647,N_4676);
nand U4803 (N_4803,N_4711,N_4696);
nor U4804 (N_4804,N_4717,N_4680);
or U4805 (N_4805,N_4691,N_4677);
xnor U4806 (N_4806,N_4681,N_4746);
xor U4807 (N_4807,N_4666,N_4701);
and U4808 (N_4808,N_4706,N_4627);
or U4809 (N_4809,N_4695,N_4654);
or U4810 (N_4810,N_4727,N_4733);
nand U4811 (N_4811,N_4631,N_4645);
or U4812 (N_4812,N_4690,N_4625);
xor U4813 (N_4813,N_4733,N_4626);
nand U4814 (N_4814,N_4739,N_4658);
nor U4815 (N_4815,N_4686,N_4726);
or U4816 (N_4816,N_4697,N_4628);
nor U4817 (N_4817,N_4741,N_4629);
and U4818 (N_4818,N_4709,N_4707);
xor U4819 (N_4819,N_4734,N_4650);
nor U4820 (N_4820,N_4670,N_4651);
nand U4821 (N_4821,N_4643,N_4641);
and U4822 (N_4822,N_4632,N_4702);
xnor U4823 (N_4823,N_4663,N_4714);
xor U4824 (N_4824,N_4710,N_4708);
and U4825 (N_4825,N_4680,N_4684);
nor U4826 (N_4826,N_4708,N_4694);
and U4827 (N_4827,N_4710,N_4676);
or U4828 (N_4828,N_4700,N_4669);
or U4829 (N_4829,N_4628,N_4641);
and U4830 (N_4830,N_4646,N_4706);
nor U4831 (N_4831,N_4697,N_4690);
nor U4832 (N_4832,N_4683,N_4625);
and U4833 (N_4833,N_4631,N_4691);
and U4834 (N_4834,N_4681,N_4715);
and U4835 (N_4835,N_4714,N_4641);
xnor U4836 (N_4836,N_4627,N_4722);
nor U4837 (N_4837,N_4666,N_4737);
and U4838 (N_4838,N_4652,N_4663);
xor U4839 (N_4839,N_4724,N_4693);
xnor U4840 (N_4840,N_4724,N_4732);
nand U4841 (N_4841,N_4724,N_4648);
xor U4842 (N_4842,N_4733,N_4655);
or U4843 (N_4843,N_4672,N_4644);
and U4844 (N_4844,N_4742,N_4727);
nor U4845 (N_4845,N_4685,N_4731);
nor U4846 (N_4846,N_4688,N_4721);
nand U4847 (N_4847,N_4713,N_4710);
nor U4848 (N_4848,N_4629,N_4745);
or U4849 (N_4849,N_4641,N_4733);
and U4850 (N_4850,N_4669,N_4741);
or U4851 (N_4851,N_4707,N_4685);
nand U4852 (N_4852,N_4637,N_4716);
xor U4853 (N_4853,N_4669,N_4724);
nand U4854 (N_4854,N_4652,N_4656);
and U4855 (N_4855,N_4729,N_4684);
xor U4856 (N_4856,N_4734,N_4711);
nor U4857 (N_4857,N_4733,N_4734);
nand U4858 (N_4858,N_4646,N_4629);
nand U4859 (N_4859,N_4628,N_4742);
xor U4860 (N_4860,N_4692,N_4672);
xnor U4861 (N_4861,N_4658,N_4735);
or U4862 (N_4862,N_4697,N_4661);
and U4863 (N_4863,N_4701,N_4676);
or U4864 (N_4864,N_4656,N_4702);
xor U4865 (N_4865,N_4739,N_4705);
or U4866 (N_4866,N_4678,N_4632);
and U4867 (N_4867,N_4702,N_4645);
xnor U4868 (N_4868,N_4698,N_4669);
and U4869 (N_4869,N_4626,N_4730);
and U4870 (N_4870,N_4698,N_4655);
and U4871 (N_4871,N_4635,N_4638);
xor U4872 (N_4872,N_4722,N_4675);
or U4873 (N_4873,N_4628,N_4726);
and U4874 (N_4874,N_4656,N_4739);
xnor U4875 (N_4875,N_4817,N_4821);
nand U4876 (N_4876,N_4856,N_4837);
nand U4877 (N_4877,N_4829,N_4780);
and U4878 (N_4878,N_4771,N_4756);
and U4879 (N_4879,N_4870,N_4792);
or U4880 (N_4880,N_4782,N_4861);
and U4881 (N_4881,N_4820,N_4860);
and U4882 (N_4882,N_4774,N_4770);
nand U4883 (N_4883,N_4847,N_4849);
nand U4884 (N_4884,N_4810,N_4834);
nand U4885 (N_4885,N_4794,N_4825);
xor U4886 (N_4886,N_4819,N_4853);
xnor U4887 (N_4887,N_4844,N_4822);
nor U4888 (N_4888,N_4790,N_4783);
or U4889 (N_4889,N_4768,N_4809);
and U4890 (N_4890,N_4838,N_4807);
xor U4891 (N_4891,N_4773,N_4785);
xor U4892 (N_4892,N_4826,N_4754);
xor U4893 (N_4893,N_4850,N_4799);
nand U4894 (N_4894,N_4784,N_4873);
nand U4895 (N_4895,N_4872,N_4801);
xor U4896 (N_4896,N_4839,N_4833);
and U4897 (N_4897,N_4786,N_4851);
nand U4898 (N_4898,N_4812,N_4811);
nor U4899 (N_4899,N_4775,N_4805);
or U4900 (N_4900,N_4866,N_4797);
or U4901 (N_4901,N_4778,N_4869);
xor U4902 (N_4902,N_4759,N_4793);
nor U4903 (N_4903,N_4832,N_4823);
or U4904 (N_4904,N_4846,N_4766);
nor U4905 (N_4905,N_4798,N_4816);
nor U4906 (N_4906,N_4765,N_4802);
and U4907 (N_4907,N_4867,N_4814);
nand U4908 (N_4908,N_4777,N_4843);
nand U4909 (N_4909,N_4761,N_4800);
xnor U4910 (N_4910,N_4827,N_4772);
or U4911 (N_4911,N_4831,N_4767);
nand U4912 (N_4912,N_4762,N_4840);
or U4913 (N_4913,N_4789,N_4874);
nand U4914 (N_4914,N_4845,N_4760);
xor U4915 (N_4915,N_4818,N_4764);
xor U4916 (N_4916,N_4864,N_4852);
or U4917 (N_4917,N_4871,N_4758);
nor U4918 (N_4918,N_4858,N_4779);
and U4919 (N_4919,N_4755,N_4828);
and U4920 (N_4920,N_4803,N_4841);
nor U4921 (N_4921,N_4859,N_4751);
and U4922 (N_4922,N_4808,N_4842);
or U4923 (N_4923,N_4788,N_4787);
nor U4924 (N_4924,N_4815,N_4855);
nand U4925 (N_4925,N_4796,N_4824);
and U4926 (N_4926,N_4750,N_4813);
or U4927 (N_4927,N_4857,N_4868);
nand U4928 (N_4928,N_4769,N_4781);
nand U4929 (N_4929,N_4753,N_4752);
and U4930 (N_4930,N_4862,N_4776);
nand U4931 (N_4931,N_4830,N_4863);
or U4932 (N_4932,N_4791,N_4806);
nand U4933 (N_4933,N_4836,N_4795);
xor U4934 (N_4934,N_4763,N_4848);
nor U4935 (N_4935,N_4854,N_4804);
nand U4936 (N_4936,N_4757,N_4865);
and U4937 (N_4937,N_4835,N_4782);
or U4938 (N_4938,N_4770,N_4871);
and U4939 (N_4939,N_4826,N_4849);
or U4940 (N_4940,N_4874,N_4833);
nor U4941 (N_4941,N_4769,N_4755);
nand U4942 (N_4942,N_4755,N_4779);
and U4943 (N_4943,N_4775,N_4761);
or U4944 (N_4944,N_4796,N_4781);
xor U4945 (N_4945,N_4780,N_4802);
xor U4946 (N_4946,N_4776,N_4820);
and U4947 (N_4947,N_4850,N_4790);
nor U4948 (N_4948,N_4819,N_4813);
nand U4949 (N_4949,N_4866,N_4824);
nand U4950 (N_4950,N_4857,N_4760);
xor U4951 (N_4951,N_4781,N_4767);
and U4952 (N_4952,N_4849,N_4832);
xor U4953 (N_4953,N_4829,N_4755);
and U4954 (N_4954,N_4802,N_4856);
or U4955 (N_4955,N_4846,N_4809);
xor U4956 (N_4956,N_4844,N_4754);
or U4957 (N_4957,N_4861,N_4855);
nand U4958 (N_4958,N_4753,N_4870);
xnor U4959 (N_4959,N_4772,N_4825);
and U4960 (N_4960,N_4798,N_4764);
xor U4961 (N_4961,N_4758,N_4821);
nor U4962 (N_4962,N_4781,N_4822);
nand U4963 (N_4963,N_4824,N_4810);
nor U4964 (N_4964,N_4823,N_4857);
or U4965 (N_4965,N_4865,N_4842);
nor U4966 (N_4966,N_4863,N_4767);
nand U4967 (N_4967,N_4793,N_4856);
nand U4968 (N_4968,N_4836,N_4780);
nor U4969 (N_4969,N_4765,N_4785);
and U4970 (N_4970,N_4820,N_4792);
and U4971 (N_4971,N_4781,N_4826);
xor U4972 (N_4972,N_4780,N_4806);
and U4973 (N_4973,N_4831,N_4816);
nand U4974 (N_4974,N_4777,N_4852);
nand U4975 (N_4975,N_4871,N_4837);
xor U4976 (N_4976,N_4806,N_4843);
or U4977 (N_4977,N_4869,N_4844);
nand U4978 (N_4978,N_4782,N_4776);
xnor U4979 (N_4979,N_4755,N_4785);
or U4980 (N_4980,N_4841,N_4772);
xnor U4981 (N_4981,N_4791,N_4853);
or U4982 (N_4982,N_4842,N_4834);
xor U4983 (N_4983,N_4790,N_4865);
and U4984 (N_4984,N_4781,N_4762);
or U4985 (N_4985,N_4759,N_4767);
xor U4986 (N_4986,N_4830,N_4793);
or U4987 (N_4987,N_4756,N_4772);
and U4988 (N_4988,N_4787,N_4782);
and U4989 (N_4989,N_4850,N_4874);
and U4990 (N_4990,N_4765,N_4760);
or U4991 (N_4991,N_4842,N_4772);
nor U4992 (N_4992,N_4773,N_4835);
or U4993 (N_4993,N_4853,N_4798);
or U4994 (N_4994,N_4850,N_4766);
or U4995 (N_4995,N_4804,N_4848);
xor U4996 (N_4996,N_4842,N_4826);
xnor U4997 (N_4997,N_4825,N_4828);
and U4998 (N_4998,N_4782,N_4798);
and U4999 (N_4999,N_4827,N_4770);
xnor U5000 (N_5000,N_4947,N_4937);
nand U5001 (N_5001,N_4952,N_4980);
nor U5002 (N_5002,N_4953,N_4907);
and U5003 (N_5003,N_4998,N_4977);
xor U5004 (N_5004,N_4992,N_4920);
nand U5005 (N_5005,N_4964,N_4876);
and U5006 (N_5006,N_4908,N_4889);
and U5007 (N_5007,N_4979,N_4881);
nor U5008 (N_5008,N_4939,N_4912);
or U5009 (N_5009,N_4880,N_4997);
or U5010 (N_5010,N_4898,N_4884);
and U5011 (N_5011,N_4970,N_4949);
nor U5012 (N_5012,N_4891,N_4895);
nand U5013 (N_5013,N_4958,N_4990);
xnor U5014 (N_5014,N_4946,N_4951);
xnor U5015 (N_5015,N_4969,N_4906);
nand U5016 (N_5016,N_4961,N_4965);
nand U5017 (N_5017,N_4938,N_4887);
nor U5018 (N_5018,N_4924,N_4972);
or U5019 (N_5019,N_4900,N_4915);
nor U5020 (N_5020,N_4919,N_4968);
nand U5021 (N_5021,N_4918,N_4903);
or U5022 (N_5022,N_4971,N_4982);
nand U5023 (N_5023,N_4933,N_4921);
and U5024 (N_5024,N_4989,N_4996);
nor U5025 (N_5025,N_4974,N_4987);
and U5026 (N_5026,N_4999,N_4883);
xnor U5027 (N_5027,N_4988,N_4892);
nor U5028 (N_5028,N_4983,N_4934);
and U5029 (N_5029,N_4875,N_4911);
nor U5030 (N_5030,N_4950,N_4897);
xnor U5031 (N_5031,N_4986,N_4981);
and U5032 (N_5032,N_4944,N_4967);
or U5033 (N_5033,N_4956,N_4896);
nor U5034 (N_5034,N_4922,N_4917);
nand U5035 (N_5035,N_4886,N_4913);
and U5036 (N_5036,N_4929,N_4995);
nor U5037 (N_5037,N_4901,N_4962);
nand U5038 (N_5038,N_4923,N_4948);
and U5039 (N_5039,N_4878,N_4985);
xnor U5040 (N_5040,N_4941,N_4936);
and U5041 (N_5041,N_4963,N_4973);
and U5042 (N_5042,N_4926,N_4984);
and U5043 (N_5043,N_4902,N_4935);
or U5044 (N_5044,N_4991,N_4888);
and U5045 (N_5045,N_4904,N_4993);
nand U5046 (N_5046,N_4960,N_4882);
nand U5047 (N_5047,N_4975,N_4916);
and U5048 (N_5048,N_4928,N_4931);
nand U5049 (N_5049,N_4905,N_4943);
nor U5050 (N_5050,N_4932,N_4945);
or U5051 (N_5051,N_4910,N_4940);
nand U5052 (N_5052,N_4890,N_4899);
or U5053 (N_5053,N_4927,N_4955);
and U5054 (N_5054,N_4925,N_4966);
nand U5055 (N_5055,N_4976,N_4877);
and U5056 (N_5056,N_4930,N_4909);
xor U5057 (N_5057,N_4885,N_4879);
nand U5058 (N_5058,N_4957,N_4994);
nor U5059 (N_5059,N_4914,N_4978);
or U5060 (N_5060,N_4959,N_4894);
xnor U5061 (N_5061,N_4942,N_4893);
xor U5062 (N_5062,N_4954,N_4965);
nand U5063 (N_5063,N_4984,N_4961);
or U5064 (N_5064,N_4926,N_4906);
or U5065 (N_5065,N_4991,N_4920);
and U5066 (N_5066,N_4926,N_4970);
xnor U5067 (N_5067,N_4930,N_4985);
and U5068 (N_5068,N_4958,N_4984);
nor U5069 (N_5069,N_4982,N_4985);
or U5070 (N_5070,N_4933,N_4890);
and U5071 (N_5071,N_4959,N_4983);
and U5072 (N_5072,N_4950,N_4945);
nor U5073 (N_5073,N_4975,N_4915);
xor U5074 (N_5074,N_4972,N_4880);
nor U5075 (N_5075,N_4899,N_4953);
or U5076 (N_5076,N_4935,N_4962);
xor U5077 (N_5077,N_4981,N_4885);
nor U5078 (N_5078,N_4900,N_4969);
and U5079 (N_5079,N_4999,N_4997);
nor U5080 (N_5080,N_4994,N_4891);
xor U5081 (N_5081,N_4962,N_4970);
nor U5082 (N_5082,N_4879,N_4919);
nand U5083 (N_5083,N_4960,N_4895);
or U5084 (N_5084,N_4918,N_4898);
and U5085 (N_5085,N_4891,N_4981);
nor U5086 (N_5086,N_4915,N_4877);
nand U5087 (N_5087,N_4945,N_4995);
nor U5088 (N_5088,N_4944,N_4929);
nand U5089 (N_5089,N_4973,N_4954);
and U5090 (N_5090,N_4996,N_4965);
and U5091 (N_5091,N_4949,N_4996);
or U5092 (N_5092,N_4976,N_4909);
nand U5093 (N_5093,N_4986,N_4914);
and U5094 (N_5094,N_4977,N_4979);
and U5095 (N_5095,N_4958,N_4893);
nand U5096 (N_5096,N_4875,N_4923);
or U5097 (N_5097,N_4982,N_4968);
and U5098 (N_5098,N_4930,N_4944);
nor U5099 (N_5099,N_4890,N_4889);
and U5100 (N_5100,N_4963,N_4893);
xnor U5101 (N_5101,N_4910,N_4984);
nor U5102 (N_5102,N_4908,N_4947);
and U5103 (N_5103,N_4879,N_4954);
nor U5104 (N_5104,N_4973,N_4904);
xnor U5105 (N_5105,N_4968,N_4912);
or U5106 (N_5106,N_4884,N_4985);
or U5107 (N_5107,N_4937,N_4890);
or U5108 (N_5108,N_4991,N_4876);
nor U5109 (N_5109,N_4917,N_4898);
and U5110 (N_5110,N_4992,N_4917);
or U5111 (N_5111,N_4971,N_4913);
nor U5112 (N_5112,N_4923,N_4980);
and U5113 (N_5113,N_4991,N_4929);
nand U5114 (N_5114,N_4994,N_4977);
or U5115 (N_5115,N_4929,N_4948);
nor U5116 (N_5116,N_4964,N_4884);
nand U5117 (N_5117,N_4881,N_4890);
or U5118 (N_5118,N_4889,N_4952);
and U5119 (N_5119,N_4929,N_4923);
xnor U5120 (N_5120,N_4981,N_4949);
xnor U5121 (N_5121,N_4919,N_4929);
or U5122 (N_5122,N_4979,N_4952);
or U5123 (N_5123,N_4936,N_4875);
xor U5124 (N_5124,N_4994,N_4903);
nor U5125 (N_5125,N_5119,N_5082);
nor U5126 (N_5126,N_5069,N_5017);
nor U5127 (N_5127,N_5073,N_5099);
nand U5128 (N_5128,N_5085,N_5039);
xnor U5129 (N_5129,N_5092,N_5059);
nand U5130 (N_5130,N_5124,N_5031);
nor U5131 (N_5131,N_5117,N_5076);
nand U5132 (N_5132,N_5049,N_5078);
or U5133 (N_5133,N_5120,N_5024);
nand U5134 (N_5134,N_5106,N_5002);
nand U5135 (N_5135,N_5087,N_5079);
nor U5136 (N_5136,N_5003,N_5116);
or U5137 (N_5137,N_5081,N_5103);
or U5138 (N_5138,N_5025,N_5090);
nand U5139 (N_5139,N_5108,N_5072);
nor U5140 (N_5140,N_5027,N_5045);
nor U5141 (N_5141,N_5013,N_5034);
or U5142 (N_5142,N_5061,N_5041);
or U5143 (N_5143,N_5004,N_5015);
xor U5144 (N_5144,N_5068,N_5109);
nor U5145 (N_5145,N_5095,N_5000);
nand U5146 (N_5146,N_5055,N_5032);
and U5147 (N_5147,N_5104,N_5014);
xnor U5148 (N_5148,N_5113,N_5051);
nor U5149 (N_5149,N_5048,N_5084);
nor U5150 (N_5150,N_5042,N_5060);
nand U5151 (N_5151,N_5038,N_5064);
nand U5152 (N_5152,N_5026,N_5007);
xor U5153 (N_5153,N_5052,N_5100);
nand U5154 (N_5154,N_5115,N_5050);
nor U5155 (N_5155,N_5122,N_5035);
nand U5156 (N_5156,N_5029,N_5006);
nor U5157 (N_5157,N_5091,N_5043);
nor U5158 (N_5158,N_5077,N_5118);
xnor U5159 (N_5159,N_5019,N_5012);
or U5160 (N_5160,N_5096,N_5008);
nand U5161 (N_5161,N_5028,N_5018);
and U5162 (N_5162,N_5110,N_5121);
nor U5163 (N_5163,N_5062,N_5075);
nand U5164 (N_5164,N_5046,N_5023);
nand U5165 (N_5165,N_5066,N_5067);
xor U5166 (N_5166,N_5107,N_5093);
nand U5167 (N_5167,N_5047,N_5020);
or U5168 (N_5168,N_5111,N_5083);
or U5169 (N_5169,N_5114,N_5074);
or U5170 (N_5170,N_5030,N_5053);
nand U5171 (N_5171,N_5098,N_5065);
and U5172 (N_5172,N_5102,N_5009);
xor U5173 (N_5173,N_5022,N_5070);
xor U5174 (N_5174,N_5016,N_5057);
and U5175 (N_5175,N_5097,N_5063);
xnor U5176 (N_5176,N_5001,N_5040);
xnor U5177 (N_5177,N_5071,N_5112);
nor U5178 (N_5178,N_5105,N_5089);
nand U5179 (N_5179,N_5054,N_5094);
nor U5180 (N_5180,N_5088,N_5080);
and U5181 (N_5181,N_5058,N_5036);
nor U5182 (N_5182,N_5037,N_5011);
and U5183 (N_5183,N_5101,N_5044);
and U5184 (N_5184,N_5123,N_5086);
and U5185 (N_5185,N_5056,N_5021);
xnor U5186 (N_5186,N_5033,N_5010);
nand U5187 (N_5187,N_5005,N_5069);
or U5188 (N_5188,N_5124,N_5079);
or U5189 (N_5189,N_5069,N_5049);
nand U5190 (N_5190,N_5043,N_5103);
and U5191 (N_5191,N_5037,N_5052);
nand U5192 (N_5192,N_5086,N_5124);
or U5193 (N_5193,N_5094,N_5073);
nor U5194 (N_5194,N_5111,N_5084);
nand U5195 (N_5195,N_5091,N_5016);
nor U5196 (N_5196,N_5071,N_5109);
nor U5197 (N_5197,N_5120,N_5061);
nor U5198 (N_5198,N_5071,N_5088);
and U5199 (N_5199,N_5118,N_5004);
xnor U5200 (N_5200,N_5053,N_5120);
or U5201 (N_5201,N_5023,N_5039);
nand U5202 (N_5202,N_5003,N_5002);
nor U5203 (N_5203,N_5117,N_5124);
nor U5204 (N_5204,N_5082,N_5123);
xor U5205 (N_5205,N_5108,N_5092);
xor U5206 (N_5206,N_5090,N_5067);
nand U5207 (N_5207,N_5116,N_5123);
nand U5208 (N_5208,N_5119,N_5039);
and U5209 (N_5209,N_5071,N_5084);
xnor U5210 (N_5210,N_5028,N_5049);
or U5211 (N_5211,N_5075,N_5096);
nand U5212 (N_5212,N_5115,N_5022);
and U5213 (N_5213,N_5016,N_5105);
nor U5214 (N_5214,N_5010,N_5050);
or U5215 (N_5215,N_5075,N_5103);
xnor U5216 (N_5216,N_5034,N_5011);
nand U5217 (N_5217,N_5099,N_5023);
nand U5218 (N_5218,N_5034,N_5091);
or U5219 (N_5219,N_5021,N_5054);
xor U5220 (N_5220,N_5008,N_5124);
nand U5221 (N_5221,N_5083,N_5033);
xor U5222 (N_5222,N_5028,N_5047);
nor U5223 (N_5223,N_5008,N_5077);
and U5224 (N_5224,N_5075,N_5025);
xor U5225 (N_5225,N_5100,N_5024);
or U5226 (N_5226,N_5098,N_5107);
nand U5227 (N_5227,N_5018,N_5007);
nand U5228 (N_5228,N_5080,N_5084);
nand U5229 (N_5229,N_5063,N_5111);
nand U5230 (N_5230,N_5010,N_5043);
or U5231 (N_5231,N_5031,N_5082);
xor U5232 (N_5232,N_5067,N_5044);
nand U5233 (N_5233,N_5038,N_5117);
and U5234 (N_5234,N_5073,N_5019);
nand U5235 (N_5235,N_5024,N_5085);
nand U5236 (N_5236,N_5102,N_5028);
xor U5237 (N_5237,N_5010,N_5040);
nor U5238 (N_5238,N_5009,N_5063);
or U5239 (N_5239,N_5027,N_5024);
or U5240 (N_5240,N_5059,N_5084);
xnor U5241 (N_5241,N_5040,N_5017);
xnor U5242 (N_5242,N_5037,N_5061);
xnor U5243 (N_5243,N_5040,N_5111);
or U5244 (N_5244,N_5023,N_5016);
nor U5245 (N_5245,N_5091,N_5056);
and U5246 (N_5246,N_5078,N_5080);
and U5247 (N_5247,N_5035,N_5069);
and U5248 (N_5248,N_5079,N_5095);
or U5249 (N_5249,N_5008,N_5081);
and U5250 (N_5250,N_5149,N_5198);
and U5251 (N_5251,N_5216,N_5234);
nor U5252 (N_5252,N_5189,N_5184);
nor U5253 (N_5253,N_5241,N_5225);
and U5254 (N_5254,N_5223,N_5132);
nor U5255 (N_5255,N_5230,N_5148);
or U5256 (N_5256,N_5194,N_5145);
nor U5257 (N_5257,N_5219,N_5221);
or U5258 (N_5258,N_5209,N_5138);
xnor U5259 (N_5259,N_5128,N_5125);
and U5260 (N_5260,N_5229,N_5146);
xnor U5261 (N_5261,N_5188,N_5226);
and U5262 (N_5262,N_5178,N_5203);
or U5263 (N_5263,N_5152,N_5180);
or U5264 (N_5264,N_5215,N_5175);
nor U5265 (N_5265,N_5205,N_5161);
nand U5266 (N_5266,N_5160,N_5153);
or U5267 (N_5267,N_5185,N_5164);
or U5268 (N_5268,N_5135,N_5163);
nand U5269 (N_5269,N_5247,N_5237);
and U5270 (N_5270,N_5239,N_5240);
xor U5271 (N_5271,N_5143,N_5244);
xnor U5272 (N_5272,N_5157,N_5150);
and U5273 (N_5273,N_5134,N_5151);
nand U5274 (N_5274,N_5192,N_5212);
nand U5275 (N_5275,N_5182,N_5191);
xor U5276 (N_5276,N_5156,N_5139);
or U5277 (N_5277,N_5169,N_5224);
and U5278 (N_5278,N_5245,N_5144);
and U5279 (N_5279,N_5187,N_5155);
xor U5280 (N_5280,N_5222,N_5211);
and U5281 (N_5281,N_5142,N_5243);
and U5282 (N_5282,N_5217,N_5246);
nor U5283 (N_5283,N_5210,N_5158);
and U5284 (N_5284,N_5173,N_5201);
xnor U5285 (N_5285,N_5186,N_5159);
or U5286 (N_5286,N_5147,N_5227);
and U5287 (N_5287,N_5214,N_5220);
nand U5288 (N_5288,N_5193,N_5181);
and U5289 (N_5289,N_5238,N_5232);
nand U5290 (N_5290,N_5174,N_5202);
and U5291 (N_5291,N_5249,N_5200);
and U5292 (N_5292,N_5197,N_5213);
nor U5293 (N_5293,N_5129,N_5141);
nor U5294 (N_5294,N_5130,N_5167);
nor U5295 (N_5295,N_5154,N_5140);
nand U5296 (N_5296,N_5190,N_5176);
nand U5297 (N_5297,N_5204,N_5228);
nor U5298 (N_5298,N_5126,N_5171);
xnor U5299 (N_5299,N_5137,N_5207);
nor U5300 (N_5300,N_5165,N_5248);
or U5301 (N_5301,N_5218,N_5166);
xor U5302 (N_5302,N_5235,N_5179);
nand U5303 (N_5303,N_5136,N_5133);
and U5304 (N_5304,N_5236,N_5231);
and U5305 (N_5305,N_5199,N_5127);
nor U5306 (N_5306,N_5177,N_5233);
nand U5307 (N_5307,N_5183,N_5196);
xnor U5308 (N_5308,N_5172,N_5206);
nand U5309 (N_5309,N_5242,N_5195);
xnor U5310 (N_5310,N_5168,N_5170);
or U5311 (N_5311,N_5162,N_5131);
nor U5312 (N_5312,N_5208,N_5143);
and U5313 (N_5313,N_5142,N_5248);
nand U5314 (N_5314,N_5207,N_5206);
and U5315 (N_5315,N_5137,N_5214);
or U5316 (N_5316,N_5152,N_5217);
and U5317 (N_5317,N_5185,N_5203);
xnor U5318 (N_5318,N_5189,N_5154);
and U5319 (N_5319,N_5178,N_5196);
nand U5320 (N_5320,N_5182,N_5134);
nand U5321 (N_5321,N_5230,N_5195);
xor U5322 (N_5322,N_5161,N_5158);
or U5323 (N_5323,N_5165,N_5238);
and U5324 (N_5324,N_5207,N_5243);
nor U5325 (N_5325,N_5202,N_5240);
xor U5326 (N_5326,N_5232,N_5192);
and U5327 (N_5327,N_5211,N_5249);
nor U5328 (N_5328,N_5157,N_5197);
and U5329 (N_5329,N_5206,N_5132);
xnor U5330 (N_5330,N_5249,N_5236);
nor U5331 (N_5331,N_5228,N_5208);
or U5332 (N_5332,N_5215,N_5160);
or U5333 (N_5333,N_5232,N_5243);
nor U5334 (N_5334,N_5247,N_5129);
or U5335 (N_5335,N_5167,N_5157);
or U5336 (N_5336,N_5219,N_5237);
or U5337 (N_5337,N_5189,N_5168);
nor U5338 (N_5338,N_5137,N_5179);
nand U5339 (N_5339,N_5193,N_5178);
xor U5340 (N_5340,N_5135,N_5159);
xor U5341 (N_5341,N_5200,N_5230);
xnor U5342 (N_5342,N_5211,N_5201);
and U5343 (N_5343,N_5145,N_5170);
xor U5344 (N_5344,N_5155,N_5134);
or U5345 (N_5345,N_5236,N_5196);
xor U5346 (N_5346,N_5243,N_5189);
xor U5347 (N_5347,N_5131,N_5138);
nor U5348 (N_5348,N_5238,N_5146);
nand U5349 (N_5349,N_5221,N_5189);
nand U5350 (N_5350,N_5162,N_5235);
and U5351 (N_5351,N_5147,N_5169);
nor U5352 (N_5352,N_5224,N_5179);
xnor U5353 (N_5353,N_5137,N_5203);
or U5354 (N_5354,N_5211,N_5183);
and U5355 (N_5355,N_5173,N_5234);
nor U5356 (N_5356,N_5135,N_5205);
and U5357 (N_5357,N_5241,N_5197);
and U5358 (N_5358,N_5215,N_5189);
xor U5359 (N_5359,N_5151,N_5164);
and U5360 (N_5360,N_5190,N_5214);
nand U5361 (N_5361,N_5147,N_5217);
or U5362 (N_5362,N_5230,N_5170);
and U5363 (N_5363,N_5170,N_5220);
nor U5364 (N_5364,N_5193,N_5219);
or U5365 (N_5365,N_5234,N_5129);
and U5366 (N_5366,N_5246,N_5197);
nand U5367 (N_5367,N_5188,N_5241);
nor U5368 (N_5368,N_5183,N_5159);
or U5369 (N_5369,N_5155,N_5126);
nand U5370 (N_5370,N_5125,N_5127);
nor U5371 (N_5371,N_5235,N_5198);
nor U5372 (N_5372,N_5198,N_5174);
xnor U5373 (N_5373,N_5195,N_5149);
nand U5374 (N_5374,N_5195,N_5218);
or U5375 (N_5375,N_5354,N_5261);
and U5376 (N_5376,N_5262,N_5296);
or U5377 (N_5377,N_5293,N_5374);
nand U5378 (N_5378,N_5312,N_5360);
xnor U5379 (N_5379,N_5325,N_5358);
xnor U5380 (N_5380,N_5253,N_5306);
and U5381 (N_5381,N_5259,N_5353);
xor U5382 (N_5382,N_5352,N_5319);
xnor U5383 (N_5383,N_5349,N_5322);
nor U5384 (N_5384,N_5300,N_5287);
or U5385 (N_5385,N_5301,N_5336);
or U5386 (N_5386,N_5339,N_5264);
or U5387 (N_5387,N_5343,N_5272);
or U5388 (N_5388,N_5307,N_5334);
or U5389 (N_5389,N_5278,N_5303);
nand U5390 (N_5390,N_5346,N_5368);
xnor U5391 (N_5391,N_5252,N_5328);
and U5392 (N_5392,N_5276,N_5320);
and U5393 (N_5393,N_5270,N_5292);
or U5394 (N_5394,N_5317,N_5370);
xnor U5395 (N_5395,N_5348,N_5310);
or U5396 (N_5396,N_5337,N_5281);
xnor U5397 (N_5397,N_5260,N_5356);
nand U5398 (N_5398,N_5341,N_5308);
nand U5399 (N_5399,N_5316,N_5265);
xnor U5400 (N_5400,N_5280,N_5297);
nand U5401 (N_5401,N_5267,N_5277);
and U5402 (N_5402,N_5362,N_5299);
nand U5403 (N_5403,N_5290,N_5350);
nand U5404 (N_5404,N_5324,N_5351);
xor U5405 (N_5405,N_5372,N_5295);
or U5406 (N_5406,N_5283,N_5286);
nor U5407 (N_5407,N_5279,N_5314);
and U5408 (N_5408,N_5340,N_5327);
nor U5409 (N_5409,N_5332,N_5367);
xnor U5410 (N_5410,N_5284,N_5373);
nor U5411 (N_5411,N_5357,N_5335);
nor U5412 (N_5412,N_5369,N_5347);
xor U5413 (N_5413,N_5338,N_5344);
xor U5414 (N_5414,N_5269,N_5321);
or U5415 (N_5415,N_5304,N_5254);
and U5416 (N_5416,N_5288,N_5363);
nand U5417 (N_5417,N_5326,N_5291);
xnor U5418 (N_5418,N_5282,N_5361);
xnor U5419 (N_5419,N_5266,N_5313);
and U5420 (N_5420,N_5355,N_5323);
xnor U5421 (N_5421,N_5256,N_5263);
nand U5422 (N_5422,N_5255,N_5302);
nand U5423 (N_5423,N_5364,N_5371);
or U5424 (N_5424,N_5298,N_5274);
xnor U5425 (N_5425,N_5331,N_5366);
nand U5426 (N_5426,N_5289,N_5329);
nand U5427 (N_5427,N_5251,N_5268);
xnor U5428 (N_5428,N_5311,N_5333);
nor U5429 (N_5429,N_5342,N_5273);
and U5430 (N_5430,N_5365,N_5318);
or U5431 (N_5431,N_5257,N_5315);
nor U5432 (N_5432,N_5294,N_5345);
nand U5433 (N_5433,N_5258,N_5275);
nand U5434 (N_5434,N_5359,N_5330);
and U5435 (N_5435,N_5309,N_5305);
and U5436 (N_5436,N_5271,N_5250);
or U5437 (N_5437,N_5285,N_5320);
or U5438 (N_5438,N_5312,N_5329);
xnor U5439 (N_5439,N_5310,N_5364);
nor U5440 (N_5440,N_5268,N_5279);
nand U5441 (N_5441,N_5372,N_5265);
xnor U5442 (N_5442,N_5328,N_5361);
xor U5443 (N_5443,N_5256,N_5286);
nand U5444 (N_5444,N_5304,N_5298);
and U5445 (N_5445,N_5335,N_5255);
and U5446 (N_5446,N_5373,N_5331);
and U5447 (N_5447,N_5260,N_5370);
and U5448 (N_5448,N_5279,N_5257);
or U5449 (N_5449,N_5331,N_5337);
or U5450 (N_5450,N_5260,N_5362);
or U5451 (N_5451,N_5356,N_5364);
or U5452 (N_5452,N_5333,N_5334);
or U5453 (N_5453,N_5285,N_5336);
and U5454 (N_5454,N_5270,N_5312);
nor U5455 (N_5455,N_5283,N_5330);
nor U5456 (N_5456,N_5289,N_5321);
xor U5457 (N_5457,N_5300,N_5257);
nor U5458 (N_5458,N_5250,N_5269);
nor U5459 (N_5459,N_5356,N_5360);
and U5460 (N_5460,N_5296,N_5313);
nand U5461 (N_5461,N_5315,N_5366);
xnor U5462 (N_5462,N_5323,N_5299);
nand U5463 (N_5463,N_5352,N_5349);
xnor U5464 (N_5464,N_5329,N_5324);
or U5465 (N_5465,N_5273,N_5279);
nor U5466 (N_5466,N_5251,N_5264);
or U5467 (N_5467,N_5277,N_5311);
nor U5468 (N_5468,N_5357,N_5344);
and U5469 (N_5469,N_5254,N_5321);
and U5470 (N_5470,N_5300,N_5295);
nor U5471 (N_5471,N_5275,N_5306);
or U5472 (N_5472,N_5283,N_5293);
nor U5473 (N_5473,N_5270,N_5324);
and U5474 (N_5474,N_5260,N_5296);
and U5475 (N_5475,N_5371,N_5354);
xor U5476 (N_5476,N_5279,N_5344);
nor U5477 (N_5477,N_5339,N_5334);
nand U5478 (N_5478,N_5267,N_5276);
or U5479 (N_5479,N_5322,N_5324);
nand U5480 (N_5480,N_5374,N_5372);
xor U5481 (N_5481,N_5311,N_5357);
nor U5482 (N_5482,N_5262,N_5283);
nand U5483 (N_5483,N_5289,N_5345);
and U5484 (N_5484,N_5362,N_5268);
or U5485 (N_5485,N_5302,N_5252);
nor U5486 (N_5486,N_5350,N_5273);
nor U5487 (N_5487,N_5348,N_5255);
nor U5488 (N_5488,N_5321,N_5263);
xnor U5489 (N_5489,N_5284,N_5274);
or U5490 (N_5490,N_5328,N_5317);
xor U5491 (N_5491,N_5321,N_5331);
nand U5492 (N_5492,N_5329,N_5334);
nor U5493 (N_5493,N_5358,N_5275);
nor U5494 (N_5494,N_5316,N_5354);
nand U5495 (N_5495,N_5257,N_5297);
nor U5496 (N_5496,N_5317,N_5331);
or U5497 (N_5497,N_5340,N_5329);
and U5498 (N_5498,N_5270,N_5302);
and U5499 (N_5499,N_5332,N_5348);
xor U5500 (N_5500,N_5490,N_5381);
xnor U5501 (N_5501,N_5386,N_5488);
nand U5502 (N_5502,N_5426,N_5387);
nand U5503 (N_5503,N_5458,N_5440);
or U5504 (N_5504,N_5457,N_5473);
xor U5505 (N_5505,N_5447,N_5431);
nor U5506 (N_5506,N_5491,N_5406);
nand U5507 (N_5507,N_5434,N_5429);
xnor U5508 (N_5508,N_5449,N_5463);
xor U5509 (N_5509,N_5393,N_5446);
nor U5510 (N_5510,N_5489,N_5414);
nor U5511 (N_5511,N_5476,N_5401);
and U5512 (N_5512,N_5478,N_5481);
or U5513 (N_5513,N_5445,N_5485);
nor U5514 (N_5514,N_5487,N_5405);
or U5515 (N_5515,N_5479,N_5437);
nand U5516 (N_5516,N_5462,N_5395);
and U5517 (N_5517,N_5496,N_5411);
and U5518 (N_5518,N_5400,N_5483);
or U5519 (N_5519,N_5442,N_5424);
and U5520 (N_5520,N_5408,N_5389);
nand U5521 (N_5521,N_5492,N_5441);
and U5522 (N_5522,N_5435,N_5422);
or U5523 (N_5523,N_5376,N_5409);
nor U5524 (N_5524,N_5474,N_5417);
nand U5525 (N_5525,N_5421,N_5456);
nor U5526 (N_5526,N_5425,N_5494);
xnor U5527 (N_5527,N_5391,N_5423);
xor U5528 (N_5528,N_5392,N_5377);
nor U5529 (N_5529,N_5420,N_5498);
or U5530 (N_5530,N_5453,N_5428);
nand U5531 (N_5531,N_5378,N_5499);
xor U5532 (N_5532,N_5385,N_5404);
or U5533 (N_5533,N_5495,N_5465);
and U5534 (N_5534,N_5486,N_5444);
nor U5535 (N_5535,N_5477,N_5375);
xnor U5536 (N_5536,N_5451,N_5455);
nand U5537 (N_5537,N_5390,N_5493);
and U5538 (N_5538,N_5472,N_5410);
xor U5539 (N_5539,N_5397,N_5475);
or U5540 (N_5540,N_5433,N_5379);
and U5541 (N_5541,N_5454,N_5484);
and U5542 (N_5542,N_5467,N_5402);
nor U5543 (N_5543,N_5443,N_5469);
nand U5544 (N_5544,N_5461,N_5407);
xor U5545 (N_5545,N_5438,N_5383);
nor U5546 (N_5546,N_5482,N_5430);
and U5547 (N_5547,N_5418,N_5480);
or U5548 (N_5548,N_5470,N_5403);
and U5549 (N_5549,N_5466,N_5415);
nand U5550 (N_5550,N_5448,N_5460);
and U5551 (N_5551,N_5399,N_5382);
or U5552 (N_5552,N_5497,N_5380);
nor U5553 (N_5553,N_5388,N_5459);
nor U5554 (N_5554,N_5471,N_5416);
xor U5555 (N_5555,N_5436,N_5396);
and U5556 (N_5556,N_5398,N_5427);
and U5557 (N_5557,N_5464,N_5439);
or U5558 (N_5558,N_5432,N_5452);
xnor U5559 (N_5559,N_5412,N_5450);
and U5560 (N_5560,N_5419,N_5468);
or U5561 (N_5561,N_5384,N_5413);
xor U5562 (N_5562,N_5394,N_5401);
xor U5563 (N_5563,N_5385,N_5465);
or U5564 (N_5564,N_5422,N_5494);
nand U5565 (N_5565,N_5498,N_5494);
nand U5566 (N_5566,N_5475,N_5411);
nand U5567 (N_5567,N_5406,N_5449);
or U5568 (N_5568,N_5427,N_5381);
or U5569 (N_5569,N_5412,N_5456);
nor U5570 (N_5570,N_5394,N_5443);
and U5571 (N_5571,N_5483,N_5445);
nand U5572 (N_5572,N_5403,N_5389);
xor U5573 (N_5573,N_5424,N_5383);
nand U5574 (N_5574,N_5407,N_5435);
xor U5575 (N_5575,N_5478,N_5433);
and U5576 (N_5576,N_5396,N_5393);
nor U5577 (N_5577,N_5376,N_5399);
nor U5578 (N_5578,N_5430,N_5442);
xor U5579 (N_5579,N_5488,N_5477);
and U5580 (N_5580,N_5420,N_5469);
and U5581 (N_5581,N_5437,N_5495);
and U5582 (N_5582,N_5439,N_5438);
or U5583 (N_5583,N_5451,N_5475);
or U5584 (N_5584,N_5444,N_5457);
and U5585 (N_5585,N_5471,N_5460);
nor U5586 (N_5586,N_5464,N_5393);
and U5587 (N_5587,N_5410,N_5398);
nand U5588 (N_5588,N_5475,N_5464);
xor U5589 (N_5589,N_5471,N_5440);
or U5590 (N_5590,N_5412,N_5499);
nand U5591 (N_5591,N_5496,N_5414);
xor U5592 (N_5592,N_5476,N_5407);
nand U5593 (N_5593,N_5430,N_5441);
xnor U5594 (N_5594,N_5450,N_5376);
or U5595 (N_5595,N_5432,N_5490);
or U5596 (N_5596,N_5391,N_5415);
or U5597 (N_5597,N_5452,N_5424);
xnor U5598 (N_5598,N_5440,N_5479);
and U5599 (N_5599,N_5459,N_5426);
xor U5600 (N_5600,N_5409,N_5429);
xor U5601 (N_5601,N_5440,N_5429);
nand U5602 (N_5602,N_5484,N_5485);
xor U5603 (N_5603,N_5377,N_5402);
nor U5604 (N_5604,N_5412,N_5386);
nand U5605 (N_5605,N_5393,N_5445);
xor U5606 (N_5606,N_5438,N_5440);
and U5607 (N_5607,N_5460,N_5423);
nand U5608 (N_5608,N_5400,N_5441);
or U5609 (N_5609,N_5457,N_5498);
nor U5610 (N_5610,N_5415,N_5419);
nor U5611 (N_5611,N_5378,N_5409);
and U5612 (N_5612,N_5434,N_5460);
and U5613 (N_5613,N_5413,N_5459);
nand U5614 (N_5614,N_5380,N_5469);
nor U5615 (N_5615,N_5417,N_5432);
or U5616 (N_5616,N_5405,N_5387);
or U5617 (N_5617,N_5412,N_5390);
and U5618 (N_5618,N_5432,N_5448);
nand U5619 (N_5619,N_5457,N_5403);
xor U5620 (N_5620,N_5462,N_5494);
or U5621 (N_5621,N_5400,N_5375);
nor U5622 (N_5622,N_5412,N_5483);
or U5623 (N_5623,N_5480,N_5457);
nand U5624 (N_5624,N_5375,N_5426);
nand U5625 (N_5625,N_5573,N_5611);
xnor U5626 (N_5626,N_5571,N_5504);
xor U5627 (N_5627,N_5562,N_5592);
nor U5628 (N_5628,N_5512,N_5520);
or U5629 (N_5629,N_5524,N_5608);
and U5630 (N_5630,N_5583,N_5561);
and U5631 (N_5631,N_5510,N_5614);
nor U5632 (N_5632,N_5556,N_5545);
nor U5633 (N_5633,N_5526,N_5519);
or U5634 (N_5634,N_5601,N_5567);
or U5635 (N_5635,N_5506,N_5516);
xor U5636 (N_5636,N_5600,N_5525);
nor U5637 (N_5637,N_5534,N_5580);
nand U5638 (N_5638,N_5543,N_5550);
xor U5639 (N_5639,N_5589,N_5576);
or U5640 (N_5640,N_5509,N_5542);
nand U5641 (N_5641,N_5521,N_5610);
nor U5642 (N_5642,N_5586,N_5617);
nand U5643 (N_5643,N_5555,N_5574);
or U5644 (N_5644,N_5565,N_5618);
nand U5645 (N_5645,N_5619,N_5500);
xnor U5646 (N_5646,N_5606,N_5532);
or U5647 (N_5647,N_5604,N_5563);
and U5648 (N_5648,N_5541,N_5503);
xnor U5649 (N_5649,N_5622,N_5518);
and U5650 (N_5650,N_5582,N_5568);
xnor U5651 (N_5651,N_5537,N_5514);
nand U5652 (N_5652,N_5505,N_5507);
or U5653 (N_5653,N_5578,N_5624);
or U5654 (N_5654,N_5615,N_5558);
and U5655 (N_5655,N_5591,N_5533);
or U5656 (N_5656,N_5522,N_5515);
or U5657 (N_5657,N_5501,N_5536);
nand U5658 (N_5658,N_5613,N_5584);
or U5659 (N_5659,N_5513,N_5557);
xor U5660 (N_5660,N_5539,N_5595);
nand U5661 (N_5661,N_5548,N_5616);
xnor U5662 (N_5662,N_5588,N_5581);
nand U5663 (N_5663,N_5605,N_5523);
nor U5664 (N_5664,N_5529,N_5547);
xnor U5665 (N_5665,N_5566,N_5502);
nor U5666 (N_5666,N_5593,N_5544);
nand U5667 (N_5667,N_5535,N_5587);
nand U5668 (N_5668,N_5554,N_5607);
nand U5669 (N_5669,N_5572,N_5609);
nand U5670 (N_5670,N_5549,N_5597);
xnor U5671 (N_5671,N_5540,N_5531);
nor U5672 (N_5672,N_5603,N_5594);
nor U5673 (N_5673,N_5538,N_5577);
and U5674 (N_5674,N_5530,N_5585);
and U5675 (N_5675,N_5598,N_5560);
nor U5676 (N_5676,N_5527,N_5612);
and U5677 (N_5677,N_5599,N_5553);
nor U5678 (N_5678,N_5508,N_5623);
nor U5679 (N_5679,N_5596,N_5546);
nor U5680 (N_5680,N_5552,N_5602);
nand U5681 (N_5681,N_5621,N_5579);
and U5682 (N_5682,N_5575,N_5511);
or U5683 (N_5683,N_5620,N_5570);
or U5684 (N_5684,N_5590,N_5551);
or U5685 (N_5685,N_5559,N_5564);
and U5686 (N_5686,N_5517,N_5569);
nand U5687 (N_5687,N_5528,N_5592);
xnor U5688 (N_5688,N_5504,N_5561);
and U5689 (N_5689,N_5510,N_5557);
xnor U5690 (N_5690,N_5539,N_5516);
xnor U5691 (N_5691,N_5601,N_5517);
nor U5692 (N_5692,N_5532,N_5500);
and U5693 (N_5693,N_5519,N_5554);
or U5694 (N_5694,N_5618,N_5602);
or U5695 (N_5695,N_5600,N_5609);
nand U5696 (N_5696,N_5558,N_5515);
nor U5697 (N_5697,N_5582,N_5564);
and U5698 (N_5698,N_5524,N_5624);
and U5699 (N_5699,N_5580,N_5579);
or U5700 (N_5700,N_5545,N_5624);
nor U5701 (N_5701,N_5579,N_5523);
nand U5702 (N_5702,N_5503,N_5597);
and U5703 (N_5703,N_5529,N_5600);
xor U5704 (N_5704,N_5620,N_5610);
xnor U5705 (N_5705,N_5527,N_5570);
or U5706 (N_5706,N_5594,N_5566);
nand U5707 (N_5707,N_5557,N_5535);
xnor U5708 (N_5708,N_5609,N_5516);
and U5709 (N_5709,N_5551,N_5518);
and U5710 (N_5710,N_5613,N_5523);
xor U5711 (N_5711,N_5589,N_5606);
xnor U5712 (N_5712,N_5603,N_5610);
and U5713 (N_5713,N_5500,N_5576);
nor U5714 (N_5714,N_5594,N_5523);
or U5715 (N_5715,N_5580,N_5591);
nand U5716 (N_5716,N_5505,N_5535);
and U5717 (N_5717,N_5609,N_5508);
nor U5718 (N_5718,N_5619,N_5587);
or U5719 (N_5719,N_5604,N_5523);
or U5720 (N_5720,N_5614,N_5616);
nand U5721 (N_5721,N_5535,N_5577);
nand U5722 (N_5722,N_5601,N_5511);
nor U5723 (N_5723,N_5543,N_5520);
xnor U5724 (N_5724,N_5600,N_5515);
nand U5725 (N_5725,N_5604,N_5595);
and U5726 (N_5726,N_5537,N_5510);
and U5727 (N_5727,N_5560,N_5620);
or U5728 (N_5728,N_5509,N_5510);
and U5729 (N_5729,N_5575,N_5544);
nor U5730 (N_5730,N_5549,N_5587);
nor U5731 (N_5731,N_5544,N_5540);
and U5732 (N_5732,N_5619,N_5512);
nand U5733 (N_5733,N_5506,N_5620);
and U5734 (N_5734,N_5563,N_5536);
nor U5735 (N_5735,N_5567,N_5573);
xor U5736 (N_5736,N_5520,N_5506);
and U5737 (N_5737,N_5541,N_5594);
nand U5738 (N_5738,N_5623,N_5504);
xnor U5739 (N_5739,N_5598,N_5520);
or U5740 (N_5740,N_5546,N_5622);
nor U5741 (N_5741,N_5564,N_5589);
xor U5742 (N_5742,N_5517,N_5544);
nand U5743 (N_5743,N_5536,N_5545);
and U5744 (N_5744,N_5609,N_5561);
or U5745 (N_5745,N_5503,N_5548);
and U5746 (N_5746,N_5539,N_5570);
and U5747 (N_5747,N_5532,N_5554);
and U5748 (N_5748,N_5552,N_5609);
xnor U5749 (N_5749,N_5554,N_5528);
and U5750 (N_5750,N_5721,N_5717);
and U5751 (N_5751,N_5642,N_5670);
xnor U5752 (N_5752,N_5737,N_5689);
or U5753 (N_5753,N_5749,N_5703);
and U5754 (N_5754,N_5639,N_5668);
nor U5755 (N_5755,N_5650,N_5630);
or U5756 (N_5756,N_5641,N_5681);
nand U5757 (N_5757,N_5655,N_5740);
nand U5758 (N_5758,N_5708,N_5718);
and U5759 (N_5759,N_5744,N_5648);
xor U5760 (N_5760,N_5663,N_5692);
or U5761 (N_5761,N_5738,N_5646);
and U5762 (N_5762,N_5691,N_5706);
and U5763 (N_5763,N_5686,N_5707);
nand U5764 (N_5764,N_5748,N_5658);
xor U5765 (N_5765,N_5632,N_5698);
and U5766 (N_5766,N_5702,N_5634);
and U5767 (N_5767,N_5637,N_5656);
nor U5768 (N_5768,N_5661,N_5682);
and U5769 (N_5769,N_5726,N_5664);
and U5770 (N_5770,N_5627,N_5690);
xnor U5771 (N_5771,N_5635,N_5651);
and U5772 (N_5772,N_5640,N_5722);
nand U5773 (N_5773,N_5687,N_5665);
or U5774 (N_5774,N_5710,N_5678);
or U5775 (N_5775,N_5649,N_5713);
xor U5776 (N_5776,N_5735,N_5629);
xor U5777 (N_5777,N_5720,N_5747);
xnor U5778 (N_5778,N_5684,N_5643);
xnor U5779 (N_5779,N_5725,N_5679);
nor U5780 (N_5780,N_5662,N_5705);
nor U5781 (N_5781,N_5695,N_5697);
or U5782 (N_5782,N_5647,N_5666);
nor U5783 (N_5783,N_5729,N_5719);
or U5784 (N_5784,N_5714,N_5694);
and U5785 (N_5785,N_5657,N_5626);
nor U5786 (N_5786,N_5716,N_5677);
and U5787 (N_5787,N_5732,N_5715);
xnor U5788 (N_5788,N_5659,N_5709);
and U5789 (N_5789,N_5730,N_5711);
and U5790 (N_5790,N_5733,N_5685);
nor U5791 (N_5791,N_5727,N_5745);
or U5792 (N_5792,N_5746,N_5654);
xor U5793 (N_5793,N_5712,N_5674);
nand U5794 (N_5794,N_5638,N_5636);
nor U5795 (N_5795,N_5704,N_5701);
and U5796 (N_5796,N_5739,N_5743);
and U5797 (N_5797,N_5734,N_5660);
nor U5798 (N_5798,N_5672,N_5723);
xnor U5799 (N_5799,N_5741,N_5653);
nand U5800 (N_5800,N_5645,N_5667);
xnor U5801 (N_5801,N_5696,N_5628);
or U5802 (N_5802,N_5731,N_5675);
and U5803 (N_5803,N_5688,N_5699);
nand U5804 (N_5804,N_5669,N_5673);
nand U5805 (N_5805,N_5631,N_5652);
nand U5806 (N_5806,N_5736,N_5671);
nand U5807 (N_5807,N_5625,N_5700);
and U5808 (N_5808,N_5693,N_5633);
and U5809 (N_5809,N_5680,N_5724);
nand U5810 (N_5810,N_5676,N_5683);
nand U5811 (N_5811,N_5742,N_5728);
or U5812 (N_5812,N_5644,N_5701);
nor U5813 (N_5813,N_5739,N_5663);
or U5814 (N_5814,N_5714,N_5628);
nand U5815 (N_5815,N_5641,N_5638);
nand U5816 (N_5816,N_5648,N_5719);
nand U5817 (N_5817,N_5723,N_5670);
nand U5818 (N_5818,N_5708,N_5691);
xor U5819 (N_5819,N_5672,N_5730);
or U5820 (N_5820,N_5676,N_5748);
and U5821 (N_5821,N_5661,N_5712);
and U5822 (N_5822,N_5661,N_5672);
nand U5823 (N_5823,N_5737,N_5700);
nor U5824 (N_5824,N_5654,N_5644);
or U5825 (N_5825,N_5664,N_5647);
and U5826 (N_5826,N_5709,N_5689);
or U5827 (N_5827,N_5631,N_5720);
nor U5828 (N_5828,N_5640,N_5709);
or U5829 (N_5829,N_5742,N_5731);
nor U5830 (N_5830,N_5690,N_5677);
xor U5831 (N_5831,N_5696,N_5632);
xnor U5832 (N_5832,N_5673,N_5685);
xnor U5833 (N_5833,N_5632,N_5658);
or U5834 (N_5834,N_5678,N_5634);
xnor U5835 (N_5835,N_5749,N_5680);
or U5836 (N_5836,N_5656,N_5683);
nand U5837 (N_5837,N_5626,N_5699);
xnor U5838 (N_5838,N_5643,N_5727);
nand U5839 (N_5839,N_5736,N_5687);
and U5840 (N_5840,N_5634,N_5710);
xnor U5841 (N_5841,N_5687,N_5648);
nand U5842 (N_5842,N_5716,N_5685);
or U5843 (N_5843,N_5721,N_5631);
and U5844 (N_5844,N_5712,N_5642);
or U5845 (N_5845,N_5740,N_5704);
xnor U5846 (N_5846,N_5625,N_5670);
or U5847 (N_5847,N_5708,N_5682);
or U5848 (N_5848,N_5713,N_5671);
or U5849 (N_5849,N_5668,N_5691);
nor U5850 (N_5850,N_5639,N_5749);
and U5851 (N_5851,N_5706,N_5687);
and U5852 (N_5852,N_5723,N_5700);
nand U5853 (N_5853,N_5744,N_5720);
nor U5854 (N_5854,N_5698,N_5699);
xor U5855 (N_5855,N_5626,N_5718);
and U5856 (N_5856,N_5742,N_5672);
and U5857 (N_5857,N_5684,N_5665);
nor U5858 (N_5858,N_5707,N_5628);
nand U5859 (N_5859,N_5734,N_5736);
nand U5860 (N_5860,N_5749,N_5707);
xor U5861 (N_5861,N_5739,N_5661);
and U5862 (N_5862,N_5710,N_5639);
or U5863 (N_5863,N_5698,N_5648);
or U5864 (N_5864,N_5629,N_5676);
or U5865 (N_5865,N_5675,N_5721);
nor U5866 (N_5866,N_5658,N_5670);
xnor U5867 (N_5867,N_5721,N_5723);
or U5868 (N_5868,N_5721,N_5659);
xor U5869 (N_5869,N_5633,N_5659);
or U5870 (N_5870,N_5649,N_5745);
nand U5871 (N_5871,N_5683,N_5734);
and U5872 (N_5872,N_5707,N_5677);
nand U5873 (N_5873,N_5630,N_5669);
xor U5874 (N_5874,N_5743,N_5735);
nand U5875 (N_5875,N_5766,N_5848);
and U5876 (N_5876,N_5820,N_5841);
or U5877 (N_5877,N_5819,N_5829);
or U5878 (N_5878,N_5869,N_5827);
and U5879 (N_5879,N_5795,N_5811);
xor U5880 (N_5880,N_5798,N_5776);
or U5881 (N_5881,N_5810,N_5814);
or U5882 (N_5882,N_5851,N_5769);
or U5883 (N_5883,N_5854,N_5850);
nand U5884 (N_5884,N_5834,N_5754);
and U5885 (N_5885,N_5858,N_5778);
nand U5886 (N_5886,N_5785,N_5764);
and U5887 (N_5887,N_5847,N_5805);
and U5888 (N_5888,N_5797,N_5789);
nor U5889 (N_5889,N_5815,N_5765);
or U5890 (N_5890,N_5832,N_5857);
nand U5891 (N_5891,N_5817,N_5753);
and U5892 (N_5892,N_5781,N_5796);
or U5893 (N_5893,N_5763,N_5853);
xor U5894 (N_5894,N_5783,N_5801);
and U5895 (N_5895,N_5775,N_5831);
nor U5896 (N_5896,N_5755,N_5813);
xnor U5897 (N_5897,N_5821,N_5777);
and U5898 (N_5898,N_5774,N_5788);
and U5899 (N_5899,N_5790,N_5836);
nor U5900 (N_5900,N_5830,N_5823);
xor U5901 (N_5901,N_5800,N_5806);
and U5902 (N_5902,N_5818,N_5852);
nand U5903 (N_5903,N_5861,N_5828);
and U5904 (N_5904,N_5837,N_5843);
nor U5905 (N_5905,N_5825,N_5794);
nand U5906 (N_5906,N_5855,N_5874);
xnor U5907 (N_5907,N_5770,N_5842);
xnor U5908 (N_5908,N_5812,N_5856);
or U5909 (N_5909,N_5863,N_5787);
and U5910 (N_5910,N_5772,N_5784);
xor U5911 (N_5911,N_5791,N_5760);
nor U5912 (N_5912,N_5807,N_5750);
xnor U5913 (N_5913,N_5822,N_5867);
or U5914 (N_5914,N_5779,N_5840);
nor U5915 (N_5915,N_5757,N_5864);
nor U5916 (N_5916,N_5809,N_5799);
and U5917 (N_5917,N_5865,N_5756);
or U5918 (N_5918,N_5816,N_5759);
or U5919 (N_5919,N_5838,N_5803);
nand U5920 (N_5920,N_5792,N_5771);
or U5921 (N_5921,N_5793,N_5786);
or U5922 (N_5922,N_5767,N_5868);
or U5923 (N_5923,N_5873,N_5782);
xnor U5924 (N_5924,N_5768,N_5870);
nor U5925 (N_5925,N_5862,N_5844);
xnor U5926 (N_5926,N_5752,N_5871);
and U5927 (N_5927,N_5802,N_5859);
or U5928 (N_5928,N_5751,N_5804);
nand U5929 (N_5929,N_5846,N_5866);
or U5930 (N_5930,N_5835,N_5758);
and U5931 (N_5931,N_5833,N_5808);
nor U5932 (N_5932,N_5872,N_5762);
or U5933 (N_5933,N_5773,N_5860);
and U5934 (N_5934,N_5849,N_5839);
and U5935 (N_5935,N_5761,N_5826);
nand U5936 (N_5936,N_5845,N_5824);
and U5937 (N_5937,N_5780,N_5790);
nand U5938 (N_5938,N_5823,N_5756);
nor U5939 (N_5939,N_5779,N_5781);
and U5940 (N_5940,N_5783,N_5805);
nor U5941 (N_5941,N_5849,N_5831);
and U5942 (N_5942,N_5870,N_5775);
and U5943 (N_5943,N_5841,N_5848);
or U5944 (N_5944,N_5829,N_5863);
or U5945 (N_5945,N_5866,N_5858);
nor U5946 (N_5946,N_5784,N_5793);
nor U5947 (N_5947,N_5773,N_5857);
and U5948 (N_5948,N_5804,N_5835);
nor U5949 (N_5949,N_5767,N_5760);
nor U5950 (N_5950,N_5808,N_5800);
nor U5951 (N_5951,N_5803,N_5863);
xor U5952 (N_5952,N_5779,N_5860);
xor U5953 (N_5953,N_5863,N_5788);
nor U5954 (N_5954,N_5781,N_5873);
nor U5955 (N_5955,N_5803,N_5801);
nand U5956 (N_5956,N_5849,N_5808);
nand U5957 (N_5957,N_5803,N_5797);
or U5958 (N_5958,N_5872,N_5859);
nor U5959 (N_5959,N_5855,N_5831);
or U5960 (N_5960,N_5823,N_5769);
xnor U5961 (N_5961,N_5769,N_5771);
and U5962 (N_5962,N_5790,N_5852);
nor U5963 (N_5963,N_5759,N_5824);
or U5964 (N_5964,N_5819,N_5806);
xor U5965 (N_5965,N_5856,N_5769);
nor U5966 (N_5966,N_5858,N_5767);
or U5967 (N_5967,N_5774,N_5828);
nor U5968 (N_5968,N_5869,N_5757);
nand U5969 (N_5969,N_5863,N_5759);
and U5970 (N_5970,N_5766,N_5784);
nor U5971 (N_5971,N_5788,N_5853);
nand U5972 (N_5972,N_5753,N_5767);
and U5973 (N_5973,N_5841,N_5831);
nand U5974 (N_5974,N_5845,N_5856);
nand U5975 (N_5975,N_5839,N_5830);
nand U5976 (N_5976,N_5795,N_5813);
nand U5977 (N_5977,N_5787,N_5776);
nand U5978 (N_5978,N_5769,N_5874);
nor U5979 (N_5979,N_5754,N_5760);
and U5980 (N_5980,N_5810,N_5766);
nand U5981 (N_5981,N_5788,N_5846);
and U5982 (N_5982,N_5780,N_5814);
xnor U5983 (N_5983,N_5763,N_5865);
or U5984 (N_5984,N_5866,N_5795);
nor U5985 (N_5985,N_5857,N_5872);
xor U5986 (N_5986,N_5825,N_5821);
or U5987 (N_5987,N_5839,N_5817);
or U5988 (N_5988,N_5785,N_5754);
nor U5989 (N_5989,N_5764,N_5795);
and U5990 (N_5990,N_5846,N_5814);
or U5991 (N_5991,N_5798,N_5867);
and U5992 (N_5992,N_5800,N_5874);
nand U5993 (N_5993,N_5777,N_5824);
or U5994 (N_5994,N_5868,N_5847);
nand U5995 (N_5995,N_5755,N_5790);
and U5996 (N_5996,N_5798,N_5782);
or U5997 (N_5997,N_5772,N_5794);
and U5998 (N_5998,N_5758,N_5828);
xnor U5999 (N_5999,N_5799,N_5817);
and U6000 (N_6000,N_5949,N_5913);
nand U6001 (N_6001,N_5984,N_5914);
nand U6002 (N_6002,N_5940,N_5965);
or U6003 (N_6003,N_5973,N_5935);
or U6004 (N_6004,N_5939,N_5921);
xnor U6005 (N_6005,N_5999,N_5968);
nor U6006 (N_6006,N_5922,N_5900);
and U6007 (N_6007,N_5946,N_5964);
xor U6008 (N_6008,N_5891,N_5896);
or U6009 (N_6009,N_5976,N_5928);
or U6010 (N_6010,N_5972,N_5986);
nand U6011 (N_6011,N_5993,N_5992);
or U6012 (N_6012,N_5907,N_5967);
and U6013 (N_6013,N_5994,N_5969);
nor U6014 (N_6014,N_5987,N_5941);
or U6015 (N_6015,N_5944,N_5953);
nor U6016 (N_6016,N_5897,N_5936);
or U6017 (N_6017,N_5954,N_5945);
nor U6018 (N_6018,N_5962,N_5925);
or U6019 (N_6019,N_5981,N_5929);
and U6020 (N_6020,N_5957,N_5924);
nand U6021 (N_6021,N_5917,N_5885);
xor U6022 (N_6022,N_5876,N_5956);
or U6023 (N_6023,N_5980,N_5899);
nand U6024 (N_6024,N_5923,N_5970);
and U6025 (N_6025,N_5995,N_5892);
and U6026 (N_6026,N_5966,N_5895);
and U6027 (N_6027,N_5943,N_5938);
xor U6028 (N_6028,N_5958,N_5880);
or U6029 (N_6029,N_5979,N_5988);
and U6030 (N_6030,N_5877,N_5911);
or U6031 (N_6031,N_5983,N_5961);
xor U6032 (N_6032,N_5991,N_5950);
nand U6033 (N_6033,N_5919,N_5898);
and U6034 (N_6034,N_5893,N_5906);
nor U6035 (N_6035,N_5916,N_5878);
nor U6036 (N_6036,N_5989,N_5875);
nand U6037 (N_6037,N_5930,N_5932);
and U6038 (N_6038,N_5890,N_5975);
nand U6039 (N_6039,N_5998,N_5977);
xnor U6040 (N_6040,N_5902,N_5905);
nor U6041 (N_6041,N_5951,N_5886);
and U6042 (N_6042,N_5934,N_5909);
xnor U6043 (N_6043,N_5971,N_5910);
or U6044 (N_6044,N_5948,N_5974);
xnor U6045 (N_6045,N_5927,N_5912);
or U6046 (N_6046,N_5920,N_5888);
or U6047 (N_6047,N_5889,N_5997);
and U6048 (N_6048,N_5894,N_5879);
nand U6049 (N_6049,N_5996,N_5963);
xnor U6050 (N_6050,N_5959,N_5887);
xnor U6051 (N_6051,N_5882,N_5908);
and U6052 (N_6052,N_5955,N_5904);
nor U6053 (N_6053,N_5881,N_5903);
and U6054 (N_6054,N_5931,N_5937);
xor U6055 (N_6055,N_5982,N_5942);
or U6056 (N_6056,N_5978,N_5901);
xnor U6057 (N_6057,N_5933,N_5947);
nand U6058 (N_6058,N_5915,N_5990);
nand U6059 (N_6059,N_5960,N_5985);
xor U6060 (N_6060,N_5952,N_5918);
xor U6061 (N_6061,N_5883,N_5926);
and U6062 (N_6062,N_5884,N_5998);
xor U6063 (N_6063,N_5883,N_5880);
or U6064 (N_6064,N_5973,N_5946);
or U6065 (N_6065,N_5887,N_5875);
nor U6066 (N_6066,N_5980,N_5910);
and U6067 (N_6067,N_5954,N_5903);
nand U6068 (N_6068,N_5881,N_5955);
or U6069 (N_6069,N_5896,N_5895);
or U6070 (N_6070,N_5943,N_5910);
nand U6071 (N_6071,N_5998,N_5883);
and U6072 (N_6072,N_5969,N_5998);
xnor U6073 (N_6073,N_5937,N_5990);
nor U6074 (N_6074,N_5971,N_5989);
nor U6075 (N_6075,N_5905,N_5889);
or U6076 (N_6076,N_5916,N_5942);
nor U6077 (N_6077,N_5976,N_5978);
and U6078 (N_6078,N_5954,N_5942);
xnor U6079 (N_6079,N_5981,N_5978);
or U6080 (N_6080,N_5896,N_5978);
nand U6081 (N_6081,N_5911,N_5906);
and U6082 (N_6082,N_5931,N_5903);
nor U6083 (N_6083,N_5932,N_5903);
or U6084 (N_6084,N_5921,N_5879);
and U6085 (N_6085,N_5906,N_5947);
nor U6086 (N_6086,N_5935,N_5942);
or U6087 (N_6087,N_5960,N_5905);
or U6088 (N_6088,N_5992,N_5970);
nand U6089 (N_6089,N_5976,N_5879);
nand U6090 (N_6090,N_5903,N_5875);
and U6091 (N_6091,N_5992,N_5902);
or U6092 (N_6092,N_5922,N_5928);
nand U6093 (N_6093,N_5945,N_5972);
nand U6094 (N_6094,N_5952,N_5980);
and U6095 (N_6095,N_5947,N_5910);
nor U6096 (N_6096,N_5931,N_5924);
and U6097 (N_6097,N_5915,N_5913);
nor U6098 (N_6098,N_5926,N_5970);
nand U6099 (N_6099,N_5966,N_5949);
or U6100 (N_6100,N_5878,N_5881);
nand U6101 (N_6101,N_5917,N_5902);
and U6102 (N_6102,N_5900,N_5989);
or U6103 (N_6103,N_5994,N_5885);
or U6104 (N_6104,N_5908,N_5984);
and U6105 (N_6105,N_5962,N_5973);
or U6106 (N_6106,N_5976,N_5895);
nand U6107 (N_6107,N_5980,N_5945);
xnor U6108 (N_6108,N_5893,N_5923);
xor U6109 (N_6109,N_5917,N_5931);
or U6110 (N_6110,N_5955,N_5936);
nand U6111 (N_6111,N_5922,N_5982);
xor U6112 (N_6112,N_5913,N_5937);
xnor U6113 (N_6113,N_5972,N_5974);
or U6114 (N_6114,N_5945,N_5947);
nand U6115 (N_6115,N_5921,N_5906);
xnor U6116 (N_6116,N_5888,N_5909);
nand U6117 (N_6117,N_5906,N_5922);
nor U6118 (N_6118,N_5980,N_5999);
and U6119 (N_6119,N_5922,N_5974);
xor U6120 (N_6120,N_5881,N_5947);
nor U6121 (N_6121,N_5994,N_5907);
and U6122 (N_6122,N_5898,N_5986);
or U6123 (N_6123,N_5881,N_5884);
nand U6124 (N_6124,N_5944,N_5931);
xor U6125 (N_6125,N_6054,N_6006);
or U6126 (N_6126,N_6059,N_6041);
nand U6127 (N_6127,N_6107,N_6042);
and U6128 (N_6128,N_6077,N_6075);
xnor U6129 (N_6129,N_6114,N_6087);
xor U6130 (N_6130,N_6074,N_6035);
xnor U6131 (N_6131,N_6031,N_6089);
or U6132 (N_6132,N_6033,N_6084);
nor U6133 (N_6133,N_6000,N_6108);
nor U6134 (N_6134,N_6009,N_6069);
and U6135 (N_6135,N_6039,N_6081);
or U6136 (N_6136,N_6121,N_6021);
or U6137 (N_6137,N_6123,N_6044);
and U6138 (N_6138,N_6118,N_6051);
and U6139 (N_6139,N_6063,N_6097);
nand U6140 (N_6140,N_6112,N_6022);
and U6141 (N_6141,N_6115,N_6113);
and U6142 (N_6142,N_6048,N_6028);
xor U6143 (N_6143,N_6030,N_6052);
and U6144 (N_6144,N_6017,N_6018);
nand U6145 (N_6145,N_6082,N_6090);
nor U6146 (N_6146,N_6080,N_6029);
nand U6147 (N_6147,N_6057,N_6116);
or U6148 (N_6148,N_6124,N_6046);
nand U6149 (N_6149,N_6014,N_6008);
or U6150 (N_6150,N_6070,N_6056);
nand U6151 (N_6151,N_6076,N_6013);
or U6152 (N_6152,N_6037,N_6104);
and U6153 (N_6153,N_6105,N_6010);
or U6154 (N_6154,N_6064,N_6120);
and U6155 (N_6155,N_6117,N_6004);
nand U6156 (N_6156,N_6012,N_6060);
xor U6157 (N_6157,N_6002,N_6110);
nor U6158 (N_6158,N_6016,N_6055);
nand U6159 (N_6159,N_6065,N_6111);
nand U6160 (N_6160,N_6071,N_6019);
xor U6161 (N_6161,N_6091,N_6062);
and U6162 (N_6162,N_6106,N_6027);
and U6163 (N_6163,N_6015,N_6047);
and U6164 (N_6164,N_6026,N_6045);
nand U6165 (N_6165,N_6073,N_6086);
nand U6166 (N_6166,N_6020,N_6061);
nor U6167 (N_6167,N_6066,N_6102);
nor U6168 (N_6168,N_6109,N_6122);
nand U6169 (N_6169,N_6001,N_6023);
xnor U6170 (N_6170,N_6058,N_6085);
xnor U6171 (N_6171,N_6053,N_6093);
nor U6172 (N_6172,N_6005,N_6100);
xnor U6173 (N_6173,N_6043,N_6103);
xor U6174 (N_6174,N_6101,N_6068);
or U6175 (N_6175,N_6119,N_6096);
and U6176 (N_6176,N_6007,N_6050);
xnor U6177 (N_6177,N_6079,N_6094);
nor U6178 (N_6178,N_6049,N_6036);
nor U6179 (N_6179,N_6088,N_6078);
nand U6180 (N_6180,N_6003,N_6072);
nand U6181 (N_6181,N_6038,N_6099);
nor U6182 (N_6182,N_6098,N_6092);
and U6183 (N_6183,N_6011,N_6067);
and U6184 (N_6184,N_6083,N_6040);
nand U6185 (N_6185,N_6025,N_6024);
or U6186 (N_6186,N_6095,N_6032);
or U6187 (N_6187,N_6034,N_6110);
xnor U6188 (N_6188,N_6115,N_6118);
or U6189 (N_6189,N_6056,N_6013);
nor U6190 (N_6190,N_6113,N_6016);
nor U6191 (N_6191,N_6054,N_6025);
nor U6192 (N_6192,N_6018,N_6013);
or U6193 (N_6193,N_6097,N_6105);
nand U6194 (N_6194,N_6000,N_6085);
nor U6195 (N_6195,N_6057,N_6071);
and U6196 (N_6196,N_6069,N_6078);
or U6197 (N_6197,N_6013,N_6082);
or U6198 (N_6198,N_6031,N_6096);
nor U6199 (N_6199,N_6077,N_6038);
or U6200 (N_6200,N_6071,N_6056);
nand U6201 (N_6201,N_6046,N_6063);
and U6202 (N_6202,N_6058,N_6011);
and U6203 (N_6203,N_6069,N_6008);
or U6204 (N_6204,N_6037,N_6103);
and U6205 (N_6205,N_6083,N_6018);
nor U6206 (N_6206,N_6099,N_6095);
nor U6207 (N_6207,N_6060,N_6041);
nand U6208 (N_6208,N_6095,N_6008);
or U6209 (N_6209,N_6061,N_6021);
or U6210 (N_6210,N_6009,N_6097);
and U6211 (N_6211,N_6052,N_6005);
xor U6212 (N_6212,N_6055,N_6046);
nand U6213 (N_6213,N_6108,N_6003);
xnor U6214 (N_6214,N_6073,N_6113);
nand U6215 (N_6215,N_6057,N_6123);
and U6216 (N_6216,N_6013,N_6120);
nand U6217 (N_6217,N_6043,N_6023);
xnor U6218 (N_6218,N_6018,N_6108);
nor U6219 (N_6219,N_6018,N_6045);
or U6220 (N_6220,N_6073,N_6060);
and U6221 (N_6221,N_6014,N_6090);
and U6222 (N_6222,N_6065,N_6106);
nor U6223 (N_6223,N_6015,N_6068);
xnor U6224 (N_6224,N_6001,N_6005);
and U6225 (N_6225,N_6024,N_6049);
and U6226 (N_6226,N_6115,N_6044);
nor U6227 (N_6227,N_6098,N_6089);
or U6228 (N_6228,N_6073,N_6001);
and U6229 (N_6229,N_6058,N_6121);
nor U6230 (N_6230,N_6084,N_6094);
nand U6231 (N_6231,N_6076,N_6043);
nand U6232 (N_6232,N_6075,N_6048);
nor U6233 (N_6233,N_6001,N_6041);
nand U6234 (N_6234,N_6031,N_6012);
nor U6235 (N_6235,N_6085,N_6042);
or U6236 (N_6236,N_6072,N_6109);
nor U6237 (N_6237,N_6105,N_6025);
nand U6238 (N_6238,N_6053,N_6089);
and U6239 (N_6239,N_6120,N_6105);
and U6240 (N_6240,N_6030,N_6095);
xor U6241 (N_6241,N_6118,N_6092);
nor U6242 (N_6242,N_6046,N_6071);
nand U6243 (N_6243,N_6122,N_6044);
nor U6244 (N_6244,N_6017,N_6004);
or U6245 (N_6245,N_6117,N_6091);
nor U6246 (N_6246,N_6003,N_6050);
or U6247 (N_6247,N_6011,N_6030);
nor U6248 (N_6248,N_6109,N_6096);
nand U6249 (N_6249,N_6027,N_6073);
or U6250 (N_6250,N_6126,N_6202);
and U6251 (N_6251,N_6154,N_6169);
xor U6252 (N_6252,N_6177,N_6148);
nand U6253 (N_6253,N_6240,N_6193);
nand U6254 (N_6254,N_6179,N_6164);
xor U6255 (N_6255,N_6231,N_6138);
nor U6256 (N_6256,N_6132,N_6173);
nor U6257 (N_6257,N_6158,N_6221);
xor U6258 (N_6258,N_6199,N_6232);
nor U6259 (N_6259,N_6207,N_6224);
xor U6260 (N_6260,N_6215,N_6239);
nand U6261 (N_6261,N_6189,N_6166);
nor U6262 (N_6262,N_6219,N_6162);
xor U6263 (N_6263,N_6180,N_6181);
or U6264 (N_6264,N_6128,N_6156);
and U6265 (N_6265,N_6139,N_6125);
xor U6266 (N_6266,N_6212,N_6135);
nand U6267 (N_6267,N_6178,N_6238);
nor U6268 (N_6268,N_6220,N_6229);
nor U6269 (N_6269,N_6226,N_6137);
and U6270 (N_6270,N_6203,N_6161);
nand U6271 (N_6271,N_6140,N_6144);
or U6272 (N_6272,N_6210,N_6227);
nand U6273 (N_6273,N_6223,N_6211);
and U6274 (N_6274,N_6142,N_6172);
xnor U6275 (N_6275,N_6242,N_6194);
and U6276 (N_6276,N_6206,N_6133);
and U6277 (N_6277,N_6213,N_6191);
or U6278 (N_6278,N_6136,N_6197);
nand U6279 (N_6279,N_6237,N_6217);
and U6280 (N_6280,N_6149,N_6205);
xnor U6281 (N_6281,N_6170,N_6186);
xnor U6282 (N_6282,N_6190,N_6235);
xnor U6283 (N_6283,N_6160,N_6214);
and U6284 (N_6284,N_6188,N_6152);
xnor U6285 (N_6285,N_6146,N_6150);
xor U6286 (N_6286,N_6228,N_6168);
nand U6287 (N_6287,N_6244,N_6183);
nand U6288 (N_6288,N_6187,N_6155);
xnor U6289 (N_6289,N_6167,N_6165);
or U6290 (N_6290,N_6241,N_6182);
and U6291 (N_6291,N_6176,N_6233);
or U6292 (N_6292,N_6201,N_6245);
or U6293 (N_6293,N_6174,N_6209);
nand U6294 (N_6294,N_6196,N_6218);
nor U6295 (N_6295,N_6200,N_6157);
nor U6296 (N_6296,N_6243,N_6130);
xnor U6297 (N_6297,N_6192,N_6127);
nand U6298 (N_6298,N_6195,N_6225);
nor U6299 (N_6299,N_6141,N_6184);
and U6300 (N_6300,N_6131,N_6175);
and U6301 (N_6301,N_6222,N_6153);
or U6302 (N_6302,N_6145,N_6230);
xnor U6303 (N_6303,N_6151,N_6159);
or U6304 (N_6304,N_6134,N_6185);
xnor U6305 (N_6305,N_6143,N_6249);
nor U6306 (N_6306,N_6147,N_6246);
or U6307 (N_6307,N_6247,N_6204);
nor U6308 (N_6308,N_6198,N_6216);
nand U6309 (N_6309,N_6236,N_6234);
and U6310 (N_6310,N_6208,N_6171);
nand U6311 (N_6311,N_6129,N_6163);
xor U6312 (N_6312,N_6248,N_6145);
and U6313 (N_6313,N_6135,N_6131);
nand U6314 (N_6314,N_6228,N_6235);
nand U6315 (N_6315,N_6237,N_6172);
nor U6316 (N_6316,N_6168,N_6181);
nand U6317 (N_6317,N_6234,N_6209);
and U6318 (N_6318,N_6127,N_6243);
or U6319 (N_6319,N_6130,N_6197);
nor U6320 (N_6320,N_6223,N_6131);
or U6321 (N_6321,N_6126,N_6215);
nand U6322 (N_6322,N_6159,N_6168);
nor U6323 (N_6323,N_6160,N_6223);
nor U6324 (N_6324,N_6189,N_6134);
or U6325 (N_6325,N_6177,N_6247);
nand U6326 (N_6326,N_6125,N_6162);
or U6327 (N_6327,N_6191,N_6155);
nor U6328 (N_6328,N_6220,N_6200);
and U6329 (N_6329,N_6128,N_6242);
nand U6330 (N_6330,N_6232,N_6176);
nor U6331 (N_6331,N_6195,N_6169);
or U6332 (N_6332,N_6234,N_6215);
and U6333 (N_6333,N_6171,N_6201);
nand U6334 (N_6334,N_6133,N_6182);
and U6335 (N_6335,N_6236,N_6135);
nand U6336 (N_6336,N_6129,N_6136);
or U6337 (N_6337,N_6174,N_6211);
nand U6338 (N_6338,N_6186,N_6171);
xor U6339 (N_6339,N_6132,N_6127);
xnor U6340 (N_6340,N_6140,N_6137);
nor U6341 (N_6341,N_6229,N_6199);
xor U6342 (N_6342,N_6227,N_6129);
xnor U6343 (N_6343,N_6236,N_6241);
xor U6344 (N_6344,N_6173,N_6214);
xor U6345 (N_6345,N_6147,N_6142);
nor U6346 (N_6346,N_6243,N_6201);
or U6347 (N_6347,N_6213,N_6200);
and U6348 (N_6348,N_6216,N_6134);
or U6349 (N_6349,N_6219,N_6221);
and U6350 (N_6350,N_6155,N_6197);
or U6351 (N_6351,N_6195,N_6176);
xor U6352 (N_6352,N_6232,N_6182);
xor U6353 (N_6353,N_6222,N_6231);
xnor U6354 (N_6354,N_6170,N_6227);
nor U6355 (N_6355,N_6234,N_6187);
xor U6356 (N_6356,N_6139,N_6191);
nor U6357 (N_6357,N_6237,N_6242);
and U6358 (N_6358,N_6213,N_6125);
nor U6359 (N_6359,N_6181,N_6220);
or U6360 (N_6360,N_6228,N_6245);
xor U6361 (N_6361,N_6175,N_6215);
and U6362 (N_6362,N_6200,N_6242);
nand U6363 (N_6363,N_6247,N_6205);
nor U6364 (N_6364,N_6178,N_6235);
nand U6365 (N_6365,N_6247,N_6145);
nor U6366 (N_6366,N_6191,N_6175);
or U6367 (N_6367,N_6181,N_6245);
or U6368 (N_6368,N_6129,N_6210);
nor U6369 (N_6369,N_6131,N_6232);
nor U6370 (N_6370,N_6138,N_6142);
nand U6371 (N_6371,N_6142,N_6127);
nor U6372 (N_6372,N_6237,N_6164);
nand U6373 (N_6373,N_6157,N_6245);
nand U6374 (N_6374,N_6229,N_6166);
nor U6375 (N_6375,N_6374,N_6360);
and U6376 (N_6376,N_6266,N_6340);
and U6377 (N_6377,N_6313,N_6322);
nor U6378 (N_6378,N_6263,N_6350);
or U6379 (N_6379,N_6287,N_6304);
and U6380 (N_6380,N_6272,N_6297);
or U6381 (N_6381,N_6311,N_6283);
nor U6382 (N_6382,N_6326,N_6342);
and U6383 (N_6383,N_6300,N_6286);
nand U6384 (N_6384,N_6367,N_6373);
or U6385 (N_6385,N_6332,N_6250);
nor U6386 (N_6386,N_6267,N_6278);
and U6387 (N_6387,N_6294,N_6336);
or U6388 (N_6388,N_6292,N_6371);
nor U6389 (N_6389,N_6252,N_6254);
and U6390 (N_6390,N_6259,N_6366);
and U6391 (N_6391,N_6256,N_6329);
nor U6392 (N_6392,N_6344,N_6302);
and U6393 (N_6393,N_6265,N_6312);
nor U6394 (N_6394,N_6273,N_6368);
xor U6395 (N_6395,N_6306,N_6330);
nand U6396 (N_6396,N_6298,N_6264);
xnor U6397 (N_6397,N_6347,N_6277);
xnor U6398 (N_6398,N_6321,N_6258);
xor U6399 (N_6399,N_6372,N_6318);
nor U6400 (N_6400,N_6315,N_6310);
nor U6401 (N_6401,N_6349,N_6276);
and U6402 (N_6402,N_6328,N_6325);
and U6403 (N_6403,N_6357,N_6285);
nor U6404 (N_6404,N_6296,N_6324);
nor U6405 (N_6405,N_6274,N_6290);
nand U6406 (N_6406,N_6337,N_6316);
nand U6407 (N_6407,N_6345,N_6269);
and U6408 (N_6408,N_6320,N_6352);
nand U6409 (N_6409,N_6295,N_6308);
and U6410 (N_6410,N_6351,N_6335);
or U6411 (N_6411,N_6370,N_6288);
nor U6412 (N_6412,N_6281,N_6359);
and U6413 (N_6413,N_6339,N_6251);
and U6414 (N_6414,N_6334,N_6364);
nand U6415 (N_6415,N_6346,N_6305);
or U6416 (N_6416,N_6343,N_6279);
xor U6417 (N_6417,N_6282,N_6307);
nand U6418 (N_6418,N_6365,N_6356);
and U6419 (N_6419,N_6323,N_6341);
nor U6420 (N_6420,N_6319,N_6253);
or U6421 (N_6421,N_6301,N_6348);
or U6422 (N_6422,N_6363,N_6280);
nand U6423 (N_6423,N_6262,N_6333);
and U6424 (N_6424,N_6314,N_6255);
nand U6425 (N_6425,N_6362,N_6353);
or U6426 (N_6426,N_6369,N_6293);
nand U6427 (N_6427,N_6338,N_6358);
and U6428 (N_6428,N_6309,N_6317);
xnor U6429 (N_6429,N_6260,N_6299);
and U6430 (N_6430,N_6257,N_6284);
and U6431 (N_6431,N_6271,N_6261);
or U6432 (N_6432,N_6270,N_6275);
xnor U6433 (N_6433,N_6331,N_6289);
nor U6434 (N_6434,N_6355,N_6354);
xnor U6435 (N_6435,N_6361,N_6327);
xnor U6436 (N_6436,N_6303,N_6291);
nor U6437 (N_6437,N_6268,N_6275);
or U6438 (N_6438,N_6348,N_6290);
and U6439 (N_6439,N_6331,N_6346);
or U6440 (N_6440,N_6339,N_6304);
or U6441 (N_6441,N_6322,N_6261);
or U6442 (N_6442,N_6323,N_6302);
xor U6443 (N_6443,N_6336,N_6305);
and U6444 (N_6444,N_6363,N_6318);
nor U6445 (N_6445,N_6336,N_6346);
xnor U6446 (N_6446,N_6372,N_6317);
nand U6447 (N_6447,N_6327,N_6308);
nand U6448 (N_6448,N_6360,N_6334);
or U6449 (N_6449,N_6336,N_6258);
xnor U6450 (N_6450,N_6326,N_6252);
nand U6451 (N_6451,N_6307,N_6326);
or U6452 (N_6452,N_6267,N_6344);
or U6453 (N_6453,N_6252,N_6315);
or U6454 (N_6454,N_6344,N_6292);
nand U6455 (N_6455,N_6337,N_6299);
or U6456 (N_6456,N_6348,N_6261);
nand U6457 (N_6457,N_6256,N_6361);
nor U6458 (N_6458,N_6323,N_6250);
nand U6459 (N_6459,N_6333,N_6294);
xnor U6460 (N_6460,N_6273,N_6374);
or U6461 (N_6461,N_6357,N_6360);
xor U6462 (N_6462,N_6297,N_6319);
or U6463 (N_6463,N_6365,N_6315);
nor U6464 (N_6464,N_6370,N_6374);
nand U6465 (N_6465,N_6284,N_6330);
xor U6466 (N_6466,N_6252,N_6363);
and U6467 (N_6467,N_6271,N_6317);
nor U6468 (N_6468,N_6351,N_6259);
or U6469 (N_6469,N_6309,N_6329);
nand U6470 (N_6470,N_6298,N_6289);
nand U6471 (N_6471,N_6368,N_6304);
xnor U6472 (N_6472,N_6352,N_6316);
or U6473 (N_6473,N_6264,N_6291);
or U6474 (N_6474,N_6337,N_6279);
nand U6475 (N_6475,N_6365,N_6374);
nor U6476 (N_6476,N_6346,N_6256);
xor U6477 (N_6477,N_6255,N_6362);
or U6478 (N_6478,N_6265,N_6267);
nand U6479 (N_6479,N_6350,N_6339);
and U6480 (N_6480,N_6343,N_6367);
and U6481 (N_6481,N_6310,N_6291);
nand U6482 (N_6482,N_6258,N_6293);
nand U6483 (N_6483,N_6288,N_6368);
or U6484 (N_6484,N_6250,N_6296);
xnor U6485 (N_6485,N_6254,N_6293);
nand U6486 (N_6486,N_6322,N_6352);
nor U6487 (N_6487,N_6275,N_6353);
nor U6488 (N_6488,N_6313,N_6265);
nor U6489 (N_6489,N_6355,N_6353);
and U6490 (N_6490,N_6269,N_6284);
or U6491 (N_6491,N_6298,N_6332);
xnor U6492 (N_6492,N_6286,N_6313);
xnor U6493 (N_6493,N_6370,N_6310);
nand U6494 (N_6494,N_6333,N_6373);
nor U6495 (N_6495,N_6357,N_6321);
nand U6496 (N_6496,N_6359,N_6268);
and U6497 (N_6497,N_6309,N_6336);
and U6498 (N_6498,N_6348,N_6292);
nand U6499 (N_6499,N_6256,N_6260);
or U6500 (N_6500,N_6381,N_6379);
or U6501 (N_6501,N_6499,N_6462);
or U6502 (N_6502,N_6495,N_6424);
or U6503 (N_6503,N_6484,N_6392);
nor U6504 (N_6504,N_6446,N_6464);
nor U6505 (N_6505,N_6498,N_6399);
nor U6506 (N_6506,N_6445,N_6442);
nor U6507 (N_6507,N_6489,N_6454);
nor U6508 (N_6508,N_6453,N_6376);
xnor U6509 (N_6509,N_6401,N_6444);
nand U6510 (N_6510,N_6459,N_6476);
xor U6511 (N_6511,N_6490,N_6428);
nor U6512 (N_6512,N_6429,N_6452);
and U6513 (N_6513,N_6477,N_6485);
or U6514 (N_6514,N_6410,N_6440);
and U6515 (N_6515,N_6411,N_6397);
and U6516 (N_6516,N_6467,N_6417);
and U6517 (N_6517,N_6449,N_6405);
nor U6518 (N_6518,N_6390,N_6393);
or U6519 (N_6519,N_6472,N_6481);
nand U6520 (N_6520,N_6461,N_6385);
nor U6521 (N_6521,N_6422,N_6407);
or U6522 (N_6522,N_6404,N_6395);
or U6523 (N_6523,N_6427,N_6387);
or U6524 (N_6524,N_6473,N_6434);
or U6525 (N_6525,N_6491,N_6415);
or U6526 (N_6526,N_6488,N_6466);
and U6527 (N_6527,N_6469,N_6460);
nor U6528 (N_6528,N_6403,N_6439);
xnor U6529 (N_6529,N_6497,N_6419);
and U6530 (N_6530,N_6414,N_6377);
or U6531 (N_6531,N_6447,N_6443);
nand U6532 (N_6532,N_6420,N_6425);
nand U6533 (N_6533,N_6430,N_6475);
xnor U6534 (N_6534,N_6435,N_6400);
or U6535 (N_6535,N_6451,N_6386);
nand U6536 (N_6536,N_6431,N_6486);
nand U6537 (N_6537,N_6436,N_6474);
or U6538 (N_6538,N_6450,N_6480);
nor U6539 (N_6539,N_6478,N_6383);
xor U6540 (N_6540,N_6468,N_6413);
or U6541 (N_6541,N_6388,N_6406);
and U6542 (N_6542,N_6448,N_6412);
nand U6543 (N_6543,N_6426,N_6441);
xnor U6544 (N_6544,N_6384,N_6375);
nand U6545 (N_6545,N_6457,N_6437);
and U6546 (N_6546,N_6487,N_6391);
xor U6547 (N_6547,N_6432,N_6380);
and U6548 (N_6548,N_6394,N_6389);
xor U6549 (N_6549,N_6409,N_6479);
nor U6550 (N_6550,N_6493,N_6416);
and U6551 (N_6551,N_6455,N_6421);
or U6552 (N_6552,N_6458,N_6496);
and U6553 (N_6553,N_6456,N_6396);
nand U6554 (N_6554,N_6470,N_6382);
nor U6555 (N_6555,N_6378,N_6492);
or U6556 (N_6556,N_6465,N_6408);
nor U6557 (N_6557,N_6471,N_6482);
nor U6558 (N_6558,N_6463,N_6402);
and U6559 (N_6559,N_6423,N_6494);
xnor U6560 (N_6560,N_6398,N_6438);
nor U6561 (N_6561,N_6418,N_6483);
or U6562 (N_6562,N_6433,N_6444);
nand U6563 (N_6563,N_6457,N_6408);
and U6564 (N_6564,N_6420,N_6484);
or U6565 (N_6565,N_6459,N_6472);
or U6566 (N_6566,N_6399,N_6450);
nand U6567 (N_6567,N_6486,N_6492);
and U6568 (N_6568,N_6499,N_6406);
nand U6569 (N_6569,N_6413,N_6387);
and U6570 (N_6570,N_6474,N_6482);
and U6571 (N_6571,N_6396,N_6415);
or U6572 (N_6572,N_6416,N_6391);
and U6573 (N_6573,N_6432,N_6480);
and U6574 (N_6574,N_6375,N_6416);
nand U6575 (N_6575,N_6428,N_6394);
xnor U6576 (N_6576,N_6379,N_6429);
and U6577 (N_6577,N_6422,N_6409);
nor U6578 (N_6578,N_6490,N_6397);
xnor U6579 (N_6579,N_6415,N_6384);
nand U6580 (N_6580,N_6397,N_6473);
or U6581 (N_6581,N_6453,N_6472);
xnor U6582 (N_6582,N_6431,N_6394);
nand U6583 (N_6583,N_6418,N_6432);
nand U6584 (N_6584,N_6405,N_6444);
xor U6585 (N_6585,N_6497,N_6415);
nor U6586 (N_6586,N_6377,N_6407);
nand U6587 (N_6587,N_6437,N_6458);
or U6588 (N_6588,N_6431,N_6424);
nand U6589 (N_6589,N_6420,N_6437);
and U6590 (N_6590,N_6407,N_6472);
or U6591 (N_6591,N_6400,N_6484);
or U6592 (N_6592,N_6496,N_6414);
xor U6593 (N_6593,N_6404,N_6396);
or U6594 (N_6594,N_6430,N_6465);
and U6595 (N_6595,N_6459,N_6417);
nand U6596 (N_6596,N_6398,N_6417);
nor U6597 (N_6597,N_6418,N_6480);
or U6598 (N_6598,N_6391,N_6494);
nor U6599 (N_6599,N_6378,N_6403);
nor U6600 (N_6600,N_6485,N_6431);
or U6601 (N_6601,N_6488,N_6431);
xor U6602 (N_6602,N_6453,N_6450);
and U6603 (N_6603,N_6393,N_6499);
and U6604 (N_6604,N_6424,N_6483);
nor U6605 (N_6605,N_6478,N_6428);
nor U6606 (N_6606,N_6375,N_6491);
or U6607 (N_6607,N_6455,N_6407);
xnor U6608 (N_6608,N_6432,N_6419);
nor U6609 (N_6609,N_6423,N_6393);
or U6610 (N_6610,N_6493,N_6377);
nor U6611 (N_6611,N_6390,N_6447);
or U6612 (N_6612,N_6385,N_6453);
nor U6613 (N_6613,N_6406,N_6383);
or U6614 (N_6614,N_6479,N_6383);
xnor U6615 (N_6615,N_6443,N_6476);
nand U6616 (N_6616,N_6440,N_6473);
nor U6617 (N_6617,N_6415,N_6431);
and U6618 (N_6618,N_6401,N_6402);
and U6619 (N_6619,N_6438,N_6442);
xor U6620 (N_6620,N_6411,N_6392);
or U6621 (N_6621,N_6397,N_6499);
and U6622 (N_6622,N_6485,N_6451);
and U6623 (N_6623,N_6480,N_6453);
and U6624 (N_6624,N_6380,N_6456);
and U6625 (N_6625,N_6522,N_6574);
nand U6626 (N_6626,N_6605,N_6548);
or U6627 (N_6627,N_6551,N_6577);
and U6628 (N_6628,N_6545,N_6569);
nor U6629 (N_6629,N_6536,N_6599);
or U6630 (N_6630,N_6552,N_6521);
xnor U6631 (N_6631,N_6512,N_6510);
xor U6632 (N_6632,N_6612,N_6591);
and U6633 (N_6633,N_6554,N_6576);
or U6634 (N_6634,N_6558,N_6567);
nand U6635 (N_6635,N_6543,N_6562);
or U6636 (N_6636,N_6553,N_6618);
xnor U6637 (N_6637,N_6582,N_6578);
or U6638 (N_6638,N_6525,N_6570);
and U6639 (N_6639,N_6517,N_6595);
and U6640 (N_6640,N_6531,N_6624);
xor U6641 (N_6641,N_6559,N_6520);
nand U6642 (N_6642,N_6541,N_6588);
or U6643 (N_6643,N_6568,N_6593);
xnor U6644 (N_6644,N_6544,N_6565);
nor U6645 (N_6645,N_6523,N_6519);
xor U6646 (N_6646,N_6502,N_6583);
or U6647 (N_6647,N_6561,N_6623);
or U6648 (N_6648,N_6604,N_6547);
and U6649 (N_6649,N_6530,N_6613);
nand U6650 (N_6650,N_6563,N_6571);
nand U6651 (N_6651,N_6550,N_6617);
nor U6652 (N_6652,N_6556,N_6518);
and U6653 (N_6653,N_6513,N_6597);
and U6654 (N_6654,N_6590,N_6560);
and U6655 (N_6655,N_6608,N_6514);
nand U6656 (N_6656,N_6538,N_6616);
and U6657 (N_6657,N_6615,N_6620);
and U6658 (N_6658,N_6566,N_6603);
nor U6659 (N_6659,N_6506,N_6526);
and U6660 (N_6660,N_6508,N_6509);
nor U6661 (N_6661,N_6537,N_6528);
or U6662 (N_6662,N_6592,N_6533);
nand U6663 (N_6663,N_6622,N_6532);
xnor U6664 (N_6664,N_6580,N_6587);
xor U6665 (N_6665,N_6589,N_6607);
or U6666 (N_6666,N_6515,N_6542);
xor U6667 (N_6667,N_6579,N_6546);
nand U6668 (N_6668,N_6524,N_6572);
nand U6669 (N_6669,N_6606,N_6534);
and U6670 (N_6670,N_6564,N_6601);
nor U6671 (N_6671,N_6555,N_6602);
nand U6672 (N_6672,N_6507,N_6540);
xor U6673 (N_6673,N_6539,N_6619);
and U6674 (N_6674,N_6621,N_6557);
or U6675 (N_6675,N_6504,N_6600);
nand U6676 (N_6676,N_6611,N_6503);
or U6677 (N_6677,N_6575,N_6596);
nand U6678 (N_6678,N_6610,N_6535);
xor U6679 (N_6679,N_6584,N_6581);
xor U6680 (N_6680,N_6529,N_6549);
nand U6681 (N_6681,N_6501,N_6585);
nor U6682 (N_6682,N_6594,N_6516);
nor U6683 (N_6683,N_6586,N_6573);
and U6684 (N_6684,N_6614,N_6505);
nor U6685 (N_6685,N_6598,N_6511);
and U6686 (N_6686,N_6609,N_6500);
nor U6687 (N_6687,N_6527,N_6521);
xor U6688 (N_6688,N_6512,N_6550);
xor U6689 (N_6689,N_6583,N_6544);
xnor U6690 (N_6690,N_6622,N_6580);
xnor U6691 (N_6691,N_6622,N_6525);
nand U6692 (N_6692,N_6605,N_6621);
and U6693 (N_6693,N_6546,N_6607);
or U6694 (N_6694,N_6582,N_6552);
and U6695 (N_6695,N_6601,N_6566);
xor U6696 (N_6696,N_6573,N_6504);
xnor U6697 (N_6697,N_6608,N_6538);
nand U6698 (N_6698,N_6590,N_6539);
nand U6699 (N_6699,N_6523,N_6614);
and U6700 (N_6700,N_6507,N_6568);
and U6701 (N_6701,N_6583,N_6541);
xor U6702 (N_6702,N_6552,N_6567);
or U6703 (N_6703,N_6598,N_6610);
xnor U6704 (N_6704,N_6600,N_6610);
and U6705 (N_6705,N_6619,N_6576);
nor U6706 (N_6706,N_6554,N_6613);
nor U6707 (N_6707,N_6575,N_6604);
or U6708 (N_6708,N_6603,N_6576);
xnor U6709 (N_6709,N_6578,N_6618);
nand U6710 (N_6710,N_6569,N_6505);
nor U6711 (N_6711,N_6507,N_6604);
nand U6712 (N_6712,N_6622,N_6552);
nand U6713 (N_6713,N_6583,N_6564);
and U6714 (N_6714,N_6590,N_6575);
xnor U6715 (N_6715,N_6571,N_6516);
and U6716 (N_6716,N_6527,N_6544);
and U6717 (N_6717,N_6596,N_6598);
xor U6718 (N_6718,N_6553,N_6609);
xor U6719 (N_6719,N_6608,N_6521);
xor U6720 (N_6720,N_6615,N_6613);
xor U6721 (N_6721,N_6569,N_6534);
or U6722 (N_6722,N_6561,N_6537);
nand U6723 (N_6723,N_6535,N_6555);
nand U6724 (N_6724,N_6533,N_6505);
nor U6725 (N_6725,N_6538,N_6577);
or U6726 (N_6726,N_6562,N_6585);
nand U6727 (N_6727,N_6596,N_6537);
xnor U6728 (N_6728,N_6550,N_6557);
and U6729 (N_6729,N_6597,N_6518);
nor U6730 (N_6730,N_6529,N_6576);
and U6731 (N_6731,N_6558,N_6527);
or U6732 (N_6732,N_6570,N_6566);
and U6733 (N_6733,N_6597,N_6552);
nand U6734 (N_6734,N_6512,N_6504);
nand U6735 (N_6735,N_6525,N_6559);
and U6736 (N_6736,N_6547,N_6609);
and U6737 (N_6737,N_6564,N_6559);
nand U6738 (N_6738,N_6548,N_6538);
and U6739 (N_6739,N_6623,N_6597);
or U6740 (N_6740,N_6602,N_6612);
nor U6741 (N_6741,N_6530,N_6520);
and U6742 (N_6742,N_6622,N_6530);
nor U6743 (N_6743,N_6500,N_6610);
and U6744 (N_6744,N_6519,N_6587);
or U6745 (N_6745,N_6503,N_6578);
nor U6746 (N_6746,N_6543,N_6591);
nand U6747 (N_6747,N_6595,N_6525);
or U6748 (N_6748,N_6562,N_6500);
or U6749 (N_6749,N_6601,N_6583);
and U6750 (N_6750,N_6641,N_6685);
nor U6751 (N_6751,N_6742,N_6705);
and U6752 (N_6752,N_6730,N_6694);
nand U6753 (N_6753,N_6650,N_6647);
and U6754 (N_6754,N_6630,N_6663);
xnor U6755 (N_6755,N_6662,N_6632);
nor U6756 (N_6756,N_6717,N_6748);
xnor U6757 (N_6757,N_6639,N_6655);
and U6758 (N_6758,N_6683,N_6688);
nor U6759 (N_6759,N_6687,N_6723);
and U6760 (N_6760,N_6698,N_6657);
nor U6761 (N_6761,N_6674,N_6697);
nor U6762 (N_6762,N_6669,N_6733);
xnor U6763 (N_6763,N_6671,N_6625);
and U6764 (N_6764,N_6649,N_6704);
nor U6765 (N_6765,N_6651,N_6713);
or U6766 (N_6766,N_6666,N_6749);
or U6767 (N_6767,N_6719,N_6696);
nor U6768 (N_6768,N_6736,N_6677);
xor U6769 (N_6769,N_6721,N_6627);
and U6770 (N_6770,N_6729,N_6712);
or U6771 (N_6771,N_6682,N_6728);
or U6772 (N_6772,N_6737,N_6680);
nand U6773 (N_6773,N_6628,N_6692);
or U6774 (N_6774,N_6701,N_6673);
and U6775 (N_6775,N_6700,N_6686);
and U6776 (N_6776,N_6722,N_6660);
or U6777 (N_6777,N_6714,N_6731);
or U6778 (N_6778,N_6732,N_6661);
and U6779 (N_6779,N_6726,N_6633);
and U6780 (N_6780,N_6653,N_6743);
nand U6781 (N_6781,N_6747,N_6646);
or U6782 (N_6782,N_6715,N_6645);
xnor U6783 (N_6783,N_6699,N_6690);
nor U6784 (N_6784,N_6739,N_6631);
or U6785 (N_6785,N_6711,N_6718);
nor U6786 (N_6786,N_6693,N_6635);
xnor U6787 (N_6787,N_6740,N_6695);
nand U6788 (N_6788,N_6707,N_6710);
or U6789 (N_6789,N_6702,N_6652);
nor U6790 (N_6790,N_6658,N_6643);
xor U6791 (N_6791,N_6744,N_6708);
or U6792 (N_6792,N_6706,N_6665);
and U6793 (N_6793,N_6637,N_6664);
or U6794 (N_6794,N_6640,N_6727);
xnor U6795 (N_6795,N_6745,N_6716);
xnor U6796 (N_6796,N_6738,N_6644);
nand U6797 (N_6797,N_6676,N_6654);
xor U6798 (N_6798,N_6629,N_6725);
and U6799 (N_6799,N_6668,N_6691);
nand U6800 (N_6800,N_6638,N_6675);
and U6801 (N_6801,N_6703,N_6720);
or U6802 (N_6802,N_6642,N_6681);
and U6803 (N_6803,N_6684,N_6741);
or U6804 (N_6804,N_6656,N_6746);
and U6805 (N_6805,N_6679,N_6667);
nand U6806 (N_6806,N_6626,N_6670);
xor U6807 (N_6807,N_6709,N_6659);
and U6808 (N_6808,N_6678,N_6648);
nor U6809 (N_6809,N_6735,N_6724);
and U6810 (N_6810,N_6634,N_6734);
nor U6811 (N_6811,N_6636,N_6672);
nor U6812 (N_6812,N_6689,N_6718);
nor U6813 (N_6813,N_6649,N_6687);
nand U6814 (N_6814,N_6641,N_6625);
or U6815 (N_6815,N_6723,N_6715);
nand U6816 (N_6816,N_6644,N_6627);
and U6817 (N_6817,N_6684,N_6747);
or U6818 (N_6818,N_6722,N_6645);
or U6819 (N_6819,N_6642,N_6722);
and U6820 (N_6820,N_6660,N_6733);
and U6821 (N_6821,N_6669,N_6667);
and U6822 (N_6822,N_6684,N_6636);
and U6823 (N_6823,N_6676,N_6736);
nor U6824 (N_6824,N_6737,N_6679);
nor U6825 (N_6825,N_6715,N_6681);
or U6826 (N_6826,N_6625,N_6638);
nor U6827 (N_6827,N_6679,N_6680);
xor U6828 (N_6828,N_6668,N_6625);
and U6829 (N_6829,N_6698,N_6712);
nor U6830 (N_6830,N_6672,N_6682);
nand U6831 (N_6831,N_6625,N_6635);
or U6832 (N_6832,N_6717,N_6660);
nor U6833 (N_6833,N_6721,N_6629);
xor U6834 (N_6834,N_6677,N_6659);
or U6835 (N_6835,N_6681,N_6645);
nor U6836 (N_6836,N_6667,N_6659);
xor U6837 (N_6837,N_6645,N_6686);
or U6838 (N_6838,N_6674,N_6656);
or U6839 (N_6839,N_6699,N_6728);
and U6840 (N_6840,N_6699,N_6629);
and U6841 (N_6841,N_6712,N_6630);
xor U6842 (N_6842,N_6703,N_6671);
xor U6843 (N_6843,N_6728,N_6660);
nor U6844 (N_6844,N_6732,N_6733);
nor U6845 (N_6845,N_6698,N_6629);
or U6846 (N_6846,N_6654,N_6733);
or U6847 (N_6847,N_6696,N_6665);
nor U6848 (N_6848,N_6669,N_6744);
and U6849 (N_6849,N_6721,N_6737);
xor U6850 (N_6850,N_6710,N_6626);
nor U6851 (N_6851,N_6632,N_6733);
xor U6852 (N_6852,N_6637,N_6670);
nor U6853 (N_6853,N_6723,N_6665);
xor U6854 (N_6854,N_6744,N_6707);
xor U6855 (N_6855,N_6727,N_6728);
or U6856 (N_6856,N_6638,N_6714);
xnor U6857 (N_6857,N_6686,N_6689);
nand U6858 (N_6858,N_6729,N_6716);
xor U6859 (N_6859,N_6743,N_6637);
and U6860 (N_6860,N_6650,N_6629);
xor U6861 (N_6861,N_6728,N_6702);
nor U6862 (N_6862,N_6680,N_6667);
xor U6863 (N_6863,N_6725,N_6667);
or U6864 (N_6864,N_6696,N_6728);
and U6865 (N_6865,N_6653,N_6651);
nor U6866 (N_6866,N_6749,N_6677);
nand U6867 (N_6867,N_6654,N_6659);
and U6868 (N_6868,N_6626,N_6695);
nand U6869 (N_6869,N_6663,N_6678);
or U6870 (N_6870,N_6674,N_6746);
xor U6871 (N_6871,N_6673,N_6689);
nand U6872 (N_6872,N_6637,N_6693);
or U6873 (N_6873,N_6648,N_6731);
or U6874 (N_6874,N_6674,N_6732);
and U6875 (N_6875,N_6770,N_6754);
and U6876 (N_6876,N_6861,N_6813);
nand U6877 (N_6877,N_6753,N_6871);
xnor U6878 (N_6878,N_6820,N_6817);
or U6879 (N_6879,N_6818,N_6785);
nand U6880 (N_6880,N_6759,N_6869);
nor U6881 (N_6881,N_6814,N_6862);
xnor U6882 (N_6882,N_6835,N_6844);
or U6883 (N_6883,N_6865,N_6838);
nand U6884 (N_6884,N_6804,N_6842);
xor U6885 (N_6885,N_6868,N_6764);
nor U6886 (N_6886,N_6827,N_6874);
nand U6887 (N_6887,N_6858,N_6803);
nand U6888 (N_6888,N_6833,N_6758);
or U6889 (N_6889,N_6812,N_6789);
nand U6890 (N_6890,N_6853,N_6851);
or U6891 (N_6891,N_6873,N_6830);
nor U6892 (N_6892,N_6773,N_6811);
xnor U6893 (N_6893,N_6782,N_6850);
nand U6894 (N_6894,N_6778,N_6761);
or U6895 (N_6895,N_6866,N_6780);
or U6896 (N_6896,N_6756,N_6849);
nand U6897 (N_6897,N_6769,N_6774);
nand U6898 (N_6898,N_6777,N_6826);
xor U6899 (N_6899,N_6797,N_6857);
nand U6900 (N_6900,N_6808,N_6809);
nor U6901 (N_6901,N_6779,N_6757);
xnor U6902 (N_6902,N_6860,N_6791);
or U6903 (N_6903,N_6792,N_6872);
nand U6904 (N_6904,N_6767,N_6867);
and U6905 (N_6905,N_6837,N_6772);
xnor U6906 (N_6906,N_6768,N_6794);
xor U6907 (N_6907,N_6828,N_6787);
xnor U6908 (N_6908,N_6786,N_6839);
xor U6909 (N_6909,N_6840,N_6810);
or U6910 (N_6910,N_6836,N_6781);
nor U6911 (N_6911,N_6799,N_6831);
nand U6912 (N_6912,N_6806,N_6816);
nor U6913 (N_6913,N_6819,N_6790);
or U6914 (N_6914,N_6750,N_6805);
xnor U6915 (N_6915,N_6841,N_6752);
nor U6916 (N_6916,N_6775,N_6760);
nor U6917 (N_6917,N_6762,N_6795);
nand U6918 (N_6918,N_6776,N_6800);
nor U6919 (N_6919,N_6854,N_6824);
or U6920 (N_6920,N_6771,N_6823);
nand U6921 (N_6921,N_6798,N_6796);
and U6922 (N_6922,N_6834,N_6784);
nand U6923 (N_6923,N_6751,N_6793);
nand U6924 (N_6924,N_6783,N_6802);
and U6925 (N_6925,N_6807,N_6765);
xor U6926 (N_6926,N_6822,N_6848);
or U6927 (N_6927,N_6766,N_6815);
and U6928 (N_6928,N_6870,N_6788);
or U6929 (N_6929,N_6832,N_6801);
xnor U6930 (N_6930,N_6821,N_6852);
xnor U6931 (N_6931,N_6843,N_6829);
or U6932 (N_6932,N_6864,N_6845);
and U6933 (N_6933,N_6755,N_6847);
nand U6934 (N_6934,N_6863,N_6855);
xor U6935 (N_6935,N_6763,N_6846);
nor U6936 (N_6936,N_6856,N_6825);
nand U6937 (N_6937,N_6859,N_6804);
nand U6938 (N_6938,N_6863,N_6825);
or U6939 (N_6939,N_6863,N_6786);
xnor U6940 (N_6940,N_6825,N_6872);
xnor U6941 (N_6941,N_6813,N_6846);
or U6942 (N_6942,N_6798,N_6851);
nor U6943 (N_6943,N_6862,N_6846);
nor U6944 (N_6944,N_6853,N_6856);
or U6945 (N_6945,N_6865,N_6847);
or U6946 (N_6946,N_6850,N_6841);
xor U6947 (N_6947,N_6874,N_6825);
nor U6948 (N_6948,N_6843,N_6777);
and U6949 (N_6949,N_6838,N_6770);
xnor U6950 (N_6950,N_6811,N_6758);
nor U6951 (N_6951,N_6861,N_6759);
nor U6952 (N_6952,N_6751,N_6766);
or U6953 (N_6953,N_6836,N_6814);
nor U6954 (N_6954,N_6859,N_6844);
nand U6955 (N_6955,N_6776,N_6771);
nor U6956 (N_6956,N_6775,N_6786);
and U6957 (N_6957,N_6844,N_6837);
nand U6958 (N_6958,N_6800,N_6819);
nand U6959 (N_6959,N_6765,N_6849);
nand U6960 (N_6960,N_6762,N_6781);
and U6961 (N_6961,N_6799,N_6849);
nand U6962 (N_6962,N_6852,N_6873);
xnor U6963 (N_6963,N_6837,N_6806);
nand U6964 (N_6964,N_6822,N_6784);
and U6965 (N_6965,N_6853,N_6828);
nand U6966 (N_6966,N_6849,N_6805);
or U6967 (N_6967,N_6855,N_6787);
nand U6968 (N_6968,N_6775,N_6798);
and U6969 (N_6969,N_6855,N_6758);
xor U6970 (N_6970,N_6779,N_6815);
or U6971 (N_6971,N_6865,N_6794);
nand U6972 (N_6972,N_6805,N_6801);
xor U6973 (N_6973,N_6768,N_6754);
nand U6974 (N_6974,N_6776,N_6767);
xnor U6975 (N_6975,N_6834,N_6870);
xnor U6976 (N_6976,N_6766,N_6759);
nand U6977 (N_6977,N_6780,N_6863);
xnor U6978 (N_6978,N_6821,N_6801);
nand U6979 (N_6979,N_6808,N_6807);
xnor U6980 (N_6980,N_6829,N_6868);
and U6981 (N_6981,N_6866,N_6781);
and U6982 (N_6982,N_6758,N_6822);
xor U6983 (N_6983,N_6771,N_6824);
or U6984 (N_6984,N_6788,N_6854);
nor U6985 (N_6985,N_6872,N_6858);
and U6986 (N_6986,N_6752,N_6859);
nand U6987 (N_6987,N_6859,N_6819);
or U6988 (N_6988,N_6788,N_6856);
nor U6989 (N_6989,N_6775,N_6782);
or U6990 (N_6990,N_6841,N_6864);
and U6991 (N_6991,N_6765,N_6771);
or U6992 (N_6992,N_6855,N_6792);
or U6993 (N_6993,N_6750,N_6795);
or U6994 (N_6994,N_6785,N_6825);
or U6995 (N_6995,N_6761,N_6774);
nand U6996 (N_6996,N_6870,N_6847);
or U6997 (N_6997,N_6774,N_6816);
or U6998 (N_6998,N_6791,N_6770);
or U6999 (N_6999,N_6820,N_6839);
or U7000 (N_7000,N_6965,N_6921);
and U7001 (N_7001,N_6914,N_6954);
or U7002 (N_7002,N_6988,N_6953);
and U7003 (N_7003,N_6949,N_6946);
nor U7004 (N_7004,N_6892,N_6942);
nand U7005 (N_7005,N_6901,N_6906);
or U7006 (N_7006,N_6959,N_6945);
nand U7007 (N_7007,N_6919,N_6935);
nor U7008 (N_7008,N_6924,N_6966);
or U7009 (N_7009,N_6899,N_6926);
xnor U7010 (N_7010,N_6983,N_6979);
nand U7011 (N_7011,N_6950,N_6888);
nand U7012 (N_7012,N_6976,N_6894);
and U7013 (N_7013,N_6904,N_6916);
nor U7014 (N_7014,N_6877,N_6875);
and U7015 (N_7015,N_6986,N_6891);
xor U7016 (N_7016,N_6980,N_6967);
or U7017 (N_7017,N_6992,N_6882);
nor U7018 (N_7018,N_6927,N_6881);
nand U7019 (N_7019,N_6905,N_6978);
xor U7020 (N_7020,N_6896,N_6947);
or U7021 (N_7021,N_6913,N_6883);
and U7022 (N_7022,N_6981,N_6876);
nand U7023 (N_7023,N_6900,N_6895);
nand U7024 (N_7024,N_6898,N_6907);
nor U7025 (N_7025,N_6937,N_6889);
and U7026 (N_7026,N_6878,N_6893);
and U7027 (N_7027,N_6922,N_6996);
xnor U7028 (N_7028,N_6925,N_6970);
or U7029 (N_7029,N_6961,N_6991);
and U7030 (N_7030,N_6990,N_6903);
nand U7031 (N_7031,N_6912,N_6985);
xor U7032 (N_7032,N_6960,N_6884);
and U7033 (N_7033,N_6987,N_6938);
nor U7034 (N_7034,N_6930,N_6890);
or U7035 (N_7035,N_6940,N_6964);
xor U7036 (N_7036,N_6948,N_6932);
or U7037 (N_7037,N_6952,N_6972);
nand U7038 (N_7038,N_6909,N_6918);
nor U7039 (N_7039,N_6939,N_6971);
and U7040 (N_7040,N_6910,N_6880);
nand U7041 (N_7041,N_6968,N_6933);
nor U7042 (N_7042,N_6977,N_6943);
xor U7043 (N_7043,N_6944,N_6975);
xor U7044 (N_7044,N_6998,N_6958);
and U7045 (N_7045,N_6969,N_6951);
and U7046 (N_7046,N_6902,N_6897);
nand U7047 (N_7047,N_6999,N_6997);
xor U7048 (N_7048,N_6934,N_6929);
nor U7049 (N_7049,N_6920,N_6957);
and U7050 (N_7050,N_6923,N_6973);
and U7051 (N_7051,N_6887,N_6936);
or U7052 (N_7052,N_6974,N_6885);
xnor U7053 (N_7053,N_6928,N_6911);
nand U7054 (N_7054,N_6982,N_6879);
nor U7055 (N_7055,N_6931,N_6956);
and U7056 (N_7056,N_6886,N_6994);
nor U7057 (N_7057,N_6962,N_6993);
and U7058 (N_7058,N_6955,N_6941);
and U7059 (N_7059,N_6908,N_6995);
or U7060 (N_7060,N_6963,N_6989);
xnor U7061 (N_7061,N_6984,N_6915);
and U7062 (N_7062,N_6917,N_6962);
or U7063 (N_7063,N_6967,N_6894);
xnor U7064 (N_7064,N_6999,N_6973);
nand U7065 (N_7065,N_6956,N_6897);
xnor U7066 (N_7066,N_6961,N_6940);
nor U7067 (N_7067,N_6946,N_6973);
xnor U7068 (N_7068,N_6937,N_6979);
xnor U7069 (N_7069,N_6995,N_6888);
or U7070 (N_7070,N_6906,N_6923);
or U7071 (N_7071,N_6889,N_6918);
or U7072 (N_7072,N_6934,N_6876);
xnor U7073 (N_7073,N_6941,N_6890);
nand U7074 (N_7074,N_6992,N_6877);
nand U7075 (N_7075,N_6966,N_6976);
xnor U7076 (N_7076,N_6909,N_6880);
and U7077 (N_7077,N_6903,N_6922);
nor U7078 (N_7078,N_6930,N_6906);
xnor U7079 (N_7079,N_6992,N_6916);
nor U7080 (N_7080,N_6918,N_6936);
nand U7081 (N_7081,N_6875,N_6915);
xor U7082 (N_7082,N_6904,N_6923);
xnor U7083 (N_7083,N_6968,N_6972);
nand U7084 (N_7084,N_6958,N_6956);
and U7085 (N_7085,N_6886,N_6893);
or U7086 (N_7086,N_6912,N_6947);
nand U7087 (N_7087,N_6916,N_6991);
nand U7088 (N_7088,N_6939,N_6928);
or U7089 (N_7089,N_6990,N_6977);
xnor U7090 (N_7090,N_6977,N_6934);
and U7091 (N_7091,N_6985,N_6876);
and U7092 (N_7092,N_6996,N_6914);
nand U7093 (N_7093,N_6904,N_6889);
nand U7094 (N_7094,N_6993,N_6890);
and U7095 (N_7095,N_6991,N_6984);
nor U7096 (N_7096,N_6934,N_6948);
nor U7097 (N_7097,N_6913,N_6891);
and U7098 (N_7098,N_6898,N_6919);
and U7099 (N_7099,N_6957,N_6901);
xnor U7100 (N_7100,N_6887,N_6946);
nand U7101 (N_7101,N_6905,N_6917);
nor U7102 (N_7102,N_6980,N_6889);
and U7103 (N_7103,N_6922,N_6882);
and U7104 (N_7104,N_6966,N_6903);
nor U7105 (N_7105,N_6949,N_6968);
and U7106 (N_7106,N_6999,N_6948);
nand U7107 (N_7107,N_6887,N_6885);
nand U7108 (N_7108,N_6939,N_6997);
nand U7109 (N_7109,N_6944,N_6940);
nand U7110 (N_7110,N_6887,N_6918);
or U7111 (N_7111,N_6985,N_6941);
xor U7112 (N_7112,N_6948,N_6993);
or U7113 (N_7113,N_6968,N_6900);
nor U7114 (N_7114,N_6887,N_6919);
nor U7115 (N_7115,N_6951,N_6922);
nor U7116 (N_7116,N_6934,N_6919);
and U7117 (N_7117,N_6993,N_6947);
or U7118 (N_7118,N_6913,N_6892);
nand U7119 (N_7119,N_6934,N_6905);
and U7120 (N_7120,N_6892,N_6974);
nor U7121 (N_7121,N_6889,N_6930);
nor U7122 (N_7122,N_6915,N_6935);
or U7123 (N_7123,N_6962,N_6972);
xor U7124 (N_7124,N_6991,N_6924);
and U7125 (N_7125,N_7035,N_7015);
nand U7126 (N_7126,N_7012,N_7008);
or U7127 (N_7127,N_7077,N_7096);
xor U7128 (N_7128,N_7110,N_7004);
or U7129 (N_7129,N_7074,N_7034);
and U7130 (N_7130,N_7010,N_7117);
nor U7131 (N_7131,N_7018,N_7007);
or U7132 (N_7132,N_7002,N_7083);
nor U7133 (N_7133,N_7062,N_7092);
xnor U7134 (N_7134,N_7085,N_7021);
and U7135 (N_7135,N_7041,N_7044);
and U7136 (N_7136,N_7111,N_7017);
or U7137 (N_7137,N_7106,N_7121);
nor U7138 (N_7138,N_7090,N_7072);
nor U7139 (N_7139,N_7027,N_7039);
nand U7140 (N_7140,N_7102,N_7032);
nor U7141 (N_7141,N_7037,N_7000);
xnor U7142 (N_7142,N_7095,N_7038);
nand U7143 (N_7143,N_7024,N_7064);
nor U7144 (N_7144,N_7100,N_7023);
nand U7145 (N_7145,N_7116,N_7047);
nand U7146 (N_7146,N_7060,N_7001);
or U7147 (N_7147,N_7063,N_7114);
or U7148 (N_7148,N_7059,N_7099);
xnor U7149 (N_7149,N_7079,N_7011);
and U7150 (N_7150,N_7051,N_7068);
or U7151 (N_7151,N_7104,N_7086);
nand U7152 (N_7152,N_7108,N_7065);
and U7153 (N_7153,N_7013,N_7066);
xor U7154 (N_7154,N_7061,N_7054);
xnor U7155 (N_7155,N_7016,N_7115);
nor U7156 (N_7156,N_7022,N_7123);
and U7157 (N_7157,N_7025,N_7003);
nor U7158 (N_7158,N_7097,N_7030);
or U7159 (N_7159,N_7109,N_7014);
nor U7160 (N_7160,N_7120,N_7122);
and U7161 (N_7161,N_7124,N_7028);
and U7162 (N_7162,N_7081,N_7026);
and U7163 (N_7163,N_7088,N_7036);
xor U7164 (N_7164,N_7113,N_7055);
and U7165 (N_7165,N_7087,N_7050);
nor U7166 (N_7166,N_7112,N_7107);
xor U7167 (N_7167,N_7020,N_7073);
and U7168 (N_7168,N_7019,N_7029);
or U7169 (N_7169,N_7119,N_7045);
and U7170 (N_7170,N_7005,N_7084);
xnor U7171 (N_7171,N_7048,N_7049);
nand U7172 (N_7172,N_7031,N_7089);
xnor U7173 (N_7173,N_7082,N_7105);
or U7174 (N_7174,N_7103,N_7042);
and U7175 (N_7175,N_7057,N_7094);
xnor U7176 (N_7176,N_7009,N_7043);
and U7177 (N_7177,N_7056,N_7053);
or U7178 (N_7178,N_7006,N_7046);
or U7179 (N_7179,N_7091,N_7075);
and U7180 (N_7180,N_7076,N_7033);
xor U7181 (N_7181,N_7101,N_7098);
or U7182 (N_7182,N_7070,N_7080);
xor U7183 (N_7183,N_7118,N_7067);
nand U7184 (N_7184,N_7040,N_7052);
nor U7185 (N_7185,N_7071,N_7078);
nor U7186 (N_7186,N_7058,N_7093);
nor U7187 (N_7187,N_7069,N_7042);
or U7188 (N_7188,N_7041,N_7118);
xor U7189 (N_7189,N_7018,N_7014);
nor U7190 (N_7190,N_7052,N_7007);
and U7191 (N_7191,N_7005,N_7029);
nand U7192 (N_7192,N_7011,N_7063);
or U7193 (N_7193,N_7085,N_7006);
and U7194 (N_7194,N_7002,N_7000);
and U7195 (N_7195,N_7020,N_7102);
and U7196 (N_7196,N_7016,N_7073);
nand U7197 (N_7197,N_7052,N_7044);
and U7198 (N_7198,N_7094,N_7012);
xor U7199 (N_7199,N_7040,N_7109);
nand U7200 (N_7200,N_7103,N_7001);
xor U7201 (N_7201,N_7034,N_7067);
nor U7202 (N_7202,N_7113,N_7023);
xor U7203 (N_7203,N_7043,N_7025);
and U7204 (N_7204,N_7051,N_7008);
or U7205 (N_7205,N_7010,N_7106);
and U7206 (N_7206,N_7011,N_7004);
and U7207 (N_7207,N_7081,N_7019);
and U7208 (N_7208,N_7089,N_7075);
and U7209 (N_7209,N_7024,N_7077);
or U7210 (N_7210,N_7068,N_7114);
xor U7211 (N_7211,N_7010,N_7055);
or U7212 (N_7212,N_7100,N_7045);
xor U7213 (N_7213,N_7118,N_7101);
nor U7214 (N_7214,N_7065,N_7113);
xor U7215 (N_7215,N_7003,N_7120);
or U7216 (N_7216,N_7084,N_7059);
xnor U7217 (N_7217,N_7091,N_7098);
and U7218 (N_7218,N_7068,N_7072);
nand U7219 (N_7219,N_7001,N_7049);
and U7220 (N_7220,N_7124,N_7006);
xnor U7221 (N_7221,N_7115,N_7091);
and U7222 (N_7222,N_7047,N_7023);
or U7223 (N_7223,N_7059,N_7081);
nor U7224 (N_7224,N_7111,N_7104);
nand U7225 (N_7225,N_7038,N_7083);
xnor U7226 (N_7226,N_7011,N_7029);
nor U7227 (N_7227,N_7067,N_7081);
and U7228 (N_7228,N_7025,N_7115);
nor U7229 (N_7229,N_7065,N_7103);
and U7230 (N_7230,N_7120,N_7117);
or U7231 (N_7231,N_7109,N_7079);
and U7232 (N_7232,N_7026,N_7097);
or U7233 (N_7233,N_7068,N_7115);
and U7234 (N_7234,N_7101,N_7108);
xor U7235 (N_7235,N_7087,N_7082);
or U7236 (N_7236,N_7025,N_7104);
or U7237 (N_7237,N_7117,N_7105);
and U7238 (N_7238,N_7115,N_7107);
nand U7239 (N_7239,N_7116,N_7050);
nor U7240 (N_7240,N_7033,N_7089);
nor U7241 (N_7241,N_7053,N_7019);
nand U7242 (N_7242,N_7062,N_7001);
and U7243 (N_7243,N_7109,N_7113);
nor U7244 (N_7244,N_7112,N_7095);
nand U7245 (N_7245,N_7027,N_7124);
nor U7246 (N_7246,N_7071,N_7052);
and U7247 (N_7247,N_7080,N_7037);
xnor U7248 (N_7248,N_7009,N_7008);
or U7249 (N_7249,N_7052,N_7117);
xnor U7250 (N_7250,N_7189,N_7149);
nand U7251 (N_7251,N_7231,N_7223);
and U7252 (N_7252,N_7220,N_7199);
nor U7253 (N_7253,N_7136,N_7215);
xor U7254 (N_7254,N_7138,N_7132);
or U7255 (N_7255,N_7217,N_7178);
nand U7256 (N_7256,N_7222,N_7248);
and U7257 (N_7257,N_7202,N_7137);
nor U7258 (N_7258,N_7171,N_7183);
nand U7259 (N_7259,N_7161,N_7157);
and U7260 (N_7260,N_7131,N_7224);
xor U7261 (N_7261,N_7181,N_7249);
xnor U7262 (N_7262,N_7143,N_7206);
or U7263 (N_7263,N_7144,N_7160);
and U7264 (N_7264,N_7150,N_7221);
or U7265 (N_7265,N_7201,N_7169);
nor U7266 (N_7266,N_7162,N_7147);
and U7267 (N_7267,N_7246,N_7165);
nand U7268 (N_7268,N_7173,N_7126);
nor U7269 (N_7269,N_7164,N_7242);
xor U7270 (N_7270,N_7129,N_7226);
and U7271 (N_7271,N_7210,N_7205);
or U7272 (N_7272,N_7140,N_7172);
xor U7273 (N_7273,N_7167,N_7185);
and U7274 (N_7274,N_7233,N_7125);
xor U7275 (N_7275,N_7247,N_7241);
xor U7276 (N_7276,N_7151,N_7158);
xor U7277 (N_7277,N_7135,N_7176);
or U7278 (N_7278,N_7200,N_7163);
xor U7279 (N_7279,N_7211,N_7148);
nor U7280 (N_7280,N_7182,N_7196);
or U7281 (N_7281,N_7237,N_7190);
xor U7282 (N_7282,N_7203,N_7216);
xnor U7283 (N_7283,N_7180,N_7228);
nor U7284 (N_7284,N_7187,N_7193);
nand U7285 (N_7285,N_7128,N_7235);
xor U7286 (N_7286,N_7184,N_7168);
or U7287 (N_7287,N_7186,N_7154);
or U7288 (N_7288,N_7127,N_7139);
nor U7289 (N_7289,N_7153,N_7207);
nand U7290 (N_7290,N_7227,N_7243);
or U7291 (N_7291,N_7239,N_7159);
or U7292 (N_7292,N_7232,N_7230);
xor U7293 (N_7293,N_7240,N_7234);
nor U7294 (N_7294,N_7197,N_7225);
nand U7295 (N_7295,N_7245,N_7170);
nand U7296 (N_7296,N_7188,N_7194);
nor U7297 (N_7297,N_7156,N_7195);
nand U7298 (N_7298,N_7166,N_7177);
nor U7299 (N_7299,N_7229,N_7134);
or U7300 (N_7300,N_7133,N_7192);
nand U7301 (N_7301,N_7208,N_7209);
and U7302 (N_7302,N_7236,N_7238);
or U7303 (N_7303,N_7155,N_7152);
nand U7304 (N_7304,N_7244,N_7146);
nor U7305 (N_7305,N_7218,N_7212);
nand U7306 (N_7306,N_7130,N_7145);
nor U7307 (N_7307,N_7191,N_7179);
and U7308 (N_7308,N_7175,N_7141);
nand U7309 (N_7309,N_7214,N_7219);
or U7310 (N_7310,N_7142,N_7204);
nand U7311 (N_7311,N_7174,N_7198);
xnor U7312 (N_7312,N_7213,N_7246);
nor U7313 (N_7313,N_7208,N_7142);
nand U7314 (N_7314,N_7223,N_7136);
xnor U7315 (N_7315,N_7188,N_7149);
nand U7316 (N_7316,N_7157,N_7171);
nand U7317 (N_7317,N_7221,N_7177);
xor U7318 (N_7318,N_7189,N_7228);
nor U7319 (N_7319,N_7219,N_7179);
xor U7320 (N_7320,N_7183,N_7182);
nor U7321 (N_7321,N_7211,N_7230);
xor U7322 (N_7322,N_7204,N_7165);
xor U7323 (N_7323,N_7126,N_7182);
xor U7324 (N_7324,N_7199,N_7146);
nor U7325 (N_7325,N_7197,N_7139);
and U7326 (N_7326,N_7149,N_7175);
nand U7327 (N_7327,N_7224,N_7229);
xor U7328 (N_7328,N_7159,N_7181);
nand U7329 (N_7329,N_7133,N_7130);
xnor U7330 (N_7330,N_7172,N_7181);
nand U7331 (N_7331,N_7230,N_7169);
xnor U7332 (N_7332,N_7149,N_7132);
and U7333 (N_7333,N_7191,N_7149);
nor U7334 (N_7334,N_7211,N_7141);
and U7335 (N_7335,N_7234,N_7127);
nor U7336 (N_7336,N_7153,N_7200);
or U7337 (N_7337,N_7208,N_7225);
xor U7338 (N_7338,N_7218,N_7162);
nor U7339 (N_7339,N_7194,N_7161);
nand U7340 (N_7340,N_7204,N_7202);
or U7341 (N_7341,N_7128,N_7173);
nor U7342 (N_7342,N_7228,N_7147);
and U7343 (N_7343,N_7220,N_7229);
xor U7344 (N_7344,N_7133,N_7163);
and U7345 (N_7345,N_7222,N_7134);
nor U7346 (N_7346,N_7236,N_7134);
or U7347 (N_7347,N_7138,N_7209);
or U7348 (N_7348,N_7157,N_7193);
and U7349 (N_7349,N_7200,N_7201);
nor U7350 (N_7350,N_7206,N_7162);
and U7351 (N_7351,N_7198,N_7136);
or U7352 (N_7352,N_7130,N_7134);
nand U7353 (N_7353,N_7165,N_7223);
and U7354 (N_7354,N_7228,N_7187);
xnor U7355 (N_7355,N_7164,N_7170);
and U7356 (N_7356,N_7176,N_7177);
xnor U7357 (N_7357,N_7155,N_7158);
xor U7358 (N_7358,N_7198,N_7152);
xor U7359 (N_7359,N_7145,N_7227);
nor U7360 (N_7360,N_7210,N_7140);
or U7361 (N_7361,N_7241,N_7193);
nor U7362 (N_7362,N_7236,N_7175);
nand U7363 (N_7363,N_7176,N_7148);
nand U7364 (N_7364,N_7141,N_7178);
and U7365 (N_7365,N_7132,N_7206);
and U7366 (N_7366,N_7190,N_7186);
and U7367 (N_7367,N_7237,N_7136);
xnor U7368 (N_7368,N_7224,N_7194);
and U7369 (N_7369,N_7220,N_7148);
xnor U7370 (N_7370,N_7185,N_7179);
nor U7371 (N_7371,N_7208,N_7137);
nand U7372 (N_7372,N_7157,N_7207);
nand U7373 (N_7373,N_7207,N_7208);
nand U7374 (N_7374,N_7235,N_7206);
xor U7375 (N_7375,N_7301,N_7328);
or U7376 (N_7376,N_7300,N_7314);
xor U7377 (N_7377,N_7315,N_7275);
or U7378 (N_7378,N_7304,N_7320);
or U7379 (N_7379,N_7346,N_7252);
or U7380 (N_7380,N_7279,N_7265);
and U7381 (N_7381,N_7339,N_7319);
nand U7382 (N_7382,N_7312,N_7307);
xnor U7383 (N_7383,N_7283,N_7311);
or U7384 (N_7384,N_7355,N_7363);
or U7385 (N_7385,N_7353,N_7257);
nor U7386 (N_7386,N_7282,N_7250);
or U7387 (N_7387,N_7256,N_7270);
xor U7388 (N_7388,N_7286,N_7288);
nor U7389 (N_7389,N_7362,N_7368);
nand U7390 (N_7390,N_7369,N_7268);
and U7391 (N_7391,N_7318,N_7266);
nor U7392 (N_7392,N_7297,N_7326);
nor U7393 (N_7393,N_7287,N_7277);
xor U7394 (N_7394,N_7367,N_7334);
or U7395 (N_7395,N_7251,N_7267);
xnor U7396 (N_7396,N_7335,N_7309);
xor U7397 (N_7397,N_7269,N_7351);
or U7398 (N_7398,N_7329,N_7263);
xnor U7399 (N_7399,N_7313,N_7338);
xor U7400 (N_7400,N_7281,N_7273);
nand U7401 (N_7401,N_7254,N_7271);
nor U7402 (N_7402,N_7325,N_7373);
or U7403 (N_7403,N_7323,N_7259);
or U7404 (N_7404,N_7340,N_7343);
nand U7405 (N_7405,N_7295,N_7274);
nand U7406 (N_7406,N_7280,N_7276);
or U7407 (N_7407,N_7321,N_7258);
and U7408 (N_7408,N_7345,N_7357);
and U7409 (N_7409,N_7324,N_7347);
or U7410 (N_7410,N_7365,N_7302);
nor U7411 (N_7411,N_7356,N_7289);
and U7412 (N_7412,N_7296,N_7371);
nand U7413 (N_7413,N_7360,N_7308);
nor U7414 (N_7414,N_7291,N_7361);
xnor U7415 (N_7415,N_7278,N_7253);
xor U7416 (N_7416,N_7372,N_7262);
or U7417 (N_7417,N_7348,N_7290);
or U7418 (N_7418,N_7298,N_7294);
xor U7419 (N_7419,N_7370,N_7330);
or U7420 (N_7420,N_7264,N_7285);
xor U7421 (N_7421,N_7331,N_7332);
nand U7422 (N_7422,N_7284,N_7342);
nor U7423 (N_7423,N_7293,N_7352);
nand U7424 (N_7424,N_7366,N_7354);
and U7425 (N_7425,N_7303,N_7327);
nor U7426 (N_7426,N_7322,N_7349);
nand U7427 (N_7427,N_7350,N_7305);
nor U7428 (N_7428,N_7374,N_7341);
nor U7429 (N_7429,N_7358,N_7364);
nor U7430 (N_7430,N_7336,N_7316);
and U7431 (N_7431,N_7260,N_7306);
nor U7432 (N_7432,N_7255,N_7310);
xnor U7433 (N_7433,N_7292,N_7261);
nor U7434 (N_7434,N_7299,N_7272);
and U7435 (N_7435,N_7359,N_7317);
or U7436 (N_7436,N_7333,N_7344);
and U7437 (N_7437,N_7337,N_7366);
nor U7438 (N_7438,N_7336,N_7353);
nand U7439 (N_7439,N_7363,N_7272);
or U7440 (N_7440,N_7360,N_7305);
xnor U7441 (N_7441,N_7280,N_7277);
and U7442 (N_7442,N_7353,N_7314);
or U7443 (N_7443,N_7304,N_7335);
or U7444 (N_7444,N_7251,N_7353);
and U7445 (N_7445,N_7356,N_7373);
and U7446 (N_7446,N_7270,N_7290);
nor U7447 (N_7447,N_7251,N_7292);
and U7448 (N_7448,N_7279,N_7303);
or U7449 (N_7449,N_7332,N_7359);
or U7450 (N_7450,N_7311,N_7341);
nor U7451 (N_7451,N_7368,N_7364);
or U7452 (N_7452,N_7290,N_7343);
nor U7453 (N_7453,N_7351,N_7309);
and U7454 (N_7454,N_7314,N_7275);
xnor U7455 (N_7455,N_7308,N_7276);
nand U7456 (N_7456,N_7292,N_7316);
nand U7457 (N_7457,N_7321,N_7269);
or U7458 (N_7458,N_7264,N_7354);
xnor U7459 (N_7459,N_7343,N_7307);
xnor U7460 (N_7460,N_7372,N_7305);
nand U7461 (N_7461,N_7254,N_7256);
and U7462 (N_7462,N_7340,N_7365);
nor U7463 (N_7463,N_7345,N_7289);
or U7464 (N_7464,N_7355,N_7273);
nand U7465 (N_7465,N_7360,N_7279);
nand U7466 (N_7466,N_7306,N_7374);
nand U7467 (N_7467,N_7320,N_7366);
nand U7468 (N_7468,N_7329,N_7256);
or U7469 (N_7469,N_7319,N_7311);
nor U7470 (N_7470,N_7327,N_7333);
nand U7471 (N_7471,N_7325,N_7292);
and U7472 (N_7472,N_7287,N_7364);
or U7473 (N_7473,N_7373,N_7341);
nor U7474 (N_7474,N_7358,N_7374);
xnor U7475 (N_7475,N_7250,N_7370);
xor U7476 (N_7476,N_7329,N_7367);
xor U7477 (N_7477,N_7369,N_7302);
xor U7478 (N_7478,N_7300,N_7365);
xnor U7479 (N_7479,N_7302,N_7353);
nand U7480 (N_7480,N_7341,N_7267);
or U7481 (N_7481,N_7258,N_7266);
nor U7482 (N_7482,N_7313,N_7286);
and U7483 (N_7483,N_7289,N_7299);
or U7484 (N_7484,N_7252,N_7313);
or U7485 (N_7485,N_7364,N_7317);
and U7486 (N_7486,N_7253,N_7277);
nor U7487 (N_7487,N_7342,N_7334);
xnor U7488 (N_7488,N_7259,N_7346);
or U7489 (N_7489,N_7293,N_7280);
xor U7490 (N_7490,N_7296,N_7323);
or U7491 (N_7491,N_7282,N_7374);
or U7492 (N_7492,N_7328,N_7322);
xnor U7493 (N_7493,N_7335,N_7331);
and U7494 (N_7494,N_7324,N_7372);
and U7495 (N_7495,N_7283,N_7355);
or U7496 (N_7496,N_7313,N_7324);
nand U7497 (N_7497,N_7337,N_7355);
nand U7498 (N_7498,N_7370,N_7308);
or U7499 (N_7499,N_7348,N_7359);
nor U7500 (N_7500,N_7416,N_7447);
and U7501 (N_7501,N_7392,N_7445);
and U7502 (N_7502,N_7443,N_7440);
xnor U7503 (N_7503,N_7451,N_7432);
xor U7504 (N_7504,N_7397,N_7485);
or U7505 (N_7505,N_7466,N_7479);
nand U7506 (N_7506,N_7458,N_7461);
nor U7507 (N_7507,N_7477,N_7469);
or U7508 (N_7508,N_7395,N_7384);
and U7509 (N_7509,N_7473,N_7476);
or U7510 (N_7510,N_7424,N_7483);
xnor U7511 (N_7511,N_7462,N_7460);
and U7512 (N_7512,N_7378,N_7436);
and U7513 (N_7513,N_7421,N_7399);
or U7514 (N_7514,N_7382,N_7389);
nor U7515 (N_7515,N_7412,N_7454);
or U7516 (N_7516,N_7413,N_7449);
or U7517 (N_7517,N_7381,N_7426);
or U7518 (N_7518,N_7434,N_7448);
nor U7519 (N_7519,N_7401,N_7415);
or U7520 (N_7520,N_7396,N_7463);
nand U7521 (N_7521,N_7410,N_7379);
nand U7522 (N_7522,N_7422,N_7380);
xnor U7523 (N_7523,N_7430,N_7474);
and U7524 (N_7524,N_7388,N_7488);
xnor U7525 (N_7525,N_7452,N_7482);
or U7526 (N_7526,N_7375,N_7438);
and U7527 (N_7527,N_7475,N_7453);
xor U7528 (N_7528,N_7492,N_7394);
and U7529 (N_7529,N_7457,N_7446);
xnor U7530 (N_7530,N_7468,N_7499);
xor U7531 (N_7531,N_7387,N_7402);
xnor U7532 (N_7532,N_7406,N_7393);
nand U7533 (N_7533,N_7472,N_7433);
nor U7534 (N_7534,N_7464,N_7411);
nand U7535 (N_7535,N_7450,N_7465);
nor U7536 (N_7536,N_7481,N_7431);
nand U7537 (N_7537,N_7437,N_7405);
nor U7538 (N_7538,N_7385,N_7398);
or U7539 (N_7539,N_7497,N_7442);
nor U7540 (N_7540,N_7489,N_7456);
nor U7541 (N_7541,N_7498,N_7383);
and U7542 (N_7542,N_7403,N_7390);
nand U7543 (N_7543,N_7471,N_7386);
xor U7544 (N_7544,N_7377,N_7417);
xor U7545 (N_7545,N_7487,N_7409);
xnor U7546 (N_7546,N_7376,N_7441);
nand U7547 (N_7547,N_7478,N_7429);
or U7548 (N_7548,N_7455,N_7420);
nand U7549 (N_7549,N_7414,N_7491);
and U7550 (N_7550,N_7435,N_7391);
and U7551 (N_7551,N_7480,N_7407);
nand U7552 (N_7552,N_7495,N_7444);
nand U7553 (N_7553,N_7459,N_7484);
nor U7554 (N_7554,N_7467,N_7419);
xor U7555 (N_7555,N_7494,N_7408);
and U7556 (N_7556,N_7400,N_7470);
nand U7557 (N_7557,N_7486,N_7423);
or U7558 (N_7558,N_7490,N_7427);
nor U7559 (N_7559,N_7496,N_7418);
nand U7560 (N_7560,N_7425,N_7404);
or U7561 (N_7561,N_7439,N_7428);
or U7562 (N_7562,N_7493,N_7410);
or U7563 (N_7563,N_7462,N_7491);
and U7564 (N_7564,N_7390,N_7436);
nand U7565 (N_7565,N_7470,N_7479);
or U7566 (N_7566,N_7392,N_7409);
nand U7567 (N_7567,N_7416,N_7391);
xor U7568 (N_7568,N_7404,N_7499);
nand U7569 (N_7569,N_7446,N_7377);
nand U7570 (N_7570,N_7484,N_7395);
nand U7571 (N_7571,N_7388,N_7442);
or U7572 (N_7572,N_7383,N_7478);
or U7573 (N_7573,N_7377,N_7414);
xor U7574 (N_7574,N_7400,N_7399);
nor U7575 (N_7575,N_7479,N_7486);
nor U7576 (N_7576,N_7392,N_7468);
or U7577 (N_7577,N_7387,N_7397);
and U7578 (N_7578,N_7403,N_7435);
xnor U7579 (N_7579,N_7405,N_7377);
xor U7580 (N_7580,N_7446,N_7416);
nand U7581 (N_7581,N_7455,N_7473);
nand U7582 (N_7582,N_7458,N_7434);
xor U7583 (N_7583,N_7430,N_7487);
or U7584 (N_7584,N_7487,N_7402);
nand U7585 (N_7585,N_7392,N_7396);
nor U7586 (N_7586,N_7421,N_7396);
nor U7587 (N_7587,N_7488,N_7456);
nand U7588 (N_7588,N_7445,N_7375);
xnor U7589 (N_7589,N_7483,N_7452);
or U7590 (N_7590,N_7384,N_7460);
xor U7591 (N_7591,N_7385,N_7441);
or U7592 (N_7592,N_7465,N_7426);
or U7593 (N_7593,N_7491,N_7486);
xor U7594 (N_7594,N_7386,N_7389);
and U7595 (N_7595,N_7472,N_7496);
xnor U7596 (N_7596,N_7484,N_7381);
nor U7597 (N_7597,N_7425,N_7471);
and U7598 (N_7598,N_7474,N_7455);
nor U7599 (N_7599,N_7492,N_7448);
nor U7600 (N_7600,N_7482,N_7405);
and U7601 (N_7601,N_7410,N_7395);
or U7602 (N_7602,N_7434,N_7393);
nand U7603 (N_7603,N_7403,N_7432);
and U7604 (N_7604,N_7487,N_7390);
xor U7605 (N_7605,N_7452,N_7406);
nand U7606 (N_7606,N_7432,N_7443);
or U7607 (N_7607,N_7478,N_7406);
and U7608 (N_7608,N_7485,N_7434);
or U7609 (N_7609,N_7474,N_7426);
xnor U7610 (N_7610,N_7404,N_7485);
and U7611 (N_7611,N_7493,N_7401);
or U7612 (N_7612,N_7440,N_7492);
and U7613 (N_7613,N_7464,N_7487);
nand U7614 (N_7614,N_7466,N_7399);
nand U7615 (N_7615,N_7395,N_7425);
nor U7616 (N_7616,N_7388,N_7493);
nand U7617 (N_7617,N_7467,N_7499);
nor U7618 (N_7618,N_7382,N_7393);
and U7619 (N_7619,N_7417,N_7418);
xor U7620 (N_7620,N_7386,N_7459);
or U7621 (N_7621,N_7384,N_7378);
xor U7622 (N_7622,N_7438,N_7465);
and U7623 (N_7623,N_7414,N_7473);
nor U7624 (N_7624,N_7430,N_7409);
nor U7625 (N_7625,N_7606,N_7603);
nor U7626 (N_7626,N_7564,N_7543);
or U7627 (N_7627,N_7541,N_7620);
nor U7628 (N_7628,N_7598,N_7624);
and U7629 (N_7629,N_7547,N_7526);
and U7630 (N_7630,N_7568,N_7514);
nand U7631 (N_7631,N_7559,N_7531);
nor U7632 (N_7632,N_7506,N_7509);
xor U7633 (N_7633,N_7503,N_7551);
nor U7634 (N_7634,N_7540,N_7530);
xnor U7635 (N_7635,N_7544,N_7621);
xnor U7636 (N_7636,N_7604,N_7574);
or U7637 (N_7637,N_7539,N_7508);
or U7638 (N_7638,N_7583,N_7532);
or U7639 (N_7639,N_7584,N_7556);
nand U7640 (N_7640,N_7591,N_7554);
or U7641 (N_7641,N_7533,N_7571);
and U7642 (N_7642,N_7513,N_7579);
or U7643 (N_7643,N_7572,N_7505);
and U7644 (N_7644,N_7596,N_7610);
nor U7645 (N_7645,N_7565,N_7600);
or U7646 (N_7646,N_7537,N_7507);
or U7647 (N_7647,N_7511,N_7608);
nor U7648 (N_7648,N_7553,N_7504);
nand U7649 (N_7649,N_7599,N_7535);
nand U7650 (N_7650,N_7536,N_7573);
or U7651 (N_7651,N_7592,N_7561);
nor U7652 (N_7652,N_7575,N_7521);
xor U7653 (N_7653,N_7609,N_7619);
nand U7654 (N_7654,N_7585,N_7570);
and U7655 (N_7655,N_7548,N_7607);
xnor U7656 (N_7656,N_7522,N_7560);
and U7657 (N_7657,N_7613,N_7557);
or U7658 (N_7658,N_7520,N_7594);
xnor U7659 (N_7659,N_7588,N_7510);
or U7660 (N_7660,N_7595,N_7529);
nand U7661 (N_7661,N_7517,N_7616);
xor U7662 (N_7662,N_7549,N_7623);
or U7663 (N_7663,N_7545,N_7538);
and U7664 (N_7664,N_7500,N_7581);
and U7665 (N_7665,N_7558,N_7525);
or U7666 (N_7666,N_7587,N_7612);
nand U7667 (N_7667,N_7542,N_7550);
and U7668 (N_7668,N_7569,N_7515);
nand U7669 (N_7669,N_7580,N_7589);
and U7670 (N_7670,N_7502,N_7501);
nor U7671 (N_7671,N_7578,N_7524);
xor U7672 (N_7672,N_7622,N_7512);
and U7673 (N_7673,N_7618,N_7601);
or U7674 (N_7674,N_7615,N_7555);
and U7675 (N_7675,N_7617,N_7562);
nand U7676 (N_7676,N_7614,N_7577);
and U7677 (N_7677,N_7523,N_7518);
or U7678 (N_7678,N_7546,N_7528);
nand U7679 (N_7679,N_7563,N_7567);
nand U7680 (N_7680,N_7527,N_7534);
or U7681 (N_7681,N_7552,N_7516);
and U7682 (N_7682,N_7519,N_7593);
xor U7683 (N_7683,N_7602,N_7586);
or U7684 (N_7684,N_7582,N_7605);
nand U7685 (N_7685,N_7566,N_7576);
or U7686 (N_7686,N_7597,N_7611);
xnor U7687 (N_7687,N_7590,N_7523);
or U7688 (N_7688,N_7604,N_7619);
nand U7689 (N_7689,N_7502,N_7564);
xor U7690 (N_7690,N_7605,N_7559);
or U7691 (N_7691,N_7534,N_7604);
xor U7692 (N_7692,N_7529,N_7508);
nor U7693 (N_7693,N_7577,N_7542);
and U7694 (N_7694,N_7579,N_7559);
and U7695 (N_7695,N_7570,N_7572);
or U7696 (N_7696,N_7590,N_7592);
nand U7697 (N_7697,N_7558,N_7566);
nor U7698 (N_7698,N_7584,N_7621);
and U7699 (N_7699,N_7521,N_7560);
or U7700 (N_7700,N_7531,N_7538);
and U7701 (N_7701,N_7559,N_7530);
xnor U7702 (N_7702,N_7526,N_7619);
or U7703 (N_7703,N_7597,N_7574);
xor U7704 (N_7704,N_7552,N_7610);
or U7705 (N_7705,N_7533,N_7538);
nor U7706 (N_7706,N_7569,N_7542);
and U7707 (N_7707,N_7549,N_7541);
or U7708 (N_7708,N_7585,N_7567);
and U7709 (N_7709,N_7610,N_7572);
nand U7710 (N_7710,N_7522,N_7563);
and U7711 (N_7711,N_7504,N_7608);
xor U7712 (N_7712,N_7598,N_7608);
nor U7713 (N_7713,N_7533,N_7606);
and U7714 (N_7714,N_7572,N_7554);
xnor U7715 (N_7715,N_7587,N_7575);
nor U7716 (N_7716,N_7509,N_7571);
nand U7717 (N_7717,N_7504,N_7622);
or U7718 (N_7718,N_7598,N_7603);
nor U7719 (N_7719,N_7511,N_7508);
and U7720 (N_7720,N_7561,N_7597);
nor U7721 (N_7721,N_7588,N_7521);
xnor U7722 (N_7722,N_7517,N_7614);
xnor U7723 (N_7723,N_7531,N_7624);
nor U7724 (N_7724,N_7589,N_7610);
nor U7725 (N_7725,N_7608,N_7565);
nor U7726 (N_7726,N_7532,N_7563);
nand U7727 (N_7727,N_7562,N_7594);
nand U7728 (N_7728,N_7592,N_7572);
or U7729 (N_7729,N_7572,N_7593);
or U7730 (N_7730,N_7538,N_7601);
or U7731 (N_7731,N_7503,N_7579);
or U7732 (N_7732,N_7513,N_7599);
nor U7733 (N_7733,N_7586,N_7507);
xnor U7734 (N_7734,N_7576,N_7549);
or U7735 (N_7735,N_7508,N_7515);
and U7736 (N_7736,N_7519,N_7532);
xor U7737 (N_7737,N_7506,N_7535);
nor U7738 (N_7738,N_7585,N_7532);
nor U7739 (N_7739,N_7568,N_7619);
nor U7740 (N_7740,N_7612,N_7601);
xnor U7741 (N_7741,N_7515,N_7555);
or U7742 (N_7742,N_7524,N_7534);
nand U7743 (N_7743,N_7583,N_7543);
or U7744 (N_7744,N_7571,N_7609);
nand U7745 (N_7745,N_7606,N_7602);
or U7746 (N_7746,N_7585,N_7515);
and U7747 (N_7747,N_7506,N_7515);
or U7748 (N_7748,N_7530,N_7618);
or U7749 (N_7749,N_7614,N_7520);
nand U7750 (N_7750,N_7740,N_7666);
xor U7751 (N_7751,N_7744,N_7697);
and U7752 (N_7752,N_7689,N_7626);
nor U7753 (N_7753,N_7717,N_7728);
nand U7754 (N_7754,N_7673,N_7655);
nor U7755 (N_7755,N_7690,N_7631);
or U7756 (N_7756,N_7683,N_7727);
or U7757 (N_7757,N_7661,N_7639);
or U7758 (N_7758,N_7701,N_7732);
nand U7759 (N_7759,N_7694,N_7720);
or U7760 (N_7760,N_7675,N_7714);
nor U7761 (N_7761,N_7660,N_7638);
and U7762 (N_7762,N_7721,N_7633);
nand U7763 (N_7763,N_7684,N_7678);
and U7764 (N_7764,N_7676,N_7748);
nand U7765 (N_7765,N_7708,N_7702);
nand U7766 (N_7766,N_7698,N_7693);
and U7767 (N_7767,N_7667,N_7632);
nor U7768 (N_7768,N_7656,N_7709);
or U7769 (N_7769,N_7649,N_7723);
xnor U7770 (N_7770,N_7718,N_7731);
nand U7771 (N_7771,N_7733,N_7674);
or U7772 (N_7772,N_7695,N_7687);
and U7773 (N_7773,N_7700,N_7692);
xnor U7774 (N_7774,N_7634,N_7625);
and U7775 (N_7775,N_7654,N_7637);
nor U7776 (N_7776,N_7651,N_7657);
xor U7777 (N_7777,N_7664,N_7688);
nand U7778 (N_7778,N_7652,N_7743);
nor U7779 (N_7779,N_7668,N_7627);
nor U7780 (N_7780,N_7713,N_7705);
or U7781 (N_7781,N_7716,N_7648);
or U7782 (N_7782,N_7707,N_7682);
and U7783 (N_7783,N_7730,N_7669);
nand U7784 (N_7784,N_7738,N_7671);
xnor U7785 (N_7785,N_7628,N_7665);
nand U7786 (N_7786,N_7724,N_7642);
and U7787 (N_7787,N_7715,N_7711);
xor U7788 (N_7788,N_7712,N_7629);
nor U7789 (N_7789,N_7706,N_7736);
nor U7790 (N_7790,N_7734,N_7726);
and U7791 (N_7791,N_7686,N_7749);
nor U7792 (N_7792,N_7737,N_7662);
and U7793 (N_7793,N_7635,N_7640);
and U7794 (N_7794,N_7650,N_7685);
and U7795 (N_7795,N_7645,N_7653);
and U7796 (N_7796,N_7710,N_7670);
nor U7797 (N_7797,N_7725,N_7672);
or U7798 (N_7798,N_7691,N_7746);
and U7799 (N_7799,N_7735,N_7742);
xnor U7800 (N_7800,N_7630,N_7696);
xnor U7801 (N_7801,N_7704,N_7646);
nor U7802 (N_7802,N_7703,N_7719);
and U7803 (N_7803,N_7636,N_7680);
and U7804 (N_7804,N_7722,N_7643);
and U7805 (N_7805,N_7659,N_7739);
xor U7806 (N_7806,N_7745,N_7741);
nor U7807 (N_7807,N_7681,N_7677);
or U7808 (N_7808,N_7663,N_7641);
xnor U7809 (N_7809,N_7679,N_7699);
or U7810 (N_7810,N_7647,N_7658);
or U7811 (N_7811,N_7644,N_7729);
or U7812 (N_7812,N_7747,N_7671);
or U7813 (N_7813,N_7634,N_7684);
xnor U7814 (N_7814,N_7696,N_7721);
and U7815 (N_7815,N_7667,N_7625);
xnor U7816 (N_7816,N_7730,N_7625);
or U7817 (N_7817,N_7727,N_7675);
nor U7818 (N_7818,N_7641,N_7648);
and U7819 (N_7819,N_7696,N_7738);
nand U7820 (N_7820,N_7694,N_7663);
or U7821 (N_7821,N_7725,N_7671);
xor U7822 (N_7822,N_7745,N_7744);
and U7823 (N_7823,N_7672,N_7671);
or U7824 (N_7824,N_7630,N_7674);
nand U7825 (N_7825,N_7723,N_7674);
nor U7826 (N_7826,N_7733,N_7711);
nand U7827 (N_7827,N_7737,N_7646);
xor U7828 (N_7828,N_7629,N_7714);
nand U7829 (N_7829,N_7709,N_7666);
nor U7830 (N_7830,N_7633,N_7737);
xnor U7831 (N_7831,N_7719,N_7644);
xor U7832 (N_7832,N_7693,N_7688);
and U7833 (N_7833,N_7679,N_7717);
or U7834 (N_7834,N_7725,N_7636);
and U7835 (N_7835,N_7707,N_7714);
xnor U7836 (N_7836,N_7719,N_7681);
and U7837 (N_7837,N_7638,N_7695);
or U7838 (N_7838,N_7680,N_7714);
xor U7839 (N_7839,N_7630,N_7704);
nor U7840 (N_7840,N_7715,N_7646);
and U7841 (N_7841,N_7705,N_7733);
and U7842 (N_7842,N_7637,N_7743);
nor U7843 (N_7843,N_7692,N_7645);
nor U7844 (N_7844,N_7667,N_7720);
and U7845 (N_7845,N_7673,N_7748);
nand U7846 (N_7846,N_7631,N_7625);
xor U7847 (N_7847,N_7653,N_7643);
or U7848 (N_7848,N_7629,N_7641);
xnor U7849 (N_7849,N_7696,N_7715);
nor U7850 (N_7850,N_7666,N_7700);
or U7851 (N_7851,N_7687,N_7696);
xnor U7852 (N_7852,N_7733,N_7640);
or U7853 (N_7853,N_7647,N_7724);
xnor U7854 (N_7854,N_7723,N_7647);
nor U7855 (N_7855,N_7648,N_7636);
nor U7856 (N_7856,N_7667,N_7703);
or U7857 (N_7857,N_7739,N_7660);
nor U7858 (N_7858,N_7686,N_7747);
nor U7859 (N_7859,N_7688,N_7726);
or U7860 (N_7860,N_7670,N_7744);
and U7861 (N_7861,N_7702,N_7677);
or U7862 (N_7862,N_7699,N_7747);
or U7863 (N_7863,N_7667,N_7653);
nor U7864 (N_7864,N_7680,N_7728);
nor U7865 (N_7865,N_7653,N_7671);
nor U7866 (N_7866,N_7668,N_7667);
and U7867 (N_7867,N_7674,N_7680);
and U7868 (N_7868,N_7739,N_7633);
xor U7869 (N_7869,N_7641,N_7732);
nor U7870 (N_7870,N_7637,N_7698);
nand U7871 (N_7871,N_7653,N_7669);
xnor U7872 (N_7872,N_7747,N_7654);
xnor U7873 (N_7873,N_7632,N_7727);
nor U7874 (N_7874,N_7719,N_7729);
xnor U7875 (N_7875,N_7858,N_7782);
xnor U7876 (N_7876,N_7857,N_7752);
or U7877 (N_7877,N_7814,N_7812);
nor U7878 (N_7878,N_7789,N_7781);
nand U7879 (N_7879,N_7855,N_7830);
xnor U7880 (N_7880,N_7848,N_7768);
nand U7881 (N_7881,N_7784,N_7839);
or U7882 (N_7882,N_7793,N_7755);
nand U7883 (N_7883,N_7798,N_7777);
nor U7884 (N_7884,N_7824,N_7758);
nor U7885 (N_7885,N_7811,N_7813);
nand U7886 (N_7886,N_7849,N_7874);
xor U7887 (N_7887,N_7827,N_7820);
nand U7888 (N_7888,N_7836,N_7826);
nor U7889 (N_7889,N_7818,N_7791);
and U7890 (N_7890,N_7764,N_7823);
nand U7891 (N_7891,N_7834,N_7801);
and U7892 (N_7892,N_7799,N_7804);
or U7893 (N_7893,N_7792,N_7800);
nor U7894 (N_7894,N_7845,N_7772);
and U7895 (N_7895,N_7775,N_7867);
or U7896 (N_7896,N_7866,N_7754);
and U7897 (N_7897,N_7817,N_7847);
xnor U7898 (N_7898,N_7795,N_7788);
or U7899 (N_7899,N_7842,N_7751);
or U7900 (N_7900,N_7770,N_7802);
and U7901 (N_7901,N_7825,N_7864);
nand U7902 (N_7902,N_7861,N_7816);
nor U7903 (N_7903,N_7872,N_7821);
and U7904 (N_7904,N_7765,N_7769);
nor U7905 (N_7905,N_7794,N_7869);
or U7906 (N_7906,N_7837,N_7860);
nor U7907 (N_7907,N_7806,N_7865);
or U7908 (N_7908,N_7829,N_7862);
xor U7909 (N_7909,N_7846,N_7773);
xor U7910 (N_7910,N_7854,N_7835);
and U7911 (N_7911,N_7760,N_7756);
nand U7912 (N_7912,N_7808,N_7763);
nor U7913 (N_7913,N_7852,N_7831);
and U7914 (N_7914,N_7805,N_7856);
xnor U7915 (N_7915,N_7844,N_7779);
or U7916 (N_7916,N_7766,N_7873);
nand U7917 (N_7917,N_7780,N_7762);
or U7918 (N_7918,N_7832,N_7778);
nor U7919 (N_7919,N_7753,N_7828);
nor U7920 (N_7920,N_7843,N_7850);
and U7921 (N_7921,N_7786,N_7822);
and U7922 (N_7922,N_7767,N_7809);
nand U7923 (N_7923,N_7797,N_7783);
and U7924 (N_7924,N_7776,N_7851);
and U7925 (N_7925,N_7833,N_7859);
nand U7926 (N_7926,N_7790,N_7840);
or U7927 (N_7927,N_7787,N_7838);
nor U7928 (N_7928,N_7871,N_7870);
xnor U7929 (N_7929,N_7863,N_7750);
xnor U7930 (N_7930,N_7803,N_7771);
xnor U7931 (N_7931,N_7796,N_7761);
nand U7932 (N_7932,N_7853,N_7815);
or U7933 (N_7933,N_7819,N_7868);
nand U7934 (N_7934,N_7785,N_7757);
and U7935 (N_7935,N_7807,N_7841);
nor U7936 (N_7936,N_7759,N_7810);
nand U7937 (N_7937,N_7774,N_7816);
nor U7938 (N_7938,N_7822,N_7792);
nor U7939 (N_7939,N_7785,N_7863);
and U7940 (N_7940,N_7813,N_7770);
nand U7941 (N_7941,N_7770,N_7868);
nand U7942 (N_7942,N_7834,N_7821);
nand U7943 (N_7943,N_7784,N_7867);
and U7944 (N_7944,N_7786,N_7860);
or U7945 (N_7945,N_7791,N_7872);
or U7946 (N_7946,N_7775,N_7786);
or U7947 (N_7947,N_7774,N_7834);
xnor U7948 (N_7948,N_7760,N_7844);
and U7949 (N_7949,N_7829,N_7784);
or U7950 (N_7950,N_7838,N_7830);
nor U7951 (N_7951,N_7802,N_7846);
nor U7952 (N_7952,N_7861,N_7764);
or U7953 (N_7953,N_7805,N_7822);
nand U7954 (N_7954,N_7783,N_7792);
and U7955 (N_7955,N_7854,N_7840);
and U7956 (N_7956,N_7791,N_7841);
xnor U7957 (N_7957,N_7768,N_7853);
nor U7958 (N_7958,N_7841,N_7850);
xor U7959 (N_7959,N_7821,N_7758);
xnor U7960 (N_7960,N_7750,N_7854);
or U7961 (N_7961,N_7793,N_7813);
and U7962 (N_7962,N_7816,N_7854);
or U7963 (N_7963,N_7869,N_7776);
xor U7964 (N_7964,N_7804,N_7848);
and U7965 (N_7965,N_7838,N_7848);
nor U7966 (N_7966,N_7779,N_7773);
nor U7967 (N_7967,N_7808,N_7863);
xor U7968 (N_7968,N_7832,N_7795);
xnor U7969 (N_7969,N_7806,N_7871);
nor U7970 (N_7970,N_7852,N_7800);
xnor U7971 (N_7971,N_7770,N_7853);
and U7972 (N_7972,N_7780,N_7833);
xnor U7973 (N_7973,N_7847,N_7820);
nand U7974 (N_7974,N_7824,N_7802);
and U7975 (N_7975,N_7839,N_7827);
or U7976 (N_7976,N_7800,N_7858);
xnor U7977 (N_7977,N_7856,N_7853);
and U7978 (N_7978,N_7837,N_7764);
nand U7979 (N_7979,N_7835,N_7813);
nand U7980 (N_7980,N_7839,N_7789);
nor U7981 (N_7981,N_7795,N_7834);
or U7982 (N_7982,N_7781,N_7870);
nand U7983 (N_7983,N_7831,N_7753);
nand U7984 (N_7984,N_7766,N_7835);
nand U7985 (N_7985,N_7847,N_7845);
xnor U7986 (N_7986,N_7842,N_7817);
nand U7987 (N_7987,N_7767,N_7806);
nand U7988 (N_7988,N_7832,N_7769);
or U7989 (N_7989,N_7799,N_7821);
xor U7990 (N_7990,N_7835,N_7800);
nor U7991 (N_7991,N_7775,N_7785);
nor U7992 (N_7992,N_7759,N_7873);
and U7993 (N_7993,N_7796,N_7768);
and U7994 (N_7994,N_7755,N_7828);
and U7995 (N_7995,N_7827,N_7869);
or U7996 (N_7996,N_7765,N_7821);
or U7997 (N_7997,N_7792,N_7791);
and U7998 (N_7998,N_7862,N_7817);
xor U7999 (N_7999,N_7851,N_7786);
nor U8000 (N_8000,N_7997,N_7945);
nor U8001 (N_8001,N_7957,N_7949);
xor U8002 (N_8002,N_7907,N_7956);
xnor U8003 (N_8003,N_7977,N_7995);
and U8004 (N_8004,N_7928,N_7994);
nor U8005 (N_8005,N_7989,N_7937);
nor U8006 (N_8006,N_7887,N_7881);
and U8007 (N_8007,N_7953,N_7976);
nor U8008 (N_8008,N_7894,N_7938);
xnor U8009 (N_8009,N_7983,N_7886);
nor U8010 (N_8010,N_7958,N_7923);
nor U8011 (N_8011,N_7925,N_7988);
or U8012 (N_8012,N_7939,N_7934);
nand U8013 (N_8013,N_7991,N_7932);
and U8014 (N_8014,N_7965,N_7884);
nor U8015 (N_8015,N_7968,N_7936);
and U8016 (N_8016,N_7924,N_7890);
and U8017 (N_8017,N_7975,N_7900);
xnor U8018 (N_8018,N_7926,N_7960);
and U8019 (N_8019,N_7996,N_7972);
and U8020 (N_8020,N_7948,N_7973);
and U8021 (N_8021,N_7969,N_7930);
nor U8022 (N_8022,N_7971,N_7911);
and U8023 (N_8023,N_7979,N_7878);
and U8024 (N_8024,N_7875,N_7920);
nor U8025 (N_8025,N_7889,N_7891);
or U8026 (N_8026,N_7947,N_7974);
xor U8027 (N_8027,N_7944,N_7966);
xnor U8028 (N_8028,N_7877,N_7897);
and U8029 (N_8029,N_7915,N_7914);
and U8030 (N_8030,N_7964,N_7987);
xnor U8031 (N_8031,N_7982,N_7961);
xor U8032 (N_8032,N_7980,N_7883);
nor U8033 (N_8033,N_7910,N_7908);
xor U8034 (N_8034,N_7888,N_7992);
or U8035 (N_8035,N_7963,N_7954);
and U8036 (N_8036,N_7893,N_7892);
nand U8037 (N_8037,N_7985,N_7902);
nand U8038 (N_8038,N_7896,N_7913);
or U8039 (N_8039,N_7921,N_7919);
and U8040 (N_8040,N_7998,N_7955);
and U8041 (N_8041,N_7999,N_7901);
nor U8042 (N_8042,N_7927,N_7912);
xor U8043 (N_8043,N_7993,N_7904);
nor U8044 (N_8044,N_7918,N_7940);
nand U8045 (N_8045,N_7962,N_7906);
or U8046 (N_8046,N_7880,N_7984);
xnor U8047 (N_8047,N_7935,N_7950);
xor U8048 (N_8048,N_7946,N_7942);
xor U8049 (N_8049,N_7895,N_7952);
nor U8050 (N_8050,N_7898,N_7990);
nor U8051 (N_8051,N_7876,N_7951);
xnor U8052 (N_8052,N_7882,N_7903);
nand U8053 (N_8053,N_7967,N_7981);
and U8054 (N_8054,N_7917,N_7959);
nand U8055 (N_8055,N_7899,N_7933);
xnor U8056 (N_8056,N_7943,N_7929);
and U8057 (N_8057,N_7885,N_7879);
xnor U8058 (N_8058,N_7922,N_7978);
and U8059 (N_8059,N_7905,N_7986);
or U8060 (N_8060,N_7941,N_7916);
or U8061 (N_8061,N_7931,N_7970);
or U8062 (N_8062,N_7909,N_7967);
nand U8063 (N_8063,N_7910,N_7985);
nor U8064 (N_8064,N_7953,N_7973);
xor U8065 (N_8065,N_7894,N_7945);
and U8066 (N_8066,N_7941,N_7926);
and U8067 (N_8067,N_7924,N_7995);
and U8068 (N_8068,N_7991,N_7950);
xnor U8069 (N_8069,N_7971,N_7882);
nand U8070 (N_8070,N_7933,N_7995);
nand U8071 (N_8071,N_7940,N_7989);
and U8072 (N_8072,N_7898,N_7949);
xor U8073 (N_8073,N_7884,N_7960);
and U8074 (N_8074,N_7952,N_7963);
and U8075 (N_8075,N_7891,N_7963);
xnor U8076 (N_8076,N_7923,N_7983);
nand U8077 (N_8077,N_7903,N_7907);
and U8078 (N_8078,N_7958,N_7957);
or U8079 (N_8079,N_7965,N_7957);
xnor U8080 (N_8080,N_7881,N_7925);
or U8081 (N_8081,N_7939,N_7930);
xnor U8082 (N_8082,N_7963,N_7971);
nand U8083 (N_8083,N_7935,N_7944);
nand U8084 (N_8084,N_7932,N_7970);
nand U8085 (N_8085,N_7894,N_7915);
nor U8086 (N_8086,N_7877,N_7886);
nand U8087 (N_8087,N_7946,N_7897);
nand U8088 (N_8088,N_7960,N_7980);
xor U8089 (N_8089,N_7961,N_7888);
nand U8090 (N_8090,N_7901,N_7895);
nor U8091 (N_8091,N_7912,N_7977);
xor U8092 (N_8092,N_7897,N_7942);
and U8093 (N_8093,N_7929,N_7991);
xor U8094 (N_8094,N_7876,N_7878);
nor U8095 (N_8095,N_7958,N_7898);
nor U8096 (N_8096,N_7883,N_7952);
xnor U8097 (N_8097,N_7980,N_7998);
or U8098 (N_8098,N_7895,N_7987);
and U8099 (N_8099,N_7911,N_7959);
or U8100 (N_8100,N_7892,N_7935);
nor U8101 (N_8101,N_7997,N_7960);
xor U8102 (N_8102,N_7876,N_7875);
nor U8103 (N_8103,N_7951,N_7972);
nor U8104 (N_8104,N_7927,N_7941);
and U8105 (N_8105,N_7968,N_7992);
nor U8106 (N_8106,N_7958,N_7908);
nand U8107 (N_8107,N_7940,N_7921);
nor U8108 (N_8108,N_7931,N_7980);
nand U8109 (N_8109,N_7929,N_7888);
nand U8110 (N_8110,N_7926,N_7993);
xnor U8111 (N_8111,N_7906,N_7954);
and U8112 (N_8112,N_7889,N_7958);
and U8113 (N_8113,N_7988,N_7920);
nand U8114 (N_8114,N_7951,N_7944);
nor U8115 (N_8115,N_7949,N_7876);
xor U8116 (N_8116,N_7951,N_7883);
xor U8117 (N_8117,N_7922,N_7985);
nor U8118 (N_8118,N_7940,N_7933);
nand U8119 (N_8119,N_7967,N_7889);
nor U8120 (N_8120,N_7975,N_7921);
nand U8121 (N_8121,N_7878,N_7926);
and U8122 (N_8122,N_7910,N_7994);
nor U8123 (N_8123,N_7945,N_7980);
or U8124 (N_8124,N_7909,N_7919);
nor U8125 (N_8125,N_8107,N_8098);
xnor U8126 (N_8126,N_8058,N_8005);
nand U8127 (N_8127,N_8026,N_8104);
nor U8128 (N_8128,N_8113,N_8096);
and U8129 (N_8129,N_8059,N_8081);
nand U8130 (N_8130,N_8067,N_8031);
nor U8131 (N_8131,N_8063,N_8011);
and U8132 (N_8132,N_8003,N_8043);
or U8133 (N_8133,N_8123,N_8124);
nand U8134 (N_8134,N_8013,N_8055);
or U8135 (N_8135,N_8066,N_8080);
and U8136 (N_8136,N_8040,N_8045);
nand U8137 (N_8137,N_8074,N_8052);
nor U8138 (N_8138,N_8101,N_8097);
or U8139 (N_8139,N_8054,N_8092);
nand U8140 (N_8140,N_8023,N_8103);
and U8141 (N_8141,N_8072,N_8088);
nor U8142 (N_8142,N_8000,N_8093);
xnor U8143 (N_8143,N_8118,N_8051);
xnor U8144 (N_8144,N_8095,N_8114);
xnor U8145 (N_8145,N_8062,N_8071);
or U8146 (N_8146,N_8086,N_8065);
xnor U8147 (N_8147,N_8120,N_8090);
nor U8148 (N_8148,N_8057,N_8001);
or U8149 (N_8149,N_8010,N_8102);
and U8150 (N_8150,N_8046,N_8060);
nor U8151 (N_8151,N_8047,N_8079);
nor U8152 (N_8152,N_8024,N_8091);
and U8153 (N_8153,N_8006,N_8110);
or U8154 (N_8154,N_8056,N_8068);
nand U8155 (N_8155,N_8094,N_8069);
nor U8156 (N_8156,N_8077,N_8112);
and U8157 (N_8157,N_8004,N_8082);
xor U8158 (N_8158,N_8034,N_8032);
xnor U8159 (N_8159,N_8012,N_8035);
and U8160 (N_8160,N_8119,N_8087);
or U8161 (N_8161,N_8108,N_8050);
xnor U8162 (N_8162,N_8117,N_8076);
and U8163 (N_8163,N_8021,N_8027);
and U8164 (N_8164,N_8100,N_8075);
nor U8165 (N_8165,N_8029,N_8044);
and U8166 (N_8166,N_8033,N_8030);
and U8167 (N_8167,N_8041,N_8121);
and U8168 (N_8168,N_8115,N_8038);
xnor U8169 (N_8169,N_8070,N_8016);
nand U8170 (N_8170,N_8020,N_8002);
nor U8171 (N_8171,N_8022,N_8036);
or U8172 (N_8172,N_8019,N_8078);
or U8173 (N_8173,N_8008,N_8009);
xnor U8174 (N_8174,N_8015,N_8039);
nor U8175 (N_8175,N_8099,N_8014);
nor U8176 (N_8176,N_8028,N_8105);
nand U8177 (N_8177,N_8111,N_8083);
or U8178 (N_8178,N_8049,N_8089);
nand U8179 (N_8179,N_8061,N_8064);
nand U8180 (N_8180,N_8109,N_8018);
nand U8181 (N_8181,N_8007,N_8084);
and U8182 (N_8182,N_8048,N_8025);
xnor U8183 (N_8183,N_8116,N_8122);
nor U8184 (N_8184,N_8042,N_8037);
nor U8185 (N_8185,N_8106,N_8017);
or U8186 (N_8186,N_8085,N_8053);
xnor U8187 (N_8187,N_8073,N_8054);
or U8188 (N_8188,N_8078,N_8055);
and U8189 (N_8189,N_8025,N_8100);
xnor U8190 (N_8190,N_8076,N_8080);
nand U8191 (N_8191,N_8091,N_8030);
and U8192 (N_8192,N_8055,N_8056);
nand U8193 (N_8193,N_8016,N_8063);
and U8194 (N_8194,N_8043,N_8076);
or U8195 (N_8195,N_8070,N_8105);
or U8196 (N_8196,N_8058,N_8012);
and U8197 (N_8197,N_8061,N_8070);
nor U8198 (N_8198,N_8059,N_8070);
nand U8199 (N_8199,N_8005,N_8101);
xor U8200 (N_8200,N_8112,N_8036);
xnor U8201 (N_8201,N_8101,N_8036);
nand U8202 (N_8202,N_8099,N_8074);
nand U8203 (N_8203,N_8086,N_8108);
nor U8204 (N_8204,N_8009,N_8114);
nor U8205 (N_8205,N_8001,N_8015);
or U8206 (N_8206,N_8118,N_8109);
nand U8207 (N_8207,N_8009,N_8010);
nor U8208 (N_8208,N_8022,N_8094);
xnor U8209 (N_8209,N_8091,N_8124);
nand U8210 (N_8210,N_8019,N_8030);
xor U8211 (N_8211,N_8018,N_8099);
or U8212 (N_8212,N_8040,N_8042);
nor U8213 (N_8213,N_8076,N_8113);
or U8214 (N_8214,N_8006,N_8075);
nand U8215 (N_8215,N_8108,N_8062);
nand U8216 (N_8216,N_8121,N_8033);
xnor U8217 (N_8217,N_8049,N_8041);
nor U8218 (N_8218,N_8117,N_8070);
or U8219 (N_8219,N_8087,N_8001);
and U8220 (N_8220,N_8051,N_8087);
nand U8221 (N_8221,N_8071,N_8102);
and U8222 (N_8222,N_8075,N_8110);
or U8223 (N_8223,N_8030,N_8000);
or U8224 (N_8224,N_8000,N_8096);
nor U8225 (N_8225,N_8035,N_8092);
or U8226 (N_8226,N_8013,N_8088);
or U8227 (N_8227,N_8079,N_8086);
nor U8228 (N_8228,N_8060,N_8095);
nor U8229 (N_8229,N_8057,N_8120);
and U8230 (N_8230,N_8082,N_8006);
nor U8231 (N_8231,N_8004,N_8099);
xor U8232 (N_8232,N_8061,N_8119);
and U8233 (N_8233,N_8059,N_8080);
or U8234 (N_8234,N_8091,N_8066);
or U8235 (N_8235,N_8112,N_8054);
nand U8236 (N_8236,N_8054,N_8067);
and U8237 (N_8237,N_8071,N_8113);
or U8238 (N_8238,N_8009,N_8108);
nor U8239 (N_8239,N_8053,N_8063);
nand U8240 (N_8240,N_8069,N_8087);
xnor U8241 (N_8241,N_8114,N_8056);
and U8242 (N_8242,N_8011,N_8100);
or U8243 (N_8243,N_8037,N_8033);
nand U8244 (N_8244,N_8101,N_8006);
nor U8245 (N_8245,N_8112,N_8081);
nand U8246 (N_8246,N_8046,N_8054);
nor U8247 (N_8247,N_8079,N_8089);
nor U8248 (N_8248,N_8073,N_8089);
or U8249 (N_8249,N_8002,N_8028);
nand U8250 (N_8250,N_8194,N_8243);
and U8251 (N_8251,N_8162,N_8132);
nor U8252 (N_8252,N_8128,N_8181);
nand U8253 (N_8253,N_8158,N_8240);
xor U8254 (N_8254,N_8157,N_8223);
xor U8255 (N_8255,N_8153,N_8142);
xnor U8256 (N_8256,N_8166,N_8236);
nor U8257 (N_8257,N_8148,N_8228);
nand U8258 (N_8258,N_8202,N_8195);
or U8259 (N_8259,N_8186,N_8156);
nand U8260 (N_8260,N_8245,N_8238);
nor U8261 (N_8261,N_8174,N_8214);
or U8262 (N_8262,N_8159,N_8190);
or U8263 (N_8263,N_8141,N_8231);
or U8264 (N_8264,N_8176,N_8237);
nand U8265 (N_8265,N_8163,N_8150);
xor U8266 (N_8266,N_8139,N_8248);
xor U8267 (N_8267,N_8161,N_8241);
xnor U8268 (N_8268,N_8235,N_8143);
nor U8269 (N_8269,N_8191,N_8232);
nand U8270 (N_8270,N_8199,N_8183);
nor U8271 (N_8271,N_8178,N_8207);
nand U8272 (N_8272,N_8219,N_8145);
xor U8273 (N_8273,N_8244,N_8217);
or U8274 (N_8274,N_8220,N_8213);
nand U8275 (N_8275,N_8180,N_8247);
or U8276 (N_8276,N_8221,N_8184);
or U8277 (N_8277,N_8135,N_8204);
or U8278 (N_8278,N_8222,N_8133);
or U8279 (N_8279,N_8125,N_8179);
xnor U8280 (N_8280,N_8138,N_8226);
nand U8281 (N_8281,N_8154,N_8215);
nand U8282 (N_8282,N_8177,N_8234);
and U8283 (N_8283,N_8149,N_8146);
nand U8284 (N_8284,N_8196,N_8227);
and U8285 (N_8285,N_8209,N_8151);
nand U8286 (N_8286,N_8144,N_8140);
or U8287 (N_8287,N_8185,N_8165);
nand U8288 (N_8288,N_8224,N_8246);
or U8289 (N_8289,N_8167,N_8208);
nor U8290 (N_8290,N_8193,N_8187);
or U8291 (N_8291,N_8200,N_8160);
nor U8292 (N_8292,N_8155,N_8233);
or U8293 (N_8293,N_8225,N_8172);
nand U8294 (N_8294,N_8203,N_8127);
and U8295 (N_8295,N_8218,N_8188);
nand U8296 (N_8296,N_8189,N_8130);
and U8297 (N_8297,N_8152,N_8212);
xor U8298 (N_8298,N_8249,N_8216);
nand U8299 (N_8299,N_8229,N_8173);
and U8300 (N_8300,N_8129,N_8175);
xor U8301 (N_8301,N_8134,N_8201);
nand U8302 (N_8302,N_8192,N_8197);
nand U8303 (N_8303,N_8169,N_8171);
or U8304 (N_8304,N_8170,N_8182);
and U8305 (N_8305,N_8242,N_8205);
and U8306 (N_8306,N_8198,N_8131);
and U8307 (N_8307,N_8126,N_8230);
or U8308 (N_8308,N_8164,N_8239);
nand U8309 (N_8309,N_8206,N_8147);
nand U8310 (N_8310,N_8136,N_8168);
or U8311 (N_8311,N_8137,N_8210);
nand U8312 (N_8312,N_8211,N_8166);
and U8313 (N_8313,N_8170,N_8237);
or U8314 (N_8314,N_8198,N_8141);
nand U8315 (N_8315,N_8174,N_8240);
nand U8316 (N_8316,N_8189,N_8157);
or U8317 (N_8317,N_8216,N_8158);
nor U8318 (N_8318,N_8237,N_8245);
xnor U8319 (N_8319,N_8149,N_8158);
xor U8320 (N_8320,N_8217,N_8208);
nand U8321 (N_8321,N_8138,N_8220);
nor U8322 (N_8322,N_8171,N_8220);
or U8323 (N_8323,N_8184,N_8189);
nor U8324 (N_8324,N_8203,N_8231);
nor U8325 (N_8325,N_8211,N_8210);
xnor U8326 (N_8326,N_8205,N_8176);
and U8327 (N_8327,N_8132,N_8200);
nand U8328 (N_8328,N_8198,N_8219);
or U8329 (N_8329,N_8171,N_8179);
nand U8330 (N_8330,N_8189,N_8190);
xnor U8331 (N_8331,N_8220,N_8142);
and U8332 (N_8332,N_8207,N_8127);
and U8333 (N_8333,N_8244,N_8183);
nor U8334 (N_8334,N_8128,N_8195);
nor U8335 (N_8335,N_8155,N_8220);
or U8336 (N_8336,N_8128,N_8193);
nand U8337 (N_8337,N_8192,N_8128);
or U8338 (N_8338,N_8145,N_8137);
xor U8339 (N_8339,N_8194,N_8241);
nor U8340 (N_8340,N_8228,N_8218);
nor U8341 (N_8341,N_8166,N_8126);
nor U8342 (N_8342,N_8128,N_8194);
nand U8343 (N_8343,N_8185,N_8218);
and U8344 (N_8344,N_8214,N_8141);
nor U8345 (N_8345,N_8199,N_8152);
or U8346 (N_8346,N_8242,N_8178);
or U8347 (N_8347,N_8161,N_8249);
and U8348 (N_8348,N_8165,N_8237);
or U8349 (N_8349,N_8141,N_8136);
or U8350 (N_8350,N_8222,N_8201);
nand U8351 (N_8351,N_8142,N_8150);
xnor U8352 (N_8352,N_8218,N_8191);
and U8353 (N_8353,N_8191,N_8192);
and U8354 (N_8354,N_8149,N_8142);
nor U8355 (N_8355,N_8236,N_8149);
or U8356 (N_8356,N_8213,N_8237);
and U8357 (N_8357,N_8204,N_8206);
and U8358 (N_8358,N_8152,N_8241);
or U8359 (N_8359,N_8228,N_8235);
or U8360 (N_8360,N_8167,N_8195);
nand U8361 (N_8361,N_8167,N_8185);
or U8362 (N_8362,N_8161,N_8177);
and U8363 (N_8363,N_8226,N_8127);
nor U8364 (N_8364,N_8151,N_8183);
nor U8365 (N_8365,N_8166,N_8173);
nand U8366 (N_8366,N_8158,N_8230);
nor U8367 (N_8367,N_8172,N_8215);
nor U8368 (N_8368,N_8234,N_8205);
or U8369 (N_8369,N_8192,N_8209);
or U8370 (N_8370,N_8165,N_8186);
nor U8371 (N_8371,N_8185,N_8228);
and U8372 (N_8372,N_8131,N_8210);
nor U8373 (N_8373,N_8142,N_8174);
or U8374 (N_8374,N_8248,N_8213);
or U8375 (N_8375,N_8289,N_8327);
nor U8376 (N_8376,N_8262,N_8269);
and U8377 (N_8377,N_8285,N_8311);
nor U8378 (N_8378,N_8310,N_8314);
xnor U8379 (N_8379,N_8374,N_8330);
and U8380 (N_8380,N_8290,N_8312);
nand U8381 (N_8381,N_8363,N_8305);
or U8382 (N_8382,N_8278,N_8292);
xnor U8383 (N_8383,N_8287,N_8264);
nor U8384 (N_8384,N_8325,N_8326);
nor U8385 (N_8385,N_8291,N_8303);
nand U8386 (N_8386,N_8301,N_8293);
nand U8387 (N_8387,N_8283,N_8274);
xor U8388 (N_8388,N_8324,N_8257);
xor U8389 (N_8389,N_8347,N_8344);
or U8390 (N_8390,N_8373,N_8254);
nand U8391 (N_8391,N_8268,N_8252);
xor U8392 (N_8392,N_8365,N_8260);
and U8393 (N_8393,N_8353,N_8317);
and U8394 (N_8394,N_8309,N_8250);
and U8395 (N_8395,N_8313,N_8316);
nand U8396 (N_8396,N_8367,N_8259);
nor U8397 (N_8397,N_8261,N_8315);
nand U8398 (N_8398,N_8286,N_8271);
nand U8399 (N_8399,N_8362,N_8369);
and U8400 (N_8400,N_8253,N_8323);
nor U8401 (N_8401,N_8280,N_8336);
and U8402 (N_8402,N_8334,N_8361);
nand U8403 (N_8403,N_8308,N_8277);
or U8404 (N_8404,N_8318,N_8299);
or U8405 (N_8405,N_8339,N_8349);
nor U8406 (N_8406,N_8300,N_8284);
nand U8407 (N_8407,N_8302,N_8256);
or U8408 (N_8408,N_8272,N_8343);
and U8409 (N_8409,N_8304,N_8298);
or U8410 (N_8410,N_8354,N_8360);
or U8411 (N_8411,N_8306,N_8333);
nor U8412 (N_8412,N_8281,N_8279);
or U8413 (N_8413,N_8251,N_8267);
nor U8414 (N_8414,N_8351,N_8342);
nand U8415 (N_8415,N_8258,N_8255);
and U8416 (N_8416,N_8357,N_8337);
and U8417 (N_8417,N_8359,N_8341);
nor U8418 (N_8418,N_8370,N_8358);
and U8419 (N_8419,N_8335,N_8366);
and U8420 (N_8420,N_8295,N_8294);
or U8421 (N_8421,N_8331,N_8273);
or U8422 (N_8422,N_8332,N_8282);
or U8423 (N_8423,N_8322,N_8346);
nor U8424 (N_8424,N_8364,N_8372);
or U8425 (N_8425,N_8328,N_8266);
and U8426 (N_8426,N_8276,N_8270);
nor U8427 (N_8427,N_8296,N_8368);
and U8428 (N_8428,N_8340,N_8352);
nor U8429 (N_8429,N_8345,N_8275);
xor U8430 (N_8430,N_8350,N_8319);
and U8431 (N_8431,N_8329,N_8288);
xor U8432 (N_8432,N_8355,N_8265);
and U8433 (N_8433,N_8307,N_8371);
or U8434 (N_8434,N_8297,N_8338);
nor U8435 (N_8435,N_8356,N_8320);
xor U8436 (N_8436,N_8321,N_8263);
nor U8437 (N_8437,N_8348,N_8351);
or U8438 (N_8438,N_8301,N_8264);
or U8439 (N_8439,N_8258,N_8294);
or U8440 (N_8440,N_8305,N_8278);
nand U8441 (N_8441,N_8332,N_8256);
xor U8442 (N_8442,N_8321,N_8346);
or U8443 (N_8443,N_8303,N_8316);
and U8444 (N_8444,N_8256,N_8314);
xnor U8445 (N_8445,N_8259,N_8323);
or U8446 (N_8446,N_8330,N_8284);
nor U8447 (N_8447,N_8370,N_8273);
nor U8448 (N_8448,N_8310,N_8371);
nand U8449 (N_8449,N_8259,N_8261);
xnor U8450 (N_8450,N_8254,N_8316);
xor U8451 (N_8451,N_8335,N_8305);
nand U8452 (N_8452,N_8334,N_8370);
nor U8453 (N_8453,N_8359,N_8269);
nor U8454 (N_8454,N_8255,N_8250);
or U8455 (N_8455,N_8264,N_8307);
xor U8456 (N_8456,N_8258,N_8363);
nor U8457 (N_8457,N_8265,N_8325);
nand U8458 (N_8458,N_8254,N_8279);
or U8459 (N_8459,N_8312,N_8366);
or U8460 (N_8460,N_8306,N_8307);
xnor U8461 (N_8461,N_8256,N_8297);
xor U8462 (N_8462,N_8358,N_8292);
nand U8463 (N_8463,N_8330,N_8370);
xor U8464 (N_8464,N_8289,N_8365);
and U8465 (N_8465,N_8362,N_8371);
and U8466 (N_8466,N_8299,N_8305);
xnor U8467 (N_8467,N_8284,N_8267);
nor U8468 (N_8468,N_8336,N_8267);
nand U8469 (N_8469,N_8340,N_8263);
nor U8470 (N_8470,N_8305,N_8294);
or U8471 (N_8471,N_8331,N_8371);
nor U8472 (N_8472,N_8317,N_8361);
xor U8473 (N_8473,N_8368,N_8274);
or U8474 (N_8474,N_8341,N_8303);
nor U8475 (N_8475,N_8309,N_8278);
xnor U8476 (N_8476,N_8362,N_8281);
and U8477 (N_8477,N_8259,N_8354);
nand U8478 (N_8478,N_8319,N_8337);
xnor U8479 (N_8479,N_8282,N_8257);
or U8480 (N_8480,N_8282,N_8258);
nor U8481 (N_8481,N_8268,N_8287);
xnor U8482 (N_8482,N_8311,N_8310);
nand U8483 (N_8483,N_8348,N_8282);
nor U8484 (N_8484,N_8274,N_8252);
xnor U8485 (N_8485,N_8260,N_8262);
xnor U8486 (N_8486,N_8359,N_8342);
nor U8487 (N_8487,N_8334,N_8292);
nand U8488 (N_8488,N_8287,N_8312);
xor U8489 (N_8489,N_8289,N_8321);
or U8490 (N_8490,N_8341,N_8306);
and U8491 (N_8491,N_8317,N_8273);
nand U8492 (N_8492,N_8275,N_8325);
nand U8493 (N_8493,N_8254,N_8256);
nor U8494 (N_8494,N_8334,N_8312);
nor U8495 (N_8495,N_8349,N_8268);
xnor U8496 (N_8496,N_8354,N_8337);
or U8497 (N_8497,N_8281,N_8288);
or U8498 (N_8498,N_8369,N_8319);
xnor U8499 (N_8499,N_8366,N_8313);
and U8500 (N_8500,N_8401,N_8408);
and U8501 (N_8501,N_8416,N_8464);
nor U8502 (N_8502,N_8398,N_8460);
xor U8503 (N_8503,N_8425,N_8466);
and U8504 (N_8504,N_8428,N_8410);
nand U8505 (N_8505,N_8493,N_8494);
nand U8506 (N_8506,N_8394,N_8459);
and U8507 (N_8507,N_8400,N_8442);
nor U8508 (N_8508,N_8386,N_8472);
nand U8509 (N_8509,N_8420,N_8499);
nand U8510 (N_8510,N_8443,N_8387);
xnor U8511 (N_8511,N_8430,N_8393);
nand U8512 (N_8512,N_8414,N_8432);
or U8513 (N_8513,N_8429,N_8462);
nand U8514 (N_8514,N_8457,N_8470);
xor U8515 (N_8515,N_8488,N_8446);
and U8516 (N_8516,N_8439,N_8495);
or U8517 (N_8517,N_8406,N_8437);
nand U8518 (N_8518,N_8385,N_8407);
and U8519 (N_8519,N_8456,N_8378);
xor U8520 (N_8520,N_8476,N_8424);
and U8521 (N_8521,N_8423,N_8480);
nand U8522 (N_8522,N_8461,N_8389);
xnor U8523 (N_8523,N_8375,N_8399);
or U8524 (N_8524,N_8452,N_8477);
and U8525 (N_8525,N_8433,N_8403);
nor U8526 (N_8526,N_8463,N_8479);
xor U8527 (N_8527,N_8381,N_8483);
and U8528 (N_8528,N_8421,N_8413);
nor U8529 (N_8529,N_8418,N_8497);
nand U8530 (N_8530,N_8447,N_8434);
nand U8531 (N_8531,N_8467,N_8390);
nand U8532 (N_8532,N_8475,N_8422);
nor U8533 (N_8533,N_8445,N_8468);
nand U8534 (N_8534,N_8485,N_8496);
xor U8535 (N_8535,N_8454,N_8379);
or U8536 (N_8536,N_8486,N_8478);
nand U8537 (N_8537,N_8473,N_8491);
nand U8538 (N_8538,N_8487,N_8490);
xnor U8539 (N_8539,N_8427,N_8431);
and U8540 (N_8540,N_8382,N_8380);
nor U8541 (N_8541,N_8458,N_8384);
and U8542 (N_8542,N_8409,N_8396);
or U8543 (N_8543,N_8397,N_8383);
nand U8544 (N_8544,N_8469,N_8426);
or U8545 (N_8545,N_8444,N_8405);
nand U8546 (N_8546,N_8484,N_8489);
nor U8547 (N_8547,N_8436,N_8419);
xnor U8548 (N_8548,N_8417,N_8481);
and U8549 (N_8549,N_8455,N_8498);
or U8550 (N_8550,N_8492,N_8474);
xor U8551 (N_8551,N_8448,N_8402);
nor U8552 (N_8552,N_8411,N_8377);
nand U8553 (N_8553,N_8435,N_8388);
xnor U8554 (N_8554,N_8412,N_8465);
nand U8555 (N_8555,N_8404,N_8453);
or U8556 (N_8556,N_8438,N_8415);
nand U8557 (N_8557,N_8392,N_8376);
or U8558 (N_8558,N_8450,N_8440);
and U8559 (N_8559,N_8441,N_8391);
or U8560 (N_8560,N_8395,N_8449);
or U8561 (N_8561,N_8471,N_8451);
xor U8562 (N_8562,N_8482,N_8403);
or U8563 (N_8563,N_8438,N_8419);
or U8564 (N_8564,N_8451,N_8482);
nand U8565 (N_8565,N_8458,N_8414);
or U8566 (N_8566,N_8376,N_8492);
or U8567 (N_8567,N_8398,N_8479);
and U8568 (N_8568,N_8439,N_8454);
nor U8569 (N_8569,N_8461,N_8428);
nor U8570 (N_8570,N_8497,N_8375);
or U8571 (N_8571,N_8467,N_8481);
nand U8572 (N_8572,N_8479,N_8452);
or U8573 (N_8573,N_8431,N_8496);
and U8574 (N_8574,N_8454,N_8456);
and U8575 (N_8575,N_8383,N_8418);
and U8576 (N_8576,N_8411,N_8479);
or U8577 (N_8577,N_8401,N_8457);
and U8578 (N_8578,N_8492,N_8484);
nor U8579 (N_8579,N_8458,N_8383);
nand U8580 (N_8580,N_8486,N_8376);
or U8581 (N_8581,N_8496,N_8494);
and U8582 (N_8582,N_8455,N_8402);
nor U8583 (N_8583,N_8491,N_8384);
nand U8584 (N_8584,N_8448,N_8451);
xor U8585 (N_8585,N_8462,N_8379);
nand U8586 (N_8586,N_8461,N_8397);
and U8587 (N_8587,N_8434,N_8495);
or U8588 (N_8588,N_8415,N_8471);
or U8589 (N_8589,N_8398,N_8475);
nand U8590 (N_8590,N_8425,N_8491);
xor U8591 (N_8591,N_8417,N_8387);
and U8592 (N_8592,N_8469,N_8408);
xor U8593 (N_8593,N_8426,N_8412);
nor U8594 (N_8594,N_8387,N_8382);
and U8595 (N_8595,N_8382,N_8407);
nand U8596 (N_8596,N_8395,N_8413);
and U8597 (N_8597,N_8480,N_8394);
xnor U8598 (N_8598,N_8493,N_8466);
or U8599 (N_8599,N_8386,N_8394);
nand U8600 (N_8600,N_8393,N_8444);
and U8601 (N_8601,N_8470,N_8449);
nand U8602 (N_8602,N_8425,N_8378);
nor U8603 (N_8603,N_8409,N_8498);
xnor U8604 (N_8604,N_8444,N_8375);
nand U8605 (N_8605,N_8475,N_8498);
or U8606 (N_8606,N_8393,N_8399);
nand U8607 (N_8607,N_8490,N_8421);
or U8608 (N_8608,N_8437,N_8476);
or U8609 (N_8609,N_8451,N_8489);
nor U8610 (N_8610,N_8418,N_8441);
nor U8611 (N_8611,N_8404,N_8398);
or U8612 (N_8612,N_8421,N_8395);
nor U8613 (N_8613,N_8478,N_8416);
or U8614 (N_8614,N_8418,N_8394);
xnor U8615 (N_8615,N_8391,N_8490);
nor U8616 (N_8616,N_8478,N_8396);
nand U8617 (N_8617,N_8398,N_8441);
or U8618 (N_8618,N_8475,N_8429);
nand U8619 (N_8619,N_8494,N_8456);
nor U8620 (N_8620,N_8456,N_8434);
xnor U8621 (N_8621,N_8383,N_8376);
or U8622 (N_8622,N_8450,N_8376);
xnor U8623 (N_8623,N_8406,N_8443);
nor U8624 (N_8624,N_8427,N_8488);
nor U8625 (N_8625,N_8520,N_8581);
xor U8626 (N_8626,N_8594,N_8598);
nand U8627 (N_8627,N_8572,N_8624);
nor U8628 (N_8628,N_8558,N_8605);
nand U8629 (N_8629,N_8523,N_8620);
and U8630 (N_8630,N_8585,N_8573);
and U8631 (N_8631,N_8569,N_8515);
xor U8632 (N_8632,N_8593,N_8544);
or U8633 (N_8633,N_8533,N_8513);
and U8634 (N_8634,N_8553,N_8583);
or U8635 (N_8635,N_8562,N_8565);
xor U8636 (N_8636,N_8621,N_8552);
or U8637 (N_8637,N_8619,N_8516);
nor U8638 (N_8638,N_8545,N_8507);
xnor U8639 (N_8639,N_8576,N_8578);
nor U8640 (N_8640,N_8503,N_8556);
nand U8641 (N_8641,N_8525,N_8616);
and U8642 (N_8642,N_8518,N_8604);
xnor U8643 (N_8643,N_8568,N_8577);
and U8644 (N_8644,N_8591,N_8574);
nand U8645 (N_8645,N_8509,N_8606);
or U8646 (N_8646,N_8575,N_8623);
and U8647 (N_8647,N_8590,N_8579);
or U8648 (N_8648,N_8596,N_8511);
nor U8649 (N_8649,N_8506,N_8597);
nand U8650 (N_8650,N_8532,N_8549);
and U8651 (N_8651,N_8550,N_8521);
or U8652 (N_8652,N_8517,N_8524);
and U8653 (N_8653,N_8536,N_8526);
or U8654 (N_8654,N_8530,N_8519);
and U8655 (N_8655,N_8512,N_8618);
nor U8656 (N_8656,N_8551,N_8601);
xnor U8657 (N_8657,N_8534,N_8539);
or U8658 (N_8658,N_8609,N_8502);
and U8659 (N_8659,N_8510,N_8540);
xnor U8660 (N_8660,N_8563,N_8508);
and U8661 (N_8661,N_8610,N_8564);
nor U8662 (N_8662,N_8559,N_8560);
or U8663 (N_8663,N_8622,N_8548);
and U8664 (N_8664,N_8543,N_8613);
and U8665 (N_8665,N_8542,N_8586);
and U8666 (N_8666,N_8541,N_8614);
xnor U8667 (N_8667,N_8504,N_8612);
or U8668 (N_8668,N_8547,N_8603);
and U8669 (N_8669,N_8602,N_8580);
nand U8670 (N_8670,N_8514,N_8588);
nor U8671 (N_8671,N_8505,N_8584);
nor U8672 (N_8672,N_8615,N_8611);
nand U8673 (N_8673,N_8531,N_8567);
or U8674 (N_8674,N_8607,N_8554);
xnor U8675 (N_8675,N_8538,N_8555);
xor U8676 (N_8676,N_8582,N_8608);
and U8677 (N_8677,N_8561,N_8600);
nand U8678 (N_8678,N_8527,N_8528);
nand U8679 (N_8679,N_8522,N_8501);
nor U8680 (N_8680,N_8571,N_8537);
nand U8681 (N_8681,N_8595,N_8500);
xor U8682 (N_8682,N_8546,N_8617);
and U8683 (N_8683,N_8587,N_8589);
nand U8684 (N_8684,N_8566,N_8592);
nand U8685 (N_8685,N_8535,N_8570);
xor U8686 (N_8686,N_8599,N_8529);
nand U8687 (N_8687,N_8557,N_8547);
xor U8688 (N_8688,N_8616,N_8554);
nand U8689 (N_8689,N_8584,N_8574);
nand U8690 (N_8690,N_8523,N_8574);
nor U8691 (N_8691,N_8589,N_8598);
or U8692 (N_8692,N_8567,N_8598);
nor U8693 (N_8693,N_8615,N_8543);
and U8694 (N_8694,N_8564,N_8583);
and U8695 (N_8695,N_8608,N_8564);
xnor U8696 (N_8696,N_8615,N_8530);
nand U8697 (N_8697,N_8528,N_8546);
xnor U8698 (N_8698,N_8586,N_8522);
xor U8699 (N_8699,N_8500,N_8559);
nor U8700 (N_8700,N_8620,N_8596);
and U8701 (N_8701,N_8614,N_8507);
or U8702 (N_8702,N_8597,N_8547);
or U8703 (N_8703,N_8619,N_8580);
xor U8704 (N_8704,N_8588,N_8555);
xnor U8705 (N_8705,N_8523,N_8536);
xor U8706 (N_8706,N_8586,N_8509);
and U8707 (N_8707,N_8538,N_8530);
xor U8708 (N_8708,N_8574,N_8518);
xor U8709 (N_8709,N_8588,N_8594);
nand U8710 (N_8710,N_8503,N_8570);
and U8711 (N_8711,N_8597,N_8585);
xor U8712 (N_8712,N_8516,N_8612);
nor U8713 (N_8713,N_8513,N_8518);
nand U8714 (N_8714,N_8546,N_8603);
xnor U8715 (N_8715,N_8594,N_8617);
nor U8716 (N_8716,N_8621,N_8549);
xnor U8717 (N_8717,N_8616,N_8559);
nand U8718 (N_8718,N_8547,N_8578);
or U8719 (N_8719,N_8511,N_8565);
or U8720 (N_8720,N_8541,N_8517);
and U8721 (N_8721,N_8559,N_8572);
nor U8722 (N_8722,N_8523,N_8509);
and U8723 (N_8723,N_8588,N_8616);
and U8724 (N_8724,N_8552,N_8558);
and U8725 (N_8725,N_8592,N_8598);
or U8726 (N_8726,N_8529,N_8539);
xor U8727 (N_8727,N_8590,N_8585);
nor U8728 (N_8728,N_8519,N_8550);
nand U8729 (N_8729,N_8525,N_8527);
or U8730 (N_8730,N_8569,N_8527);
xnor U8731 (N_8731,N_8553,N_8601);
or U8732 (N_8732,N_8548,N_8507);
nor U8733 (N_8733,N_8540,N_8582);
nor U8734 (N_8734,N_8609,N_8554);
xnor U8735 (N_8735,N_8515,N_8617);
nand U8736 (N_8736,N_8526,N_8624);
nor U8737 (N_8737,N_8587,N_8592);
xnor U8738 (N_8738,N_8526,N_8587);
nand U8739 (N_8739,N_8514,N_8613);
and U8740 (N_8740,N_8570,N_8621);
or U8741 (N_8741,N_8568,N_8598);
or U8742 (N_8742,N_8540,N_8557);
or U8743 (N_8743,N_8608,N_8583);
nand U8744 (N_8744,N_8563,N_8505);
nor U8745 (N_8745,N_8586,N_8506);
and U8746 (N_8746,N_8533,N_8504);
nand U8747 (N_8747,N_8503,N_8577);
or U8748 (N_8748,N_8617,N_8529);
xor U8749 (N_8749,N_8602,N_8518);
nor U8750 (N_8750,N_8648,N_8645);
or U8751 (N_8751,N_8710,N_8658);
nor U8752 (N_8752,N_8721,N_8675);
xor U8753 (N_8753,N_8722,N_8684);
or U8754 (N_8754,N_8679,N_8741);
nand U8755 (N_8755,N_8719,N_8729);
or U8756 (N_8756,N_8716,N_8651);
nor U8757 (N_8757,N_8701,N_8732);
nor U8758 (N_8758,N_8728,N_8738);
and U8759 (N_8759,N_8692,N_8657);
and U8760 (N_8760,N_8724,N_8625);
xor U8761 (N_8761,N_8674,N_8672);
nand U8762 (N_8762,N_8694,N_8681);
nand U8763 (N_8763,N_8659,N_8703);
xor U8764 (N_8764,N_8632,N_8642);
nand U8765 (N_8765,N_8697,N_8673);
nand U8766 (N_8766,N_8714,N_8631);
or U8767 (N_8767,N_8650,N_8737);
nand U8768 (N_8768,N_8706,N_8636);
nand U8769 (N_8769,N_8748,N_8671);
nor U8770 (N_8770,N_8717,N_8709);
and U8771 (N_8771,N_8713,N_8705);
nor U8772 (N_8772,N_8740,N_8654);
or U8773 (N_8773,N_8702,N_8646);
xnor U8774 (N_8774,N_8634,N_8736);
or U8775 (N_8775,N_8667,N_8744);
xor U8776 (N_8776,N_8734,N_8640);
nor U8777 (N_8777,N_8685,N_8656);
or U8778 (N_8778,N_8669,N_8637);
or U8779 (N_8779,N_8628,N_8639);
and U8780 (N_8780,N_8693,N_8688);
nor U8781 (N_8781,N_8689,N_8723);
xnor U8782 (N_8782,N_8660,N_8718);
nand U8783 (N_8783,N_8635,N_8735);
nor U8784 (N_8784,N_8731,N_8727);
and U8785 (N_8785,N_8686,N_8743);
nand U8786 (N_8786,N_8664,N_8653);
and U8787 (N_8787,N_8696,N_8739);
nor U8788 (N_8788,N_8661,N_8643);
xnor U8789 (N_8789,N_8627,N_8691);
and U8790 (N_8790,N_8677,N_8720);
xor U8791 (N_8791,N_8708,N_8690);
and U8792 (N_8792,N_8678,N_8733);
and U8793 (N_8793,N_8655,N_8730);
and U8794 (N_8794,N_8630,N_8680);
and U8795 (N_8795,N_8629,N_8749);
or U8796 (N_8796,N_8711,N_8695);
and U8797 (N_8797,N_8668,N_8699);
or U8798 (N_8798,N_8700,N_8707);
or U8799 (N_8799,N_8670,N_8652);
and U8800 (N_8800,N_8662,N_8633);
nor U8801 (N_8801,N_8682,N_8687);
xnor U8802 (N_8802,N_8725,N_8626);
or U8803 (N_8803,N_8665,N_8663);
nor U8804 (N_8804,N_8698,N_8712);
and U8805 (N_8805,N_8745,N_8742);
xor U8806 (N_8806,N_8746,N_8647);
nand U8807 (N_8807,N_8676,N_8644);
or U8808 (N_8808,N_8641,N_8726);
xnor U8809 (N_8809,N_8638,N_8683);
and U8810 (N_8810,N_8715,N_8666);
nor U8811 (N_8811,N_8704,N_8747);
nor U8812 (N_8812,N_8649,N_8630);
and U8813 (N_8813,N_8640,N_8701);
nand U8814 (N_8814,N_8685,N_8687);
and U8815 (N_8815,N_8665,N_8673);
nor U8816 (N_8816,N_8681,N_8728);
or U8817 (N_8817,N_8699,N_8715);
nor U8818 (N_8818,N_8682,N_8706);
xnor U8819 (N_8819,N_8726,N_8651);
xor U8820 (N_8820,N_8631,N_8634);
xnor U8821 (N_8821,N_8746,N_8676);
xnor U8822 (N_8822,N_8719,N_8651);
xor U8823 (N_8823,N_8681,N_8645);
or U8824 (N_8824,N_8705,N_8637);
or U8825 (N_8825,N_8725,N_8746);
xor U8826 (N_8826,N_8680,N_8707);
and U8827 (N_8827,N_8733,N_8638);
and U8828 (N_8828,N_8646,N_8730);
or U8829 (N_8829,N_8740,N_8625);
nor U8830 (N_8830,N_8688,N_8737);
xor U8831 (N_8831,N_8680,N_8692);
or U8832 (N_8832,N_8721,N_8699);
nor U8833 (N_8833,N_8695,N_8665);
and U8834 (N_8834,N_8641,N_8735);
and U8835 (N_8835,N_8690,N_8749);
and U8836 (N_8836,N_8694,N_8676);
nand U8837 (N_8837,N_8628,N_8736);
and U8838 (N_8838,N_8678,N_8727);
and U8839 (N_8839,N_8666,N_8699);
xnor U8840 (N_8840,N_8658,N_8747);
and U8841 (N_8841,N_8629,N_8627);
nor U8842 (N_8842,N_8637,N_8708);
or U8843 (N_8843,N_8652,N_8711);
and U8844 (N_8844,N_8654,N_8681);
nor U8845 (N_8845,N_8680,N_8685);
nand U8846 (N_8846,N_8642,N_8647);
or U8847 (N_8847,N_8745,N_8704);
nand U8848 (N_8848,N_8692,N_8649);
or U8849 (N_8849,N_8743,N_8728);
nor U8850 (N_8850,N_8687,N_8678);
or U8851 (N_8851,N_8679,N_8659);
and U8852 (N_8852,N_8707,N_8649);
and U8853 (N_8853,N_8672,N_8679);
or U8854 (N_8854,N_8708,N_8744);
xnor U8855 (N_8855,N_8659,N_8692);
nand U8856 (N_8856,N_8735,N_8670);
nand U8857 (N_8857,N_8716,N_8677);
nor U8858 (N_8858,N_8702,N_8666);
or U8859 (N_8859,N_8662,N_8708);
and U8860 (N_8860,N_8649,N_8720);
or U8861 (N_8861,N_8723,N_8715);
nand U8862 (N_8862,N_8697,N_8690);
nor U8863 (N_8863,N_8647,N_8659);
nand U8864 (N_8864,N_8728,N_8633);
nand U8865 (N_8865,N_8636,N_8630);
and U8866 (N_8866,N_8738,N_8641);
or U8867 (N_8867,N_8690,N_8716);
xor U8868 (N_8868,N_8740,N_8656);
or U8869 (N_8869,N_8733,N_8735);
or U8870 (N_8870,N_8676,N_8695);
xor U8871 (N_8871,N_8720,N_8713);
xnor U8872 (N_8872,N_8706,N_8625);
nand U8873 (N_8873,N_8691,N_8670);
xnor U8874 (N_8874,N_8683,N_8710);
nor U8875 (N_8875,N_8796,N_8814);
or U8876 (N_8876,N_8791,N_8806);
nand U8877 (N_8877,N_8761,N_8837);
xnor U8878 (N_8878,N_8817,N_8823);
and U8879 (N_8879,N_8778,N_8789);
nand U8880 (N_8880,N_8861,N_8832);
nor U8881 (N_8881,N_8753,N_8781);
nand U8882 (N_8882,N_8838,N_8822);
and U8883 (N_8883,N_8805,N_8862);
or U8884 (N_8884,N_8760,N_8809);
nor U8885 (N_8885,N_8810,N_8775);
and U8886 (N_8886,N_8818,N_8850);
nor U8887 (N_8887,N_8820,N_8754);
xor U8888 (N_8888,N_8864,N_8839);
and U8889 (N_8889,N_8844,N_8854);
and U8890 (N_8890,N_8757,N_8851);
or U8891 (N_8891,N_8776,N_8849);
and U8892 (N_8892,N_8801,N_8858);
nor U8893 (N_8893,N_8859,N_8834);
nor U8894 (N_8894,N_8803,N_8774);
xnor U8895 (N_8895,N_8764,N_8765);
nand U8896 (N_8896,N_8779,N_8759);
or U8897 (N_8897,N_8797,N_8783);
nor U8898 (N_8898,N_8856,N_8786);
xnor U8899 (N_8899,N_8813,N_8867);
xor U8900 (N_8900,N_8768,N_8842);
nor U8901 (N_8901,N_8752,N_8827);
nand U8902 (N_8902,N_8784,N_8807);
and U8903 (N_8903,N_8835,N_8804);
nor U8904 (N_8904,N_8798,N_8865);
and U8905 (N_8905,N_8808,N_8770);
or U8906 (N_8906,N_8771,N_8762);
xor U8907 (N_8907,N_8785,N_8815);
and U8908 (N_8908,N_8763,N_8780);
or U8909 (N_8909,N_8866,N_8843);
or U8910 (N_8910,N_8872,N_8852);
and U8911 (N_8911,N_8799,N_8767);
nor U8912 (N_8912,N_8819,N_8845);
and U8913 (N_8913,N_8870,N_8829);
xor U8914 (N_8914,N_8869,N_8812);
or U8915 (N_8915,N_8795,N_8792);
or U8916 (N_8916,N_8816,N_8750);
or U8917 (N_8917,N_8830,N_8821);
or U8918 (N_8918,N_8840,N_8833);
and U8919 (N_8919,N_8868,N_8836);
nand U8920 (N_8920,N_8863,N_8848);
nor U8921 (N_8921,N_8755,N_8794);
nand U8922 (N_8922,N_8873,N_8788);
nand U8923 (N_8923,N_8825,N_8790);
or U8924 (N_8924,N_8811,N_8846);
nand U8925 (N_8925,N_8828,N_8857);
and U8926 (N_8926,N_8782,N_8841);
and U8927 (N_8927,N_8773,N_8853);
nor U8928 (N_8928,N_8777,N_8793);
or U8929 (N_8929,N_8826,N_8800);
nand U8930 (N_8930,N_8766,N_8847);
nor U8931 (N_8931,N_8824,N_8751);
xnor U8932 (N_8932,N_8860,N_8874);
and U8933 (N_8933,N_8831,N_8756);
nand U8934 (N_8934,N_8871,N_8769);
and U8935 (N_8935,N_8855,N_8787);
and U8936 (N_8936,N_8772,N_8758);
and U8937 (N_8937,N_8802,N_8760);
xor U8938 (N_8938,N_8831,N_8780);
and U8939 (N_8939,N_8758,N_8873);
or U8940 (N_8940,N_8819,N_8764);
nand U8941 (N_8941,N_8872,N_8791);
and U8942 (N_8942,N_8804,N_8765);
xnor U8943 (N_8943,N_8867,N_8816);
or U8944 (N_8944,N_8797,N_8820);
nor U8945 (N_8945,N_8765,N_8809);
nand U8946 (N_8946,N_8874,N_8811);
or U8947 (N_8947,N_8753,N_8774);
or U8948 (N_8948,N_8851,N_8758);
nor U8949 (N_8949,N_8843,N_8783);
or U8950 (N_8950,N_8830,N_8858);
or U8951 (N_8951,N_8863,N_8874);
and U8952 (N_8952,N_8781,N_8818);
and U8953 (N_8953,N_8874,N_8826);
and U8954 (N_8954,N_8770,N_8768);
and U8955 (N_8955,N_8761,N_8849);
nor U8956 (N_8956,N_8752,N_8842);
nand U8957 (N_8957,N_8846,N_8802);
or U8958 (N_8958,N_8774,N_8788);
nand U8959 (N_8959,N_8870,N_8831);
nor U8960 (N_8960,N_8863,N_8790);
or U8961 (N_8961,N_8833,N_8816);
nor U8962 (N_8962,N_8754,N_8843);
and U8963 (N_8963,N_8837,N_8790);
nand U8964 (N_8964,N_8817,N_8842);
nor U8965 (N_8965,N_8818,N_8809);
and U8966 (N_8966,N_8847,N_8763);
nor U8967 (N_8967,N_8863,N_8858);
and U8968 (N_8968,N_8821,N_8817);
nor U8969 (N_8969,N_8791,N_8759);
nand U8970 (N_8970,N_8777,N_8769);
or U8971 (N_8971,N_8818,N_8860);
and U8972 (N_8972,N_8787,N_8829);
or U8973 (N_8973,N_8870,N_8756);
xor U8974 (N_8974,N_8774,N_8797);
nor U8975 (N_8975,N_8841,N_8852);
or U8976 (N_8976,N_8819,N_8851);
and U8977 (N_8977,N_8836,N_8778);
or U8978 (N_8978,N_8850,N_8822);
or U8979 (N_8979,N_8762,N_8823);
xor U8980 (N_8980,N_8873,N_8791);
and U8981 (N_8981,N_8814,N_8872);
nor U8982 (N_8982,N_8874,N_8845);
nand U8983 (N_8983,N_8828,N_8812);
and U8984 (N_8984,N_8778,N_8846);
xnor U8985 (N_8985,N_8784,N_8787);
nor U8986 (N_8986,N_8755,N_8776);
xor U8987 (N_8987,N_8753,N_8831);
or U8988 (N_8988,N_8778,N_8768);
and U8989 (N_8989,N_8758,N_8871);
xor U8990 (N_8990,N_8778,N_8818);
xnor U8991 (N_8991,N_8865,N_8815);
xor U8992 (N_8992,N_8873,N_8854);
nand U8993 (N_8993,N_8812,N_8786);
nand U8994 (N_8994,N_8860,N_8866);
nor U8995 (N_8995,N_8778,N_8773);
nand U8996 (N_8996,N_8827,N_8756);
nor U8997 (N_8997,N_8751,N_8757);
nand U8998 (N_8998,N_8767,N_8795);
nor U8999 (N_8999,N_8770,N_8818);
nand U9000 (N_9000,N_8899,N_8906);
nor U9001 (N_9001,N_8971,N_8957);
nor U9002 (N_9002,N_8892,N_8967);
nand U9003 (N_9003,N_8919,N_8909);
or U9004 (N_9004,N_8953,N_8915);
or U9005 (N_9005,N_8960,N_8897);
xnor U9006 (N_9006,N_8962,N_8879);
or U9007 (N_9007,N_8894,N_8961);
nand U9008 (N_9008,N_8969,N_8956);
and U9009 (N_9009,N_8937,N_8977);
nand U9010 (N_9010,N_8941,N_8930);
and U9011 (N_9011,N_8889,N_8951);
xnor U9012 (N_9012,N_8954,N_8947);
and U9013 (N_9013,N_8935,N_8997);
or U9014 (N_9014,N_8890,N_8938);
nand U9015 (N_9015,N_8986,N_8900);
and U9016 (N_9016,N_8989,N_8907);
nand U9017 (N_9017,N_8995,N_8904);
and U9018 (N_9018,N_8917,N_8931);
or U9019 (N_9019,N_8985,N_8928);
xor U9020 (N_9020,N_8885,N_8981);
xor U9021 (N_9021,N_8948,N_8875);
xor U9022 (N_9022,N_8877,N_8910);
or U9023 (N_9023,N_8911,N_8987);
xor U9024 (N_9024,N_8946,N_8896);
or U9025 (N_9025,N_8992,N_8998);
and U9026 (N_9026,N_8993,N_8955);
xor U9027 (N_9027,N_8925,N_8940);
nand U9028 (N_9028,N_8942,N_8983);
xor U9029 (N_9029,N_8999,N_8936);
nand U9030 (N_9030,N_8945,N_8918);
and U9031 (N_9031,N_8878,N_8923);
or U9032 (N_9032,N_8965,N_8884);
nand U9033 (N_9033,N_8994,N_8891);
and U9034 (N_9034,N_8881,N_8933);
or U9035 (N_9035,N_8929,N_8883);
and U9036 (N_9036,N_8876,N_8927);
or U9037 (N_9037,N_8914,N_8982);
and U9038 (N_9038,N_8979,N_8916);
or U9039 (N_9039,N_8950,N_8880);
or U9040 (N_9040,N_8990,N_8973);
xor U9041 (N_9041,N_8966,N_8975);
xor U9042 (N_9042,N_8978,N_8959);
nand U9043 (N_9043,N_8924,N_8952);
xnor U9044 (N_9044,N_8903,N_8920);
xor U9045 (N_9045,N_8912,N_8980);
or U9046 (N_9046,N_8939,N_8949);
nor U9047 (N_9047,N_8964,N_8963);
nand U9048 (N_9048,N_8943,N_8988);
xnor U9049 (N_9049,N_8976,N_8913);
or U9050 (N_9050,N_8902,N_8972);
or U9051 (N_9051,N_8984,N_8898);
nand U9052 (N_9052,N_8895,N_8974);
or U9053 (N_9053,N_8921,N_8996);
and U9054 (N_9054,N_8893,N_8886);
and U9055 (N_9055,N_8958,N_8887);
or U9056 (N_9056,N_8932,N_8934);
nor U9057 (N_9057,N_8922,N_8968);
and U9058 (N_9058,N_8905,N_8901);
or U9059 (N_9059,N_8944,N_8991);
nand U9060 (N_9060,N_8882,N_8970);
xor U9061 (N_9061,N_8908,N_8926);
or U9062 (N_9062,N_8888,N_8968);
and U9063 (N_9063,N_8886,N_8965);
nor U9064 (N_9064,N_8888,N_8889);
nand U9065 (N_9065,N_8900,N_8961);
and U9066 (N_9066,N_8910,N_8957);
xor U9067 (N_9067,N_8914,N_8991);
nor U9068 (N_9068,N_8934,N_8930);
xnor U9069 (N_9069,N_8884,N_8901);
xor U9070 (N_9070,N_8976,N_8929);
or U9071 (N_9071,N_8971,N_8964);
and U9072 (N_9072,N_8944,N_8883);
or U9073 (N_9073,N_8891,N_8888);
and U9074 (N_9074,N_8954,N_8929);
nand U9075 (N_9075,N_8893,N_8972);
and U9076 (N_9076,N_8971,N_8893);
xor U9077 (N_9077,N_8879,N_8948);
or U9078 (N_9078,N_8919,N_8927);
and U9079 (N_9079,N_8909,N_8936);
or U9080 (N_9080,N_8913,N_8877);
nand U9081 (N_9081,N_8890,N_8945);
and U9082 (N_9082,N_8958,N_8895);
xnor U9083 (N_9083,N_8942,N_8966);
and U9084 (N_9084,N_8914,N_8936);
and U9085 (N_9085,N_8923,N_8922);
nor U9086 (N_9086,N_8886,N_8929);
or U9087 (N_9087,N_8891,N_8903);
xnor U9088 (N_9088,N_8949,N_8914);
xnor U9089 (N_9089,N_8905,N_8893);
or U9090 (N_9090,N_8905,N_8969);
xor U9091 (N_9091,N_8880,N_8885);
xor U9092 (N_9092,N_8981,N_8884);
nand U9093 (N_9093,N_8913,N_8927);
nor U9094 (N_9094,N_8900,N_8960);
or U9095 (N_9095,N_8883,N_8922);
or U9096 (N_9096,N_8891,N_8922);
nand U9097 (N_9097,N_8981,N_8907);
or U9098 (N_9098,N_8956,N_8915);
nor U9099 (N_9099,N_8916,N_8935);
nand U9100 (N_9100,N_8914,N_8878);
and U9101 (N_9101,N_8880,N_8939);
and U9102 (N_9102,N_8940,N_8893);
nand U9103 (N_9103,N_8945,N_8885);
or U9104 (N_9104,N_8965,N_8934);
nor U9105 (N_9105,N_8965,N_8960);
nor U9106 (N_9106,N_8965,N_8926);
or U9107 (N_9107,N_8930,N_8917);
or U9108 (N_9108,N_8888,N_8950);
nor U9109 (N_9109,N_8905,N_8955);
xor U9110 (N_9110,N_8935,N_8949);
xnor U9111 (N_9111,N_8967,N_8931);
or U9112 (N_9112,N_8973,N_8946);
xnor U9113 (N_9113,N_8999,N_8986);
and U9114 (N_9114,N_8924,N_8898);
and U9115 (N_9115,N_8983,N_8929);
xnor U9116 (N_9116,N_8956,N_8925);
and U9117 (N_9117,N_8961,N_8926);
or U9118 (N_9118,N_8887,N_8886);
xnor U9119 (N_9119,N_8938,N_8907);
nor U9120 (N_9120,N_8994,N_8995);
nand U9121 (N_9121,N_8917,N_8932);
nand U9122 (N_9122,N_8937,N_8916);
xnor U9123 (N_9123,N_8901,N_8968);
and U9124 (N_9124,N_8940,N_8916);
nand U9125 (N_9125,N_9084,N_9116);
or U9126 (N_9126,N_9024,N_9112);
and U9127 (N_9127,N_9089,N_9053);
or U9128 (N_9128,N_9006,N_9058);
nand U9129 (N_9129,N_9030,N_9088);
nor U9130 (N_9130,N_9079,N_9097);
and U9131 (N_9131,N_9062,N_9080);
and U9132 (N_9132,N_9044,N_9020);
or U9133 (N_9133,N_9073,N_9121);
nand U9134 (N_9134,N_9048,N_9105);
nand U9135 (N_9135,N_9110,N_9122);
xor U9136 (N_9136,N_9066,N_9119);
or U9137 (N_9137,N_9047,N_9081);
or U9138 (N_9138,N_9077,N_9094);
xor U9139 (N_9139,N_9106,N_9007);
and U9140 (N_9140,N_9015,N_9017);
and U9141 (N_9141,N_9046,N_9001);
and U9142 (N_9142,N_9018,N_9032);
xor U9143 (N_9143,N_9102,N_9108);
nor U9144 (N_9144,N_9010,N_9035);
xor U9145 (N_9145,N_9107,N_9064);
nand U9146 (N_9146,N_9123,N_9042);
and U9147 (N_9147,N_9114,N_9031);
nor U9148 (N_9148,N_9022,N_9099);
and U9149 (N_9149,N_9011,N_9041);
nand U9150 (N_9150,N_9072,N_9085);
or U9151 (N_9151,N_9040,N_9019);
xnor U9152 (N_9152,N_9023,N_9016);
nor U9153 (N_9153,N_9009,N_9027);
nor U9154 (N_9154,N_9067,N_9060);
nand U9155 (N_9155,N_9039,N_9091);
nand U9156 (N_9156,N_9050,N_9059);
nor U9157 (N_9157,N_9075,N_9095);
and U9158 (N_9158,N_9096,N_9005);
and U9159 (N_9159,N_9093,N_9029);
xor U9160 (N_9160,N_9120,N_9056);
xor U9161 (N_9161,N_9071,N_9003);
and U9162 (N_9162,N_9098,N_9082);
and U9163 (N_9163,N_9100,N_9124);
nor U9164 (N_9164,N_9013,N_9045);
nand U9165 (N_9165,N_9008,N_9086);
xnor U9166 (N_9166,N_9068,N_9090);
xor U9167 (N_9167,N_9036,N_9026);
xor U9168 (N_9168,N_9087,N_9002);
or U9169 (N_9169,N_9061,N_9063);
nor U9170 (N_9170,N_9000,N_9101);
nand U9171 (N_9171,N_9070,N_9115);
nand U9172 (N_9172,N_9076,N_9038);
xor U9173 (N_9173,N_9118,N_9021);
nor U9174 (N_9174,N_9012,N_9037);
xnor U9175 (N_9175,N_9074,N_9014);
nor U9176 (N_9176,N_9103,N_9092);
or U9177 (N_9177,N_9057,N_9117);
and U9178 (N_9178,N_9028,N_9055);
nor U9179 (N_9179,N_9083,N_9109);
and U9180 (N_9180,N_9043,N_9049);
nor U9181 (N_9181,N_9004,N_9034);
nor U9182 (N_9182,N_9078,N_9054);
xnor U9183 (N_9183,N_9033,N_9111);
xor U9184 (N_9184,N_9051,N_9069);
and U9185 (N_9185,N_9052,N_9065);
xor U9186 (N_9186,N_9104,N_9025);
or U9187 (N_9187,N_9113,N_9030);
nor U9188 (N_9188,N_9019,N_9042);
and U9189 (N_9189,N_9042,N_9002);
or U9190 (N_9190,N_9066,N_9004);
xor U9191 (N_9191,N_9007,N_9054);
xnor U9192 (N_9192,N_9060,N_9038);
nand U9193 (N_9193,N_9036,N_9112);
and U9194 (N_9194,N_9075,N_9070);
nand U9195 (N_9195,N_9013,N_9010);
or U9196 (N_9196,N_9089,N_9034);
nor U9197 (N_9197,N_9004,N_9067);
and U9198 (N_9198,N_9092,N_9078);
and U9199 (N_9199,N_9001,N_9107);
and U9200 (N_9200,N_9018,N_9014);
or U9201 (N_9201,N_9057,N_9071);
and U9202 (N_9202,N_9014,N_9094);
xor U9203 (N_9203,N_9067,N_9014);
xnor U9204 (N_9204,N_9087,N_9048);
and U9205 (N_9205,N_9010,N_9102);
nand U9206 (N_9206,N_9057,N_9124);
and U9207 (N_9207,N_9075,N_9042);
nand U9208 (N_9208,N_9067,N_9093);
nor U9209 (N_9209,N_9075,N_9019);
nand U9210 (N_9210,N_9002,N_9031);
xnor U9211 (N_9211,N_9015,N_9045);
and U9212 (N_9212,N_9060,N_9119);
or U9213 (N_9213,N_9087,N_9084);
and U9214 (N_9214,N_9047,N_9010);
and U9215 (N_9215,N_9020,N_9024);
and U9216 (N_9216,N_9078,N_9014);
and U9217 (N_9217,N_9082,N_9089);
or U9218 (N_9218,N_9066,N_9005);
and U9219 (N_9219,N_9117,N_9010);
xor U9220 (N_9220,N_9106,N_9011);
or U9221 (N_9221,N_9025,N_9096);
and U9222 (N_9222,N_9070,N_9065);
or U9223 (N_9223,N_9081,N_9026);
and U9224 (N_9224,N_9002,N_9034);
nand U9225 (N_9225,N_9069,N_9092);
nor U9226 (N_9226,N_9008,N_9017);
and U9227 (N_9227,N_9089,N_9116);
nand U9228 (N_9228,N_9035,N_9058);
or U9229 (N_9229,N_9061,N_9105);
and U9230 (N_9230,N_9086,N_9047);
xor U9231 (N_9231,N_9033,N_9116);
xor U9232 (N_9232,N_9069,N_9008);
nor U9233 (N_9233,N_9026,N_9009);
and U9234 (N_9234,N_9084,N_9086);
nor U9235 (N_9235,N_9059,N_9077);
nand U9236 (N_9236,N_9032,N_9037);
or U9237 (N_9237,N_9072,N_9053);
and U9238 (N_9238,N_9018,N_9109);
nor U9239 (N_9239,N_9068,N_9073);
or U9240 (N_9240,N_9069,N_9085);
nand U9241 (N_9241,N_9025,N_9052);
or U9242 (N_9242,N_9089,N_9016);
nor U9243 (N_9243,N_9080,N_9060);
nor U9244 (N_9244,N_9084,N_9092);
nand U9245 (N_9245,N_9098,N_9000);
nor U9246 (N_9246,N_9098,N_9075);
and U9247 (N_9247,N_9099,N_9020);
nand U9248 (N_9248,N_9078,N_9116);
and U9249 (N_9249,N_9047,N_9025);
or U9250 (N_9250,N_9140,N_9163);
nor U9251 (N_9251,N_9218,N_9200);
xor U9252 (N_9252,N_9168,N_9188);
and U9253 (N_9253,N_9205,N_9247);
or U9254 (N_9254,N_9177,N_9225);
or U9255 (N_9255,N_9142,N_9182);
nor U9256 (N_9256,N_9212,N_9241);
nand U9257 (N_9257,N_9244,N_9207);
and U9258 (N_9258,N_9175,N_9153);
or U9259 (N_9259,N_9176,N_9125);
nand U9260 (N_9260,N_9210,N_9185);
nor U9261 (N_9261,N_9221,N_9230);
xnor U9262 (N_9262,N_9211,N_9136);
and U9263 (N_9263,N_9186,N_9228);
or U9264 (N_9264,N_9242,N_9137);
xor U9265 (N_9265,N_9170,N_9224);
and U9266 (N_9266,N_9158,N_9239);
nor U9267 (N_9267,N_9130,N_9198);
xor U9268 (N_9268,N_9223,N_9203);
nand U9269 (N_9269,N_9214,N_9246);
nor U9270 (N_9270,N_9245,N_9189);
and U9271 (N_9271,N_9161,N_9159);
and U9272 (N_9272,N_9193,N_9184);
xnor U9273 (N_9273,N_9248,N_9169);
nor U9274 (N_9274,N_9236,N_9166);
and U9275 (N_9275,N_9147,N_9178);
or U9276 (N_9276,N_9172,N_9209);
nor U9277 (N_9277,N_9148,N_9199);
or U9278 (N_9278,N_9206,N_9173);
and U9279 (N_9279,N_9139,N_9227);
or U9280 (N_9280,N_9165,N_9249);
nand U9281 (N_9281,N_9160,N_9233);
and U9282 (N_9282,N_9216,N_9171);
xnor U9283 (N_9283,N_9197,N_9195);
and U9284 (N_9284,N_9126,N_9167);
and U9285 (N_9285,N_9192,N_9141);
xnor U9286 (N_9286,N_9129,N_9149);
or U9287 (N_9287,N_9155,N_9131);
nor U9288 (N_9288,N_9164,N_9143);
nand U9289 (N_9289,N_9133,N_9179);
or U9290 (N_9290,N_9243,N_9181);
and U9291 (N_9291,N_9235,N_9240);
or U9292 (N_9292,N_9146,N_9231);
xor U9293 (N_9293,N_9157,N_9187);
nor U9294 (N_9294,N_9220,N_9190);
and U9295 (N_9295,N_9196,N_9204);
and U9296 (N_9296,N_9150,N_9201);
nor U9297 (N_9297,N_9132,N_9202);
and U9298 (N_9298,N_9156,N_9151);
nand U9299 (N_9299,N_9217,N_9138);
and U9300 (N_9300,N_9219,N_9194);
or U9301 (N_9301,N_9180,N_9183);
and U9302 (N_9302,N_9215,N_9232);
nor U9303 (N_9303,N_9237,N_9152);
nand U9304 (N_9304,N_9229,N_9144);
and U9305 (N_9305,N_9222,N_9145);
nor U9306 (N_9306,N_9174,N_9154);
xnor U9307 (N_9307,N_9191,N_9128);
or U9308 (N_9308,N_9213,N_9226);
nor U9309 (N_9309,N_9234,N_9162);
and U9310 (N_9310,N_9127,N_9134);
and U9311 (N_9311,N_9208,N_9135);
nor U9312 (N_9312,N_9238,N_9164);
or U9313 (N_9313,N_9216,N_9166);
or U9314 (N_9314,N_9237,N_9193);
nand U9315 (N_9315,N_9246,N_9127);
and U9316 (N_9316,N_9157,N_9198);
xor U9317 (N_9317,N_9217,N_9193);
and U9318 (N_9318,N_9130,N_9144);
and U9319 (N_9319,N_9206,N_9170);
xnor U9320 (N_9320,N_9144,N_9242);
nand U9321 (N_9321,N_9224,N_9184);
xnor U9322 (N_9322,N_9245,N_9141);
or U9323 (N_9323,N_9225,N_9211);
xnor U9324 (N_9324,N_9140,N_9153);
nand U9325 (N_9325,N_9149,N_9164);
nand U9326 (N_9326,N_9245,N_9204);
nand U9327 (N_9327,N_9187,N_9246);
xor U9328 (N_9328,N_9136,N_9128);
or U9329 (N_9329,N_9152,N_9249);
xnor U9330 (N_9330,N_9215,N_9187);
nor U9331 (N_9331,N_9136,N_9224);
nor U9332 (N_9332,N_9235,N_9177);
nor U9333 (N_9333,N_9131,N_9154);
and U9334 (N_9334,N_9238,N_9236);
nor U9335 (N_9335,N_9148,N_9184);
and U9336 (N_9336,N_9133,N_9172);
or U9337 (N_9337,N_9177,N_9242);
xnor U9338 (N_9338,N_9131,N_9192);
nor U9339 (N_9339,N_9211,N_9197);
or U9340 (N_9340,N_9160,N_9140);
nand U9341 (N_9341,N_9178,N_9135);
or U9342 (N_9342,N_9172,N_9147);
nor U9343 (N_9343,N_9142,N_9172);
nor U9344 (N_9344,N_9180,N_9162);
nand U9345 (N_9345,N_9130,N_9194);
and U9346 (N_9346,N_9184,N_9164);
nand U9347 (N_9347,N_9147,N_9225);
nor U9348 (N_9348,N_9229,N_9241);
and U9349 (N_9349,N_9169,N_9192);
nor U9350 (N_9350,N_9200,N_9130);
nor U9351 (N_9351,N_9131,N_9167);
nor U9352 (N_9352,N_9128,N_9240);
or U9353 (N_9353,N_9140,N_9169);
or U9354 (N_9354,N_9225,N_9239);
or U9355 (N_9355,N_9244,N_9167);
and U9356 (N_9356,N_9246,N_9140);
nor U9357 (N_9357,N_9216,N_9237);
xor U9358 (N_9358,N_9221,N_9132);
and U9359 (N_9359,N_9173,N_9204);
nor U9360 (N_9360,N_9198,N_9177);
or U9361 (N_9361,N_9207,N_9144);
or U9362 (N_9362,N_9209,N_9219);
or U9363 (N_9363,N_9174,N_9185);
or U9364 (N_9364,N_9234,N_9212);
or U9365 (N_9365,N_9139,N_9229);
nand U9366 (N_9366,N_9219,N_9237);
nor U9367 (N_9367,N_9146,N_9249);
or U9368 (N_9368,N_9235,N_9186);
xor U9369 (N_9369,N_9208,N_9245);
nand U9370 (N_9370,N_9204,N_9155);
nor U9371 (N_9371,N_9204,N_9161);
and U9372 (N_9372,N_9128,N_9147);
xnor U9373 (N_9373,N_9233,N_9125);
or U9374 (N_9374,N_9159,N_9204);
and U9375 (N_9375,N_9275,N_9257);
nand U9376 (N_9376,N_9294,N_9251);
nor U9377 (N_9377,N_9293,N_9253);
nand U9378 (N_9378,N_9357,N_9324);
xor U9379 (N_9379,N_9301,N_9288);
xnor U9380 (N_9380,N_9366,N_9323);
xor U9381 (N_9381,N_9363,N_9254);
and U9382 (N_9382,N_9278,N_9259);
and U9383 (N_9383,N_9312,N_9277);
nand U9384 (N_9384,N_9348,N_9285);
xnor U9385 (N_9385,N_9269,N_9341);
or U9386 (N_9386,N_9373,N_9307);
nor U9387 (N_9387,N_9315,N_9308);
or U9388 (N_9388,N_9252,N_9276);
nor U9389 (N_9389,N_9317,N_9267);
and U9390 (N_9390,N_9271,N_9347);
nor U9391 (N_9391,N_9302,N_9329);
nor U9392 (N_9392,N_9361,N_9325);
xor U9393 (N_9393,N_9292,N_9371);
and U9394 (N_9394,N_9356,N_9295);
nand U9395 (N_9395,N_9343,N_9334);
and U9396 (N_9396,N_9313,N_9328);
or U9397 (N_9397,N_9352,N_9320);
xor U9398 (N_9398,N_9309,N_9330);
nor U9399 (N_9399,N_9338,N_9296);
nor U9400 (N_9400,N_9369,N_9322);
and U9401 (N_9401,N_9346,N_9284);
nor U9402 (N_9402,N_9300,N_9306);
xnor U9403 (N_9403,N_9368,N_9256);
nor U9404 (N_9404,N_9290,N_9342);
xnor U9405 (N_9405,N_9281,N_9298);
and U9406 (N_9406,N_9266,N_9349);
and U9407 (N_9407,N_9333,N_9274);
nor U9408 (N_9408,N_9250,N_9297);
nor U9409 (N_9409,N_9310,N_9344);
nand U9410 (N_9410,N_9283,N_9316);
nand U9411 (N_9411,N_9289,N_9305);
nor U9412 (N_9412,N_9364,N_9258);
nand U9413 (N_9413,N_9270,N_9314);
nor U9414 (N_9414,N_9265,N_9358);
nor U9415 (N_9415,N_9370,N_9365);
nor U9416 (N_9416,N_9279,N_9304);
nand U9417 (N_9417,N_9345,N_9282);
or U9418 (N_9418,N_9299,N_9351);
and U9419 (N_9419,N_9339,N_9260);
and U9420 (N_9420,N_9272,N_9362);
xnor U9421 (N_9421,N_9340,N_9255);
nor U9422 (N_9422,N_9321,N_9264);
or U9423 (N_9423,N_9367,N_9268);
or U9424 (N_9424,N_9350,N_9359);
or U9425 (N_9425,N_9291,N_9319);
or U9426 (N_9426,N_9273,N_9327);
and U9427 (N_9427,N_9335,N_9354);
or U9428 (N_9428,N_9355,N_9336);
or U9429 (N_9429,N_9318,N_9286);
nor U9430 (N_9430,N_9353,N_9287);
xor U9431 (N_9431,N_9261,N_9372);
and U9432 (N_9432,N_9360,N_9332);
xnor U9433 (N_9433,N_9326,N_9311);
nor U9434 (N_9434,N_9331,N_9303);
xor U9435 (N_9435,N_9374,N_9337);
or U9436 (N_9436,N_9262,N_9263);
nor U9437 (N_9437,N_9280,N_9328);
nor U9438 (N_9438,N_9315,N_9362);
nand U9439 (N_9439,N_9370,N_9311);
nand U9440 (N_9440,N_9346,N_9283);
or U9441 (N_9441,N_9319,N_9325);
nor U9442 (N_9442,N_9273,N_9304);
xnor U9443 (N_9443,N_9371,N_9357);
nor U9444 (N_9444,N_9368,N_9312);
and U9445 (N_9445,N_9307,N_9299);
nand U9446 (N_9446,N_9311,N_9372);
nand U9447 (N_9447,N_9287,N_9273);
nand U9448 (N_9448,N_9304,N_9297);
or U9449 (N_9449,N_9295,N_9302);
or U9450 (N_9450,N_9316,N_9310);
nand U9451 (N_9451,N_9325,N_9311);
nand U9452 (N_9452,N_9327,N_9325);
nor U9453 (N_9453,N_9263,N_9354);
xor U9454 (N_9454,N_9301,N_9285);
nand U9455 (N_9455,N_9264,N_9369);
nor U9456 (N_9456,N_9294,N_9307);
nor U9457 (N_9457,N_9308,N_9312);
nor U9458 (N_9458,N_9254,N_9257);
and U9459 (N_9459,N_9265,N_9344);
nor U9460 (N_9460,N_9267,N_9370);
nand U9461 (N_9461,N_9364,N_9263);
nor U9462 (N_9462,N_9260,N_9262);
nand U9463 (N_9463,N_9283,N_9303);
nand U9464 (N_9464,N_9260,N_9361);
and U9465 (N_9465,N_9331,N_9374);
xnor U9466 (N_9466,N_9292,N_9325);
nor U9467 (N_9467,N_9330,N_9372);
nor U9468 (N_9468,N_9320,N_9343);
xnor U9469 (N_9469,N_9342,N_9338);
or U9470 (N_9470,N_9360,N_9367);
nand U9471 (N_9471,N_9259,N_9279);
xor U9472 (N_9472,N_9260,N_9340);
and U9473 (N_9473,N_9287,N_9310);
nand U9474 (N_9474,N_9365,N_9367);
nor U9475 (N_9475,N_9283,N_9251);
and U9476 (N_9476,N_9359,N_9291);
nor U9477 (N_9477,N_9322,N_9339);
or U9478 (N_9478,N_9311,N_9352);
nand U9479 (N_9479,N_9351,N_9264);
nor U9480 (N_9480,N_9309,N_9275);
nand U9481 (N_9481,N_9349,N_9252);
and U9482 (N_9482,N_9305,N_9354);
or U9483 (N_9483,N_9332,N_9374);
nand U9484 (N_9484,N_9254,N_9361);
xor U9485 (N_9485,N_9279,N_9289);
nand U9486 (N_9486,N_9288,N_9337);
xor U9487 (N_9487,N_9295,N_9285);
xnor U9488 (N_9488,N_9252,N_9312);
or U9489 (N_9489,N_9320,N_9370);
or U9490 (N_9490,N_9314,N_9348);
and U9491 (N_9491,N_9326,N_9317);
xnor U9492 (N_9492,N_9291,N_9320);
nand U9493 (N_9493,N_9277,N_9296);
and U9494 (N_9494,N_9292,N_9369);
nand U9495 (N_9495,N_9254,N_9311);
and U9496 (N_9496,N_9330,N_9326);
and U9497 (N_9497,N_9361,N_9267);
xnor U9498 (N_9498,N_9301,N_9334);
xor U9499 (N_9499,N_9326,N_9319);
nand U9500 (N_9500,N_9392,N_9460);
and U9501 (N_9501,N_9411,N_9497);
and U9502 (N_9502,N_9453,N_9480);
nor U9503 (N_9503,N_9389,N_9386);
xor U9504 (N_9504,N_9398,N_9408);
xor U9505 (N_9505,N_9462,N_9491);
nand U9506 (N_9506,N_9397,N_9452);
xnor U9507 (N_9507,N_9481,N_9484);
or U9508 (N_9508,N_9387,N_9454);
xnor U9509 (N_9509,N_9432,N_9384);
and U9510 (N_9510,N_9383,N_9416);
xnor U9511 (N_9511,N_9475,N_9494);
xnor U9512 (N_9512,N_9378,N_9412);
xor U9513 (N_9513,N_9464,N_9492);
and U9514 (N_9514,N_9451,N_9424);
or U9515 (N_9515,N_9466,N_9434);
or U9516 (N_9516,N_9393,N_9425);
and U9517 (N_9517,N_9449,N_9465);
or U9518 (N_9518,N_9470,N_9382);
nand U9519 (N_9519,N_9380,N_9489);
xnor U9520 (N_9520,N_9485,N_9429);
xnor U9521 (N_9521,N_9455,N_9450);
xnor U9522 (N_9522,N_9396,N_9433);
or U9523 (N_9523,N_9446,N_9423);
xor U9524 (N_9524,N_9391,N_9395);
nor U9525 (N_9525,N_9456,N_9413);
and U9526 (N_9526,N_9415,N_9376);
and U9527 (N_9527,N_9459,N_9410);
and U9528 (N_9528,N_9390,N_9473);
nand U9529 (N_9529,N_9399,N_9468);
nor U9530 (N_9530,N_9404,N_9379);
nand U9531 (N_9531,N_9388,N_9405);
nor U9532 (N_9532,N_9439,N_9377);
nand U9533 (N_9533,N_9463,N_9417);
and U9534 (N_9534,N_9483,N_9422);
and U9535 (N_9535,N_9486,N_9487);
nand U9536 (N_9536,N_9385,N_9445);
or U9537 (N_9537,N_9442,N_9472);
nor U9538 (N_9538,N_9447,N_9407);
and U9539 (N_9539,N_9381,N_9419);
xor U9540 (N_9540,N_9498,N_9437);
nand U9541 (N_9541,N_9409,N_9426);
nand U9542 (N_9542,N_9474,N_9495);
nor U9543 (N_9543,N_9428,N_9414);
nand U9544 (N_9544,N_9431,N_9394);
or U9545 (N_9545,N_9421,N_9493);
nor U9546 (N_9546,N_9469,N_9427);
xnor U9547 (N_9547,N_9458,N_9479);
and U9548 (N_9548,N_9418,N_9482);
or U9549 (N_9549,N_9488,N_9435);
or U9550 (N_9550,N_9467,N_9436);
nand U9551 (N_9551,N_9441,N_9420);
nor U9552 (N_9552,N_9478,N_9476);
and U9553 (N_9553,N_9403,N_9499);
nand U9554 (N_9554,N_9406,N_9443);
nand U9555 (N_9555,N_9490,N_9457);
xor U9556 (N_9556,N_9440,N_9448);
xnor U9557 (N_9557,N_9400,N_9430);
and U9558 (N_9558,N_9444,N_9438);
xnor U9559 (N_9559,N_9401,N_9461);
nand U9560 (N_9560,N_9471,N_9477);
nor U9561 (N_9561,N_9375,N_9496);
and U9562 (N_9562,N_9402,N_9463);
nor U9563 (N_9563,N_9390,N_9469);
or U9564 (N_9564,N_9412,N_9433);
or U9565 (N_9565,N_9432,N_9389);
and U9566 (N_9566,N_9490,N_9484);
nand U9567 (N_9567,N_9476,N_9394);
nor U9568 (N_9568,N_9410,N_9490);
and U9569 (N_9569,N_9414,N_9390);
or U9570 (N_9570,N_9459,N_9392);
xor U9571 (N_9571,N_9400,N_9486);
or U9572 (N_9572,N_9458,N_9404);
and U9573 (N_9573,N_9474,N_9381);
nand U9574 (N_9574,N_9451,N_9397);
or U9575 (N_9575,N_9488,N_9400);
or U9576 (N_9576,N_9493,N_9471);
nor U9577 (N_9577,N_9417,N_9410);
xor U9578 (N_9578,N_9384,N_9394);
or U9579 (N_9579,N_9481,N_9447);
nand U9580 (N_9580,N_9407,N_9498);
nand U9581 (N_9581,N_9412,N_9410);
nor U9582 (N_9582,N_9443,N_9384);
nand U9583 (N_9583,N_9499,N_9434);
or U9584 (N_9584,N_9461,N_9441);
and U9585 (N_9585,N_9491,N_9446);
nand U9586 (N_9586,N_9405,N_9436);
nand U9587 (N_9587,N_9402,N_9468);
xnor U9588 (N_9588,N_9383,N_9396);
and U9589 (N_9589,N_9457,N_9439);
nor U9590 (N_9590,N_9461,N_9386);
or U9591 (N_9591,N_9490,N_9486);
nand U9592 (N_9592,N_9444,N_9383);
nand U9593 (N_9593,N_9391,N_9464);
xor U9594 (N_9594,N_9457,N_9485);
or U9595 (N_9595,N_9408,N_9421);
xor U9596 (N_9596,N_9408,N_9457);
or U9597 (N_9597,N_9381,N_9406);
nor U9598 (N_9598,N_9438,N_9443);
or U9599 (N_9599,N_9451,N_9442);
xor U9600 (N_9600,N_9484,N_9496);
xor U9601 (N_9601,N_9431,N_9452);
nor U9602 (N_9602,N_9439,N_9451);
and U9603 (N_9603,N_9442,N_9487);
or U9604 (N_9604,N_9496,N_9420);
and U9605 (N_9605,N_9382,N_9473);
nor U9606 (N_9606,N_9444,N_9388);
nor U9607 (N_9607,N_9375,N_9493);
or U9608 (N_9608,N_9454,N_9458);
nor U9609 (N_9609,N_9427,N_9384);
and U9610 (N_9610,N_9415,N_9446);
xnor U9611 (N_9611,N_9453,N_9433);
and U9612 (N_9612,N_9499,N_9404);
nor U9613 (N_9613,N_9376,N_9385);
and U9614 (N_9614,N_9433,N_9375);
nand U9615 (N_9615,N_9388,N_9384);
nor U9616 (N_9616,N_9495,N_9382);
or U9617 (N_9617,N_9394,N_9442);
or U9618 (N_9618,N_9468,N_9384);
and U9619 (N_9619,N_9461,N_9483);
nand U9620 (N_9620,N_9493,N_9409);
xnor U9621 (N_9621,N_9440,N_9386);
or U9622 (N_9622,N_9411,N_9478);
or U9623 (N_9623,N_9469,N_9424);
or U9624 (N_9624,N_9393,N_9470);
xnor U9625 (N_9625,N_9582,N_9580);
xnor U9626 (N_9626,N_9512,N_9589);
and U9627 (N_9627,N_9562,N_9597);
and U9628 (N_9628,N_9612,N_9584);
nand U9629 (N_9629,N_9555,N_9518);
xnor U9630 (N_9630,N_9617,N_9621);
or U9631 (N_9631,N_9576,N_9604);
xnor U9632 (N_9632,N_9514,N_9611);
nand U9633 (N_9633,N_9606,N_9574);
xor U9634 (N_9634,N_9502,N_9546);
nor U9635 (N_9635,N_9587,N_9524);
nor U9636 (N_9636,N_9581,N_9609);
nor U9637 (N_9637,N_9526,N_9547);
nor U9638 (N_9638,N_9540,N_9575);
and U9639 (N_9639,N_9601,N_9619);
nand U9640 (N_9640,N_9552,N_9553);
nand U9641 (N_9641,N_9500,N_9595);
xor U9642 (N_9642,N_9599,N_9620);
nand U9643 (N_9643,N_9564,N_9515);
nor U9644 (N_9644,N_9531,N_9566);
and U9645 (N_9645,N_9541,N_9537);
xnor U9646 (N_9646,N_9571,N_9600);
and U9647 (N_9647,N_9527,N_9525);
nor U9648 (N_9648,N_9593,N_9623);
and U9649 (N_9649,N_9585,N_9577);
and U9650 (N_9650,N_9569,N_9602);
and U9651 (N_9651,N_9570,N_9513);
nor U9652 (N_9652,N_9603,N_9545);
xnor U9653 (N_9653,N_9554,N_9578);
xor U9654 (N_9654,N_9536,N_9523);
or U9655 (N_9655,N_9586,N_9590);
nor U9656 (N_9656,N_9544,N_9529);
xnor U9657 (N_9657,N_9610,N_9542);
nand U9658 (N_9658,N_9594,N_9522);
xor U9659 (N_9659,N_9507,N_9615);
or U9660 (N_9660,N_9539,N_9506);
nand U9661 (N_9661,N_9596,N_9549);
xnor U9662 (N_9662,N_9557,N_9561);
or U9663 (N_9663,N_9605,N_9551);
nor U9664 (N_9664,N_9572,N_9509);
xnor U9665 (N_9665,N_9505,N_9583);
nand U9666 (N_9666,N_9579,N_9501);
and U9667 (N_9667,N_9548,N_9588);
or U9668 (N_9668,N_9613,N_9533);
nor U9669 (N_9669,N_9521,N_9510);
nor U9670 (N_9670,N_9503,N_9543);
nor U9671 (N_9671,N_9624,N_9622);
nand U9672 (N_9672,N_9573,N_9558);
and U9673 (N_9673,N_9608,N_9568);
or U9674 (N_9674,N_9538,N_9528);
nand U9675 (N_9675,N_9618,N_9560);
nand U9676 (N_9676,N_9532,N_9607);
nand U9677 (N_9677,N_9519,N_9565);
nor U9678 (N_9678,N_9511,N_9508);
or U9679 (N_9679,N_9530,N_9559);
nor U9680 (N_9680,N_9534,N_9516);
nand U9681 (N_9681,N_9614,N_9535);
and U9682 (N_9682,N_9598,N_9616);
nor U9683 (N_9683,N_9563,N_9592);
and U9684 (N_9684,N_9556,N_9520);
and U9685 (N_9685,N_9504,N_9550);
or U9686 (N_9686,N_9567,N_9517);
or U9687 (N_9687,N_9591,N_9501);
xnor U9688 (N_9688,N_9581,N_9570);
nand U9689 (N_9689,N_9509,N_9579);
and U9690 (N_9690,N_9619,N_9604);
nand U9691 (N_9691,N_9527,N_9500);
or U9692 (N_9692,N_9585,N_9606);
nor U9693 (N_9693,N_9596,N_9610);
and U9694 (N_9694,N_9562,N_9611);
nand U9695 (N_9695,N_9533,N_9599);
nand U9696 (N_9696,N_9587,N_9535);
xnor U9697 (N_9697,N_9610,N_9619);
nand U9698 (N_9698,N_9579,N_9604);
xor U9699 (N_9699,N_9514,N_9531);
or U9700 (N_9700,N_9567,N_9590);
or U9701 (N_9701,N_9545,N_9602);
and U9702 (N_9702,N_9623,N_9612);
or U9703 (N_9703,N_9580,N_9589);
nor U9704 (N_9704,N_9574,N_9522);
xnor U9705 (N_9705,N_9568,N_9514);
or U9706 (N_9706,N_9549,N_9577);
nor U9707 (N_9707,N_9512,N_9610);
or U9708 (N_9708,N_9549,N_9584);
or U9709 (N_9709,N_9537,N_9562);
nor U9710 (N_9710,N_9541,N_9571);
nand U9711 (N_9711,N_9560,N_9503);
and U9712 (N_9712,N_9540,N_9597);
and U9713 (N_9713,N_9586,N_9508);
nor U9714 (N_9714,N_9526,N_9620);
or U9715 (N_9715,N_9565,N_9620);
and U9716 (N_9716,N_9586,N_9534);
nand U9717 (N_9717,N_9538,N_9616);
xor U9718 (N_9718,N_9589,N_9615);
nand U9719 (N_9719,N_9511,N_9590);
nand U9720 (N_9720,N_9500,N_9594);
or U9721 (N_9721,N_9613,N_9583);
or U9722 (N_9722,N_9552,N_9610);
or U9723 (N_9723,N_9544,N_9615);
and U9724 (N_9724,N_9508,N_9577);
nand U9725 (N_9725,N_9609,N_9535);
or U9726 (N_9726,N_9528,N_9529);
xor U9727 (N_9727,N_9581,N_9565);
xor U9728 (N_9728,N_9507,N_9596);
xnor U9729 (N_9729,N_9541,N_9544);
nor U9730 (N_9730,N_9586,N_9546);
and U9731 (N_9731,N_9549,N_9611);
nand U9732 (N_9732,N_9535,N_9578);
nor U9733 (N_9733,N_9550,N_9549);
or U9734 (N_9734,N_9609,N_9580);
or U9735 (N_9735,N_9525,N_9516);
nor U9736 (N_9736,N_9611,N_9583);
and U9737 (N_9737,N_9613,N_9597);
and U9738 (N_9738,N_9508,N_9548);
nor U9739 (N_9739,N_9566,N_9582);
xor U9740 (N_9740,N_9552,N_9519);
nor U9741 (N_9741,N_9557,N_9500);
xor U9742 (N_9742,N_9577,N_9551);
xnor U9743 (N_9743,N_9592,N_9500);
or U9744 (N_9744,N_9624,N_9570);
nand U9745 (N_9745,N_9527,N_9535);
or U9746 (N_9746,N_9621,N_9540);
nor U9747 (N_9747,N_9581,N_9608);
nand U9748 (N_9748,N_9558,N_9574);
xnor U9749 (N_9749,N_9559,N_9510);
nand U9750 (N_9750,N_9730,N_9715);
and U9751 (N_9751,N_9634,N_9649);
nor U9752 (N_9752,N_9698,N_9723);
nand U9753 (N_9753,N_9693,N_9647);
nor U9754 (N_9754,N_9727,N_9652);
xnor U9755 (N_9755,N_9678,N_9714);
nor U9756 (N_9756,N_9718,N_9685);
and U9757 (N_9757,N_9712,N_9692);
nand U9758 (N_9758,N_9661,N_9696);
nor U9759 (N_9759,N_9677,N_9695);
and U9760 (N_9760,N_9710,N_9707);
xor U9761 (N_9761,N_9667,N_9673);
nor U9762 (N_9762,N_9689,N_9665);
nor U9763 (N_9763,N_9739,N_9740);
nor U9764 (N_9764,N_9668,N_9719);
and U9765 (N_9765,N_9644,N_9669);
nand U9766 (N_9766,N_9721,N_9641);
nand U9767 (N_9767,N_9684,N_9681);
and U9768 (N_9768,N_9738,N_9703);
nor U9769 (N_9769,N_9706,N_9650);
nand U9770 (N_9770,N_9713,N_9709);
and U9771 (N_9771,N_9691,N_9645);
nand U9772 (N_9772,N_9734,N_9690);
and U9773 (N_9773,N_9662,N_9749);
nor U9774 (N_9774,N_9686,N_9670);
xnor U9775 (N_9775,N_9720,N_9631);
or U9776 (N_9776,N_9642,N_9716);
and U9777 (N_9777,N_9651,N_9737);
nand U9778 (N_9778,N_9679,N_9656);
xnor U9779 (N_9779,N_9672,N_9748);
nand U9780 (N_9780,N_9711,N_9674);
xnor U9781 (N_9781,N_9663,N_9683);
xnor U9782 (N_9782,N_9700,N_9638);
and U9783 (N_9783,N_9648,N_9688);
xnor U9784 (N_9784,N_9701,N_9635);
xnor U9785 (N_9785,N_9653,N_9728);
xor U9786 (N_9786,N_9705,N_9732);
xor U9787 (N_9787,N_9666,N_9743);
xnor U9788 (N_9788,N_9708,N_9659);
xnor U9789 (N_9789,N_9722,N_9725);
or U9790 (N_9790,N_9736,N_9675);
xor U9791 (N_9791,N_9747,N_9630);
nor U9792 (N_9792,N_9660,N_9625);
or U9793 (N_9793,N_9629,N_9729);
nand U9794 (N_9794,N_9633,N_9682);
nor U9795 (N_9795,N_9627,N_9628);
and U9796 (N_9796,N_9741,N_9676);
or U9797 (N_9797,N_9640,N_9654);
or U9798 (N_9798,N_9704,N_9702);
xnor U9799 (N_9799,N_9637,N_9742);
nor U9800 (N_9800,N_9639,N_9632);
and U9801 (N_9801,N_9636,N_9735);
nor U9802 (N_9802,N_9643,N_9694);
nor U9803 (N_9803,N_9658,N_9697);
nor U9804 (N_9804,N_9731,N_9646);
or U9805 (N_9805,N_9626,N_9664);
and U9806 (N_9806,N_9745,N_9717);
nand U9807 (N_9807,N_9726,N_9699);
and U9808 (N_9808,N_9680,N_9687);
xnor U9809 (N_9809,N_9671,N_9744);
and U9810 (N_9810,N_9657,N_9746);
nor U9811 (N_9811,N_9655,N_9724);
nor U9812 (N_9812,N_9733,N_9707);
and U9813 (N_9813,N_9732,N_9713);
and U9814 (N_9814,N_9728,N_9727);
and U9815 (N_9815,N_9673,N_9655);
or U9816 (N_9816,N_9715,N_9731);
xnor U9817 (N_9817,N_9745,N_9679);
nand U9818 (N_9818,N_9667,N_9749);
xnor U9819 (N_9819,N_9721,N_9712);
nor U9820 (N_9820,N_9680,N_9739);
xor U9821 (N_9821,N_9713,N_9677);
or U9822 (N_9822,N_9729,N_9631);
nand U9823 (N_9823,N_9723,N_9690);
xor U9824 (N_9824,N_9677,N_9745);
nand U9825 (N_9825,N_9712,N_9644);
nor U9826 (N_9826,N_9636,N_9701);
and U9827 (N_9827,N_9716,N_9732);
nor U9828 (N_9828,N_9660,N_9748);
and U9829 (N_9829,N_9664,N_9691);
and U9830 (N_9830,N_9703,N_9682);
and U9831 (N_9831,N_9725,N_9710);
and U9832 (N_9832,N_9701,N_9675);
xor U9833 (N_9833,N_9693,N_9643);
or U9834 (N_9834,N_9650,N_9690);
or U9835 (N_9835,N_9674,N_9726);
or U9836 (N_9836,N_9654,N_9659);
or U9837 (N_9837,N_9743,N_9731);
and U9838 (N_9838,N_9724,N_9640);
or U9839 (N_9839,N_9668,N_9746);
xnor U9840 (N_9840,N_9689,N_9637);
or U9841 (N_9841,N_9709,N_9693);
and U9842 (N_9842,N_9640,N_9677);
or U9843 (N_9843,N_9654,N_9696);
nand U9844 (N_9844,N_9681,N_9728);
nor U9845 (N_9845,N_9643,N_9704);
or U9846 (N_9846,N_9678,N_9749);
xnor U9847 (N_9847,N_9667,N_9631);
or U9848 (N_9848,N_9701,N_9710);
xor U9849 (N_9849,N_9719,N_9628);
xnor U9850 (N_9850,N_9674,N_9690);
and U9851 (N_9851,N_9696,N_9708);
nand U9852 (N_9852,N_9699,N_9674);
or U9853 (N_9853,N_9651,N_9725);
xnor U9854 (N_9854,N_9630,N_9671);
nor U9855 (N_9855,N_9661,N_9748);
xnor U9856 (N_9856,N_9627,N_9632);
and U9857 (N_9857,N_9709,N_9742);
nand U9858 (N_9858,N_9642,N_9674);
xnor U9859 (N_9859,N_9732,N_9671);
nand U9860 (N_9860,N_9706,N_9664);
and U9861 (N_9861,N_9644,N_9733);
and U9862 (N_9862,N_9723,N_9687);
or U9863 (N_9863,N_9690,N_9688);
and U9864 (N_9864,N_9649,N_9726);
xor U9865 (N_9865,N_9683,N_9674);
nor U9866 (N_9866,N_9676,N_9685);
and U9867 (N_9867,N_9684,N_9706);
nand U9868 (N_9868,N_9662,N_9660);
and U9869 (N_9869,N_9670,N_9743);
xnor U9870 (N_9870,N_9630,N_9628);
nor U9871 (N_9871,N_9716,N_9703);
nor U9872 (N_9872,N_9637,N_9731);
nand U9873 (N_9873,N_9647,N_9654);
nor U9874 (N_9874,N_9651,N_9663);
nand U9875 (N_9875,N_9771,N_9750);
nand U9876 (N_9876,N_9842,N_9818);
and U9877 (N_9877,N_9787,N_9819);
nand U9878 (N_9878,N_9753,N_9846);
nor U9879 (N_9879,N_9853,N_9817);
or U9880 (N_9880,N_9761,N_9812);
xor U9881 (N_9881,N_9830,N_9825);
or U9882 (N_9882,N_9781,N_9852);
nand U9883 (N_9883,N_9808,N_9834);
nor U9884 (N_9884,N_9826,N_9799);
nand U9885 (N_9885,N_9780,N_9833);
or U9886 (N_9886,N_9828,N_9861);
nor U9887 (N_9887,N_9868,N_9863);
or U9888 (N_9888,N_9837,N_9768);
and U9889 (N_9889,N_9785,N_9758);
and U9890 (N_9890,N_9769,N_9792);
xnor U9891 (N_9891,N_9858,N_9800);
nand U9892 (N_9892,N_9831,N_9789);
nor U9893 (N_9893,N_9822,N_9848);
nor U9894 (N_9894,N_9856,N_9773);
xnor U9895 (N_9895,N_9855,N_9803);
xor U9896 (N_9896,N_9766,N_9849);
nor U9897 (N_9897,N_9804,N_9757);
and U9898 (N_9898,N_9836,N_9824);
nor U9899 (N_9899,N_9864,N_9838);
and U9900 (N_9900,N_9791,N_9859);
xnor U9901 (N_9901,N_9778,N_9866);
nor U9902 (N_9902,N_9847,N_9851);
xnor U9903 (N_9903,N_9786,N_9827);
nor U9904 (N_9904,N_9839,N_9867);
or U9905 (N_9905,N_9870,N_9807);
xnor U9906 (N_9906,N_9810,N_9821);
or U9907 (N_9907,N_9860,N_9790);
xor U9908 (N_9908,N_9871,N_9772);
nor U9909 (N_9909,N_9843,N_9850);
and U9910 (N_9910,N_9811,N_9865);
or U9911 (N_9911,N_9806,N_9823);
nand U9912 (N_9912,N_9755,N_9832);
or U9913 (N_9913,N_9857,N_9844);
or U9914 (N_9914,N_9793,N_9775);
nand U9915 (N_9915,N_9759,N_9776);
nand U9916 (N_9916,N_9777,N_9797);
or U9917 (N_9917,N_9816,N_9774);
and U9918 (N_9918,N_9873,N_9801);
or U9919 (N_9919,N_9835,N_9763);
and U9920 (N_9920,N_9796,N_9829);
nor U9921 (N_9921,N_9854,N_9862);
and U9922 (N_9922,N_9760,N_9820);
and U9923 (N_9923,N_9752,N_9872);
xor U9924 (N_9924,N_9813,N_9762);
xor U9925 (N_9925,N_9765,N_9874);
xnor U9926 (N_9926,N_9840,N_9798);
nor U9927 (N_9927,N_9783,N_9756);
and U9928 (N_9928,N_9869,N_9782);
or U9929 (N_9929,N_9751,N_9841);
xnor U9930 (N_9930,N_9814,N_9845);
nor U9931 (N_9931,N_9795,N_9764);
xor U9932 (N_9932,N_9794,N_9784);
xor U9933 (N_9933,N_9802,N_9767);
xor U9934 (N_9934,N_9770,N_9815);
nand U9935 (N_9935,N_9809,N_9779);
nor U9936 (N_9936,N_9788,N_9754);
nor U9937 (N_9937,N_9805,N_9790);
xor U9938 (N_9938,N_9810,N_9763);
xor U9939 (N_9939,N_9752,N_9871);
and U9940 (N_9940,N_9852,N_9858);
nand U9941 (N_9941,N_9849,N_9831);
and U9942 (N_9942,N_9798,N_9818);
and U9943 (N_9943,N_9849,N_9752);
or U9944 (N_9944,N_9771,N_9752);
and U9945 (N_9945,N_9853,N_9847);
or U9946 (N_9946,N_9802,N_9824);
xnor U9947 (N_9947,N_9784,N_9778);
and U9948 (N_9948,N_9792,N_9763);
xnor U9949 (N_9949,N_9784,N_9753);
nor U9950 (N_9950,N_9830,N_9815);
and U9951 (N_9951,N_9796,N_9751);
nand U9952 (N_9952,N_9760,N_9752);
and U9953 (N_9953,N_9853,N_9789);
xor U9954 (N_9954,N_9848,N_9868);
nand U9955 (N_9955,N_9834,N_9858);
xor U9956 (N_9956,N_9843,N_9807);
nand U9957 (N_9957,N_9795,N_9770);
nor U9958 (N_9958,N_9867,N_9816);
nand U9959 (N_9959,N_9759,N_9842);
xnor U9960 (N_9960,N_9760,N_9810);
nand U9961 (N_9961,N_9816,N_9869);
nor U9962 (N_9962,N_9870,N_9816);
nor U9963 (N_9963,N_9866,N_9804);
xnor U9964 (N_9964,N_9815,N_9800);
or U9965 (N_9965,N_9812,N_9776);
nand U9966 (N_9966,N_9762,N_9869);
nand U9967 (N_9967,N_9803,N_9811);
and U9968 (N_9968,N_9790,N_9782);
nand U9969 (N_9969,N_9758,N_9797);
and U9970 (N_9970,N_9774,N_9786);
or U9971 (N_9971,N_9784,N_9820);
or U9972 (N_9972,N_9873,N_9789);
or U9973 (N_9973,N_9827,N_9823);
xor U9974 (N_9974,N_9844,N_9788);
or U9975 (N_9975,N_9799,N_9767);
or U9976 (N_9976,N_9756,N_9861);
nor U9977 (N_9977,N_9775,N_9785);
or U9978 (N_9978,N_9762,N_9817);
and U9979 (N_9979,N_9752,N_9862);
or U9980 (N_9980,N_9794,N_9824);
nand U9981 (N_9981,N_9871,N_9783);
xnor U9982 (N_9982,N_9874,N_9802);
nand U9983 (N_9983,N_9827,N_9841);
or U9984 (N_9984,N_9804,N_9850);
xor U9985 (N_9985,N_9794,N_9799);
nor U9986 (N_9986,N_9809,N_9761);
or U9987 (N_9987,N_9762,N_9780);
and U9988 (N_9988,N_9846,N_9798);
nor U9989 (N_9989,N_9793,N_9825);
nor U9990 (N_9990,N_9820,N_9764);
nor U9991 (N_9991,N_9813,N_9782);
xnor U9992 (N_9992,N_9809,N_9776);
xnor U9993 (N_9993,N_9872,N_9831);
nor U9994 (N_9994,N_9778,N_9788);
or U9995 (N_9995,N_9858,N_9817);
xor U9996 (N_9996,N_9762,N_9765);
and U9997 (N_9997,N_9857,N_9792);
or U9998 (N_9998,N_9833,N_9872);
nor U9999 (N_9999,N_9811,N_9828);
or U10000 (N_10000,N_9999,N_9954);
and U10001 (N_10001,N_9948,N_9926);
and U10002 (N_10002,N_9924,N_9947);
and U10003 (N_10003,N_9884,N_9987);
nor U10004 (N_10004,N_9919,N_9977);
and U10005 (N_10005,N_9962,N_9934);
or U10006 (N_10006,N_9878,N_9998);
nor U10007 (N_10007,N_9985,N_9951);
nor U10008 (N_10008,N_9901,N_9913);
or U10009 (N_10009,N_9993,N_9983);
xnor U10010 (N_10010,N_9904,N_9970);
nor U10011 (N_10011,N_9880,N_9905);
nand U10012 (N_10012,N_9902,N_9988);
or U10013 (N_10013,N_9911,N_9927);
xnor U10014 (N_10014,N_9912,N_9898);
nand U10015 (N_10015,N_9994,N_9939);
xor U10016 (N_10016,N_9995,N_9923);
or U10017 (N_10017,N_9889,N_9937);
nand U10018 (N_10018,N_9917,N_9925);
and U10019 (N_10019,N_9950,N_9943);
or U10020 (N_10020,N_9891,N_9965);
nor U10021 (N_10021,N_9933,N_9940);
nand U10022 (N_10022,N_9936,N_9959);
and U10023 (N_10023,N_9938,N_9928);
xnor U10024 (N_10024,N_9899,N_9941);
nor U10025 (N_10025,N_9979,N_9966);
or U10026 (N_10026,N_9978,N_9946);
nor U10027 (N_10027,N_9918,N_9976);
nand U10028 (N_10028,N_9982,N_9960);
and U10029 (N_10029,N_9921,N_9920);
nor U10030 (N_10030,N_9932,N_9929);
or U10031 (N_10031,N_9885,N_9984);
nand U10032 (N_10032,N_9916,N_9955);
nand U10033 (N_10033,N_9930,N_9968);
nand U10034 (N_10034,N_9877,N_9907);
xnor U10035 (N_10035,N_9882,N_9949);
nor U10036 (N_10036,N_9956,N_9879);
nand U10037 (N_10037,N_9893,N_9886);
xnor U10038 (N_10038,N_9974,N_9989);
nand U10039 (N_10039,N_9888,N_9892);
and U10040 (N_10040,N_9961,N_9895);
xor U10041 (N_10041,N_9997,N_9945);
and U10042 (N_10042,N_9981,N_9883);
xor U10043 (N_10043,N_9908,N_9910);
or U10044 (N_10044,N_9991,N_9942);
or U10045 (N_10045,N_9971,N_9935);
nor U10046 (N_10046,N_9914,N_9958);
nand U10047 (N_10047,N_9876,N_9897);
or U10048 (N_10048,N_9922,N_9969);
or U10049 (N_10049,N_9957,N_9964);
xor U10050 (N_10050,N_9986,N_9881);
and U10051 (N_10051,N_9931,N_9992);
nor U10052 (N_10052,N_9973,N_9953);
or U10053 (N_10053,N_9963,N_9896);
or U10054 (N_10054,N_9990,N_9980);
nor U10055 (N_10055,N_9887,N_9975);
and U10056 (N_10056,N_9909,N_9972);
nand U10057 (N_10057,N_9875,N_9890);
or U10058 (N_10058,N_9903,N_9996);
or U10059 (N_10059,N_9906,N_9894);
or U10060 (N_10060,N_9952,N_9915);
nand U10061 (N_10061,N_9900,N_9944);
and U10062 (N_10062,N_9967,N_9974);
nand U10063 (N_10063,N_9973,N_9960);
nor U10064 (N_10064,N_9994,N_9936);
xnor U10065 (N_10065,N_9993,N_9879);
nand U10066 (N_10066,N_9881,N_9943);
xor U10067 (N_10067,N_9892,N_9964);
xnor U10068 (N_10068,N_9968,N_9891);
nand U10069 (N_10069,N_9968,N_9995);
nor U10070 (N_10070,N_9987,N_9890);
or U10071 (N_10071,N_9935,N_9980);
nand U10072 (N_10072,N_9883,N_9936);
and U10073 (N_10073,N_9901,N_9934);
nor U10074 (N_10074,N_9976,N_9911);
xnor U10075 (N_10075,N_9902,N_9916);
xor U10076 (N_10076,N_9940,N_9883);
nor U10077 (N_10077,N_9904,N_9952);
xor U10078 (N_10078,N_9969,N_9980);
xnor U10079 (N_10079,N_9995,N_9954);
or U10080 (N_10080,N_9929,N_9996);
nand U10081 (N_10081,N_9931,N_9912);
nor U10082 (N_10082,N_9952,N_9997);
and U10083 (N_10083,N_9892,N_9940);
or U10084 (N_10084,N_9919,N_9982);
or U10085 (N_10085,N_9900,N_9974);
xor U10086 (N_10086,N_9900,N_9981);
and U10087 (N_10087,N_9894,N_9914);
nor U10088 (N_10088,N_9991,N_9884);
nand U10089 (N_10089,N_9915,N_9983);
xor U10090 (N_10090,N_9885,N_9875);
and U10091 (N_10091,N_9975,N_9926);
xnor U10092 (N_10092,N_9884,N_9909);
nor U10093 (N_10093,N_9928,N_9968);
and U10094 (N_10094,N_9948,N_9922);
xnor U10095 (N_10095,N_9913,N_9959);
nand U10096 (N_10096,N_9909,N_9885);
and U10097 (N_10097,N_9999,N_9906);
nor U10098 (N_10098,N_9894,N_9893);
or U10099 (N_10099,N_9886,N_9909);
nor U10100 (N_10100,N_9890,N_9881);
and U10101 (N_10101,N_9924,N_9983);
and U10102 (N_10102,N_9917,N_9985);
nor U10103 (N_10103,N_9880,N_9930);
nor U10104 (N_10104,N_9878,N_9929);
and U10105 (N_10105,N_9935,N_9968);
and U10106 (N_10106,N_9976,N_9999);
and U10107 (N_10107,N_9966,N_9957);
and U10108 (N_10108,N_9966,N_9911);
xor U10109 (N_10109,N_9930,N_9876);
and U10110 (N_10110,N_9987,N_9965);
and U10111 (N_10111,N_9932,N_9944);
xor U10112 (N_10112,N_9896,N_9921);
or U10113 (N_10113,N_9969,N_9932);
xnor U10114 (N_10114,N_9988,N_9963);
nor U10115 (N_10115,N_9906,N_9994);
xnor U10116 (N_10116,N_9996,N_9973);
nor U10117 (N_10117,N_9942,N_9982);
and U10118 (N_10118,N_9932,N_9889);
and U10119 (N_10119,N_9944,N_9963);
xnor U10120 (N_10120,N_9957,N_9970);
xor U10121 (N_10121,N_9878,N_9942);
and U10122 (N_10122,N_9944,N_9914);
nand U10123 (N_10123,N_9887,N_9922);
nor U10124 (N_10124,N_9977,N_9950);
and U10125 (N_10125,N_10022,N_10015);
nand U10126 (N_10126,N_10094,N_10061);
nor U10127 (N_10127,N_10120,N_10004);
and U10128 (N_10128,N_10019,N_10081);
xor U10129 (N_10129,N_10107,N_10075);
nor U10130 (N_10130,N_10012,N_10085);
and U10131 (N_10131,N_10102,N_10123);
nor U10132 (N_10132,N_10080,N_10083);
and U10133 (N_10133,N_10059,N_10103);
and U10134 (N_10134,N_10096,N_10065);
xnor U10135 (N_10135,N_10113,N_10068);
and U10136 (N_10136,N_10024,N_10079);
nor U10137 (N_10137,N_10051,N_10115);
nor U10138 (N_10138,N_10055,N_10052);
or U10139 (N_10139,N_10027,N_10111);
and U10140 (N_10140,N_10099,N_10087);
or U10141 (N_10141,N_10033,N_10044);
nand U10142 (N_10142,N_10008,N_10023);
or U10143 (N_10143,N_10098,N_10063);
xor U10144 (N_10144,N_10045,N_10070);
nor U10145 (N_10145,N_10071,N_10025);
or U10146 (N_10146,N_10000,N_10108);
nor U10147 (N_10147,N_10042,N_10020);
xnor U10148 (N_10148,N_10016,N_10069);
nand U10149 (N_10149,N_10046,N_10040);
xnor U10150 (N_10150,N_10072,N_10034);
or U10151 (N_10151,N_10109,N_10005);
nor U10152 (N_10152,N_10088,N_10037);
nand U10153 (N_10153,N_10014,N_10104);
nor U10154 (N_10154,N_10076,N_10029);
or U10155 (N_10155,N_10074,N_10058);
nand U10156 (N_10156,N_10122,N_10017);
or U10157 (N_10157,N_10032,N_10053);
or U10158 (N_10158,N_10117,N_10090);
nand U10159 (N_10159,N_10048,N_10036);
and U10160 (N_10160,N_10060,N_10092);
or U10161 (N_10161,N_10124,N_10062);
nand U10162 (N_10162,N_10119,N_10110);
nand U10163 (N_10163,N_10031,N_10077);
and U10164 (N_10164,N_10009,N_10095);
or U10165 (N_10165,N_10097,N_10038);
and U10166 (N_10166,N_10112,N_10047);
nor U10167 (N_10167,N_10116,N_10101);
nor U10168 (N_10168,N_10013,N_10067);
xnor U10169 (N_10169,N_10026,N_10043);
xor U10170 (N_10170,N_10039,N_10003);
nand U10171 (N_10171,N_10078,N_10011);
nor U10172 (N_10172,N_10073,N_10118);
nor U10173 (N_10173,N_10018,N_10028);
xor U10174 (N_10174,N_10054,N_10089);
nand U10175 (N_10175,N_10050,N_10086);
nand U10176 (N_10176,N_10106,N_10021);
nand U10177 (N_10177,N_10093,N_10057);
or U10178 (N_10178,N_10100,N_10056);
and U10179 (N_10179,N_10002,N_10084);
xnor U10180 (N_10180,N_10066,N_10049);
nand U10181 (N_10181,N_10091,N_10041);
xor U10182 (N_10182,N_10001,N_10030);
and U10183 (N_10183,N_10121,N_10082);
and U10184 (N_10184,N_10064,N_10007);
nand U10185 (N_10185,N_10114,N_10105);
nand U10186 (N_10186,N_10006,N_10010);
xor U10187 (N_10187,N_10035,N_10069);
nand U10188 (N_10188,N_10003,N_10000);
nor U10189 (N_10189,N_10057,N_10013);
nand U10190 (N_10190,N_10038,N_10037);
or U10191 (N_10191,N_10033,N_10005);
and U10192 (N_10192,N_10063,N_10000);
nor U10193 (N_10193,N_10117,N_10084);
and U10194 (N_10194,N_10020,N_10006);
and U10195 (N_10195,N_10048,N_10117);
nand U10196 (N_10196,N_10011,N_10087);
and U10197 (N_10197,N_10104,N_10061);
nor U10198 (N_10198,N_10091,N_10029);
and U10199 (N_10199,N_10115,N_10109);
xnor U10200 (N_10200,N_10009,N_10017);
nor U10201 (N_10201,N_10090,N_10122);
and U10202 (N_10202,N_10041,N_10086);
or U10203 (N_10203,N_10097,N_10029);
and U10204 (N_10204,N_10031,N_10061);
or U10205 (N_10205,N_10098,N_10075);
nor U10206 (N_10206,N_10057,N_10036);
or U10207 (N_10207,N_10015,N_10021);
xor U10208 (N_10208,N_10124,N_10092);
or U10209 (N_10209,N_10022,N_10010);
or U10210 (N_10210,N_10116,N_10088);
nor U10211 (N_10211,N_10121,N_10048);
nor U10212 (N_10212,N_10081,N_10034);
or U10213 (N_10213,N_10083,N_10041);
nand U10214 (N_10214,N_10049,N_10099);
nand U10215 (N_10215,N_10122,N_10119);
or U10216 (N_10216,N_10068,N_10004);
nor U10217 (N_10217,N_10070,N_10094);
nor U10218 (N_10218,N_10002,N_10109);
xor U10219 (N_10219,N_10002,N_10066);
nor U10220 (N_10220,N_10051,N_10004);
nand U10221 (N_10221,N_10002,N_10010);
nor U10222 (N_10222,N_10114,N_10120);
or U10223 (N_10223,N_10009,N_10075);
xor U10224 (N_10224,N_10102,N_10056);
or U10225 (N_10225,N_10047,N_10004);
xor U10226 (N_10226,N_10122,N_10075);
nor U10227 (N_10227,N_10062,N_10053);
nand U10228 (N_10228,N_10103,N_10104);
or U10229 (N_10229,N_10110,N_10085);
xor U10230 (N_10230,N_10042,N_10005);
xor U10231 (N_10231,N_10076,N_10116);
and U10232 (N_10232,N_10015,N_10052);
xor U10233 (N_10233,N_10093,N_10011);
nor U10234 (N_10234,N_10022,N_10042);
xnor U10235 (N_10235,N_10113,N_10081);
or U10236 (N_10236,N_10042,N_10093);
nand U10237 (N_10237,N_10099,N_10112);
and U10238 (N_10238,N_10031,N_10110);
or U10239 (N_10239,N_10005,N_10029);
nand U10240 (N_10240,N_10108,N_10099);
nor U10241 (N_10241,N_10107,N_10094);
nand U10242 (N_10242,N_10110,N_10058);
nor U10243 (N_10243,N_10100,N_10116);
nor U10244 (N_10244,N_10081,N_10036);
nand U10245 (N_10245,N_10066,N_10024);
nand U10246 (N_10246,N_10070,N_10000);
and U10247 (N_10247,N_10092,N_10067);
or U10248 (N_10248,N_10011,N_10007);
or U10249 (N_10249,N_10017,N_10049);
nand U10250 (N_10250,N_10163,N_10148);
or U10251 (N_10251,N_10194,N_10186);
nor U10252 (N_10252,N_10172,N_10175);
xor U10253 (N_10253,N_10167,N_10236);
xnor U10254 (N_10254,N_10203,N_10151);
xnor U10255 (N_10255,N_10229,N_10219);
nor U10256 (N_10256,N_10249,N_10182);
xnor U10257 (N_10257,N_10143,N_10130);
xnor U10258 (N_10258,N_10189,N_10240);
or U10259 (N_10259,N_10214,N_10232);
or U10260 (N_10260,N_10131,N_10140);
and U10261 (N_10261,N_10139,N_10216);
nor U10262 (N_10262,N_10193,N_10132);
nor U10263 (N_10263,N_10196,N_10181);
and U10264 (N_10264,N_10192,N_10244);
nor U10265 (N_10265,N_10171,N_10180);
xor U10266 (N_10266,N_10187,N_10212);
or U10267 (N_10267,N_10165,N_10125);
or U10268 (N_10268,N_10239,N_10217);
and U10269 (N_10269,N_10184,N_10224);
nor U10270 (N_10270,N_10210,N_10199);
or U10271 (N_10271,N_10170,N_10220);
nor U10272 (N_10272,N_10176,N_10227);
or U10273 (N_10273,N_10178,N_10204);
nor U10274 (N_10274,N_10134,N_10174);
or U10275 (N_10275,N_10198,N_10188);
xnor U10276 (N_10276,N_10222,N_10195);
and U10277 (N_10277,N_10213,N_10215);
nor U10278 (N_10278,N_10226,N_10233);
nand U10279 (N_10279,N_10142,N_10248);
xor U10280 (N_10280,N_10133,N_10166);
xor U10281 (N_10281,N_10230,N_10185);
xnor U10282 (N_10282,N_10206,N_10150);
xnor U10283 (N_10283,N_10238,N_10153);
or U10284 (N_10284,N_10129,N_10160);
xor U10285 (N_10285,N_10202,N_10234);
xnor U10286 (N_10286,N_10247,N_10177);
or U10287 (N_10287,N_10155,N_10162);
or U10288 (N_10288,N_10207,N_10228);
nand U10289 (N_10289,N_10159,N_10127);
xnor U10290 (N_10290,N_10225,N_10179);
or U10291 (N_10291,N_10149,N_10168);
xnor U10292 (N_10292,N_10231,N_10197);
or U10293 (N_10293,N_10164,N_10243);
nand U10294 (N_10294,N_10209,N_10144);
nand U10295 (N_10295,N_10191,N_10138);
nand U10296 (N_10296,N_10245,N_10128);
and U10297 (N_10297,N_10221,N_10135);
xor U10298 (N_10298,N_10241,N_10235);
xor U10299 (N_10299,N_10173,N_10237);
nand U10300 (N_10300,N_10183,N_10126);
nand U10301 (N_10301,N_10161,N_10147);
nor U10302 (N_10302,N_10246,N_10157);
nor U10303 (N_10303,N_10154,N_10146);
or U10304 (N_10304,N_10169,N_10156);
xnor U10305 (N_10305,N_10190,N_10211);
xnor U10306 (N_10306,N_10158,N_10136);
xnor U10307 (N_10307,N_10218,N_10201);
nor U10308 (N_10308,N_10141,N_10223);
and U10309 (N_10309,N_10145,N_10208);
or U10310 (N_10310,N_10200,N_10137);
nor U10311 (N_10311,N_10152,N_10242);
and U10312 (N_10312,N_10205,N_10141);
or U10313 (N_10313,N_10162,N_10126);
and U10314 (N_10314,N_10217,N_10171);
or U10315 (N_10315,N_10195,N_10168);
nor U10316 (N_10316,N_10219,N_10142);
or U10317 (N_10317,N_10154,N_10219);
xor U10318 (N_10318,N_10222,N_10151);
xor U10319 (N_10319,N_10202,N_10130);
and U10320 (N_10320,N_10152,N_10193);
and U10321 (N_10321,N_10224,N_10247);
or U10322 (N_10322,N_10192,N_10221);
nand U10323 (N_10323,N_10130,N_10186);
nor U10324 (N_10324,N_10248,N_10160);
or U10325 (N_10325,N_10201,N_10146);
or U10326 (N_10326,N_10182,N_10244);
and U10327 (N_10327,N_10201,N_10158);
nand U10328 (N_10328,N_10193,N_10217);
xnor U10329 (N_10329,N_10207,N_10229);
nand U10330 (N_10330,N_10229,N_10128);
nand U10331 (N_10331,N_10241,N_10129);
nand U10332 (N_10332,N_10245,N_10218);
and U10333 (N_10333,N_10247,N_10132);
or U10334 (N_10334,N_10170,N_10181);
xor U10335 (N_10335,N_10226,N_10216);
nand U10336 (N_10336,N_10228,N_10183);
and U10337 (N_10337,N_10142,N_10212);
nor U10338 (N_10338,N_10153,N_10156);
nor U10339 (N_10339,N_10228,N_10178);
or U10340 (N_10340,N_10201,N_10132);
nor U10341 (N_10341,N_10132,N_10217);
or U10342 (N_10342,N_10249,N_10211);
xnor U10343 (N_10343,N_10249,N_10146);
nand U10344 (N_10344,N_10163,N_10202);
or U10345 (N_10345,N_10172,N_10234);
or U10346 (N_10346,N_10167,N_10141);
and U10347 (N_10347,N_10198,N_10144);
or U10348 (N_10348,N_10233,N_10138);
nor U10349 (N_10349,N_10139,N_10165);
or U10350 (N_10350,N_10144,N_10147);
xnor U10351 (N_10351,N_10232,N_10220);
or U10352 (N_10352,N_10173,N_10188);
or U10353 (N_10353,N_10229,N_10162);
or U10354 (N_10354,N_10189,N_10137);
nor U10355 (N_10355,N_10184,N_10200);
and U10356 (N_10356,N_10249,N_10130);
nor U10357 (N_10357,N_10152,N_10244);
xor U10358 (N_10358,N_10140,N_10249);
xor U10359 (N_10359,N_10216,N_10201);
and U10360 (N_10360,N_10137,N_10180);
and U10361 (N_10361,N_10217,N_10138);
and U10362 (N_10362,N_10153,N_10222);
nor U10363 (N_10363,N_10239,N_10187);
xnor U10364 (N_10364,N_10225,N_10130);
and U10365 (N_10365,N_10220,N_10199);
xor U10366 (N_10366,N_10173,N_10192);
xnor U10367 (N_10367,N_10129,N_10154);
or U10368 (N_10368,N_10217,N_10205);
or U10369 (N_10369,N_10147,N_10136);
and U10370 (N_10370,N_10187,N_10154);
or U10371 (N_10371,N_10220,N_10192);
xor U10372 (N_10372,N_10195,N_10227);
nor U10373 (N_10373,N_10237,N_10160);
nand U10374 (N_10374,N_10127,N_10204);
nand U10375 (N_10375,N_10303,N_10358);
or U10376 (N_10376,N_10300,N_10267);
xor U10377 (N_10377,N_10352,N_10338);
xor U10378 (N_10378,N_10366,N_10281);
xor U10379 (N_10379,N_10269,N_10283);
nand U10380 (N_10380,N_10297,N_10355);
xnor U10381 (N_10381,N_10345,N_10365);
nor U10382 (N_10382,N_10275,N_10284);
or U10383 (N_10383,N_10346,N_10337);
and U10384 (N_10384,N_10354,N_10367);
or U10385 (N_10385,N_10279,N_10371);
and U10386 (N_10386,N_10285,N_10288);
xnor U10387 (N_10387,N_10335,N_10286);
xor U10388 (N_10388,N_10259,N_10298);
nand U10389 (N_10389,N_10321,N_10328);
xor U10390 (N_10390,N_10276,N_10262);
nand U10391 (N_10391,N_10252,N_10363);
nor U10392 (N_10392,N_10315,N_10356);
or U10393 (N_10393,N_10336,N_10339);
nand U10394 (N_10394,N_10319,N_10290);
xnor U10395 (N_10395,N_10314,N_10268);
or U10396 (N_10396,N_10316,N_10250);
and U10397 (N_10397,N_10313,N_10312);
and U10398 (N_10398,N_10282,N_10353);
nand U10399 (N_10399,N_10263,N_10272);
xnor U10400 (N_10400,N_10260,N_10359);
or U10401 (N_10401,N_10324,N_10370);
nor U10402 (N_10402,N_10331,N_10333);
nand U10403 (N_10403,N_10301,N_10280);
or U10404 (N_10404,N_10294,N_10317);
xor U10405 (N_10405,N_10349,N_10350);
nor U10406 (N_10406,N_10320,N_10369);
xor U10407 (N_10407,N_10264,N_10256);
nor U10408 (N_10408,N_10287,N_10296);
nor U10409 (N_10409,N_10347,N_10332);
xor U10410 (N_10410,N_10357,N_10330);
or U10411 (N_10411,N_10325,N_10255);
or U10412 (N_10412,N_10341,N_10311);
and U10413 (N_10413,N_10273,N_10342);
nand U10414 (N_10414,N_10310,N_10306);
or U10415 (N_10415,N_10253,N_10254);
or U10416 (N_10416,N_10304,N_10278);
xnor U10417 (N_10417,N_10322,N_10309);
and U10418 (N_10418,N_10270,N_10343);
nor U10419 (N_10419,N_10308,N_10372);
and U10420 (N_10420,N_10302,N_10305);
and U10421 (N_10421,N_10271,N_10295);
or U10422 (N_10422,N_10307,N_10289);
xor U10423 (N_10423,N_10251,N_10327);
nand U10424 (N_10424,N_10265,N_10361);
xnor U10425 (N_10425,N_10368,N_10257);
or U10426 (N_10426,N_10261,N_10258);
xnor U10427 (N_10427,N_10291,N_10299);
nand U10428 (N_10428,N_10334,N_10326);
xnor U10429 (N_10429,N_10293,N_10374);
nand U10430 (N_10430,N_10373,N_10266);
nor U10431 (N_10431,N_10292,N_10329);
nor U10432 (N_10432,N_10340,N_10362);
xor U10433 (N_10433,N_10323,N_10364);
xnor U10434 (N_10434,N_10351,N_10274);
xnor U10435 (N_10435,N_10360,N_10318);
or U10436 (N_10436,N_10348,N_10344);
nand U10437 (N_10437,N_10277,N_10268);
or U10438 (N_10438,N_10367,N_10277);
nand U10439 (N_10439,N_10291,N_10328);
and U10440 (N_10440,N_10310,N_10305);
nor U10441 (N_10441,N_10342,N_10255);
nor U10442 (N_10442,N_10304,N_10254);
and U10443 (N_10443,N_10297,N_10274);
nand U10444 (N_10444,N_10372,N_10361);
xnor U10445 (N_10445,N_10339,N_10313);
nand U10446 (N_10446,N_10369,N_10316);
nor U10447 (N_10447,N_10289,N_10342);
or U10448 (N_10448,N_10253,N_10315);
nand U10449 (N_10449,N_10281,N_10373);
or U10450 (N_10450,N_10276,N_10326);
xnor U10451 (N_10451,N_10311,N_10366);
xnor U10452 (N_10452,N_10367,N_10265);
nor U10453 (N_10453,N_10262,N_10345);
or U10454 (N_10454,N_10317,N_10337);
or U10455 (N_10455,N_10321,N_10326);
and U10456 (N_10456,N_10309,N_10297);
or U10457 (N_10457,N_10251,N_10322);
nand U10458 (N_10458,N_10313,N_10269);
nand U10459 (N_10459,N_10340,N_10365);
or U10460 (N_10460,N_10353,N_10311);
nand U10461 (N_10461,N_10272,N_10313);
xor U10462 (N_10462,N_10368,N_10293);
and U10463 (N_10463,N_10270,N_10302);
xnor U10464 (N_10464,N_10367,N_10318);
or U10465 (N_10465,N_10264,N_10317);
nor U10466 (N_10466,N_10353,N_10342);
nand U10467 (N_10467,N_10339,N_10332);
nor U10468 (N_10468,N_10354,N_10333);
xor U10469 (N_10469,N_10286,N_10352);
xnor U10470 (N_10470,N_10284,N_10267);
nor U10471 (N_10471,N_10351,N_10296);
and U10472 (N_10472,N_10305,N_10275);
and U10473 (N_10473,N_10318,N_10353);
nor U10474 (N_10474,N_10350,N_10359);
and U10475 (N_10475,N_10289,N_10330);
nand U10476 (N_10476,N_10350,N_10355);
nand U10477 (N_10477,N_10363,N_10341);
nor U10478 (N_10478,N_10268,N_10261);
and U10479 (N_10479,N_10307,N_10326);
and U10480 (N_10480,N_10256,N_10260);
nand U10481 (N_10481,N_10330,N_10331);
nor U10482 (N_10482,N_10367,N_10349);
and U10483 (N_10483,N_10303,N_10373);
nor U10484 (N_10484,N_10356,N_10308);
or U10485 (N_10485,N_10324,N_10313);
nand U10486 (N_10486,N_10374,N_10288);
xnor U10487 (N_10487,N_10276,N_10322);
and U10488 (N_10488,N_10334,N_10258);
or U10489 (N_10489,N_10359,N_10313);
nor U10490 (N_10490,N_10366,N_10347);
nor U10491 (N_10491,N_10323,N_10269);
nand U10492 (N_10492,N_10313,N_10347);
or U10493 (N_10493,N_10350,N_10332);
xnor U10494 (N_10494,N_10365,N_10317);
nor U10495 (N_10495,N_10321,N_10317);
xor U10496 (N_10496,N_10372,N_10340);
nor U10497 (N_10497,N_10360,N_10368);
nor U10498 (N_10498,N_10268,N_10336);
or U10499 (N_10499,N_10252,N_10356);
or U10500 (N_10500,N_10405,N_10391);
or U10501 (N_10501,N_10477,N_10411);
nor U10502 (N_10502,N_10453,N_10381);
or U10503 (N_10503,N_10422,N_10390);
or U10504 (N_10504,N_10485,N_10430);
or U10505 (N_10505,N_10406,N_10408);
nor U10506 (N_10506,N_10488,N_10475);
xor U10507 (N_10507,N_10494,N_10483);
nor U10508 (N_10508,N_10443,N_10441);
or U10509 (N_10509,N_10393,N_10435);
and U10510 (N_10510,N_10461,N_10471);
or U10511 (N_10511,N_10487,N_10442);
nor U10512 (N_10512,N_10382,N_10478);
or U10513 (N_10513,N_10432,N_10458);
and U10514 (N_10514,N_10482,N_10493);
nand U10515 (N_10515,N_10379,N_10473);
and U10516 (N_10516,N_10459,N_10476);
or U10517 (N_10517,N_10395,N_10462);
and U10518 (N_10518,N_10469,N_10383);
and U10519 (N_10519,N_10437,N_10492);
xnor U10520 (N_10520,N_10456,N_10385);
or U10521 (N_10521,N_10479,N_10447);
and U10522 (N_10522,N_10467,N_10399);
or U10523 (N_10523,N_10397,N_10491);
or U10524 (N_10524,N_10424,N_10413);
nor U10525 (N_10525,N_10433,N_10389);
or U10526 (N_10526,N_10486,N_10468);
nor U10527 (N_10527,N_10420,N_10410);
and U10528 (N_10528,N_10449,N_10412);
or U10529 (N_10529,N_10415,N_10429);
nor U10530 (N_10530,N_10484,N_10466);
nand U10531 (N_10531,N_10444,N_10431);
nor U10532 (N_10532,N_10452,N_10384);
nand U10533 (N_10533,N_10434,N_10451);
nor U10534 (N_10534,N_10448,N_10398);
nor U10535 (N_10535,N_10463,N_10465);
nor U10536 (N_10536,N_10427,N_10438);
xnor U10537 (N_10537,N_10470,N_10409);
nor U10538 (N_10538,N_10455,N_10436);
nand U10539 (N_10539,N_10380,N_10394);
and U10540 (N_10540,N_10499,N_10472);
nor U10541 (N_10541,N_10376,N_10489);
nand U10542 (N_10542,N_10401,N_10497);
nor U10543 (N_10543,N_10414,N_10419);
nand U10544 (N_10544,N_10387,N_10450);
nor U10545 (N_10545,N_10392,N_10423);
nor U10546 (N_10546,N_10403,N_10425);
xor U10547 (N_10547,N_10426,N_10498);
xor U10548 (N_10548,N_10439,N_10490);
and U10549 (N_10549,N_10480,N_10386);
and U10550 (N_10550,N_10375,N_10457);
nand U10551 (N_10551,N_10445,N_10496);
nor U10552 (N_10552,N_10421,N_10396);
and U10553 (N_10553,N_10417,N_10474);
nor U10554 (N_10554,N_10418,N_10440);
xnor U10555 (N_10555,N_10416,N_10481);
xor U10556 (N_10556,N_10454,N_10402);
or U10557 (N_10557,N_10377,N_10428);
or U10558 (N_10558,N_10407,N_10388);
or U10559 (N_10559,N_10404,N_10378);
and U10560 (N_10560,N_10464,N_10400);
nor U10561 (N_10561,N_10495,N_10460);
or U10562 (N_10562,N_10446,N_10409);
nor U10563 (N_10563,N_10487,N_10397);
nor U10564 (N_10564,N_10431,N_10426);
xor U10565 (N_10565,N_10432,N_10411);
and U10566 (N_10566,N_10433,N_10415);
or U10567 (N_10567,N_10439,N_10468);
nand U10568 (N_10568,N_10408,N_10436);
and U10569 (N_10569,N_10433,N_10453);
nand U10570 (N_10570,N_10487,N_10432);
or U10571 (N_10571,N_10425,N_10490);
nor U10572 (N_10572,N_10462,N_10446);
nor U10573 (N_10573,N_10477,N_10443);
xnor U10574 (N_10574,N_10417,N_10389);
and U10575 (N_10575,N_10406,N_10377);
xnor U10576 (N_10576,N_10441,N_10436);
nand U10577 (N_10577,N_10419,N_10498);
or U10578 (N_10578,N_10427,N_10399);
or U10579 (N_10579,N_10377,N_10410);
and U10580 (N_10580,N_10432,N_10415);
and U10581 (N_10581,N_10482,N_10421);
nand U10582 (N_10582,N_10419,N_10443);
or U10583 (N_10583,N_10389,N_10448);
nand U10584 (N_10584,N_10483,N_10447);
xnor U10585 (N_10585,N_10376,N_10404);
nand U10586 (N_10586,N_10462,N_10466);
and U10587 (N_10587,N_10469,N_10480);
nor U10588 (N_10588,N_10452,N_10405);
and U10589 (N_10589,N_10450,N_10483);
and U10590 (N_10590,N_10432,N_10482);
or U10591 (N_10591,N_10451,N_10459);
and U10592 (N_10592,N_10392,N_10443);
nand U10593 (N_10593,N_10497,N_10491);
nor U10594 (N_10594,N_10393,N_10414);
and U10595 (N_10595,N_10398,N_10417);
or U10596 (N_10596,N_10414,N_10461);
and U10597 (N_10597,N_10449,N_10469);
nand U10598 (N_10598,N_10426,N_10397);
and U10599 (N_10599,N_10423,N_10410);
nand U10600 (N_10600,N_10451,N_10415);
nor U10601 (N_10601,N_10420,N_10439);
or U10602 (N_10602,N_10439,N_10419);
and U10603 (N_10603,N_10451,N_10463);
nand U10604 (N_10604,N_10390,N_10395);
or U10605 (N_10605,N_10418,N_10484);
or U10606 (N_10606,N_10400,N_10392);
xor U10607 (N_10607,N_10475,N_10431);
or U10608 (N_10608,N_10443,N_10415);
nand U10609 (N_10609,N_10449,N_10411);
and U10610 (N_10610,N_10381,N_10471);
nor U10611 (N_10611,N_10447,N_10489);
and U10612 (N_10612,N_10478,N_10496);
or U10613 (N_10613,N_10428,N_10423);
xor U10614 (N_10614,N_10388,N_10405);
nand U10615 (N_10615,N_10424,N_10474);
or U10616 (N_10616,N_10437,N_10412);
xnor U10617 (N_10617,N_10445,N_10476);
nand U10618 (N_10618,N_10389,N_10453);
nand U10619 (N_10619,N_10449,N_10448);
xor U10620 (N_10620,N_10407,N_10394);
and U10621 (N_10621,N_10486,N_10376);
xor U10622 (N_10622,N_10454,N_10469);
or U10623 (N_10623,N_10486,N_10497);
and U10624 (N_10624,N_10461,N_10380);
xor U10625 (N_10625,N_10605,N_10594);
or U10626 (N_10626,N_10511,N_10623);
xor U10627 (N_10627,N_10555,N_10566);
nand U10628 (N_10628,N_10571,N_10614);
xor U10629 (N_10629,N_10569,N_10548);
xnor U10630 (N_10630,N_10570,N_10535);
xnor U10631 (N_10631,N_10516,N_10596);
nor U10632 (N_10632,N_10556,N_10509);
nand U10633 (N_10633,N_10531,N_10601);
and U10634 (N_10634,N_10587,N_10619);
nand U10635 (N_10635,N_10504,N_10501);
or U10636 (N_10636,N_10550,N_10540);
xnor U10637 (N_10637,N_10591,N_10545);
nor U10638 (N_10638,N_10595,N_10567);
or U10639 (N_10639,N_10607,N_10512);
nand U10640 (N_10640,N_10522,N_10558);
xnor U10641 (N_10641,N_10563,N_10518);
xor U10642 (N_10642,N_10582,N_10617);
nand U10643 (N_10643,N_10610,N_10553);
nand U10644 (N_10644,N_10616,N_10624);
nand U10645 (N_10645,N_10515,N_10552);
nor U10646 (N_10646,N_10621,N_10519);
nand U10647 (N_10647,N_10593,N_10580);
or U10648 (N_10648,N_10573,N_10537);
nand U10649 (N_10649,N_10592,N_10602);
xor U10650 (N_10650,N_10599,N_10529);
nor U10651 (N_10651,N_10579,N_10604);
xnor U10652 (N_10652,N_10603,N_10554);
or U10653 (N_10653,N_10508,N_10533);
nand U10654 (N_10654,N_10576,N_10564);
xor U10655 (N_10655,N_10547,N_10517);
nor U10656 (N_10656,N_10588,N_10532);
and U10657 (N_10657,N_10559,N_10520);
and U10658 (N_10658,N_10590,N_10551);
nor U10659 (N_10659,N_10530,N_10542);
or U10660 (N_10660,N_10502,N_10544);
nand U10661 (N_10661,N_10572,N_10557);
xnor U10662 (N_10662,N_10608,N_10565);
xor U10663 (N_10663,N_10507,N_10525);
nand U10664 (N_10664,N_10612,N_10597);
or U10665 (N_10665,N_10541,N_10589);
xor U10666 (N_10666,N_10514,N_10503);
nor U10667 (N_10667,N_10513,N_10549);
and U10668 (N_10668,N_10534,N_10620);
nand U10669 (N_10669,N_10584,N_10618);
xnor U10670 (N_10670,N_10613,N_10598);
nor U10671 (N_10671,N_10505,N_10609);
nand U10672 (N_10672,N_10561,N_10536);
nor U10673 (N_10673,N_10606,N_10560);
nor U10674 (N_10674,N_10562,N_10615);
xor U10675 (N_10675,N_10586,N_10506);
xnor U10676 (N_10676,N_10543,N_10538);
nor U10677 (N_10677,N_10600,N_10546);
nand U10678 (N_10678,N_10581,N_10575);
xnor U10679 (N_10679,N_10524,N_10521);
or U10680 (N_10680,N_10583,N_10578);
and U10681 (N_10681,N_10568,N_10527);
and U10682 (N_10682,N_10611,N_10526);
nor U10683 (N_10683,N_10585,N_10510);
nor U10684 (N_10684,N_10574,N_10539);
and U10685 (N_10685,N_10577,N_10523);
nand U10686 (N_10686,N_10528,N_10622);
nand U10687 (N_10687,N_10500,N_10591);
or U10688 (N_10688,N_10501,N_10534);
nand U10689 (N_10689,N_10587,N_10518);
xor U10690 (N_10690,N_10540,N_10595);
or U10691 (N_10691,N_10522,N_10518);
nand U10692 (N_10692,N_10542,N_10585);
xor U10693 (N_10693,N_10554,N_10593);
nor U10694 (N_10694,N_10560,N_10615);
nor U10695 (N_10695,N_10620,N_10606);
nand U10696 (N_10696,N_10600,N_10511);
or U10697 (N_10697,N_10559,N_10582);
and U10698 (N_10698,N_10600,N_10517);
nand U10699 (N_10699,N_10548,N_10576);
nor U10700 (N_10700,N_10514,N_10521);
nor U10701 (N_10701,N_10585,N_10562);
nor U10702 (N_10702,N_10548,N_10607);
and U10703 (N_10703,N_10598,N_10510);
xor U10704 (N_10704,N_10506,N_10587);
xor U10705 (N_10705,N_10585,N_10596);
xor U10706 (N_10706,N_10591,N_10515);
nor U10707 (N_10707,N_10562,N_10593);
and U10708 (N_10708,N_10509,N_10615);
or U10709 (N_10709,N_10578,N_10604);
nor U10710 (N_10710,N_10517,N_10561);
and U10711 (N_10711,N_10617,N_10572);
nand U10712 (N_10712,N_10532,N_10524);
xor U10713 (N_10713,N_10511,N_10526);
nand U10714 (N_10714,N_10582,N_10524);
nand U10715 (N_10715,N_10545,N_10602);
or U10716 (N_10716,N_10501,N_10605);
nor U10717 (N_10717,N_10550,N_10530);
xor U10718 (N_10718,N_10589,N_10587);
xor U10719 (N_10719,N_10543,N_10595);
and U10720 (N_10720,N_10598,N_10579);
nor U10721 (N_10721,N_10595,N_10547);
nor U10722 (N_10722,N_10509,N_10603);
and U10723 (N_10723,N_10513,N_10592);
xor U10724 (N_10724,N_10517,N_10540);
or U10725 (N_10725,N_10506,N_10562);
or U10726 (N_10726,N_10616,N_10587);
and U10727 (N_10727,N_10614,N_10560);
or U10728 (N_10728,N_10524,N_10523);
nor U10729 (N_10729,N_10569,N_10564);
nand U10730 (N_10730,N_10545,N_10615);
and U10731 (N_10731,N_10568,N_10604);
xnor U10732 (N_10732,N_10556,N_10618);
xor U10733 (N_10733,N_10538,N_10592);
xnor U10734 (N_10734,N_10597,N_10501);
or U10735 (N_10735,N_10515,N_10599);
or U10736 (N_10736,N_10581,N_10559);
or U10737 (N_10737,N_10504,N_10603);
xnor U10738 (N_10738,N_10560,N_10503);
nor U10739 (N_10739,N_10555,N_10546);
nor U10740 (N_10740,N_10571,N_10530);
or U10741 (N_10741,N_10586,N_10513);
nor U10742 (N_10742,N_10582,N_10560);
xor U10743 (N_10743,N_10525,N_10573);
and U10744 (N_10744,N_10550,N_10570);
xor U10745 (N_10745,N_10511,N_10619);
nor U10746 (N_10746,N_10526,N_10514);
nor U10747 (N_10747,N_10606,N_10596);
xor U10748 (N_10748,N_10566,N_10586);
nand U10749 (N_10749,N_10598,N_10609);
or U10750 (N_10750,N_10676,N_10736);
nor U10751 (N_10751,N_10698,N_10718);
nand U10752 (N_10752,N_10641,N_10679);
nor U10753 (N_10753,N_10643,N_10715);
nand U10754 (N_10754,N_10663,N_10633);
and U10755 (N_10755,N_10658,N_10652);
xor U10756 (N_10756,N_10694,N_10727);
nor U10757 (N_10757,N_10640,N_10739);
xnor U10758 (N_10758,N_10659,N_10677);
xor U10759 (N_10759,N_10725,N_10699);
and U10760 (N_10760,N_10723,N_10668);
nor U10761 (N_10761,N_10701,N_10651);
and U10762 (N_10762,N_10706,N_10708);
and U10763 (N_10763,N_10747,N_10724);
or U10764 (N_10764,N_10630,N_10733);
xnor U10765 (N_10765,N_10683,N_10729);
and U10766 (N_10766,N_10741,N_10732);
and U10767 (N_10767,N_10737,N_10654);
or U10768 (N_10768,N_10673,N_10684);
nor U10769 (N_10769,N_10689,N_10682);
or U10770 (N_10770,N_10656,N_10711);
and U10771 (N_10771,N_10700,N_10707);
and U10772 (N_10772,N_10749,N_10628);
and U10773 (N_10773,N_10647,N_10704);
xnor U10774 (N_10774,N_10692,N_10691);
and U10775 (N_10775,N_10665,N_10639);
xor U10776 (N_10776,N_10657,N_10666);
or U10777 (N_10777,N_10670,N_10645);
and U10778 (N_10778,N_10735,N_10695);
and U10779 (N_10779,N_10710,N_10742);
xor U10780 (N_10780,N_10632,N_10712);
or U10781 (N_10781,N_10703,N_10731);
xnor U10782 (N_10782,N_10675,N_10705);
and U10783 (N_10783,N_10716,N_10728);
or U10784 (N_10784,N_10743,N_10681);
nor U10785 (N_10785,N_10688,N_10746);
and U10786 (N_10786,N_10740,N_10696);
xor U10787 (N_10787,N_10650,N_10713);
nor U10788 (N_10788,N_10634,N_10655);
and U10789 (N_10789,N_10722,N_10672);
and U10790 (N_10790,N_10631,N_10664);
xor U10791 (N_10791,N_10648,N_10626);
xor U10792 (N_10792,N_10636,N_10680);
or U10793 (N_10793,N_10744,N_10669);
nand U10794 (N_10794,N_10745,N_10662);
or U10795 (N_10795,N_10627,N_10660);
xnor U10796 (N_10796,N_10638,N_10720);
xnor U10797 (N_10797,N_10687,N_10748);
nor U10798 (N_10798,N_10674,N_10686);
and U10799 (N_10799,N_10730,N_10693);
xor U10800 (N_10800,N_10709,N_10685);
or U10801 (N_10801,N_10671,N_10667);
xor U10802 (N_10802,N_10629,N_10649);
or U10803 (N_10803,N_10678,N_10635);
nor U10804 (N_10804,N_10726,N_10637);
or U10805 (N_10805,N_10690,N_10734);
and U10806 (N_10806,N_10719,N_10646);
nor U10807 (N_10807,N_10661,N_10697);
or U10808 (N_10808,N_10653,N_10714);
nand U10809 (N_10809,N_10625,N_10642);
nor U10810 (N_10810,N_10721,N_10717);
and U10811 (N_10811,N_10644,N_10702);
and U10812 (N_10812,N_10738,N_10648);
and U10813 (N_10813,N_10745,N_10655);
or U10814 (N_10814,N_10661,N_10724);
xor U10815 (N_10815,N_10692,N_10746);
nor U10816 (N_10816,N_10709,N_10638);
nor U10817 (N_10817,N_10627,N_10625);
nor U10818 (N_10818,N_10680,N_10719);
or U10819 (N_10819,N_10705,N_10708);
nand U10820 (N_10820,N_10743,N_10674);
xor U10821 (N_10821,N_10742,N_10645);
xor U10822 (N_10822,N_10728,N_10735);
nor U10823 (N_10823,N_10666,N_10689);
xor U10824 (N_10824,N_10707,N_10684);
xnor U10825 (N_10825,N_10740,N_10737);
or U10826 (N_10826,N_10714,N_10718);
and U10827 (N_10827,N_10698,N_10703);
nor U10828 (N_10828,N_10731,N_10690);
and U10829 (N_10829,N_10709,N_10732);
or U10830 (N_10830,N_10687,N_10665);
or U10831 (N_10831,N_10740,N_10690);
or U10832 (N_10832,N_10625,N_10740);
nor U10833 (N_10833,N_10666,N_10626);
xor U10834 (N_10834,N_10681,N_10720);
nand U10835 (N_10835,N_10680,N_10707);
and U10836 (N_10836,N_10629,N_10630);
nand U10837 (N_10837,N_10694,N_10698);
xor U10838 (N_10838,N_10730,N_10713);
nand U10839 (N_10839,N_10626,N_10661);
xor U10840 (N_10840,N_10629,N_10719);
or U10841 (N_10841,N_10700,N_10647);
nand U10842 (N_10842,N_10637,N_10657);
nor U10843 (N_10843,N_10661,N_10730);
nor U10844 (N_10844,N_10626,N_10636);
xnor U10845 (N_10845,N_10738,N_10686);
xnor U10846 (N_10846,N_10738,N_10662);
and U10847 (N_10847,N_10734,N_10726);
nor U10848 (N_10848,N_10695,N_10642);
nor U10849 (N_10849,N_10721,N_10742);
nor U10850 (N_10850,N_10653,N_10667);
nand U10851 (N_10851,N_10659,N_10736);
or U10852 (N_10852,N_10726,N_10700);
and U10853 (N_10853,N_10628,N_10684);
nor U10854 (N_10854,N_10662,N_10739);
or U10855 (N_10855,N_10651,N_10644);
nand U10856 (N_10856,N_10638,N_10625);
nor U10857 (N_10857,N_10636,N_10724);
nand U10858 (N_10858,N_10626,N_10659);
nand U10859 (N_10859,N_10733,N_10714);
nor U10860 (N_10860,N_10649,N_10698);
and U10861 (N_10861,N_10740,N_10708);
or U10862 (N_10862,N_10704,N_10742);
xnor U10863 (N_10863,N_10656,N_10747);
nor U10864 (N_10864,N_10695,N_10663);
nor U10865 (N_10865,N_10678,N_10713);
or U10866 (N_10866,N_10734,N_10642);
nand U10867 (N_10867,N_10717,N_10697);
or U10868 (N_10868,N_10742,N_10667);
nand U10869 (N_10869,N_10656,N_10676);
xnor U10870 (N_10870,N_10641,N_10724);
and U10871 (N_10871,N_10696,N_10723);
xor U10872 (N_10872,N_10736,N_10687);
xnor U10873 (N_10873,N_10694,N_10724);
nand U10874 (N_10874,N_10723,N_10660);
nor U10875 (N_10875,N_10846,N_10784);
nor U10876 (N_10876,N_10851,N_10778);
xnor U10877 (N_10877,N_10759,N_10762);
nand U10878 (N_10878,N_10870,N_10869);
xor U10879 (N_10879,N_10837,N_10764);
nand U10880 (N_10880,N_10821,N_10841);
nand U10881 (N_10881,N_10753,N_10835);
or U10882 (N_10882,N_10838,N_10810);
and U10883 (N_10883,N_10751,N_10771);
nor U10884 (N_10884,N_10830,N_10871);
nand U10885 (N_10885,N_10789,N_10832);
and U10886 (N_10886,N_10772,N_10842);
nand U10887 (N_10887,N_10807,N_10786);
or U10888 (N_10888,N_10819,N_10858);
nand U10889 (N_10889,N_10791,N_10792);
nand U10890 (N_10890,N_10813,N_10844);
nor U10891 (N_10891,N_10783,N_10775);
and U10892 (N_10892,N_10845,N_10864);
and U10893 (N_10893,N_10754,N_10800);
nand U10894 (N_10894,N_10794,N_10799);
nor U10895 (N_10895,N_10782,N_10822);
or U10896 (N_10896,N_10849,N_10809);
xnor U10897 (N_10897,N_10761,N_10826);
nand U10898 (N_10898,N_10797,N_10860);
and U10899 (N_10899,N_10866,N_10769);
xnor U10900 (N_10900,N_10820,N_10863);
nor U10901 (N_10901,N_10779,N_10833);
nor U10902 (N_10902,N_10755,N_10847);
and U10903 (N_10903,N_10834,N_10788);
or U10904 (N_10904,N_10859,N_10867);
and U10905 (N_10905,N_10758,N_10768);
and U10906 (N_10906,N_10812,N_10806);
or U10907 (N_10907,N_10840,N_10774);
nand U10908 (N_10908,N_10750,N_10767);
xor U10909 (N_10909,N_10843,N_10781);
nand U10910 (N_10910,N_10857,N_10852);
and U10911 (N_10911,N_10773,N_10856);
or U10912 (N_10912,N_10823,N_10793);
xor U10913 (N_10913,N_10829,N_10831);
nor U10914 (N_10914,N_10802,N_10785);
and U10915 (N_10915,N_10872,N_10865);
nand U10916 (N_10916,N_10853,N_10763);
nand U10917 (N_10917,N_10854,N_10874);
xnor U10918 (N_10918,N_10776,N_10862);
nor U10919 (N_10919,N_10868,N_10825);
or U10920 (N_10920,N_10795,N_10796);
nor U10921 (N_10921,N_10836,N_10766);
xor U10922 (N_10922,N_10815,N_10839);
xor U10923 (N_10923,N_10818,N_10805);
and U10924 (N_10924,N_10855,N_10765);
and U10925 (N_10925,N_10752,N_10780);
nand U10926 (N_10926,N_10801,N_10848);
or U10927 (N_10927,N_10811,N_10824);
and U10928 (N_10928,N_10787,N_10828);
nand U10929 (N_10929,N_10816,N_10861);
nor U10930 (N_10930,N_10777,N_10756);
nor U10931 (N_10931,N_10817,N_10827);
nand U10932 (N_10932,N_10790,N_10804);
nand U10933 (N_10933,N_10808,N_10814);
xor U10934 (N_10934,N_10760,N_10850);
xor U10935 (N_10935,N_10770,N_10798);
nor U10936 (N_10936,N_10757,N_10803);
or U10937 (N_10937,N_10873,N_10772);
xnor U10938 (N_10938,N_10815,N_10819);
nand U10939 (N_10939,N_10837,N_10754);
nor U10940 (N_10940,N_10795,N_10791);
nand U10941 (N_10941,N_10777,N_10770);
and U10942 (N_10942,N_10750,N_10764);
xor U10943 (N_10943,N_10859,N_10813);
nor U10944 (N_10944,N_10771,N_10823);
or U10945 (N_10945,N_10775,N_10820);
nor U10946 (N_10946,N_10770,N_10750);
xor U10947 (N_10947,N_10831,N_10827);
xor U10948 (N_10948,N_10868,N_10797);
xor U10949 (N_10949,N_10836,N_10871);
nor U10950 (N_10950,N_10765,N_10851);
or U10951 (N_10951,N_10774,N_10805);
or U10952 (N_10952,N_10787,N_10842);
nor U10953 (N_10953,N_10873,N_10836);
and U10954 (N_10954,N_10859,N_10796);
or U10955 (N_10955,N_10865,N_10861);
nor U10956 (N_10956,N_10753,N_10807);
xor U10957 (N_10957,N_10814,N_10765);
xnor U10958 (N_10958,N_10850,N_10827);
or U10959 (N_10959,N_10782,N_10846);
nand U10960 (N_10960,N_10792,N_10865);
nor U10961 (N_10961,N_10778,N_10772);
xor U10962 (N_10962,N_10812,N_10864);
or U10963 (N_10963,N_10827,N_10759);
nand U10964 (N_10964,N_10869,N_10813);
nand U10965 (N_10965,N_10773,N_10822);
or U10966 (N_10966,N_10874,N_10780);
nand U10967 (N_10967,N_10869,N_10799);
and U10968 (N_10968,N_10874,N_10830);
xnor U10969 (N_10969,N_10760,N_10845);
nand U10970 (N_10970,N_10841,N_10796);
xor U10971 (N_10971,N_10861,N_10780);
xnor U10972 (N_10972,N_10816,N_10763);
xor U10973 (N_10973,N_10778,N_10850);
xnor U10974 (N_10974,N_10870,N_10834);
nand U10975 (N_10975,N_10768,N_10770);
xor U10976 (N_10976,N_10806,N_10765);
or U10977 (N_10977,N_10762,N_10754);
nor U10978 (N_10978,N_10854,N_10758);
or U10979 (N_10979,N_10767,N_10851);
xnor U10980 (N_10980,N_10872,N_10820);
and U10981 (N_10981,N_10867,N_10803);
xor U10982 (N_10982,N_10863,N_10762);
nand U10983 (N_10983,N_10867,N_10872);
nand U10984 (N_10984,N_10787,N_10798);
and U10985 (N_10985,N_10845,N_10865);
and U10986 (N_10986,N_10819,N_10804);
or U10987 (N_10987,N_10762,N_10831);
and U10988 (N_10988,N_10840,N_10788);
and U10989 (N_10989,N_10765,N_10860);
xor U10990 (N_10990,N_10870,N_10824);
xnor U10991 (N_10991,N_10811,N_10791);
nor U10992 (N_10992,N_10799,N_10808);
or U10993 (N_10993,N_10802,N_10831);
nor U10994 (N_10994,N_10847,N_10799);
xnor U10995 (N_10995,N_10822,N_10789);
nand U10996 (N_10996,N_10820,N_10833);
and U10997 (N_10997,N_10800,N_10855);
and U10998 (N_10998,N_10780,N_10787);
nand U10999 (N_10999,N_10771,N_10816);
nor U11000 (N_11000,N_10965,N_10962);
and U11001 (N_11001,N_10890,N_10998);
nand U11002 (N_11002,N_10981,N_10925);
xor U11003 (N_11003,N_10964,N_10944);
nor U11004 (N_11004,N_10875,N_10967);
nor U11005 (N_11005,N_10909,N_10969);
or U11006 (N_11006,N_10942,N_10896);
nand U11007 (N_11007,N_10882,N_10899);
and U11008 (N_11008,N_10958,N_10968);
nor U11009 (N_11009,N_10892,N_10986);
and U11010 (N_11010,N_10917,N_10881);
nand U11011 (N_11011,N_10966,N_10889);
and U11012 (N_11012,N_10979,N_10976);
nor U11013 (N_11013,N_10915,N_10898);
or U11014 (N_11014,N_10949,N_10959);
nand U11015 (N_11015,N_10895,N_10891);
xnor U11016 (N_11016,N_10930,N_10888);
or U11017 (N_11017,N_10957,N_10975);
nor U11018 (N_11018,N_10938,N_10940);
nor U11019 (N_11019,N_10948,N_10877);
or U11020 (N_11020,N_10906,N_10950);
or U11021 (N_11021,N_10912,N_10982);
nand U11022 (N_11022,N_10903,N_10947);
nand U11023 (N_11023,N_10955,N_10920);
nor U11024 (N_11024,N_10910,N_10988);
xor U11025 (N_11025,N_10902,N_10886);
xor U11026 (N_11026,N_10914,N_10887);
nor U11027 (N_11027,N_10922,N_10943);
nand U11028 (N_11028,N_10946,N_10921);
and U11029 (N_11029,N_10876,N_10977);
nor U11030 (N_11030,N_10913,N_10945);
nor U11031 (N_11031,N_10901,N_10960);
nand U11032 (N_11032,N_10918,N_10932);
and U11033 (N_11033,N_10991,N_10905);
and U11034 (N_11034,N_10992,N_10908);
nand U11035 (N_11035,N_10941,N_10884);
and U11036 (N_11036,N_10973,N_10936);
nor U11037 (N_11037,N_10924,N_10972);
and U11038 (N_11038,N_10935,N_10984);
xnor U11039 (N_11039,N_10907,N_10993);
and U11040 (N_11040,N_10983,N_10927);
nor U11041 (N_11041,N_10954,N_10971);
xnor U11042 (N_11042,N_10897,N_10952);
xnor U11043 (N_11043,N_10923,N_10963);
nor U11044 (N_11044,N_10926,N_10961);
and U11045 (N_11045,N_10995,N_10880);
and U11046 (N_11046,N_10893,N_10919);
nor U11047 (N_11047,N_10997,N_10900);
and U11048 (N_11048,N_10994,N_10974);
nand U11049 (N_11049,N_10934,N_10970);
and U11050 (N_11050,N_10980,N_10937);
nand U11051 (N_11051,N_10883,N_10951);
nor U11052 (N_11052,N_10878,N_10987);
nand U11053 (N_11053,N_10928,N_10916);
and U11054 (N_11054,N_10879,N_10989);
nor U11055 (N_11055,N_10985,N_10904);
and U11056 (N_11056,N_10911,N_10929);
xnor U11057 (N_11057,N_10956,N_10978);
or U11058 (N_11058,N_10885,N_10999);
nor U11059 (N_11059,N_10939,N_10894);
nor U11060 (N_11060,N_10953,N_10931);
nand U11061 (N_11061,N_10990,N_10996);
or U11062 (N_11062,N_10933,N_10927);
nor U11063 (N_11063,N_10971,N_10992);
nor U11064 (N_11064,N_10910,N_10904);
and U11065 (N_11065,N_10960,N_10972);
and U11066 (N_11066,N_10950,N_10991);
nand U11067 (N_11067,N_10960,N_10917);
nor U11068 (N_11068,N_10909,N_10985);
nor U11069 (N_11069,N_10961,N_10899);
nor U11070 (N_11070,N_10994,N_10937);
or U11071 (N_11071,N_10918,N_10911);
or U11072 (N_11072,N_10987,N_10972);
and U11073 (N_11073,N_10929,N_10932);
and U11074 (N_11074,N_10913,N_10924);
xnor U11075 (N_11075,N_10920,N_10960);
xor U11076 (N_11076,N_10918,N_10927);
xnor U11077 (N_11077,N_10931,N_10963);
or U11078 (N_11078,N_10996,N_10973);
nand U11079 (N_11079,N_10953,N_10876);
nor U11080 (N_11080,N_10880,N_10922);
or U11081 (N_11081,N_10970,N_10936);
nand U11082 (N_11082,N_10962,N_10993);
nand U11083 (N_11083,N_10977,N_10933);
and U11084 (N_11084,N_10916,N_10935);
nor U11085 (N_11085,N_10983,N_10948);
nor U11086 (N_11086,N_10895,N_10888);
and U11087 (N_11087,N_10994,N_10990);
nor U11088 (N_11088,N_10948,N_10911);
xnor U11089 (N_11089,N_10970,N_10883);
and U11090 (N_11090,N_10983,N_10884);
xnor U11091 (N_11091,N_10940,N_10892);
nand U11092 (N_11092,N_10994,N_10880);
and U11093 (N_11093,N_10958,N_10885);
nor U11094 (N_11094,N_10997,N_10975);
or U11095 (N_11095,N_10883,N_10888);
xnor U11096 (N_11096,N_10914,N_10969);
nor U11097 (N_11097,N_10915,N_10978);
nor U11098 (N_11098,N_10959,N_10937);
and U11099 (N_11099,N_10921,N_10934);
and U11100 (N_11100,N_10885,N_10978);
and U11101 (N_11101,N_10910,N_10995);
and U11102 (N_11102,N_10928,N_10990);
and U11103 (N_11103,N_10878,N_10904);
nor U11104 (N_11104,N_10934,N_10982);
xnor U11105 (N_11105,N_10967,N_10937);
and U11106 (N_11106,N_10888,N_10973);
and U11107 (N_11107,N_10948,N_10941);
nor U11108 (N_11108,N_10942,N_10959);
nor U11109 (N_11109,N_10984,N_10932);
nor U11110 (N_11110,N_10949,N_10974);
xor U11111 (N_11111,N_10965,N_10892);
or U11112 (N_11112,N_10933,N_10931);
and U11113 (N_11113,N_10936,N_10952);
and U11114 (N_11114,N_10895,N_10973);
or U11115 (N_11115,N_10982,N_10956);
xnor U11116 (N_11116,N_10990,N_10893);
and U11117 (N_11117,N_10888,N_10897);
and U11118 (N_11118,N_10994,N_10919);
and U11119 (N_11119,N_10913,N_10903);
xor U11120 (N_11120,N_10905,N_10943);
nor U11121 (N_11121,N_10952,N_10913);
nor U11122 (N_11122,N_10984,N_10900);
nor U11123 (N_11123,N_10988,N_10941);
and U11124 (N_11124,N_10894,N_10922);
or U11125 (N_11125,N_11077,N_11032);
and U11126 (N_11126,N_11062,N_11084);
xor U11127 (N_11127,N_11031,N_11116);
nor U11128 (N_11128,N_11118,N_11010);
nor U11129 (N_11129,N_11053,N_11028);
nor U11130 (N_11130,N_11026,N_11042);
nor U11131 (N_11131,N_11112,N_11021);
nor U11132 (N_11132,N_11078,N_11067);
nor U11133 (N_11133,N_11117,N_11040);
xnor U11134 (N_11134,N_11074,N_11041);
nand U11135 (N_11135,N_11047,N_11065);
nand U11136 (N_11136,N_11049,N_11098);
nor U11137 (N_11137,N_11099,N_11105);
nand U11138 (N_11138,N_11064,N_11106);
or U11139 (N_11139,N_11001,N_11109);
xnor U11140 (N_11140,N_11006,N_11070);
nand U11141 (N_11141,N_11058,N_11017);
nand U11142 (N_11142,N_11072,N_11056);
and U11143 (N_11143,N_11079,N_11073);
nor U11144 (N_11144,N_11108,N_11027);
xnor U11145 (N_11145,N_11124,N_11055);
and U11146 (N_11146,N_11060,N_11110);
nor U11147 (N_11147,N_11013,N_11069);
xnor U11148 (N_11148,N_11014,N_11089);
xnor U11149 (N_11149,N_11059,N_11083);
and U11150 (N_11150,N_11051,N_11066);
xor U11151 (N_11151,N_11095,N_11046);
nand U11152 (N_11152,N_11113,N_11029);
or U11153 (N_11153,N_11020,N_11088);
nand U11154 (N_11154,N_11091,N_11024);
and U11155 (N_11155,N_11087,N_11075);
xnor U11156 (N_11156,N_11121,N_11008);
nand U11157 (N_11157,N_11036,N_11022);
or U11158 (N_11158,N_11016,N_11096);
nor U11159 (N_11159,N_11018,N_11103);
nor U11160 (N_11160,N_11035,N_11052);
and U11161 (N_11161,N_11063,N_11044);
and U11162 (N_11162,N_11080,N_11054);
nand U11163 (N_11163,N_11033,N_11114);
and U11164 (N_11164,N_11115,N_11025);
xnor U11165 (N_11165,N_11005,N_11094);
nand U11166 (N_11166,N_11002,N_11071);
nand U11167 (N_11167,N_11043,N_11004);
nand U11168 (N_11168,N_11011,N_11107);
nand U11169 (N_11169,N_11097,N_11038);
or U11170 (N_11170,N_11102,N_11061);
or U11171 (N_11171,N_11023,N_11076);
xor U11172 (N_11172,N_11050,N_11122);
nand U11173 (N_11173,N_11086,N_11068);
nand U11174 (N_11174,N_11093,N_11048);
and U11175 (N_11175,N_11120,N_11003);
xnor U11176 (N_11176,N_11009,N_11101);
xor U11177 (N_11177,N_11037,N_11034);
nand U11178 (N_11178,N_11039,N_11100);
and U11179 (N_11179,N_11019,N_11012);
xor U11180 (N_11180,N_11085,N_11000);
or U11181 (N_11181,N_11030,N_11092);
xor U11182 (N_11182,N_11111,N_11007);
or U11183 (N_11183,N_11104,N_11015);
nand U11184 (N_11184,N_11081,N_11045);
or U11185 (N_11185,N_11123,N_11119);
nor U11186 (N_11186,N_11090,N_11057);
nand U11187 (N_11187,N_11082,N_11081);
or U11188 (N_11188,N_11050,N_11106);
nand U11189 (N_11189,N_11111,N_11084);
nand U11190 (N_11190,N_11113,N_11058);
or U11191 (N_11191,N_11114,N_11059);
nand U11192 (N_11192,N_11109,N_11014);
nor U11193 (N_11193,N_11003,N_11022);
xnor U11194 (N_11194,N_11010,N_11042);
xnor U11195 (N_11195,N_11113,N_11112);
xnor U11196 (N_11196,N_11002,N_11093);
nand U11197 (N_11197,N_11040,N_11092);
or U11198 (N_11198,N_11068,N_11028);
xor U11199 (N_11199,N_11036,N_11099);
and U11200 (N_11200,N_11066,N_11077);
and U11201 (N_11201,N_11043,N_11058);
or U11202 (N_11202,N_11008,N_11123);
or U11203 (N_11203,N_11001,N_11008);
xor U11204 (N_11204,N_11003,N_11068);
nor U11205 (N_11205,N_11102,N_11085);
nor U11206 (N_11206,N_11007,N_11041);
nand U11207 (N_11207,N_11065,N_11021);
and U11208 (N_11208,N_11004,N_11061);
or U11209 (N_11209,N_11042,N_11066);
xnor U11210 (N_11210,N_11102,N_11119);
and U11211 (N_11211,N_11033,N_11022);
and U11212 (N_11212,N_11121,N_11097);
and U11213 (N_11213,N_11081,N_11095);
xor U11214 (N_11214,N_11025,N_11026);
or U11215 (N_11215,N_11097,N_11004);
nand U11216 (N_11216,N_11020,N_11081);
xnor U11217 (N_11217,N_11028,N_11083);
and U11218 (N_11218,N_11083,N_11085);
nor U11219 (N_11219,N_11062,N_11053);
nor U11220 (N_11220,N_11114,N_11049);
nor U11221 (N_11221,N_11071,N_11094);
and U11222 (N_11222,N_11061,N_11076);
nor U11223 (N_11223,N_11092,N_11036);
nor U11224 (N_11224,N_11025,N_11102);
nand U11225 (N_11225,N_11087,N_11092);
xnor U11226 (N_11226,N_11121,N_11116);
and U11227 (N_11227,N_11004,N_11036);
or U11228 (N_11228,N_11094,N_11054);
and U11229 (N_11229,N_11078,N_11028);
nor U11230 (N_11230,N_11053,N_11080);
nand U11231 (N_11231,N_11108,N_11012);
nand U11232 (N_11232,N_11103,N_11005);
and U11233 (N_11233,N_11065,N_11040);
and U11234 (N_11234,N_11040,N_11024);
nand U11235 (N_11235,N_11060,N_11001);
and U11236 (N_11236,N_11017,N_11075);
xor U11237 (N_11237,N_11121,N_11102);
xor U11238 (N_11238,N_11083,N_11008);
and U11239 (N_11239,N_11080,N_11068);
or U11240 (N_11240,N_11018,N_11005);
xnor U11241 (N_11241,N_11101,N_11051);
nand U11242 (N_11242,N_11118,N_11039);
nor U11243 (N_11243,N_11064,N_11107);
xor U11244 (N_11244,N_11068,N_11090);
or U11245 (N_11245,N_11094,N_11084);
or U11246 (N_11246,N_11030,N_11038);
or U11247 (N_11247,N_11117,N_11048);
xor U11248 (N_11248,N_11003,N_11093);
nand U11249 (N_11249,N_11096,N_11075);
nor U11250 (N_11250,N_11249,N_11133);
or U11251 (N_11251,N_11242,N_11233);
xnor U11252 (N_11252,N_11140,N_11135);
or U11253 (N_11253,N_11162,N_11223);
or U11254 (N_11254,N_11149,N_11218);
xnor U11255 (N_11255,N_11136,N_11211);
and U11256 (N_11256,N_11175,N_11198);
or U11257 (N_11257,N_11232,N_11195);
xor U11258 (N_11258,N_11204,N_11182);
and U11259 (N_11259,N_11156,N_11125);
xnor U11260 (N_11260,N_11222,N_11200);
and U11261 (N_11261,N_11164,N_11228);
nor U11262 (N_11262,N_11235,N_11247);
and U11263 (N_11263,N_11188,N_11181);
xor U11264 (N_11264,N_11146,N_11152);
xor U11265 (N_11265,N_11183,N_11141);
nand U11266 (N_11266,N_11214,N_11206);
and U11267 (N_11267,N_11166,N_11194);
and U11268 (N_11268,N_11209,N_11159);
and U11269 (N_11269,N_11187,N_11173);
nor U11270 (N_11270,N_11155,N_11126);
or U11271 (N_11271,N_11150,N_11216);
or U11272 (N_11272,N_11205,N_11158);
nand U11273 (N_11273,N_11170,N_11132);
or U11274 (N_11274,N_11229,N_11221);
nand U11275 (N_11275,N_11134,N_11192);
xnor U11276 (N_11276,N_11178,N_11203);
or U11277 (N_11277,N_11227,N_11189);
and U11278 (N_11278,N_11185,N_11210);
and U11279 (N_11279,N_11163,N_11193);
xnor U11280 (N_11280,N_11239,N_11202);
nor U11281 (N_11281,N_11236,N_11248);
nor U11282 (N_11282,N_11245,N_11143);
or U11283 (N_11283,N_11246,N_11190);
xnor U11284 (N_11284,N_11168,N_11167);
xnor U11285 (N_11285,N_11176,N_11213);
or U11286 (N_11286,N_11180,N_11174);
and U11287 (N_11287,N_11244,N_11196);
xnor U11288 (N_11288,N_11240,N_11197);
xor U11289 (N_11289,N_11231,N_11160);
and U11290 (N_11290,N_11165,N_11142);
xor U11291 (N_11291,N_11243,N_11148);
and U11292 (N_11292,N_11208,N_11238);
and U11293 (N_11293,N_11147,N_11138);
nand U11294 (N_11294,N_11230,N_11207);
nand U11295 (N_11295,N_11220,N_11130);
xnor U11296 (N_11296,N_11169,N_11153);
or U11297 (N_11297,N_11241,N_11226);
or U11298 (N_11298,N_11217,N_11128);
xnor U11299 (N_11299,N_11199,N_11131);
or U11300 (N_11300,N_11144,N_11215);
xor U11301 (N_11301,N_11219,N_11137);
xnor U11302 (N_11302,N_11139,N_11129);
xnor U11303 (N_11303,N_11184,N_11145);
or U11304 (N_11304,N_11186,N_11191);
and U11305 (N_11305,N_11237,N_11212);
and U11306 (N_11306,N_11161,N_11225);
and U11307 (N_11307,N_11224,N_11201);
xnor U11308 (N_11308,N_11154,N_11151);
xor U11309 (N_11309,N_11234,N_11177);
and U11310 (N_11310,N_11171,N_11172);
nand U11311 (N_11311,N_11127,N_11179);
nor U11312 (N_11312,N_11157,N_11247);
xor U11313 (N_11313,N_11223,N_11246);
nand U11314 (N_11314,N_11179,N_11130);
nand U11315 (N_11315,N_11160,N_11165);
nor U11316 (N_11316,N_11137,N_11181);
xnor U11317 (N_11317,N_11141,N_11247);
and U11318 (N_11318,N_11218,N_11165);
and U11319 (N_11319,N_11227,N_11147);
xnor U11320 (N_11320,N_11190,N_11154);
nor U11321 (N_11321,N_11181,N_11189);
or U11322 (N_11322,N_11162,N_11220);
xor U11323 (N_11323,N_11145,N_11179);
xor U11324 (N_11324,N_11165,N_11246);
xor U11325 (N_11325,N_11177,N_11219);
and U11326 (N_11326,N_11220,N_11238);
and U11327 (N_11327,N_11141,N_11245);
or U11328 (N_11328,N_11232,N_11179);
and U11329 (N_11329,N_11220,N_11185);
or U11330 (N_11330,N_11203,N_11143);
nor U11331 (N_11331,N_11222,N_11205);
nand U11332 (N_11332,N_11125,N_11146);
or U11333 (N_11333,N_11223,N_11242);
or U11334 (N_11334,N_11147,N_11136);
or U11335 (N_11335,N_11173,N_11127);
nor U11336 (N_11336,N_11241,N_11221);
nand U11337 (N_11337,N_11132,N_11202);
nand U11338 (N_11338,N_11195,N_11230);
and U11339 (N_11339,N_11247,N_11161);
nor U11340 (N_11340,N_11145,N_11183);
nand U11341 (N_11341,N_11131,N_11126);
xnor U11342 (N_11342,N_11211,N_11194);
or U11343 (N_11343,N_11174,N_11221);
xnor U11344 (N_11344,N_11184,N_11151);
nand U11345 (N_11345,N_11165,N_11239);
nand U11346 (N_11346,N_11148,N_11168);
xor U11347 (N_11347,N_11233,N_11138);
xor U11348 (N_11348,N_11187,N_11127);
and U11349 (N_11349,N_11177,N_11235);
nor U11350 (N_11350,N_11235,N_11237);
nand U11351 (N_11351,N_11221,N_11237);
or U11352 (N_11352,N_11163,N_11126);
and U11353 (N_11353,N_11196,N_11182);
nor U11354 (N_11354,N_11210,N_11169);
nand U11355 (N_11355,N_11246,N_11243);
xnor U11356 (N_11356,N_11227,N_11156);
nor U11357 (N_11357,N_11128,N_11245);
or U11358 (N_11358,N_11141,N_11225);
nor U11359 (N_11359,N_11126,N_11147);
or U11360 (N_11360,N_11220,N_11151);
nor U11361 (N_11361,N_11142,N_11213);
or U11362 (N_11362,N_11249,N_11179);
nor U11363 (N_11363,N_11148,N_11245);
and U11364 (N_11364,N_11159,N_11244);
xor U11365 (N_11365,N_11169,N_11199);
and U11366 (N_11366,N_11180,N_11205);
nand U11367 (N_11367,N_11198,N_11150);
or U11368 (N_11368,N_11220,N_11232);
or U11369 (N_11369,N_11178,N_11226);
nand U11370 (N_11370,N_11249,N_11136);
or U11371 (N_11371,N_11208,N_11135);
nand U11372 (N_11372,N_11187,N_11167);
nor U11373 (N_11373,N_11149,N_11181);
or U11374 (N_11374,N_11172,N_11203);
and U11375 (N_11375,N_11267,N_11252);
nand U11376 (N_11376,N_11262,N_11305);
xor U11377 (N_11377,N_11329,N_11296);
or U11378 (N_11378,N_11328,N_11338);
or U11379 (N_11379,N_11359,N_11287);
nor U11380 (N_11380,N_11302,N_11347);
xor U11381 (N_11381,N_11276,N_11318);
nor U11382 (N_11382,N_11278,N_11324);
and U11383 (N_11383,N_11350,N_11259);
and U11384 (N_11384,N_11360,N_11367);
nand U11385 (N_11385,N_11283,N_11269);
xor U11386 (N_11386,N_11357,N_11321);
or U11387 (N_11387,N_11280,N_11343);
and U11388 (N_11388,N_11340,N_11342);
xnor U11389 (N_11389,N_11313,N_11284);
nand U11390 (N_11390,N_11282,N_11348);
xor U11391 (N_11391,N_11295,N_11326);
xor U11392 (N_11392,N_11257,N_11277);
or U11393 (N_11393,N_11286,N_11292);
or U11394 (N_11394,N_11306,N_11251);
and U11395 (N_11395,N_11345,N_11346);
or U11396 (N_11396,N_11341,N_11304);
and U11397 (N_11397,N_11355,N_11322);
nand U11398 (N_11398,N_11311,N_11250);
nor U11399 (N_11399,N_11288,N_11331);
nor U11400 (N_11400,N_11279,N_11281);
xnor U11401 (N_11401,N_11291,N_11319);
xnor U11402 (N_11402,N_11293,N_11330);
and U11403 (N_11403,N_11371,N_11351);
nor U11404 (N_11404,N_11364,N_11316);
or U11405 (N_11405,N_11258,N_11320);
and U11406 (N_11406,N_11356,N_11374);
or U11407 (N_11407,N_11264,N_11323);
xor U11408 (N_11408,N_11307,N_11294);
nand U11409 (N_11409,N_11298,N_11362);
xor U11410 (N_11410,N_11266,N_11370);
nand U11411 (N_11411,N_11361,N_11336);
nor U11412 (N_11412,N_11312,N_11349);
and U11413 (N_11413,N_11285,N_11272);
or U11414 (N_11414,N_11315,N_11301);
nor U11415 (N_11415,N_11274,N_11344);
and U11416 (N_11416,N_11325,N_11354);
or U11417 (N_11417,N_11337,N_11365);
nor U11418 (N_11418,N_11297,N_11373);
or U11419 (N_11419,N_11372,N_11309);
and U11420 (N_11420,N_11308,N_11368);
nor U11421 (N_11421,N_11335,N_11260);
xor U11422 (N_11422,N_11256,N_11273);
nand U11423 (N_11423,N_11314,N_11339);
and U11424 (N_11424,N_11299,N_11363);
and U11425 (N_11425,N_11333,N_11327);
nand U11426 (N_11426,N_11369,N_11263);
nand U11427 (N_11427,N_11268,N_11265);
and U11428 (N_11428,N_11270,N_11366);
nand U11429 (N_11429,N_11303,N_11253);
xor U11430 (N_11430,N_11271,N_11254);
nor U11431 (N_11431,N_11332,N_11289);
and U11432 (N_11432,N_11255,N_11300);
xnor U11433 (N_11433,N_11310,N_11275);
and U11434 (N_11434,N_11317,N_11358);
nand U11435 (N_11435,N_11353,N_11334);
or U11436 (N_11436,N_11290,N_11261);
nor U11437 (N_11437,N_11352,N_11274);
xnor U11438 (N_11438,N_11334,N_11369);
nor U11439 (N_11439,N_11373,N_11306);
xor U11440 (N_11440,N_11358,N_11366);
nor U11441 (N_11441,N_11288,N_11268);
or U11442 (N_11442,N_11334,N_11288);
and U11443 (N_11443,N_11258,N_11310);
nand U11444 (N_11444,N_11253,N_11346);
and U11445 (N_11445,N_11347,N_11355);
nor U11446 (N_11446,N_11300,N_11374);
nor U11447 (N_11447,N_11346,N_11357);
and U11448 (N_11448,N_11320,N_11279);
xnor U11449 (N_11449,N_11335,N_11323);
and U11450 (N_11450,N_11346,N_11372);
or U11451 (N_11451,N_11344,N_11254);
xnor U11452 (N_11452,N_11364,N_11363);
nand U11453 (N_11453,N_11344,N_11315);
or U11454 (N_11454,N_11310,N_11306);
nor U11455 (N_11455,N_11351,N_11302);
nor U11456 (N_11456,N_11251,N_11298);
and U11457 (N_11457,N_11347,N_11273);
and U11458 (N_11458,N_11320,N_11351);
nor U11459 (N_11459,N_11339,N_11352);
nand U11460 (N_11460,N_11358,N_11348);
xor U11461 (N_11461,N_11259,N_11320);
nor U11462 (N_11462,N_11323,N_11289);
xnor U11463 (N_11463,N_11309,N_11259);
xor U11464 (N_11464,N_11354,N_11369);
nand U11465 (N_11465,N_11359,N_11367);
or U11466 (N_11466,N_11284,N_11267);
nand U11467 (N_11467,N_11342,N_11250);
and U11468 (N_11468,N_11364,N_11303);
or U11469 (N_11469,N_11353,N_11333);
or U11470 (N_11470,N_11330,N_11326);
nand U11471 (N_11471,N_11288,N_11359);
xnor U11472 (N_11472,N_11291,N_11283);
or U11473 (N_11473,N_11281,N_11292);
nor U11474 (N_11474,N_11274,N_11272);
and U11475 (N_11475,N_11286,N_11342);
nor U11476 (N_11476,N_11261,N_11319);
or U11477 (N_11477,N_11321,N_11256);
nor U11478 (N_11478,N_11265,N_11325);
xor U11479 (N_11479,N_11367,N_11364);
and U11480 (N_11480,N_11374,N_11304);
or U11481 (N_11481,N_11274,N_11321);
nand U11482 (N_11482,N_11300,N_11317);
xnor U11483 (N_11483,N_11335,N_11272);
nor U11484 (N_11484,N_11347,N_11374);
or U11485 (N_11485,N_11324,N_11251);
nor U11486 (N_11486,N_11343,N_11294);
xor U11487 (N_11487,N_11258,N_11287);
nand U11488 (N_11488,N_11263,N_11326);
xnor U11489 (N_11489,N_11310,N_11340);
or U11490 (N_11490,N_11270,N_11340);
nand U11491 (N_11491,N_11322,N_11349);
or U11492 (N_11492,N_11279,N_11261);
and U11493 (N_11493,N_11290,N_11352);
nor U11494 (N_11494,N_11263,N_11287);
xnor U11495 (N_11495,N_11309,N_11317);
xor U11496 (N_11496,N_11288,N_11314);
or U11497 (N_11497,N_11276,N_11321);
or U11498 (N_11498,N_11346,N_11307);
and U11499 (N_11499,N_11344,N_11266);
and U11500 (N_11500,N_11404,N_11387);
and U11501 (N_11501,N_11455,N_11451);
nor U11502 (N_11502,N_11446,N_11495);
and U11503 (N_11503,N_11435,N_11478);
xor U11504 (N_11504,N_11411,N_11497);
and U11505 (N_11505,N_11479,N_11381);
nor U11506 (N_11506,N_11484,N_11471);
nand U11507 (N_11507,N_11469,N_11406);
nand U11508 (N_11508,N_11481,N_11475);
and U11509 (N_11509,N_11379,N_11419);
nand U11510 (N_11510,N_11492,N_11499);
xnor U11511 (N_11511,N_11483,N_11383);
nand U11512 (N_11512,N_11456,N_11422);
xnor U11513 (N_11513,N_11498,N_11477);
and U11514 (N_11514,N_11449,N_11377);
nor U11515 (N_11515,N_11382,N_11418);
or U11516 (N_11516,N_11460,N_11450);
and U11517 (N_11517,N_11392,N_11413);
nand U11518 (N_11518,N_11417,N_11488);
or U11519 (N_11519,N_11490,N_11416);
or U11520 (N_11520,N_11496,N_11453);
nor U11521 (N_11521,N_11423,N_11461);
xnor U11522 (N_11522,N_11428,N_11421);
xnor U11523 (N_11523,N_11427,N_11468);
and U11524 (N_11524,N_11443,N_11409);
nand U11525 (N_11525,N_11440,N_11396);
nand U11526 (N_11526,N_11486,N_11410);
nand U11527 (N_11527,N_11459,N_11414);
and U11528 (N_11528,N_11431,N_11425);
nand U11529 (N_11529,N_11395,N_11401);
or U11530 (N_11530,N_11437,N_11480);
nor U11531 (N_11531,N_11407,N_11494);
or U11532 (N_11532,N_11393,N_11452);
and U11533 (N_11533,N_11433,N_11402);
xnor U11534 (N_11534,N_11465,N_11397);
nor U11535 (N_11535,N_11391,N_11476);
nor U11536 (N_11536,N_11442,N_11487);
nand U11537 (N_11537,N_11415,N_11438);
and U11538 (N_11538,N_11462,N_11420);
and U11539 (N_11539,N_11493,N_11444);
or U11540 (N_11540,N_11464,N_11485);
xnor U11541 (N_11541,N_11445,N_11386);
xor U11542 (N_11542,N_11489,N_11458);
or U11543 (N_11543,N_11388,N_11491);
nand U11544 (N_11544,N_11454,N_11482);
or U11545 (N_11545,N_11412,N_11424);
or U11546 (N_11546,N_11405,N_11472);
xor U11547 (N_11547,N_11463,N_11394);
nand U11548 (N_11548,N_11408,N_11448);
nand U11549 (N_11549,N_11474,N_11441);
nand U11550 (N_11550,N_11384,N_11439);
and U11551 (N_11551,N_11426,N_11430);
nand U11552 (N_11552,N_11429,N_11467);
or U11553 (N_11553,N_11447,N_11403);
nand U11554 (N_11554,N_11385,N_11389);
xor U11555 (N_11555,N_11376,N_11399);
or U11556 (N_11556,N_11434,N_11473);
and U11557 (N_11557,N_11432,N_11436);
nor U11558 (N_11558,N_11470,N_11375);
or U11559 (N_11559,N_11378,N_11380);
nor U11560 (N_11560,N_11400,N_11457);
nor U11561 (N_11561,N_11398,N_11466);
and U11562 (N_11562,N_11390,N_11419);
nor U11563 (N_11563,N_11430,N_11494);
and U11564 (N_11564,N_11452,N_11499);
nor U11565 (N_11565,N_11389,N_11432);
and U11566 (N_11566,N_11415,N_11384);
or U11567 (N_11567,N_11486,N_11467);
nand U11568 (N_11568,N_11385,N_11416);
or U11569 (N_11569,N_11460,N_11386);
xnor U11570 (N_11570,N_11467,N_11379);
and U11571 (N_11571,N_11425,N_11420);
or U11572 (N_11572,N_11420,N_11466);
nor U11573 (N_11573,N_11398,N_11499);
nand U11574 (N_11574,N_11405,N_11499);
nor U11575 (N_11575,N_11483,N_11441);
nor U11576 (N_11576,N_11488,N_11456);
and U11577 (N_11577,N_11437,N_11396);
xnor U11578 (N_11578,N_11497,N_11474);
nor U11579 (N_11579,N_11455,N_11424);
nand U11580 (N_11580,N_11469,N_11462);
nand U11581 (N_11581,N_11387,N_11398);
nand U11582 (N_11582,N_11491,N_11401);
and U11583 (N_11583,N_11497,N_11441);
xnor U11584 (N_11584,N_11385,N_11409);
and U11585 (N_11585,N_11490,N_11445);
nor U11586 (N_11586,N_11485,N_11412);
or U11587 (N_11587,N_11415,N_11469);
or U11588 (N_11588,N_11475,N_11495);
xor U11589 (N_11589,N_11437,N_11401);
xor U11590 (N_11590,N_11430,N_11402);
and U11591 (N_11591,N_11422,N_11472);
xnor U11592 (N_11592,N_11480,N_11389);
or U11593 (N_11593,N_11493,N_11429);
or U11594 (N_11594,N_11456,N_11429);
nand U11595 (N_11595,N_11418,N_11436);
or U11596 (N_11596,N_11439,N_11452);
xnor U11597 (N_11597,N_11404,N_11496);
and U11598 (N_11598,N_11463,N_11473);
xnor U11599 (N_11599,N_11417,N_11391);
and U11600 (N_11600,N_11405,N_11404);
xnor U11601 (N_11601,N_11427,N_11482);
xnor U11602 (N_11602,N_11471,N_11428);
and U11603 (N_11603,N_11451,N_11432);
nor U11604 (N_11604,N_11466,N_11465);
xnor U11605 (N_11605,N_11422,N_11439);
xnor U11606 (N_11606,N_11399,N_11444);
or U11607 (N_11607,N_11429,N_11397);
nand U11608 (N_11608,N_11469,N_11471);
xor U11609 (N_11609,N_11458,N_11421);
xor U11610 (N_11610,N_11455,N_11443);
and U11611 (N_11611,N_11460,N_11409);
and U11612 (N_11612,N_11478,N_11420);
xnor U11613 (N_11613,N_11389,N_11471);
and U11614 (N_11614,N_11386,N_11381);
nor U11615 (N_11615,N_11462,N_11486);
or U11616 (N_11616,N_11479,N_11430);
nand U11617 (N_11617,N_11474,N_11465);
nand U11618 (N_11618,N_11420,N_11429);
or U11619 (N_11619,N_11497,N_11486);
nand U11620 (N_11620,N_11468,N_11477);
nand U11621 (N_11621,N_11395,N_11435);
xor U11622 (N_11622,N_11460,N_11462);
nor U11623 (N_11623,N_11497,N_11391);
xor U11624 (N_11624,N_11376,N_11395);
xnor U11625 (N_11625,N_11621,N_11619);
nor U11626 (N_11626,N_11540,N_11557);
nor U11627 (N_11627,N_11567,N_11580);
or U11628 (N_11628,N_11556,N_11591);
xor U11629 (N_11629,N_11585,N_11510);
or U11630 (N_11630,N_11520,N_11608);
or U11631 (N_11631,N_11562,N_11614);
or U11632 (N_11632,N_11541,N_11530);
xnor U11633 (N_11633,N_11572,N_11565);
nand U11634 (N_11634,N_11561,N_11583);
xnor U11635 (N_11635,N_11515,N_11535);
or U11636 (N_11636,N_11620,N_11555);
xor U11637 (N_11637,N_11613,N_11563);
and U11638 (N_11638,N_11597,N_11551);
xnor U11639 (N_11639,N_11539,N_11624);
nand U11640 (N_11640,N_11616,N_11516);
nor U11641 (N_11641,N_11564,N_11586);
or U11642 (N_11642,N_11596,N_11553);
and U11643 (N_11643,N_11582,N_11511);
and U11644 (N_11644,N_11545,N_11595);
xnor U11645 (N_11645,N_11513,N_11606);
or U11646 (N_11646,N_11618,N_11592);
xor U11647 (N_11647,N_11594,N_11612);
nand U11648 (N_11648,N_11604,N_11528);
xor U11649 (N_11649,N_11501,N_11536);
xnor U11650 (N_11650,N_11527,N_11506);
and U11651 (N_11651,N_11525,N_11599);
and U11652 (N_11652,N_11610,N_11503);
xnor U11653 (N_11653,N_11500,N_11578);
and U11654 (N_11654,N_11532,N_11601);
nand U11655 (N_11655,N_11609,N_11543);
or U11656 (N_11656,N_11598,N_11508);
or U11657 (N_11657,N_11622,N_11569);
nand U11658 (N_11658,N_11589,N_11603);
nor U11659 (N_11659,N_11537,N_11544);
xnor U11660 (N_11660,N_11579,N_11573);
nand U11661 (N_11661,N_11611,N_11552);
nor U11662 (N_11662,N_11605,N_11574);
nand U11663 (N_11663,N_11542,N_11623);
nand U11664 (N_11664,N_11559,N_11521);
nor U11665 (N_11665,N_11607,N_11547);
xor U11666 (N_11666,N_11522,N_11554);
nand U11667 (N_11667,N_11517,N_11588);
and U11668 (N_11668,N_11507,N_11526);
or U11669 (N_11669,N_11584,N_11549);
and U11670 (N_11670,N_11581,N_11519);
and U11671 (N_11671,N_11576,N_11512);
nand U11672 (N_11672,N_11514,N_11502);
xnor U11673 (N_11673,N_11602,N_11593);
or U11674 (N_11674,N_11575,N_11550);
xnor U11675 (N_11675,N_11615,N_11523);
nand U11676 (N_11676,N_11577,N_11509);
and U11677 (N_11677,N_11504,N_11617);
nor U11678 (N_11678,N_11558,N_11587);
nor U11679 (N_11679,N_11571,N_11560);
or U11680 (N_11680,N_11568,N_11546);
nor U11681 (N_11681,N_11590,N_11524);
xor U11682 (N_11682,N_11529,N_11548);
and U11683 (N_11683,N_11566,N_11518);
nor U11684 (N_11684,N_11531,N_11533);
and U11685 (N_11685,N_11534,N_11538);
nand U11686 (N_11686,N_11505,N_11570);
nor U11687 (N_11687,N_11600,N_11567);
nand U11688 (N_11688,N_11522,N_11503);
nor U11689 (N_11689,N_11615,N_11514);
nand U11690 (N_11690,N_11570,N_11566);
nor U11691 (N_11691,N_11583,N_11533);
or U11692 (N_11692,N_11532,N_11562);
nor U11693 (N_11693,N_11610,N_11502);
xor U11694 (N_11694,N_11524,N_11548);
and U11695 (N_11695,N_11580,N_11559);
or U11696 (N_11696,N_11574,N_11505);
nand U11697 (N_11697,N_11624,N_11557);
and U11698 (N_11698,N_11616,N_11555);
or U11699 (N_11699,N_11608,N_11592);
nor U11700 (N_11700,N_11559,N_11508);
nand U11701 (N_11701,N_11518,N_11603);
nor U11702 (N_11702,N_11586,N_11531);
nand U11703 (N_11703,N_11621,N_11572);
nand U11704 (N_11704,N_11527,N_11617);
or U11705 (N_11705,N_11609,N_11603);
xor U11706 (N_11706,N_11507,N_11505);
nor U11707 (N_11707,N_11510,N_11598);
nand U11708 (N_11708,N_11513,N_11622);
xnor U11709 (N_11709,N_11597,N_11580);
nand U11710 (N_11710,N_11571,N_11588);
nor U11711 (N_11711,N_11600,N_11561);
nand U11712 (N_11712,N_11534,N_11610);
nor U11713 (N_11713,N_11546,N_11620);
nor U11714 (N_11714,N_11529,N_11556);
xnor U11715 (N_11715,N_11509,N_11522);
nor U11716 (N_11716,N_11563,N_11597);
or U11717 (N_11717,N_11596,N_11607);
nand U11718 (N_11718,N_11588,N_11581);
and U11719 (N_11719,N_11613,N_11513);
xnor U11720 (N_11720,N_11508,N_11576);
nand U11721 (N_11721,N_11520,N_11624);
nand U11722 (N_11722,N_11520,N_11566);
nand U11723 (N_11723,N_11525,N_11518);
nor U11724 (N_11724,N_11526,N_11548);
xnor U11725 (N_11725,N_11564,N_11594);
and U11726 (N_11726,N_11506,N_11542);
and U11727 (N_11727,N_11595,N_11572);
or U11728 (N_11728,N_11537,N_11605);
xnor U11729 (N_11729,N_11615,N_11534);
nor U11730 (N_11730,N_11574,N_11547);
and U11731 (N_11731,N_11546,N_11598);
nand U11732 (N_11732,N_11531,N_11577);
or U11733 (N_11733,N_11570,N_11539);
or U11734 (N_11734,N_11585,N_11584);
xor U11735 (N_11735,N_11520,N_11564);
xnor U11736 (N_11736,N_11552,N_11620);
or U11737 (N_11737,N_11541,N_11519);
or U11738 (N_11738,N_11559,N_11527);
and U11739 (N_11739,N_11501,N_11603);
xor U11740 (N_11740,N_11616,N_11603);
nand U11741 (N_11741,N_11609,N_11559);
and U11742 (N_11742,N_11616,N_11566);
or U11743 (N_11743,N_11586,N_11566);
and U11744 (N_11744,N_11507,N_11503);
nor U11745 (N_11745,N_11551,N_11581);
or U11746 (N_11746,N_11597,N_11603);
or U11747 (N_11747,N_11570,N_11606);
and U11748 (N_11748,N_11584,N_11597);
nor U11749 (N_11749,N_11561,N_11516);
nand U11750 (N_11750,N_11731,N_11677);
or U11751 (N_11751,N_11660,N_11658);
nand U11752 (N_11752,N_11635,N_11662);
and U11753 (N_11753,N_11730,N_11683);
nor U11754 (N_11754,N_11630,N_11627);
and U11755 (N_11755,N_11723,N_11734);
and U11756 (N_11756,N_11652,N_11742);
nand U11757 (N_11757,N_11674,N_11636);
or U11758 (N_11758,N_11712,N_11640);
and U11759 (N_11759,N_11699,N_11705);
and U11760 (N_11760,N_11643,N_11680);
or U11761 (N_11761,N_11682,N_11721);
and U11762 (N_11762,N_11725,N_11696);
nor U11763 (N_11763,N_11719,N_11664);
and U11764 (N_11764,N_11633,N_11675);
or U11765 (N_11765,N_11678,N_11737);
xor U11766 (N_11766,N_11746,N_11728);
and U11767 (N_11767,N_11628,N_11727);
and U11768 (N_11768,N_11676,N_11685);
or U11769 (N_11769,N_11668,N_11669);
nand U11770 (N_11770,N_11661,N_11641);
nor U11771 (N_11771,N_11702,N_11659);
and U11772 (N_11772,N_11629,N_11681);
or U11773 (N_11773,N_11644,N_11694);
and U11774 (N_11774,N_11703,N_11647);
and U11775 (N_11775,N_11706,N_11645);
nand U11776 (N_11776,N_11743,N_11722);
and U11777 (N_11777,N_11736,N_11749);
nor U11778 (N_11778,N_11666,N_11655);
nand U11779 (N_11779,N_11716,N_11740);
nor U11780 (N_11780,N_11670,N_11687);
or U11781 (N_11781,N_11626,N_11708);
nor U11782 (N_11782,N_11657,N_11711);
or U11783 (N_11783,N_11689,N_11744);
nor U11784 (N_11784,N_11729,N_11654);
nor U11785 (N_11785,N_11724,N_11646);
nor U11786 (N_11786,N_11748,N_11671);
xnor U11787 (N_11787,N_11733,N_11710);
nor U11788 (N_11788,N_11747,N_11638);
nand U11789 (N_11789,N_11713,N_11632);
and U11790 (N_11790,N_11648,N_11714);
nand U11791 (N_11791,N_11693,N_11686);
or U11792 (N_11792,N_11738,N_11720);
or U11793 (N_11793,N_11665,N_11717);
nor U11794 (N_11794,N_11715,N_11697);
or U11795 (N_11795,N_11739,N_11698);
nand U11796 (N_11796,N_11663,N_11634);
xor U11797 (N_11797,N_11679,N_11735);
xnor U11798 (N_11798,N_11631,N_11691);
xor U11799 (N_11799,N_11745,N_11692);
nand U11800 (N_11800,N_11700,N_11667);
nand U11801 (N_11801,N_11704,N_11701);
nor U11802 (N_11802,N_11649,N_11690);
xnor U11803 (N_11803,N_11709,N_11718);
and U11804 (N_11804,N_11732,N_11639);
and U11805 (N_11805,N_11642,N_11688);
nand U11806 (N_11806,N_11650,N_11625);
nand U11807 (N_11807,N_11707,N_11637);
xor U11808 (N_11808,N_11656,N_11651);
xor U11809 (N_11809,N_11672,N_11741);
xor U11810 (N_11810,N_11653,N_11684);
xor U11811 (N_11811,N_11695,N_11673);
nand U11812 (N_11812,N_11726,N_11709);
and U11813 (N_11813,N_11695,N_11682);
nand U11814 (N_11814,N_11685,N_11663);
nor U11815 (N_11815,N_11688,N_11715);
or U11816 (N_11816,N_11628,N_11679);
or U11817 (N_11817,N_11664,N_11731);
xnor U11818 (N_11818,N_11635,N_11668);
nor U11819 (N_11819,N_11664,N_11699);
nand U11820 (N_11820,N_11671,N_11678);
nand U11821 (N_11821,N_11717,N_11746);
xnor U11822 (N_11822,N_11725,N_11633);
nand U11823 (N_11823,N_11648,N_11703);
xnor U11824 (N_11824,N_11674,N_11661);
nand U11825 (N_11825,N_11668,N_11702);
xor U11826 (N_11826,N_11650,N_11747);
nor U11827 (N_11827,N_11698,N_11747);
or U11828 (N_11828,N_11664,N_11633);
and U11829 (N_11829,N_11709,N_11749);
nor U11830 (N_11830,N_11727,N_11728);
nand U11831 (N_11831,N_11715,N_11628);
nand U11832 (N_11832,N_11657,N_11675);
nand U11833 (N_11833,N_11745,N_11739);
xnor U11834 (N_11834,N_11662,N_11730);
nand U11835 (N_11835,N_11727,N_11643);
and U11836 (N_11836,N_11729,N_11671);
and U11837 (N_11837,N_11707,N_11632);
nand U11838 (N_11838,N_11705,N_11663);
nor U11839 (N_11839,N_11649,N_11721);
and U11840 (N_11840,N_11641,N_11695);
nand U11841 (N_11841,N_11712,N_11660);
nand U11842 (N_11842,N_11727,N_11748);
nand U11843 (N_11843,N_11653,N_11686);
nor U11844 (N_11844,N_11741,N_11737);
nor U11845 (N_11845,N_11627,N_11696);
or U11846 (N_11846,N_11704,N_11694);
or U11847 (N_11847,N_11652,N_11712);
or U11848 (N_11848,N_11658,N_11693);
xnor U11849 (N_11849,N_11720,N_11682);
xnor U11850 (N_11850,N_11720,N_11665);
nor U11851 (N_11851,N_11658,N_11682);
xor U11852 (N_11852,N_11655,N_11673);
or U11853 (N_11853,N_11636,N_11628);
nor U11854 (N_11854,N_11744,N_11682);
nor U11855 (N_11855,N_11661,N_11630);
and U11856 (N_11856,N_11695,N_11739);
xnor U11857 (N_11857,N_11680,N_11722);
nand U11858 (N_11858,N_11703,N_11747);
nor U11859 (N_11859,N_11725,N_11729);
nor U11860 (N_11860,N_11687,N_11664);
xnor U11861 (N_11861,N_11701,N_11640);
nand U11862 (N_11862,N_11721,N_11742);
and U11863 (N_11863,N_11744,N_11721);
xor U11864 (N_11864,N_11724,N_11642);
or U11865 (N_11865,N_11697,N_11727);
nor U11866 (N_11866,N_11721,N_11741);
or U11867 (N_11867,N_11696,N_11670);
and U11868 (N_11868,N_11747,N_11636);
and U11869 (N_11869,N_11732,N_11694);
nor U11870 (N_11870,N_11659,N_11719);
and U11871 (N_11871,N_11696,N_11743);
or U11872 (N_11872,N_11687,N_11697);
nor U11873 (N_11873,N_11703,N_11717);
nand U11874 (N_11874,N_11694,N_11734);
nand U11875 (N_11875,N_11866,N_11831);
nand U11876 (N_11876,N_11856,N_11836);
nor U11877 (N_11877,N_11859,N_11796);
nor U11878 (N_11878,N_11754,N_11782);
xnor U11879 (N_11879,N_11751,N_11784);
xnor U11880 (N_11880,N_11765,N_11766);
xnor U11881 (N_11881,N_11826,N_11872);
and U11882 (N_11882,N_11799,N_11750);
and U11883 (N_11883,N_11824,N_11862);
or U11884 (N_11884,N_11756,N_11844);
or U11885 (N_11885,N_11760,N_11833);
nor U11886 (N_11886,N_11803,N_11812);
or U11887 (N_11887,N_11864,N_11809);
nand U11888 (N_11888,N_11768,N_11755);
nor U11889 (N_11889,N_11835,N_11753);
or U11890 (N_11890,N_11790,N_11817);
nand U11891 (N_11891,N_11811,N_11802);
and U11892 (N_11892,N_11763,N_11752);
or U11893 (N_11893,N_11792,N_11814);
nor U11894 (N_11894,N_11853,N_11810);
nor U11895 (N_11895,N_11818,N_11785);
nor U11896 (N_11896,N_11845,N_11771);
nor U11897 (N_11897,N_11804,N_11834);
nand U11898 (N_11898,N_11773,N_11794);
xor U11899 (N_11899,N_11851,N_11789);
nand U11900 (N_11900,N_11837,N_11828);
nand U11901 (N_11901,N_11776,N_11863);
xnor U11902 (N_11902,N_11798,N_11758);
xnor U11903 (N_11903,N_11778,N_11767);
xnor U11904 (N_11904,N_11779,N_11858);
or U11905 (N_11905,N_11820,N_11827);
xor U11906 (N_11906,N_11813,N_11840);
or U11907 (N_11907,N_11762,N_11838);
or U11908 (N_11908,N_11781,N_11852);
nor U11909 (N_11909,N_11865,N_11816);
xnor U11910 (N_11910,N_11860,N_11801);
xor U11911 (N_11911,N_11775,N_11842);
and U11912 (N_11912,N_11757,N_11857);
and U11913 (N_11913,N_11806,N_11832);
nand U11914 (N_11914,N_11780,N_11867);
nand U11915 (N_11915,N_11839,N_11871);
or U11916 (N_11916,N_11874,N_11791);
nand U11917 (N_11917,N_11772,N_11759);
or U11918 (N_11918,N_11761,N_11787);
xor U11919 (N_11919,N_11823,N_11870);
or U11920 (N_11920,N_11800,N_11769);
nor U11921 (N_11921,N_11830,N_11770);
nand U11922 (N_11922,N_11795,N_11841);
or U11923 (N_11923,N_11808,N_11821);
nor U11924 (N_11924,N_11849,N_11843);
nor U11925 (N_11925,N_11819,N_11847);
or U11926 (N_11926,N_11869,N_11873);
or U11927 (N_11927,N_11846,N_11783);
xnor U11928 (N_11928,N_11807,N_11786);
nand U11929 (N_11929,N_11764,N_11848);
or U11930 (N_11930,N_11854,N_11855);
nor U11931 (N_11931,N_11825,N_11861);
xor U11932 (N_11932,N_11868,N_11850);
nand U11933 (N_11933,N_11815,N_11805);
or U11934 (N_11934,N_11777,N_11829);
xor U11935 (N_11935,N_11774,N_11822);
nand U11936 (N_11936,N_11788,N_11793);
or U11937 (N_11937,N_11797,N_11773);
nand U11938 (N_11938,N_11789,N_11751);
xor U11939 (N_11939,N_11769,N_11820);
nor U11940 (N_11940,N_11842,N_11793);
or U11941 (N_11941,N_11858,N_11831);
nor U11942 (N_11942,N_11814,N_11848);
or U11943 (N_11943,N_11837,N_11755);
nor U11944 (N_11944,N_11761,N_11789);
nand U11945 (N_11945,N_11843,N_11765);
or U11946 (N_11946,N_11772,N_11818);
and U11947 (N_11947,N_11852,N_11842);
nor U11948 (N_11948,N_11862,N_11774);
xnor U11949 (N_11949,N_11840,N_11805);
and U11950 (N_11950,N_11871,N_11826);
nand U11951 (N_11951,N_11786,N_11799);
nor U11952 (N_11952,N_11806,N_11844);
xnor U11953 (N_11953,N_11864,N_11771);
and U11954 (N_11954,N_11817,N_11792);
nand U11955 (N_11955,N_11834,N_11866);
and U11956 (N_11956,N_11812,N_11835);
or U11957 (N_11957,N_11843,N_11809);
and U11958 (N_11958,N_11792,N_11868);
nor U11959 (N_11959,N_11819,N_11777);
and U11960 (N_11960,N_11803,N_11801);
nand U11961 (N_11961,N_11831,N_11872);
or U11962 (N_11962,N_11857,N_11816);
nor U11963 (N_11963,N_11765,N_11830);
nand U11964 (N_11964,N_11812,N_11822);
or U11965 (N_11965,N_11799,N_11783);
xor U11966 (N_11966,N_11826,N_11766);
xor U11967 (N_11967,N_11843,N_11761);
xor U11968 (N_11968,N_11801,N_11815);
and U11969 (N_11969,N_11785,N_11845);
or U11970 (N_11970,N_11873,N_11865);
or U11971 (N_11971,N_11792,N_11801);
or U11972 (N_11972,N_11821,N_11752);
or U11973 (N_11973,N_11871,N_11852);
nor U11974 (N_11974,N_11831,N_11809);
or U11975 (N_11975,N_11784,N_11839);
or U11976 (N_11976,N_11806,N_11762);
xor U11977 (N_11977,N_11869,N_11862);
nand U11978 (N_11978,N_11795,N_11809);
and U11979 (N_11979,N_11858,N_11846);
nand U11980 (N_11980,N_11833,N_11802);
xor U11981 (N_11981,N_11761,N_11846);
nor U11982 (N_11982,N_11796,N_11845);
and U11983 (N_11983,N_11796,N_11820);
and U11984 (N_11984,N_11795,N_11763);
and U11985 (N_11985,N_11826,N_11854);
and U11986 (N_11986,N_11826,N_11800);
nand U11987 (N_11987,N_11864,N_11800);
nand U11988 (N_11988,N_11807,N_11809);
nor U11989 (N_11989,N_11852,N_11858);
nand U11990 (N_11990,N_11750,N_11847);
nand U11991 (N_11991,N_11786,N_11754);
nand U11992 (N_11992,N_11830,N_11761);
xnor U11993 (N_11993,N_11761,N_11829);
nand U11994 (N_11994,N_11777,N_11769);
nand U11995 (N_11995,N_11849,N_11760);
and U11996 (N_11996,N_11798,N_11840);
and U11997 (N_11997,N_11861,N_11849);
nand U11998 (N_11998,N_11771,N_11848);
xnor U11999 (N_11999,N_11843,N_11866);
xnor U12000 (N_12000,N_11997,N_11875);
nor U12001 (N_12001,N_11935,N_11956);
xor U12002 (N_12002,N_11911,N_11905);
or U12003 (N_12003,N_11890,N_11916);
and U12004 (N_12004,N_11985,N_11925);
nor U12005 (N_12005,N_11970,N_11975);
and U12006 (N_12006,N_11895,N_11965);
nor U12007 (N_12007,N_11938,N_11969);
nor U12008 (N_12008,N_11885,N_11964);
xnor U12009 (N_12009,N_11884,N_11981);
nor U12010 (N_12010,N_11908,N_11949);
or U12011 (N_12011,N_11974,N_11951);
and U12012 (N_12012,N_11966,N_11927);
and U12013 (N_12013,N_11992,N_11896);
xnor U12014 (N_12014,N_11947,N_11990);
nand U12015 (N_12015,N_11957,N_11883);
and U12016 (N_12016,N_11960,N_11919);
xnor U12017 (N_12017,N_11915,N_11941);
nor U12018 (N_12018,N_11978,N_11891);
nand U12019 (N_12019,N_11936,N_11893);
or U12020 (N_12020,N_11886,N_11902);
and U12021 (N_12021,N_11904,N_11879);
or U12022 (N_12022,N_11993,N_11994);
nor U12023 (N_12023,N_11914,N_11898);
nor U12024 (N_12024,N_11900,N_11906);
or U12025 (N_12025,N_11918,N_11972);
and U12026 (N_12026,N_11940,N_11892);
nor U12027 (N_12027,N_11920,N_11922);
nor U12028 (N_12028,N_11948,N_11942);
nor U12029 (N_12029,N_11979,N_11894);
or U12030 (N_12030,N_11931,N_11967);
nand U12031 (N_12031,N_11986,N_11962);
nor U12032 (N_12032,N_11945,N_11977);
nor U12033 (N_12033,N_11880,N_11932);
nand U12034 (N_12034,N_11988,N_11955);
nand U12035 (N_12035,N_11996,N_11943);
nor U12036 (N_12036,N_11921,N_11995);
or U12037 (N_12037,N_11953,N_11881);
or U12038 (N_12038,N_11934,N_11954);
nor U12039 (N_12039,N_11917,N_11878);
nand U12040 (N_12040,N_11933,N_11959);
nand U12041 (N_12041,N_11971,N_11897);
and U12042 (N_12042,N_11998,N_11888);
nand U12043 (N_12043,N_11923,N_11913);
and U12044 (N_12044,N_11929,N_11930);
or U12045 (N_12045,N_11877,N_11889);
and U12046 (N_12046,N_11924,N_11983);
and U12047 (N_12047,N_11991,N_11982);
or U12048 (N_12048,N_11910,N_11989);
nand U12049 (N_12049,N_11976,N_11984);
nor U12050 (N_12050,N_11973,N_11876);
xnor U12051 (N_12051,N_11963,N_11912);
xnor U12052 (N_12052,N_11944,N_11958);
nor U12053 (N_12053,N_11952,N_11907);
and U12054 (N_12054,N_11980,N_11961);
nor U12055 (N_12055,N_11926,N_11968);
and U12056 (N_12056,N_11909,N_11901);
xnor U12057 (N_12057,N_11887,N_11937);
nor U12058 (N_12058,N_11987,N_11899);
nand U12059 (N_12059,N_11903,N_11939);
or U12060 (N_12060,N_11950,N_11999);
nor U12061 (N_12061,N_11882,N_11928);
nor U12062 (N_12062,N_11946,N_11898);
and U12063 (N_12063,N_11952,N_11963);
or U12064 (N_12064,N_11901,N_11937);
or U12065 (N_12065,N_11901,N_11954);
nand U12066 (N_12066,N_11970,N_11954);
xnor U12067 (N_12067,N_11929,N_11935);
nand U12068 (N_12068,N_11950,N_11953);
and U12069 (N_12069,N_11890,N_11987);
nand U12070 (N_12070,N_11986,N_11928);
nand U12071 (N_12071,N_11999,N_11984);
and U12072 (N_12072,N_11965,N_11904);
xnor U12073 (N_12073,N_11922,N_11954);
and U12074 (N_12074,N_11893,N_11981);
nand U12075 (N_12075,N_11970,N_11930);
xnor U12076 (N_12076,N_11995,N_11907);
and U12077 (N_12077,N_11928,N_11941);
nand U12078 (N_12078,N_11982,N_11891);
xor U12079 (N_12079,N_11967,N_11961);
or U12080 (N_12080,N_11970,N_11916);
nand U12081 (N_12081,N_11932,N_11937);
nor U12082 (N_12082,N_11917,N_11945);
or U12083 (N_12083,N_11988,N_11901);
nand U12084 (N_12084,N_11933,N_11971);
xnor U12085 (N_12085,N_11935,N_11902);
and U12086 (N_12086,N_11950,N_11933);
xnor U12087 (N_12087,N_11899,N_11895);
nand U12088 (N_12088,N_11990,N_11902);
and U12089 (N_12089,N_11992,N_11933);
nor U12090 (N_12090,N_11917,N_11944);
nor U12091 (N_12091,N_11969,N_11925);
and U12092 (N_12092,N_11972,N_11878);
or U12093 (N_12093,N_11952,N_11976);
nor U12094 (N_12094,N_11921,N_11892);
xor U12095 (N_12095,N_11980,N_11971);
or U12096 (N_12096,N_11997,N_11876);
and U12097 (N_12097,N_11947,N_11935);
or U12098 (N_12098,N_11925,N_11960);
xor U12099 (N_12099,N_11968,N_11925);
or U12100 (N_12100,N_11966,N_11910);
nor U12101 (N_12101,N_11925,N_11935);
nor U12102 (N_12102,N_11931,N_11927);
nor U12103 (N_12103,N_11938,N_11932);
nand U12104 (N_12104,N_11950,N_11895);
and U12105 (N_12105,N_11887,N_11941);
nor U12106 (N_12106,N_11968,N_11957);
xnor U12107 (N_12107,N_11975,N_11916);
nand U12108 (N_12108,N_11884,N_11928);
nand U12109 (N_12109,N_11995,N_11915);
or U12110 (N_12110,N_11953,N_11935);
nand U12111 (N_12111,N_11972,N_11961);
nor U12112 (N_12112,N_11887,N_11885);
xor U12113 (N_12113,N_11957,N_11967);
and U12114 (N_12114,N_11916,N_11918);
nor U12115 (N_12115,N_11951,N_11947);
nand U12116 (N_12116,N_11930,N_11947);
nor U12117 (N_12117,N_11923,N_11940);
nor U12118 (N_12118,N_11892,N_11875);
xnor U12119 (N_12119,N_11923,N_11971);
xnor U12120 (N_12120,N_11988,N_11994);
xnor U12121 (N_12121,N_11921,N_11944);
xor U12122 (N_12122,N_11967,N_11913);
nand U12123 (N_12123,N_11911,N_11942);
or U12124 (N_12124,N_11956,N_11997);
nor U12125 (N_12125,N_12065,N_12076);
and U12126 (N_12126,N_12011,N_12005);
nor U12127 (N_12127,N_12097,N_12075);
nor U12128 (N_12128,N_12022,N_12112);
nor U12129 (N_12129,N_12120,N_12053);
nand U12130 (N_12130,N_12042,N_12012);
and U12131 (N_12131,N_12092,N_12108);
and U12132 (N_12132,N_12121,N_12028);
nand U12133 (N_12133,N_12032,N_12072);
nor U12134 (N_12134,N_12098,N_12007);
and U12135 (N_12135,N_12000,N_12059);
nor U12136 (N_12136,N_12113,N_12067);
and U12137 (N_12137,N_12013,N_12055);
nand U12138 (N_12138,N_12044,N_12054);
nor U12139 (N_12139,N_12045,N_12002);
nor U12140 (N_12140,N_12026,N_12100);
nor U12141 (N_12141,N_12020,N_12001);
nand U12142 (N_12142,N_12089,N_12094);
and U12143 (N_12143,N_12118,N_12062);
nand U12144 (N_12144,N_12095,N_12087);
or U12145 (N_12145,N_12102,N_12106);
nand U12146 (N_12146,N_12099,N_12082);
and U12147 (N_12147,N_12030,N_12039);
xnor U12148 (N_12148,N_12037,N_12058);
or U12149 (N_12149,N_12085,N_12096);
nand U12150 (N_12150,N_12014,N_12016);
or U12151 (N_12151,N_12071,N_12025);
or U12152 (N_12152,N_12086,N_12029);
and U12153 (N_12153,N_12035,N_12043);
nand U12154 (N_12154,N_12056,N_12079);
and U12155 (N_12155,N_12049,N_12077);
xor U12156 (N_12156,N_12115,N_12040);
nor U12157 (N_12157,N_12051,N_12060);
xor U12158 (N_12158,N_12111,N_12006);
xnor U12159 (N_12159,N_12122,N_12124);
nor U12160 (N_12160,N_12080,N_12031);
or U12161 (N_12161,N_12047,N_12010);
nand U12162 (N_12162,N_12063,N_12048);
nor U12163 (N_12163,N_12078,N_12069);
xor U12164 (N_12164,N_12041,N_12009);
nand U12165 (N_12165,N_12114,N_12105);
nand U12166 (N_12166,N_12081,N_12117);
nand U12167 (N_12167,N_12066,N_12064);
nand U12168 (N_12168,N_12091,N_12083);
xor U12169 (N_12169,N_12110,N_12034);
nand U12170 (N_12170,N_12119,N_12090);
xor U12171 (N_12171,N_12004,N_12123);
nand U12172 (N_12172,N_12103,N_12107);
or U12173 (N_12173,N_12050,N_12068);
xor U12174 (N_12174,N_12038,N_12104);
nand U12175 (N_12175,N_12070,N_12023);
xor U12176 (N_12176,N_12057,N_12088);
and U12177 (N_12177,N_12046,N_12074);
and U12178 (N_12178,N_12109,N_12061);
nand U12179 (N_12179,N_12093,N_12015);
or U12180 (N_12180,N_12017,N_12052);
xnor U12181 (N_12181,N_12084,N_12024);
xnor U12182 (N_12182,N_12116,N_12019);
xnor U12183 (N_12183,N_12021,N_12008);
nor U12184 (N_12184,N_12003,N_12027);
xor U12185 (N_12185,N_12073,N_12018);
nand U12186 (N_12186,N_12036,N_12033);
nand U12187 (N_12187,N_12101,N_12070);
nand U12188 (N_12188,N_12050,N_12044);
and U12189 (N_12189,N_12120,N_12081);
nor U12190 (N_12190,N_12115,N_12013);
nand U12191 (N_12191,N_12030,N_12070);
or U12192 (N_12192,N_12102,N_12094);
nor U12193 (N_12193,N_12024,N_12124);
nor U12194 (N_12194,N_12114,N_12027);
xor U12195 (N_12195,N_12117,N_12027);
nand U12196 (N_12196,N_12062,N_12092);
xor U12197 (N_12197,N_12024,N_12062);
nand U12198 (N_12198,N_12121,N_12058);
nor U12199 (N_12199,N_12101,N_12081);
nand U12200 (N_12200,N_12018,N_12037);
nor U12201 (N_12201,N_12103,N_12124);
nand U12202 (N_12202,N_12074,N_12081);
nor U12203 (N_12203,N_12081,N_12100);
nand U12204 (N_12204,N_12049,N_12105);
xor U12205 (N_12205,N_12013,N_12095);
nor U12206 (N_12206,N_12034,N_12071);
nor U12207 (N_12207,N_12076,N_12006);
and U12208 (N_12208,N_12113,N_12018);
and U12209 (N_12209,N_12005,N_12081);
or U12210 (N_12210,N_12059,N_12054);
nor U12211 (N_12211,N_12076,N_12068);
nand U12212 (N_12212,N_12095,N_12045);
and U12213 (N_12213,N_12115,N_12046);
or U12214 (N_12214,N_12042,N_12076);
or U12215 (N_12215,N_12036,N_12025);
and U12216 (N_12216,N_12023,N_12007);
xnor U12217 (N_12217,N_12016,N_12100);
nand U12218 (N_12218,N_12016,N_12086);
and U12219 (N_12219,N_12101,N_12098);
xor U12220 (N_12220,N_12111,N_12093);
nand U12221 (N_12221,N_12074,N_12097);
and U12222 (N_12222,N_12017,N_12065);
or U12223 (N_12223,N_12104,N_12116);
nand U12224 (N_12224,N_12043,N_12016);
and U12225 (N_12225,N_12097,N_12106);
and U12226 (N_12226,N_12046,N_12099);
and U12227 (N_12227,N_12001,N_12026);
nand U12228 (N_12228,N_12020,N_12011);
or U12229 (N_12229,N_12077,N_12044);
and U12230 (N_12230,N_12091,N_12060);
or U12231 (N_12231,N_12011,N_12112);
xnor U12232 (N_12232,N_12000,N_12102);
xnor U12233 (N_12233,N_12043,N_12081);
xnor U12234 (N_12234,N_12026,N_12090);
nor U12235 (N_12235,N_12055,N_12032);
or U12236 (N_12236,N_12091,N_12113);
xor U12237 (N_12237,N_12089,N_12085);
xnor U12238 (N_12238,N_12107,N_12072);
xor U12239 (N_12239,N_12090,N_12118);
nand U12240 (N_12240,N_12086,N_12036);
or U12241 (N_12241,N_12023,N_12065);
xnor U12242 (N_12242,N_12074,N_12079);
and U12243 (N_12243,N_12019,N_12099);
nand U12244 (N_12244,N_12079,N_12060);
or U12245 (N_12245,N_12079,N_12033);
and U12246 (N_12246,N_12071,N_12115);
nor U12247 (N_12247,N_12013,N_12027);
nand U12248 (N_12248,N_12109,N_12033);
nor U12249 (N_12249,N_12060,N_12047);
xnor U12250 (N_12250,N_12143,N_12205);
xor U12251 (N_12251,N_12220,N_12188);
and U12252 (N_12252,N_12181,N_12179);
nor U12253 (N_12253,N_12195,N_12231);
and U12254 (N_12254,N_12154,N_12168);
nor U12255 (N_12255,N_12129,N_12238);
nand U12256 (N_12256,N_12130,N_12157);
and U12257 (N_12257,N_12128,N_12127);
or U12258 (N_12258,N_12236,N_12156);
and U12259 (N_12259,N_12159,N_12165);
xnor U12260 (N_12260,N_12227,N_12237);
nor U12261 (N_12261,N_12246,N_12166);
nand U12262 (N_12262,N_12164,N_12225);
xor U12263 (N_12263,N_12241,N_12162);
or U12264 (N_12264,N_12173,N_12219);
xor U12265 (N_12265,N_12229,N_12247);
xnor U12266 (N_12266,N_12136,N_12183);
or U12267 (N_12267,N_12145,N_12134);
or U12268 (N_12268,N_12208,N_12224);
or U12269 (N_12269,N_12178,N_12153);
nand U12270 (N_12270,N_12193,N_12199);
nand U12271 (N_12271,N_12203,N_12170);
and U12272 (N_12272,N_12244,N_12222);
xnor U12273 (N_12273,N_12243,N_12135);
xnor U12274 (N_12274,N_12189,N_12240);
and U12275 (N_12275,N_12215,N_12198);
and U12276 (N_12276,N_12239,N_12191);
xnor U12277 (N_12277,N_12138,N_12144);
nand U12278 (N_12278,N_12126,N_12147);
nand U12279 (N_12279,N_12155,N_12211);
nor U12280 (N_12280,N_12207,N_12148);
nor U12281 (N_12281,N_12194,N_12230);
nand U12282 (N_12282,N_12206,N_12172);
nand U12283 (N_12283,N_12160,N_12146);
and U12284 (N_12284,N_12152,N_12151);
and U12285 (N_12285,N_12218,N_12187);
nand U12286 (N_12286,N_12158,N_12192);
xnor U12287 (N_12287,N_12248,N_12137);
nor U12288 (N_12288,N_12201,N_12167);
and U12289 (N_12289,N_12200,N_12142);
or U12290 (N_12290,N_12226,N_12235);
xor U12291 (N_12291,N_12174,N_12185);
nand U12292 (N_12292,N_12161,N_12223);
nand U12293 (N_12293,N_12182,N_12249);
xor U12294 (N_12294,N_12175,N_12197);
xor U12295 (N_12295,N_12133,N_12214);
nand U12296 (N_12296,N_12196,N_12210);
and U12297 (N_12297,N_12149,N_12190);
xnor U12298 (N_12298,N_12209,N_12184);
xnor U12299 (N_12299,N_12132,N_12202);
nor U12300 (N_12300,N_12169,N_12131);
xor U12301 (N_12301,N_12150,N_12212);
xnor U12302 (N_12302,N_12221,N_12216);
xor U12303 (N_12303,N_12125,N_12141);
nor U12304 (N_12304,N_12139,N_12140);
or U12305 (N_12305,N_12163,N_12176);
and U12306 (N_12306,N_12228,N_12171);
nor U12307 (N_12307,N_12217,N_12242);
or U12308 (N_12308,N_12233,N_12180);
xor U12309 (N_12309,N_12213,N_12232);
nor U12310 (N_12310,N_12186,N_12234);
nor U12311 (N_12311,N_12245,N_12177);
or U12312 (N_12312,N_12204,N_12138);
xor U12313 (N_12313,N_12182,N_12172);
xnor U12314 (N_12314,N_12149,N_12204);
nor U12315 (N_12315,N_12190,N_12228);
nand U12316 (N_12316,N_12163,N_12194);
nor U12317 (N_12317,N_12137,N_12136);
nand U12318 (N_12318,N_12179,N_12215);
nor U12319 (N_12319,N_12228,N_12131);
and U12320 (N_12320,N_12162,N_12168);
xnor U12321 (N_12321,N_12166,N_12224);
xnor U12322 (N_12322,N_12183,N_12190);
xor U12323 (N_12323,N_12238,N_12234);
and U12324 (N_12324,N_12132,N_12164);
nor U12325 (N_12325,N_12141,N_12144);
nor U12326 (N_12326,N_12182,N_12229);
xor U12327 (N_12327,N_12161,N_12191);
xor U12328 (N_12328,N_12201,N_12166);
nor U12329 (N_12329,N_12213,N_12165);
and U12330 (N_12330,N_12185,N_12139);
nor U12331 (N_12331,N_12169,N_12160);
and U12332 (N_12332,N_12146,N_12180);
nand U12333 (N_12333,N_12248,N_12184);
and U12334 (N_12334,N_12209,N_12234);
and U12335 (N_12335,N_12231,N_12142);
and U12336 (N_12336,N_12246,N_12234);
nand U12337 (N_12337,N_12185,N_12191);
xor U12338 (N_12338,N_12206,N_12152);
and U12339 (N_12339,N_12197,N_12129);
or U12340 (N_12340,N_12154,N_12149);
or U12341 (N_12341,N_12194,N_12211);
and U12342 (N_12342,N_12126,N_12162);
nand U12343 (N_12343,N_12220,N_12234);
xor U12344 (N_12344,N_12233,N_12158);
and U12345 (N_12345,N_12245,N_12192);
and U12346 (N_12346,N_12194,N_12135);
or U12347 (N_12347,N_12169,N_12164);
nand U12348 (N_12348,N_12244,N_12199);
or U12349 (N_12349,N_12242,N_12221);
or U12350 (N_12350,N_12187,N_12232);
and U12351 (N_12351,N_12140,N_12131);
xnor U12352 (N_12352,N_12223,N_12166);
nor U12353 (N_12353,N_12181,N_12172);
and U12354 (N_12354,N_12237,N_12142);
nand U12355 (N_12355,N_12243,N_12147);
xnor U12356 (N_12356,N_12241,N_12150);
nand U12357 (N_12357,N_12135,N_12187);
nand U12358 (N_12358,N_12245,N_12230);
or U12359 (N_12359,N_12213,N_12160);
and U12360 (N_12360,N_12190,N_12153);
or U12361 (N_12361,N_12136,N_12176);
xnor U12362 (N_12362,N_12136,N_12146);
nor U12363 (N_12363,N_12172,N_12235);
xnor U12364 (N_12364,N_12225,N_12179);
nor U12365 (N_12365,N_12214,N_12128);
xnor U12366 (N_12366,N_12146,N_12127);
nand U12367 (N_12367,N_12226,N_12133);
xor U12368 (N_12368,N_12216,N_12170);
nor U12369 (N_12369,N_12170,N_12134);
or U12370 (N_12370,N_12154,N_12178);
nor U12371 (N_12371,N_12153,N_12221);
nor U12372 (N_12372,N_12222,N_12194);
nand U12373 (N_12373,N_12236,N_12244);
nor U12374 (N_12374,N_12206,N_12220);
and U12375 (N_12375,N_12260,N_12354);
nand U12376 (N_12376,N_12346,N_12353);
xor U12377 (N_12377,N_12258,N_12361);
and U12378 (N_12378,N_12293,N_12302);
nand U12379 (N_12379,N_12298,N_12290);
and U12380 (N_12380,N_12333,N_12283);
or U12381 (N_12381,N_12308,N_12277);
nand U12382 (N_12382,N_12292,N_12296);
nand U12383 (N_12383,N_12366,N_12307);
and U12384 (N_12384,N_12356,N_12287);
or U12385 (N_12385,N_12310,N_12278);
xor U12386 (N_12386,N_12259,N_12320);
nand U12387 (N_12387,N_12364,N_12316);
nand U12388 (N_12388,N_12312,N_12301);
xor U12389 (N_12389,N_12317,N_12358);
and U12390 (N_12390,N_12299,N_12251);
nand U12391 (N_12391,N_12348,N_12282);
nor U12392 (N_12392,N_12315,N_12355);
and U12393 (N_12393,N_12265,N_12264);
nand U12394 (N_12394,N_12340,N_12322);
nand U12395 (N_12395,N_12373,N_12369);
nand U12396 (N_12396,N_12344,N_12327);
nand U12397 (N_12397,N_12274,N_12347);
or U12398 (N_12398,N_12365,N_12332);
and U12399 (N_12399,N_12257,N_12367);
nor U12400 (N_12400,N_12319,N_12313);
nor U12401 (N_12401,N_12279,N_12271);
nor U12402 (N_12402,N_12374,N_12255);
xnor U12403 (N_12403,N_12281,N_12276);
or U12404 (N_12404,N_12280,N_12331);
or U12405 (N_12405,N_12330,N_12306);
or U12406 (N_12406,N_12342,N_12311);
nand U12407 (N_12407,N_12334,N_12250);
nand U12408 (N_12408,N_12272,N_12341);
nand U12409 (N_12409,N_12323,N_12352);
nor U12410 (N_12410,N_12305,N_12350);
nor U12411 (N_12411,N_12338,N_12309);
xor U12412 (N_12412,N_12351,N_12289);
or U12413 (N_12413,N_12253,N_12371);
xor U12414 (N_12414,N_12314,N_12303);
and U12415 (N_12415,N_12261,N_12268);
xnor U12416 (N_12416,N_12262,N_12325);
xor U12417 (N_12417,N_12273,N_12357);
and U12418 (N_12418,N_12337,N_12329);
or U12419 (N_12419,N_12339,N_12295);
nor U12420 (N_12420,N_12336,N_12345);
nor U12421 (N_12421,N_12363,N_12266);
nand U12422 (N_12422,N_12288,N_12324);
and U12423 (N_12423,N_12267,N_12318);
nor U12424 (N_12424,N_12291,N_12269);
or U12425 (N_12425,N_12300,N_12362);
or U12426 (N_12426,N_12349,N_12359);
xor U12427 (N_12427,N_12263,N_12370);
xnor U12428 (N_12428,N_12297,N_12335);
nor U12429 (N_12429,N_12304,N_12368);
and U12430 (N_12430,N_12286,N_12328);
nor U12431 (N_12431,N_12254,N_12275);
xnor U12432 (N_12432,N_12360,N_12294);
xor U12433 (N_12433,N_12285,N_12270);
or U12434 (N_12434,N_12256,N_12321);
nand U12435 (N_12435,N_12326,N_12284);
nor U12436 (N_12436,N_12372,N_12343);
and U12437 (N_12437,N_12252,N_12368);
nand U12438 (N_12438,N_12371,N_12281);
nand U12439 (N_12439,N_12344,N_12333);
xnor U12440 (N_12440,N_12341,N_12372);
xnor U12441 (N_12441,N_12372,N_12337);
xnor U12442 (N_12442,N_12270,N_12363);
xnor U12443 (N_12443,N_12259,N_12315);
nor U12444 (N_12444,N_12357,N_12347);
and U12445 (N_12445,N_12335,N_12251);
nand U12446 (N_12446,N_12341,N_12321);
or U12447 (N_12447,N_12302,N_12351);
or U12448 (N_12448,N_12298,N_12308);
nor U12449 (N_12449,N_12361,N_12273);
nor U12450 (N_12450,N_12357,N_12295);
or U12451 (N_12451,N_12347,N_12303);
nor U12452 (N_12452,N_12309,N_12288);
and U12453 (N_12453,N_12336,N_12272);
and U12454 (N_12454,N_12283,N_12256);
or U12455 (N_12455,N_12329,N_12294);
xnor U12456 (N_12456,N_12324,N_12291);
nor U12457 (N_12457,N_12365,N_12311);
or U12458 (N_12458,N_12319,N_12338);
and U12459 (N_12459,N_12365,N_12324);
or U12460 (N_12460,N_12313,N_12263);
and U12461 (N_12461,N_12312,N_12366);
or U12462 (N_12462,N_12289,N_12334);
nand U12463 (N_12463,N_12327,N_12328);
nor U12464 (N_12464,N_12348,N_12354);
nor U12465 (N_12465,N_12330,N_12296);
or U12466 (N_12466,N_12289,N_12283);
xor U12467 (N_12467,N_12352,N_12267);
or U12468 (N_12468,N_12268,N_12269);
nand U12469 (N_12469,N_12332,N_12369);
nand U12470 (N_12470,N_12374,N_12254);
nand U12471 (N_12471,N_12355,N_12359);
and U12472 (N_12472,N_12311,N_12318);
xnor U12473 (N_12473,N_12292,N_12283);
nor U12474 (N_12474,N_12292,N_12330);
or U12475 (N_12475,N_12291,N_12295);
nor U12476 (N_12476,N_12307,N_12365);
xnor U12477 (N_12477,N_12293,N_12330);
nor U12478 (N_12478,N_12264,N_12266);
xnor U12479 (N_12479,N_12345,N_12285);
and U12480 (N_12480,N_12253,N_12274);
nand U12481 (N_12481,N_12353,N_12298);
nor U12482 (N_12482,N_12368,N_12328);
nor U12483 (N_12483,N_12366,N_12287);
nand U12484 (N_12484,N_12272,N_12358);
xor U12485 (N_12485,N_12272,N_12357);
or U12486 (N_12486,N_12287,N_12277);
nand U12487 (N_12487,N_12276,N_12309);
nor U12488 (N_12488,N_12284,N_12338);
nor U12489 (N_12489,N_12312,N_12300);
nand U12490 (N_12490,N_12294,N_12352);
xnor U12491 (N_12491,N_12313,N_12300);
xnor U12492 (N_12492,N_12347,N_12362);
nor U12493 (N_12493,N_12319,N_12252);
and U12494 (N_12494,N_12294,N_12262);
and U12495 (N_12495,N_12356,N_12339);
and U12496 (N_12496,N_12349,N_12339);
or U12497 (N_12497,N_12328,N_12319);
and U12498 (N_12498,N_12346,N_12296);
or U12499 (N_12499,N_12303,N_12370);
xnor U12500 (N_12500,N_12385,N_12493);
xor U12501 (N_12501,N_12459,N_12478);
nand U12502 (N_12502,N_12436,N_12416);
xnor U12503 (N_12503,N_12384,N_12454);
xnor U12504 (N_12504,N_12442,N_12488);
and U12505 (N_12505,N_12407,N_12461);
xor U12506 (N_12506,N_12393,N_12420);
nor U12507 (N_12507,N_12499,N_12379);
nand U12508 (N_12508,N_12441,N_12470);
nor U12509 (N_12509,N_12380,N_12398);
nor U12510 (N_12510,N_12490,N_12446);
or U12511 (N_12511,N_12494,N_12415);
nor U12512 (N_12512,N_12486,N_12422);
and U12513 (N_12513,N_12472,N_12451);
or U12514 (N_12514,N_12438,N_12432);
nor U12515 (N_12515,N_12390,N_12444);
and U12516 (N_12516,N_12387,N_12408);
xor U12517 (N_12517,N_12411,N_12391);
nor U12518 (N_12518,N_12464,N_12491);
nor U12519 (N_12519,N_12463,N_12437);
and U12520 (N_12520,N_12495,N_12401);
xor U12521 (N_12521,N_12456,N_12397);
nor U12522 (N_12522,N_12419,N_12435);
nor U12523 (N_12523,N_12487,N_12479);
nand U12524 (N_12524,N_12378,N_12413);
xnor U12525 (N_12525,N_12458,N_12429);
and U12526 (N_12526,N_12377,N_12400);
and U12527 (N_12527,N_12434,N_12439);
xor U12528 (N_12528,N_12484,N_12498);
nor U12529 (N_12529,N_12383,N_12445);
or U12530 (N_12530,N_12403,N_12406);
nor U12531 (N_12531,N_12449,N_12404);
or U12532 (N_12532,N_12427,N_12424);
nor U12533 (N_12533,N_12417,N_12430);
xnor U12534 (N_12534,N_12423,N_12389);
xor U12535 (N_12535,N_12447,N_12410);
or U12536 (N_12536,N_12497,N_12381);
nor U12537 (N_12537,N_12477,N_12496);
xor U12538 (N_12538,N_12482,N_12450);
nand U12539 (N_12539,N_12448,N_12409);
and U12540 (N_12540,N_12376,N_12460);
or U12541 (N_12541,N_12375,N_12428);
and U12542 (N_12542,N_12467,N_12412);
and U12543 (N_12543,N_12426,N_12433);
and U12544 (N_12544,N_12457,N_12485);
or U12545 (N_12545,N_12453,N_12402);
or U12546 (N_12546,N_12462,N_12476);
xor U12547 (N_12547,N_12471,N_12392);
xnor U12548 (N_12548,N_12431,N_12394);
nand U12549 (N_12549,N_12396,N_12468);
nor U12550 (N_12550,N_12421,N_12483);
nor U12551 (N_12551,N_12474,N_12388);
or U12552 (N_12552,N_12405,N_12399);
nor U12553 (N_12553,N_12443,N_12466);
xor U12554 (N_12554,N_12418,N_12425);
or U12555 (N_12555,N_12452,N_12440);
nor U12556 (N_12556,N_12489,N_12492);
nor U12557 (N_12557,N_12386,N_12480);
nand U12558 (N_12558,N_12475,N_12473);
nor U12559 (N_12559,N_12455,N_12481);
nor U12560 (N_12560,N_12382,N_12414);
xnor U12561 (N_12561,N_12395,N_12465);
nand U12562 (N_12562,N_12469,N_12399);
xor U12563 (N_12563,N_12410,N_12407);
and U12564 (N_12564,N_12430,N_12386);
and U12565 (N_12565,N_12392,N_12462);
and U12566 (N_12566,N_12423,N_12492);
xor U12567 (N_12567,N_12471,N_12448);
nor U12568 (N_12568,N_12456,N_12376);
nor U12569 (N_12569,N_12420,N_12412);
nor U12570 (N_12570,N_12401,N_12399);
and U12571 (N_12571,N_12412,N_12489);
nand U12572 (N_12572,N_12457,N_12483);
and U12573 (N_12573,N_12489,N_12440);
nand U12574 (N_12574,N_12446,N_12480);
or U12575 (N_12575,N_12446,N_12489);
nand U12576 (N_12576,N_12407,N_12390);
nor U12577 (N_12577,N_12496,N_12406);
and U12578 (N_12578,N_12382,N_12412);
nor U12579 (N_12579,N_12499,N_12397);
or U12580 (N_12580,N_12457,N_12382);
nand U12581 (N_12581,N_12440,N_12487);
or U12582 (N_12582,N_12422,N_12378);
nand U12583 (N_12583,N_12470,N_12396);
nor U12584 (N_12584,N_12420,N_12410);
xor U12585 (N_12585,N_12413,N_12431);
or U12586 (N_12586,N_12481,N_12482);
or U12587 (N_12587,N_12411,N_12432);
nand U12588 (N_12588,N_12457,N_12477);
and U12589 (N_12589,N_12451,N_12407);
xor U12590 (N_12590,N_12439,N_12444);
xor U12591 (N_12591,N_12478,N_12420);
nand U12592 (N_12592,N_12379,N_12389);
xnor U12593 (N_12593,N_12435,N_12376);
xnor U12594 (N_12594,N_12488,N_12417);
nand U12595 (N_12595,N_12379,N_12405);
or U12596 (N_12596,N_12489,N_12425);
nor U12597 (N_12597,N_12492,N_12482);
xnor U12598 (N_12598,N_12482,N_12457);
or U12599 (N_12599,N_12481,N_12389);
xnor U12600 (N_12600,N_12471,N_12381);
and U12601 (N_12601,N_12471,N_12493);
nor U12602 (N_12602,N_12447,N_12443);
nand U12603 (N_12603,N_12489,N_12480);
xor U12604 (N_12604,N_12493,N_12466);
nor U12605 (N_12605,N_12488,N_12441);
nand U12606 (N_12606,N_12406,N_12437);
nand U12607 (N_12607,N_12474,N_12429);
nand U12608 (N_12608,N_12439,N_12468);
xor U12609 (N_12609,N_12493,N_12404);
or U12610 (N_12610,N_12443,N_12378);
or U12611 (N_12611,N_12499,N_12458);
xnor U12612 (N_12612,N_12398,N_12393);
nand U12613 (N_12613,N_12411,N_12441);
and U12614 (N_12614,N_12427,N_12421);
nor U12615 (N_12615,N_12392,N_12432);
xor U12616 (N_12616,N_12377,N_12424);
or U12617 (N_12617,N_12447,N_12480);
and U12618 (N_12618,N_12381,N_12398);
and U12619 (N_12619,N_12407,N_12413);
and U12620 (N_12620,N_12444,N_12430);
nand U12621 (N_12621,N_12391,N_12430);
and U12622 (N_12622,N_12390,N_12425);
nand U12623 (N_12623,N_12438,N_12404);
nand U12624 (N_12624,N_12412,N_12437);
xnor U12625 (N_12625,N_12537,N_12525);
and U12626 (N_12626,N_12538,N_12571);
nand U12627 (N_12627,N_12556,N_12569);
or U12628 (N_12628,N_12588,N_12585);
and U12629 (N_12629,N_12591,N_12518);
nand U12630 (N_12630,N_12531,N_12532);
nor U12631 (N_12631,N_12545,N_12511);
or U12632 (N_12632,N_12586,N_12610);
and U12633 (N_12633,N_12616,N_12582);
nand U12634 (N_12634,N_12554,N_12590);
xor U12635 (N_12635,N_12611,N_12551);
and U12636 (N_12636,N_12622,N_12606);
or U12637 (N_12637,N_12614,N_12512);
nand U12638 (N_12638,N_12523,N_12605);
nor U12639 (N_12639,N_12504,N_12548);
nand U12640 (N_12640,N_12509,N_12557);
xnor U12641 (N_12641,N_12516,N_12562);
or U12642 (N_12642,N_12520,N_12597);
and U12643 (N_12643,N_12600,N_12553);
nand U12644 (N_12644,N_12593,N_12601);
xnor U12645 (N_12645,N_12564,N_12552);
nand U12646 (N_12646,N_12527,N_12533);
nor U12647 (N_12647,N_12607,N_12570);
and U12648 (N_12648,N_12535,N_12596);
or U12649 (N_12649,N_12568,N_12623);
nor U12650 (N_12650,N_12580,N_12617);
xor U12651 (N_12651,N_12608,N_12624);
or U12652 (N_12652,N_12508,N_12522);
xor U12653 (N_12653,N_12543,N_12526);
nand U12654 (N_12654,N_12502,N_12542);
or U12655 (N_12655,N_12540,N_12565);
or U12656 (N_12656,N_12618,N_12621);
nor U12657 (N_12657,N_12544,N_12576);
nor U12658 (N_12658,N_12575,N_12592);
and U12659 (N_12659,N_12501,N_12589);
nand U12660 (N_12660,N_12563,N_12581);
and U12661 (N_12661,N_12587,N_12549);
xnor U12662 (N_12662,N_12620,N_12609);
nor U12663 (N_12663,N_12612,N_12615);
or U12664 (N_12664,N_12559,N_12574);
xor U12665 (N_12665,N_12602,N_12524);
nand U12666 (N_12666,N_12536,N_12547);
or U12667 (N_12667,N_12555,N_12546);
nor U12668 (N_12668,N_12503,N_12550);
and U12669 (N_12669,N_12573,N_12579);
xnor U12670 (N_12670,N_12519,N_12595);
nand U12671 (N_12671,N_12515,N_12594);
nand U12672 (N_12672,N_12500,N_12513);
xnor U12673 (N_12673,N_12584,N_12521);
nand U12674 (N_12674,N_12507,N_12541);
nand U12675 (N_12675,N_12599,N_12530);
xnor U12676 (N_12676,N_12510,N_12572);
nor U12677 (N_12677,N_12567,N_12514);
and U12678 (N_12678,N_12558,N_12517);
xnor U12679 (N_12679,N_12577,N_12528);
xnor U12680 (N_12680,N_12603,N_12560);
or U12681 (N_12681,N_12566,N_12506);
xnor U12682 (N_12682,N_12598,N_12613);
and U12683 (N_12683,N_12534,N_12505);
nor U12684 (N_12684,N_12583,N_12539);
and U12685 (N_12685,N_12604,N_12561);
nor U12686 (N_12686,N_12578,N_12619);
nand U12687 (N_12687,N_12529,N_12592);
nor U12688 (N_12688,N_12554,N_12514);
nor U12689 (N_12689,N_12609,N_12611);
xor U12690 (N_12690,N_12556,N_12571);
and U12691 (N_12691,N_12528,N_12621);
or U12692 (N_12692,N_12511,N_12601);
and U12693 (N_12693,N_12579,N_12570);
and U12694 (N_12694,N_12623,N_12560);
nor U12695 (N_12695,N_12581,N_12582);
and U12696 (N_12696,N_12525,N_12618);
xor U12697 (N_12697,N_12529,N_12564);
or U12698 (N_12698,N_12578,N_12524);
and U12699 (N_12699,N_12582,N_12617);
nor U12700 (N_12700,N_12525,N_12602);
or U12701 (N_12701,N_12541,N_12609);
xnor U12702 (N_12702,N_12567,N_12589);
and U12703 (N_12703,N_12601,N_12615);
nand U12704 (N_12704,N_12583,N_12529);
or U12705 (N_12705,N_12588,N_12593);
or U12706 (N_12706,N_12606,N_12572);
or U12707 (N_12707,N_12531,N_12613);
nand U12708 (N_12708,N_12552,N_12502);
xor U12709 (N_12709,N_12608,N_12619);
and U12710 (N_12710,N_12602,N_12568);
and U12711 (N_12711,N_12508,N_12587);
or U12712 (N_12712,N_12575,N_12605);
nor U12713 (N_12713,N_12525,N_12579);
or U12714 (N_12714,N_12500,N_12608);
and U12715 (N_12715,N_12537,N_12520);
nor U12716 (N_12716,N_12558,N_12554);
nand U12717 (N_12717,N_12527,N_12559);
nor U12718 (N_12718,N_12577,N_12578);
nand U12719 (N_12719,N_12587,N_12615);
nand U12720 (N_12720,N_12568,N_12603);
or U12721 (N_12721,N_12504,N_12522);
and U12722 (N_12722,N_12524,N_12598);
nor U12723 (N_12723,N_12584,N_12562);
and U12724 (N_12724,N_12561,N_12614);
nand U12725 (N_12725,N_12531,N_12519);
or U12726 (N_12726,N_12553,N_12518);
nor U12727 (N_12727,N_12606,N_12620);
xnor U12728 (N_12728,N_12547,N_12598);
nor U12729 (N_12729,N_12617,N_12594);
and U12730 (N_12730,N_12611,N_12583);
nand U12731 (N_12731,N_12511,N_12594);
and U12732 (N_12732,N_12594,N_12574);
and U12733 (N_12733,N_12515,N_12538);
nand U12734 (N_12734,N_12593,N_12542);
nand U12735 (N_12735,N_12522,N_12523);
or U12736 (N_12736,N_12562,N_12597);
nor U12737 (N_12737,N_12583,N_12580);
nand U12738 (N_12738,N_12535,N_12563);
nor U12739 (N_12739,N_12613,N_12570);
nor U12740 (N_12740,N_12530,N_12531);
nor U12741 (N_12741,N_12553,N_12610);
nor U12742 (N_12742,N_12573,N_12606);
nand U12743 (N_12743,N_12623,N_12500);
or U12744 (N_12744,N_12612,N_12560);
nor U12745 (N_12745,N_12508,N_12590);
and U12746 (N_12746,N_12525,N_12521);
xor U12747 (N_12747,N_12550,N_12552);
nand U12748 (N_12748,N_12541,N_12532);
or U12749 (N_12749,N_12503,N_12607);
or U12750 (N_12750,N_12661,N_12662);
or U12751 (N_12751,N_12694,N_12649);
and U12752 (N_12752,N_12627,N_12660);
nand U12753 (N_12753,N_12748,N_12744);
nor U12754 (N_12754,N_12680,N_12646);
nand U12755 (N_12755,N_12665,N_12645);
xor U12756 (N_12756,N_12650,N_12629);
nand U12757 (N_12757,N_12667,N_12656);
and U12758 (N_12758,N_12709,N_12677);
xnor U12759 (N_12759,N_12632,N_12685);
nor U12760 (N_12760,N_12676,N_12653);
nor U12761 (N_12761,N_12711,N_12712);
xor U12762 (N_12762,N_12700,N_12637);
nand U12763 (N_12763,N_12643,N_12733);
nor U12764 (N_12764,N_12657,N_12678);
nand U12765 (N_12765,N_12719,N_12738);
or U12766 (N_12766,N_12701,N_12647);
or U12767 (N_12767,N_12716,N_12683);
xor U12768 (N_12768,N_12745,N_12681);
and U12769 (N_12769,N_12742,N_12729);
xor U12770 (N_12770,N_12731,N_12724);
or U12771 (N_12771,N_12707,N_12634);
and U12772 (N_12772,N_12651,N_12655);
or U12773 (N_12773,N_12674,N_12723);
or U12774 (N_12774,N_12628,N_12699);
or U12775 (N_12775,N_12713,N_12704);
or U12776 (N_12776,N_12644,N_12743);
and U12777 (N_12777,N_12717,N_12714);
xor U12778 (N_12778,N_12664,N_12659);
and U12779 (N_12779,N_12725,N_12691);
xor U12780 (N_12780,N_12720,N_12641);
or U12781 (N_12781,N_12675,N_12658);
or U12782 (N_12782,N_12706,N_12630);
or U12783 (N_12783,N_12692,N_12715);
and U12784 (N_12784,N_12626,N_12746);
and U12785 (N_12785,N_12687,N_12686);
nor U12786 (N_12786,N_12696,N_12631);
nand U12787 (N_12787,N_12741,N_12654);
nor U12788 (N_12788,N_12633,N_12652);
or U12789 (N_12789,N_12670,N_12672);
nor U12790 (N_12790,N_12684,N_12697);
nand U12791 (N_12791,N_12702,N_12727);
nand U12792 (N_12792,N_12705,N_12673);
xor U12793 (N_12793,N_12668,N_12639);
or U12794 (N_12794,N_12726,N_12747);
xor U12795 (N_12795,N_12749,N_12737);
and U12796 (N_12796,N_12735,N_12690);
or U12797 (N_12797,N_12636,N_12635);
or U12798 (N_12798,N_12642,N_12703);
nor U12799 (N_12799,N_12679,N_12698);
or U12800 (N_12800,N_12734,N_12638);
xnor U12801 (N_12801,N_12722,N_12671);
or U12802 (N_12802,N_12739,N_12689);
and U12803 (N_12803,N_12669,N_12718);
and U12804 (N_12804,N_12736,N_12732);
and U12805 (N_12805,N_12648,N_12640);
and U12806 (N_12806,N_12740,N_12730);
nor U12807 (N_12807,N_12688,N_12663);
nand U12808 (N_12808,N_12682,N_12666);
and U12809 (N_12809,N_12728,N_12710);
or U12810 (N_12810,N_12708,N_12693);
and U12811 (N_12811,N_12625,N_12721);
or U12812 (N_12812,N_12695,N_12647);
nor U12813 (N_12813,N_12697,N_12681);
xnor U12814 (N_12814,N_12702,N_12638);
and U12815 (N_12815,N_12700,N_12716);
nand U12816 (N_12816,N_12719,N_12706);
and U12817 (N_12817,N_12713,N_12675);
and U12818 (N_12818,N_12731,N_12734);
nor U12819 (N_12819,N_12694,N_12628);
nor U12820 (N_12820,N_12714,N_12646);
nor U12821 (N_12821,N_12677,N_12625);
nor U12822 (N_12822,N_12627,N_12691);
and U12823 (N_12823,N_12749,N_12643);
nand U12824 (N_12824,N_12749,N_12668);
nor U12825 (N_12825,N_12637,N_12730);
xor U12826 (N_12826,N_12636,N_12696);
xnor U12827 (N_12827,N_12706,N_12670);
or U12828 (N_12828,N_12691,N_12704);
and U12829 (N_12829,N_12712,N_12652);
and U12830 (N_12830,N_12682,N_12687);
nand U12831 (N_12831,N_12741,N_12721);
xor U12832 (N_12832,N_12644,N_12713);
nand U12833 (N_12833,N_12659,N_12749);
nand U12834 (N_12834,N_12685,N_12660);
xor U12835 (N_12835,N_12631,N_12727);
nor U12836 (N_12836,N_12730,N_12710);
nand U12837 (N_12837,N_12746,N_12660);
xor U12838 (N_12838,N_12681,N_12685);
or U12839 (N_12839,N_12695,N_12632);
and U12840 (N_12840,N_12712,N_12726);
xor U12841 (N_12841,N_12684,N_12688);
and U12842 (N_12842,N_12738,N_12636);
or U12843 (N_12843,N_12680,N_12748);
and U12844 (N_12844,N_12720,N_12634);
nor U12845 (N_12845,N_12716,N_12631);
nand U12846 (N_12846,N_12702,N_12678);
nand U12847 (N_12847,N_12652,N_12655);
or U12848 (N_12848,N_12745,N_12630);
nand U12849 (N_12849,N_12676,N_12714);
nor U12850 (N_12850,N_12707,N_12670);
nand U12851 (N_12851,N_12662,N_12749);
or U12852 (N_12852,N_12734,N_12745);
and U12853 (N_12853,N_12695,N_12713);
nor U12854 (N_12854,N_12691,N_12733);
nand U12855 (N_12855,N_12633,N_12666);
nor U12856 (N_12856,N_12663,N_12666);
nand U12857 (N_12857,N_12688,N_12654);
nor U12858 (N_12858,N_12725,N_12741);
or U12859 (N_12859,N_12667,N_12724);
xor U12860 (N_12860,N_12644,N_12645);
xor U12861 (N_12861,N_12675,N_12649);
or U12862 (N_12862,N_12671,N_12704);
and U12863 (N_12863,N_12709,N_12676);
and U12864 (N_12864,N_12725,N_12695);
xnor U12865 (N_12865,N_12643,N_12728);
nor U12866 (N_12866,N_12733,N_12709);
nor U12867 (N_12867,N_12737,N_12663);
xnor U12868 (N_12868,N_12668,N_12632);
xor U12869 (N_12869,N_12740,N_12670);
xnor U12870 (N_12870,N_12709,N_12726);
and U12871 (N_12871,N_12742,N_12712);
and U12872 (N_12872,N_12741,N_12681);
nor U12873 (N_12873,N_12628,N_12686);
nor U12874 (N_12874,N_12713,N_12721);
nor U12875 (N_12875,N_12865,N_12873);
and U12876 (N_12876,N_12780,N_12851);
nand U12877 (N_12877,N_12765,N_12850);
or U12878 (N_12878,N_12868,N_12824);
xor U12879 (N_12879,N_12769,N_12825);
nor U12880 (N_12880,N_12821,N_12786);
nand U12881 (N_12881,N_12866,N_12844);
xnor U12882 (N_12882,N_12760,N_12797);
nand U12883 (N_12883,N_12814,N_12764);
xor U12884 (N_12884,N_12842,N_12826);
nand U12885 (N_12885,N_12773,N_12855);
nor U12886 (N_12886,N_12833,N_12792);
and U12887 (N_12887,N_12794,N_12830);
nor U12888 (N_12888,N_12864,N_12858);
nor U12889 (N_12889,N_12854,N_12845);
or U12890 (N_12890,N_12766,N_12785);
nand U12891 (N_12891,N_12860,N_12770);
nor U12892 (N_12892,N_12812,N_12846);
or U12893 (N_12893,N_12840,N_12781);
nor U12894 (N_12894,N_12822,N_12799);
and U12895 (N_12895,N_12782,N_12834);
xnor U12896 (N_12896,N_12798,N_12872);
and U12897 (N_12897,N_12828,N_12807);
nor U12898 (N_12898,N_12863,N_12784);
and U12899 (N_12899,N_12874,N_12813);
xnor U12900 (N_12900,N_12837,N_12835);
and U12901 (N_12901,N_12832,N_12790);
nand U12902 (N_12902,N_12804,N_12771);
and U12903 (N_12903,N_12796,N_12757);
and U12904 (N_12904,N_12778,N_12817);
nor U12905 (N_12905,N_12809,N_12820);
nand U12906 (N_12906,N_12831,N_12843);
nor U12907 (N_12907,N_12827,N_12777);
nand U12908 (N_12908,N_12756,N_12763);
and U12909 (N_12909,N_12801,N_12779);
or U12910 (N_12910,N_12839,N_12793);
nor U12911 (N_12911,N_12788,N_12762);
and U12912 (N_12912,N_12767,N_12751);
or U12913 (N_12913,N_12852,N_12759);
or U12914 (N_12914,N_12774,N_12823);
or U12915 (N_12915,N_12805,N_12768);
or U12916 (N_12916,N_12847,N_12857);
nand U12917 (N_12917,N_12811,N_12836);
and U12918 (N_12918,N_12841,N_12856);
xor U12919 (N_12919,N_12867,N_12861);
nor U12920 (N_12920,N_12829,N_12808);
and U12921 (N_12921,N_12815,N_12870);
nand U12922 (N_12922,N_12871,N_12753);
or U12923 (N_12923,N_12819,N_12806);
or U12924 (N_12924,N_12810,N_12750);
nor U12925 (N_12925,N_12818,N_12848);
nor U12926 (N_12926,N_12791,N_12816);
and U12927 (N_12927,N_12758,N_12783);
nand U12928 (N_12928,N_12789,N_12853);
nor U12929 (N_12929,N_12800,N_12849);
and U12930 (N_12930,N_12869,N_12795);
nor U12931 (N_12931,N_12838,N_12787);
nor U12932 (N_12932,N_12752,N_12862);
nor U12933 (N_12933,N_12761,N_12775);
or U12934 (N_12934,N_12776,N_12802);
or U12935 (N_12935,N_12859,N_12803);
xor U12936 (N_12936,N_12755,N_12754);
nand U12937 (N_12937,N_12772,N_12872);
nor U12938 (N_12938,N_12751,N_12857);
nor U12939 (N_12939,N_12764,N_12758);
and U12940 (N_12940,N_12812,N_12760);
xor U12941 (N_12941,N_12803,N_12844);
and U12942 (N_12942,N_12854,N_12783);
nor U12943 (N_12943,N_12843,N_12861);
nand U12944 (N_12944,N_12820,N_12784);
or U12945 (N_12945,N_12871,N_12782);
xnor U12946 (N_12946,N_12786,N_12849);
or U12947 (N_12947,N_12847,N_12831);
and U12948 (N_12948,N_12796,N_12774);
nand U12949 (N_12949,N_12801,N_12768);
nand U12950 (N_12950,N_12765,N_12754);
or U12951 (N_12951,N_12854,N_12792);
nor U12952 (N_12952,N_12764,N_12809);
nand U12953 (N_12953,N_12785,N_12802);
nand U12954 (N_12954,N_12812,N_12763);
xnor U12955 (N_12955,N_12781,N_12832);
xnor U12956 (N_12956,N_12800,N_12873);
and U12957 (N_12957,N_12773,N_12759);
or U12958 (N_12958,N_12787,N_12847);
or U12959 (N_12959,N_12837,N_12859);
and U12960 (N_12960,N_12863,N_12868);
or U12961 (N_12961,N_12756,N_12846);
nor U12962 (N_12962,N_12849,N_12790);
or U12963 (N_12963,N_12753,N_12812);
and U12964 (N_12964,N_12752,N_12753);
and U12965 (N_12965,N_12811,N_12788);
nand U12966 (N_12966,N_12853,N_12846);
or U12967 (N_12967,N_12870,N_12800);
nor U12968 (N_12968,N_12826,N_12805);
nand U12969 (N_12969,N_12831,N_12797);
and U12970 (N_12970,N_12785,N_12774);
or U12971 (N_12971,N_12842,N_12846);
xor U12972 (N_12972,N_12751,N_12799);
nor U12973 (N_12973,N_12794,N_12759);
nand U12974 (N_12974,N_12826,N_12751);
xor U12975 (N_12975,N_12841,N_12851);
or U12976 (N_12976,N_12820,N_12854);
and U12977 (N_12977,N_12867,N_12871);
nor U12978 (N_12978,N_12811,N_12813);
nor U12979 (N_12979,N_12769,N_12802);
or U12980 (N_12980,N_12798,N_12800);
and U12981 (N_12981,N_12796,N_12840);
or U12982 (N_12982,N_12756,N_12812);
or U12983 (N_12983,N_12862,N_12777);
or U12984 (N_12984,N_12799,N_12859);
nor U12985 (N_12985,N_12847,N_12779);
and U12986 (N_12986,N_12866,N_12869);
nand U12987 (N_12987,N_12834,N_12751);
xnor U12988 (N_12988,N_12751,N_12873);
or U12989 (N_12989,N_12836,N_12848);
nor U12990 (N_12990,N_12792,N_12799);
xnor U12991 (N_12991,N_12798,N_12777);
xor U12992 (N_12992,N_12866,N_12771);
nand U12993 (N_12993,N_12807,N_12858);
nand U12994 (N_12994,N_12766,N_12801);
and U12995 (N_12995,N_12791,N_12770);
and U12996 (N_12996,N_12853,N_12834);
nor U12997 (N_12997,N_12818,N_12759);
nand U12998 (N_12998,N_12837,N_12870);
or U12999 (N_12999,N_12836,N_12862);
nor U13000 (N_13000,N_12887,N_12877);
xor U13001 (N_13001,N_12938,N_12906);
nor U13002 (N_13002,N_12921,N_12935);
and U13003 (N_13003,N_12946,N_12965);
or U13004 (N_13004,N_12949,N_12882);
xor U13005 (N_13005,N_12988,N_12976);
xnor U13006 (N_13006,N_12914,N_12987);
xnor U13007 (N_13007,N_12876,N_12964);
nand U13008 (N_13008,N_12885,N_12968);
nor U13009 (N_13009,N_12951,N_12929);
and U13010 (N_13010,N_12989,N_12958);
and U13011 (N_13011,N_12923,N_12904);
xor U13012 (N_13012,N_12960,N_12886);
nor U13013 (N_13013,N_12970,N_12902);
and U13014 (N_13014,N_12937,N_12966);
xor U13015 (N_13015,N_12894,N_12920);
nor U13016 (N_13016,N_12974,N_12953);
nor U13017 (N_13017,N_12930,N_12878);
xor U13018 (N_13018,N_12925,N_12909);
xnor U13019 (N_13019,N_12950,N_12985);
nor U13020 (N_13020,N_12880,N_12944);
and U13021 (N_13021,N_12997,N_12924);
and U13022 (N_13022,N_12912,N_12900);
nor U13023 (N_13023,N_12922,N_12978);
xor U13024 (N_13024,N_12954,N_12995);
nand U13025 (N_13025,N_12975,N_12895);
xnor U13026 (N_13026,N_12969,N_12948);
nand U13027 (N_13027,N_12963,N_12907);
nor U13028 (N_13028,N_12955,N_12959);
xnor U13029 (N_13029,N_12986,N_12957);
or U13030 (N_13030,N_12883,N_12984);
or U13031 (N_13031,N_12961,N_12996);
nor U13032 (N_13032,N_12947,N_12982);
nor U13033 (N_13033,N_12992,N_12967);
nor U13034 (N_13034,N_12980,N_12896);
and U13035 (N_13035,N_12939,N_12956);
and U13036 (N_13036,N_12940,N_12893);
xor U13037 (N_13037,N_12915,N_12875);
nand U13038 (N_13038,N_12898,N_12927);
xnor U13039 (N_13039,N_12881,N_12983);
nor U13040 (N_13040,N_12903,N_12932);
nor U13041 (N_13041,N_12981,N_12977);
or U13042 (N_13042,N_12879,N_12919);
and U13043 (N_13043,N_12962,N_12998);
nor U13044 (N_13044,N_12941,N_12891);
nand U13045 (N_13045,N_12918,N_12908);
and U13046 (N_13046,N_12942,N_12926);
and U13047 (N_13047,N_12979,N_12972);
nand U13048 (N_13048,N_12936,N_12931);
and U13049 (N_13049,N_12911,N_12934);
xnor U13050 (N_13050,N_12913,N_12892);
xor U13051 (N_13051,N_12916,N_12917);
nand U13052 (N_13052,N_12890,N_12897);
nor U13053 (N_13053,N_12952,N_12999);
and U13054 (N_13054,N_12905,N_12884);
xnor U13055 (N_13055,N_12973,N_12910);
nor U13056 (N_13056,N_12945,N_12971);
nor U13057 (N_13057,N_12888,N_12889);
nor U13058 (N_13058,N_12928,N_12991);
nor U13059 (N_13059,N_12993,N_12899);
nor U13060 (N_13060,N_12933,N_12994);
xor U13061 (N_13061,N_12901,N_12990);
nor U13062 (N_13062,N_12943,N_12919);
nor U13063 (N_13063,N_12903,N_12975);
xor U13064 (N_13064,N_12980,N_12970);
and U13065 (N_13065,N_12923,N_12896);
nand U13066 (N_13066,N_12999,N_12879);
xor U13067 (N_13067,N_12957,N_12917);
and U13068 (N_13068,N_12952,N_12888);
nor U13069 (N_13069,N_12990,N_12979);
nor U13070 (N_13070,N_12960,N_12984);
or U13071 (N_13071,N_12931,N_12891);
nand U13072 (N_13072,N_12887,N_12898);
xor U13073 (N_13073,N_12899,N_12915);
nand U13074 (N_13074,N_12978,N_12966);
or U13075 (N_13075,N_12929,N_12902);
or U13076 (N_13076,N_12968,N_12986);
xor U13077 (N_13077,N_12975,N_12915);
or U13078 (N_13078,N_12931,N_12976);
xnor U13079 (N_13079,N_12884,N_12978);
nand U13080 (N_13080,N_12944,N_12966);
nor U13081 (N_13081,N_12902,N_12999);
or U13082 (N_13082,N_12881,N_12918);
and U13083 (N_13083,N_12970,N_12968);
and U13084 (N_13084,N_12973,N_12905);
or U13085 (N_13085,N_12877,N_12937);
and U13086 (N_13086,N_12878,N_12904);
nand U13087 (N_13087,N_12911,N_12930);
or U13088 (N_13088,N_12995,N_12955);
or U13089 (N_13089,N_12920,N_12992);
or U13090 (N_13090,N_12997,N_12990);
nand U13091 (N_13091,N_12916,N_12989);
and U13092 (N_13092,N_12958,N_12915);
or U13093 (N_13093,N_12993,N_12898);
nor U13094 (N_13094,N_12884,N_12915);
nand U13095 (N_13095,N_12895,N_12954);
and U13096 (N_13096,N_12928,N_12987);
nor U13097 (N_13097,N_12983,N_12928);
xnor U13098 (N_13098,N_12946,N_12910);
nor U13099 (N_13099,N_12918,N_12914);
nand U13100 (N_13100,N_12959,N_12896);
and U13101 (N_13101,N_12875,N_12926);
nand U13102 (N_13102,N_12883,N_12911);
nor U13103 (N_13103,N_12997,N_12917);
nand U13104 (N_13104,N_12945,N_12878);
and U13105 (N_13105,N_12903,N_12944);
xnor U13106 (N_13106,N_12889,N_12902);
or U13107 (N_13107,N_12917,N_12908);
nor U13108 (N_13108,N_12938,N_12901);
nor U13109 (N_13109,N_12902,N_12995);
nor U13110 (N_13110,N_12926,N_12972);
or U13111 (N_13111,N_12904,N_12884);
xnor U13112 (N_13112,N_12877,N_12996);
xnor U13113 (N_13113,N_12996,N_12941);
nand U13114 (N_13114,N_12911,N_12880);
nand U13115 (N_13115,N_12956,N_12894);
nand U13116 (N_13116,N_12985,N_12884);
or U13117 (N_13117,N_12931,N_12879);
or U13118 (N_13118,N_12977,N_12955);
nor U13119 (N_13119,N_12887,N_12933);
nand U13120 (N_13120,N_12882,N_12969);
and U13121 (N_13121,N_12908,N_12915);
xnor U13122 (N_13122,N_12882,N_12905);
and U13123 (N_13123,N_12974,N_12977);
xor U13124 (N_13124,N_12912,N_12941);
xor U13125 (N_13125,N_13119,N_13065);
nand U13126 (N_13126,N_13075,N_13063);
nand U13127 (N_13127,N_13034,N_13019);
and U13128 (N_13128,N_13056,N_13047);
nand U13129 (N_13129,N_13016,N_13078);
and U13130 (N_13130,N_13071,N_13114);
and U13131 (N_13131,N_13074,N_13030);
and U13132 (N_13132,N_13124,N_13069);
or U13133 (N_13133,N_13102,N_13046);
or U13134 (N_13134,N_13032,N_13039);
or U13135 (N_13135,N_13120,N_13084);
and U13136 (N_13136,N_13038,N_13023);
or U13137 (N_13137,N_13080,N_13054);
and U13138 (N_13138,N_13011,N_13089);
xnor U13139 (N_13139,N_13113,N_13051);
nor U13140 (N_13140,N_13007,N_13029);
and U13141 (N_13141,N_13108,N_13042);
or U13142 (N_13142,N_13015,N_13024);
xnor U13143 (N_13143,N_13053,N_13044);
nand U13144 (N_13144,N_13123,N_13076);
and U13145 (N_13145,N_13107,N_13027);
xor U13146 (N_13146,N_13079,N_13087);
and U13147 (N_13147,N_13021,N_13101);
or U13148 (N_13148,N_13048,N_13122);
nor U13149 (N_13149,N_13090,N_13104);
nor U13150 (N_13150,N_13064,N_13000);
xor U13151 (N_13151,N_13018,N_13014);
xnor U13152 (N_13152,N_13073,N_13070);
or U13153 (N_13153,N_13105,N_13055);
or U13154 (N_13154,N_13068,N_13095);
and U13155 (N_13155,N_13077,N_13092);
nand U13156 (N_13156,N_13012,N_13111);
nor U13157 (N_13157,N_13002,N_13022);
xnor U13158 (N_13158,N_13058,N_13109);
or U13159 (N_13159,N_13020,N_13086);
and U13160 (N_13160,N_13040,N_13017);
or U13161 (N_13161,N_13088,N_13043);
nand U13162 (N_13162,N_13062,N_13010);
and U13163 (N_13163,N_13049,N_13085);
or U13164 (N_13164,N_13033,N_13094);
nand U13165 (N_13165,N_13091,N_13118);
xor U13166 (N_13166,N_13110,N_13083);
xnor U13167 (N_13167,N_13061,N_13060);
or U13168 (N_13168,N_13045,N_13041);
nand U13169 (N_13169,N_13117,N_13100);
nor U13170 (N_13170,N_13005,N_13006);
nor U13171 (N_13171,N_13099,N_13115);
xnor U13172 (N_13172,N_13004,N_13052);
nor U13173 (N_13173,N_13112,N_13096);
nor U13174 (N_13174,N_13066,N_13001);
and U13175 (N_13175,N_13003,N_13036);
or U13176 (N_13176,N_13028,N_13057);
and U13177 (N_13177,N_13031,N_13106);
xnor U13178 (N_13178,N_13026,N_13025);
and U13179 (N_13179,N_13008,N_13037);
and U13180 (N_13180,N_13082,N_13050);
or U13181 (N_13181,N_13098,N_13081);
xnor U13182 (N_13182,N_13097,N_13121);
nand U13183 (N_13183,N_13116,N_13093);
xor U13184 (N_13184,N_13059,N_13103);
xnor U13185 (N_13185,N_13013,N_13072);
nor U13186 (N_13186,N_13035,N_13067);
xnor U13187 (N_13187,N_13009,N_13066);
and U13188 (N_13188,N_13044,N_13027);
xor U13189 (N_13189,N_13028,N_13043);
nor U13190 (N_13190,N_13117,N_13024);
or U13191 (N_13191,N_13071,N_13031);
xor U13192 (N_13192,N_13032,N_13094);
xnor U13193 (N_13193,N_13046,N_13098);
and U13194 (N_13194,N_13020,N_13017);
nand U13195 (N_13195,N_13042,N_13123);
or U13196 (N_13196,N_13084,N_13074);
nand U13197 (N_13197,N_13006,N_13121);
xor U13198 (N_13198,N_13116,N_13020);
nor U13199 (N_13199,N_13065,N_13071);
xnor U13200 (N_13200,N_13092,N_13097);
or U13201 (N_13201,N_13089,N_13008);
xor U13202 (N_13202,N_13074,N_13039);
nand U13203 (N_13203,N_13095,N_13079);
nor U13204 (N_13204,N_13101,N_13070);
and U13205 (N_13205,N_13064,N_13103);
nor U13206 (N_13206,N_13114,N_13073);
and U13207 (N_13207,N_13106,N_13078);
and U13208 (N_13208,N_13059,N_13053);
nand U13209 (N_13209,N_13106,N_13117);
and U13210 (N_13210,N_13080,N_13010);
or U13211 (N_13211,N_13063,N_13000);
nand U13212 (N_13212,N_13100,N_13074);
or U13213 (N_13213,N_13019,N_13092);
xor U13214 (N_13214,N_13073,N_13048);
xnor U13215 (N_13215,N_13000,N_13093);
or U13216 (N_13216,N_13094,N_13000);
nor U13217 (N_13217,N_13029,N_13024);
xor U13218 (N_13218,N_13080,N_13111);
nand U13219 (N_13219,N_13047,N_13108);
and U13220 (N_13220,N_13056,N_13039);
or U13221 (N_13221,N_13044,N_13101);
nor U13222 (N_13222,N_13054,N_13108);
xor U13223 (N_13223,N_13106,N_13013);
nor U13224 (N_13224,N_13077,N_13033);
and U13225 (N_13225,N_13015,N_13075);
nand U13226 (N_13226,N_13067,N_13010);
nand U13227 (N_13227,N_13058,N_13100);
xor U13228 (N_13228,N_13105,N_13114);
and U13229 (N_13229,N_13088,N_13119);
xnor U13230 (N_13230,N_13050,N_13119);
nand U13231 (N_13231,N_13102,N_13072);
or U13232 (N_13232,N_13121,N_13068);
and U13233 (N_13233,N_13005,N_13042);
and U13234 (N_13234,N_13038,N_13081);
xnor U13235 (N_13235,N_13010,N_13070);
nand U13236 (N_13236,N_13020,N_13070);
or U13237 (N_13237,N_13001,N_13028);
or U13238 (N_13238,N_13029,N_13110);
and U13239 (N_13239,N_13000,N_13066);
xor U13240 (N_13240,N_13001,N_13083);
or U13241 (N_13241,N_13077,N_13108);
nand U13242 (N_13242,N_13086,N_13065);
nor U13243 (N_13243,N_13042,N_13100);
xor U13244 (N_13244,N_13054,N_13120);
nand U13245 (N_13245,N_13038,N_13073);
and U13246 (N_13246,N_13037,N_13062);
xor U13247 (N_13247,N_13046,N_13034);
nor U13248 (N_13248,N_13073,N_13087);
nand U13249 (N_13249,N_13003,N_13077);
or U13250 (N_13250,N_13182,N_13152);
nand U13251 (N_13251,N_13212,N_13213);
nand U13252 (N_13252,N_13181,N_13136);
nand U13253 (N_13253,N_13126,N_13241);
nand U13254 (N_13254,N_13141,N_13155);
nor U13255 (N_13255,N_13164,N_13157);
and U13256 (N_13256,N_13166,N_13177);
or U13257 (N_13257,N_13151,N_13145);
xnor U13258 (N_13258,N_13154,N_13185);
xor U13259 (N_13259,N_13129,N_13156);
nand U13260 (N_13260,N_13134,N_13147);
xor U13261 (N_13261,N_13191,N_13178);
xnor U13262 (N_13262,N_13190,N_13195);
or U13263 (N_13263,N_13243,N_13173);
nor U13264 (N_13264,N_13209,N_13172);
or U13265 (N_13265,N_13219,N_13138);
nor U13266 (N_13266,N_13174,N_13169);
nand U13267 (N_13267,N_13218,N_13170);
xor U13268 (N_13268,N_13208,N_13148);
nor U13269 (N_13269,N_13167,N_13226);
nor U13270 (N_13270,N_13201,N_13240);
nor U13271 (N_13271,N_13228,N_13140);
nor U13272 (N_13272,N_13131,N_13242);
nor U13273 (N_13273,N_13222,N_13133);
nor U13274 (N_13274,N_13239,N_13128);
nand U13275 (N_13275,N_13130,N_13163);
xnor U13276 (N_13276,N_13238,N_13162);
nor U13277 (N_13277,N_13229,N_13184);
nor U13278 (N_13278,N_13203,N_13143);
xor U13279 (N_13279,N_13180,N_13168);
or U13280 (N_13280,N_13230,N_13206);
xnor U13281 (N_13281,N_13245,N_13231);
nand U13282 (N_13282,N_13246,N_13189);
nor U13283 (N_13283,N_13199,N_13144);
or U13284 (N_13284,N_13192,N_13204);
nand U13285 (N_13285,N_13216,N_13153);
and U13286 (N_13286,N_13223,N_13176);
nand U13287 (N_13287,N_13150,N_13217);
and U13288 (N_13288,N_13220,N_13132);
or U13289 (N_13289,N_13234,N_13249);
or U13290 (N_13290,N_13214,N_13187);
nand U13291 (N_13291,N_13202,N_13188);
nor U13292 (N_13292,N_13193,N_13227);
nand U13293 (N_13293,N_13139,N_13232);
nor U13294 (N_13294,N_13135,N_13142);
or U13295 (N_13295,N_13194,N_13159);
nand U13296 (N_13296,N_13221,N_13196);
nand U13297 (N_13297,N_13127,N_13247);
xnor U13298 (N_13298,N_13137,N_13186);
nand U13299 (N_13299,N_13183,N_13205);
or U13300 (N_13300,N_13179,N_13125);
nor U13301 (N_13301,N_13244,N_13149);
xnor U13302 (N_13302,N_13158,N_13233);
xnor U13303 (N_13303,N_13207,N_13165);
nor U13304 (N_13304,N_13225,N_13175);
nand U13305 (N_13305,N_13160,N_13235);
nor U13306 (N_13306,N_13210,N_13211);
nand U13307 (N_13307,N_13200,N_13198);
xnor U13308 (N_13308,N_13197,N_13161);
xnor U13309 (N_13309,N_13237,N_13236);
nand U13310 (N_13310,N_13171,N_13215);
nor U13311 (N_13311,N_13146,N_13248);
xor U13312 (N_13312,N_13224,N_13203);
or U13313 (N_13313,N_13230,N_13171);
nand U13314 (N_13314,N_13154,N_13207);
and U13315 (N_13315,N_13190,N_13159);
or U13316 (N_13316,N_13183,N_13190);
nand U13317 (N_13317,N_13174,N_13222);
nor U13318 (N_13318,N_13164,N_13181);
nand U13319 (N_13319,N_13226,N_13195);
or U13320 (N_13320,N_13154,N_13198);
nand U13321 (N_13321,N_13222,N_13216);
nand U13322 (N_13322,N_13192,N_13139);
xnor U13323 (N_13323,N_13156,N_13224);
nor U13324 (N_13324,N_13242,N_13163);
nor U13325 (N_13325,N_13147,N_13242);
xor U13326 (N_13326,N_13238,N_13233);
or U13327 (N_13327,N_13189,N_13223);
nor U13328 (N_13328,N_13204,N_13165);
nor U13329 (N_13329,N_13194,N_13224);
xor U13330 (N_13330,N_13206,N_13234);
or U13331 (N_13331,N_13144,N_13171);
or U13332 (N_13332,N_13153,N_13205);
or U13333 (N_13333,N_13135,N_13126);
nor U13334 (N_13334,N_13208,N_13170);
and U13335 (N_13335,N_13221,N_13142);
and U13336 (N_13336,N_13215,N_13186);
nand U13337 (N_13337,N_13231,N_13203);
and U13338 (N_13338,N_13140,N_13156);
and U13339 (N_13339,N_13222,N_13163);
nand U13340 (N_13340,N_13181,N_13209);
or U13341 (N_13341,N_13221,N_13235);
and U13342 (N_13342,N_13198,N_13162);
and U13343 (N_13343,N_13219,N_13125);
or U13344 (N_13344,N_13209,N_13239);
nor U13345 (N_13345,N_13193,N_13236);
or U13346 (N_13346,N_13202,N_13128);
xor U13347 (N_13347,N_13243,N_13198);
nor U13348 (N_13348,N_13200,N_13176);
and U13349 (N_13349,N_13246,N_13249);
or U13350 (N_13350,N_13182,N_13212);
or U13351 (N_13351,N_13230,N_13198);
or U13352 (N_13352,N_13174,N_13226);
xnor U13353 (N_13353,N_13184,N_13134);
xor U13354 (N_13354,N_13150,N_13126);
nor U13355 (N_13355,N_13154,N_13178);
nor U13356 (N_13356,N_13137,N_13152);
nand U13357 (N_13357,N_13141,N_13199);
nor U13358 (N_13358,N_13157,N_13165);
and U13359 (N_13359,N_13128,N_13248);
xor U13360 (N_13360,N_13216,N_13172);
and U13361 (N_13361,N_13199,N_13185);
nor U13362 (N_13362,N_13130,N_13147);
or U13363 (N_13363,N_13245,N_13243);
xnor U13364 (N_13364,N_13184,N_13196);
or U13365 (N_13365,N_13248,N_13221);
xor U13366 (N_13366,N_13247,N_13246);
or U13367 (N_13367,N_13214,N_13177);
and U13368 (N_13368,N_13226,N_13168);
xnor U13369 (N_13369,N_13164,N_13188);
nor U13370 (N_13370,N_13218,N_13175);
nand U13371 (N_13371,N_13182,N_13143);
and U13372 (N_13372,N_13187,N_13155);
nor U13373 (N_13373,N_13228,N_13178);
nand U13374 (N_13374,N_13207,N_13225);
xnor U13375 (N_13375,N_13295,N_13284);
nor U13376 (N_13376,N_13268,N_13309);
nand U13377 (N_13377,N_13348,N_13275);
and U13378 (N_13378,N_13285,N_13270);
and U13379 (N_13379,N_13308,N_13281);
nor U13380 (N_13380,N_13333,N_13304);
or U13381 (N_13381,N_13360,N_13367);
and U13382 (N_13382,N_13278,N_13356);
nor U13383 (N_13383,N_13326,N_13297);
or U13384 (N_13384,N_13324,N_13250);
and U13385 (N_13385,N_13263,N_13343);
or U13386 (N_13386,N_13274,N_13260);
xor U13387 (N_13387,N_13305,N_13266);
and U13388 (N_13388,N_13342,N_13323);
xor U13389 (N_13389,N_13282,N_13344);
nor U13390 (N_13390,N_13346,N_13277);
nand U13391 (N_13391,N_13338,N_13369);
and U13392 (N_13392,N_13265,N_13253);
nand U13393 (N_13393,N_13276,N_13372);
xor U13394 (N_13394,N_13289,N_13349);
or U13395 (N_13395,N_13310,N_13279);
xnor U13396 (N_13396,N_13320,N_13303);
xnor U13397 (N_13397,N_13273,N_13302);
or U13398 (N_13398,N_13359,N_13292);
xnor U13399 (N_13399,N_13353,N_13350);
or U13400 (N_13400,N_13298,N_13255);
nor U13401 (N_13401,N_13325,N_13311);
nor U13402 (N_13402,N_13294,N_13341);
and U13403 (N_13403,N_13252,N_13366);
or U13404 (N_13404,N_13269,N_13327);
nand U13405 (N_13405,N_13261,N_13352);
nor U13406 (N_13406,N_13331,N_13317);
and U13407 (N_13407,N_13370,N_13307);
and U13408 (N_13408,N_13336,N_13354);
or U13409 (N_13409,N_13328,N_13259);
and U13410 (N_13410,N_13365,N_13287);
and U13411 (N_13411,N_13288,N_13293);
nor U13412 (N_13412,N_13335,N_13371);
or U13413 (N_13413,N_13364,N_13363);
and U13414 (N_13414,N_13339,N_13322);
nand U13415 (N_13415,N_13361,N_13267);
nand U13416 (N_13416,N_13262,N_13306);
and U13417 (N_13417,N_13301,N_13351);
xnor U13418 (N_13418,N_13258,N_13337);
nand U13419 (N_13419,N_13347,N_13264);
nand U13420 (N_13420,N_13362,N_13280);
xnor U13421 (N_13421,N_13312,N_13286);
nor U13422 (N_13422,N_13321,N_13345);
and U13423 (N_13423,N_13313,N_13315);
nand U13424 (N_13424,N_13358,N_13283);
xor U13425 (N_13425,N_13340,N_13272);
or U13426 (N_13426,N_13290,N_13271);
and U13427 (N_13427,N_13318,N_13254);
xor U13428 (N_13428,N_13334,N_13296);
xor U13429 (N_13429,N_13374,N_13257);
or U13430 (N_13430,N_13314,N_13256);
nand U13431 (N_13431,N_13291,N_13299);
nor U13432 (N_13432,N_13357,N_13332);
and U13433 (N_13433,N_13251,N_13368);
or U13434 (N_13434,N_13319,N_13316);
nand U13435 (N_13435,N_13329,N_13300);
or U13436 (N_13436,N_13355,N_13373);
and U13437 (N_13437,N_13330,N_13313);
or U13438 (N_13438,N_13342,N_13264);
or U13439 (N_13439,N_13360,N_13264);
or U13440 (N_13440,N_13298,N_13332);
and U13441 (N_13441,N_13328,N_13334);
and U13442 (N_13442,N_13281,N_13252);
or U13443 (N_13443,N_13362,N_13295);
xor U13444 (N_13444,N_13285,N_13363);
nand U13445 (N_13445,N_13284,N_13359);
xor U13446 (N_13446,N_13349,N_13352);
xnor U13447 (N_13447,N_13347,N_13337);
nand U13448 (N_13448,N_13319,N_13274);
nor U13449 (N_13449,N_13311,N_13359);
nor U13450 (N_13450,N_13347,N_13295);
nor U13451 (N_13451,N_13363,N_13329);
or U13452 (N_13452,N_13301,N_13326);
xnor U13453 (N_13453,N_13258,N_13344);
and U13454 (N_13454,N_13292,N_13310);
nand U13455 (N_13455,N_13363,N_13295);
or U13456 (N_13456,N_13374,N_13290);
and U13457 (N_13457,N_13267,N_13367);
or U13458 (N_13458,N_13298,N_13352);
nand U13459 (N_13459,N_13253,N_13267);
and U13460 (N_13460,N_13266,N_13372);
xnor U13461 (N_13461,N_13280,N_13281);
xnor U13462 (N_13462,N_13297,N_13274);
xnor U13463 (N_13463,N_13277,N_13316);
xnor U13464 (N_13464,N_13326,N_13352);
or U13465 (N_13465,N_13312,N_13304);
and U13466 (N_13466,N_13257,N_13337);
and U13467 (N_13467,N_13298,N_13275);
xor U13468 (N_13468,N_13351,N_13308);
and U13469 (N_13469,N_13298,N_13301);
or U13470 (N_13470,N_13371,N_13302);
xor U13471 (N_13471,N_13261,N_13299);
nand U13472 (N_13472,N_13371,N_13309);
nor U13473 (N_13473,N_13277,N_13321);
or U13474 (N_13474,N_13340,N_13330);
nand U13475 (N_13475,N_13331,N_13347);
or U13476 (N_13476,N_13338,N_13286);
and U13477 (N_13477,N_13344,N_13260);
nor U13478 (N_13478,N_13324,N_13265);
and U13479 (N_13479,N_13344,N_13250);
nand U13480 (N_13480,N_13357,N_13316);
and U13481 (N_13481,N_13372,N_13286);
nand U13482 (N_13482,N_13351,N_13291);
nor U13483 (N_13483,N_13299,N_13251);
nand U13484 (N_13484,N_13284,N_13285);
nand U13485 (N_13485,N_13269,N_13297);
nor U13486 (N_13486,N_13323,N_13348);
nand U13487 (N_13487,N_13346,N_13260);
xnor U13488 (N_13488,N_13341,N_13252);
nand U13489 (N_13489,N_13357,N_13326);
and U13490 (N_13490,N_13263,N_13279);
and U13491 (N_13491,N_13250,N_13308);
nand U13492 (N_13492,N_13367,N_13310);
nor U13493 (N_13493,N_13283,N_13343);
and U13494 (N_13494,N_13328,N_13349);
or U13495 (N_13495,N_13319,N_13370);
xnor U13496 (N_13496,N_13312,N_13278);
nor U13497 (N_13497,N_13251,N_13334);
and U13498 (N_13498,N_13251,N_13327);
xnor U13499 (N_13499,N_13279,N_13300);
xor U13500 (N_13500,N_13449,N_13394);
and U13501 (N_13501,N_13477,N_13413);
nor U13502 (N_13502,N_13414,N_13464);
nand U13503 (N_13503,N_13425,N_13428);
and U13504 (N_13504,N_13388,N_13462);
or U13505 (N_13505,N_13377,N_13441);
and U13506 (N_13506,N_13438,N_13384);
xor U13507 (N_13507,N_13440,N_13451);
and U13508 (N_13508,N_13475,N_13397);
xnor U13509 (N_13509,N_13390,N_13379);
or U13510 (N_13510,N_13403,N_13442);
xnor U13511 (N_13511,N_13426,N_13433);
nor U13512 (N_13512,N_13454,N_13380);
or U13513 (N_13513,N_13412,N_13448);
xnor U13514 (N_13514,N_13495,N_13445);
nand U13515 (N_13515,N_13490,N_13427);
and U13516 (N_13516,N_13436,N_13409);
and U13517 (N_13517,N_13431,N_13443);
xor U13518 (N_13518,N_13457,N_13437);
nor U13519 (N_13519,N_13396,N_13439);
xor U13520 (N_13520,N_13498,N_13494);
xnor U13521 (N_13521,N_13472,N_13401);
nand U13522 (N_13522,N_13411,N_13417);
or U13523 (N_13523,N_13455,N_13382);
or U13524 (N_13524,N_13468,N_13398);
and U13525 (N_13525,N_13410,N_13402);
and U13526 (N_13526,N_13444,N_13435);
nor U13527 (N_13527,N_13421,N_13432);
xor U13528 (N_13528,N_13453,N_13491);
or U13529 (N_13529,N_13466,N_13389);
nand U13530 (N_13530,N_13486,N_13470);
or U13531 (N_13531,N_13473,N_13420);
nor U13532 (N_13532,N_13383,N_13408);
nand U13533 (N_13533,N_13430,N_13456);
xnor U13534 (N_13534,N_13497,N_13476);
xor U13535 (N_13535,N_13469,N_13423);
and U13536 (N_13536,N_13493,N_13458);
nor U13537 (N_13537,N_13496,N_13418);
or U13538 (N_13538,N_13407,N_13460);
or U13539 (N_13539,N_13481,N_13404);
nand U13540 (N_13540,N_13483,N_13422);
nand U13541 (N_13541,N_13465,N_13461);
xnor U13542 (N_13542,N_13387,N_13447);
nand U13543 (N_13543,N_13499,N_13446);
xnor U13544 (N_13544,N_13406,N_13395);
nand U13545 (N_13545,N_13376,N_13487);
nand U13546 (N_13546,N_13463,N_13392);
and U13547 (N_13547,N_13400,N_13429);
or U13548 (N_13548,N_13488,N_13419);
xor U13549 (N_13549,N_13450,N_13482);
nand U13550 (N_13550,N_13385,N_13467);
nand U13551 (N_13551,N_13415,N_13399);
nand U13552 (N_13552,N_13492,N_13391);
xor U13553 (N_13553,N_13424,N_13459);
or U13554 (N_13554,N_13434,N_13375);
nor U13555 (N_13555,N_13471,N_13378);
xnor U13556 (N_13556,N_13405,N_13478);
or U13557 (N_13557,N_13393,N_13474);
nor U13558 (N_13558,N_13484,N_13479);
xor U13559 (N_13559,N_13480,N_13485);
xnor U13560 (N_13560,N_13416,N_13489);
and U13561 (N_13561,N_13386,N_13452);
nand U13562 (N_13562,N_13381,N_13489);
and U13563 (N_13563,N_13460,N_13479);
xnor U13564 (N_13564,N_13400,N_13499);
xor U13565 (N_13565,N_13382,N_13435);
xnor U13566 (N_13566,N_13410,N_13409);
xnor U13567 (N_13567,N_13440,N_13398);
or U13568 (N_13568,N_13428,N_13410);
xnor U13569 (N_13569,N_13466,N_13490);
or U13570 (N_13570,N_13443,N_13418);
and U13571 (N_13571,N_13386,N_13458);
and U13572 (N_13572,N_13494,N_13396);
nor U13573 (N_13573,N_13430,N_13471);
nand U13574 (N_13574,N_13413,N_13394);
xor U13575 (N_13575,N_13379,N_13487);
nor U13576 (N_13576,N_13494,N_13436);
or U13577 (N_13577,N_13439,N_13487);
and U13578 (N_13578,N_13433,N_13385);
xor U13579 (N_13579,N_13458,N_13439);
nand U13580 (N_13580,N_13431,N_13393);
nor U13581 (N_13581,N_13405,N_13434);
and U13582 (N_13582,N_13383,N_13417);
nand U13583 (N_13583,N_13398,N_13394);
nor U13584 (N_13584,N_13497,N_13392);
and U13585 (N_13585,N_13479,N_13433);
nor U13586 (N_13586,N_13450,N_13479);
and U13587 (N_13587,N_13476,N_13385);
nand U13588 (N_13588,N_13392,N_13435);
and U13589 (N_13589,N_13479,N_13426);
or U13590 (N_13590,N_13412,N_13473);
xnor U13591 (N_13591,N_13375,N_13494);
or U13592 (N_13592,N_13464,N_13495);
nand U13593 (N_13593,N_13383,N_13495);
nand U13594 (N_13594,N_13395,N_13425);
nand U13595 (N_13595,N_13442,N_13409);
and U13596 (N_13596,N_13404,N_13482);
nor U13597 (N_13597,N_13461,N_13432);
nor U13598 (N_13598,N_13415,N_13482);
nor U13599 (N_13599,N_13390,N_13460);
nor U13600 (N_13600,N_13460,N_13484);
xor U13601 (N_13601,N_13456,N_13453);
or U13602 (N_13602,N_13498,N_13459);
and U13603 (N_13603,N_13461,N_13437);
nor U13604 (N_13604,N_13497,N_13401);
nor U13605 (N_13605,N_13391,N_13463);
nand U13606 (N_13606,N_13417,N_13450);
nand U13607 (N_13607,N_13376,N_13390);
nand U13608 (N_13608,N_13396,N_13409);
nor U13609 (N_13609,N_13411,N_13489);
and U13610 (N_13610,N_13446,N_13381);
nand U13611 (N_13611,N_13464,N_13455);
and U13612 (N_13612,N_13428,N_13395);
and U13613 (N_13613,N_13416,N_13449);
nand U13614 (N_13614,N_13393,N_13483);
or U13615 (N_13615,N_13429,N_13487);
or U13616 (N_13616,N_13476,N_13445);
nand U13617 (N_13617,N_13444,N_13402);
xnor U13618 (N_13618,N_13492,N_13392);
or U13619 (N_13619,N_13418,N_13393);
and U13620 (N_13620,N_13487,N_13448);
nor U13621 (N_13621,N_13491,N_13427);
nor U13622 (N_13622,N_13454,N_13439);
xnor U13623 (N_13623,N_13420,N_13461);
and U13624 (N_13624,N_13495,N_13454);
nor U13625 (N_13625,N_13514,N_13600);
or U13626 (N_13626,N_13585,N_13530);
xor U13627 (N_13627,N_13522,N_13584);
xnor U13628 (N_13628,N_13542,N_13617);
xnor U13629 (N_13629,N_13565,N_13623);
xor U13630 (N_13630,N_13572,N_13539);
nand U13631 (N_13631,N_13544,N_13557);
nor U13632 (N_13632,N_13541,N_13543);
and U13633 (N_13633,N_13540,N_13521);
nand U13634 (N_13634,N_13501,N_13520);
xnor U13635 (N_13635,N_13576,N_13590);
xnor U13636 (N_13636,N_13560,N_13608);
nand U13637 (N_13637,N_13609,N_13620);
or U13638 (N_13638,N_13561,N_13523);
and U13639 (N_13639,N_13622,N_13519);
nor U13640 (N_13640,N_13556,N_13594);
nor U13641 (N_13641,N_13583,N_13554);
nand U13642 (N_13642,N_13563,N_13533);
xor U13643 (N_13643,N_13507,N_13589);
or U13644 (N_13644,N_13569,N_13527);
xor U13645 (N_13645,N_13612,N_13578);
or U13646 (N_13646,N_13615,N_13528);
or U13647 (N_13647,N_13619,N_13599);
nand U13648 (N_13648,N_13537,N_13579);
and U13649 (N_13649,N_13515,N_13580);
xor U13650 (N_13650,N_13564,N_13506);
xor U13651 (N_13651,N_13503,N_13593);
nand U13652 (N_13652,N_13545,N_13509);
or U13653 (N_13653,N_13577,N_13508);
or U13654 (N_13654,N_13621,N_13513);
nand U13655 (N_13655,N_13536,N_13595);
nand U13656 (N_13656,N_13552,N_13575);
xnor U13657 (N_13657,N_13548,N_13558);
or U13658 (N_13658,N_13547,N_13551);
and U13659 (N_13659,N_13525,N_13610);
xnor U13660 (N_13660,N_13526,N_13587);
xor U13661 (N_13661,N_13511,N_13553);
nand U13662 (N_13662,N_13562,N_13532);
and U13663 (N_13663,N_13567,N_13516);
and U13664 (N_13664,N_13592,N_13510);
nor U13665 (N_13665,N_13574,N_13524);
xnor U13666 (N_13666,N_13598,N_13624);
nor U13667 (N_13667,N_13604,N_13611);
nand U13668 (N_13668,N_13555,N_13568);
or U13669 (N_13669,N_13573,N_13616);
xor U13670 (N_13670,N_13588,N_13618);
nor U13671 (N_13671,N_13550,N_13546);
or U13672 (N_13672,N_13591,N_13613);
nand U13673 (N_13673,N_13559,N_13602);
and U13674 (N_13674,N_13606,N_13512);
nand U13675 (N_13675,N_13534,N_13517);
nor U13676 (N_13676,N_13549,N_13607);
nand U13677 (N_13677,N_13518,N_13505);
xor U13678 (N_13678,N_13535,N_13586);
and U13679 (N_13679,N_13601,N_13570);
and U13680 (N_13680,N_13582,N_13596);
xnor U13681 (N_13681,N_13603,N_13502);
or U13682 (N_13682,N_13566,N_13571);
xor U13683 (N_13683,N_13605,N_13538);
and U13684 (N_13684,N_13597,N_13614);
or U13685 (N_13685,N_13531,N_13581);
nor U13686 (N_13686,N_13504,N_13500);
nor U13687 (N_13687,N_13529,N_13615);
nand U13688 (N_13688,N_13624,N_13617);
and U13689 (N_13689,N_13568,N_13524);
and U13690 (N_13690,N_13613,N_13589);
or U13691 (N_13691,N_13616,N_13507);
xnor U13692 (N_13692,N_13616,N_13559);
nand U13693 (N_13693,N_13616,N_13572);
nor U13694 (N_13694,N_13615,N_13521);
or U13695 (N_13695,N_13618,N_13560);
or U13696 (N_13696,N_13568,N_13603);
and U13697 (N_13697,N_13581,N_13522);
nand U13698 (N_13698,N_13577,N_13602);
and U13699 (N_13699,N_13613,N_13585);
or U13700 (N_13700,N_13525,N_13566);
nand U13701 (N_13701,N_13610,N_13599);
nor U13702 (N_13702,N_13540,N_13608);
nor U13703 (N_13703,N_13552,N_13534);
xnor U13704 (N_13704,N_13591,N_13601);
xor U13705 (N_13705,N_13539,N_13620);
nor U13706 (N_13706,N_13586,N_13543);
or U13707 (N_13707,N_13558,N_13561);
or U13708 (N_13708,N_13617,N_13598);
and U13709 (N_13709,N_13582,N_13618);
nand U13710 (N_13710,N_13569,N_13516);
xnor U13711 (N_13711,N_13501,N_13617);
xnor U13712 (N_13712,N_13605,N_13594);
nor U13713 (N_13713,N_13611,N_13568);
and U13714 (N_13714,N_13526,N_13562);
and U13715 (N_13715,N_13604,N_13520);
xor U13716 (N_13716,N_13574,N_13613);
and U13717 (N_13717,N_13564,N_13592);
or U13718 (N_13718,N_13529,N_13590);
and U13719 (N_13719,N_13586,N_13575);
xnor U13720 (N_13720,N_13576,N_13558);
nor U13721 (N_13721,N_13560,N_13573);
nor U13722 (N_13722,N_13578,N_13556);
xor U13723 (N_13723,N_13583,N_13601);
nor U13724 (N_13724,N_13574,N_13600);
or U13725 (N_13725,N_13607,N_13618);
nor U13726 (N_13726,N_13609,N_13502);
or U13727 (N_13727,N_13570,N_13553);
or U13728 (N_13728,N_13557,N_13610);
and U13729 (N_13729,N_13617,N_13513);
or U13730 (N_13730,N_13594,N_13507);
and U13731 (N_13731,N_13551,N_13505);
or U13732 (N_13732,N_13506,N_13530);
nand U13733 (N_13733,N_13586,N_13612);
and U13734 (N_13734,N_13617,N_13522);
or U13735 (N_13735,N_13504,N_13624);
nor U13736 (N_13736,N_13525,N_13533);
nor U13737 (N_13737,N_13565,N_13505);
and U13738 (N_13738,N_13576,N_13579);
xor U13739 (N_13739,N_13601,N_13612);
nor U13740 (N_13740,N_13557,N_13611);
nand U13741 (N_13741,N_13506,N_13568);
nor U13742 (N_13742,N_13505,N_13568);
or U13743 (N_13743,N_13531,N_13543);
nand U13744 (N_13744,N_13548,N_13571);
nor U13745 (N_13745,N_13567,N_13535);
xor U13746 (N_13746,N_13586,N_13592);
xor U13747 (N_13747,N_13615,N_13580);
or U13748 (N_13748,N_13605,N_13568);
nor U13749 (N_13749,N_13596,N_13624);
and U13750 (N_13750,N_13728,N_13686);
xnor U13751 (N_13751,N_13733,N_13747);
xnor U13752 (N_13752,N_13690,N_13681);
nand U13753 (N_13753,N_13691,N_13678);
and U13754 (N_13754,N_13668,N_13742);
xor U13755 (N_13755,N_13727,N_13656);
xnor U13756 (N_13756,N_13630,N_13674);
and U13757 (N_13757,N_13726,N_13694);
nor U13758 (N_13758,N_13683,N_13697);
nand U13759 (N_13759,N_13663,N_13721);
nor U13760 (N_13760,N_13722,N_13698);
and U13761 (N_13761,N_13659,N_13632);
nor U13762 (N_13762,N_13640,N_13643);
xnor U13763 (N_13763,N_13702,N_13736);
nor U13764 (N_13764,N_13741,N_13700);
or U13765 (N_13765,N_13705,N_13744);
nand U13766 (N_13766,N_13735,N_13650);
or U13767 (N_13767,N_13713,N_13696);
nand U13768 (N_13768,N_13706,N_13679);
nor U13769 (N_13769,N_13749,N_13636);
and U13770 (N_13770,N_13671,N_13664);
nand U13771 (N_13771,N_13718,N_13685);
nor U13772 (N_13772,N_13657,N_13672);
xnor U13773 (N_13773,N_13661,N_13711);
or U13774 (N_13774,N_13626,N_13653);
or U13775 (N_13775,N_13689,N_13652);
xor U13776 (N_13776,N_13645,N_13748);
nor U13777 (N_13777,N_13707,N_13745);
nand U13778 (N_13778,N_13720,N_13688);
or U13779 (N_13779,N_13731,N_13699);
nand U13780 (N_13780,N_13716,N_13725);
xnor U13781 (N_13781,N_13692,N_13660);
nand U13782 (N_13782,N_13641,N_13627);
xnor U13783 (N_13783,N_13740,N_13649);
nor U13784 (N_13784,N_13644,N_13684);
and U13785 (N_13785,N_13631,N_13695);
nor U13786 (N_13786,N_13655,N_13732);
nor U13787 (N_13787,N_13719,N_13670);
xnor U13788 (N_13788,N_13701,N_13647);
nor U13789 (N_13789,N_13665,N_13738);
and U13790 (N_13790,N_13666,N_13669);
nor U13791 (N_13791,N_13625,N_13737);
xor U13792 (N_13792,N_13743,N_13673);
nor U13793 (N_13793,N_13628,N_13675);
and U13794 (N_13794,N_13717,N_13677);
and U13795 (N_13795,N_13646,N_13676);
xor U13796 (N_13796,N_13680,N_13739);
and U13797 (N_13797,N_13637,N_13704);
or U13798 (N_13798,N_13635,N_13634);
xnor U13799 (N_13799,N_13724,N_13642);
and U13800 (N_13800,N_13667,N_13709);
xor U13801 (N_13801,N_13639,N_13710);
and U13802 (N_13802,N_13662,N_13658);
xnor U13803 (N_13803,N_13633,N_13682);
or U13804 (N_13804,N_13648,N_13734);
xor U13805 (N_13805,N_13651,N_13746);
and U13806 (N_13806,N_13703,N_13715);
nor U13807 (N_13807,N_13714,N_13730);
xnor U13808 (N_13808,N_13708,N_13723);
xnor U13809 (N_13809,N_13693,N_13629);
and U13810 (N_13810,N_13687,N_13729);
nand U13811 (N_13811,N_13638,N_13712);
nor U13812 (N_13812,N_13654,N_13671);
xor U13813 (N_13813,N_13665,N_13684);
xor U13814 (N_13814,N_13672,N_13681);
or U13815 (N_13815,N_13654,N_13641);
or U13816 (N_13816,N_13718,N_13719);
nor U13817 (N_13817,N_13735,N_13670);
and U13818 (N_13818,N_13719,N_13686);
and U13819 (N_13819,N_13647,N_13664);
or U13820 (N_13820,N_13629,N_13682);
nand U13821 (N_13821,N_13716,N_13720);
nand U13822 (N_13822,N_13693,N_13745);
and U13823 (N_13823,N_13636,N_13632);
or U13824 (N_13824,N_13732,N_13685);
xnor U13825 (N_13825,N_13706,N_13715);
or U13826 (N_13826,N_13633,N_13742);
or U13827 (N_13827,N_13671,N_13694);
xnor U13828 (N_13828,N_13732,N_13720);
nor U13829 (N_13829,N_13625,N_13627);
xnor U13830 (N_13830,N_13645,N_13653);
and U13831 (N_13831,N_13636,N_13674);
and U13832 (N_13832,N_13705,N_13628);
xnor U13833 (N_13833,N_13655,N_13688);
nand U13834 (N_13834,N_13736,N_13705);
nor U13835 (N_13835,N_13677,N_13665);
xor U13836 (N_13836,N_13702,N_13710);
and U13837 (N_13837,N_13682,N_13710);
xnor U13838 (N_13838,N_13647,N_13698);
xnor U13839 (N_13839,N_13686,N_13743);
and U13840 (N_13840,N_13662,N_13697);
and U13841 (N_13841,N_13673,N_13645);
xor U13842 (N_13842,N_13716,N_13682);
nand U13843 (N_13843,N_13685,N_13701);
xor U13844 (N_13844,N_13668,N_13663);
nor U13845 (N_13845,N_13693,N_13732);
xor U13846 (N_13846,N_13648,N_13626);
and U13847 (N_13847,N_13634,N_13707);
xnor U13848 (N_13848,N_13729,N_13665);
nor U13849 (N_13849,N_13659,N_13679);
xor U13850 (N_13850,N_13707,N_13688);
and U13851 (N_13851,N_13641,N_13647);
and U13852 (N_13852,N_13742,N_13736);
nand U13853 (N_13853,N_13683,N_13653);
and U13854 (N_13854,N_13741,N_13660);
and U13855 (N_13855,N_13692,N_13735);
xnor U13856 (N_13856,N_13746,N_13678);
xor U13857 (N_13857,N_13739,N_13725);
xor U13858 (N_13858,N_13697,N_13747);
nand U13859 (N_13859,N_13717,N_13638);
and U13860 (N_13860,N_13723,N_13701);
or U13861 (N_13861,N_13633,N_13658);
nor U13862 (N_13862,N_13689,N_13684);
or U13863 (N_13863,N_13657,N_13653);
xor U13864 (N_13864,N_13676,N_13634);
nand U13865 (N_13865,N_13742,N_13630);
or U13866 (N_13866,N_13746,N_13711);
nand U13867 (N_13867,N_13675,N_13705);
and U13868 (N_13868,N_13670,N_13743);
nor U13869 (N_13869,N_13738,N_13692);
nor U13870 (N_13870,N_13708,N_13658);
and U13871 (N_13871,N_13643,N_13683);
nor U13872 (N_13872,N_13708,N_13648);
xnor U13873 (N_13873,N_13682,N_13671);
nor U13874 (N_13874,N_13686,N_13631);
or U13875 (N_13875,N_13815,N_13854);
xnor U13876 (N_13876,N_13760,N_13782);
xor U13877 (N_13877,N_13752,N_13751);
nor U13878 (N_13878,N_13852,N_13857);
xor U13879 (N_13879,N_13853,N_13835);
or U13880 (N_13880,N_13873,N_13803);
xnor U13881 (N_13881,N_13799,N_13781);
and U13882 (N_13882,N_13757,N_13798);
nand U13883 (N_13883,N_13813,N_13778);
nor U13884 (N_13884,N_13833,N_13753);
nor U13885 (N_13885,N_13824,N_13776);
nand U13886 (N_13886,N_13823,N_13868);
and U13887 (N_13887,N_13805,N_13827);
or U13888 (N_13888,N_13844,N_13790);
xnor U13889 (N_13889,N_13860,N_13851);
and U13890 (N_13890,N_13838,N_13750);
or U13891 (N_13891,N_13842,N_13763);
nand U13892 (N_13892,N_13874,N_13819);
nor U13893 (N_13893,N_13786,N_13820);
nand U13894 (N_13894,N_13765,N_13867);
nor U13895 (N_13895,N_13758,N_13858);
nor U13896 (N_13896,N_13795,N_13834);
nor U13897 (N_13897,N_13871,N_13843);
nor U13898 (N_13898,N_13869,N_13837);
and U13899 (N_13899,N_13772,N_13780);
and U13900 (N_13900,N_13862,N_13774);
and U13901 (N_13901,N_13850,N_13825);
or U13902 (N_13902,N_13863,N_13811);
and U13903 (N_13903,N_13800,N_13783);
xor U13904 (N_13904,N_13826,N_13859);
or U13905 (N_13905,N_13866,N_13831);
or U13906 (N_13906,N_13787,N_13832);
xnor U13907 (N_13907,N_13804,N_13848);
and U13908 (N_13908,N_13808,N_13789);
nand U13909 (N_13909,N_13773,N_13816);
and U13910 (N_13910,N_13766,N_13796);
nor U13911 (N_13911,N_13788,N_13767);
nand U13912 (N_13912,N_13771,N_13841);
and U13913 (N_13913,N_13797,N_13791);
xor U13914 (N_13914,N_13792,N_13847);
nor U13915 (N_13915,N_13840,N_13755);
nor U13916 (N_13916,N_13775,N_13818);
nand U13917 (N_13917,N_13754,N_13762);
or U13918 (N_13918,N_13809,N_13836);
or U13919 (N_13919,N_13814,N_13865);
and U13920 (N_13920,N_13768,N_13870);
and U13921 (N_13921,N_13830,N_13846);
xnor U13922 (N_13922,N_13761,N_13801);
and U13923 (N_13923,N_13802,N_13828);
xnor U13924 (N_13924,N_13861,N_13810);
nor U13925 (N_13925,N_13821,N_13794);
nor U13926 (N_13926,N_13872,N_13769);
nor U13927 (N_13927,N_13764,N_13849);
and U13928 (N_13928,N_13784,N_13807);
xnor U13929 (N_13929,N_13759,N_13855);
and U13930 (N_13930,N_13779,N_13845);
nand U13931 (N_13931,N_13777,N_13785);
nand U13932 (N_13932,N_13756,N_13812);
nor U13933 (N_13933,N_13839,N_13770);
and U13934 (N_13934,N_13856,N_13806);
nand U13935 (N_13935,N_13793,N_13864);
nand U13936 (N_13936,N_13822,N_13817);
or U13937 (N_13937,N_13829,N_13840);
nor U13938 (N_13938,N_13843,N_13794);
and U13939 (N_13939,N_13793,N_13794);
nand U13940 (N_13940,N_13863,N_13810);
or U13941 (N_13941,N_13821,N_13852);
xnor U13942 (N_13942,N_13768,N_13835);
nor U13943 (N_13943,N_13817,N_13808);
and U13944 (N_13944,N_13826,N_13810);
and U13945 (N_13945,N_13785,N_13831);
or U13946 (N_13946,N_13799,N_13815);
or U13947 (N_13947,N_13766,N_13839);
nor U13948 (N_13948,N_13829,N_13762);
nand U13949 (N_13949,N_13864,N_13802);
and U13950 (N_13950,N_13838,N_13752);
xnor U13951 (N_13951,N_13755,N_13873);
xnor U13952 (N_13952,N_13793,N_13814);
nand U13953 (N_13953,N_13818,N_13829);
nor U13954 (N_13954,N_13868,N_13835);
xor U13955 (N_13955,N_13873,N_13763);
nor U13956 (N_13956,N_13802,N_13773);
xnor U13957 (N_13957,N_13786,N_13787);
nand U13958 (N_13958,N_13807,N_13792);
nand U13959 (N_13959,N_13810,N_13839);
nand U13960 (N_13960,N_13856,N_13802);
nand U13961 (N_13961,N_13801,N_13777);
and U13962 (N_13962,N_13763,N_13778);
xor U13963 (N_13963,N_13840,N_13816);
and U13964 (N_13964,N_13840,N_13861);
nand U13965 (N_13965,N_13753,N_13809);
nand U13966 (N_13966,N_13763,N_13776);
or U13967 (N_13967,N_13860,N_13829);
or U13968 (N_13968,N_13838,N_13780);
and U13969 (N_13969,N_13825,N_13809);
and U13970 (N_13970,N_13799,N_13854);
nor U13971 (N_13971,N_13817,N_13786);
and U13972 (N_13972,N_13806,N_13759);
nor U13973 (N_13973,N_13773,N_13858);
or U13974 (N_13974,N_13812,N_13794);
or U13975 (N_13975,N_13789,N_13859);
and U13976 (N_13976,N_13870,N_13752);
and U13977 (N_13977,N_13766,N_13781);
xor U13978 (N_13978,N_13840,N_13758);
and U13979 (N_13979,N_13771,N_13800);
nand U13980 (N_13980,N_13855,N_13837);
nor U13981 (N_13981,N_13820,N_13752);
and U13982 (N_13982,N_13853,N_13817);
and U13983 (N_13983,N_13812,N_13814);
nor U13984 (N_13984,N_13827,N_13865);
nand U13985 (N_13985,N_13856,N_13852);
nand U13986 (N_13986,N_13802,N_13817);
and U13987 (N_13987,N_13868,N_13798);
nand U13988 (N_13988,N_13829,N_13791);
and U13989 (N_13989,N_13802,N_13764);
xor U13990 (N_13990,N_13778,N_13850);
and U13991 (N_13991,N_13824,N_13832);
or U13992 (N_13992,N_13797,N_13852);
or U13993 (N_13993,N_13758,N_13780);
xor U13994 (N_13994,N_13849,N_13814);
xor U13995 (N_13995,N_13806,N_13847);
and U13996 (N_13996,N_13806,N_13797);
nor U13997 (N_13997,N_13764,N_13858);
and U13998 (N_13998,N_13840,N_13857);
nand U13999 (N_13999,N_13828,N_13846);
nand U14000 (N_14000,N_13989,N_13899);
nand U14001 (N_14001,N_13997,N_13981);
nand U14002 (N_14002,N_13939,N_13935);
and U14003 (N_14003,N_13921,N_13957);
xnor U14004 (N_14004,N_13886,N_13894);
nor U14005 (N_14005,N_13927,N_13902);
nor U14006 (N_14006,N_13909,N_13940);
and U14007 (N_14007,N_13889,N_13922);
nand U14008 (N_14008,N_13919,N_13930);
nand U14009 (N_14009,N_13916,N_13954);
xnor U14010 (N_14010,N_13943,N_13908);
nand U14011 (N_14011,N_13915,N_13906);
xnor U14012 (N_14012,N_13880,N_13882);
and U14013 (N_14013,N_13926,N_13956);
and U14014 (N_14014,N_13877,N_13958);
and U14015 (N_14015,N_13992,N_13875);
and U14016 (N_14016,N_13895,N_13976);
nor U14017 (N_14017,N_13980,N_13897);
xor U14018 (N_14018,N_13962,N_13955);
xnor U14019 (N_14019,N_13912,N_13934);
or U14020 (N_14020,N_13969,N_13931);
and U14021 (N_14021,N_13901,N_13968);
xnor U14022 (N_14022,N_13914,N_13999);
nor U14023 (N_14023,N_13885,N_13900);
or U14024 (N_14024,N_13946,N_13911);
xnor U14025 (N_14025,N_13974,N_13944);
xor U14026 (N_14026,N_13947,N_13887);
xor U14027 (N_14027,N_13892,N_13948);
and U14028 (N_14028,N_13950,N_13971);
nand U14029 (N_14029,N_13984,N_13932);
or U14030 (N_14030,N_13978,N_13959);
nand U14031 (N_14031,N_13993,N_13878);
and U14032 (N_14032,N_13924,N_13928);
nand U14033 (N_14033,N_13991,N_13972);
xnor U14034 (N_14034,N_13942,N_13963);
nor U14035 (N_14035,N_13907,N_13890);
nor U14036 (N_14036,N_13961,N_13913);
and U14037 (N_14037,N_13891,N_13905);
nand U14038 (N_14038,N_13898,N_13888);
nand U14039 (N_14039,N_13937,N_13918);
nor U14040 (N_14040,N_13994,N_13973);
or U14041 (N_14041,N_13986,N_13945);
or U14042 (N_14042,N_13996,N_13938);
nor U14043 (N_14043,N_13929,N_13951);
xnor U14044 (N_14044,N_13941,N_13988);
and U14045 (N_14045,N_13970,N_13903);
or U14046 (N_14046,N_13949,N_13977);
or U14047 (N_14047,N_13982,N_13904);
or U14048 (N_14048,N_13879,N_13893);
nand U14049 (N_14049,N_13990,N_13883);
nor U14050 (N_14050,N_13933,N_13983);
nor U14051 (N_14051,N_13925,N_13923);
or U14052 (N_14052,N_13952,N_13995);
or U14053 (N_14053,N_13964,N_13987);
nand U14054 (N_14054,N_13960,N_13917);
xor U14055 (N_14055,N_13975,N_13910);
nand U14056 (N_14056,N_13979,N_13965);
nand U14057 (N_14057,N_13881,N_13936);
nor U14058 (N_14058,N_13896,N_13966);
nor U14059 (N_14059,N_13967,N_13920);
nand U14060 (N_14060,N_13953,N_13884);
nand U14061 (N_14061,N_13998,N_13985);
xor U14062 (N_14062,N_13876,N_13880);
or U14063 (N_14063,N_13932,N_13970);
nor U14064 (N_14064,N_13887,N_13903);
or U14065 (N_14065,N_13970,N_13960);
nand U14066 (N_14066,N_13951,N_13965);
nand U14067 (N_14067,N_13895,N_13890);
xnor U14068 (N_14068,N_13995,N_13980);
xnor U14069 (N_14069,N_13994,N_13886);
xor U14070 (N_14070,N_13912,N_13977);
and U14071 (N_14071,N_13998,N_13909);
and U14072 (N_14072,N_13957,N_13985);
and U14073 (N_14073,N_13954,N_13875);
nor U14074 (N_14074,N_13944,N_13943);
nand U14075 (N_14075,N_13963,N_13984);
xor U14076 (N_14076,N_13887,N_13913);
or U14077 (N_14077,N_13942,N_13978);
xor U14078 (N_14078,N_13881,N_13993);
nand U14079 (N_14079,N_13938,N_13897);
nand U14080 (N_14080,N_13885,N_13904);
nand U14081 (N_14081,N_13937,N_13912);
xnor U14082 (N_14082,N_13926,N_13876);
xnor U14083 (N_14083,N_13992,N_13883);
or U14084 (N_14084,N_13971,N_13991);
and U14085 (N_14085,N_13974,N_13878);
nor U14086 (N_14086,N_13986,N_13919);
xnor U14087 (N_14087,N_13976,N_13941);
xor U14088 (N_14088,N_13956,N_13948);
or U14089 (N_14089,N_13922,N_13947);
and U14090 (N_14090,N_13934,N_13937);
and U14091 (N_14091,N_13976,N_13999);
nor U14092 (N_14092,N_13926,N_13877);
and U14093 (N_14093,N_13968,N_13934);
and U14094 (N_14094,N_13913,N_13919);
nor U14095 (N_14095,N_13875,N_13910);
and U14096 (N_14096,N_13885,N_13954);
nor U14097 (N_14097,N_13919,N_13933);
and U14098 (N_14098,N_13908,N_13923);
and U14099 (N_14099,N_13969,N_13911);
or U14100 (N_14100,N_13878,N_13997);
nand U14101 (N_14101,N_13906,N_13926);
xor U14102 (N_14102,N_13913,N_13987);
and U14103 (N_14103,N_13907,N_13973);
and U14104 (N_14104,N_13880,N_13973);
nor U14105 (N_14105,N_13882,N_13993);
xor U14106 (N_14106,N_13970,N_13919);
and U14107 (N_14107,N_13991,N_13959);
xor U14108 (N_14108,N_13896,N_13968);
xnor U14109 (N_14109,N_13972,N_13891);
and U14110 (N_14110,N_13973,N_13979);
nor U14111 (N_14111,N_13996,N_13963);
or U14112 (N_14112,N_13938,N_13940);
and U14113 (N_14113,N_13901,N_13992);
xor U14114 (N_14114,N_13935,N_13898);
or U14115 (N_14115,N_13978,N_13918);
xor U14116 (N_14116,N_13897,N_13926);
nand U14117 (N_14117,N_13904,N_13958);
xor U14118 (N_14118,N_13919,N_13932);
or U14119 (N_14119,N_13888,N_13918);
nand U14120 (N_14120,N_13973,N_13954);
xor U14121 (N_14121,N_13947,N_13937);
nand U14122 (N_14122,N_13990,N_13941);
nor U14123 (N_14123,N_13902,N_13881);
nor U14124 (N_14124,N_13911,N_13960);
nor U14125 (N_14125,N_14066,N_14100);
or U14126 (N_14126,N_14106,N_14006);
nand U14127 (N_14127,N_14071,N_14097);
nand U14128 (N_14128,N_14114,N_14069);
xnor U14129 (N_14129,N_14107,N_14054);
nand U14130 (N_14130,N_14079,N_14012);
nand U14131 (N_14131,N_14074,N_14095);
and U14132 (N_14132,N_14109,N_14029);
and U14133 (N_14133,N_14049,N_14008);
nand U14134 (N_14134,N_14021,N_14042);
nor U14135 (N_14135,N_14009,N_14034);
and U14136 (N_14136,N_14113,N_14058);
nor U14137 (N_14137,N_14031,N_14033);
and U14138 (N_14138,N_14086,N_14002);
or U14139 (N_14139,N_14035,N_14048);
nand U14140 (N_14140,N_14024,N_14055);
or U14141 (N_14141,N_14124,N_14121);
and U14142 (N_14142,N_14115,N_14019);
nor U14143 (N_14143,N_14089,N_14045);
nand U14144 (N_14144,N_14120,N_14040);
or U14145 (N_14145,N_14085,N_14038);
nor U14146 (N_14146,N_14015,N_14025);
nand U14147 (N_14147,N_14117,N_14087);
nand U14148 (N_14148,N_14057,N_14083);
and U14149 (N_14149,N_14103,N_14112);
and U14150 (N_14150,N_14123,N_14119);
or U14151 (N_14151,N_14047,N_14014);
nand U14152 (N_14152,N_14070,N_14023);
and U14153 (N_14153,N_14041,N_14059);
nand U14154 (N_14154,N_14007,N_14108);
and U14155 (N_14155,N_14068,N_14090);
and U14156 (N_14156,N_14036,N_14032);
nor U14157 (N_14157,N_14030,N_14018);
xor U14158 (N_14158,N_14000,N_14111);
nand U14159 (N_14159,N_14118,N_14122);
and U14160 (N_14160,N_14056,N_14026);
nand U14161 (N_14161,N_14078,N_14016);
xor U14162 (N_14162,N_14064,N_14062);
nor U14163 (N_14163,N_14094,N_14099);
nand U14164 (N_14164,N_14101,N_14005);
or U14165 (N_14165,N_14098,N_14053);
xor U14166 (N_14166,N_14081,N_14076);
and U14167 (N_14167,N_14017,N_14116);
xnor U14168 (N_14168,N_14088,N_14096);
xnor U14169 (N_14169,N_14067,N_14065);
or U14170 (N_14170,N_14104,N_14050);
xor U14171 (N_14171,N_14011,N_14072);
xnor U14172 (N_14172,N_14080,N_14051);
and U14173 (N_14173,N_14102,N_14020);
nand U14174 (N_14174,N_14075,N_14046);
and U14175 (N_14175,N_14077,N_14022);
nor U14176 (N_14176,N_14060,N_14039);
nor U14177 (N_14177,N_14091,N_14084);
or U14178 (N_14178,N_14043,N_14013);
nand U14179 (N_14179,N_14105,N_14010);
nand U14180 (N_14180,N_14110,N_14003);
nor U14181 (N_14181,N_14001,N_14044);
xor U14182 (N_14182,N_14037,N_14027);
and U14183 (N_14183,N_14073,N_14063);
nand U14184 (N_14184,N_14052,N_14028);
or U14185 (N_14185,N_14004,N_14082);
or U14186 (N_14186,N_14093,N_14061);
xor U14187 (N_14187,N_14092,N_14022);
xor U14188 (N_14188,N_14081,N_14008);
nand U14189 (N_14189,N_14045,N_14051);
or U14190 (N_14190,N_14119,N_14023);
nand U14191 (N_14191,N_14083,N_14093);
or U14192 (N_14192,N_14063,N_14019);
xnor U14193 (N_14193,N_14038,N_14065);
nor U14194 (N_14194,N_14067,N_14020);
xnor U14195 (N_14195,N_14058,N_14077);
or U14196 (N_14196,N_14114,N_14088);
or U14197 (N_14197,N_14014,N_14082);
xnor U14198 (N_14198,N_14018,N_14015);
or U14199 (N_14199,N_14031,N_14112);
nand U14200 (N_14200,N_14064,N_14047);
and U14201 (N_14201,N_14054,N_14029);
nor U14202 (N_14202,N_14099,N_14013);
nor U14203 (N_14203,N_14013,N_14122);
or U14204 (N_14204,N_14084,N_14103);
and U14205 (N_14205,N_14056,N_14117);
or U14206 (N_14206,N_14045,N_14026);
xor U14207 (N_14207,N_14070,N_14039);
nand U14208 (N_14208,N_14091,N_14046);
and U14209 (N_14209,N_14010,N_14007);
or U14210 (N_14210,N_14009,N_14036);
and U14211 (N_14211,N_14039,N_14065);
and U14212 (N_14212,N_14119,N_14071);
nand U14213 (N_14213,N_14079,N_14054);
nand U14214 (N_14214,N_14051,N_14026);
nand U14215 (N_14215,N_14070,N_14095);
nor U14216 (N_14216,N_14085,N_14071);
or U14217 (N_14217,N_14057,N_14120);
or U14218 (N_14218,N_14030,N_14062);
or U14219 (N_14219,N_14092,N_14091);
and U14220 (N_14220,N_14088,N_14070);
nand U14221 (N_14221,N_14066,N_14031);
xor U14222 (N_14222,N_14057,N_14077);
and U14223 (N_14223,N_14062,N_14039);
xor U14224 (N_14224,N_14088,N_14068);
and U14225 (N_14225,N_14055,N_14061);
nand U14226 (N_14226,N_14006,N_14054);
nand U14227 (N_14227,N_14121,N_14083);
and U14228 (N_14228,N_14104,N_14089);
and U14229 (N_14229,N_14073,N_14082);
and U14230 (N_14230,N_14057,N_14075);
and U14231 (N_14231,N_14068,N_14054);
nor U14232 (N_14232,N_14068,N_14077);
nor U14233 (N_14233,N_14098,N_14012);
and U14234 (N_14234,N_14083,N_14054);
nor U14235 (N_14235,N_14115,N_14067);
xor U14236 (N_14236,N_14059,N_14056);
xnor U14237 (N_14237,N_14002,N_14107);
and U14238 (N_14238,N_14052,N_14069);
nor U14239 (N_14239,N_14049,N_14000);
xor U14240 (N_14240,N_14060,N_14041);
nor U14241 (N_14241,N_14053,N_14121);
or U14242 (N_14242,N_14041,N_14056);
nand U14243 (N_14243,N_14056,N_14079);
or U14244 (N_14244,N_14064,N_14099);
nand U14245 (N_14245,N_14048,N_14021);
and U14246 (N_14246,N_14058,N_14019);
xnor U14247 (N_14247,N_14121,N_14097);
or U14248 (N_14248,N_14080,N_14006);
xnor U14249 (N_14249,N_14071,N_14007);
nand U14250 (N_14250,N_14192,N_14186);
nand U14251 (N_14251,N_14137,N_14188);
nor U14252 (N_14252,N_14162,N_14206);
and U14253 (N_14253,N_14177,N_14190);
xnor U14254 (N_14254,N_14242,N_14146);
nor U14255 (N_14255,N_14141,N_14163);
and U14256 (N_14256,N_14182,N_14194);
or U14257 (N_14257,N_14208,N_14169);
or U14258 (N_14258,N_14241,N_14143);
and U14259 (N_14259,N_14217,N_14213);
xor U14260 (N_14260,N_14126,N_14157);
nor U14261 (N_14261,N_14136,N_14171);
xor U14262 (N_14262,N_14230,N_14138);
and U14263 (N_14263,N_14127,N_14214);
or U14264 (N_14264,N_14215,N_14153);
xnor U14265 (N_14265,N_14232,N_14203);
and U14266 (N_14266,N_14142,N_14202);
nor U14267 (N_14267,N_14246,N_14201);
xor U14268 (N_14268,N_14140,N_14174);
and U14269 (N_14269,N_14160,N_14204);
or U14270 (N_14270,N_14187,N_14147);
and U14271 (N_14271,N_14144,N_14245);
or U14272 (N_14272,N_14235,N_14132);
nor U14273 (N_14273,N_14210,N_14154);
nor U14274 (N_14274,N_14229,N_14216);
nor U14275 (N_14275,N_14133,N_14191);
xor U14276 (N_14276,N_14185,N_14247);
xor U14277 (N_14277,N_14244,N_14239);
or U14278 (N_14278,N_14131,N_14149);
nand U14279 (N_14279,N_14172,N_14207);
nand U14280 (N_14280,N_14195,N_14128);
xnor U14281 (N_14281,N_14180,N_14234);
nand U14282 (N_14282,N_14205,N_14218);
nand U14283 (N_14283,N_14223,N_14167);
nand U14284 (N_14284,N_14130,N_14184);
and U14285 (N_14285,N_14166,N_14220);
and U14286 (N_14286,N_14225,N_14139);
nor U14287 (N_14287,N_14237,N_14240);
and U14288 (N_14288,N_14145,N_14125);
nor U14289 (N_14289,N_14156,N_14151);
xor U14290 (N_14290,N_14159,N_14212);
xnor U14291 (N_14291,N_14238,N_14152);
xor U14292 (N_14292,N_14189,N_14134);
or U14293 (N_14293,N_14209,N_14211);
and U14294 (N_14294,N_14228,N_14227);
nor U14295 (N_14295,N_14249,N_14179);
or U14296 (N_14296,N_14193,N_14231);
nand U14297 (N_14297,N_14135,N_14197);
nand U14298 (N_14298,N_14183,N_14221);
and U14299 (N_14299,N_14178,N_14173);
nand U14300 (N_14300,N_14155,N_14181);
nor U14301 (N_14301,N_14224,N_14226);
nand U14302 (N_14302,N_14219,N_14148);
and U14303 (N_14303,N_14199,N_14161);
xnor U14304 (N_14304,N_14175,N_14158);
nor U14305 (N_14305,N_14129,N_14222);
and U14306 (N_14306,N_14196,N_14248);
nor U14307 (N_14307,N_14168,N_14170);
or U14308 (N_14308,N_14198,N_14164);
xor U14309 (N_14309,N_14150,N_14243);
nand U14310 (N_14310,N_14236,N_14165);
or U14311 (N_14311,N_14176,N_14233);
nand U14312 (N_14312,N_14200,N_14131);
xnor U14313 (N_14313,N_14228,N_14191);
and U14314 (N_14314,N_14133,N_14242);
xnor U14315 (N_14315,N_14153,N_14191);
or U14316 (N_14316,N_14163,N_14130);
nor U14317 (N_14317,N_14176,N_14203);
nor U14318 (N_14318,N_14193,N_14239);
and U14319 (N_14319,N_14243,N_14192);
and U14320 (N_14320,N_14132,N_14178);
or U14321 (N_14321,N_14216,N_14142);
nor U14322 (N_14322,N_14223,N_14215);
xor U14323 (N_14323,N_14228,N_14169);
xnor U14324 (N_14324,N_14213,N_14176);
and U14325 (N_14325,N_14179,N_14234);
nand U14326 (N_14326,N_14176,N_14247);
nand U14327 (N_14327,N_14216,N_14219);
and U14328 (N_14328,N_14138,N_14187);
nand U14329 (N_14329,N_14151,N_14134);
nor U14330 (N_14330,N_14172,N_14126);
nand U14331 (N_14331,N_14227,N_14173);
nor U14332 (N_14332,N_14125,N_14186);
nor U14333 (N_14333,N_14145,N_14155);
nand U14334 (N_14334,N_14135,N_14153);
xnor U14335 (N_14335,N_14161,N_14128);
nand U14336 (N_14336,N_14211,N_14200);
and U14337 (N_14337,N_14136,N_14227);
nand U14338 (N_14338,N_14225,N_14133);
and U14339 (N_14339,N_14131,N_14144);
nor U14340 (N_14340,N_14155,N_14137);
nand U14341 (N_14341,N_14194,N_14165);
and U14342 (N_14342,N_14194,N_14128);
or U14343 (N_14343,N_14127,N_14233);
nand U14344 (N_14344,N_14206,N_14221);
xnor U14345 (N_14345,N_14157,N_14200);
xnor U14346 (N_14346,N_14221,N_14189);
nand U14347 (N_14347,N_14176,N_14133);
or U14348 (N_14348,N_14152,N_14191);
nor U14349 (N_14349,N_14162,N_14132);
or U14350 (N_14350,N_14232,N_14205);
nor U14351 (N_14351,N_14248,N_14221);
nor U14352 (N_14352,N_14232,N_14127);
and U14353 (N_14353,N_14151,N_14147);
nor U14354 (N_14354,N_14224,N_14185);
nand U14355 (N_14355,N_14208,N_14220);
and U14356 (N_14356,N_14249,N_14156);
and U14357 (N_14357,N_14239,N_14232);
nand U14358 (N_14358,N_14248,N_14134);
or U14359 (N_14359,N_14157,N_14179);
and U14360 (N_14360,N_14227,N_14245);
xnor U14361 (N_14361,N_14213,N_14195);
or U14362 (N_14362,N_14235,N_14202);
xor U14363 (N_14363,N_14235,N_14179);
xnor U14364 (N_14364,N_14229,N_14219);
or U14365 (N_14365,N_14200,N_14221);
nor U14366 (N_14366,N_14173,N_14139);
xnor U14367 (N_14367,N_14189,N_14196);
nand U14368 (N_14368,N_14236,N_14187);
or U14369 (N_14369,N_14221,N_14139);
nor U14370 (N_14370,N_14176,N_14236);
nand U14371 (N_14371,N_14239,N_14209);
xnor U14372 (N_14372,N_14125,N_14176);
nor U14373 (N_14373,N_14209,N_14127);
xnor U14374 (N_14374,N_14222,N_14210);
xor U14375 (N_14375,N_14356,N_14366);
nand U14376 (N_14376,N_14266,N_14348);
xor U14377 (N_14377,N_14273,N_14373);
xor U14378 (N_14378,N_14260,N_14309);
and U14379 (N_14379,N_14311,N_14335);
xor U14380 (N_14380,N_14364,N_14282);
nor U14381 (N_14381,N_14359,N_14265);
or U14382 (N_14382,N_14275,N_14302);
nor U14383 (N_14383,N_14325,N_14319);
and U14384 (N_14384,N_14299,N_14308);
and U14385 (N_14385,N_14307,N_14271);
nor U14386 (N_14386,N_14353,N_14339);
nor U14387 (N_14387,N_14341,N_14284);
or U14388 (N_14388,N_14371,N_14327);
xnor U14389 (N_14389,N_14368,N_14262);
or U14390 (N_14390,N_14357,N_14297);
nand U14391 (N_14391,N_14355,N_14318);
nor U14392 (N_14392,N_14343,N_14369);
and U14393 (N_14393,N_14291,N_14306);
or U14394 (N_14394,N_14250,N_14362);
nand U14395 (N_14395,N_14283,N_14269);
nor U14396 (N_14396,N_14293,N_14290);
nand U14397 (N_14397,N_14324,N_14314);
nand U14398 (N_14398,N_14360,N_14257);
and U14399 (N_14399,N_14258,N_14298);
xnor U14400 (N_14400,N_14288,N_14286);
nor U14401 (N_14401,N_14281,N_14331);
and U14402 (N_14402,N_14345,N_14256);
or U14403 (N_14403,N_14321,N_14304);
nand U14404 (N_14404,N_14268,N_14278);
xor U14405 (N_14405,N_14323,N_14361);
nor U14406 (N_14406,N_14363,N_14253);
and U14407 (N_14407,N_14365,N_14277);
xor U14408 (N_14408,N_14350,N_14251);
xnor U14409 (N_14409,N_14329,N_14272);
nand U14410 (N_14410,N_14270,N_14263);
nor U14411 (N_14411,N_14276,N_14274);
and U14412 (N_14412,N_14374,N_14316);
nor U14413 (N_14413,N_14344,N_14349);
or U14414 (N_14414,N_14295,N_14328);
xor U14415 (N_14415,N_14342,N_14254);
nand U14416 (N_14416,N_14322,N_14338);
or U14417 (N_14417,N_14303,N_14351);
and U14418 (N_14418,N_14354,N_14313);
xnor U14419 (N_14419,N_14336,N_14333);
nor U14420 (N_14420,N_14301,N_14315);
or U14421 (N_14421,N_14264,N_14358);
and U14422 (N_14422,N_14280,N_14261);
xor U14423 (N_14423,N_14255,N_14317);
or U14424 (N_14424,N_14372,N_14305);
xnor U14425 (N_14425,N_14346,N_14289);
or U14426 (N_14426,N_14370,N_14285);
or U14427 (N_14427,N_14330,N_14337);
xnor U14428 (N_14428,N_14326,N_14294);
and U14429 (N_14429,N_14334,N_14252);
and U14430 (N_14430,N_14340,N_14347);
or U14431 (N_14431,N_14292,N_14332);
nand U14432 (N_14432,N_14259,N_14352);
nand U14433 (N_14433,N_14367,N_14300);
nor U14434 (N_14434,N_14296,N_14310);
xnor U14435 (N_14435,N_14267,N_14287);
xnor U14436 (N_14436,N_14320,N_14279);
nand U14437 (N_14437,N_14312,N_14303);
nor U14438 (N_14438,N_14259,N_14294);
and U14439 (N_14439,N_14292,N_14323);
xnor U14440 (N_14440,N_14364,N_14266);
nor U14441 (N_14441,N_14351,N_14305);
and U14442 (N_14442,N_14266,N_14353);
nor U14443 (N_14443,N_14374,N_14285);
nor U14444 (N_14444,N_14361,N_14371);
and U14445 (N_14445,N_14253,N_14312);
nand U14446 (N_14446,N_14297,N_14271);
nand U14447 (N_14447,N_14347,N_14360);
nand U14448 (N_14448,N_14328,N_14348);
or U14449 (N_14449,N_14262,N_14270);
and U14450 (N_14450,N_14322,N_14264);
and U14451 (N_14451,N_14289,N_14372);
xor U14452 (N_14452,N_14347,N_14313);
nor U14453 (N_14453,N_14257,N_14300);
nand U14454 (N_14454,N_14337,N_14287);
and U14455 (N_14455,N_14318,N_14344);
and U14456 (N_14456,N_14328,N_14314);
and U14457 (N_14457,N_14364,N_14320);
nor U14458 (N_14458,N_14251,N_14339);
xnor U14459 (N_14459,N_14252,N_14270);
nand U14460 (N_14460,N_14371,N_14330);
nand U14461 (N_14461,N_14330,N_14302);
nor U14462 (N_14462,N_14335,N_14352);
and U14463 (N_14463,N_14335,N_14369);
and U14464 (N_14464,N_14311,N_14250);
or U14465 (N_14465,N_14340,N_14265);
or U14466 (N_14466,N_14366,N_14369);
xnor U14467 (N_14467,N_14348,N_14361);
nor U14468 (N_14468,N_14304,N_14325);
nor U14469 (N_14469,N_14359,N_14336);
nand U14470 (N_14470,N_14283,N_14320);
xor U14471 (N_14471,N_14313,N_14309);
or U14472 (N_14472,N_14351,N_14372);
nor U14473 (N_14473,N_14283,N_14303);
nor U14474 (N_14474,N_14366,N_14275);
nor U14475 (N_14475,N_14266,N_14317);
or U14476 (N_14476,N_14287,N_14320);
nand U14477 (N_14477,N_14255,N_14304);
xor U14478 (N_14478,N_14370,N_14366);
nand U14479 (N_14479,N_14359,N_14320);
and U14480 (N_14480,N_14298,N_14327);
xor U14481 (N_14481,N_14350,N_14282);
nand U14482 (N_14482,N_14310,N_14325);
or U14483 (N_14483,N_14297,N_14339);
xnor U14484 (N_14484,N_14363,N_14329);
or U14485 (N_14485,N_14289,N_14252);
and U14486 (N_14486,N_14285,N_14310);
xnor U14487 (N_14487,N_14374,N_14256);
nand U14488 (N_14488,N_14294,N_14296);
and U14489 (N_14489,N_14315,N_14286);
nor U14490 (N_14490,N_14313,N_14336);
nor U14491 (N_14491,N_14337,N_14267);
or U14492 (N_14492,N_14351,N_14360);
and U14493 (N_14493,N_14261,N_14312);
nand U14494 (N_14494,N_14284,N_14310);
or U14495 (N_14495,N_14352,N_14336);
nand U14496 (N_14496,N_14269,N_14373);
and U14497 (N_14497,N_14335,N_14371);
nor U14498 (N_14498,N_14264,N_14362);
xnor U14499 (N_14499,N_14343,N_14256);
nor U14500 (N_14500,N_14453,N_14477);
nor U14501 (N_14501,N_14486,N_14387);
or U14502 (N_14502,N_14417,N_14424);
xnor U14503 (N_14503,N_14400,N_14393);
nand U14504 (N_14504,N_14420,N_14497);
xnor U14505 (N_14505,N_14415,N_14383);
nor U14506 (N_14506,N_14457,N_14391);
and U14507 (N_14507,N_14482,N_14448);
and U14508 (N_14508,N_14459,N_14480);
nor U14509 (N_14509,N_14499,N_14432);
or U14510 (N_14510,N_14474,N_14398);
or U14511 (N_14511,N_14469,N_14454);
and U14512 (N_14512,N_14492,N_14450);
nand U14513 (N_14513,N_14407,N_14449);
nand U14514 (N_14514,N_14413,N_14498);
nor U14515 (N_14515,N_14433,N_14409);
or U14516 (N_14516,N_14378,N_14485);
xnor U14517 (N_14517,N_14496,N_14389);
nor U14518 (N_14518,N_14472,N_14437);
nand U14519 (N_14519,N_14476,N_14428);
nand U14520 (N_14520,N_14458,N_14452);
xor U14521 (N_14521,N_14468,N_14402);
nor U14522 (N_14522,N_14431,N_14401);
nand U14523 (N_14523,N_14456,N_14435);
and U14524 (N_14524,N_14466,N_14444);
or U14525 (N_14525,N_14399,N_14426);
and U14526 (N_14526,N_14479,N_14385);
and U14527 (N_14527,N_14493,N_14462);
nand U14528 (N_14528,N_14390,N_14436);
nor U14529 (N_14529,N_14441,N_14404);
and U14530 (N_14530,N_14487,N_14419);
nor U14531 (N_14531,N_14429,N_14384);
or U14532 (N_14532,N_14397,N_14381);
or U14533 (N_14533,N_14425,N_14447);
nand U14534 (N_14534,N_14460,N_14408);
nand U14535 (N_14535,N_14388,N_14395);
nand U14536 (N_14536,N_14489,N_14396);
or U14537 (N_14537,N_14438,N_14494);
xnor U14538 (N_14538,N_14434,N_14377);
nor U14539 (N_14539,N_14386,N_14430);
and U14540 (N_14540,N_14427,N_14392);
or U14541 (N_14541,N_14481,N_14475);
nor U14542 (N_14542,N_14414,N_14418);
and U14543 (N_14543,N_14446,N_14406);
nand U14544 (N_14544,N_14464,N_14440);
xnor U14545 (N_14545,N_14490,N_14412);
and U14546 (N_14546,N_14423,N_14445);
or U14547 (N_14547,N_14484,N_14376);
and U14548 (N_14548,N_14394,N_14411);
nand U14549 (N_14549,N_14491,N_14461);
nand U14550 (N_14550,N_14442,N_14421);
and U14551 (N_14551,N_14478,N_14467);
and U14552 (N_14552,N_14379,N_14439);
and U14553 (N_14553,N_14375,N_14483);
or U14554 (N_14554,N_14465,N_14470);
or U14555 (N_14555,N_14455,N_14382);
and U14556 (N_14556,N_14416,N_14463);
and U14557 (N_14557,N_14422,N_14471);
and U14558 (N_14558,N_14380,N_14488);
or U14559 (N_14559,N_14495,N_14451);
nor U14560 (N_14560,N_14410,N_14473);
xnor U14561 (N_14561,N_14403,N_14443);
xor U14562 (N_14562,N_14405,N_14439);
and U14563 (N_14563,N_14467,N_14377);
nor U14564 (N_14564,N_14462,N_14440);
xnor U14565 (N_14565,N_14416,N_14486);
xor U14566 (N_14566,N_14480,N_14452);
and U14567 (N_14567,N_14414,N_14438);
or U14568 (N_14568,N_14476,N_14497);
nand U14569 (N_14569,N_14489,N_14494);
or U14570 (N_14570,N_14447,N_14453);
xnor U14571 (N_14571,N_14407,N_14404);
or U14572 (N_14572,N_14421,N_14431);
nand U14573 (N_14573,N_14464,N_14384);
nand U14574 (N_14574,N_14485,N_14480);
or U14575 (N_14575,N_14444,N_14393);
nand U14576 (N_14576,N_14495,N_14461);
and U14577 (N_14577,N_14475,N_14454);
or U14578 (N_14578,N_14377,N_14490);
nand U14579 (N_14579,N_14402,N_14401);
or U14580 (N_14580,N_14417,N_14438);
nor U14581 (N_14581,N_14466,N_14464);
xnor U14582 (N_14582,N_14484,N_14463);
nor U14583 (N_14583,N_14448,N_14399);
nand U14584 (N_14584,N_14465,N_14426);
xor U14585 (N_14585,N_14475,N_14417);
and U14586 (N_14586,N_14410,N_14425);
nand U14587 (N_14587,N_14485,N_14432);
xnor U14588 (N_14588,N_14498,N_14478);
nor U14589 (N_14589,N_14497,N_14474);
xnor U14590 (N_14590,N_14473,N_14455);
and U14591 (N_14591,N_14378,N_14423);
and U14592 (N_14592,N_14477,N_14440);
nor U14593 (N_14593,N_14429,N_14463);
nor U14594 (N_14594,N_14388,N_14377);
and U14595 (N_14595,N_14472,N_14474);
nor U14596 (N_14596,N_14426,N_14411);
xnor U14597 (N_14597,N_14394,N_14425);
xnor U14598 (N_14598,N_14494,N_14389);
xor U14599 (N_14599,N_14455,N_14468);
nor U14600 (N_14600,N_14469,N_14470);
nand U14601 (N_14601,N_14398,N_14380);
nand U14602 (N_14602,N_14403,N_14385);
nand U14603 (N_14603,N_14391,N_14406);
and U14604 (N_14604,N_14480,N_14466);
nor U14605 (N_14605,N_14418,N_14387);
and U14606 (N_14606,N_14462,N_14424);
nand U14607 (N_14607,N_14429,N_14415);
xor U14608 (N_14608,N_14407,N_14428);
xnor U14609 (N_14609,N_14465,N_14405);
xnor U14610 (N_14610,N_14425,N_14380);
nor U14611 (N_14611,N_14413,N_14414);
and U14612 (N_14612,N_14478,N_14416);
nor U14613 (N_14613,N_14465,N_14393);
nand U14614 (N_14614,N_14380,N_14446);
nor U14615 (N_14615,N_14477,N_14446);
nor U14616 (N_14616,N_14439,N_14489);
nor U14617 (N_14617,N_14392,N_14486);
and U14618 (N_14618,N_14468,N_14400);
or U14619 (N_14619,N_14414,N_14411);
xnor U14620 (N_14620,N_14485,N_14426);
or U14621 (N_14621,N_14394,N_14473);
nand U14622 (N_14622,N_14390,N_14388);
and U14623 (N_14623,N_14416,N_14468);
xnor U14624 (N_14624,N_14412,N_14481);
and U14625 (N_14625,N_14605,N_14580);
nand U14626 (N_14626,N_14570,N_14608);
nand U14627 (N_14627,N_14573,N_14622);
and U14628 (N_14628,N_14613,N_14597);
or U14629 (N_14629,N_14583,N_14504);
nand U14630 (N_14630,N_14530,N_14609);
xor U14631 (N_14631,N_14552,N_14546);
nand U14632 (N_14632,N_14562,N_14617);
or U14633 (N_14633,N_14620,N_14574);
nand U14634 (N_14634,N_14558,N_14533);
xnor U14635 (N_14635,N_14621,N_14528);
xor U14636 (N_14636,N_14551,N_14518);
or U14637 (N_14637,N_14611,N_14598);
xnor U14638 (N_14638,N_14579,N_14590);
or U14639 (N_14639,N_14523,N_14601);
nand U14640 (N_14640,N_14526,N_14501);
xnor U14641 (N_14641,N_14584,N_14527);
nor U14642 (N_14642,N_14540,N_14503);
or U14643 (N_14643,N_14596,N_14511);
or U14644 (N_14644,N_14522,N_14535);
or U14645 (N_14645,N_14624,N_14588);
nor U14646 (N_14646,N_14532,N_14578);
and U14647 (N_14647,N_14568,N_14543);
xor U14648 (N_14648,N_14560,N_14555);
or U14649 (N_14649,N_14525,N_14582);
nor U14650 (N_14650,N_14614,N_14615);
xor U14651 (N_14651,N_14564,N_14516);
or U14652 (N_14652,N_14524,N_14505);
or U14653 (N_14653,N_14542,N_14548);
and U14654 (N_14654,N_14545,N_14619);
nand U14655 (N_14655,N_14571,N_14592);
or U14656 (N_14656,N_14586,N_14616);
and U14657 (N_14657,N_14514,N_14610);
and U14658 (N_14658,N_14618,N_14581);
nand U14659 (N_14659,N_14506,N_14607);
nor U14660 (N_14660,N_14509,N_14572);
xnor U14661 (N_14661,N_14539,N_14512);
xor U14662 (N_14662,N_14561,N_14566);
xnor U14663 (N_14663,N_14623,N_14585);
and U14664 (N_14664,N_14591,N_14553);
or U14665 (N_14665,N_14577,N_14536);
or U14666 (N_14666,N_14565,N_14517);
xnor U14667 (N_14667,N_14569,N_14507);
nor U14668 (N_14668,N_14547,N_14554);
nor U14669 (N_14669,N_14567,N_14531);
or U14670 (N_14670,N_14550,N_14500);
and U14671 (N_14671,N_14576,N_14603);
and U14672 (N_14672,N_14515,N_14602);
or U14673 (N_14673,N_14556,N_14595);
xor U14674 (N_14674,N_14529,N_14541);
xnor U14675 (N_14675,N_14508,N_14519);
nor U14676 (N_14676,N_14612,N_14589);
xnor U14677 (N_14677,N_14606,N_14513);
nand U14678 (N_14678,N_14600,N_14549);
and U14679 (N_14679,N_14537,N_14594);
xor U14680 (N_14680,N_14557,N_14563);
xor U14681 (N_14681,N_14599,N_14544);
nand U14682 (N_14682,N_14502,N_14604);
nor U14683 (N_14683,N_14521,N_14510);
nand U14684 (N_14684,N_14559,N_14520);
or U14685 (N_14685,N_14575,N_14593);
or U14686 (N_14686,N_14587,N_14534);
nor U14687 (N_14687,N_14538,N_14576);
nand U14688 (N_14688,N_14592,N_14572);
xor U14689 (N_14689,N_14593,N_14580);
nor U14690 (N_14690,N_14607,N_14578);
or U14691 (N_14691,N_14590,N_14551);
nand U14692 (N_14692,N_14616,N_14596);
xnor U14693 (N_14693,N_14514,N_14501);
or U14694 (N_14694,N_14585,N_14580);
and U14695 (N_14695,N_14529,N_14510);
nand U14696 (N_14696,N_14577,N_14507);
nand U14697 (N_14697,N_14583,N_14518);
and U14698 (N_14698,N_14603,N_14513);
nor U14699 (N_14699,N_14589,N_14536);
and U14700 (N_14700,N_14550,N_14524);
nand U14701 (N_14701,N_14524,N_14620);
or U14702 (N_14702,N_14580,N_14596);
and U14703 (N_14703,N_14538,N_14522);
xnor U14704 (N_14704,N_14602,N_14592);
xnor U14705 (N_14705,N_14557,N_14624);
nand U14706 (N_14706,N_14505,N_14513);
nor U14707 (N_14707,N_14515,N_14598);
and U14708 (N_14708,N_14553,N_14500);
and U14709 (N_14709,N_14519,N_14558);
or U14710 (N_14710,N_14558,N_14568);
nand U14711 (N_14711,N_14518,N_14592);
nand U14712 (N_14712,N_14523,N_14610);
nor U14713 (N_14713,N_14579,N_14593);
nor U14714 (N_14714,N_14614,N_14523);
and U14715 (N_14715,N_14521,N_14503);
xnor U14716 (N_14716,N_14567,N_14521);
or U14717 (N_14717,N_14591,N_14559);
or U14718 (N_14718,N_14599,N_14611);
and U14719 (N_14719,N_14595,N_14603);
or U14720 (N_14720,N_14554,N_14561);
and U14721 (N_14721,N_14599,N_14543);
xnor U14722 (N_14722,N_14610,N_14593);
or U14723 (N_14723,N_14570,N_14621);
or U14724 (N_14724,N_14507,N_14605);
xnor U14725 (N_14725,N_14558,N_14508);
and U14726 (N_14726,N_14542,N_14588);
nor U14727 (N_14727,N_14568,N_14583);
and U14728 (N_14728,N_14504,N_14551);
nor U14729 (N_14729,N_14545,N_14610);
or U14730 (N_14730,N_14594,N_14519);
xnor U14731 (N_14731,N_14538,N_14563);
nor U14732 (N_14732,N_14578,N_14521);
or U14733 (N_14733,N_14532,N_14593);
nand U14734 (N_14734,N_14589,N_14543);
and U14735 (N_14735,N_14574,N_14575);
nand U14736 (N_14736,N_14553,N_14573);
and U14737 (N_14737,N_14594,N_14500);
nand U14738 (N_14738,N_14525,N_14607);
nor U14739 (N_14739,N_14616,N_14568);
and U14740 (N_14740,N_14554,N_14566);
or U14741 (N_14741,N_14525,N_14601);
nor U14742 (N_14742,N_14610,N_14525);
xor U14743 (N_14743,N_14569,N_14512);
and U14744 (N_14744,N_14557,N_14503);
nor U14745 (N_14745,N_14503,N_14559);
nand U14746 (N_14746,N_14514,N_14597);
xor U14747 (N_14747,N_14551,N_14588);
nor U14748 (N_14748,N_14572,N_14515);
nor U14749 (N_14749,N_14506,N_14610);
nor U14750 (N_14750,N_14722,N_14627);
and U14751 (N_14751,N_14637,N_14736);
and U14752 (N_14752,N_14672,N_14701);
nor U14753 (N_14753,N_14679,N_14636);
or U14754 (N_14754,N_14694,N_14646);
or U14755 (N_14755,N_14669,N_14697);
nor U14756 (N_14756,N_14690,N_14630);
nor U14757 (N_14757,N_14700,N_14642);
and U14758 (N_14758,N_14717,N_14635);
or U14759 (N_14759,N_14665,N_14725);
and U14760 (N_14760,N_14683,N_14698);
and U14761 (N_14761,N_14654,N_14734);
nor U14762 (N_14762,N_14675,N_14677);
xor U14763 (N_14763,N_14703,N_14656);
nor U14764 (N_14764,N_14727,N_14664);
nand U14765 (N_14765,N_14631,N_14738);
nand U14766 (N_14766,N_14680,N_14660);
xnor U14767 (N_14767,N_14641,N_14744);
xor U14768 (N_14768,N_14692,N_14709);
xor U14769 (N_14769,N_14671,N_14676);
xnor U14770 (N_14770,N_14657,N_14640);
and U14771 (N_14771,N_14720,N_14684);
xnor U14772 (N_14772,N_14745,N_14643);
nor U14773 (N_14773,N_14693,N_14714);
or U14774 (N_14774,N_14749,N_14689);
xnor U14775 (N_14775,N_14748,N_14723);
xnor U14776 (N_14776,N_14696,N_14634);
nor U14777 (N_14777,N_14726,N_14702);
xor U14778 (N_14778,N_14710,N_14741);
and U14779 (N_14779,N_14663,N_14705);
and U14780 (N_14780,N_14712,N_14649);
nor U14781 (N_14781,N_14629,N_14678);
xor U14782 (N_14782,N_14668,N_14733);
and U14783 (N_14783,N_14732,N_14651);
and U14784 (N_14784,N_14713,N_14666);
and U14785 (N_14785,N_14674,N_14719);
nor U14786 (N_14786,N_14721,N_14648);
and U14787 (N_14787,N_14687,N_14718);
and U14788 (N_14788,N_14743,N_14708);
nand U14789 (N_14789,N_14673,N_14633);
nand U14790 (N_14790,N_14658,N_14729);
nor U14791 (N_14791,N_14706,N_14670);
nand U14792 (N_14792,N_14638,N_14695);
nand U14793 (N_14793,N_14711,N_14647);
nand U14794 (N_14794,N_14691,N_14681);
nor U14795 (N_14795,N_14661,N_14728);
nand U14796 (N_14796,N_14626,N_14682);
nand U14797 (N_14797,N_14662,N_14655);
or U14798 (N_14798,N_14716,N_14686);
and U14799 (N_14799,N_14735,N_14652);
or U14800 (N_14800,N_14685,N_14731);
xor U14801 (N_14801,N_14659,N_14740);
xor U14802 (N_14802,N_14704,N_14653);
nand U14803 (N_14803,N_14639,N_14747);
nand U14804 (N_14804,N_14632,N_14739);
xnor U14805 (N_14805,N_14742,N_14644);
and U14806 (N_14806,N_14724,N_14737);
and U14807 (N_14807,N_14628,N_14699);
nor U14808 (N_14808,N_14707,N_14715);
nor U14809 (N_14809,N_14730,N_14625);
and U14810 (N_14810,N_14667,N_14645);
xnor U14811 (N_14811,N_14688,N_14746);
xor U14812 (N_14812,N_14650,N_14716);
or U14813 (N_14813,N_14707,N_14723);
or U14814 (N_14814,N_14677,N_14732);
nand U14815 (N_14815,N_14636,N_14736);
nor U14816 (N_14816,N_14746,N_14660);
nand U14817 (N_14817,N_14741,N_14742);
xnor U14818 (N_14818,N_14671,N_14744);
nor U14819 (N_14819,N_14743,N_14644);
and U14820 (N_14820,N_14641,N_14735);
or U14821 (N_14821,N_14627,N_14641);
or U14822 (N_14822,N_14694,N_14727);
and U14823 (N_14823,N_14711,N_14671);
and U14824 (N_14824,N_14696,N_14719);
and U14825 (N_14825,N_14728,N_14748);
xor U14826 (N_14826,N_14731,N_14719);
nor U14827 (N_14827,N_14625,N_14639);
nand U14828 (N_14828,N_14679,N_14709);
nor U14829 (N_14829,N_14663,N_14643);
and U14830 (N_14830,N_14706,N_14667);
xor U14831 (N_14831,N_14720,N_14700);
nor U14832 (N_14832,N_14687,N_14702);
xor U14833 (N_14833,N_14628,N_14629);
or U14834 (N_14834,N_14686,N_14676);
nor U14835 (N_14835,N_14654,N_14702);
xnor U14836 (N_14836,N_14681,N_14644);
or U14837 (N_14837,N_14689,N_14703);
or U14838 (N_14838,N_14687,N_14744);
or U14839 (N_14839,N_14660,N_14669);
or U14840 (N_14840,N_14681,N_14709);
xor U14841 (N_14841,N_14701,N_14691);
and U14842 (N_14842,N_14735,N_14633);
nor U14843 (N_14843,N_14695,N_14707);
nor U14844 (N_14844,N_14713,N_14689);
and U14845 (N_14845,N_14748,N_14626);
or U14846 (N_14846,N_14721,N_14746);
or U14847 (N_14847,N_14722,N_14708);
and U14848 (N_14848,N_14650,N_14689);
nor U14849 (N_14849,N_14688,N_14629);
or U14850 (N_14850,N_14698,N_14630);
and U14851 (N_14851,N_14733,N_14734);
nand U14852 (N_14852,N_14665,N_14702);
and U14853 (N_14853,N_14693,N_14635);
xnor U14854 (N_14854,N_14729,N_14663);
or U14855 (N_14855,N_14630,N_14686);
nand U14856 (N_14856,N_14636,N_14642);
or U14857 (N_14857,N_14657,N_14729);
nor U14858 (N_14858,N_14665,N_14636);
xnor U14859 (N_14859,N_14735,N_14711);
xnor U14860 (N_14860,N_14721,N_14666);
nor U14861 (N_14861,N_14707,N_14658);
xor U14862 (N_14862,N_14646,N_14655);
and U14863 (N_14863,N_14649,N_14638);
or U14864 (N_14864,N_14725,N_14663);
nand U14865 (N_14865,N_14628,N_14666);
nor U14866 (N_14866,N_14625,N_14718);
xor U14867 (N_14867,N_14697,N_14688);
nand U14868 (N_14868,N_14678,N_14635);
or U14869 (N_14869,N_14705,N_14722);
nor U14870 (N_14870,N_14724,N_14707);
nand U14871 (N_14871,N_14647,N_14735);
xor U14872 (N_14872,N_14649,N_14735);
or U14873 (N_14873,N_14726,N_14732);
and U14874 (N_14874,N_14684,N_14666);
xnor U14875 (N_14875,N_14767,N_14790);
nor U14876 (N_14876,N_14820,N_14870);
and U14877 (N_14877,N_14801,N_14832);
nand U14878 (N_14878,N_14854,N_14798);
or U14879 (N_14879,N_14780,N_14822);
or U14880 (N_14880,N_14789,N_14837);
xor U14881 (N_14881,N_14824,N_14812);
or U14882 (N_14882,N_14873,N_14852);
and U14883 (N_14883,N_14813,N_14842);
nor U14884 (N_14884,N_14754,N_14771);
or U14885 (N_14885,N_14860,N_14847);
or U14886 (N_14886,N_14751,N_14773);
and U14887 (N_14887,N_14809,N_14840);
nor U14888 (N_14888,N_14757,N_14846);
or U14889 (N_14889,N_14831,N_14803);
nor U14890 (N_14890,N_14843,N_14755);
or U14891 (N_14891,N_14844,N_14808);
xnor U14892 (N_14892,N_14806,N_14768);
xor U14893 (N_14893,N_14792,N_14800);
xnor U14894 (N_14894,N_14821,N_14769);
or U14895 (N_14895,N_14815,N_14759);
nand U14896 (N_14896,N_14779,N_14848);
or U14897 (N_14897,N_14811,N_14807);
and U14898 (N_14898,N_14794,N_14774);
nor U14899 (N_14899,N_14845,N_14869);
or U14900 (N_14900,N_14752,N_14825);
or U14901 (N_14901,N_14851,N_14787);
nor U14902 (N_14902,N_14797,N_14859);
and U14903 (N_14903,N_14853,N_14863);
and U14904 (N_14904,N_14753,N_14758);
xnor U14905 (N_14905,N_14810,N_14857);
and U14906 (N_14906,N_14850,N_14872);
nor U14907 (N_14907,N_14839,N_14783);
xnor U14908 (N_14908,N_14817,N_14778);
nand U14909 (N_14909,N_14793,N_14855);
nand U14910 (N_14910,N_14761,N_14827);
xnor U14911 (N_14911,N_14796,N_14823);
xnor U14912 (N_14912,N_14805,N_14838);
nor U14913 (N_14913,N_14874,N_14816);
and U14914 (N_14914,N_14802,N_14781);
nor U14915 (N_14915,N_14777,N_14782);
and U14916 (N_14916,N_14829,N_14826);
or U14917 (N_14917,N_14772,N_14764);
nor U14918 (N_14918,N_14833,N_14763);
and U14919 (N_14919,N_14841,N_14865);
or U14920 (N_14920,N_14819,N_14864);
and U14921 (N_14921,N_14814,N_14835);
xor U14922 (N_14922,N_14849,N_14858);
and U14923 (N_14923,N_14775,N_14856);
xor U14924 (N_14924,N_14786,N_14868);
nand U14925 (N_14925,N_14862,N_14760);
or U14926 (N_14926,N_14866,N_14788);
and U14927 (N_14927,N_14861,N_14791);
or U14928 (N_14928,N_14834,N_14766);
and U14929 (N_14929,N_14784,N_14867);
nor U14930 (N_14930,N_14762,N_14871);
and U14931 (N_14931,N_14830,N_14795);
and U14932 (N_14932,N_14799,N_14770);
nor U14933 (N_14933,N_14756,N_14836);
nor U14934 (N_14934,N_14776,N_14818);
or U14935 (N_14935,N_14750,N_14804);
or U14936 (N_14936,N_14785,N_14765);
nand U14937 (N_14937,N_14828,N_14793);
xor U14938 (N_14938,N_14770,N_14871);
or U14939 (N_14939,N_14772,N_14780);
or U14940 (N_14940,N_14780,N_14779);
nand U14941 (N_14941,N_14770,N_14808);
nor U14942 (N_14942,N_14822,N_14848);
nand U14943 (N_14943,N_14841,N_14792);
or U14944 (N_14944,N_14829,N_14802);
nor U14945 (N_14945,N_14752,N_14780);
and U14946 (N_14946,N_14773,N_14782);
xnor U14947 (N_14947,N_14819,N_14846);
and U14948 (N_14948,N_14791,N_14763);
nor U14949 (N_14949,N_14854,N_14800);
nand U14950 (N_14950,N_14751,N_14861);
nor U14951 (N_14951,N_14812,N_14781);
nor U14952 (N_14952,N_14836,N_14754);
and U14953 (N_14953,N_14768,N_14869);
or U14954 (N_14954,N_14847,N_14818);
or U14955 (N_14955,N_14781,N_14862);
nand U14956 (N_14956,N_14765,N_14776);
or U14957 (N_14957,N_14833,N_14776);
or U14958 (N_14958,N_14843,N_14764);
and U14959 (N_14959,N_14823,N_14805);
xor U14960 (N_14960,N_14847,N_14756);
nor U14961 (N_14961,N_14831,N_14771);
and U14962 (N_14962,N_14780,N_14750);
or U14963 (N_14963,N_14763,N_14761);
nor U14964 (N_14964,N_14799,N_14849);
and U14965 (N_14965,N_14771,N_14843);
and U14966 (N_14966,N_14860,N_14796);
and U14967 (N_14967,N_14869,N_14764);
nand U14968 (N_14968,N_14791,N_14795);
nor U14969 (N_14969,N_14756,N_14857);
or U14970 (N_14970,N_14840,N_14849);
nor U14971 (N_14971,N_14759,N_14828);
nand U14972 (N_14972,N_14794,N_14757);
xor U14973 (N_14973,N_14772,N_14777);
and U14974 (N_14974,N_14785,N_14800);
xnor U14975 (N_14975,N_14834,N_14820);
nand U14976 (N_14976,N_14802,N_14796);
xor U14977 (N_14977,N_14824,N_14826);
or U14978 (N_14978,N_14873,N_14822);
or U14979 (N_14979,N_14829,N_14842);
nor U14980 (N_14980,N_14764,N_14832);
xor U14981 (N_14981,N_14755,N_14819);
xnor U14982 (N_14982,N_14822,N_14834);
nor U14983 (N_14983,N_14828,N_14757);
nand U14984 (N_14984,N_14780,N_14758);
nand U14985 (N_14985,N_14792,N_14785);
xnor U14986 (N_14986,N_14759,N_14858);
or U14987 (N_14987,N_14812,N_14789);
nor U14988 (N_14988,N_14874,N_14800);
nor U14989 (N_14989,N_14837,N_14868);
and U14990 (N_14990,N_14854,N_14846);
or U14991 (N_14991,N_14853,N_14759);
xnor U14992 (N_14992,N_14856,N_14830);
xnor U14993 (N_14993,N_14760,N_14800);
or U14994 (N_14994,N_14791,N_14803);
xor U14995 (N_14995,N_14796,N_14826);
xnor U14996 (N_14996,N_14860,N_14780);
xor U14997 (N_14997,N_14812,N_14813);
or U14998 (N_14998,N_14758,N_14859);
nand U14999 (N_14999,N_14809,N_14859);
or UO_0 (O_0,N_14889,N_14940);
xnor UO_1 (O_1,N_14947,N_14967);
and UO_2 (O_2,N_14893,N_14952);
nor UO_3 (O_3,N_14941,N_14966);
nor UO_4 (O_4,N_14953,N_14922);
nand UO_5 (O_5,N_14980,N_14897);
or UO_6 (O_6,N_14903,N_14934);
xor UO_7 (O_7,N_14951,N_14883);
nand UO_8 (O_8,N_14907,N_14987);
and UO_9 (O_9,N_14898,N_14994);
nor UO_10 (O_10,N_14964,N_14971);
xor UO_11 (O_11,N_14975,N_14976);
nand UO_12 (O_12,N_14901,N_14942);
and UO_13 (O_13,N_14880,N_14991);
and UO_14 (O_14,N_14943,N_14914);
nor UO_15 (O_15,N_14879,N_14930);
xnor UO_16 (O_16,N_14896,N_14892);
nor UO_17 (O_17,N_14918,N_14904);
nor UO_18 (O_18,N_14902,N_14977);
xor UO_19 (O_19,N_14890,N_14956);
or UO_20 (O_20,N_14959,N_14905);
nor UO_21 (O_21,N_14895,N_14950);
nor UO_22 (O_22,N_14981,N_14984);
nor UO_23 (O_23,N_14884,N_14970);
nand UO_24 (O_24,N_14995,N_14937);
nor UO_25 (O_25,N_14948,N_14972);
and UO_26 (O_26,N_14962,N_14908);
xor UO_27 (O_27,N_14891,N_14917);
or UO_28 (O_28,N_14931,N_14986);
nand UO_29 (O_29,N_14900,N_14916);
nor UO_30 (O_30,N_14978,N_14888);
and UO_31 (O_31,N_14911,N_14939);
and UO_32 (O_32,N_14965,N_14906);
or UO_33 (O_33,N_14915,N_14921);
nand UO_34 (O_34,N_14920,N_14979);
xor UO_35 (O_35,N_14909,N_14924);
nand UO_36 (O_36,N_14957,N_14945);
xnor UO_37 (O_37,N_14985,N_14919);
nor UO_38 (O_38,N_14973,N_14993);
and UO_39 (O_39,N_14946,N_14927);
or UO_40 (O_40,N_14938,N_14875);
nor UO_41 (O_41,N_14877,N_14989);
nand UO_42 (O_42,N_14899,N_14992);
or UO_43 (O_43,N_14928,N_14882);
xnor UO_44 (O_44,N_14881,N_14913);
and UO_45 (O_45,N_14960,N_14990);
or UO_46 (O_46,N_14955,N_14936);
or UO_47 (O_47,N_14998,N_14954);
nor UO_48 (O_48,N_14887,N_14969);
nor UO_49 (O_49,N_14933,N_14926);
or UO_50 (O_50,N_14983,N_14885);
or UO_51 (O_51,N_14963,N_14961);
nor UO_52 (O_52,N_14944,N_14949);
nor UO_53 (O_53,N_14912,N_14968);
xnor UO_54 (O_54,N_14878,N_14886);
xor UO_55 (O_55,N_14988,N_14932);
xor UO_56 (O_56,N_14997,N_14974);
nand UO_57 (O_57,N_14910,N_14958);
nor UO_58 (O_58,N_14999,N_14923);
and UO_59 (O_59,N_14982,N_14925);
nor UO_60 (O_60,N_14929,N_14935);
nand UO_61 (O_61,N_14894,N_14996);
xnor UO_62 (O_62,N_14876,N_14955);
xnor UO_63 (O_63,N_14927,N_14888);
or UO_64 (O_64,N_14914,N_14931);
nand UO_65 (O_65,N_14927,N_14977);
nand UO_66 (O_66,N_14906,N_14918);
nor UO_67 (O_67,N_14915,N_14908);
or UO_68 (O_68,N_14992,N_14993);
nor UO_69 (O_69,N_14895,N_14915);
or UO_70 (O_70,N_14888,N_14957);
nor UO_71 (O_71,N_14947,N_14954);
xnor UO_72 (O_72,N_14963,N_14957);
nor UO_73 (O_73,N_14995,N_14885);
nand UO_74 (O_74,N_14987,N_14966);
nand UO_75 (O_75,N_14899,N_14910);
nor UO_76 (O_76,N_14875,N_14935);
or UO_77 (O_77,N_14996,N_14895);
and UO_78 (O_78,N_14983,N_14886);
or UO_79 (O_79,N_14974,N_14947);
xnor UO_80 (O_80,N_14880,N_14905);
nand UO_81 (O_81,N_14881,N_14922);
or UO_82 (O_82,N_14964,N_14960);
and UO_83 (O_83,N_14986,N_14946);
and UO_84 (O_84,N_14898,N_14928);
xor UO_85 (O_85,N_14960,N_14995);
nor UO_86 (O_86,N_14886,N_14955);
or UO_87 (O_87,N_14991,N_14922);
nand UO_88 (O_88,N_14983,N_14907);
and UO_89 (O_89,N_14898,N_14885);
xor UO_90 (O_90,N_14876,N_14941);
xnor UO_91 (O_91,N_14982,N_14947);
nand UO_92 (O_92,N_14893,N_14899);
xor UO_93 (O_93,N_14969,N_14951);
nor UO_94 (O_94,N_14878,N_14929);
nand UO_95 (O_95,N_14903,N_14879);
nor UO_96 (O_96,N_14934,N_14964);
xor UO_97 (O_97,N_14915,N_14918);
nor UO_98 (O_98,N_14961,N_14910);
nand UO_99 (O_99,N_14985,N_14978);
nor UO_100 (O_100,N_14922,N_14983);
nand UO_101 (O_101,N_14880,N_14897);
xor UO_102 (O_102,N_14971,N_14909);
nor UO_103 (O_103,N_14973,N_14934);
nor UO_104 (O_104,N_14993,N_14919);
and UO_105 (O_105,N_14998,N_14952);
xor UO_106 (O_106,N_14943,N_14920);
xor UO_107 (O_107,N_14987,N_14973);
nor UO_108 (O_108,N_14882,N_14990);
or UO_109 (O_109,N_14980,N_14923);
nand UO_110 (O_110,N_14897,N_14999);
nand UO_111 (O_111,N_14995,N_14898);
xnor UO_112 (O_112,N_14885,N_14918);
nor UO_113 (O_113,N_14932,N_14875);
nor UO_114 (O_114,N_14903,N_14915);
and UO_115 (O_115,N_14968,N_14880);
nor UO_116 (O_116,N_14970,N_14909);
xnor UO_117 (O_117,N_14879,N_14906);
nand UO_118 (O_118,N_14935,N_14956);
and UO_119 (O_119,N_14887,N_14910);
and UO_120 (O_120,N_14923,N_14881);
xnor UO_121 (O_121,N_14897,N_14895);
or UO_122 (O_122,N_14981,N_14998);
nand UO_123 (O_123,N_14996,N_14897);
nor UO_124 (O_124,N_14901,N_14908);
nand UO_125 (O_125,N_14929,N_14915);
nand UO_126 (O_126,N_14882,N_14886);
and UO_127 (O_127,N_14894,N_14978);
nand UO_128 (O_128,N_14935,N_14907);
xnor UO_129 (O_129,N_14952,N_14928);
nor UO_130 (O_130,N_14898,N_14900);
xnor UO_131 (O_131,N_14957,N_14969);
or UO_132 (O_132,N_14889,N_14983);
xor UO_133 (O_133,N_14936,N_14966);
or UO_134 (O_134,N_14954,N_14923);
nor UO_135 (O_135,N_14958,N_14885);
nand UO_136 (O_136,N_14934,N_14937);
nand UO_137 (O_137,N_14882,N_14993);
and UO_138 (O_138,N_14877,N_14974);
nor UO_139 (O_139,N_14898,N_14923);
xnor UO_140 (O_140,N_14977,N_14886);
nor UO_141 (O_141,N_14995,N_14975);
xnor UO_142 (O_142,N_14892,N_14997);
nand UO_143 (O_143,N_14878,N_14940);
nor UO_144 (O_144,N_14936,N_14911);
nor UO_145 (O_145,N_14939,N_14964);
nand UO_146 (O_146,N_14979,N_14899);
or UO_147 (O_147,N_14996,N_14931);
and UO_148 (O_148,N_14955,N_14883);
and UO_149 (O_149,N_14889,N_14906);
nor UO_150 (O_150,N_14945,N_14974);
or UO_151 (O_151,N_14981,N_14987);
or UO_152 (O_152,N_14964,N_14998);
and UO_153 (O_153,N_14916,N_14976);
xor UO_154 (O_154,N_14900,N_14930);
and UO_155 (O_155,N_14907,N_14877);
xnor UO_156 (O_156,N_14984,N_14975);
and UO_157 (O_157,N_14893,N_14926);
and UO_158 (O_158,N_14998,N_14875);
nor UO_159 (O_159,N_14962,N_14928);
xnor UO_160 (O_160,N_14922,N_14979);
nor UO_161 (O_161,N_14893,N_14911);
xor UO_162 (O_162,N_14882,N_14973);
nor UO_163 (O_163,N_14898,N_14983);
xor UO_164 (O_164,N_14979,N_14934);
nand UO_165 (O_165,N_14891,N_14926);
or UO_166 (O_166,N_14891,N_14887);
nor UO_167 (O_167,N_14920,N_14905);
or UO_168 (O_168,N_14950,N_14923);
xnor UO_169 (O_169,N_14926,N_14964);
and UO_170 (O_170,N_14878,N_14891);
nor UO_171 (O_171,N_14877,N_14900);
xor UO_172 (O_172,N_14967,N_14997);
or UO_173 (O_173,N_14943,N_14902);
nor UO_174 (O_174,N_14886,N_14972);
or UO_175 (O_175,N_14899,N_14926);
xor UO_176 (O_176,N_14900,N_14951);
nor UO_177 (O_177,N_14915,N_14961);
nand UO_178 (O_178,N_14891,N_14935);
or UO_179 (O_179,N_14983,N_14969);
and UO_180 (O_180,N_14880,N_14921);
nor UO_181 (O_181,N_14990,N_14928);
xnor UO_182 (O_182,N_14956,N_14996);
or UO_183 (O_183,N_14898,N_14958);
or UO_184 (O_184,N_14924,N_14878);
xor UO_185 (O_185,N_14979,N_14982);
or UO_186 (O_186,N_14913,N_14905);
and UO_187 (O_187,N_14990,N_14959);
and UO_188 (O_188,N_14976,N_14908);
or UO_189 (O_189,N_14952,N_14897);
and UO_190 (O_190,N_14881,N_14996);
or UO_191 (O_191,N_14912,N_14937);
or UO_192 (O_192,N_14940,N_14990);
and UO_193 (O_193,N_14946,N_14948);
nand UO_194 (O_194,N_14977,N_14878);
nand UO_195 (O_195,N_14935,N_14883);
xnor UO_196 (O_196,N_14973,N_14899);
and UO_197 (O_197,N_14881,N_14941);
nand UO_198 (O_198,N_14883,N_14905);
nand UO_199 (O_199,N_14943,N_14936);
nor UO_200 (O_200,N_14958,N_14914);
xnor UO_201 (O_201,N_14934,N_14989);
xnor UO_202 (O_202,N_14913,N_14962);
nand UO_203 (O_203,N_14900,N_14907);
or UO_204 (O_204,N_14885,N_14985);
and UO_205 (O_205,N_14918,N_14971);
xnor UO_206 (O_206,N_14919,N_14960);
nand UO_207 (O_207,N_14957,N_14901);
xor UO_208 (O_208,N_14944,N_14895);
nor UO_209 (O_209,N_14927,N_14883);
nor UO_210 (O_210,N_14936,N_14877);
or UO_211 (O_211,N_14943,N_14963);
or UO_212 (O_212,N_14876,N_14881);
and UO_213 (O_213,N_14876,N_14978);
nor UO_214 (O_214,N_14905,N_14929);
and UO_215 (O_215,N_14964,N_14925);
nor UO_216 (O_216,N_14970,N_14887);
or UO_217 (O_217,N_14939,N_14904);
and UO_218 (O_218,N_14993,N_14924);
and UO_219 (O_219,N_14944,N_14982);
nor UO_220 (O_220,N_14910,N_14946);
xor UO_221 (O_221,N_14982,N_14891);
nand UO_222 (O_222,N_14925,N_14875);
xnor UO_223 (O_223,N_14931,N_14921);
nand UO_224 (O_224,N_14988,N_14882);
xnor UO_225 (O_225,N_14959,N_14885);
or UO_226 (O_226,N_14920,N_14938);
and UO_227 (O_227,N_14878,N_14974);
nor UO_228 (O_228,N_14939,N_14986);
or UO_229 (O_229,N_14991,N_14944);
nor UO_230 (O_230,N_14922,N_14902);
and UO_231 (O_231,N_14998,N_14885);
xnor UO_232 (O_232,N_14890,N_14951);
and UO_233 (O_233,N_14950,N_14970);
and UO_234 (O_234,N_14901,N_14879);
xnor UO_235 (O_235,N_14957,N_14984);
nor UO_236 (O_236,N_14945,N_14953);
nor UO_237 (O_237,N_14934,N_14995);
or UO_238 (O_238,N_14995,N_14925);
nor UO_239 (O_239,N_14896,N_14911);
and UO_240 (O_240,N_14974,N_14936);
nand UO_241 (O_241,N_14924,N_14996);
nor UO_242 (O_242,N_14924,N_14998);
and UO_243 (O_243,N_14901,N_14932);
nand UO_244 (O_244,N_14958,N_14899);
and UO_245 (O_245,N_14974,N_14968);
and UO_246 (O_246,N_14907,N_14955);
nand UO_247 (O_247,N_14963,N_14946);
nor UO_248 (O_248,N_14955,N_14994);
xor UO_249 (O_249,N_14919,N_14894);
nand UO_250 (O_250,N_14927,N_14923);
xor UO_251 (O_251,N_14955,N_14995);
and UO_252 (O_252,N_14902,N_14951);
or UO_253 (O_253,N_14956,N_14925);
and UO_254 (O_254,N_14906,N_14877);
and UO_255 (O_255,N_14950,N_14977);
and UO_256 (O_256,N_14944,N_14967);
or UO_257 (O_257,N_14927,N_14996);
nor UO_258 (O_258,N_14995,N_14913);
nor UO_259 (O_259,N_14958,N_14937);
nor UO_260 (O_260,N_14947,N_14887);
xor UO_261 (O_261,N_14963,N_14949);
or UO_262 (O_262,N_14975,N_14889);
nor UO_263 (O_263,N_14875,N_14939);
nor UO_264 (O_264,N_14956,N_14954);
or UO_265 (O_265,N_14953,N_14915);
nor UO_266 (O_266,N_14992,N_14909);
and UO_267 (O_267,N_14947,N_14884);
xor UO_268 (O_268,N_14975,N_14916);
nor UO_269 (O_269,N_14921,N_14908);
nand UO_270 (O_270,N_14898,N_14924);
or UO_271 (O_271,N_14922,N_14908);
or UO_272 (O_272,N_14974,N_14914);
or UO_273 (O_273,N_14924,N_14901);
nor UO_274 (O_274,N_14965,N_14936);
nor UO_275 (O_275,N_14924,N_14980);
and UO_276 (O_276,N_14961,N_14914);
xnor UO_277 (O_277,N_14971,N_14892);
xor UO_278 (O_278,N_14977,N_14962);
nor UO_279 (O_279,N_14998,N_14890);
nor UO_280 (O_280,N_14955,N_14898);
or UO_281 (O_281,N_14995,N_14921);
xnor UO_282 (O_282,N_14959,N_14943);
or UO_283 (O_283,N_14920,N_14946);
and UO_284 (O_284,N_14974,N_14889);
nor UO_285 (O_285,N_14938,N_14925);
xnor UO_286 (O_286,N_14940,N_14985);
or UO_287 (O_287,N_14940,N_14879);
nor UO_288 (O_288,N_14962,N_14999);
xor UO_289 (O_289,N_14898,N_14992);
nor UO_290 (O_290,N_14988,N_14936);
nor UO_291 (O_291,N_14885,N_14929);
and UO_292 (O_292,N_14919,N_14955);
nor UO_293 (O_293,N_14964,N_14962);
nand UO_294 (O_294,N_14920,N_14966);
nor UO_295 (O_295,N_14927,N_14898);
xor UO_296 (O_296,N_14923,N_14935);
or UO_297 (O_297,N_14924,N_14995);
nand UO_298 (O_298,N_14952,N_14990);
xnor UO_299 (O_299,N_14981,N_14920);
nand UO_300 (O_300,N_14991,N_14905);
or UO_301 (O_301,N_14906,N_14959);
xnor UO_302 (O_302,N_14891,N_14924);
xor UO_303 (O_303,N_14928,N_14902);
and UO_304 (O_304,N_14943,N_14931);
or UO_305 (O_305,N_14967,N_14981);
xnor UO_306 (O_306,N_14939,N_14929);
or UO_307 (O_307,N_14957,N_14917);
nand UO_308 (O_308,N_14930,N_14944);
or UO_309 (O_309,N_14960,N_14938);
or UO_310 (O_310,N_14982,N_14905);
and UO_311 (O_311,N_14960,N_14884);
nand UO_312 (O_312,N_14896,N_14987);
nor UO_313 (O_313,N_14927,N_14924);
nand UO_314 (O_314,N_14984,N_14911);
nand UO_315 (O_315,N_14936,N_14918);
nor UO_316 (O_316,N_14910,N_14990);
xor UO_317 (O_317,N_14948,N_14950);
and UO_318 (O_318,N_14909,N_14877);
nor UO_319 (O_319,N_14893,N_14966);
nor UO_320 (O_320,N_14992,N_14947);
nand UO_321 (O_321,N_14943,N_14925);
nor UO_322 (O_322,N_14886,N_14936);
xnor UO_323 (O_323,N_14914,N_14948);
nor UO_324 (O_324,N_14909,N_14879);
xor UO_325 (O_325,N_14896,N_14976);
and UO_326 (O_326,N_14882,N_14889);
nor UO_327 (O_327,N_14942,N_14928);
and UO_328 (O_328,N_14979,N_14967);
nand UO_329 (O_329,N_14917,N_14934);
nor UO_330 (O_330,N_14925,N_14915);
and UO_331 (O_331,N_14987,N_14893);
and UO_332 (O_332,N_14943,N_14878);
or UO_333 (O_333,N_14948,N_14894);
nand UO_334 (O_334,N_14981,N_14914);
nor UO_335 (O_335,N_14948,N_14932);
nand UO_336 (O_336,N_14916,N_14891);
nand UO_337 (O_337,N_14948,N_14944);
and UO_338 (O_338,N_14936,N_14987);
or UO_339 (O_339,N_14981,N_14915);
nand UO_340 (O_340,N_14902,N_14954);
or UO_341 (O_341,N_14958,N_14941);
nor UO_342 (O_342,N_14979,N_14970);
nand UO_343 (O_343,N_14907,N_14890);
or UO_344 (O_344,N_14959,N_14896);
and UO_345 (O_345,N_14915,N_14993);
nand UO_346 (O_346,N_14905,N_14985);
nand UO_347 (O_347,N_14957,N_14928);
or UO_348 (O_348,N_14966,N_14887);
xnor UO_349 (O_349,N_14886,N_14887);
and UO_350 (O_350,N_14978,N_14972);
nand UO_351 (O_351,N_14907,N_14966);
xor UO_352 (O_352,N_14890,N_14937);
or UO_353 (O_353,N_14987,N_14926);
nand UO_354 (O_354,N_14920,N_14881);
nor UO_355 (O_355,N_14985,N_14936);
or UO_356 (O_356,N_14990,N_14895);
xnor UO_357 (O_357,N_14944,N_14886);
nand UO_358 (O_358,N_14966,N_14969);
nand UO_359 (O_359,N_14886,N_14885);
nor UO_360 (O_360,N_14991,N_14881);
nor UO_361 (O_361,N_14909,N_14939);
nor UO_362 (O_362,N_14973,N_14944);
nor UO_363 (O_363,N_14973,N_14908);
nand UO_364 (O_364,N_14966,N_14997);
nand UO_365 (O_365,N_14895,N_14948);
or UO_366 (O_366,N_14892,N_14911);
or UO_367 (O_367,N_14959,N_14917);
nor UO_368 (O_368,N_14897,N_14944);
xnor UO_369 (O_369,N_14916,N_14960);
and UO_370 (O_370,N_14921,N_14946);
and UO_371 (O_371,N_14971,N_14967);
or UO_372 (O_372,N_14960,N_14891);
or UO_373 (O_373,N_14933,N_14997);
and UO_374 (O_374,N_14952,N_14888);
xnor UO_375 (O_375,N_14890,N_14909);
or UO_376 (O_376,N_14890,N_14961);
xor UO_377 (O_377,N_14887,N_14994);
and UO_378 (O_378,N_14996,N_14883);
nand UO_379 (O_379,N_14955,N_14904);
or UO_380 (O_380,N_14966,N_14882);
nand UO_381 (O_381,N_14935,N_14980);
and UO_382 (O_382,N_14970,N_14905);
nor UO_383 (O_383,N_14923,N_14983);
xor UO_384 (O_384,N_14944,N_14912);
or UO_385 (O_385,N_14952,N_14931);
xnor UO_386 (O_386,N_14983,N_14974);
xor UO_387 (O_387,N_14936,N_14954);
and UO_388 (O_388,N_14890,N_14901);
or UO_389 (O_389,N_14959,N_14972);
or UO_390 (O_390,N_14915,N_14946);
nand UO_391 (O_391,N_14980,N_14999);
or UO_392 (O_392,N_14901,N_14887);
and UO_393 (O_393,N_14968,N_14892);
and UO_394 (O_394,N_14951,N_14880);
nand UO_395 (O_395,N_14968,N_14910);
nor UO_396 (O_396,N_14885,N_14903);
and UO_397 (O_397,N_14997,N_14964);
or UO_398 (O_398,N_14943,N_14945);
nor UO_399 (O_399,N_14953,N_14973);
or UO_400 (O_400,N_14954,N_14990);
nor UO_401 (O_401,N_14915,N_14917);
and UO_402 (O_402,N_14971,N_14999);
nor UO_403 (O_403,N_14996,N_14950);
or UO_404 (O_404,N_14922,N_14937);
nand UO_405 (O_405,N_14981,N_14882);
or UO_406 (O_406,N_14929,N_14942);
nand UO_407 (O_407,N_14912,N_14907);
nor UO_408 (O_408,N_14943,N_14986);
or UO_409 (O_409,N_14998,N_14990);
or UO_410 (O_410,N_14878,N_14991);
nand UO_411 (O_411,N_14996,N_14964);
xnor UO_412 (O_412,N_14940,N_14986);
and UO_413 (O_413,N_14940,N_14944);
or UO_414 (O_414,N_14892,N_14951);
xor UO_415 (O_415,N_14925,N_14979);
and UO_416 (O_416,N_14941,N_14882);
xnor UO_417 (O_417,N_14887,N_14895);
xor UO_418 (O_418,N_14923,N_14971);
xor UO_419 (O_419,N_14883,N_14895);
nand UO_420 (O_420,N_14984,N_14900);
or UO_421 (O_421,N_14932,N_14981);
or UO_422 (O_422,N_14926,N_14929);
xnor UO_423 (O_423,N_14924,N_14950);
nand UO_424 (O_424,N_14923,N_14968);
and UO_425 (O_425,N_14956,N_14957);
nor UO_426 (O_426,N_14941,N_14901);
nand UO_427 (O_427,N_14878,N_14915);
nand UO_428 (O_428,N_14882,N_14914);
nand UO_429 (O_429,N_14970,N_14916);
or UO_430 (O_430,N_14978,N_14944);
xor UO_431 (O_431,N_14901,N_14954);
nor UO_432 (O_432,N_14896,N_14928);
or UO_433 (O_433,N_14911,N_14975);
nor UO_434 (O_434,N_14944,N_14955);
nor UO_435 (O_435,N_14986,N_14976);
nor UO_436 (O_436,N_14983,N_14892);
nor UO_437 (O_437,N_14879,N_14908);
xnor UO_438 (O_438,N_14985,N_14901);
nor UO_439 (O_439,N_14920,N_14909);
xor UO_440 (O_440,N_14919,N_14942);
nor UO_441 (O_441,N_14947,N_14879);
xor UO_442 (O_442,N_14891,N_14880);
and UO_443 (O_443,N_14914,N_14909);
nand UO_444 (O_444,N_14941,N_14924);
and UO_445 (O_445,N_14925,N_14883);
or UO_446 (O_446,N_14894,N_14981);
nor UO_447 (O_447,N_14901,N_14917);
nor UO_448 (O_448,N_14888,N_14948);
or UO_449 (O_449,N_14916,N_14947);
nand UO_450 (O_450,N_14942,N_14898);
nand UO_451 (O_451,N_14994,N_14925);
xor UO_452 (O_452,N_14945,N_14891);
xor UO_453 (O_453,N_14996,N_14887);
nor UO_454 (O_454,N_14893,N_14994);
and UO_455 (O_455,N_14960,N_14899);
xnor UO_456 (O_456,N_14986,N_14995);
nand UO_457 (O_457,N_14954,N_14881);
and UO_458 (O_458,N_14949,N_14918);
nand UO_459 (O_459,N_14902,N_14879);
xor UO_460 (O_460,N_14921,N_14964);
or UO_461 (O_461,N_14960,N_14994);
nand UO_462 (O_462,N_14967,N_14949);
or UO_463 (O_463,N_14949,N_14990);
xor UO_464 (O_464,N_14959,N_14999);
and UO_465 (O_465,N_14983,N_14964);
or UO_466 (O_466,N_14948,N_14929);
and UO_467 (O_467,N_14992,N_14982);
and UO_468 (O_468,N_14958,N_14903);
and UO_469 (O_469,N_14927,N_14942);
xnor UO_470 (O_470,N_14923,N_14945);
and UO_471 (O_471,N_14996,N_14946);
xnor UO_472 (O_472,N_14897,N_14979);
nand UO_473 (O_473,N_14911,N_14876);
nand UO_474 (O_474,N_14959,N_14928);
nor UO_475 (O_475,N_14900,N_14931);
and UO_476 (O_476,N_14977,N_14941);
xnor UO_477 (O_477,N_14895,N_14911);
xnor UO_478 (O_478,N_14929,N_14938);
xor UO_479 (O_479,N_14882,N_14989);
xnor UO_480 (O_480,N_14981,N_14892);
and UO_481 (O_481,N_14904,N_14949);
xnor UO_482 (O_482,N_14904,N_14896);
nand UO_483 (O_483,N_14953,N_14963);
and UO_484 (O_484,N_14909,N_14896);
nand UO_485 (O_485,N_14978,N_14892);
xor UO_486 (O_486,N_14988,N_14917);
xor UO_487 (O_487,N_14903,N_14881);
xor UO_488 (O_488,N_14892,N_14930);
or UO_489 (O_489,N_14990,N_14936);
nand UO_490 (O_490,N_14878,N_14926);
or UO_491 (O_491,N_14918,N_14907);
nor UO_492 (O_492,N_14941,N_14940);
xor UO_493 (O_493,N_14947,N_14929);
xnor UO_494 (O_494,N_14922,N_14928);
xnor UO_495 (O_495,N_14989,N_14953);
xnor UO_496 (O_496,N_14884,N_14998);
or UO_497 (O_497,N_14976,N_14990);
xnor UO_498 (O_498,N_14999,N_14889);
xor UO_499 (O_499,N_14953,N_14954);
nor UO_500 (O_500,N_14957,N_14909);
xnor UO_501 (O_501,N_14955,N_14916);
or UO_502 (O_502,N_14941,N_14975);
nor UO_503 (O_503,N_14900,N_14954);
or UO_504 (O_504,N_14909,N_14933);
or UO_505 (O_505,N_14891,N_14993);
or UO_506 (O_506,N_14969,N_14960);
nand UO_507 (O_507,N_14883,N_14924);
xnor UO_508 (O_508,N_14899,N_14879);
nand UO_509 (O_509,N_14969,N_14885);
nand UO_510 (O_510,N_14978,N_14907);
nor UO_511 (O_511,N_14955,N_14947);
xor UO_512 (O_512,N_14895,N_14884);
or UO_513 (O_513,N_14965,N_14898);
nor UO_514 (O_514,N_14980,N_14986);
or UO_515 (O_515,N_14879,N_14917);
nor UO_516 (O_516,N_14928,N_14991);
or UO_517 (O_517,N_14999,N_14992);
nand UO_518 (O_518,N_14922,N_14959);
xor UO_519 (O_519,N_14981,N_14959);
or UO_520 (O_520,N_14921,N_14976);
xnor UO_521 (O_521,N_14994,N_14892);
xnor UO_522 (O_522,N_14942,N_14973);
nand UO_523 (O_523,N_14887,N_14933);
nor UO_524 (O_524,N_14914,N_14902);
nand UO_525 (O_525,N_14964,N_14912);
nor UO_526 (O_526,N_14877,N_14982);
nor UO_527 (O_527,N_14928,N_14935);
xor UO_528 (O_528,N_14999,N_14894);
or UO_529 (O_529,N_14918,N_14961);
nand UO_530 (O_530,N_14963,N_14875);
nand UO_531 (O_531,N_14979,N_14972);
or UO_532 (O_532,N_14931,N_14993);
nand UO_533 (O_533,N_14897,N_14883);
nand UO_534 (O_534,N_14934,N_14911);
or UO_535 (O_535,N_14955,N_14960);
and UO_536 (O_536,N_14976,N_14968);
or UO_537 (O_537,N_14879,N_14935);
nand UO_538 (O_538,N_14966,N_14914);
and UO_539 (O_539,N_14959,N_14888);
or UO_540 (O_540,N_14890,N_14976);
and UO_541 (O_541,N_14921,N_14977);
nand UO_542 (O_542,N_14913,N_14992);
or UO_543 (O_543,N_14972,N_14974);
nand UO_544 (O_544,N_14970,N_14888);
and UO_545 (O_545,N_14943,N_14897);
or UO_546 (O_546,N_14992,N_14908);
nand UO_547 (O_547,N_14917,N_14966);
nor UO_548 (O_548,N_14964,N_14988);
nand UO_549 (O_549,N_14884,N_14964);
and UO_550 (O_550,N_14991,N_14926);
nor UO_551 (O_551,N_14964,N_14876);
nand UO_552 (O_552,N_14889,N_14925);
xor UO_553 (O_553,N_14990,N_14993);
or UO_554 (O_554,N_14997,N_14940);
nand UO_555 (O_555,N_14991,N_14986);
or UO_556 (O_556,N_14938,N_14936);
nor UO_557 (O_557,N_14937,N_14969);
xor UO_558 (O_558,N_14986,N_14993);
xor UO_559 (O_559,N_14905,N_14939);
nand UO_560 (O_560,N_14961,N_14977);
nand UO_561 (O_561,N_14998,N_14938);
nor UO_562 (O_562,N_14966,N_14886);
nand UO_563 (O_563,N_14943,N_14998);
nand UO_564 (O_564,N_14943,N_14996);
xor UO_565 (O_565,N_14957,N_14878);
nor UO_566 (O_566,N_14998,N_14927);
or UO_567 (O_567,N_14889,N_14945);
and UO_568 (O_568,N_14881,N_14905);
nor UO_569 (O_569,N_14887,N_14955);
nor UO_570 (O_570,N_14901,N_14905);
nand UO_571 (O_571,N_14916,N_14935);
and UO_572 (O_572,N_14908,N_14913);
xnor UO_573 (O_573,N_14924,N_14965);
or UO_574 (O_574,N_14934,N_14935);
xor UO_575 (O_575,N_14971,N_14933);
nor UO_576 (O_576,N_14916,N_14988);
nor UO_577 (O_577,N_14915,N_14877);
or UO_578 (O_578,N_14914,N_14946);
xor UO_579 (O_579,N_14912,N_14946);
xor UO_580 (O_580,N_14954,N_14913);
nand UO_581 (O_581,N_14925,N_14983);
nand UO_582 (O_582,N_14945,N_14881);
and UO_583 (O_583,N_14980,N_14964);
xnor UO_584 (O_584,N_14876,N_14961);
and UO_585 (O_585,N_14960,N_14929);
or UO_586 (O_586,N_14915,N_14911);
nor UO_587 (O_587,N_14896,N_14900);
or UO_588 (O_588,N_14884,N_14885);
or UO_589 (O_589,N_14932,N_14942);
or UO_590 (O_590,N_14994,N_14952);
xnor UO_591 (O_591,N_14897,N_14992);
or UO_592 (O_592,N_14875,N_14934);
or UO_593 (O_593,N_14966,N_14921);
xnor UO_594 (O_594,N_14929,N_14877);
nor UO_595 (O_595,N_14920,N_14944);
xnor UO_596 (O_596,N_14952,N_14937);
or UO_597 (O_597,N_14953,N_14959);
and UO_598 (O_598,N_14935,N_14925);
xnor UO_599 (O_599,N_14915,N_14932);
nand UO_600 (O_600,N_14929,N_14930);
or UO_601 (O_601,N_14940,N_14979);
nor UO_602 (O_602,N_14983,N_14989);
or UO_603 (O_603,N_14919,N_14906);
or UO_604 (O_604,N_14993,N_14975);
xnor UO_605 (O_605,N_14952,N_14956);
nand UO_606 (O_606,N_14876,N_14896);
xnor UO_607 (O_607,N_14971,N_14982);
nor UO_608 (O_608,N_14970,N_14920);
nor UO_609 (O_609,N_14914,N_14890);
nand UO_610 (O_610,N_14928,N_14999);
nand UO_611 (O_611,N_14893,N_14971);
nand UO_612 (O_612,N_14878,N_14986);
xnor UO_613 (O_613,N_14997,N_14878);
nand UO_614 (O_614,N_14907,N_14928);
nand UO_615 (O_615,N_14914,N_14979);
and UO_616 (O_616,N_14945,N_14998);
nand UO_617 (O_617,N_14935,N_14932);
and UO_618 (O_618,N_14974,N_14955);
xnor UO_619 (O_619,N_14884,N_14951);
nor UO_620 (O_620,N_14980,N_14896);
nor UO_621 (O_621,N_14921,N_14889);
nor UO_622 (O_622,N_14920,N_14993);
xor UO_623 (O_623,N_14897,N_14960);
nand UO_624 (O_624,N_14968,N_14969);
or UO_625 (O_625,N_14961,N_14886);
or UO_626 (O_626,N_14958,N_14882);
nand UO_627 (O_627,N_14901,N_14923);
or UO_628 (O_628,N_14921,N_14982);
nand UO_629 (O_629,N_14978,N_14965);
or UO_630 (O_630,N_14988,N_14883);
nor UO_631 (O_631,N_14893,N_14922);
nand UO_632 (O_632,N_14999,N_14877);
xor UO_633 (O_633,N_14958,N_14994);
xor UO_634 (O_634,N_14975,N_14992);
nor UO_635 (O_635,N_14933,N_14984);
nor UO_636 (O_636,N_14888,N_14914);
and UO_637 (O_637,N_14990,N_14968);
nand UO_638 (O_638,N_14991,N_14893);
and UO_639 (O_639,N_14979,N_14951);
and UO_640 (O_640,N_14945,N_14902);
xnor UO_641 (O_641,N_14914,N_14920);
xor UO_642 (O_642,N_14949,N_14919);
and UO_643 (O_643,N_14988,N_14908);
nand UO_644 (O_644,N_14923,N_14948);
nand UO_645 (O_645,N_14971,N_14884);
nand UO_646 (O_646,N_14918,N_14920);
nor UO_647 (O_647,N_14990,N_14884);
nor UO_648 (O_648,N_14898,N_14926);
or UO_649 (O_649,N_14910,N_14976);
or UO_650 (O_650,N_14971,N_14885);
xor UO_651 (O_651,N_14989,N_14945);
and UO_652 (O_652,N_14881,N_14937);
and UO_653 (O_653,N_14884,N_14972);
or UO_654 (O_654,N_14922,N_14995);
xnor UO_655 (O_655,N_14897,N_14910);
and UO_656 (O_656,N_14979,N_14905);
xor UO_657 (O_657,N_14960,N_14885);
nand UO_658 (O_658,N_14900,N_14976);
nor UO_659 (O_659,N_14885,N_14954);
xor UO_660 (O_660,N_14890,N_14943);
nor UO_661 (O_661,N_14938,N_14979);
nand UO_662 (O_662,N_14887,N_14937);
and UO_663 (O_663,N_14934,N_14893);
or UO_664 (O_664,N_14980,N_14977);
or UO_665 (O_665,N_14999,N_14932);
and UO_666 (O_666,N_14922,N_14986);
xor UO_667 (O_667,N_14927,N_14943);
nor UO_668 (O_668,N_14943,N_14974);
xor UO_669 (O_669,N_14948,N_14884);
and UO_670 (O_670,N_14957,N_14875);
nor UO_671 (O_671,N_14976,N_14901);
and UO_672 (O_672,N_14920,N_14932);
and UO_673 (O_673,N_14978,N_14923);
and UO_674 (O_674,N_14878,N_14934);
nand UO_675 (O_675,N_14986,N_14973);
and UO_676 (O_676,N_14973,N_14877);
or UO_677 (O_677,N_14951,N_14988);
nor UO_678 (O_678,N_14953,N_14925);
nand UO_679 (O_679,N_14958,N_14952);
or UO_680 (O_680,N_14960,N_14987);
nand UO_681 (O_681,N_14927,N_14901);
or UO_682 (O_682,N_14988,N_14893);
xnor UO_683 (O_683,N_14891,N_14931);
and UO_684 (O_684,N_14989,N_14888);
or UO_685 (O_685,N_14959,N_14919);
nor UO_686 (O_686,N_14935,N_14993);
or UO_687 (O_687,N_14937,N_14907);
or UO_688 (O_688,N_14880,N_14995);
nor UO_689 (O_689,N_14945,N_14968);
or UO_690 (O_690,N_14928,N_14890);
or UO_691 (O_691,N_14918,N_14990);
or UO_692 (O_692,N_14887,N_14903);
nor UO_693 (O_693,N_14915,N_14979);
and UO_694 (O_694,N_14945,N_14886);
nand UO_695 (O_695,N_14928,N_14911);
or UO_696 (O_696,N_14978,N_14947);
nand UO_697 (O_697,N_14928,N_14973);
nand UO_698 (O_698,N_14964,N_14935);
nand UO_699 (O_699,N_14949,N_14923);
nor UO_700 (O_700,N_14985,N_14948);
nand UO_701 (O_701,N_14966,N_14967);
nand UO_702 (O_702,N_14879,N_14963);
nand UO_703 (O_703,N_14994,N_14957);
nand UO_704 (O_704,N_14928,N_14905);
or UO_705 (O_705,N_14948,N_14986);
and UO_706 (O_706,N_14897,N_14902);
and UO_707 (O_707,N_14878,N_14944);
and UO_708 (O_708,N_14999,N_14979);
and UO_709 (O_709,N_14902,N_14895);
nand UO_710 (O_710,N_14975,N_14971);
or UO_711 (O_711,N_14966,N_14982);
xnor UO_712 (O_712,N_14966,N_14877);
nor UO_713 (O_713,N_14950,N_14908);
or UO_714 (O_714,N_14934,N_14952);
and UO_715 (O_715,N_14981,N_14930);
or UO_716 (O_716,N_14975,N_14974);
nand UO_717 (O_717,N_14978,N_14936);
xor UO_718 (O_718,N_14973,N_14965);
xor UO_719 (O_719,N_14919,N_14913);
xor UO_720 (O_720,N_14926,N_14995);
nor UO_721 (O_721,N_14972,N_14945);
nand UO_722 (O_722,N_14896,N_14964);
nand UO_723 (O_723,N_14882,N_14951);
xor UO_724 (O_724,N_14994,N_14986);
xor UO_725 (O_725,N_14992,N_14921);
and UO_726 (O_726,N_14939,N_14982);
and UO_727 (O_727,N_14996,N_14906);
xnor UO_728 (O_728,N_14958,N_14955);
nand UO_729 (O_729,N_14955,N_14914);
and UO_730 (O_730,N_14981,N_14891);
nand UO_731 (O_731,N_14968,N_14998);
xor UO_732 (O_732,N_14994,N_14932);
xor UO_733 (O_733,N_14904,N_14888);
xnor UO_734 (O_734,N_14887,N_14876);
nor UO_735 (O_735,N_14949,N_14940);
xor UO_736 (O_736,N_14907,N_14959);
nor UO_737 (O_737,N_14951,N_14898);
or UO_738 (O_738,N_14916,N_14920);
or UO_739 (O_739,N_14884,N_14969);
and UO_740 (O_740,N_14889,N_14963);
or UO_741 (O_741,N_14983,N_14913);
xor UO_742 (O_742,N_14963,N_14974);
and UO_743 (O_743,N_14916,N_14980);
xor UO_744 (O_744,N_14967,N_14924);
nor UO_745 (O_745,N_14957,N_14886);
and UO_746 (O_746,N_14948,N_14916);
or UO_747 (O_747,N_14937,N_14999);
xor UO_748 (O_748,N_14985,N_14875);
and UO_749 (O_749,N_14994,N_14976);
xor UO_750 (O_750,N_14979,N_14963);
and UO_751 (O_751,N_14998,N_14911);
xnor UO_752 (O_752,N_14946,N_14940);
nor UO_753 (O_753,N_14968,N_14951);
nand UO_754 (O_754,N_14875,N_14883);
nand UO_755 (O_755,N_14986,N_14985);
nand UO_756 (O_756,N_14876,N_14894);
nor UO_757 (O_757,N_14882,N_14899);
xnor UO_758 (O_758,N_14981,N_14951);
and UO_759 (O_759,N_14955,N_14875);
or UO_760 (O_760,N_14888,N_14971);
or UO_761 (O_761,N_14901,N_14937);
xnor UO_762 (O_762,N_14933,N_14912);
and UO_763 (O_763,N_14876,N_14982);
nand UO_764 (O_764,N_14902,N_14933);
and UO_765 (O_765,N_14959,N_14931);
nand UO_766 (O_766,N_14991,N_14983);
and UO_767 (O_767,N_14925,N_14976);
xnor UO_768 (O_768,N_14905,N_14897);
or UO_769 (O_769,N_14920,N_14995);
nor UO_770 (O_770,N_14918,N_14930);
or UO_771 (O_771,N_14875,N_14961);
or UO_772 (O_772,N_14929,N_14976);
xor UO_773 (O_773,N_14997,N_14882);
or UO_774 (O_774,N_14968,N_14953);
or UO_775 (O_775,N_14902,N_14996);
nor UO_776 (O_776,N_14965,N_14985);
xnor UO_777 (O_777,N_14887,N_14951);
or UO_778 (O_778,N_14985,N_14912);
or UO_779 (O_779,N_14887,N_14923);
and UO_780 (O_780,N_14927,N_14955);
xnor UO_781 (O_781,N_14973,N_14959);
xnor UO_782 (O_782,N_14904,N_14962);
nand UO_783 (O_783,N_14894,N_14995);
nor UO_784 (O_784,N_14890,N_14989);
or UO_785 (O_785,N_14898,N_14939);
nand UO_786 (O_786,N_14989,N_14893);
and UO_787 (O_787,N_14985,N_14951);
xor UO_788 (O_788,N_14908,N_14914);
or UO_789 (O_789,N_14978,N_14975);
xor UO_790 (O_790,N_14890,N_14965);
xnor UO_791 (O_791,N_14922,N_14949);
nor UO_792 (O_792,N_14944,N_14989);
nor UO_793 (O_793,N_14907,N_14936);
nand UO_794 (O_794,N_14916,N_14929);
nand UO_795 (O_795,N_14947,N_14892);
and UO_796 (O_796,N_14973,N_14946);
nor UO_797 (O_797,N_14950,N_14903);
nor UO_798 (O_798,N_14969,N_14875);
xnor UO_799 (O_799,N_14958,N_14925);
nand UO_800 (O_800,N_14898,N_14974);
nand UO_801 (O_801,N_14989,N_14936);
or UO_802 (O_802,N_14906,N_14927);
and UO_803 (O_803,N_14943,N_14918);
nand UO_804 (O_804,N_14945,N_14962);
or UO_805 (O_805,N_14972,N_14891);
xnor UO_806 (O_806,N_14903,N_14904);
and UO_807 (O_807,N_14891,N_14950);
and UO_808 (O_808,N_14984,N_14919);
xor UO_809 (O_809,N_14956,N_14965);
and UO_810 (O_810,N_14935,N_14933);
and UO_811 (O_811,N_14945,N_14879);
xnor UO_812 (O_812,N_14935,N_14952);
nor UO_813 (O_813,N_14949,N_14978);
nand UO_814 (O_814,N_14942,N_14984);
or UO_815 (O_815,N_14897,N_14970);
nor UO_816 (O_816,N_14977,N_14964);
nand UO_817 (O_817,N_14880,N_14912);
or UO_818 (O_818,N_14982,N_14940);
and UO_819 (O_819,N_14951,N_14942);
xnor UO_820 (O_820,N_14979,N_14880);
or UO_821 (O_821,N_14897,N_14957);
nor UO_822 (O_822,N_14945,N_14977);
or UO_823 (O_823,N_14894,N_14925);
nor UO_824 (O_824,N_14904,N_14934);
nand UO_825 (O_825,N_14889,N_14998);
and UO_826 (O_826,N_14967,N_14887);
nor UO_827 (O_827,N_14902,N_14912);
or UO_828 (O_828,N_14928,N_14951);
or UO_829 (O_829,N_14940,N_14976);
nand UO_830 (O_830,N_14982,N_14930);
xor UO_831 (O_831,N_14984,N_14966);
and UO_832 (O_832,N_14895,N_14940);
xor UO_833 (O_833,N_14952,N_14988);
and UO_834 (O_834,N_14926,N_14930);
nor UO_835 (O_835,N_14988,N_14990);
or UO_836 (O_836,N_14987,N_14991);
nor UO_837 (O_837,N_14963,N_14997);
nand UO_838 (O_838,N_14941,N_14923);
or UO_839 (O_839,N_14881,N_14994);
nor UO_840 (O_840,N_14961,N_14940);
nor UO_841 (O_841,N_14981,N_14895);
xor UO_842 (O_842,N_14882,N_14930);
and UO_843 (O_843,N_14967,N_14895);
and UO_844 (O_844,N_14947,N_14938);
xor UO_845 (O_845,N_14930,N_14978);
nand UO_846 (O_846,N_14936,N_14913);
and UO_847 (O_847,N_14875,N_14897);
and UO_848 (O_848,N_14974,N_14967);
xor UO_849 (O_849,N_14985,N_14989);
nor UO_850 (O_850,N_14939,N_14903);
nand UO_851 (O_851,N_14931,N_14893);
xnor UO_852 (O_852,N_14968,N_14957);
or UO_853 (O_853,N_14982,N_14963);
nor UO_854 (O_854,N_14897,N_14958);
xor UO_855 (O_855,N_14999,N_14975);
nand UO_856 (O_856,N_14896,N_14943);
xnor UO_857 (O_857,N_14925,N_14927);
nand UO_858 (O_858,N_14988,N_14999);
and UO_859 (O_859,N_14931,N_14894);
and UO_860 (O_860,N_14888,N_14886);
nand UO_861 (O_861,N_14943,N_14988);
nor UO_862 (O_862,N_14940,N_14992);
and UO_863 (O_863,N_14943,N_14926);
xor UO_864 (O_864,N_14909,N_14881);
xor UO_865 (O_865,N_14984,N_14938);
nor UO_866 (O_866,N_14926,N_14971);
nand UO_867 (O_867,N_14967,N_14892);
nor UO_868 (O_868,N_14957,N_14936);
or UO_869 (O_869,N_14883,N_14916);
xnor UO_870 (O_870,N_14953,N_14918);
nor UO_871 (O_871,N_14937,N_14886);
nor UO_872 (O_872,N_14932,N_14907);
xor UO_873 (O_873,N_14978,N_14883);
and UO_874 (O_874,N_14961,N_14879);
nand UO_875 (O_875,N_14969,N_14964);
and UO_876 (O_876,N_14908,N_14923);
xnor UO_877 (O_877,N_14875,N_14876);
xnor UO_878 (O_878,N_14944,N_14909);
nor UO_879 (O_879,N_14914,N_14947);
or UO_880 (O_880,N_14919,N_14897);
nor UO_881 (O_881,N_14991,N_14887);
or UO_882 (O_882,N_14958,N_14984);
or UO_883 (O_883,N_14909,N_14910);
or UO_884 (O_884,N_14887,N_14892);
nor UO_885 (O_885,N_14940,N_14994);
xnor UO_886 (O_886,N_14903,N_14897);
nand UO_887 (O_887,N_14995,N_14957);
and UO_888 (O_888,N_14967,N_14945);
nor UO_889 (O_889,N_14892,N_14938);
or UO_890 (O_890,N_14997,N_14962);
nor UO_891 (O_891,N_14895,N_14935);
and UO_892 (O_892,N_14935,N_14887);
nor UO_893 (O_893,N_14990,N_14943);
nand UO_894 (O_894,N_14883,N_14997);
nand UO_895 (O_895,N_14955,N_14899);
or UO_896 (O_896,N_14951,N_14915);
or UO_897 (O_897,N_14889,N_14903);
and UO_898 (O_898,N_14896,N_14932);
nor UO_899 (O_899,N_14961,N_14970);
xor UO_900 (O_900,N_14901,N_14892);
nand UO_901 (O_901,N_14918,N_14934);
and UO_902 (O_902,N_14943,N_14966);
xor UO_903 (O_903,N_14995,N_14883);
nand UO_904 (O_904,N_14945,N_14922);
and UO_905 (O_905,N_14927,N_14899);
nor UO_906 (O_906,N_14958,N_14912);
and UO_907 (O_907,N_14912,N_14896);
nor UO_908 (O_908,N_14909,N_14916);
nor UO_909 (O_909,N_14955,N_14943);
or UO_910 (O_910,N_14919,N_14990);
xnor UO_911 (O_911,N_14906,N_14993);
xnor UO_912 (O_912,N_14892,N_14904);
or UO_913 (O_913,N_14937,N_14988);
or UO_914 (O_914,N_14956,N_14983);
nand UO_915 (O_915,N_14911,N_14966);
or UO_916 (O_916,N_14991,N_14955);
or UO_917 (O_917,N_14989,N_14991);
and UO_918 (O_918,N_14938,N_14948);
or UO_919 (O_919,N_14890,N_14875);
and UO_920 (O_920,N_14886,N_14942);
xnor UO_921 (O_921,N_14930,N_14972);
xor UO_922 (O_922,N_14905,N_14927);
xnor UO_923 (O_923,N_14984,N_14885);
xor UO_924 (O_924,N_14954,N_14937);
nand UO_925 (O_925,N_14887,N_14984);
or UO_926 (O_926,N_14878,N_14911);
and UO_927 (O_927,N_14923,N_14958);
xor UO_928 (O_928,N_14947,N_14919);
nor UO_929 (O_929,N_14994,N_14890);
nand UO_930 (O_930,N_14957,N_14882);
nand UO_931 (O_931,N_14919,N_14917);
or UO_932 (O_932,N_14949,N_14924);
nand UO_933 (O_933,N_14958,N_14906);
nor UO_934 (O_934,N_14913,N_14948);
and UO_935 (O_935,N_14921,N_14975);
and UO_936 (O_936,N_14879,N_14894);
and UO_937 (O_937,N_14953,N_14996);
and UO_938 (O_938,N_14944,N_14942);
nor UO_939 (O_939,N_14921,N_14881);
or UO_940 (O_940,N_14949,N_14929);
and UO_941 (O_941,N_14953,N_14912);
or UO_942 (O_942,N_14888,N_14912);
nor UO_943 (O_943,N_14953,N_14877);
nor UO_944 (O_944,N_14949,N_14887);
and UO_945 (O_945,N_14983,N_14897);
nor UO_946 (O_946,N_14898,N_14931);
nand UO_947 (O_947,N_14974,N_14944);
xnor UO_948 (O_948,N_14904,N_14991);
nor UO_949 (O_949,N_14983,N_14981);
xnor UO_950 (O_950,N_14876,N_14992);
nor UO_951 (O_951,N_14974,N_14908);
nor UO_952 (O_952,N_14973,N_14878);
and UO_953 (O_953,N_14877,N_14962);
xnor UO_954 (O_954,N_14931,N_14937);
nand UO_955 (O_955,N_14896,N_14915);
and UO_956 (O_956,N_14984,N_14962);
nand UO_957 (O_957,N_14970,N_14902);
xnor UO_958 (O_958,N_14909,N_14973);
xor UO_959 (O_959,N_14997,N_14899);
or UO_960 (O_960,N_14880,N_14973);
nor UO_961 (O_961,N_14885,N_14911);
nor UO_962 (O_962,N_14904,N_14986);
nor UO_963 (O_963,N_14966,N_14952);
nor UO_964 (O_964,N_14927,N_14884);
nor UO_965 (O_965,N_14951,N_14955);
and UO_966 (O_966,N_14906,N_14925);
xor UO_967 (O_967,N_14924,N_14987);
or UO_968 (O_968,N_14937,N_14998);
or UO_969 (O_969,N_14978,N_14979);
xnor UO_970 (O_970,N_14970,N_14988);
and UO_971 (O_971,N_14994,N_14901);
and UO_972 (O_972,N_14890,N_14887);
and UO_973 (O_973,N_14978,N_14958);
nor UO_974 (O_974,N_14949,N_14917);
and UO_975 (O_975,N_14891,N_14918);
nor UO_976 (O_976,N_14885,N_14940);
nor UO_977 (O_977,N_14915,N_14883);
xnor UO_978 (O_978,N_14899,N_14987);
or UO_979 (O_979,N_14888,N_14889);
nand UO_980 (O_980,N_14925,N_14930);
xnor UO_981 (O_981,N_14971,N_14879);
or UO_982 (O_982,N_14977,N_14894);
nor UO_983 (O_983,N_14945,N_14936);
and UO_984 (O_984,N_14911,N_14962);
nor UO_985 (O_985,N_14975,N_14891);
or UO_986 (O_986,N_14920,N_14994);
or UO_987 (O_987,N_14897,N_14973);
and UO_988 (O_988,N_14961,N_14986);
xor UO_989 (O_989,N_14883,N_14982);
or UO_990 (O_990,N_14911,N_14927);
nor UO_991 (O_991,N_14901,N_14993);
nor UO_992 (O_992,N_14998,N_14886);
nand UO_993 (O_993,N_14890,N_14908);
and UO_994 (O_994,N_14894,N_14904);
and UO_995 (O_995,N_14989,N_14958);
xor UO_996 (O_996,N_14885,N_14991);
and UO_997 (O_997,N_14953,N_14974);
nor UO_998 (O_998,N_14884,N_14968);
nor UO_999 (O_999,N_14930,N_14878);
nand UO_1000 (O_1000,N_14966,N_14975);
nor UO_1001 (O_1001,N_14945,N_14908);
nand UO_1002 (O_1002,N_14938,N_14940);
and UO_1003 (O_1003,N_14902,N_14901);
or UO_1004 (O_1004,N_14993,N_14929);
or UO_1005 (O_1005,N_14964,N_14944);
nor UO_1006 (O_1006,N_14903,N_14898);
xnor UO_1007 (O_1007,N_14899,N_14908);
nor UO_1008 (O_1008,N_14922,N_14994);
nor UO_1009 (O_1009,N_14977,N_14997);
nor UO_1010 (O_1010,N_14891,N_14921);
xor UO_1011 (O_1011,N_14924,N_14889);
or UO_1012 (O_1012,N_14940,N_14943);
nand UO_1013 (O_1013,N_14883,N_14975);
or UO_1014 (O_1014,N_14927,N_14919);
nand UO_1015 (O_1015,N_14904,N_14883);
nand UO_1016 (O_1016,N_14927,N_14910);
nand UO_1017 (O_1017,N_14899,N_14900);
nor UO_1018 (O_1018,N_14904,N_14911);
and UO_1019 (O_1019,N_14987,N_14920);
and UO_1020 (O_1020,N_14974,N_14920);
and UO_1021 (O_1021,N_14882,N_14927);
nand UO_1022 (O_1022,N_14889,N_14976);
nand UO_1023 (O_1023,N_14911,N_14955);
nor UO_1024 (O_1024,N_14906,N_14900);
nand UO_1025 (O_1025,N_14909,N_14898);
and UO_1026 (O_1026,N_14959,N_14904);
nand UO_1027 (O_1027,N_14994,N_14926);
nand UO_1028 (O_1028,N_14916,N_14880);
and UO_1029 (O_1029,N_14882,N_14891);
nor UO_1030 (O_1030,N_14875,N_14933);
xor UO_1031 (O_1031,N_14938,N_14890);
or UO_1032 (O_1032,N_14887,N_14963);
nand UO_1033 (O_1033,N_14888,N_14933);
and UO_1034 (O_1034,N_14933,N_14962);
or UO_1035 (O_1035,N_14917,N_14882);
nor UO_1036 (O_1036,N_14931,N_14897);
nand UO_1037 (O_1037,N_14991,N_14908);
xor UO_1038 (O_1038,N_14876,N_14990);
nand UO_1039 (O_1039,N_14972,N_14997);
xnor UO_1040 (O_1040,N_14973,N_14979);
nor UO_1041 (O_1041,N_14953,N_14990);
or UO_1042 (O_1042,N_14892,N_14987);
xnor UO_1043 (O_1043,N_14937,N_14965);
nand UO_1044 (O_1044,N_14974,N_14984);
or UO_1045 (O_1045,N_14958,N_14929);
nand UO_1046 (O_1046,N_14897,N_14930);
nor UO_1047 (O_1047,N_14939,N_14922);
and UO_1048 (O_1048,N_14904,N_14964);
and UO_1049 (O_1049,N_14884,N_14877);
nor UO_1050 (O_1050,N_14990,N_14966);
nor UO_1051 (O_1051,N_14914,N_14977);
nand UO_1052 (O_1052,N_14887,N_14954);
and UO_1053 (O_1053,N_14906,N_14945);
nand UO_1054 (O_1054,N_14879,N_14941);
xnor UO_1055 (O_1055,N_14984,N_14976);
and UO_1056 (O_1056,N_14892,N_14963);
and UO_1057 (O_1057,N_14999,N_14902);
nor UO_1058 (O_1058,N_14979,N_14989);
nor UO_1059 (O_1059,N_14879,N_14904);
and UO_1060 (O_1060,N_14894,N_14905);
xor UO_1061 (O_1061,N_14959,N_14923);
or UO_1062 (O_1062,N_14930,N_14884);
and UO_1063 (O_1063,N_14998,N_14950);
or UO_1064 (O_1064,N_14961,N_14928);
xnor UO_1065 (O_1065,N_14879,N_14890);
xor UO_1066 (O_1066,N_14899,N_14982);
nor UO_1067 (O_1067,N_14934,N_14884);
nand UO_1068 (O_1068,N_14972,N_14885);
and UO_1069 (O_1069,N_14943,N_14909);
xor UO_1070 (O_1070,N_14939,N_14924);
and UO_1071 (O_1071,N_14967,N_14899);
or UO_1072 (O_1072,N_14985,N_14911);
xor UO_1073 (O_1073,N_14912,N_14924);
nor UO_1074 (O_1074,N_14909,N_14878);
nand UO_1075 (O_1075,N_14895,N_14937);
and UO_1076 (O_1076,N_14918,N_14967);
nand UO_1077 (O_1077,N_14908,N_14937);
nand UO_1078 (O_1078,N_14906,N_14921);
xnor UO_1079 (O_1079,N_14946,N_14899);
xor UO_1080 (O_1080,N_14909,N_14903);
or UO_1081 (O_1081,N_14944,N_14889);
xor UO_1082 (O_1082,N_14938,N_14954);
nor UO_1083 (O_1083,N_14886,N_14975);
or UO_1084 (O_1084,N_14914,N_14892);
nor UO_1085 (O_1085,N_14889,N_14909);
nor UO_1086 (O_1086,N_14954,N_14909);
nand UO_1087 (O_1087,N_14903,N_14979);
nor UO_1088 (O_1088,N_14976,N_14954);
nor UO_1089 (O_1089,N_14992,N_14903);
xor UO_1090 (O_1090,N_14952,N_14916);
nor UO_1091 (O_1091,N_14936,N_14882);
nor UO_1092 (O_1092,N_14996,N_14967);
nor UO_1093 (O_1093,N_14982,N_14886);
nand UO_1094 (O_1094,N_14913,N_14947);
xnor UO_1095 (O_1095,N_14944,N_14932);
and UO_1096 (O_1096,N_14921,N_14962);
nor UO_1097 (O_1097,N_14970,N_14906);
and UO_1098 (O_1098,N_14952,N_14875);
nand UO_1099 (O_1099,N_14933,N_14972);
nor UO_1100 (O_1100,N_14908,N_14893);
nand UO_1101 (O_1101,N_14967,N_14913);
nand UO_1102 (O_1102,N_14979,N_14892);
and UO_1103 (O_1103,N_14991,N_14953);
or UO_1104 (O_1104,N_14993,N_14884);
xor UO_1105 (O_1105,N_14899,N_14989);
nor UO_1106 (O_1106,N_14914,N_14939);
xnor UO_1107 (O_1107,N_14987,N_14940);
and UO_1108 (O_1108,N_14919,N_14956);
xor UO_1109 (O_1109,N_14954,N_14999);
nor UO_1110 (O_1110,N_14908,N_14895);
or UO_1111 (O_1111,N_14971,N_14903);
or UO_1112 (O_1112,N_14943,N_14919);
and UO_1113 (O_1113,N_14996,N_14962);
nand UO_1114 (O_1114,N_14926,N_14938);
nor UO_1115 (O_1115,N_14930,N_14988);
and UO_1116 (O_1116,N_14916,N_14895);
nor UO_1117 (O_1117,N_14990,N_14982);
nand UO_1118 (O_1118,N_14888,N_14993);
xor UO_1119 (O_1119,N_14955,N_14967);
xor UO_1120 (O_1120,N_14962,N_14940);
nor UO_1121 (O_1121,N_14948,N_14994);
or UO_1122 (O_1122,N_14875,N_14914);
nor UO_1123 (O_1123,N_14924,N_14914);
nand UO_1124 (O_1124,N_14992,N_14948);
nand UO_1125 (O_1125,N_14934,N_14951);
xor UO_1126 (O_1126,N_14883,N_14998);
xnor UO_1127 (O_1127,N_14922,N_14906);
and UO_1128 (O_1128,N_14954,N_14899);
nor UO_1129 (O_1129,N_14974,N_14965);
nand UO_1130 (O_1130,N_14904,N_14965);
and UO_1131 (O_1131,N_14997,N_14903);
xnor UO_1132 (O_1132,N_14974,N_14976);
and UO_1133 (O_1133,N_14931,N_14932);
xor UO_1134 (O_1134,N_14973,N_14960);
nand UO_1135 (O_1135,N_14888,N_14975);
xor UO_1136 (O_1136,N_14975,N_14943);
and UO_1137 (O_1137,N_14893,N_14914);
or UO_1138 (O_1138,N_14980,N_14885);
nand UO_1139 (O_1139,N_14910,N_14997);
and UO_1140 (O_1140,N_14900,N_14914);
nand UO_1141 (O_1141,N_14945,N_14899);
xnor UO_1142 (O_1142,N_14892,N_14937);
and UO_1143 (O_1143,N_14967,N_14998);
xor UO_1144 (O_1144,N_14962,N_14966);
nor UO_1145 (O_1145,N_14987,N_14958);
nor UO_1146 (O_1146,N_14950,N_14921);
nand UO_1147 (O_1147,N_14982,N_14885);
or UO_1148 (O_1148,N_14953,N_14947);
and UO_1149 (O_1149,N_14886,N_14967);
or UO_1150 (O_1150,N_14976,N_14938);
or UO_1151 (O_1151,N_14910,N_14898);
or UO_1152 (O_1152,N_14989,N_14968);
xnor UO_1153 (O_1153,N_14943,N_14949);
nor UO_1154 (O_1154,N_14922,N_14954);
nor UO_1155 (O_1155,N_14932,N_14985);
xor UO_1156 (O_1156,N_14998,N_14887);
nand UO_1157 (O_1157,N_14984,N_14950);
nor UO_1158 (O_1158,N_14991,N_14959);
or UO_1159 (O_1159,N_14927,N_14929);
nor UO_1160 (O_1160,N_14978,N_14926);
and UO_1161 (O_1161,N_14881,N_14890);
nor UO_1162 (O_1162,N_14990,N_14996);
and UO_1163 (O_1163,N_14886,N_14880);
or UO_1164 (O_1164,N_14983,N_14939);
xnor UO_1165 (O_1165,N_14900,N_14901);
or UO_1166 (O_1166,N_14919,N_14950);
and UO_1167 (O_1167,N_14997,N_14887);
and UO_1168 (O_1168,N_14947,N_14979);
xnor UO_1169 (O_1169,N_14988,N_14887);
nand UO_1170 (O_1170,N_14900,N_14881);
nor UO_1171 (O_1171,N_14917,N_14922);
nor UO_1172 (O_1172,N_14971,N_14968);
nor UO_1173 (O_1173,N_14935,N_14982);
or UO_1174 (O_1174,N_14984,N_14918);
xor UO_1175 (O_1175,N_14938,N_14910);
nor UO_1176 (O_1176,N_14947,N_14939);
nand UO_1177 (O_1177,N_14916,N_14915);
nand UO_1178 (O_1178,N_14979,N_14968);
nor UO_1179 (O_1179,N_14978,N_14934);
and UO_1180 (O_1180,N_14992,N_14954);
and UO_1181 (O_1181,N_14939,N_14930);
or UO_1182 (O_1182,N_14969,N_14999);
nor UO_1183 (O_1183,N_14881,N_14977);
nand UO_1184 (O_1184,N_14920,N_14988);
nand UO_1185 (O_1185,N_14930,N_14961);
nor UO_1186 (O_1186,N_14902,N_14967);
nor UO_1187 (O_1187,N_14894,N_14918);
or UO_1188 (O_1188,N_14897,N_14998);
or UO_1189 (O_1189,N_14901,N_14893);
and UO_1190 (O_1190,N_14935,N_14947);
and UO_1191 (O_1191,N_14892,N_14969);
xnor UO_1192 (O_1192,N_14883,N_14881);
xnor UO_1193 (O_1193,N_14969,N_14882);
nor UO_1194 (O_1194,N_14972,N_14977);
or UO_1195 (O_1195,N_14911,N_14916);
nor UO_1196 (O_1196,N_14877,N_14903);
nor UO_1197 (O_1197,N_14926,N_14986);
xor UO_1198 (O_1198,N_14879,N_14931);
nand UO_1199 (O_1199,N_14983,N_14945);
nand UO_1200 (O_1200,N_14929,N_14937);
nor UO_1201 (O_1201,N_14994,N_14903);
xor UO_1202 (O_1202,N_14943,N_14910);
xor UO_1203 (O_1203,N_14921,N_14925);
xnor UO_1204 (O_1204,N_14988,N_14993);
or UO_1205 (O_1205,N_14975,N_14876);
and UO_1206 (O_1206,N_14923,N_14878);
nand UO_1207 (O_1207,N_14974,N_14882);
nor UO_1208 (O_1208,N_14916,N_14882);
nor UO_1209 (O_1209,N_14987,N_14978);
xnor UO_1210 (O_1210,N_14881,N_14929);
xnor UO_1211 (O_1211,N_14990,N_14911);
nor UO_1212 (O_1212,N_14987,N_14964);
nand UO_1213 (O_1213,N_14965,N_14947);
nor UO_1214 (O_1214,N_14960,N_14961);
nor UO_1215 (O_1215,N_14990,N_14890);
nor UO_1216 (O_1216,N_14921,N_14943);
xor UO_1217 (O_1217,N_14996,N_14936);
nand UO_1218 (O_1218,N_14907,N_14952);
xnor UO_1219 (O_1219,N_14881,N_14878);
xor UO_1220 (O_1220,N_14911,N_14925);
and UO_1221 (O_1221,N_14879,N_14892);
or UO_1222 (O_1222,N_14895,N_14934);
and UO_1223 (O_1223,N_14920,N_14935);
nor UO_1224 (O_1224,N_14923,N_14989);
and UO_1225 (O_1225,N_14899,N_14950);
nor UO_1226 (O_1226,N_14968,N_14934);
nand UO_1227 (O_1227,N_14884,N_14925);
nor UO_1228 (O_1228,N_14926,N_14894);
or UO_1229 (O_1229,N_14990,N_14889);
nor UO_1230 (O_1230,N_14908,N_14977);
or UO_1231 (O_1231,N_14979,N_14910);
nor UO_1232 (O_1232,N_14891,N_14995);
and UO_1233 (O_1233,N_14912,N_14999);
and UO_1234 (O_1234,N_14970,N_14883);
nand UO_1235 (O_1235,N_14972,N_14918);
or UO_1236 (O_1236,N_14971,N_14991);
and UO_1237 (O_1237,N_14937,N_14927);
and UO_1238 (O_1238,N_14972,N_14917);
nor UO_1239 (O_1239,N_14934,N_14939);
nor UO_1240 (O_1240,N_14914,N_14880);
nand UO_1241 (O_1241,N_14921,N_14903);
or UO_1242 (O_1242,N_14955,N_14993);
or UO_1243 (O_1243,N_14885,N_14974);
nor UO_1244 (O_1244,N_14887,N_14902);
xor UO_1245 (O_1245,N_14959,N_14963);
nor UO_1246 (O_1246,N_14943,N_14979);
xor UO_1247 (O_1247,N_14954,N_14894);
xnor UO_1248 (O_1248,N_14989,N_14975);
xnor UO_1249 (O_1249,N_14924,N_14975);
xor UO_1250 (O_1250,N_14936,N_14884);
and UO_1251 (O_1251,N_14913,N_14997);
or UO_1252 (O_1252,N_14958,N_14934);
xor UO_1253 (O_1253,N_14908,N_14882);
xnor UO_1254 (O_1254,N_14938,N_14991);
and UO_1255 (O_1255,N_14940,N_14918);
nand UO_1256 (O_1256,N_14994,N_14992);
or UO_1257 (O_1257,N_14934,N_14907);
or UO_1258 (O_1258,N_14967,N_14946);
nand UO_1259 (O_1259,N_14914,N_14929);
xor UO_1260 (O_1260,N_14964,N_14968);
and UO_1261 (O_1261,N_14979,N_14998);
nor UO_1262 (O_1262,N_14983,N_14996);
and UO_1263 (O_1263,N_14882,N_14975);
and UO_1264 (O_1264,N_14983,N_14908);
and UO_1265 (O_1265,N_14968,N_14897);
and UO_1266 (O_1266,N_14958,N_14947);
xnor UO_1267 (O_1267,N_14937,N_14948);
xnor UO_1268 (O_1268,N_14952,N_14890);
nand UO_1269 (O_1269,N_14902,N_14905);
and UO_1270 (O_1270,N_14946,N_14995);
xor UO_1271 (O_1271,N_14979,N_14898);
nand UO_1272 (O_1272,N_14951,N_14916);
and UO_1273 (O_1273,N_14966,N_14998);
and UO_1274 (O_1274,N_14995,N_14900);
nor UO_1275 (O_1275,N_14925,N_14901);
xor UO_1276 (O_1276,N_14915,N_14948);
and UO_1277 (O_1277,N_14985,N_14973);
nor UO_1278 (O_1278,N_14951,N_14965);
or UO_1279 (O_1279,N_14950,N_14991);
xnor UO_1280 (O_1280,N_14901,N_14949);
and UO_1281 (O_1281,N_14931,N_14976);
and UO_1282 (O_1282,N_14939,N_14962);
and UO_1283 (O_1283,N_14988,N_14927);
nor UO_1284 (O_1284,N_14918,N_14924);
and UO_1285 (O_1285,N_14999,N_14917);
xor UO_1286 (O_1286,N_14959,N_14966);
nand UO_1287 (O_1287,N_14995,N_14999);
and UO_1288 (O_1288,N_14912,N_14919);
nor UO_1289 (O_1289,N_14983,N_14952);
nand UO_1290 (O_1290,N_14948,N_14973);
nor UO_1291 (O_1291,N_14960,N_14912);
or UO_1292 (O_1292,N_14899,N_14995);
nand UO_1293 (O_1293,N_14986,N_14935);
or UO_1294 (O_1294,N_14913,N_14906);
nand UO_1295 (O_1295,N_14883,N_14966);
or UO_1296 (O_1296,N_14985,N_14946);
and UO_1297 (O_1297,N_14938,N_14883);
nand UO_1298 (O_1298,N_14914,N_14889);
xor UO_1299 (O_1299,N_14892,N_14961);
or UO_1300 (O_1300,N_14976,N_14951);
nor UO_1301 (O_1301,N_14985,N_14889);
nor UO_1302 (O_1302,N_14934,N_14954);
xnor UO_1303 (O_1303,N_14980,N_14942);
or UO_1304 (O_1304,N_14993,N_14972);
xnor UO_1305 (O_1305,N_14979,N_14944);
xor UO_1306 (O_1306,N_14959,N_14960);
and UO_1307 (O_1307,N_14967,N_14879);
xnor UO_1308 (O_1308,N_14904,N_14985);
nand UO_1309 (O_1309,N_14905,N_14931);
and UO_1310 (O_1310,N_14963,N_14888);
xor UO_1311 (O_1311,N_14952,N_14938);
xnor UO_1312 (O_1312,N_14913,N_14941);
nand UO_1313 (O_1313,N_14913,N_14885);
or UO_1314 (O_1314,N_14893,N_14919);
xnor UO_1315 (O_1315,N_14973,N_14924);
nor UO_1316 (O_1316,N_14887,N_14897);
xor UO_1317 (O_1317,N_14890,N_14944);
or UO_1318 (O_1318,N_14968,N_14933);
nand UO_1319 (O_1319,N_14989,N_14889);
or UO_1320 (O_1320,N_14908,N_14978);
nand UO_1321 (O_1321,N_14943,N_14977);
nor UO_1322 (O_1322,N_14893,N_14938);
nor UO_1323 (O_1323,N_14877,N_14998);
or UO_1324 (O_1324,N_14947,N_14952);
and UO_1325 (O_1325,N_14891,N_14936);
nor UO_1326 (O_1326,N_14926,N_14911);
nor UO_1327 (O_1327,N_14990,N_14922);
nor UO_1328 (O_1328,N_14949,N_14880);
nor UO_1329 (O_1329,N_14878,N_14905);
nor UO_1330 (O_1330,N_14924,N_14968);
nor UO_1331 (O_1331,N_14940,N_14945);
xor UO_1332 (O_1332,N_14958,N_14900);
nand UO_1333 (O_1333,N_14994,N_14945);
xnor UO_1334 (O_1334,N_14888,N_14995);
nor UO_1335 (O_1335,N_14981,N_14939);
nand UO_1336 (O_1336,N_14879,N_14944);
and UO_1337 (O_1337,N_14954,N_14939);
xor UO_1338 (O_1338,N_14983,N_14877);
nor UO_1339 (O_1339,N_14928,N_14996);
or UO_1340 (O_1340,N_14906,N_14997);
and UO_1341 (O_1341,N_14975,N_14913);
and UO_1342 (O_1342,N_14928,N_14975);
or UO_1343 (O_1343,N_14933,N_14882);
nand UO_1344 (O_1344,N_14902,N_14950);
nand UO_1345 (O_1345,N_14919,N_14925);
nor UO_1346 (O_1346,N_14983,N_14893);
and UO_1347 (O_1347,N_14992,N_14979);
or UO_1348 (O_1348,N_14930,N_14888);
nor UO_1349 (O_1349,N_14910,N_14888);
and UO_1350 (O_1350,N_14933,N_14886);
and UO_1351 (O_1351,N_14982,N_14967);
nand UO_1352 (O_1352,N_14960,N_14922);
nor UO_1353 (O_1353,N_14959,N_14961);
and UO_1354 (O_1354,N_14926,N_14983);
nor UO_1355 (O_1355,N_14970,N_14892);
and UO_1356 (O_1356,N_14894,N_14903);
xor UO_1357 (O_1357,N_14912,N_14975);
and UO_1358 (O_1358,N_14916,N_14965);
or UO_1359 (O_1359,N_14899,N_14890);
and UO_1360 (O_1360,N_14934,N_14926);
nand UO_1361 (O_1361,N_14916,N_14984);
and UO_1362 (O_1362,N_14996,N_14976);
xor UO_1363 (O_1363,N_14918,N_14896);
nand UO_1364 (O_1364,N_14951,N_14894);
xor UO_1365 (O_1365,N_14921,N_14902);
nand UO_1366 (O_1366,N_14897,N_14914);
nor UO_1367 (O_1367,N_14938,N_14922);
or UO_1368 (O_1368,N_14903,N_14935);
and UO_1369 (O_1369,N_14897,N_14906);
xnor UO_1370 (O_1370,N_14921,N_14893);
nand UO_1371 (O_1371,N_14878,N_14876);
xor UO_1372 (O_1372,N_14892,N_14932);
and UO_1373 (O_1373,N_14969,N_14988);
or UO_1374 (O_1374,N_14953,N_14902);
or UO_1375 (O_1375,N_14987,N_14945);
xnor UO_1376 (O_1376,N_14889,N_14982);
xnor UO_1377 (O_1377,N_14935,N_14927);
or UO_1378 (O_1378,N_14893,N_14960);
nor UO_1379 (O_1379,N_14924,N_14986);
or UO_1380 (O_1380,N_14921,N_14920);
or UO_1381 (O_1381,N_14878,N_14996);
and UO_1382 (O_1382,N_14887,N_14981);
nor UO_1383 (O_1383,N_14966,N_14929);
and UO_1384 (O_1384,N_14910,N_14920);
nor UO_1385 (O_1385,N_14888,N_14991);
nand UO_1386 (O_1386,N_14981,N_14969);
nand UO_1387 (O_1387,N_14969,N_14977);
nor UO_1388 (O_1388,N_14968,N_14949);
nand UO_1389 (O_1389,N_14970,N_14966);
xor UO_1390 (O_1390,N_14898,N_14882);
xor UO_1391 (O_1391,N_14944,N_14941);
xnor UO_1392 (O_1392,N_14961,N_14981);
or UO_1393 (O_1393,N_14953,N_14976);
xor UO_1394 (O_1394,N_14990,N_14989);
or UO_1395 (O_1395,N_14958,N_14976);
nor UO_1396 (O_1396,N_14978,N_14995);
nor UO_1397 (O_1397,N_14942,N_14912);
xor UO_1398 (O_1398,N_14943,N_14887);
nand UO_1399 (O_1399,N_14943,N_14999);
xnor UO_1400 (O_1400,N_14993,N_14956);
xnor UO_1401 (O_1401,N_14948,N_14998);
xnor UO_1402 (O_1402,N_14956,N_14881);
nand UO_1403 (O_1403,N_14911,N_14963);
nor UO_1404 (O_1404,N_14937,N_14949);
and UO_1405 (O_1405,N_14926,N_14974);
nor UO_1406 (O_1406,N_14964,N_14886);
nor UO_1407 (O_1407,N_14978,N_14875);
or UO_1408 (O_1408,N_14937,N_14963);
or UO_1409 (O_1409,N_14978,N_14970);
nor UO_1410 (O_1410,N_14912,N_14925);
xor UO_1411 (O_1411,N_14911,N_14942);
and UO_1412 (O_1412,N_14972,N_14876);
xnor UO_1413 (O_1413,N_14952,N_14879);
or UO_1414 (O_1414,N_14967,N_14894);
nor UO_1415 (O_1415,N_14914,N_14937);
or UO_1416 (O_1416,N_14986,N_14955);
nand UO_1417 (O_1417,N_14959,N_14894);
or UO_1418 (O_1418,N_14956,N_14942);
and UO_1419 (O_1419,N_14889,N_14896);
or UO_1420 (O_1420,N_14896,N_14875);
nand UO_1421 (O_1421,N_14920,N_14958);
or UO_1422 (O_1422,N_14882,N_14962);
and UO_1423 (O_1423,N_14935,N_14996);
and UO_1424 (O_1424,N_14893,N_14935);
nand UO_1425 (O_1425,N_14916,N_14906);
nor UO_1426 (O_1426,N_14886,N_14891);
and UO_1427 (O_1427,N_14933,N_14895);
nand UO_1428 (O_1428,N_14877,N_14922);
nand UO_1429 (O_1429,N_14986,N_14894);
xor UO_1430 (O_1430,N_14923,N_14896);
nand UO_1431 (O_1431,N_14927,N_14950);
or UO_1432 (O_1432,N_14924,N_14989);
or UO_1433 (O_1433,N_14960,N_14908);
nand UO_1434 (O_1434,N_14999,N_14978);
xnor UO_1435 (O_1435,N_14956,N_14970);
and UO_1436 (O_1436,N_14913,N_14889);
nor UO_1437 (O_1437,N_14875,N_14992);
and UO_1438 (O_1438,N_14997,N_14908);
xor UO_1439 (O_1439,N_14878,N_14910);
xor UO_1440 (O_1440,N_14893,N_14956);
and UO_1441 (O_1441,N_14875,N_14960);
and UO_1442 (O_1442,N_14917,N_14930);
nand UO_1443 (O_1443,N_14980,N_14962);
and UO_1444 (O_1444,N_14894,N_14935);
nor UO_1445 (O_1445,N_14888,N_14877);
or UO_1446 (O_1446,N_14970,N_14927);
nor UO_1447 (O_1447,N_14894,N_14938);
and UO_1448 (O_1448,N_14903,N_14924);
nand UO_1449 (O_1449,N_14939,N_14980);
xnor UO_1450 (O_1450,N_14968,N_14954);
xor UO_1451 (O_1451,N_14988,N_14957);
xor UO_1452 (O_1452,N_14950,N_14955);
and UO_1453 (O_1453,N_14904,N_14992);
or UO_1454 (O_1454,N_14905,N_14999);
nor UO_1455 (O_1455,N_14886,N_14884);
and UO_1456 (O_1456,N_14926,N_14940);
nand UO_1457 (O_1457,N_14926,N_14959);
or UO_1458 (O_1458,N_14912,N_14938);
and UO_1459 (O_1459,N_14955,N_14925);
or UO_1460 (O_1460,N_14913,N_14884);
nand UO_1461 (O_1461,N_14971,N_14955);
or UO_1462 (O_1462,N_14926,N_14912);
nor UO_1463 (O_1463,N_14997,N_14951);
or UO_1464 (O_1464,N_14955,N_14926);
and UO_1465 (O_1465,N_14923,N_14970);
or UO_1466 (O_1466,N_14926,N_14980);
nand UO_1467 (O_1467,N_14969,N_14924);
and UO_1468 (O_1468,N_14908,N_14957);
nand UO_1469 (O_1469,N_14996,N_14974);
nand UO_1470 (O_1470,N_14902,N_14920);
or UO_1471 (O_1471,N_14958,N_14999);
xnor UO_1472 (O_1472,N_14963,N_14990);
and UO_1473 (O_1473,N_14996,N_14898);
and UO_1474 (O_1474,N_14916,N_14971);
xnor UO_1475 (O_1475,N_14875,N_14977);
and UO_1476 (O_1476,N_14966,N_14932);
xor UO_1477 (O_1477,N_14932,N_14956);
xor UO_1478 (O_1478,N_14915,N_14885);
nor UO_1479 (O_1479,N_14888,N_14951);
and UO_1480 (O_1480,N_14990,N_14888);
nand UO_1481 (O_1481,N_14958,N_14902);
nor UO_1482 (O_1482,N_14922,N_14989);
and UO_1483 (O_1483,N_14890,N_14904);
xor UO_1484 (O_1484,N_14916,N_14941);
xnor UO_1485 (O_1485,N_14997,N_14890);
and UO_1486 (O_1486,N_14931,N_14953);
or UO_1487 (O_1487,N_14947,N_14901);
nand UO_1488 (O_1488,N_14992,N_14962);
nand UO_1489 (O_1489,N_14974,N_14951);
nor UO_1490 (O_1490,N_14931,N_14892);
and UO_1491 (O_1491,N_14901,N_14986);
or UO_1492 (O_1492,N_14980,N_14970);
nand UO_1493 (O_1493,N_14988,N_14971);
xor UO_1494 (O_1494,N_14909,N_14892);
or UO_1495 (O_1495,N_14901,N_14880);
or UO_1496 (O_1496,N_14980,N_14918);
nor UO_1497 (O_1497,N_14936,N_14909);
and UO_1498 (O_1498,N_14977,N_14876);
xnor UO_1499 (O_1499,N_14949,N_14906);
xnor UO_1500 (O_1500,N_14994,N_14889);
nand UO_1501 (O_1501,N_14906,N_14924);
xor UO_1502 (O_1502,N_14905,N_14954);
and UO_1503 (O_1503,N_14947,N_14980);
xor UO_1504 (O_1504,N_14973,N_14918);
nor UO_1505 (O_1505,N_14966,N_14923);
and UO_1506 (O_1506,N_14946,N_14906);
xor UO_1507 (O_1507,N_14999,N_14882);
nor UO_1508 (O_1508,N_14930,N_14979);
xnor UO_1509 (O_1509,N_14888,N_14941);
or UO_1510 (O_1510,N_14957,N_14895);
nand UO_1511 (O_1511,N_14936,N_14893);
or UO_1512 (O_1512,N_14926,N_14976);
xnor UO_1513 (O_1513,N_14977,N_14904);
or UO_1514 (O_1514,N_14934,N_14882);
nand UO_1515 (O_1515,N_14875,N_14983);
nor UO_1516 (O_1516,N_14986,N_14959);
nor UO_1517 (O_1517,N_14951,N_14975);
and UO_1518 (O_1518,N_14970,N_14938);
nor UO_1519 (O_1519,N_14951,N_14931);
nor UO_1520 (O_1520,N_14878,N_14981);
nor UO_1521 (O_1521,N_14906,N_14983);
and UO_1522 (O_1522,N_14989,N_14897);
xor UO_1523 (O_1523,N_14942,N_14893);
nor UO_1524 (O_1524,N_14950,N_14934);
nand UO_1525 (O_1525,N_14992,N_14915);
nor UO_1526 (O_1526,N_14995,N_14971);
or UO_1527 (O_1527,N_14966,N_14976);
xnor UO_1528 (O_1528,N_14993,N_14917);
nand UO_1529 (O_1529,N_14890,N_14947);
xnor UO_1530 (O_1530,N_14900,N_14980);
nor UO_1531 (O_1531,N_14891,N_14906);
and UO_1532 (O_1532,N_14904,N_14972);
nand UO_1533 (O_1533,N_14895,N_14936);
or UO_1534 (O_1534,N_14981,N_14957);
xnor UO_1535 (O_1535,N_14994,N_14906);
xor UO_1536 (O_1536,N_14961,N_14882);
nand UO_1537 (O_1537,N_14881,N_14889);
nand UO_1538 (O_1538,N_14908,N_14946);
and UO_1539 (O_1539,N_14910,N_14948);
xor UO_1540 (O_1540,N_14950,N_14958);
nand UO_1541 (O_1541,N_14974,N_14890);
or UO_1542 (O_1542,N_14970,N_14968);
xor UO_1543 (O_1543,N_14981,N_14903);
or UO_1544 (O_1544,N_14954,N_14967);
or UO_1545 (O_1545,N_14897,N_14908);
and UO_1546 (O_1546,N_14985,N_14906);
xnor UO_1547 (O_1547,N_14918,N_14899);
nor UO_1548 (O_1548,N_14964,N_14967);
or UO_1549 (O_1549,N_14929,N_14967);
and UO_1550 (O_1550,N_14903,N_14895);
nand UO_1551 (O_1551,N_14987,N_14878);
nor UO_1552 (O_1552,N_14985,N_14982);
nand UO_1553 (O_1553,N_14943,N_14960);
or UO_1554 (O_1554,N_14997,N_14965);
nand UO_1555 (O_1555,N_14932,N_14895);
and UO_1556 (O_1556,N_14951,N_14896);
xor UO_1557 (O_1557,N_14997,N_14941);
nand UO_1558 (O_1558,N_14971,N_14998);
nand UO_1559 (O_1559,N_14995,N_14982);
xnor UO_1560 (O_1560,N_14924,N_14972);
or UO_1561 (O_1561,N_14903,N_14976);
nand UO_1562 (O_1562,N_14922,N_14921);
or UO_1563 (O_1563,N_14964,N_14970);
and UO_1564 (O_1564,N_14943,N_14950);
nor UO_1565 (O_1565,N_14935,N_14901);
nand UO_1566 (O_1566,N_14926,N_14885);
nand UO_1567 (O_1567,N_14923,N_14967);
xor UO_1568 (O_1568,N_14982,N_14977);
nand UO_1569 (O_1569,N_14904,N_14885);
nor UO_1570 (O_1570,N_14980,N_14903);
or UO_1571 (O_1571,N_14955,N_14901);
xnor UO_1572 (O_1572,N_14940,N_14915);
and UO_1573 (O_1573,N_14910,N_14913);
and UO_1574 (O_1574,N_14918,N_14959);
nand UO_1575 (O_1575,N_14913,N_14949);
or UO_1576 (O_1576,N_14911,N_14923);
xnor UO_1577 (O_1577,N_14928,N_14965);
nor UO_1578 (O_1578,N_14973,N_14996);
xnor UO_1579 (O_1579,N_14991,N_14956);
nand UO_1580 (O_1580,N_14952,N_14978);
and UO_1581 (O_1581,N_14915,N_14880);
nor UO_1582 (O_1582,N_14906,N_14917);
xnor UO_1583 (O_1583,N_14999,N_14944);
xor UO_1584 (O_1584,N_14982,N_14917);
nor UO_1585 (O_1585,N_14932,N_14955);
nand UO_1586 (O_1586,N_14988,N_14950);
or UO_1587 (O_1587,N_14977,N_14903);
nor UO_1588 (O_1588,N_14908,N_14995);
xnor UO_1589 (O_1589,N_14995,N_14996);
and UO_1590 (O_1590,N_14986,N_14944);
or UO_1591 (O_1591,N_14945,N_14958);
nor UO_1592 (O_1592,N_14994,N_14987);
or UO_1593 (O_1593,N_14934,N_14997);
and UO_1594 (O_1594,N_14920,N_14961);
or UO_1595 (O_1595,N_14903,N_14993);
or UO_1596 (O_1596,N_14976,N_14970);
nand UO_1597 (O_1597,N_14901,N_14899);
nor UO_1598 (O_1598,N_14992,N_14926);
nor UO_1599 (O_1599,N_14977,N_14968);
and UO_1600 (O_1600,N_14988,N_14976);
or UO_1601 (O_1601,N_14915,N_14886);
nor UO_1602 (O_1602,N_14931,N_14992);
nor UO_1603 (O_1603,N_14946,N_14942);
nor UO_1604 (O_1604,N_14956,N_14900);
nand UO_1605 (O_1605,N_14967,N_14973);
or UO_1606 (O_1606,N_14887,N_14938);
nand UO_1607 (O_1607,N_14883,N_14942);
or UO_1608 (O_1608,N_14992,N_14910);
nand UO_1609 (O_1609,N_14908,N_14909);
or UO_1610 (O_1610,N_14975,N_14929);
and UO_1611 (O_1611,N_14912,N_14971);
nand UO_1612 (O_1612,N_14877,N_14956);
and UO_1613 (O_1613,N_14990,N_14946);
and UO_1614 (O_1614,N_14963,N_14914);
and UO_1615 (O_1615,N_14921,N_14968);
or UO_1616 (O_1616,N_14954,N_14878);
or UO_1617 (O_1617,N_14889,N_14893);
or UO_1618 (O_1618,N_14883,N_14878);
xnor UO_1619 (O_1619,N_14875,N_14893);
nor UO_1620 (O_1620,N_14938,N_14951);
nand UO_1621 (O_1621,N_14991,N_14930);
nand UO_1622 (O_1622,N_14975,N_14910);
nand UO_1623 (O_1623,N_14912,N_14950);
and UO_1624 (O_1624,N_14891,N_14901);
nand UO_1625 (O_1625,N_14961,N_14992);
xor UO_1626 (O_1626,N_14975,N_14960);
nand UO_1627 (O_1627,N_14897,N_14971);
nor UO_1628 (O_1628,N_14963,N_14971);
and UO_1629 (O_1629,N_14919,N_14996);
nor UO_1630 (O_1630,N_14980,N_14886);
nand UO_1631 (O_1631,N_14885,N_14970);
or UO_1632 (O_1632,N_14967,N_14883);
nand UO_1633 (O_1633,N_14993,N_14913);
and UO_1634 (O_1634,N_14955,N_14959);
or UO_1635 (O_1635,N_14966,N_14933);
and UO_1636 (O_1636,N_14905,N_14892);
nand UO_1637 (O_1637,N_14897,N_14947);
nor UO_1638 (O_1638,N_14986,N_14945);
or UO_1639 (O_1639,N_14942,N_14915);
or UO_1640 (O_1640,N_14979,N_14906);
nand UO_1641 (O_1641,N_14996,N_14940);
and UO_1642 (O_1642,N_14937,N_14951);
nand UO_1643 (O_1643,N_14917,N_14905);
nand UO_1644 (O_1644,N_14929,N_14972);
nand UO_1645 (O_1645,N_14983,N_14980);
and UO_1646 (O_1646,N_14954,N_14980);
xnor UO_1647 (O_1647,N_14959,N_14983);
and UO_1648 (O_1648,N_14964,N_14992);
or UO_1649 (O_1649,N_14962,N_14893);
nor UO_1650 (O_1650,N_14895,N_14893);
nor UO_1651 (O_1651,N_14972,N_14936);
or UO_1652 (O_1652,N_14990,N_14958);
xor UO_1653 (O_1653,N_14985,N_14876);
nand UO_1654 (O_1654,N_14903,N_14922);
and UO_1655 (O_1655,N_14981,N_14927);
nor UO_1656 (O_1656,N_14941,N_14951);
nand UO_1657 (O_1657,N_14924,N_14945);
and UO_1658 (O_1658,N_14907,N_14949);
nand UO_1659 (O_1659,N_14964,N_14907);
and UO_1660 (O_1660,N_14897,N_14951);
nor UO_1661 (O_1661,N_14893,N_14912);
and UO_1662 (O_1662,N_14899,N_14937);
or UO_1663 (O_1663,N_14968,N_14886);
nor UO_1664 (O_1664,N_14938,N_14967);
nand UO_1665 (O_1665,N_14890,N_14988);
and UO_1666 (O_1666,N_14981,N_14909);
nand UO_1667 (O_1667,N_14944,N_14877);
nor UO_1668 (O_1668,N_14875,N_14988);
or UO_1669 (O_1669,N_14976,N_14977);
nand UO_1670 (O_1670,N_14918,N_14999);
and UO_1671 (O_1671,N_14875,N_14889);
and UO_1672 (O_1672,N_14972,N_14919);
nor UO_1673 (O_1673,N_14967,N_14988);
nand UO_1674 (O_1674,N_14973,N_14887);
nor UO_1675 (O_1675,N_14980,N_14968);
or UO_1676 (O_1676,N_14924,N_14913);
xnor UO_1677 (O_1677,N_14878,N_14903);
nand UO_1678 (O_1678,N_14941,N_14925);
nand UO_1679 (O_1679,N_14939,N_14997);
nand UO_1680 (O_1680,N_14920,N_14940);
and UO_1681 (O_1681,N_14929,N_14951);
xor UO_1682 (O_1682,N_14915,N_14983);
xor UO_1683 (O_1683,N_14905,N_14933);
nand UO_1684 (O_1684,N_14928,N_14955);
xor UO_1685 (O_1685,N_14929,N_14957);
nand UO_1686 (O_1686,N_14903,N_14917);
nand UO_1687 (O_1687,N_14912,N_14906);
nor UO_1688 (O_1688,N_14968,N_14902);
nor UO_1689 (O_1689,N_14893,N_14977);
or UO_1690 (O_1690,N_14962,N_14894);
or UO_1691 (O_1691,N_14970,N_14893);
nand UO_1692 (O_1692,N_14938,N_14878);
xnor UO_1693 (O_1693,N_14965,N_14970);
nor UO_1694 (O_1694,N_14940,N_14922);
and UO_1695 (O_1695,N_14887,N_14941);
or UO_1696 (O_1696,N_14884,N_14965);
nand UO_1697 (O_1697,N_14962,N_14990);
nor UO_1698 (O_1698,N_14904,N_14921);
and UO_1699 (O_1699,N_14910,N_14900);
nor UO_1700 (O_1700,N_14875,N_14906);
or UO_1701 (O_1701,N_14944,N_14923);
xnor UO_1702 (O_1702,N_14977,N_14993);
xnor UO_1703 (O_1703,N_14907,N_14941);
nor UO_1704 (O_1704,N_14931,N_14966);
and UO_1705 (O_1705,N_14970,N_14954);
nor UO_1706 (O_1706,N_14919,N_14918);
or UO_1707 (O_1707,N_14895,N_14979);
or UO_1708 (O_1708,N_14932,N_14991);
or UO_1709 (O_1709,N_14911,N_14937);
nor UO_1710 (O_1710,N_14914,N_14933);
nand UO_1711 (O_1711,N_14913,N_14986);
and UO_1712 (O_1712,N_14990,N_14914);
and UO_1713 (O_1713,N_14967,N_14912);
and UO_1714 (O_1714,N_14886,N_14889);
xor UO_1715 (O_1715,N_14944,N_14896);
nor UO_1716 (O_1716,N_14993,N_14908);
or UO_1717 (O_1717,N_14927,N_14984);
or UO_1718 (O_1718,N_14931,N_14941);
or UO_1719 (O_1719,N_14914,N_14950);
or UO_1720 (O_1720,N_14972,N_14981);
nor UO_1721 (O_1721,N_14905,N_14903);
nor UO_1722 (O_1722,N_14978,N_14990);
nor UO_1723 (O_1723,N_14883,N_14968);
nand UO_1724 (O_1724,N_14907,N_14998);
nand UO_1725 (O_1725,N_14934,N_14961);
and UO_1726 (O_1726,N_14903,N_14932);
nor UO_1727 (O_1727,N_14898,N_14975);
xnor UO_1728 (O_1728,N_14908,N_14939);
nor UO_1729 (O_1729,N_14945,N_14916);
or UO_1730 (O_1730,N_14944,N_14917);
nor UO_1731 (O_1731,N_14945,N_14984);
and UO_1732 (O_1732,N_14923,N_14964);
or UO_1733 (O_1733,N_14875,N_14948);
or UO_1734 (O_1734,N_14917,N_14912);
nor UO_1735 (O_1735,N_14913,N_14930);
and UO_1736 (O_1736,N_14877,N_14911);
and UO_1737 (O_1737,N_14940,N_14899);
xnor UO_1738 (O_1738,N_14949,N_14942);
xnor UO_1739 (O_1739,N_14939,N_14949);
nor UO_1740 (O_1740,N_14891,N_14961);
xor UO_1741 (O_1741,N_14961,N_14925);
xnor UO_1742 (O_1742,N_14996,N_14877);
or UO_1743 (O_1743,N_14882,N_14875);
nor UO_1744 (O_1744,N_14894,N_14947);
nand UO_1745 (O_1745,N_14906,N_14963);
or UO_1746 (O_1746,N_14939,N_14917);
or UO_1747 (O_1747,N_14958,N_14974);
xnor UO_1748 (O_1748,N_14921,N_14923);
nand UO_1749 (O_1749,N_14945,N_14880);
nor UO_1750 (O_1750,N_14877,N_14965);
or UO_1751 (O_1751,N_14921,N_14877);
nand UO_1752 (O_1752,N_14879,N_14955);
nand UO_1753 (O_1753,N_14885,N_14906);
or UO_1754 (O_1754,N_14908,N_14903);
nand UO_1755 (O_1755,N_14919,N_14941);
xnor UO_1756 (O_1756,N_14881,N_14965);
or UO_1757 (O_1757,N_14948,N_14951);
nand UO_1758 (O_1758,N_14921,N_14936);
xnor UO_1759 (O_1759,N_14957,N_14979);
nand UO_1760 (O_1760,N_14934,N_14942);
and UO_1761 (O_1761,N_14899,N_14990);
and UO_1762 (O_1762,N_14933,N_14923);
and UO_1763 (O_1763,N_14893,N_14997);
nor UO_1764 (O_1764,N_14944,N_14954);
nor UO_1765 (O_1765,N_14997,N_14970);
nor UO_1766 (O_1766,N_14886,N_14876);
and UO_1767 (O_1767,N_14884,N_14887);
nand UO_1768 (O_1768,N_14880,N_14952);
nand UO_1769 (O_1769,N_14944,N_14951);
xor UO_1770 (O_1770,N_14908,N_14925);
and UO_1771 (O_1771,N_14975,N_14964);
nor UO_1772 (O_1772,N_14889,N_14908);
nor UO_1773 (O_1773,N_14878,N_14914);
xor UO_1774 (O_1774,N_14894,N_14936);
nor UO_1775 (O_1775,N_14904,N_14976);
nor UO_1776 (O_1776,N_14941,N_14985);
and UO_1777 (O_1777,N_14975,N_14939);
nor UO_1778 (O_1778,N_14982,N_14945);
and UO_1779 (O_1779,N_14911,N_14938);
nor UO_1780 (O_1780,N_14971,N_14906);
or UO_1781 (O_1781,N_14994,N_14905);
nor UO_1782 (O_1782,N_14905,N_14877);
and UO_1783 (O_1783,N_14963,N_14969);
nor UO_1784 (O_1784,N_14876,N_14917);
and UO_1785 (O_1785,N_14939,N_14900);
nor UO_1786 (O_1786,N_14962,N_14963);
xnor UO_1787 (O_1787,N_14922,N_14944);
or UO_1788 (O_1788,N_14939,N_14902);
and UO_1789 (O_1789,N_14972,N_14940);
and UO_1790 (O_1790,N_14899,N_14978);
nor UO_1791 (O_1791,N_14914,N_14987);
or UO_1792 (O_1792,N_14977,N_14895);
and UO_1793 (O_1793,N_14902,N_14904);
and UO_1794 (O_1794,N_14938,N_14934);
or UO_1795 (O_1795,N_14996,N_14989);
nand UO_1796 (O_1796,N_14961,N_14975);
nand UO_1797 (O_1797,N_14920,N_14991);
nand UO_1798 (O_1798,N_14952,N_14887);
xnor UO_1799 (O_1799,N_14957,N_14907);
nor UO_1800 (O_1800,N_14950,N_14915);
nor UO_1801 (O_1801,N_14887,N_14961);
or UO_1802 (O_1802,N_14936,N_14968);
xor UO_1803 (O_1803,N_14902,N_14987);
and UO_1804 (O_1804,N_14998,N_14903);
nand UO_1805 (O_1805,N_14881,N_14963);
or UO_1806 (O_1806,N_14951,N_14875);
or UO_1807 (O_1807,N_14944,N_14992);
or UO_1808 (O_1808,N_14915,N_14995);
xnor UO_1809 (O_1809,N_14885,N_14973);
and UO_1810 (O_1810,N_14945,N_14925);
nor UO_1811 (O_1811,N_14994,N_14964);
xor UO_1812 (O_1812,N_14888,N_14986);
nor UO_1813 (O_1813,N_14894,N_14964);
xor UO_1814 (O_1814,N_14974,N_14934);
xor UO_1815 (O_1815,N_14981,N_14999);
or UO_1816 (O_1816,N_14991,N_14985);
or UO_1817 (O_1817,N_14958,N_14880);
and UO_1818 (O_1818,N_14933,N_14974);
nor UO_1819 (O_1819,N_14879,N_14989);
xor UO_1820 (O_1820,N_14964,N_14942);
and UO_1821 (O_1821,N_14887,N_14913);
xor UO_1822 (O_1822,N_14923,N_14884);
nor UO_1823 (O_1823,N_14875,N_14979);
or UO_1824 (O_1824,N_14896,N_14924);
and UO_1825 (O_1825,N_14890,N_14955);
nand UO_1826 (O_1826,N_14946,N_14949);
and UO_1827 (O_1827,N_14976,N_14957);
and UO_1828 (O_1828,N_14977,N_14924);
xor UO_1829 (O_1829,N_14918,N_14878);
xor UO_1830 (O_1830,N_14927,N_14890);
xor UO_1831 (O_1831,N_14917,N_14878);
nand UO_1832 (O_1832,N_14921,N_14905);
nand UO_1833 (O_1833,N_14884,N_14891);
or UO_1834 (O_1834,N_14876,N_14922);
or UO_1835 (O_1835,N_14922,N_14930);
or UO_1836 (O_1836,N_14876,N_14942);
xor UO_1837 (O_1837,N_14958,N_14904);
and UO_1838 (O_1838,N_14929,N_14977);
nor UO_1839 (O_1839,N_14911,N_14956);
and UO_1840 (O_1840,N_14968,N_14958);
xnor UO_1841 (O_1841,N_14998,N_14933);
nor UO_1842 (O_1842,N_14975,N_14935);
xnor UO_1843 (O_1843,N_14939,N_14925);
and UO_1844 (O_1844,N_14948,N_14990);
or UO_1845 (O_1845,N_14951,N_14954);
or UO_1846 (O_1846,N_14911,N_14949);
and UO_1847 (O_1847,N_14963,N_14895);
and UO_1848 (O_1848,N_14906,N_14969);
nor UO_1849 (O_1849,N_14929,N_14971);
and UO_1850 (O_1850,N_14976,N_14928);
or UO_1851 (O_1851,N_14929,N_14952);
nand UO_1852 (O_1852,N_14949,N_14875);
nor UO_1853 (O_1853,N_14960,N_14953);
nor UO_1854 (O_1854,N_14916,N_14956);
xnor UO_1855 (O_1855,N_14962,N_14972);
nand UO_1856 (O_1856,N_14986,N_14960);
and UO_1857 (O_1857,N_14944,N_14924);
nand UO_1858 (O_1858,N_14953,N_14986);
nor UO_1859 (O_1859,N_14909,N_14968);
or UO_1860 (O_1860,N_14890,N_14882);
nand UO_1861 (O_1861,N_14988,N_14959);
nand UO_1862 (O_1862,N_14924,N_14926);
xnor UO_1863 (O_1863,N_14882,N_14954);
or UO_1864 (O_1864,N_14908,N_14952);
xor UO_1865 (O_1865,N_14908,N_14898);
and UO_1866 (O_1866,N_14945,N_14917);
or UO_1867 (O_1867,N_14980,N_14927);
xor UO_1868 (O_1868,N_14962,N_14878);
nor UO_1869 (O_1869,N_14976,N_14944);
nor UO_1870 (O_1870,N_14905,N_14971);
xnor UO_1871 (O_1871,N_14906,N_14942);
xnor UO_1872 (O_1872,N_14999,N_14884);
or UO_1873 (O_1873,N_14896,N_14898);
and UO_1874 (O_1874,N_14977,N_14960);
nor UO_1875 (O_1875,N_14905,N_14949);
and UO_1876 (O_1876,N_14969,N_14967);
or UO_1877 (O_1877,N_14912,N_14886);
or UO_1878 (O_1878,N_14931,N_14895);
nand UO_1879 (O_1879,N_14918,N_14927);
nand UO_1880 (O_1880,N_14927,N_14967);
nand UO_1881 (O_1881,N_14904,N_14910);
nand UO_1882 (O_1882,N_14991,N_14934);
and UO_1883 (O_1883,N_14918,N_14966);
and UO_1884 (O_1884,N_14963,N_14933);
or UO_1885 (O_1885,N_14950,N_14907);
xnor UO_1886 (O_1886,N_14907,N_14960);
and UO_1887 (O_1887,N_14909,N_14955);
nor UO_1888 (O_1888,N_14907,N_14951);
and UO_1889 (O_1889,N_14890,N_14983);
or UO_1890 (O_1890,N_14996,N_14918);
nand UO_1891 (O_1891,N_14965,N_14980);
xnor UO_1892 (O_1892,N_14970,N_14994);
or UO_1893 (O_1893,N_14975,N_14907);
nor UO_1894 (O_1894,N_14892,N_14960);
or UO_1895 (O_1895,N_14993,N_14967);
or UO_1896 (O_1896,N_14936,N_14946);
and UO_1897 (O_1897,N_14970,N_14952);
or UO_1898 (O_1898,N_14985,N_14938);
nor UO_1899 (O_1899,N_14878,N_14945);
nor UO_1900 (O_1900,N_14880,N_14950);
nor UO_1901 (O_1901,N_14923,N_14922);
nand UO_1902 (O_1902,N_14990,N_14932);
or UO_1903 (O_1903,N_14908,N_14877);
nor UO_1904 (O_1904,N_14927,N_14976);
or UO_1905 (O_1905,N_14875,N_14910);
nand UO_1906 (O_1906,N_14900,N_14959);
nand UO_1907 (O_1907,N_14930,N_14924);
and UO_1908 (O_1908,N_14975,N_14967);
nor UO_1909 (O_1909,N_14975,N_14880);
and UO_1910 (O_1910,N_14956,N_14955);
xor UO_1911 (O_1911,N_14928,N_14932);
and UO_1912 (O_1912,N_14890,N_14960);
and UO_1913 (O_1913,N_14984,N_14892);
or UO_1914 (O_1914,N_14963,N_14956);
xor UO_1915 (O_1915,N_14910,N_14902);
xnor UO_1916 (O_1916,N_14884,N_14966);
xnor UO_1917 (O_1917,N_14895,N_14927);
xnor UO_1918 (O_1918,N_14923,N_14916);
and UO_1919 (O_1919,N_14889,N_14957);
nand UO_1920 (O_1920,N_14883,N_14889);
nor UO_1921 (O_1921,N_14963,N_14913);
nor UO_1922 (O_1922,N_14891,N_14962);
xor UO_1923 (O_1923,N_14925,N_14937);
nand UO_1924 (O_1924,N_14897,N_14900);
nor UO_1925 (O_1925,N_14915,N_14928);
or UO_1926 (O_1926,N_14978,N_14900);
or UO_1927 (O_1927,N_14909,N_14913);
and UO_1928 (O_1928,N_14952,N_14921);
and UO_1929 (O_1929,N_14993,N_14940);
or UO_1930 (O_1930,N_14905,N_14992);
nand UO_1931 (O_1931,N_14889,N_14951);
or UO_1932 (O_1932,N_14924,N_14981);
and UO_1933 (O_1933,N_14910,N_14964);
and UO_1934 (O_1934,N_14902,N_14961);
nand UO_1935 (O_1935,N_14906,N_14943);
nor UO_1936 (O_1936,N_14896,N_14940);
and UO_1937 (O_1937,N_14953,N_14958);
xnor UO_1938 (O_1938,N_14931,N_14945);
or UO_1939 (O_1939,N_14942,N_14962);
and UO_1940 (O_1940,N_14896,N_14962);
or UO_1941 (O_1941,N_14924,N_14899);
nand UO_1942 (O_1942,N_14902,N_14896);
and UO_1943 (O_1943,N_14952,N_14932);
nand UO_1944 (O_1944,N_14998,N_14987);
nand UO_1945 (O_1945,N_14897,N_14926);
or UO_1946 (O_1946,N_14962,N_14981);
or UO_1947 (O_1947,N_14978,N_14946);
nor UO_1948 (O_1948,N_14901,N_14876);
nor UO_1949 (O_1949,N_14986,N_14937);
or UO_1950 (O_1950,N_14997,N_14960);
or UO_1951 (O_1951,N_14976,N_14885);
and UO_1952 (O_1952,N_14971,N_14937);
nand UO_1953 (O_1953,N_14972,N_14937);
and UO_1954 (O_1954,N_14976,N_14998);
nor UO_1955 (O_1955,N_14895,N_14997);
nor UO_1956 (O_1956,N_14885,N_14891);
xor UO_1957 (O_1957,N_14914,N_14903);
and UO_1958 (O_1958,N_14916,N_14991);
nand UO_1959 (O_1959,N_14876,N_14958);
nand UO_1960 (O_1960,N_14970,N_14914);
and UO_1961 (O_1961,N_14994,N_14962);
nor UO_1962 (O_1962,N_14907,N_14927);
or UO_1963 (O_1963,N_14998,N_14958);
nand UO_1964 (O_1964,N_14917,N_14985);
nand UO_1965 (O_1965,N_14941,N_14928);
nor UO_1966 (O_1966,N_14912,N_14920);
xor UO_1967 (O_1967,N_14943,N_14976);
nor UO_1968 (O_1968,N_14882,N_14978);
or UO_1969 (O_1969,N_14895,N_14926);
xnor UO_1970 (O_1970,N_14912,N_14965);
nor UO_1971 (O_1971,N_14992,N_14911);
nand UO_1972 (O_1972,N_14888,N_14884);
xnor UO_1973 (O_1973,N_14893,N_14878);
nand UO_1974 (O_1974,N_14876,N_14892);
xor UO_1975 (O_1975,N_14878,N_14958);
xnor UO_1976 (O_1976,N_14954,N_14962);
and UO_1977 (O_1977,N_14943,N_14951);
xor UO_1978 (O_1978,N_14997,N_14982);
nand UO_1979 (O_1979,N_14953,N_14903);
nand UO_1980 (O_1980,N_14952,N_14933);
xnor UO_1981 (O_1981,N_14880,N_14903);
xnor UO_1982 (O_1982,N_14984,N_14890);
or UO_1983 (O_1983,N_14998,N_14901);
and UO_1984 (O_1984,N_14899,N_14980);
or UO_1985 (O_1985,N_14980,N_14878);
nor UO_1986 (O_1986,N_14998,N_14986);
nor UO_1987 (O_1987,N_14888,N_14887);
xor UO_1988 (O_1988,N_14980,N_14932);
or UO_1989 (O_1989,N_14955,N_14930);
and UO_1990 (O_1990,N_14924,N_14905);
and UO_1991 (O_1991,N_14920,N_14999);
nand UO_1992 (O_1992,N_14956,N_14929);
and UO_1993 (O_1993,N_14916,N_14922);
nand UO_1994 (O_1994,N_14953,N_14883);
nor UO_1995 (O_1995,N_14985,N_14983);
and UO_1996 (O_1996,N_14963,N_14917);
and UO_1997 (O_1997,N_14975,N_14977);
or UO_1998 (O_1998,N_14923,N_14931);
and UO_1999 (O_1999,N_14978,N_14881);
endmodule