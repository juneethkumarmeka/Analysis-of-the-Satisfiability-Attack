module basic_1000_10000_1500_4_levels_2xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_801,In_236);
and U1 (N_1,In_508,In_332);
and U2 (N_2,In_609,In_80);
and U3 (N_3,In_139,In_378);
nor U4 (N_4,In_754,In_631);
nand U5 (N_5,In_322,In_420);
nor U6 (N_6,In_253,In_862);
nand U7 (N_7,In_742,In_866);
nor U8 (N_8,In_169,In_324);
or U9 (N_9,In_677,In_524);
and U10 (N_10,In_611,In_816);
or U11 (N_11,In_91,In_724);
and U12 (N_12,In_585,In_164);
nand U13 (N_13,In_314,In_81);
nand U14 (N_14,In_304,In_534);
and U15 (N_15,In_851,In_713);
nor U16 (N_16,In_550,In_708);
xnor U17 (N_17,In_899,In_487);
nand U18 (N_18,In_868,In_285);
nor U19 (N_19,In_403,In_785);
or U20 (N_20,In_988,In_786);
or U21 (N_21,In_367,In_523);
and U22 (N_22,In_340,In_500);
nand U23 (N_23,In_654,In_860);
or U24 (N_24,In_728,In_835);
nand U25 (N_25,In_318,In_774);
and U26 (N_26,In_796,In_50);
or U27 (N_27,In_41,In_651);
or U28 (N_28,In_597,In_771);
nand U29 (N_29,In_592,In_414);
nor U30 (N_30,In_748,In_961);
nand U31 (N_31,In_457,In_507);
nand U32 (N_32,In_845,In_445);
and U33 (N_33,In_14,In_413);
nand U34 (N_34,In_308,In_738);
nand U35 (N_35,In_619,In_687);
or U36 (N_36,In_944,In_985);
nand U37 (N_37,In_389,In_875);
and U38 (N_38,In_973,In_642);
and U39 (N_39,In_702,In_662);
or U40 (N_40,In_813,In_810);
or U41 (N_41,In_473,In_474);
or U42 (N_42,In_426,In_995);
nor U43 (N_43,In_564,In_543);
or U44 (N_44,In_26,In_815);
and U45 (N_45,In_805,In_496);
and U46 (N_46,In_260,In_12);
nor U47 (N_47,In_760,In_512);
nand U48 (N_48,In_681,In_269);
nor U49 (N_49,In_549,In_187);
nand U50 (N_50,In_204,In_514);
nand U51 (N_51,In_522,In_369);
nand U52 (N_52,In_896,In_935);
nor U53 (N_53,In_203,In_34);
nand U54 (N_54,In_122,In_622);
nor U55 (N_55,In_69,In_215);
nor U56 (N_56,In_730,In_674);
or U57 (N_57,In_453,In_917);
nand U58 (N_58,In_154,In_115);
nor U59 (N_59,In_615,In_610);
nor U60 (N_60,In_948,In_630);
nand U61 (N_61,In_600,In_823);
or U62 (N_62,In_411,In_872);
nand U63 (N_63,In_443,In_763);
and U64 (N_64,In_104,In_562);
or U65 (N_65,In_761,In_464);
and U66 (N_66,In_53,In_979);
nand U67 (N_67,In_33,In_209);
or U68 (N_68,In_377,In_42);
or U69 (N_69,In_374,In_305);
nand U70 (N_70,In_999,In_72);
nor U71 (N_71,In_538,In_177);
xnor U72 (N_72,In_319,In_697);
nand U73 (N_73,In_804,In_497);
nand U74 (N_74,In_782,In_199);
and U75 (N_75,In_167,In_108);
and U76 (N_76,In_827,In_479);
nand U77 (N_77,In_298,In_941);
nor U78 (N_78,In_21,In_229);
nand U79 (N_79,In_31,In_808);
nand U80 (N_80,In_330,In_221);
nand U81 (N_81,In_818,In_650);
and U82 (N_82,In_223,In_297);
or U83 (N_83,In_58,In_323);
and U84 (N_84,In_879,In_688);
or U85 (N_85,In_39,In_280);
or U86 (N_86,In_36,In_670);
and U87 (N_87,In_641,In_155);
or U88 (N_88,In_248,In_405);
nor U89 (N_89,In_30,In_547);
nand U90 (N_90,In_397,In_66);
or U91 (N_91,In_235,In_894);
nor U92 (N_92,In_214,In_859);
nor U93 (N_93,In_345,In_501);
xor U94 (N_94,In_124,In_173);
nand U95 (N_95,In_238,In_387);
and U96 (N_96,In_923,In_201);
and U97 (N_97,In_275,In_869);
or U98 (N_98,In_698,In_920);
nand U99 (N_99,In_380,In_213);
nor U100 (N_100,In_532,In_711);
or U101 (N_101,In_784,In_125);
nand U102 (N_102,In_205,In_766);
nand U103 (N_103,In_942,In_998);
and U104 (N_104,In_567,In_352);
nor U105 (N_105,In_437,In_890);
nor U106 (N_106,In_188,In_829);
or U107 (N_107,In_32,In_976);
nand U108 (N_108,In_695,In_914);
and U109 (N_109,In_718,In_360);
nor U110 (N_110,In_370,In_439);
or U111 (N_111,In_165,In_373);
and U112 (N_112,In_136,In_245);
and U113 (N_113,In_661,In_44);
nand U114 (N_114,In_971,In_266);
nand U115 (N_115,In_519,In_423);
or U116 (N_116,In_858,In_166);
or U117 (N_117,In_462,In_54);
nand U118 (N_118,In_310,In_779);
and U119 (N_119,In_338,In_720);
and U120 (N_120,In_412,In_328);
nand U121 (N_121,In_753,In_329);
nor U122 (N_122,In_839,In_660);
xor U123 (N_123,In_447,In_48);
and U124 (N_124,In_85,In_398);
or U125 (N_125,In_283,In_905);
nor U126 (N_126,In_440,In_797);
xor U127 (N_127,In_406,In_157);
xnor U128 (N_128,In_780,In_545);
nand U129 (N_129,In_251,In_602);
and U130 (N_130,In_491,In_381);
or U131 (N_131,In_361,In_312);
or U132 (N_132,In_883,In_561);
nand U133 (N_133,In_530,In_581);
nand U134 (N_134,In_231,In_133);
nor U135 (N_135,In_488,In_960);
and U136 (N_136,In_655,In_832);
nand U137 (N_137,In_132,In_593);
nand U138 (N_138,In_734,In_653);
nand U139 (N_139,In_791,In_364);
and U140 (N_140,In_798,In_599);
nor U141 (N_141,In_142,In_723);
and U142 (N_142,In_901,In_13);
nand U143 (N_143,In_938,In_645);
nor U144 (N_144,In_294,In_25);
or U145 (N_145,In_475,In_395);
and U146 (N_146,In_588,In_127);
nor U147 (N_147,In_983,In_388);
or U148 (N_148,In_636,In_882);
nand U149 (N_149,In_230,In_986);
nand U150 (N_150,In_929,In_402);
and U151 (N_151,In_232,In_925);
or U152 (N_152,In_764,In_624);
nand U153 (N_153,In_924,In_20);
or U154 (N_154,In_415,In_646);
nor U155 (N_155,In_943,In_331);
or U156 (N_156,In_955,In_671);
nand U157 (N_157,In_633,In_657);
nand U158 (N_158,In_461,In_281);
nand U159 (N_159,In_239,In_277);
and U160 (N_160,In_65,In_975);
nand U161 (N_161,In_559,In_595);
nand U162 (N_162,In_958,In_151);
and U163 (N_163,In_493,In_171);
and U164 (N_164,In_162,In_981);
nand U165 (N_165,In_974,In_28);
and U166 (N_166,In_416,In_358);
nand U167 (N_167,In_504,In_994);
nand U168 (N_168,In_70,In_517);
nor U169 (N_169,In_296,In_259);
nor U170 (N_170,In_793,In_47);
or U171 (N_171,In_852,In_696);
nand U172 (N_172,In_705,In_746);
and U173 (N_173,In_825,In_563);
nor U174 (N_174,In_962,In_977);
or U175 (N_175,In_685,In_15);
nand U176 (N_176,In_997,In_385);
nand U177 (N_177,In_427,In_144);
nor U178 (N_178,In_190,In_834);
and U179 (N_179,In_227,In_152);
nand U180 (N_180,In_57,In_349);
or U181 (N_181,In_105,In_417);
nor U182 (N_182,In_356,In_964);
xnor U183 (N_183,In_638,In_972);
nor U184 (N_184,In_989,In_46);
or U185 (N_185,In_254,In_806);
nor U186 (N_186,In_98,In_116);
or U187 (N_187,In_744,In_515);
nor U188 (N_188,In_52,In_623);
or U189 (N_189,In_114,In_586);
nor U190 (N_190,In_918,In_608);
nand U191 (N_191,In_1,In_568);
nor U192 (N_192,In_438,In_126);
nand U193 (N_193,In_419,In_528);
nand U194 (N_194,In_913,In_591);
and U195 (N_195,In_811,In_196);
nand U196 (N_196,In_891,In_980);
and U197 (N_197,In_518,In_68);
or U198 (N_198,In_502,In_659);
and U199 (N_199,In_250,In_353);
and U200 (N_200,In_300,In_857);
or U201 (N_201,In_278,In_295);
and U202 (N_202,In_676,In_284);
xnor U203 (N_203,In_893,In_481);
nor U204 (N_204,In_170,In_27);
nor U205 (N_205,In_612,In_881);
and U206 (N_206,In_912,In_892);
or U207 (N_207,In_526,In_8);
or U208 (N_208,In_452,In_272);
xnor U209 (N_209,In_101,In_573);
and U210 (N_210,In_301,In_89);
or U211 (N_211,In_922,In_635);
or U212 (N_212,In_768,In_767);
and U213 (N_213,In_428,In_788);
nand U214 (N_214,In_178,In_529);
or U215 (N_215,In_191,In_510);
or U216 (N_216,In_544,In_429);
and U217 (N_217,In_197,In_366);
and U218 (N_218,In_990,In_712);
and U219 (N_219,In_148,In_978);
or U220 (N_220,In_341,In_665);
and U221 (N_221,In_343,In_97);
nand U222 (N_222,In_795,In_505);
nor U223 (N_223,In_639,In_939);
nand U224 (N_224,In_601,In_582);
nor U225 (N_225,In_625,In_926);
nor U226 (N_226,In_949,In_194);
nand U227 (N_227,In_874,In_449);
or U228 (N_228,In_480,In_172);
or U229 (N_229,In_992,In_903);
or U230 (N_230,In_828,In_790);
nor U231 (N_231,In_743,In_220);
nor U232 (N_232,In_29,In_865);
or U233 (N_233,In_119,In_287);
or U234 (N_234,In_668,In_889);
nand U235 (N_235,In_261,In_90);
nor U236 (N_236,In_919,In_404);
or U237 (N_237,In_817,In_555);
and U238 (N_238,In_193,In_431);
or U239 (N_239,In_158,In_807);
or U240 (N_240,In_679,In_478);
and U241 (N_241,In_103,In_584);
nor U242 (N_242,In_770,In_870);
xnor U243 (N_243,In_887,In_485);
or U244 (N_244,In_459,In_574);
and U245 (N_245,In_721,In_113);
nor U246 (N_246,In_598,In_489);
or U247 (N_247,In_135,In_831);
nor U248 (N_248,In_513,In_906);
or U249 (N_249,In_970,In_548);
and U250 (N_250,In_210,In_921);
and U251 (N_251,In_847,In_226);
and U252 (N_252,In_557,In_940);
and U253 (N_253,In_384,In_854);
nor U254 (N_254,In_700,In_359);
nand U255 (N_255,In_620,In_321);
nand U256 (N_256,In_762,In_930);
nor U257 (N_257,In_495,In_741);
nor U258 (N_258,In_302,In_701);
nor U259 (N_259,In_855,In_731);
nor U260 (N_260,In_690,In_430);
nor U261 (N_261,In_460,In_647);
nor U262 (N_262,In_79,In_9);
nor U263 (N_263,In_556,In_183);
or U264 (N_264,In_969,In_252);
nand U265 (N_265,In_794,In_182);
nor U266 (N_266,In_184,In_673);
and U267 (N_267,In_118,In_732);
nand U268 (N_268,In_932,In_401);
or U269 (N_269,In_535,In_327);
or U270 (N_270,In_527,In_106);
nand U271 (N_271,In_725,In_908);
nor U272 (N_272,In_993,In_552);
nand U273 (N_273,In_264,In_963);
nand U274 (N_274,In_802,In_45);
nand U275 (N_275,In_207,In_107);
and U276 (N_276,In_265,In_627);
nor U277 (N_277,In_289,In_849);
nor U278 (N_278,In_7,In_910);
and U279 (N_279,In_575,In_477);
nor U280 (N_280,In_604,In_506);
or U281 (N_281,In_216,In_957);
nor U282 (N_282,In_335,In_355);
xor U283 (N_283,In_59,In_363);
and U284 (N_284,In_717,In_709);
xnor U285 (N_285,In_76,In_863);
xnor U286 (N_286,In_451,In_803);
nor U287 (N_287,In_648,In_160);
nand U288 (N_288,In_315,In_288);
nor U289 (N_289,In_484,In_904);
nor U290 (N_290,In_886,In_463);
nor U291 (N_291,In_86,In_735);
nor U292 (N_292,In_159,In_382);
nand U293 (N_293,In_937,In_521);
nor U294 (N_294,In_982,In_407);
nand U295 (N_295,In_87,In_390);
nand U296 (N_296,In_109,In_826);
nor U297 (N_297,In_391,In_821);
nor U298 (N_298,In_234,In_987);
or U299 (N_299,In_536,In_590);
or U300 (N_300,In_640,In_628);
nor U301 (N_301,In_486,In_848);
nand U302 (N_302,In_822,In_750);
nor U303 (N_303,In_316,In_492);
nand U304 (N_304,In_306,In_82);
nor U305 (N_305,In_35,In_375);
nand U306 (N_306,In_836,In_436);
nand U307 (N_307,In_565,In_897);
and U308 (N_308,In_719,In_967);
or U309 (N_309,In_605,In_222);
nand U310 (N_310,In_773,In_634);
nor U311 (N_311,In_161,In_649);
nor U312 (N_312,In_703,In_393);
and U313 (N_313,In_11,In_120);
nor U314 (N_314,In_444,In_189);
or U315 (N_315,In_291,In_394);
nor U316 (N_316,In_455,In_928);
and U317 (N_317,In_663,In_309);
or U318 (N_318,In_837,In_200);
nor U319 (N_319,In_3,In_809);
nor U320 (N_320,In_137,In_174);
nand U321 (N_321,In_10,In_965);
nand U322 (N_322,In_511,In_800);
or U323 (N_323,In_678,In_185);
and U324 (N_324,In_344,In_606);
nor U325 (N_325,In_64,In_726);
nand U326 (N_326,In_242,In_362);
xor U327 (N_327,In_727,In_273);
or U328 (N_328,In_707,In_838);
and U329 (N_329,In_691,In_441);
nor U330 (N_330,In_243,In_596);
nand U331 (N_331,In_952,In_716);
or U332 (N_332,In_579,In_694);
or U333 (N_333,In_799,In_656);
nand U334 (N_334,In_664,In_249);
nor U335 (N_335,In_643,In_931);
nand U336 (N_336,In_617,In_885);
nand U337 (N_337,In_350,In_129);
and U338 (N_338,In_739,In_933);
or U339 (N_339,In_442,In_146);
or U340 (N_340,In_421,In_792);
and U341 (N_341,In_409,In_570);
or U342 (N_342,In_311,In_888);
or U343 (N_343,In_755,In_777);
nand U344 (N_344,In_583,In_945);
and U345 (N_345,In_299,In_757);
nand U346 (N_346,In_840,In_775);
nand U347 (N_347,In_824,In_379);
and U348 (N_348,In_372,In_386);
nand U349 (N_349,In_895,In_334);
and U350 (N_350,In_909,In_680);
and U351 (N_351,In_482,In_40);
xnor U352 (N_352,In_307,In_399);
and U353 (N_353,In_776,In_19);
or U354 (N_354,In_73,In_898);
nor U355 (N_355,In_102,In_410);
xor U356 (N_356,In_78,In_873);
nand U357 (N_357,In_141,In_286);
or U358 (N_358,In_537,In_934);
nor U359 (N_359,In_94,In_880);
and U360 (N_360,In_163,In_542);
nor U361 (N_361,In_953,In_467);
nand U362 (N_362,In_192,In_371);
nor U363 (N_363,In_326,In_589);
and U364 (N_364,In_130,In_408);
and U365 (N_365,In_594,In_469);
and U366 (N_366,In_846,In_787);
nand U367 (N_367,In_911,In_244);
or U368 (N_368,In_652,In_733);
and U369 (N_369,In_729,In_74);
nor U370 (N_370,In_186,In_333);
nor U371 (N_371,In_927,In_95);
or U372 (N_372,In_233,In_769);
or U373 (N_373,In_131,In_271);
and U374 (N_374,In_217,In_218);
or U375 (N_375,In_454,In_644);
and U376 (N_376,In_490,In_110);
nand U377 (N_377,In_268,In_684);
nand U378 (N_378,In_77,In_675);
nand U379 (N_379,In_317,In_546);
and U380 (N_380,In_348,In_56);
or U381 (N_381,In_117,In_17);
nor U382 (N_382,In_145,In_293);
nor U383 (N_383,In_458,In_722);
and U384 (N_384,In_257,In_616);
xor U385 (N_385,In_814,In_736);
nor U386 (N_386,In_476,In_580);
and U387 (N_387,In_282,In_637);
or U388 (N_388,In_554,In_339);
or U389 (N_389,In_551,In_667);
nor U390 (N_390,In_202,In_60);
nand U391 (N_391,In_448,In_621);
or U392 (N_392,In_270,In_699);
nor U393 (N_393,In_759,In_950);
and U394 (N_394,In_778,In_228);
or U395 (N_395,In_153,In_842);
or U396 (N_396,In_195,In_996);
xnor U397 (N_397,In_255,In_368);
nand U398 (N_398,In_632,In_765);
and U399 (N_399,In_258,In_710);
and U400 (N_400,In_871,In_540);
nand U401 (N_401,In_149,In_128);
and U402 (N_402,In_772,In_830);
nor U403 (N_403,In_539,In_789);
and U404 (N_404,In_751,In_181);
and U405 (N_405,In_38,In_256);
and U406 (N_406,In_470,In_351);
nand U407 (N_407,In_347,In_396);
and U408 (N_408,In_237,In_61);
or U409 (N_409,In_465,In_841);
or U410 (N_410,In_706,In_346);
or U411 (N_411,In_520,In_820);
nand U412 (N_412,In_947,In_5);
and U413 (N_413,In_587,In_576);
nor U414 (N_414,In_179,In_566);
nor U415 (N_415,In_951,In_224);
or U416 (N_416,In_629,In_686);
and U417 (N_417,In_93,In_626);
and U418 (N_418,In_867,In_320);
nand U419 (N_419,In_241,In_211);
nor U420 (N_420,In_812,In_432);
or U421 (N_421,In_6,In_92);
or U422 (N_422,In_84,In_682);
or U423 (N_423,In_422,In_499);
nor U424 (N_424,In_850,In_354);
nor U425 (N_425,In_946,In_498);
or U426 (N_426,In_915,In_614);
and U427 (N_427,In_2,In_111);
and U428 (N_428,In_666,In_737);
nor U429 (N_429,In_456,In_844);
or U430 (N_430,In_376,In_861);
and U431 (N_431,In_740,In_435);
or U432 (N_432,In_819,In_246);
nor U433 (N_433,In_365,In_569);
and U434 (N_434,In_672,In_756);
nor U435 (N_435,In_531,In_433);
nor U436 (N_436,In_541,In_0);
or U437 (N_437,In_878,In_276);
nor U438 (N_438,In_876,In_856);
or U439 (N_439,In_704,In_516);
nand U440 (N_440,In_884,In_418);
nand U441 (N_441,In_446,In_175);
nor U442 (N_442,In_150,In_279);
and U443 (N_443,In_37,In_212);
or U444 (N_444,In_247,In_24);
or U445 (N_445,In_483,In_325);
or U446 (N_446,In_22,In_83);
nand U447 (N_447,In_425,In_558);
or U448 (N_448,In_134,In_240);
nand U449 (N_449,In_864,In_168);
and U450 (N_450,In_342,In_156);
nor U451 (N_451,In_336,In_303);
nor U452 (N_452,In_900,In_603);
or U453 (N_453,In_902,In_968);
or U454 (N_454,In_121,In_553);
or U455 (N_455,In_71,In_509);
and U456 (N_456,In_745,In_400);
or U457 (N_457,In_693,In_833);
and U458 (N_458,In_466,In_607);
nand U459 (N_459,In_692,In_143);
nor U460 (N_460,In_337,In_63);
nand U461 (N_461,In_225,In_503);
nand U462 (N_462,In_262,In_494);
and U463 (N_463,In_450,In_781);
nor U464 (N_464,In_783,In_560);
or U465 (N_465,In_62,In_472);
nand U466 (N_466,In_434,In_984);
nor U467 (N_467,In_747,In_16);
nand U468 (N_468,In_267,In_18);
nor U469 (N_469,In_274,In_43);
nand U470 (N_470,In_916,In_140);
nor U471 (N_471,In_843,In_613);
nand U472 (N_472,In_424,In_689);
and U473 (N_473,In_758,In_956);
nand U474 (N_474,In_147,In_525);
nor U475 (N_475,In_715,In_96);
nor U476 (N_476,In_749,In_112);
nand U477 (N_477,In_936,In_683);
or U478 (N_478,In_138,In_577);
nor U479 (N_479,In_313,In_23);
nor U480 (N_480,In_292,In_578);
nand U481 (N_481,In_572,In_383);
nor U482 (N_482,In_714,In_180);
nand U483 (N_483,In_4,In_471);
nor U484 (N_484,In_959,In_392);
and U485 (N_485,In_954,In_571);
or U486 (N_486,In_357,In_877);
or U487 (N_487,In_658,In_206);
and U488 (N_488,In_991,In_176);
nand U489 (N_489,In_75,In_290);
nand U490 (N_490,In_67,In_100);
and U491 (N_491,In_468,In_88);
nand U492 (N_492,In_51,In_99);
and U493 (N_493,In_123,In_198);
and U494 (N_494,In_208,In_966);
and U495 (N_495,In_618,In_853);
nand U496 (N_496,In_49,In_752);
nor U497 (N_497,In_669,In_219);
nor U498 (N_498,In_533,In_55);
or U499 (N_499,In_263,In_907);
or U500 (N_500,In_976,In_85);
nand U501 (N_501,In_109,In_710);
and U502 (N_502,In_241,In_601);
nor U503 (N_503,In_342,In_811);
and U504 (N_504,In_842,In_970);
nand U505 (N_505,In_346,In_761);
xnor U506 (N_506,In_494,In_113);
nor U507 (N_507,In_39,In_630);
nand U508 (N_508,In_997,In_277);
nor U509 (N_509,In_960,In_17);
xnor U510 (N_510,In_59,In_719);
or U511 (N_511,In_854,In_201);
nor U512 (N_512,In_441,In_646);
nor U513 (N_513,In_574,In_737);
and U514 (N_514,In_409,In_671);
and U515 (N_515,In_476,In_597);
and U516 (N_516,In_87,In_232);
xor U517 (N_517,In_812,In_332);
nor U518 (N_518,In_371,In_474);
and U519 (N_519,In_358,In_633);
or U520 (N_520,In_71,In_197);
nand U521 (N_521,In_231,In_225);
or U522 (N_522,In_732,In_571);
nor U523 (N_523,In_279,In_564);
and U524 (N_524,In_757,In_567);
nor U525 (N_525,In_812,In_740);
nor U526 (N_526,In_322,In_315);
or U527 (N_527,In_62,In_142);
and U528 (N_528,In_809,In_939);
and U529 (N_529,In_661,In_611);
or U530 (N_530,In_3,In_19);
and U531 (N_531,In_260,In_90);
nand U532 (N_532,In_941,In_188);
nor U533 (N_533,In_635,In_263);
nor U534 (N_534,In_785,In_998);
nor U535 (N_535,In_119,In_990);
nor U536 (N_536,In_657,In_587);
and U537 (N_537,In_462,In_177);
nand U538 (N_538,In_853,In_539);
and U539 (N_539,In_275,In_208);
or U540 (N_540,In_415,In_533);
and U541 (N_541,In_916,In_166);
nor U542 (N_542,In_229,In_252);
nand U543 (N_543,In_942,In_943);
or U544 (N_544,In_564,In_695);
nor U545 (N_545,In_264,In_944);
and U546 (N_546,In_501,In_793);
nand U547 (N_547,In_809,In_706);
nand U548 (N_548,In_427,In_242);
nor U549 (N_549,In_422,In_905);
and U550 (N_550,In_93,In_35);
nand U551 (N_551,In_737,In_103);
or U552 (N_552,In_939,In_14);
nand U553 (N_553,In_468,In_367);
nor U554 (N_554,In_634,In_194);
or U555 (N_555,In_903,In_770);
xor U556 (N_556,In_765,In_376);
nand U557 (N_557,In_43,In_166);
or U558 (N_558,In_301,In_14);
and U559 (N_559,In_960,In_468);
and U560 (N_560,In_415,In_745);
or U561 (N_561,In_40,In_567);
and U562 (N_562,In_211,In_121);
or U563 (N_563,In_487,In_533);
and U564 (N_564,In_129,In_247);
nand U565 (N_565,In_654,In_376);
or U566 (N_566,In_666,In_202);
or U567 (N_567,In_773,In_702);
or U568 (N_568,In_578,In_352);
nand U569 (N_569,In_481,In_643);
xnor U570 (N_570,In_561,In_634);
and U571 (N_571,In_495,In_908);
and U572 (N_572,In_594,In_979);
nor U573 (N_573,In_436,In_183);
and U574 (N_574,In_986,In_456);
nand U575 (N_575,In_426,In_14);
or U576 (N_576,In_791,In_365);
or U577 (N_577,In_657,In_27);
nand U578 (N_578,In_564,In_498);
and U579 (N_579,In_154,In_101);
nand U580 (N_580,In_973,In_862);
nand U581 (N_581,In_209,In_86);
nand U582 (N_582,In_134,In_908);
nor U583 (N_583,In_373,In_784);
or U584 (N_584,In_36,In_388);
nand U585 (N_585,In_367,In_482);
nor U586 (N_586,In_668,In_569);
and U587 (N_587,In_533,In_309);
and U588 (N_588,In_993,In_352);
and U589 (N_589,In_331,In_788);
or U590 (N_590,In_102,In_480);
or U591 (N_591,In_850,In_449);
nor U592 (N_592,In_132,In_697);
nand U593 (N_593,In_658,In_485);
or U594 (N_594,In_375,In_819);
or U595 (N_595,In_475,In_206);
or U596 (N_596,In_433,In_165);
xor U597 (N_597,In_836,In_459);
xnor U598 (N_598,In_517,In_98);
nor U599 (N_599,In_432,In_72);
nor U600 (N_600,In_231,In_98);
and U601 (N_601,In_896,In_491);
and U602 (N_602,In_387,In_535);
nand U603 (N_603,In_213,In_210);
nand U604 (N_604,In_911,In_791);
or U605 (N_605,In_315,In_992);
or U606 (N_606,In_85,In_538);
nand U607 (N_607,In_850,In_807);
nor U608 (N_608,In_272,In_48);
or U609 (N_609,In_674,In_692);
nor U610 (N_610,In_501,In_231);
and U611 (N_611,In_148,In_366);
and U612 (N_612,In_963,In_747);
and U613 (N_613,In_569,In_257);
nand U614 (N_614,In_579,In_91);
nor U615 (N_615,In_118,In_901);
or U616 (N_616,In_875,In_723);
or U617 (N_617,In_127,In_276);
or U618 (N_618,In_133,In_792);
nor U619 (N_619,In_988,In_842);
and U620 (N_620,In_623,In_73);
or U621 (N_621,In_50,In_769);
and U622 (N_622,In_291,In_108);
nor U623 (N_623,In_167,In_976);
nor U624 (N_624,In_385,In_769);
nand U625 (N_625,In_116,In_890);
nor U626 (N_626,In_473,In_721);
and U627 (N_627,In_933,In_229);
or U628 (N_628,In_748,In_154);
nor U629 (N_629,In_668,In_541);
nand U630 (N_630,In_917,In_206);
and U631 (N_631,In_281,In_215);
nor U632 (N_632,In_561,In_805);
and U633 (N_633,In_335,In_71);
nor U634 (N_634,In_219,In_407);
and U635 (N_635,In_342,In_683);
nand U636 (N_636,In_538,In_286);
xnor U637 (N_637,In_379,In_487);
or U638 (N_638,In_220,In_592);
or U639 (N_639,In_150,In_788);
nor U640 (N_640,In_789,In_553);
xnor U641 (N_641,In_426,In_691);
nor U642 (N_642,In_665,In_780);
nand U643 (N_643,In_448,In_762);
nor U644 (N_644,In_840,In_550);
or U645 (N_645,In_454,In_381);
nand U646 (N_646,In_973,In_305);
nor U647 (N_647,In_807,In_354);
nand U648 (N_648,In_695,In_16);
or U649 (N_649,In_586,In_321);
or U650 (N_650,In_247,In_270);
nor U651 (N_651,In_72,In_583);
nor U652 (N_652,In_367,In_92);
nor U653 (N_653,In_605,In_247);
nor U654 (N_654,In_519,In_43);
nand U655 (N_655,In_804,In_310);
nand U656 (N_656,In_116,In_889);
or U657 (N_657,In_73,In_540);
nand U658 (N_658,In_42,In_415);
and U659 (N_659,In_141,In_240);
and U660 (N_660,In_771,In_429);
and U661 (N_661,In_50,In_423);
or U662 (N_662,In_890,In_209);
or U663 (N_663,In_873,In_502);
nand U664 (N_664,In_951,In_785);
and U665 (N_665,In_764,In_907);
nand U666 (N_666,In_447,In_457);
nor U667 (N_667,In_323,In_555);
nand U668 (N_668,In_131,In_829);
or U669 (N_669,In_73,In_455);
nand U670 (N_670,In_541,In_548);
or U671 (N_671,In_278,In_725);
or U672 (N_672,In_278,In_414);
nand U673 (N_673,In_479,In_717);
nor U674 (N_674,In_135,In_468);
nand U675 (N_675,In_742,In_920);
and U676 (N_676,In_278,In_540);
and U677 (N_677,In_754,In_972);
nor U678 (N_678,In_396,In_490);
nor U679 (N_679,In_663,In_886);
or U680 (N_680,In_457,In_703);
nand U681 (N_681,In_2,In_702);
or U682 (N_682,In_437,In_994);
and U683 (N_683,In_639,In_133);
nand U684 (N_684,In_818,In_133);
or U685 (N_685,In_756,In_987);
and U686 (N_686,In_737,In_804);
nor U687 (N_687,In_442,In_447);
nand U688 (N_688,In_994,In_764);
xnor U689 (N_689,In_820,In_921);
and U690 (N_690,In_177,In_778);
nand U691 (N_691,In_261,In_288);
nand U692 (N_692,In_725,In_839);
nor U693 (N_693,In_542,In_527);
or U694 (N_694,In_397,In_387);
nand U695 (N_695,In_443,In_793);
nand U696 (N_696,In_340,In_905);
and U697 (N_697,In_425,In_961);
and U698 (N_698,In_995,In_126);
and U699 (N_699,In_498,In_493);
and U700 (N_700,In_153,In_378);
or U701 (N_701,In_622,In_849);
or U702 (N_702,In_225,In_732);
or U703 (N_703,In_278,In_565);
nor U704 (N_704,In_691,In_918);
nor U705 (N_705,In_165,In_854);
and U706 (N_706,In_821,In_780);
nor U707 (N_707,In_229,In_40);
nor U708 (N_708,In_110,In_527);
and U709 (N_709,In_522,In_854);
or U710 (N_710,In_877,In_276);
nand U711 (N_711,In_562,In_833);
nor U712 (N_712,In_996,In_53);
or U713 (N_713,In_874,In_737);
or U714 (N_714,In_773,In_537);
or U715 (N_715,In_189,In_14);
or U716 (N_716,In_382,In_817);
nor U717 (N_717,In_752,In_744);
or U718 (N_718,In_68,In_557);
nor U719 (N_719,In_502,In_338);
and U720 (N_720,In_68,In_901);
nand U721 (N_721,In_438,In_614);
and U722 (N_722,In_827,In_708);
nand U723 (N_723,In_942,In_944);
and U724 (N_724,In_428,In_552);
nand U725 (N_725,In_446,In_821);
or U726 (N_726,In_531,In_914);
nand U727 (N_727,In_304,In_602);
or U728 (N_728,In_634,In_662);
nand U729 (N_729,In_965,In_540);
nand U730 (N_730,In_244,In_353);
nor U731 (N_731,In_933,In_829);
nand U732 (N_732,In_974,In_931);
and U733 (N_733,In_391,In_297);
nand U734 (N_734,In_110,In_572);
nor U735 (N_735,In_270,In_584);
nor U736 (N_736,In_681,In_725);
or U737 (N_737,In_126,In_889);
nor U738 (N_738,In_507,In_383);
and U739 (N_739,In_954,In_181);
or U740 (N_740,In_311,In_6);
or U741 (N_741,In_250,In_495);
nor U742 (N_742,In_990,In_738);
nand U743 (N_743,In_513,In_814);
and U744 (N_744,In_866,In_838);
nand U745 (N_745,In_730,In_354);
nor U746 (N_746,In_584,In_553);
nand U747 (N_747,In_574,In_764);
or U748 (N_748,In_411,In_846);
nor U749 (N_749,In_9,In_676);
nor U750 (N_750,In_277,In_319);
and U751 (N_751,In_249,In_650);
nor U752 (N_752,In_211,In_25);
xor U753 (N_753,In_386,In_960);
or U754 (N_754,In_865,In_70);
or U755 (N_755,In_715,In_632);
nor U756 (N_756,In_549,In_135);
xor U757 (N_757,In_939,In_587);
nand U758 (N_758,In_765,In_325);
or U759 (N_759,In_108,In_31);
nor U760 (N_760,In_677,In_562);
or U761 (N_761,In_947,In_887);
nand U762 (N_762,In_502,In_534);
or U763 (N_763,In_728,In_931);
nand U764 (N_764,In_163,In_711);
nand U765 (N_765,In_999,In_291);
or U766 (N_766,In_960,In_599);
or U767 (N_767,In_932,In_154);
and U768 (N_768,In_370,In_150);
and U769 (N_769,In_940,In_587);
nor U770 (N_770,In_3,In_907);
nand U771 (N_771,In_649,In_208);
nor U772 (N_772,In_109,In_200);
or U773 (N_773,In_412,In_303);
nor U774 (N_774,In_487,In_310);
xnor U775 (N_775,In_693,In_930);
nor U776 (N_776,In_885,In_133);
or U777 (N_777,In_207,In_686);
nand U778 (N_778,In_603,In_485);
or U779 (N_779,In_730,In_575);
nand U780 (N_780,In_388,In_316);
and U781 (N_781,In_103,In_147);
nor U782 (N_782,In_558,In_854);
or U783 (N_783,In_386,In_178);
nor U784 (N_784,In_271,In_240);
or U785 (N_785,In_343,In_205);
or U786 (N_786,In_178,In_597);
and U787 (N_787,In_327,In_898);
nor U788 (N_788,In_497,In_123);
and U789 (N_789,In_898,In_864);
or U790 (N_790,In_758,In_90);
nor U791 (N_791,In_650,In_317);
or U792 (N_792,In_785,In_654);
and U793 (N_793,In_42,In_295);
or U794 (N_794,In_409,In_418);
nor U795 (N_795,In_609,In_961);
nor U796 (N_796,In_742,In_211);
nand U797 (N_797,In_833,In_250);
or U798 (N_798,In_60,In_110);
nor U799 (N_799,In_943,In_716);
and U800 (N_800,In_163,In_76);
xnor U801 (N_801,In_987,In_509);
and U802 (N_802,In_587,In_392);
nor U803 (N_803,In_238,In_949);
and U804 (N_804,In_165,In_836);
and U805 (N_805,In_803,In_89);
nand U806 (N_806,In_301,In_715);
and U807 (N_807,In_760,In_488);
or U808 (N_808,In_965,In_389);
nand U809 (N_809,In_142,In_814);
and U810 (N_810,In_858,In_26);
nand U811 (N_811,In_807,In_907);
and U812 (N_812,In_761,In_131);
xor U813 (N_813,In_376,In_643);
or U814 (N_814,In_190,In_104);
or U815 (N_815,In_391,In_872);
or U816 (N_816,In_350,In_562);
nor U817 (N_817,In_143,In_263);
nor U818 (N_818,In_920,In_672);
and U819 (N_819,In_39,In_989);
nand U820 (N_820,In_50,In_961);
and U821 (N_821,In_282,In_572);
nor U822 (N_822,In_535,In_24);
or U823 (N_823,In_129,In_608);
and U824 (N_824,In_872,In_956);
and U825 (N_825,In_347,In_707);
and U826 (N_826,In_586,In_810);
nand U827 (N_827,In_41,In_154);
or U828 (N_828,In_107,In_22);
or U829 (N_829,In_174,In_183);
nor U830 (N_830,In_523,In_973);
or U831 (N_831,In_760,In_261);
nand U832 (N_832,In_365,In_548);
nor U833 (N_833,In_581,In_999);
nand U834 (N_834,In_179,In_633);
nand U835 (N_835,In_76,In_293);
nor U836 (N_836,In_517,In_801);
nor U837 (N_837,In_510,In_348);
nand U838 (N_838,In_870,In_822);
nand U839 (N_839,In_500,In_203);
nand U840 (N_840,In_694,In_772);
and U841 (N_841,In_612,In_264);
nand U842 (N_842,In_122,In_625);
nor U843 (N_843,In_559,In_265);
and U844 (N_844,In_66,In_700);
nand U845 (N_845,In_836,In_545);
nor U846 (N_846,In_370,In_955);
nor U847 (N_847,In_911,In_863);
nor U848 (N_848,In_615,In_748);
or U849 (N_849,In_321,In_199);
xnor U850 (N_850,In_91,In_612);
nor U851 (N_851,In_269,In_373);
nand U852 (N_852,In_864,In_50);
and U853 (N_853,In_489,In_1);
or U854 (N_854,In_805,In_66);
or U855 (N_855,In_971,In_659);
or U856 (N_856,In_817,In_595);
and U857 (N_857,In_504,In_963);
nand U858 (N_858,In_917,In_273);
nand U859 (N_859,In_771,In_983);
nor U860 (N_860,In_277,In_302);
nor U861 (N_861,In_795,In_481);
nor U862 (N_862,In_619,In_213);
nand U863 (N_863,In_6,In_849);
nand U864 (N_864,In_785,In_922);
or U865 (N_865,In_641,In_392);
and U866 (N_866,In_103,In_643);
and U867 (N_867,In_745,In_878);
and U868 (N_868,In_966,In_191);
nor U869 (N_869,In_247,In_406);
nor U870 (N_870,In_866,In_976);
or U871 (N_871,In_460,In_55);
or U872 (N_872,In_385,In_735);
nand U873 (N_873,In_429,In_879);
nand U874 (N_874,In_398,In_534);
or U875 (N_875,In_897,In_961);
nand U876 (N_876,In_819,In_539);
and U877 (N_877,In_110,In_891);
nand U878 (N_878,In_531,In_751);
or U879 (N_879,In_607,In_934);
nand U880 (N_880,In_620,In_860);
and U881 (N_881,In_161,In_139);
nand U882 (N_882,In_177,In_191);
or U883 (N_883,In_266,In_561);
and U884 (N_884,In_261,In_984);
and U885 (N_885,In_328,In_314);
nand U886 (N_886,In_476,In_609);
or U887 (N_887,In_184,In_611);
or U888 (N_888,In_655,In_213);
nand U889 (N_889,In_636,In_625);
and U890 (N_890,In_488,In_679);
nand U891 (N_891,In_823,In_192);
and U892 (N_892,In_80,In_0);
nand U893 (N_893,In_843,In_535);
nor U894 (N_894,In_700,In_472);
or U895 (N_895,In_703,In_83);
or U896 (N_896,In_706,In_307);
nand U897 (N_897,In_584,In_655);
nor U898 (N_898,In_878,In_414);
or U899 (N_899,In_96,In_953);
nor U900 (N_900,In_316,In_2);
and U901 (N_901,In_737,In_270);
nor U902 (N_902,In_505,In_678);
nand U903 (N_903,In_983,In_624);
or U904 (N_904,In_55,In_758);
nand U905 (N_905,In_849,In_263);
nand U906 (N_906,In_771,In_622);
nor U907 (N_907,In_982,In_979);
nor U908 (N_908,In_374,In_599);
and U909 (N_909,In_689,In_923);
or U910 (N_910,In_129,In_858);
or U911 (N_911,In_688,In_896);
nand U912 (N_912,In_882,In_382);
nand U913 (N_913,In_940,In_293);
and U914 (N_914,In_566,In_953);
xnor U915 (N_915,In_66,In_394);
and U916 (N_916,In_306,In_663);
and U917 (N_917,In_927,In_973);
nand U918 (N_918,In_48,In_96);
nor U919 (N_919,In_362,In_778);
xor U920 (N_920,In_542,In_704);
and U921 (N_921,In_977,In_658);
or U922 (N_922,In_334,In_454);
and U923 (N_923,In_323,In_452);
and U924 (N_924,In_912,In_248);
and U925 (N_925,In_654,In_418);
nor U926 (N_926,In_165,In_590);
nand U927 (N_927,In_931,In_349);
or U928 (N_928,In_864,In_369);
nor U929 (N_929,In_928,In_910);
nor U930 (N_930,In_165,In_687);
nor U931 (N_931,In_580,In_358);
nor U932 (N_932,In_901,In_182);
nor U933 (N_933,In_837,In_232);
nor U934 (N_934,In_815,In_699);
and U935 (N_935,In_479,In_847);
or U936 (N_936,In_792,In_892);
xnor U937 (N_937,In_962,In_282);
nor U938 (N_938,In_377,In_112);
nor U939 (N_939,In_624,In_618);
nor U940 (N_940,In_427,In_98);
nand U941 (N_941,In_799,In_681);
nand U942 (N_942,In_607,In_286);
nand U943 (N_943,In_970,In_710);
nor U944 (N_944,In_855,In_222);
or U945 (N_945,In_776,In_944);
nor U946 (N_946,In_347,In_550);
or U947 (N_947,In_833,In_741);
and U948 (N_948,In_401,In_479);
and U949 (N_949,In_821,In_887);
and U950 (N_950,In_54,In_579);
nand U951 (N_951,In_986,In_708);
nand U952 (N_952,In_48,In_149);
nor U953 (N_953,In_215,In_997);
nor U954 (N_954,In_488,In_995);
or U955 (N_955,In_308,In_227);
nor U956 (N_956,In_980,In_351);
or U957 (N_957,In_226,In_656);
nor U958 (N_958,In_697,In_335);
nand U959 (N_959,In_763,In_623);
and U960 (N_960,In_82,In_766);
nor U961 (N_961,In_68,In_1);
and U962 (N_962,In_243,In_622);
nor U963 (N_963,In_832,In_257);
nor U964 (N_964,In_772,In_171);
and U965 (N_965,In_869,In_805);
and U966 (N_966,In_810,In_144);
or U967 (N_967,In_104,In_921);
or U968 (N_968,In_546,In_100);
nand U969 (N_969,In_91,In_189);
nand U970 (N_970,In_327,In_256);
nor U971 (N_971,In_618,In_981);
nand U972 (N_972,In_154,In_770);
nor U973 (N_973,In_718,In_705);
or U974 (N_974,In_284,In_628);
nand U975 (N_975,In_991,In_33);
nor U976 (N_976,In_413,In_109);
and U977 (N_977,In_532,In_780);
and U978 (N_978,In_967,In_958);
and U979 (N_979,In_926,In_790);
xor U980 (N_980,In_485,In_767);
or U981 (N_981,In_572,In_461);
nand U982 (N_982,In_638,In_152);
and U983 (N_983,In_604,In_798);
nand U984 (N_984,In_679,In_59);
nor U985 (N_985,In_234,In_393);
nand U986 (N_986,In_793,In_966);
nor U987 (N_987,In_933,In_817);
or U988 (N_988,In_677,In_182);
nor U989 (N_989,In_764,In_27);
nand U990 (N_990,In_63,In_146);
nor U991 (N_991,In_174,In_474);
nand U992 (N_992,In_189,In_909);
nand U993 (N_993,In_592,In_316);
and U994 (N_994,In_374,In_115);
nor U995 (N_995,In_372,In_648);
and U996 (N_996,In_586,In_521);
nor U997 (N_997,In_726,In_383);
xnor U998 (N_998,In_790,In_592);
nor U999 (N_999,In_381,In_32);
nor U1000 (N_1000,In_294,In_17);
and U1001 (N_1001,In_582,In_546);
nand U1002 (N_1002,In_522,In_361);
or U1003 (N_1003,In_144,In_649);
nand U1004 (N_1004,In_599,In_975);
and U1005 (N_1005,In_482,In_176);
xor U1006 (N_1006,In_30,In_43);
or U1007 (N_1007,In_658,In_152);
nor U1008 (N_1008,In_499,In_42);
and U1009 (N_1009,In_194,In_399);
or U1010 (N_1010,In_687,In_523);
or U1011 (N_1011,In_282,In_906);
nor U1012 (N_1012,In_892,In_748);
and U1013 (N_1013,In_663,In_232);
and U1014 (N_1014,In_545,In_443);
nand U1015 (N_1015,In_50,In_887);
and U1016 (N_1016,In_930,In_232);
nor U1017 (N_1017,In_131,In_38);
nor U1018 (N_1018,In_941,In_78);
xor U1019 (N_1019,In_568,In_115);
nand U1020 (N_1020,In_292,In_183);
and U1021 (N_1021,In_746,In_789);
nor U1022 (N_1022,In_919,In_192);
or U1023 (N_1023,In_746,In_273);
or U1024 (N_1024,In_566,In_472);
or U1025 (N_1025,In_157,In_394);
nand U1026 (N_1026,In_887,In_248);
nand U1027 (N_1027,In_870,In_122);
nor U1028 (N_1028,In_120,In_648);
nand U1029 (N_1029,In_783,In_534);
or U1030 (N_1030,In_35,In_124);
and U1031 (N_1031,In_173,In_134);
or U1032 (N_1032,In_43,In_115);
nand U1033 (N_1033,In_767,In_395);
nor U1034 (N_1034,In_576,In_509);
or U1035 (N_1035,In_827,In_766);
nand U1036 (N_1036,In_865,In_234);
nor U1037 (N_1037,In_581,In_165);
nor U1038 (N_1038,In_345,In_835);
nand U1039 (N_1039,In_838,In_350);
or U1040 (N_1040,In_899,In_300);
nor U1041 (N_1041,In_294,In_84);
xor U1042 (N_1042,In_260,In_816);
or U1043 (N_1043,In_270,In_718);
or U1044 (N_1044,In_725,In_954);
or U1045 (N_1045,In_839,In_240);
and U1046 (N_1046,In_84,In_116);
or U1047 (N_1047,In_437,In_105);
nor U1048 (N_1048,In_623,In_505);
nand U1049 (N_1049,In_780,In_477);
and U1050 (N_1050,In_777,In_216);
or U1051 (N_1051,In_841,In_472);
nand U1052 (N_1052,In_767,In_50);
nor U1053 (N_1053,In_169,In_183);
nand U1054 (N_1054,In_133,In_296);
and U1055 (N_1055,In_392,In_579);
and U1056 (N_1056,In_990,In_441);
or U1057 (N_1057,In_931,In_306);
and U1058 (N_1058,In_955,In_745);
and U1059 (N_1059,In_170,In_240);
and U1060 (N_1060,In_147,In_37);
or U1061 (N_1061,In_212,In_600);
or U1062 (N_1062,In_973,In_372);
or U1063 (N_1063,In_44,In_415);
nor U1064 (N_1064,In_945,In_556);
nand U1065 (N_1065,In_347,In_170);
nand U1066 (N_1066,In_318,In_408);
nor U1067 (N_1067,In_226,In_682);
and U1068 (N_1068,In_705,In_25);
and U1069 (N_1069,In_22,In_196);
or U1070 (N_1070,In_321,In_247);
and U1071 (N_1071,In_271,In_518);
nor U1072 (N_1072,In_754,In_222);
nor U1073 (N_1073,In_484,In_533);
nand U1074 (N_1074,In_283,In_517);
or U1075 (N_1075,In_790,In_778);
and U1076 (N_1076,In_442,In_344);
nor U1077 (N_1077,In_348,In_354);
and U1078 (N_1078,In_917,In_611);
and U1079 (N_1079,In_673,In_804);
or U1080 (N_1080,In_61,In_473);
and U1081 (N_1081,In_150,In_552);
or U1082 (N_1082,In_617,In_634);
or U1083 (N_1083,In_127,In_238);
and U1084 (N_1084,In_874,In_610);
nand U1085 (N_1085,In_717,In_116);
nand U1086 (N_1086,In_411,In_921);
or U1087 (N_1087,In_468,In_704);
or U1088 (N_1088,In_138,In_516);
nor U1089 (N_1089,In_523,In_774);
xor U1090 (N_1090,In_475,In_432);
and U1091 (N_1091,In_247,In_244);
or U1092 (N_1092,In_411,In_569);
nor U1093 (N_1093,In_356,In_710);
or U1094 (N_1094,In_29,In_167);
nand U1095 (N_1095,In_168,In_66);
nor U1096 (N_1096,In_884,In_913);
xnor U1097 (N_1097,In_212,In_351);
nand U1098 (N_1098,In_500,In_10);
and U1099 (N_1099,In_11,In_697);
nand U1100 (N_1100,In_597,In_263);
nor U1101 (N_1101,In_978,In_554);
or U1102 (N_1102,In_820,In_595);
nor U1103 (N_1103,In_850,In_539);
nand U1104 (N_1104,In_927,In_65);
xnor U1105 (N_1105,In_708,In_70);
or U1106 (N_1106,In_305,In_403);
nand U1107 (N_1107,In_681,In_915);
nand U1108 (N_1108,In_81,In_635);
and U1109 (N_1109,In_915,In_548);
or U1110 (N_1110,In_752,In_358);
and U1111 (N_1111,In_983,In_593);
nor U1112 (N_1112,In_149,In_173);
and U1113 (N_1113,In_209,In_486);
or U1114 (N_1114,In_878,In_89);
xor U1115 (N_1115,In_68,In_705);
nor U1116 (N_1116,In_370,In_252);
and U1117 (N_1117,In_332,In_334);
nand U1118 (N_1118,In_716,In_968);
or U1119 (N_1119,In_348,In_903);
and U1120 (N_1120,In_590,In_505);
nand U1121 (N_1121,In_487,In_493);
nand U1122 (N_1122,In_514,In_477);
or U1123 (N_1123,In_857,In_318);
or U1124 (N_1124,In_9,In_97);
and U1125 (N_1125,In_311,In_724);
or U1126 (N_1126,In_493,In_218);
nor U1127 (N_1127,In_934,In_551);
or U1128 (N_1128,In_214,In_988);
or U1129 (N_1129,In_65,In_985);
or U1130 (N_1130,In_523,In_189);
xnor U1131 (N_1131,In_424,In_343);
nand U1132 (N_1132,In_57,In_480);
nand U1133 (N_1133,In_950,In_326);
xor U1134 (N_1134,In_187,In_923);
or U1135 (N_1135,In_791,In_176);
nor U1136 (N_1136,In_723,In_820);
nand U1137 (N_1137,In_647,In_697);
or U1138 (N_1138,In_555,In_860);
and U1139 (N_1139,In_708,In_948);
nor U1140 (N_1140,In_981,In_524);
nor U1141 (N_1141,In_794,In_340);
nand U1142 (N_1142,In_927,In_320);
nor U1143 (N_1143,In_315,In_985);
nand U1144 (N_1144,In_174,In_981);
nand U1145 (N_1145,In_483,In_699);
or U1146 (N_1146,In_789,In_361);
nor U1147 (N_1147,In_666,In_679);
nand U1148 (N_1148,In_182,In_144);
and U1149 (N_1149,In_846,In_935);
or U1150 (N_1150,In_486,In_138);
or U1151 (N_1151,In_374,In_379);
and U1152 (N_1152,In_93,In_932);
or U1153 (N_1153,In_855,In_114);
nor U1154 (N_1154,In_25,In_103);
nand U1155 (N_1155,In_875,In_24);
or U1156 (N_1156,In_55,In_691);
nand U1157 (N_1157,In_192,In_752);
nor U1158 (N_1158,In_393,In_413);
or U1159 (N_1159,In_561,In_202);
nor U1160 (N_1160,In_292,In_261);
and U1161 (N_1161,In_782,In_924);
or U1162 (N_1162,In_780,In_462);
nand U1163 (N_1163,In_907,In_735);
or U1164 (N_1164,In_325,In_595);
nand U1165 (N_1165,In_806,In_896);
and U1166 (N_1166,In_644,In_580);
nand U1167 (N_1167,In_195,In_753);
nand U1168 (N_1168,In_983,In_267);
nor U1169 (N_1169,In_952,In_946);
or U1170 (N_1170,In_33,In_74);
nor U1171 (N_1171,In_185,In_371);
and U1172 (N_1172,In_757,In_66);
and U1173 (N_1173,In_566,In_0);
or U1174 (N_1174,In_121,In_799);
nand U1175 (N_1175,In_488,In_765);
and U1176 (N_1176,In_497,In_770);
and U1177 (N_1177,In_150,In_66);
nor U1178 (N_1178,In_61,In_888);
nand U1179 (N_1179,In_243,In_245);
nor U1180 (N_1180,In_450,In_613);
xor U1181 (N_1181,In_853,In_727);
nand U1182 (N_1182,In_833,In_197);
nor U1183 (N_1183,In_644,In_154);
or U1184 (N_1184,In_154,In_207);
nand U1185 (N_1185,In_209,In_40);
or U1186 (N_1186,In_639,In_826);
nor U1187 (N_1187,In_970,In_933);
and U1188 (N_1188,In_57,In_399);
nor U1189 (N_1189,In_236,In_788);
and U1190 (N_1190,In_116,In_486);
nand U1191 (N_1191,In_311,In_208);
nand U1192 (N_1192,In_769,In_641);
and U1193 (N_1193,In_449,In_454);
nor U1194 (N_1194,In_359,In_980);
or U1195 (N_1195,In_477,In_750);
and U1196 (N_1196,In_912,In_971);
and U1197 (N_1197,In_494,In_148);
nor U1198 (N_1198,In_549,In_376);
or U1199 (N_1199,In_228,In_682);
and U1200 (N_1200,In_32,In_518);
and U1201 (N_1201,In_161,In_695);
nor U1202 (N_1202,In_93,In_682);
or U1203 (N_1203,In_532,In_585);
or U1204 (N_1204,In_358,In_74);
or U1205 (N_1205,In_851,In_143);
and U1206 (N_1206,In_58,In_513);
nand U1207 (N_1207,In_44,In_550);
and U1208 (N_1208,In_458,In_430);
and U1209 (N_1209,In_278,In_463);
and U1210 (N_1210,In_407,In_938);
nor U1211 (N_1211,In_989,In_87);
or U1212 (N_1212,In_622,In_743);
nor U1213 (N_1213,In_505,In_202);
or U1214 (N_1214,In_7,In_687);
and U1215 (N_1215,In_529,In_172);
xor U1216 (N_1216,In_357,In_61);
nor U1217 (N_1217,In_582,In_21);
nor U1218 (N_1218,In_221,In_199);
and U1219 (N_1219,In_477,In_456);
or U1220 (N_1220,In_463,In_562);
nand U1221 (N_1221,In_352,In_336);
and U1222 (N_1222,In_443,In_695);
nand U1223 (N_1223,In_211,In_496);
nand U1224 (N_1224,In_646,In_757);
nand U1225 (N_1225,In_646,In_880);
and U1226 (N_1226,In_57,In_442);
and U1227 (N_1227,In_776,In_231);
and U1228 (N_1228,In_928,In_153);
or U1229 (N_1229,In_130,In_36);
nand U1230 (N_1230,In_850,In_507);
and U1231 (N_1231,In_303,In_119);
nor U1232 (N_1232,In_130,In_621);
or U1233 (N_1233,In_792,In_205);
nand U1234 (N_1234,In_762,In_211);
nor U1235 (N_1235,In_918,In_869);
xor U1236 (N_1236,In_400,In_299);
nand U1237 (N_1237,In_101,In_922);
and U1238 (N_1238,In_596,In_587);
nor U1239 (N_1239,In_374,In_159);
or U1240 (N_1240,In_561,In_148);
or U1241 (N_1241,In_320,In_356);
nand U1242 (N_1242,In_345,In_301);
nor U1243 (N_1243,In_220,In_842);
and U1244 (N_1244,In_796,In_749);
or U1245 (N_1245,In_737,In_802);
nor U1246 (N_1246,In_241,In_791);
and U1247 (N_1247,In_42,In_636);
or U1248 (N_1248,In_826,In_830);
nor U1249 (N_1249,In_488,In_996);
nor U1250 (N_1250,In_288,In_235);
and U1251 (N_1251,In_757,In_697);
or U1252 (N_1252,In_761,In_340);
nand U1253 (N_1253,In_709,In_432);
or U1254 (N_1254,In_707,In_988);
or U1255 (N_1255,In_937,In_260);
nand U1256 (N_1256,In_698,In_391);
nand U1257 (N_1257,In_664,In_543);
nor U1258 (N_1258,In_998,In_188);
nand U1259 (N_1259,In_294,In_609);
nor U1260 (N_1260,In_185,In_950);
nor U1261 (N_1261,In_814,In_737);
and U1262 (N_1262,In_175,In_713);
or U1263 (N_1263,In_718,In_143);
nand U1264 (N_1264,In_378,In_221);
nand U1265 (N_1265,In_902,In_439);
and U1266 (N_1266,In_655,In_108);
nor U1267 (N_1267,In_200,In_915);
and U1268 (N_1268,In_699,In_882);
or U1269 (N_1269,In_635,In_512);
or U1270 (N_1270,In_333,In_264);
and U1271 (N_1271,In_640,In_350);
nand U1272 (N_1272,In_188,In_260);
and U1273 (N_1273,In_119,In_693);
or U1274 (N_1274,In_237,In_971);
nand U1275 (N_1275,In_652,In_840);
or U1276 (N_1276,In_623,In_866);
and U1277 (N_1277,In_232,In_301);
xnor U1278 (N_1278,In_124,In_906);
and U1279 (N_1279,In_68,In_928);
or U1280 (N_1280,In_510,In_943);
nor U1281 (N_1281,In_699,In_2);
or U1282 (N_1282,In_720,In_143);
and U1283 (N_1283,In_981,In_395);
nor U1284 (N_1284,In_217,In_111);
and U1285 (N_1285,In_793,In_681);
or U1286 (N_1286,In_240,In_699);
or U1287 (N_1287,In_532,In_345);
and U1288 (N_1288,In_445,In_42);
nor U1289 (N_1289,In_822,In_639);
nand U1290 (N_1290,In_393,In_37);
xnor U1291 (N_1291,In_618,In_523);
and U1292 (N_1292,In_177,In_599);
nor U1293 (N_1293,In_366,In_196);
nand U1294 (N_1294,In_77,In_421);
nand U1295 (N_1295,In_940,In_165);
and U1296 (N_1296,In_22,In_623);
and U1297 (N_1297,In_617,In_66);
and U1298 (N_1298,In_552,In_869);
and U1299 (N_1299,In_290,In_620);
nor U1300 (N_1300,In_627,In_593);
nor U1301 (N_1301,In_490,In_369);
or U1302 (N_1302,In_576,In_890);
nand U1303 (N_1303,In_705,In_702);
and U1304 (N_1304,In_388,In_595);
nor U1305 (N_1305,In_586,In_475);
nand U1306 (N_1306,In_953,In_63);
nor U1307 (N_1307,In_848,In_887);
or U1308 (N_1308,In_702,In_729);
nand U1309 (N_1309,In_388,In_883);
or U1310 (N_1310,In_127,In_983);
nand U1311 (N_1311,In_110,In_382);
and U1312 (N_1312,In_908,In_268);
or U1313 (N_1313,In_514,In_859);
nor U1314 (N_1314,In_804,In_395);
xor U1315 (N_1315,In_108,In_399);
and U1316 (N_1316,In_651,In_215);
or U1317 (N_1317,In_956,In_291);
or U1318 (N_1318,In_182,In_295);
nand U1319 (N_1319,In_136,In_69);
nor U1320 (N_1320,In_987,In_622);
or U1321 (N_1321,In_975,In_291);
nand U1322 (N_1322,In_602,In_931);
nand U1323 (N_1323,In_679,In_237);
nor U1324 (N_1324,In_858,In_472);
nor U1325 (N_1325,In_778,In_280);
or U1326 (N_1326,In_949,In_220);
nor U1327 (N_1327,In_21,In_604);
and U1328 (N_1328,In_609,In_226);
nand U1329 (N_1329,In_752,In_128);
nor U1330 (N_1330,In_394,In_311);
nor U1331 (N_1331,In_567,In_420);
nand U1332 (N_1332,In_28,In_82);
nand U1333 (N_1333,In_514,In_157);
nor U1334 (N_1334,In_637,In_115);
nand U1335 (N_1335,In_283,In_577);
and U1336 (N_1336,In_740,In_970);
and U1337 (N_1337,In_928,In_377);
and U1338 (N_1338,In_634,In_630);
and U1339 (N_1339,In_991,In_726);
nor U1340 (N_1340,In_240,In_656);
and U1341 (N_1341,In_687,In_255);
nand U1342 (N_1342,In_622,In_84);
nand U1343 (N_1343,In_433,In_204);
or U1344 (N_1344,In_292,In_687);
nand U1345 (N_1345,In_983,In_665);
or U1346 (N_1346,In_123,In_736);
and U1347 (N_1347,In_283,In_22);
nand U1348 (N_1348,In_65,In_978);
and U1349 (N_1349,In_476,In_188);
and U1350 (N_1350,In_160,In_284);
nand U1351 (N_1351,In_212,In_892);
nor U1352 (N_1352,In_245,In_422);
nor U1353 (N_1353,In_256,In_126);
nand U1354 (N_1354,In_826,In_831);
or U1355 (N_1355,In_870,In_81);
or U1356 (N_1356,In_381,In_33);
or U1357 (N_1357,In_992,In_718);
xnor U1358 (N_1358,In_349,In_284);
and U1359 (N_1359,In_242,In_107);
and U1360 (N_1360,In_929,In_115);
nor U1361 (N_1361,In_42,In_409);
nand U1362 (N_1362,In_719,In_312);
or U1363 (N_1363,In_451,In_422);
nand U1364 (N_1364,In_865,In_947);
nand U1365 (N_1365,In_133,In_236);
or U1366 (N_1366,In_985,In_494);
or U1367 (N_1367,In_30,In_859);
or U1368 (N_1368,In_339,In_645);
and U1369 (N_1369,In_575,In_382);
and U1370 (N_1370,In_90,In_602);
xnor U1371 (N_1371,In_637,In_496);
nor U1372 (N_1372,In_202,In_349);
nand U1373 (N_1373,In_789,In_545);
nor U1374 (N_1374,In_162,In_949);
nor U1375 (N_1375,In_584,In_149);
and U1376 (N_1376,In_671,In_339);
and U1377 (N_1377,In_169,In_511);
and U1378 (N_1378,In_133,In_84);
and U1379 (N_1379,In_501,In_582);
nor U1380 (N_1380,In_324,In_697);
nand U1381 (N_1381,In_710,In_916);
nand U1382 (N_1382,In_85,In_171);
nor U1383 (N_1383,In_881,In_62);
nand U1384 (N_1384,In_328,In_680);
nor U1385 (N_1385,In_714,In_84);
and U1386 (N_1386,In_722,In_507);
and U1387 (N_1387,In_583,In_9);
nand U1388 (N_1388,In_896,In_554);
or U1389 (N_1389,In_822,In_152);
or U1390 (N_1390,In_326,In_918);
or U1391 (N_1391,In_526,In_858);
and U1392 (N_1392,In_684,In_904);
nor U1393 (N_1393,In_798,In_813);
and U1394 (N_1394,In_287,In_470);
nand U1395 (N_1395,In_339,In_38);
and U1396 (N_1396,In_257,In_176);
or U1397 (N_1397,In_45,In_241);
and U1398 (N_1398,In_986,In_562);
and U1399 (N_1399,In_376,In_859);
nor U1400 (N_1400,In_723,In_553);
nand U1401 (N_1401,In_294,In_624);
or U1402 (N_1402,In_700,In_33);
or U1403 (N_1403,In_440,In_953);
nand U1404 (N_1404,In_996,In_584);
and U1405 (N_1405,In_101,In_161);
and U1406 (N_1406,In_763,In_991);
and U1407 (N_1407,In_535,In_978);
nor U1408 (N_1408,In_875,In_753);
or U1409 (N_1409,In_897,In_187);
and U1410 (N_1410,In_266,In_972);
nor U1411 (N_1411,In_126,In_736);
and U1412 (N_1412,In_84,In_624);
and U1413 (N_1413,In_841,In_957);
nand U1414 (N_1414,In_666,In_616);
nor U1415 (N_1415,In_274,In_770);
nand U1416 (N_1416,In_284,In_455);
or U1417 (N_1417,In_501,In_803);
or U1418 (N_1418,In_980,In_149);
or U1419 (N_1419,In_877,In_225);
nand U1420 (N_1420,In_443,In_349);
nor U1421 (N_1421,In_859,In_75);
and U1422 (N_1422,In_321,In_710);
and U1423 (N_1423,In_491,In_774);
nand U1424 (N_1424,In_457,In_964);
nor U1425 (N_1425,In_987,In_113);
nand U1426 (N_1426,In_801,In_146);
and U1427 (N_1427,In_772,In_532);
nand U1428 (N_1428,In_885,In_149);
nand U1429 (N_1429,In_137,In_252);
nor U1430 (N_1430,In_623,In_16);
or U1431 (N_1431,In_307,In_777);
nand U1432 (N_1432,In_912,In_322);
nor U1433 (N_1433,In_131,In_16);
or U1434 (N_1434,In_258,In_195);
nand U1435 (N_1435,In_716,In_603);
nor U1436 (N_1436,In_648,In_750);
or U1437 (N_1437,In_594,In_304);
nand U1438 (N_1438,In_970,In_642);
and U1439 (N_1439,In_760,In_7);
and U1440 (N_1440,In_838,In_517);
and U1441 (N_1441,In_370,In_467);
and U1442 (N_1442,In_598,In_968);
and U1443 (N_1443,In_895,In_673);
nand U1444 (N_1444,In_780,In_904);
nor U1445 (N_1445,In_119,In_780);
or U1446 (N_1446,In_234,In_73);
or U1447 (N_1447,In_417,In_310);
nor U1448 (N_1448,In_252,In_39);
and U1449 (N_1449,In_945,In_26);
nor U1450 (N_1450,In_827,In_832);
nand U1451 (N_1451,In_690,In_613);
nand U1452 (N_1452,In_931,In_934);
and U1453 (N_1453,In_484,In_400);
nor U1454 (N_1454,In_791,In_339);
nand U1455 (N_1455,In_431,In_199);
nand U1456 (N_1456,In_677,In_74);
nand U1457 (N_1457,In_136,In_13);
and U1458 (N_1458,In_508,In_502);
nand U1459 (N_1459,In_780,In_102);
nor U1460 (N_1460,In_42,In_977);
nand U1461 (N_1461,In_197,In_583);
or U1462 (N_1462,In_946,In_822);
nand U1463 (N_1463,In_932,In_554);
nand U1464 (N_1464,In_913,In_352);
nand U1465 (N_1465,In_107,In_525);
nor U1466 (N_1466,In_190,In_54);
and U1467 (N_1467,In_650,In_65);
nand U1468 (N_1468,In_387,In_143);
and U1469 (N_1469,In_275,In_250);
nand U1470 (N_1470,In_223,In_32);
or U1471 (N_1471,In_626,In_922);
and U1472 (N_1472,In_653,In_920);
or U1473 (N_1473,In_747,In_540);
nor U1474 (N_1474,In_333,In_501);
and U1475 (N_1475,In_247,In_825);
nand U1476 (N_1476,In_711,In_398);
and U1477 (N_1477,In_300,In_361);
or U1478 (N_1478,In_979,In_75);
nor U1479 (N_1479,In_418,In_633);
nand U1480 (N_1480,In_355,In_188);
or U1481 (N_1481,In_381,In_838);
nor U1482 (N_1482,In_721,In_186);
nand U1483 (N_1483,In_188,In_25);
nand U1484 (N_1484,In_883,In_43);
nor U1485 (N_1485,In_456,In_967);
nand U1486 (N_1486,In_303,In_608);
and U1487 (N_1487,In_872,In_61);
and U1488 (N_1488,In_935,In_463);
and U1489 (N_1489,In_46,In_332);
and U1490 (N_1490,In_588,In_1);
and U1491 (N_1491,In_198,In_30);
and U1492 (N_1492,In_605,In_648);
and U1493 (N_1493,In_372,In_432);
nor U1494 (N_1494,In_656,In_757);
nand U1495 (N_1495,In_158,In_401);
or U1496 (N_1496,In_25,In_629);
xor U1497 (N_1497,In_548,In_465);
and U1498 (N_1498,In_65,In_125);
nand U1499 (N_1499,In_874,In_158);
nand U1500 (N_1500,In_780,In_45);
nand U1501 (N_1501,In_127,In_694);
or U1502 (N_1502,In_199,In_716);
or U1503 (N_1503,In_85,In_151);
or U1504 (N_1504,In_103,In_666);
or U1505 (N_1505,In_857,In_176);
and U1506 (N_1506,In_898,In_663);
or U1507 (N_1507,In_119,In_39);
and U1508 (N_1508,In_228,In_951);
nand U1509 (N_1509,In_323,In_431);
xnor U1510 (N_1510,In_453,In_318);
nand U1511 (N_1511,In_799,In_610);
and U1512 (N_1512,In_95,In_674);
or U1513 (N_1513,In_955,In_544);
nand U1514 (N_1514,In_108,In_448);
or U1515 (N_1515,In_240,In_316);
nor U1516 (N_1516,In_301,In_290);
nand U1517 (N_1517,In_255,In_55);
nand U1518 (N_1518,In_569,In_905);
nor U1519 (N_1519,In_959,In_776);
nor U1520 (N_1520,In_56,In_604);
or U1521 (N_1521,In_794,In_815);
or U1522 (N_1522,In_171,In_215);
or U1523 (N_1523,In_662,In_412);
and U1524 (N_1524,In_336,In_188);
and U1525 (N_1525,In_849,In_125);
and U1526 (N_1526,In_160,In_738);
nor U1527 (N_1527,In_768,In_134);
nor U1528 (N_1528,In_789,In_715);
nand U1529 (N_1529,In_779,In_98);
and U1530 (N_1530,In_3,In_973);
nand U1531 (N_1531,In_20,In_702);
nand U1532 (N_1532,In_51,In_258);
or U1533 (N_1533,In_371,In_728);
and U1534 (N_1534,In_572,In_595);
nor U1535 (N_1535,In_867,In_212);
nor U1536 (N_1536,In_529,In_571);
and U1537 (N_1537,In_184,In_876);
or U1538 (N_1538,In_323,In_843);
and U1539 (N_1539,In_921,In_545);
nand U1540 (N_1540,In_338,In_641);
nand U1541 (N_1541,In_382,In_818);
or U1542 (N_1542,In_932,In_842);
and U1543 (N_1543,In_174,In_553);
and U1544 (N_1544,In_50,In_118);
or U1545 (N_1545,In_766,In_33);
or U1546 (N_1546,In_970,In_486);
and U1547 (N_1547,In_277,In_811);
or U1548 (N_1548,In_326,In_952);
nand U1549 (N_1549,In_938,In_405);
and U1550 (N_1550,In_127,In_19);
nand U1551 (N_1551,In_468,In_519);
xnor U1552 (N_1552,In_46,In_340);
nand U1553 (N_1553,In_944,In_257);
and U1554 (N_1554,In_514,In_725);
and U1555 (N_1555,In_562,In_232);
nor U1556 (N_1556,In_425,In_525);
or U1557 (N_1557,In_46,In_140);
or U1558 (N_1558,In_392,In_803);
and U1559 (N_1559,In_529,In_419);
or U1560 (N_1560,In_784,In_883);
nand U1561 (N_1561,In_970,In_265);
nor U1562 (N_1562,In_945,In_139);
and U1563 (N_1563,In_762,In_866);
and U1564 (N_1564,In_65,In_114);
and U1565 (N_1565,In_445,In_261);
and U1566 (N_1566,In_93,In_194);
and U1567 (N_1567,In_54,In_533);
or U1568 (N_1568,In_688,In_185);
nor U1569 (N_1569,In_107,In_39);
nand U1570 (N_1570,In_395,In_450);
or U1571 (N_1571,In_742,In_551);
and U1572 (N_1572,In_595,In_946);
nand U1573 (N_1573,In_118,In_484);
nor U1574 (N_1574,In_604,In_40);
and U1575 (N_1575,In_38,In_181);
nand U1576 (N_1576,In_900,In_54);
nand U1577 (N_1577,In_654,In_645);
or U1578 (N_1578,In_343,In_174);
nand U1579 (N_1579,In_829,In_775);
nor U1580 (N_1580,In_569,In_608);
nand U1581 (N_1581,In_142,In_133);
nor U1582 (N_1582,In_775,In_349);
nor U1583 (N_1583,In_808,In_731);
nor U1584 (N_1584,In_236,In_819);
nand U1585 (N_1585,In_533,In_584);
xnor U1586 (N_1586,In_30,In_650);
nor U1587 (N_1587,In_446,In_38);
or U1588 (N_1588,In_192,In_629);
nor U1589 (N_1589,In_974,In_699);
nor U1590 (N_1590,In_286,In_545);
and U1591 (N_1591,In_857,In_825);
or U1592 (N_1592,In_932,In_537);
and U1593 (N_1593,In_554,In_19);
or U1594 (N_1594,In_846,In_713);
and U1595 (N_1595,In_403,In_808);
and U1596 (N_1596,In_258,In_765);
nor U1597 (N_1597,In_613,In_68);
and U1598 (N_1598,In_742,In_576);
nor U1599 (N_1599,In_234,In_61);
nor U1600 (N_1600,In_428,In_821);
nor U1601 (N_1601,In_659,In_564);
or U1602 (N_1602,In_846,In_949);
nor U1603 (N_1603,In_639,In_443);
nor U1604 (N_1604,In_861,In_533);
nand U1605 (N_1605,In_64,In_698);
or U1606 (N_1606,In_282,In_395);
and U1607 (N_1607,In_854,In_696);
and U1608 (N_1608,In_268,In_869);
xnor U1609 (N_1609,In_516,In_587);
nor U1610 (N_1610,In_243,In_69);
xnor U1611 (N_1611,In_114,In_361);
nor U1612 (N_1612,In_138,In_511);
and U1613 (N_1613,In_317,In_887);
or U1614 (N_1614,In_673,In_207);
or U1615 (N_1615,In_123,In_920);
nand U1616 (N_1616,In_395,In_811);
and U1617 (N_1617,In_633,In_78);
nor U1618 (N_1618,In_41,In_627);
nor U1619 (N_1619,In_454,In_699);
nand U1620 (N_1620,In_778,In_197);
nor U1621 (N_1621,In_328,In_919);
and U1622 (N_1622,In_368,In_427);
nor U1623 (N_1623,In_244,In_27);
and U1624 (N_1624,In_11,In_273);
or U1625 (N_1625,In_262,In_691);
nor U1626 (N_1626,In_379,In_448);
nor U1627 (N_1627,In_74,In_171);
and U1628 (N_1628,In_392,In_708);
and U1629 (N_1629,In_422,In_405);
nand U1630 (N_1630,In_981,In_568);
nand U1631 (N_1631,In_79,In_849);
nor U1632 (N_1632,In_71,In_978);
and U1633 (N_1633,In_922,In_636);
or U1634 (N_1634,In_113,In_526);
nand U1635 (N_1635,In_590,In_494);
nand U1636 (N_1636,In_667,In_584);
nor U1637 (N_1637,In_687,In_994);
and U1638 (N_1638,In_627,In_481);
and U1639 (N_1639,In_905,In_520);
and U1640 (N_1640,In_192,In_513);
nand U1641 (N_1641,In_825,In_653);
xor U1642 (N_1642,In_498,In_711);
and U1643 (N_1643,In_866,In_377);
or U1644 (N_1644,In_287,In_190);
nor U1645 (N_1645,In_565,In_392);
nor U1646 (N_1646,In_958,In_781);
or U1647 (N_1647,In_929,In_124);
nand U1648 (N_1648,In_824,In_915);
and U1649 (N_1649,In_303,In_590);
nand U1650 (N_1650,In_433,In_140);
or U1651 (N_1651,In_205,In_829);
nand U1652 (N_1652,In_696,In_450);
and U1653 (N_1653,In_996,In_283);
nand U1654 (N_1654,In_578,In_460);
nor U1655 (N_1655,In_703,In_973);
nor U1656 (N_1656,In_687,In_343);
nor U1657 (N_1657,In_665,In_447);
and U1658 (N_1658,In_975,In_197);
or U1659 (N_1659,In_323,In_804);
nor U1660 (N_1660,In_813,In_791);
nand U1661 (N_1661,In_570,In_636);
nor U1662 (N_1662,In_912,In_212);
nand U1663 (N_1663,In_616,In_544);
nand U1664 (N_1664,In_756,In_986);
nor U1665 (N_1665,In_428,In_444);
nor U1666 (N_1666,In_307,In_221);
nand U1667 (N_1667,In_402,In_75);
nor U1668 (N_1668,In_670,In_339);
nor U1669 (N_1669,In_813,In_636);
or U1670 (N_1670,In_269,In_24);
or U1671 (N_1671,In_894,In_823);
nand U1672 (N_1672,In_687,In_340);
nand U1673 (N_1673,In_29,In_259);
or U1674 (N_1674,In_108,In_571);
and U1675 (N_1675,In_47,In_101);
nor U1676 (N_1676,In_330,In_861);
or U1677 (N_1677,In_363,In_293);
nand U1678 (N_1678,In_525,In_653);
nand U1679 (N_1679,In_881,In_761);
nor U1680 (N_1680,In_563,In_1);
and U1681 (N_1681,In_740,In_842);
xor U1682 (N_1682,In_923,In_831);
or U1683 (N_1683,In_959,In_45);
and U1684 (N_1684,In_953,In_804);
or U1685 (N_1685,In_47,In_903);
nor U1686 (N_1686,In_480,In_790);
and U1687 (N_1687,In_72,In_388);
or U1688 (N_1688,In_558,In_955);
and U1689 (N_1689,In_708,In_37);
xor U1690 (N_1690,In_668,In_728);
or U1691 (N_1691,In_176,In_72);
nand U1692 (N_1692,In_827,In_338);
or U1693 (N_1693,In_146,In_582);
nand U1694 (N_1694,In_384,In_674);
or U1695 (N_1695,In_651,In_26);
or U1696 (N_1696,In_572,In_294);
nor U1697 (N_1697,In_200,In_447);
and U1698 (N_1698,In_30,In_825);
nor U1699 (N_1699,In_242,In_393);
or U1700 (N_1700,In_759,In_210);
and U1701 (N_1701,In_534,In_715);
or U1702 (N_1702,In_661,In_966);
nor U1703 (N_1703,In_798,In_528);
nand U1704 (N_1704,In_412,In_153);
nand U1705 (N_1705,In_204,In_682);
nor U1706 (N_1706,In_204,In_616);
nand U1707 (N_1707,In_781,In_864);
nor U1708 (N_1708,In_58,In_201);
or U1709 (N_1709,In_130,In_504);
and U1710 (N_1710,In_282,In_290);
nor U1711 (N_1711,In_598,In_380);
nand U1712 (N_1712,In_624,In_922);
and U1713 (N_1713,In_368,In_888);
nand U1714 (N_1714,In_717,In_971);
or U1715 (N_1715,In_883,In_251);
xor U1716 (N_1716,In_708,In_310);
or U1717 (N_1717,In_942,In_136);
nand U1718 (N_1718,In_632,In_226);
nand U1719 (N_1719,In_460,In_124);
nor U1720 (N_1720,In_223,In_845);
or U1721 (N_1721,In_121,In_276);
nand U1722 (N_1722,In_958,In_700);
and U1723 (N_1723,In_288,In_745);
and U1724 (N_1724,In_821,In_442);
nor U1725 (N_1725,In_969,In_222);
nand U1726 (N_1726,In_447,In_837);
nand U1727 (N_1727,In_604,In_375);
or U1728 (N_1728,In_570,In_871);
nor U1729 (N_1729,In_273,In_263);
nor U1730 (N_1730,In_196,In_379);
xnor U1731 (N_1731,In_39,In_919);
nor U1732 (N_1732,In_533,In_105);
or U1733 (N_1733,In_188,In_126);
nor U1734 (N_1734,In_786,In_901);
nor U1735 (N_1735,In_127,In_61);
nand U1736 (N_1736,In_480,In_726);
and U1737 (N_1737,In_663,In_933);
nand U1738 (N_1738,In_36,In_810);
nor U1739 (N_1739,In_606,In_729);
and U1740 (N_1740,In_9,In_153);
or U1741 (N_1741,In_353,In_217);
and U1742 (N_1742,In_205,In_481);
nor U1743 (N_1743,In_468,In_155);
nor U1744 (N_1744,In_121,In_212);
and U1745 (N_1745,In_109,In_340);
nand U1746 (N_1746,In_193,In_828);
nand U1747 (N_1747,In_502,In_896);
and U1748 (N_1748,In_75,In_44);
nor U1749 (N_1749,In_166,In_742);
and U1750 (N_1750,In_60,In_132);
nand U1751 (N_1751,In_219,In_289);
nand U1752 (N_1752,In_144,In_147);
and U1753 (N_1753,In_615,In_740);
or U1754 (N_1754,In_90,In_343);
or U1755 (N_1755,In_974,In_581);
nor U1756 (N_1756,In_690,In_819);
nor U1757 (N_1757,In_546,In_139);
or U1758 (N_1758,In_354,In_699);
nand U1759 (N_1759,In_267,In_821);
or U1760 (N_1760,In_199,In_428);
or U1761 (N_1761,In_144,In_541);
nand U1762 (N_1762,In_634,In_20);
or U1763 (N_1763,In_471,In_559);
or U1764 (N_1764,In_477,In_592);
nor U1765 (N_1765,In_718,In_682);
or U1766 (N_1766,In_943,In_44);
and U1767 (N_1767,In_164,In_950);
nand U1768 (N_1768,In_453,In_475);
nor U1769 (N_1769,In_357,In_331);
or U1770 (N_1770,In_71,In_189);
or U1771 (N_1771,In_705,In_906);
xor U1772 (N_1772,In_554,In_17);
and U1773 (N_1773,In_617,In_656);
nor U1774 (N_1774,In_89,In_988);
or U1775 (N_1775,In_725,In_234);
and U1776 (N_1776,In_164,In_528);
xnor U1777 (N_1777,In_139,In_800);
nand U1778 (N_1778,In_137,In_290);
nand U1779 (N_1779,In_550,In_814);
nor U1780 (N_1780,In_722,In_844);
or U1781 (N_1781,In_242,In_282);
or U1782 (N_1782,In_49,In_949);
or U1783 (N_1783,In_50,In_993);
and U1784 (N_1784,In_13,In_637);
or U1785 (N_1785,In_473,In_371);
nand U1786 (N_1786,In_143,In_938);
or U1787 (N_1787,In_560,In_437);
and U1788 (N_1788,In_684,In_223);
or U1789 (N_1789,In_204,In_51);
and U1790 (N_1790,In_370,In_324);
nand U1791 (N_1791,In_394,In_353);
nand U1792 (N_1792,In_432,In_451);
or U1793 (N_1793,In_646,In_140);
xnor U1794 (N_1794,In_244,In_512);
nor U1795 (N_1795,In_31,In_393);
and U1796 (N_1796,In_687,In_31);
and U1797 (N_1797,In_984,In_563);
nor U1798 (N_1798,In_882,In_281);
nand U1799 (N_1799,In_216,In_711);
nand U1800 (N_1800,In_533,In_226);
and U1801 (N_1801,In_317,In_195);
nand U1802 (N_1802,In_932,In_37);
xnor U1803 (N_1803,In_197,In_429);
and U1804 (N_1804,In_437,In_656);
or U1805 (N_1805,In_877,In_625);
or U1806 (N_1806,In_616,In_484);
nor U1807 (N_1807,In_56,In_695);
or U1808 (N_1808,In_480,In_736);
or U1809 (N_1809,In_617,In_470);
or U1810 (N_1810,In_931,In_598);
or U1811 (N_1811,In_666,In_148);
and U1812 (N_1812,In_196,In_564);
nor U1813 (N_1813,In_577,In_825);
or U1814 (N_1814,In_527,In_356);
nand U1815 (N_1815,In_946,In_645);
nand U1816 (N_1816,In_149,In_291);
or U1817 (N_1817,In_589,In_177);
nor U1818 (N_1818,In_142,In_223);
nand U1819 (N_1819,In_25,In_122);
nor U1820 (N_1820,In_598,In_619);
nor U1821 (N_1821,In_19,In_701);
nor U1822 (N_1822,In_293,In_15);
and U1823 (N_1823,In_659,In_37);
nor U1824 (N_1824,In_604,In_439);
or U1825 (N_1825,In_55,In_844);
and U1826 (N_1826,In_577,In_962);
and U1827 (N_1827,In_501,In_893);
nor U1828 (N_1828,In_772,In_917);
nor U1829 (N_1829,In_508,In_527);
nor U1830 (N_1830,In_136,In_803);
and U1831 (N_1831,In_874,In_766);
and U1832 (N_1832,In_832,In_947);
or U1833 (N_1833,In_444,In_305);
nand U1834 (N_1834,In_822,In_990);
nand U1835 (N_1835,In_542,In_625);
and U1836 (N_1836,In_519,In_592);
or U1837 (N_1837,In_52,In_700);
or U1838 (N_1838,In_710,In_84);
nor U1839 (N_1839,In_182,In_805);
nand U1840 (N_1840,In_985,In_690);
nand U1841 (N_1841,In_987,In_379);
or U1842 (N_1842,In_807,In_441);
and U1843 (N_1843,In_92,In_559);
and U1844 (N_1844,In_666,In_485);
nor U1845 (N_1845,In_455,In_155);
or U1846 (N_1846,In_384,In_3);
or U1847 (N_1847,In_87,In_559);
nand U1848 (N_1848,In_561,In_486);
nor U1849 (N_1849,In_875,In_732);
and U1850 (N_1850,In_935,In_450);
nor U1851 (N_1851,In_307,In_416);
or U1852 (N_1852,In_116,In_300);
nand U1853 (N_1853,In_469,In_993);
nor U1854 (N_1854,In_338,In_219);
nand U1855 (N_1855,In_404,In_80);
or U1856 (N_1856,In_217,In_503);
and U1857 (N_1857,In_889,In_382);
and U1858 (N_1858,In_176,In_610);
nand U1859 (N_1859,In_594,In_236);
and U1860 (N_1860,In_468,In_795);
nand U1861 (N_1861,In_486,In_316);
nor U1862 (N_1862,In_282,In_389);
or U1863 (N_1863,In_497,In_548);
or U1864 (N_1864,In_178,In_758);
and U1865 (N_1865,In_335,In_669);
and U1866 (N_1866,In_356,In_408);
xnor U1867 (N_1867,In_385,In_823);
nand U1868 (N_1868,In_564,In_278);
nor U1869 (N_1869,In_472,In_639);
or U1870 (N_1870,In_763,In_145);
or U1871 (N_1871,In_977,In_301);
or U1872 (N_1872,In_647,In_862);
nor U1873 (N_1873,In_902,In_498);
xor U1874 (N_1874,In_138,In_788);
or U1875 (N_1875,In_929,In_825);
and U1876 (N_1876,In_503,In_70);
nor U1877 (N_1877,In_932,In_638);
and U1878 (N_1878,In_319,In_758);
nand U1879 (N_1879,In_203,In_858);
and U1880 (N_1880,In_456,In_944);
xor U1881 (N_1881,In_505,In_217);
or U1882 (N_1882,In_736,In_727);
and U1883 (N_1883,In_80,In_712);
nor U1884 (N_1884,In_384,In_503);
nor U1885 (N_1885,In_261,In_648);
nand U1886 (N_1886,In_886,In_875);
and U1887 (N_1887,In_390,In_199);
or U1888 (N_1888,In_553,In_111);
nand U1889 (N_1889,In_580,In_376);
nand U1890 (N_1890,In_683,In_185);
nand U1891 (N_1891,In_846,In_217);
or U1892 (N_1892,In_330,In_184);
nand U1893 (N_1893,In_923,In_310);
nand U1894 (N_1894,In_668,In_474);
nand U1895 (N_1895,In_104,In_25);
and U1896 (N_1896,In_121,In_837);
and U1897 (N_1897,In_410,In_278);
or U1898 (N_1898,In_481,In_835);
nor U1899 (N_1899,In_471,In_25);
or U1900 (N_1900,In_456,In_261);
and U1901 (N_1901,In_499,In_549);
and U1902 (N_1902,In_91,In_111);
and U1903 (N_1903,In_776,In_267);
nand U1904 (N_1904,In_952,In_816);
nand U1905 (N_1905,In_552,In_824);
or U1906 (N_1906,In_242,In_214);
or U1907 (N_1907,In_444,In_231);
nand U1908 (N_1908,In_796,In_418);
nand U1909 (N_1909,In_285,In_944);
or U1910 (N_1910,In_388,In_726);
xor U1911 (N_1911,In_325,In_623);
xnor U1912 (N_1912,In_16,In_432);
and U1913 (N_1913,In_513,In_776);
nand U1914 (N_1914,In_653,In_999);
nor U1915 (N_1915,In_817,In_123);
and U1916 (N_1916,In_133,In_660);
and U1917 (N_1917,In_614,In_642);
nor U1918 (N_1918,In_670,In_963);
nor U1919 (N_1919,In_947,In_847);
nand U1920 (N_1920,In_620,In_150);
and U1921 (N_1921,In_11,In_790);
nor U1922 (N_1922,In_68,In_824);
nor U1923 (N_1923,In_185,In_670);
nand U1924 (N_1924,In_170,In_108);
nor U1925 (N_1925,In_821,In_382);
or U1926 (N_1926,In_137,In_268);
or U1927 (N_1927,In_519,In_825);
xnor U1928 (N_1928,In_968,In_582);
nand U1929 (N_1929,In_250,In_542);
xor U1930 (N_1930,In_862,In_933);
and U1931 (N_1931,In_720,In_318);
nor U1932 (N_1932,In_937,In_41);
and U1933 (N_1933,In_955,In_35);
nand U1934 (N_1934,In_551,In_127);
nor U1935 (N_1935,In_698,In_904);
nand U1936 (N_1936,In_847,In_184);
or U1937 (N_1937,In_667,In_884);
nand U1938 (N_1938,In_660,In_73);
nor U1939 (N_1939,In_883,In_371);
nand U1940 (N_1940,In_607,In_686);
or U1941 (N_1941,In_802,In_178);
nor U1942 (N_1942,In_4,In_394);
or U1943 (N_1943,In_854,In_986);
and U1944 (N_1944,In_700,In_748);
and U1945 (N_1945,In_231,In_281);
and U1946 (N_1946,In_411,In_304);
or U1947 (N_1947,In_393,In_238);
nand U1948 (N_1948,In_57,In_424);
or U1949 (N_1949,In_219,In_222);
or U1950 (N_1950,In_513,In_991);
nor U1951 (N_1951,In_156,In_860);
nor U1952 (N_1952,In_919,In_805);
nor U1953 (N_1953,In_543,In_5);
or U1954 (N_1954,In_570,In_343);
or U1955 (N_1955,In_882,In_118);
nor U1956 (N_1956,In_592,In_728);
and U1957 (N_1957,In_786,In_450);
nand U1958 (N_1958,In_580,In_796);
nor U1959 (N_1959,In_640,In_285);
nand U1960 (N_1960,In_678,In_37);
or U1961 (N_1961,In_501,In_119);
nor U1962 (N_1962,In_240,In_65);
nand U1963 (N_1963,In_508,In_498);
or U1964 (N_1964,In_887,In_652);
nor U1965 (N_1965,In_142,In_793);
and U1966 (N_1966,In_658,In_194);
or U1967 (N_1967,In_84,In_706);
or U1968 (N_1968,In_983,In_100);
and U1969 (N_1969,In_146,In_5);
or U1970 (N_1970,In_605,In_620);
and U1971 (N_1971,In_620,In_857);
nand U1972 (N_1972,In_699,In_290);
and U1973 (N_1973,In_606,In_252);
nor U1974 (N_1974,In_111,In_289);
nand U1975 (N_1975,In_733,In_152);
or U1976 (N_1976,In_804,In_44);
and U1977 (N_1977,In_91,In_286);
nand U1978 (N_1978,In_910,In_371);
nor U1979 (N_1979,In_353,In_805);
or U1980 (N_1980,In_553,In_600);
nor U1981 (N_1981,In_182,In_313);
nand U1982 (N_1982,In_423,In_128);
nor U1983 (N_1983,In_896,In_900);
nor U1984 (N_1984,In_622,In_432);
and U1985 (N_1985,In_96,In_35);
nand U1986 (N_1986,In_241,In_55);
nand U1987 (N_1987,In_616,In_873);
nor U1988 (N_1988,In_779,In_308);
or U1989 (N_1989,In_20,In_509);
and U1990 (N_1990,In_577,In_345);
and U1991 (N_1991,In_966,In_1);
or U1992 (N_1992,In_732,In_587);
nor U1993 (N_1993,In_207,In_53);
or U1994 (N_1994,In_366,In_881);
nand U1995 (N_1995,In_565,In_393);
and U1996 (N_1996,In_336,In_17);
nand U1997 (N_1997,In_412,In_134);
and U1998 (N_1998,In_798,In_738);
nor U1999 (N_1999,In_562,In_783);
nand U2000 (N_2000,In_195,In_564);
nand U2001 (N_2001,In_584,In_147);
nand U2002 (N_2002,In_678,In_274);
nor U2003 (N_2003,In_60,In_55);
or U2004 (N_2004,In_553,In_583);
nand U2005 (N_2005,In_69,In_610);
nor U2006 (N_2006,In_316,In_173);
nand U2007 (N_2007,In_882,In_746);
or U2008 (N_2008,In_384,In_742);
or U2009 (N_2009,In_624,In_740);
nor U2010 (N_2010,In_359,In_262);
or U2011 (N_2011,In_346,In_268);
nor U2012 (N_2012,In_681,In_545);
nor U2013 (N_2013,In_783,In_185);
nand U2014 (N_2014,In_962,In_433);
and U2015 (N_2015,In_541,In_488);
nand U2016 (N_2016,In_832,In_199);
or U2017 (N_2017,In_384,In_253);
and U2018 (N_2018,In_659,In_227);
nand U2019 (N_2019,In_31,In_126);
nor U2020 (N_2020,In_281,In_324);
or U2021 (N_2021,In_427,In_307);
and U2022 (N_2022,In_612,In_827);
nor U2023 (N_2023,In_591,In_161);
nor U2024 (N_2024,In_711,In_643);
and U2025 (N_2025,In_26,In_841);
nand U2026 (N_2026,In_402,In_565);
nor U2027 (N_2027,In_12,In_955);
nor U2028 (N_2028,In_617,In_972);
nand U2029 (N_2029,In_804,In_742);
nand U2030 (N_2030,In_725,In_656);
and U2031 (N_2031,In_214,In_187);
nand U2032 (N_2032,In_824,In_956);
nor U2033 (N_2033,In_403,In_927);
or U2034 (N_2034,In_484,In_169);
nand U2035 (N_2035,In_896,In_68);
nor U2036 (N_2036,In_773,In_195);
nand U2037 (N_2037,In_12,In_638);
nor U2038 (N_2038,In_170,In_793);
nand U2039 (N_2039,In_310,In_718);
or U2040 (N_2040,In_634,In_949);
or U2041 (N_2041,In_120,In_627);
nand U2042 (N_2042,In_513,In_896);
nor U2043 (N_2043,In_775,In_620);
or U2044 (N_2044,In_852,In_74);
nor U2045 (N_2045,In_64,In_838);
nor U2046 (N_2046,In_996,In_228);
or U2047 (N_2047,In_443,In_447);
nand U2048 (N_2048,In_533,In_95);
or U2049 (N_2049,In_334,In_783);
and U2050 (N_2050,In_987,In_339);
xor U2051 (N_2051,In_59,In_292);
nand U2052 (N_2052,In_392,In_709);
nor U2053 (N_2053,In_73,In_544);
and U2054 (N_2054,In_469,In_730);
nand U2055 (N_2055,In_408,In_399);
or U2056 (N_2056,In_961,In_86);
nand U2057 (N_2057,In_986,In_941);
or U2058 (N_2058,In_41,In_437);
or U2059 (N_2059,In_154,In_503);
xnor U2060 (N_2060,In_854,In_358);
and U2061 (N_2061,In_181,In_584);
and U2062 (N_2062,In_356,In_989);
or U2063 (N_2063,In_309,In_987);
or U2064 (N_2064,In_420,In_565);
or U2065 (N_2065,In_318,In_736);
xor U2066 (N_2066,In_597,In_630);
xnor U2067 (N_2067,In_630,In_479);
nand U2068 (N_2068,In_913,In_987);
nand U2069 (N_2069,In_731,In_598);
nand U2070 (N_2070,In_437,In_153);
nor U2071 (N_2071,In_920,In_429);
or U2072 (N_2072,In_700,In_931);
or U2073 (N_2073,In_960,In_242);
or U2074 (N_2074,In_759,In_653);
and U2075 (N_2075,In_155,In_454);
nand U2076 (N_2076,In_649,In_435);
nor U2077 (N_2077,In_784,In_738);
or U2078 (N_2078,In_789,In_949);
or U2079 (N_2079,In_109,In_138);
nor U2080 (N_2080,In_509,In_304);
and U2081 (N_2081,In_986,In_58);
nand U2082 (N_2082,In_997,In_779);
or U2083 (N_2083,In_44,In_681);
or U2084 (N_2084,In_393,In_797);
nor U2085 (N_2085,In_502,In_242);
nor U2086 (N_2086,In_468,In_824);
and U2087 (N_2087,In_915,In_244);
or U2088 (N_2088,In_598,In_458);
or U2089 (N_2089,In_271,In_783);
and U2090 (N_2090,In_758,In_878);
and U2091 (N_2091,In_826,In_967);
nor U2092 (N_2092,In_98,In_715);
or U2093 (N_2093,In_799,In_88);
or U2094 (N_2094,In_207,In_523);
nor U2095 (N_2095,In_436,In_541);
or U2096 (N_2096,In_670,In_580);
and U2097 (N_2097,In_977,In_787);
or U2098 (N_2098,In_141,In_654);
nor U2099 (N_2099,In_179,In_311);
xor U2100 (N_2100,In_744,In_872);
or U2101 (N_2101,In_103,In_141);
xnor U2102 (N_2102,In_246,In_945);
nand U2103 (N_2103,In_694,In_45);
and U2104 (N_2104,In_0,In_737);
nor U2105 (N_2105,In_757,In_159);
nor U2106 (N_2106,In_3,In_778);
or U2107 (N_2107,In_886,In_600);
nand U2108 (N_2108,In_709,In_809);
nand U2109 (N_2109,In_499,In_656);
and U2110 (N_2110,In_526,In_759);
and U2111 (N_2111,In_546,In_269);
or U2112 (N_2112,In_45,In_97);
nor U2113 (N_2113,In_581,In_882);
nor U2114 (N_2114,In_181,In_841);
or U2115 (N_2115,In_871,In_487);
nor U2116 (N_2116,In_384,In_657);
or U2117 (N_2117,In_972,In_357);
or U2118 (N_2118,In_109,In_324);
xnor U2119 (N_2119,In_874,In_123);
nor U2120 (N_2120,In_910,In_248);
xor U2121 (N_2121,In_557,In_486);
nor U2122 (N_2122,In_517,In_152);
or U2123 (N_2123,In_171,In_7);
nand U2124 (N_2124,In_624,In_929);
nand U2125 (N_2125,In_559,In_790);
nand U2126 (N_2126,In_520,In_699);
nand U2127 (N_2127,In_292,In_851);
nand U2128 (N_2128,In_464,In_766);
nor U2129 (N_2129,In_215,In_969);
nor U2130 (N_2130,In_241,In_979);
xor U2131 (N_2131,In_472,In_865);
and U2132 (N_2132,In_612,In_445);
nor U2133 (N_2133,In_107,In_384);
or U2134 (N_2134,In_41,In_33);
nand U2135 (N_2135,In_133,In_406);
nor U2136 (N_2136,In_875,In_151);
nand U2137 (N_2137,In_388,In_19);
or U2138 (N_2138,In_409,In_348);
or U2139 (N_2139,In_773,In_354);
nand U2140 (N_2140,In_461,In_360);
or U2141 (N_2141,In_607,In_539);
or U2142 (N_2142,In_623,In_314);
and U2143 (N_2143,In_789,In_446);
nor U2144 (N_2144,In_411,In_968);
nand U2145 (N_2145,In_173,In_97);
or U2146 (N_2146,In_361,In_896);
nor U2147 (N_2147,In_193,In_178);
nor U2148 (N_2148,In_607,In_85);
or U2149 (N_2149,In_349,In_66);
and U2150 (N_2150,In_256,In_201);
nor U2151 (N_2151,In_763,In_731);
or U2152 (N_2152,In_721,In_914);
and U2153 (N_2153,In_685,In_728);
and U2154 (N_2154,In_400,In_705);
or U2155 (N_2155,In_290,In_13);
nand U2156 (N_2156,In_125,In_659);
and U2157 (N_2157,In_658,In_316);
and U2158 (N_2158,In_66,In_253);
nand U2159 (N_2159,In_446,In_34);
and U2160 (N_2160,In_211,In_416);
and U2161 (N_2161,In_262,In_503);
xor U2162 (N_2162,In_774,In_956);
or U2163 (N_2163,In_592,In_614);
and U2164 (N_2164,In_520,In_616);
or U2165 (N_2165,In_862,In_217);
nor U2166 (N_2166,In_486,In_564);
and U2167 (N_2167,In_158,In_191);
nor U2168 (N_2168,In_896,In_129);
nor U2169 (N_2169,In_638,In_196);
nand U2170 (N_2170,In_497,In_14);
and U2171 (N_2171,In_356,In_19);
nor U2172 (N_2172,In_560,In_211);
nor U2173 (N_2173,In_57,In_140);
and U2174 (N_2174,In_985,In_857);
and U2175 (N_2175,In_825,In_491);
nand U2176 (N_2176,In_640,In_623);
or U2177 (N_2177,In_416,In_245);
nand U2178 (N_2178,In_450,In_250);
or U2179 (N_2179,In_269,In_561);
and U2180 (N_2180,In_220,In_502);
or U2181 (N_2181,In_264,In_393);
or U2182 (N_2182,In_14,In_913);
and U2183 (N_2183,In_27,In_955);
nand U2184 (N_2184,In_460,In_355);
nand U2185 (N_2185,In_909,In_675);
nor U2186 (N_2186,In_927,In_894);
nand U2187 (N_2187,In_98,In_958);
nand U2188 (N_2188,In_754,In_580);
and U2189 (N_2189,In_179,In_14);
and U2190 (N_2190,In_117,In_919);
nand U2191 (N_2191,In_288,In_249);
nand U2192 (N_2192,In_291,In_319);
nand U2193 (N_2193,In_435,In_643);
nor U2194 (N_2194,In_910,In_572);
nor U2195 (N_2195,In_436,In_770);
or U2196 (N_2196,In_316,In_427);
nor U2197 (N_2197,In_557,In_743);
nand U2198 (N_2198,In_143,In_673);
nor U2199 (N_2199,In_583,In_411);
nand U2200 (N_2200,In_361,In_213);
and U2201 (N_2201,In_542,In_738);
or U2202 (N_2202,In_484,In_691);
xor U2203 (N_2203,In_224,In_603);
nor U2204 (N_2204,In_123,In_748);
nor U2205 (N_2205,In_280,In_2);
and U2206 (N_2206,In_726,In_286);
nand U2207 (N_2207,In_86,In_707);
nor U2208 (N_2208,In_348,In_890);
nor U2209 (N_2209,In_33,In_897);
nand U2210 (N_2210,In_33,In_525);
or U2211 (N_2211,In_10,In_630);
and U2212 (N_2212,In_324,In_223);
and U2213 (N_2213,In_268,In_988);
nand U2214 (N_2214,In_521,In_811);
and U2215 (N_2215,In_970,In_378);
and U2216 (N_2216,In_989,In_7);
or U2217 (N_2217,In_960,In_744);
nand U2218 (N_2218,In_803,In_800);
nor U2219 (N_2219,In_802,In_924);
or U2220 (N_2220,In_589,In_264);
and U2221 (N_2221,In_914,In_263);
nor U2222 (N_2222,In_795,In_275);
or U2223 (N_2223,In_513,In_957);
or U2224 (N_2224,In_833,In_381);
nand U2225 (N_2225,In_932,In_913);
or U2226 (N_2226,In_340,In_310);
nor U2227 (N_2227,In_261,In_245);
or U2228 (N_2228,In_689,In_497);
nor U2229 (N_2229,In_727,In_115);
and U2230 (N_2230,In_812,In_68);
nor U2231 (N_2231,In_238,In_956);
nor U2232 (N_2232,In_865,In_619);
or U2233 (N_2233,In_136,In_526);
and U2234 (N_2234,In_114,In_567);
or U2235 (N_2235,In_683,In_934);
nand U2236 (N_2236,In_295,In_750);
and U2237 (N_2237,In_106,In_861);
nor U2238 (N_2238,In_814,In_717);
nand U2239 (N_2239,In_544,In_281);
or U2240 (N_2240,In_94,In_321);
nor U2241 (N_2241,In_548,In_736);
and U2242 (N_2242,In_611,In_16);
nor U2243 (N_2243,In_877,In_743);
and U2244 (N_2244,In_984,In_473);
and U2245 (N_2245,In_369,In_732);
or U2246 (N_2246,In_472,In_151);
nor U2247 (N_2247,In_988,In_374);
and U2248 (N_2248,In_971,In_181);
xor U2249 (N_2249,In_318,In_72);
nor U2250 (N_2250,In_730,In_520);
nor U2251 (N_2251,In_213,In_159);
or U2252 (N_2252,In_777,In_530);
nand U2253 (N_2253,In_696,In_335);
nor U2254 (N_2254,In_222,In_820);
xor U2255 (N_2255,In_10,In_368);
nor U2256 (N_2256,In_674,In_669);
nor U2257 (N_2257,In_88,In_552);
nand U2258 (N_2258,In_399,In_763);
and U2259 (N_2259,In_737,In_975);
nor U2260 (N_2260,In_120,In_106);
nor U2261 (N_2261,In_489,In_610);
nor U2262 (N_2262,In_435,In_390);
nor U2263 (N_2263,In_36,In_864);
xnor U2264 (N_2264,In_980,In_936);
xnor U2265 (N_2265,In_613,In_850);
nand U2266 (N_2266,In_440,In_187);
or U2267 (N_2267,In_70,In_769);
and U2268 (N_2268,In_783,In_470);
or U2269 (N_2269,In_322,In_936);
nand U2270 (N_2270,In_688,In_977);
or U2271 (N_2271,In_384,In_311);
or U2272 (N_2272,In_800,In_841);
or U2273 (N_2273,In_320,In_641);
nor U2274 (N_2274,In_707,In_225);
and U2275 (N_2275,In_34,In_41);
nor U2276 (N_2276,In_823,In_786);
nand U2277 (N_2277,In_231,In_68);
nand U2278 (N_2278,In_320,In_368);
nand U2279 (N_2279,In_897,In_805);
nand U2280 (N_2280,In_185,In_25);
or U2281 (N_2281,In_249,In_290);
nor U2282 (N_2282,In_771,In_921);
and U2283 (N_2283,In_843,In_629);
or U2284 (N_2284,In_803,In_813);
xnor U2285 (N_2285,In_401,In_482);
nor U2286 (N_2286,In_81,In_101);
and U2287 (N_2287,In_582,In_132);
or U2288 (N_2288,In_118,In_704);
nor U2289 (N_2289,In_312,In_481);
or U2290 (N_2290,In_78,In_305);
nand U2291 (N_2291,In_513,In_428);
nand U2292 (N_2292,In_709,In_770);
and U2293 (N_2293,In_143,In_351);
and U2294 (N_2294,In_282,In_640);
nand U2295 (N_2295,In_475,In_97);
nor U2296 (N_2296,In_825,In_912);
nand U2297 (N_2297,In_875,In_418);
or U2298 (N_2298,In_78,In_77);
and U2299 (N_2299,In_392,In_953);
nand U2300 (N_2300,In_599,In_52);
nand U2301 (N_2301,In_678,In_965);
xnor U2302 (N_2302,In_722,In_45);
and U2303 (N_2303,In_911,In_72);
and U2304 (N_2304,In_802,In_571);
xnor U2305 (N_2305,In_757,In_848);
nand U2306 (N_2306,In_832,In_87);
nor U2307 (N_2307,In_182,In_779);
nor U2308 (N_2308,In_197,In_228);
or U2309 (N_2309,In_915,In_871);
and U2310 (N_2310,In_79,In_615);
nor U2311 (N_2311,In_850,In_351);
and U2312 (N_2312,In_429,In_304);
or U2313 (N_2313,In_838,In_264);
nor U2314 (N_2314,In_817,In_405);
or U2315 (N_2315,In_699,In_613);
nand U2316 (N_2316,In_975,In_399);
or U2317 (N_2317,In_932,In_116);
and U2318 (N_2318,In_809,In_762);
and U2319 (N_2319,In_264,In_162);
or U2320 (N_2320,In_897,In_118);
nand U2321 (N_2321,In_959,In_755);
xor U2322 (N_2322,In_666,In_351);
nand U2323 (N_2323,In_541,In_413);
and U2324 (N_2324,In_228,In_847);
nand U2325 (N_2325,In_174,In_670);
or U2326 (N_2326,In_525,In_124);
nor U2327 (N_2327,In_898,In_225);
nand U2328 (N_2328,In_676,In_558);
nand U2329 (N_2329,In_345,In_704);
and U2330 (N_2330,In_588,In_728);
and U2331 (N_2331,In_782,In_386);
or U2332 (N_2332,In_834,In_152);
xnor U2333 (N_2333,In_866,In_897);
nor U2334 (N_2334,In_412,In_951);
nand U2335 (N_2335,In_4,In_738);
and U2336 (N_2336,In_910,In_22);
and U2337 (N_2337,In_147,In_295);
nand U2338 (N_2338,In_701,In_249);
nor U2339 (N_2339,In_952,In_489);
nor U2340 (N_2340,In_327,In_659);
or U2341 (N_2341,In_210,In_365);
nor U2342 (N_2342,In_539,In_368);
and U2343 (N_2343,In_11,In_406);
and U2344 (N_2344,In_788,In_658);
or U2345 (N_2345,In_708,In_328);
or U2346 (N_2346,In_140,In_385);
nor U2347 (N_2347,In_25,In_255);
or U2348 (N_2348,In_686,In_436);
and U2349 (N_2349,In_910,In_366);
and U2350 (N_2350,In_319,In_511);
and U2351 (N_2351,In_983,In_700);
and U2352 (N_2352,In_883,In_589);
or U2353 (N_2353,In_386,In_455);
and U2354 (N_2354,In_168,In_345);
xor U2355 (N_2355,In_391,In_546);
and U2356 (N_2356,In_329,In_486);
nand U2357 (N_2357,In_195,In_704);
or U2358 (N_2358,In_494,In_127);
and U2359 (N_2359,In_55,In_529);
nor U2360 (N_2360,In_864,In_870);
nor U2361 (N_2361,In_974,In_307);
and U2362 (N_2362,In_176,In_477);
xnor U2363 (N_2363,In_130,In_523);
nor U2364 (N_2364,In_79,In_184);
and U2365 (N_2365,In_787,In_796);
nand U2366 (N_2366,In_226,In_293);
or U2367 (N_2367,In_433,In_70);
or U2368 (N_2368,In_639,In_905);
nand U2369 (N_2369,In_135,In_376);
xnor U2370 (N_2370,In_803,In_45);
and U2371 (N_2371,In_349,In_536);
nand U2372 (N_2372,In_633,In_133);
nand U2373 (N_2373,In_349,In_989);
or U2374 (N_2374,In_261,In_585);
nor U2375 (N_2375,In_289,In_25);
and U2376 (N_2376,In_549,In_538);
or U2377 (N_2377,In_755,In_849);
nor U2378 (N_2378,In_272,In_722);
and U2379 (N_2379,In_174,In_756);
nor U2380 (N_2380,In_904,In_540);
nor U2381 (N_2381,In_90,In_677);
nor U2382 (N_2382,In_757,In_715);
or U2383 (N_2383,In_169,In_600);
nand U2384 (N_2384,In_566,In_810);
nor U2385 (N_2385,In_168,In_895);
nor U2386 (N_2386,In_517,In_94);
and U2387 (N_2387,In_553,In_782);
or U2388 (N_2388,In_603,In_812);
or U2389 (N_2389,In_607,In_458);
nor U2390 (N_2390,In_837,In_552);
and U2391 (N_2391,In_308,In_737);
xor U2392 (N_2392,In_89,In_978);
nor U2393 (N_2393,In_265,In_694);
nand U2394 (N_2394,In_484,In_406);
nor U2395 (N_2395,In_435,In_661);
nor U2396 (N_2396,In_562,In_272);
nand U2397 (N_2397,In_893,In_985);
and U2398 (N_2398,In_635,In_380);
nand U2399 (N_2399,In_588,In_140);
or U2400 (N_2400,In_622,In_75);
nor U2401 (N_2401,In_113,In_511);
or U2402 (N_2402,In_184,In_151);
nand U2403 (N_2403,In_182,In_38);
and U2404 (N_2404,In_515,In_227);
or U2405 (N_2405,In_154,In_481);
nor U2406 (N_2406,In_926,In_586);
xor U2407 (N_2407,In_681,In_933);
and U2408 (N_2408,In_487,In_497);
or U2409 (N_2409,In_81,In_803);
nand U2410 (N_2410,In_952,In_738);
and U2411 (N_2411,In_225,In_979);
or U2412 (N_2412,In_371,In_669);
nand U2413 (N_2413,In_912,In_870);
nor U2414 (N_2414,In_238,In_957);
and U2415 (N_2415,In_58,In_268);
and U2416 (N_2416,In_298,In_454);
and U2417 (N_2417,In_482,In_13);
or U2418 (N_2418,In_169,In_701);
xor U2419 (N_2419,In_994,In_232);
and U2420 (N_2420,In_649,In_120);
and U2421 (N_2421,In_35,In_123);
nor U2422 (N_2422,In_24,In_445);
nand U2423 (N_2423,In_9,In_507);
nand U2424 (N_2424,In_44,In_50);
and U2425 (N_2425,In_352,In_534);
nand U2426 (N_2426,In_724,In_166);
or U2427 (N_2427,In_262,In_325);
xnor U2428 (N_2428,In_757,In_434);
nor U2429 (N_2429,In_579,In_658);
nand U2430 (N_2430,In_497,In_484);
xor U2431 (N_2431,In_613,In_300);
and U2432 (N_2432,In_362,In_131);
and U2433 (N_2433,In_106,In_17);
nor U2434 (N_2434,In_991,In_668);
nor U2435 (N_2435,In_249,In_725);
or U2436 (N_2436,In_863,In_726);
and U2437 (N_2437,In_176,In_137);
nor U2438 (N_2438,In_747,In_513);
and U2439 (N_2439,In_999,In_808);
or U2440 (N_2440,In_375,In_158);
nand U2441 (N_2441,In_381,In_245);
nor U2442 (N_2442,In_510,In_979);
nand U2443 (N_2443,In_751,In_295);
and U2444 (N_2444,In_244,In_500);
or U2445 (N_2445,In_806,In_269);
nor U2446 (N_2446,In_421,In_762);
or U2447 (N_2447,In_176,In_9);
and U2448 (N_2448,In_480,In_601);
or U2449 (N_2449,In_986,In_463);
and U2450 (N_2450,In_646,In_154);
or U2451 (N_2451,In_947,In_598);
nor U2452 (N_2452,In_67,In_696);
and U2453 (N_2453,In_115,In_89);
nor U2454 (N_2454,In_758,In_296);
nand U2455 (N_2455,In_42,In_320);
nand U2456 (N_2456,In_310,In_179);
nor U2457 (N_2457,In_702,In_559);
nor U2458 (N_2458,In_222,In_586);
nor U2459 (N_2459,In_349,In_939);
nand U2460 (N_2460,In_525,In_559);
nand U2461 (N_2461,In_383,In_674);
and U2462 (N_2462,In_683,In_460);
nor U2463 (N_2463,In_58,In_719);
nand U2464 (N_2464,In_399,In_382);
nor U2465 (N_2465,In_246,In_45);
nand U2466 (N_2466,In_41,In_998);
nand U2467 (N_2467,In_362,In_84);
nand U2468 (N_2468,In_327,In_757);
or U2469 (N_2469,In_306,In_143);
nor U2470 (N_2470,In_0,In_802);
or U2471 (N_2471,In_86,In_555);
and U2472 (N_2472,In_505,In_695);
and U2473 (N_2473,In_468,In_9);
nand U2474 (N_2474,In_346,In_861);
nor U2475 (N_2475,In_199,In_776);
or U2476 (N_2476,In_198,In_666);
and U2477 (N_2477,In_606,In_163);
nand U2478 (N_2478,In_699,In_694);
nor U2479 (N_2479,In_967,In_9);
nand U2480 (N_2480,In_134,In_403);
or U2481 (N_2481,In_225,In_995);
nor U2482 (N_2482,In_29,In_277);
or U2483 (N_2483,In_805,In_293);
or U2484 (N_2484,In_743,In_915);
or U2485 (N_2485,In_99,In_531);
nor U2486 (N_2486,In_785,In_144);
xnor U2487 (N_2487,In_490,In_308);
and U2488 (N_2488,In_556,In_822);
nand U2489 (N_2489,In_361,In_748);
nor U2490 (N_2490,In_293,In_487);
or U2491 (N_2491,In_447,In_489);
and U2492 (N_2492,In_403,In_75);
nand U2493 (N_2493,In_455,In_176);
and U2494 (N_2494,In_967,In_173);
or U2495 (N_2495,In_710,In_616);
or U2496 (N_2496,In_972,In_239);
or U2497 (N_2497,In_729,In_566);
nand U2498 (N_2498,In_780,In_325);
nand U2499 (N_2499,In_944,In_878);
and U2500 (N_2500,N_1488,N_1020);
nand U2501 (N_2501,N_1862,N_589);
or U2502 (N_2502,N_521,N_1137);
and U2503 (N_2503,N_1028,N_2342);
nor U2504 (N_2504,N_1664,N_1156);
and U2505 (N_2505,N_36,N_164);
and U2506 (N_2506,N_2222,N_91);
and U2507 (N_2507,N_33,N_1160);
or U2508 (N_2508,N_2171,N_1201);
nand U2509 (N_2509,N_388,N_30);
nor U2510 (N_2510,N_6,N_1103);
nor U2511 (N_2511,N_1049,N_1421);
and U2512 (N_2512,N_1381,N_506);
nor U2513 (N_2513,N_1024,N_2264);
nor U2514 (N_2514,N_1632,N_1852);
nor U2515 (N_2515,N_480,N_2498);
nor U2516 (N_2516,N_1346,N_145);
nor U2517 (N_2517,N_2272,N_72);
or U2518 (N_2518,N_2210,N_1431);
nand U2519 (N_2519,N_1719,N_990);
nand U2520 (N_2520,N_482,N_1974);
nor U2521 (N_2521,N_1162,N_2008);
nor U2522 (N_2522,N_1276,N_377);
and U2523 (N_2523,N_774,N_281);
and U2524 (N_2524,N_2305,N_529);
and U2525 (N_2525,N_1202,N_2485);
or U2526 (N_2526,N_2098,N_295);
nand U2527 (N_2527,N_2476,N_971);
and U2528 (N_2528,N_23,N_106);
xnor U2529 (N_2529,N_889,N_980);
or U2530 (N_2530,N_1196,N_85);
and U2531 (N_2531,N_2135,N_501);
and U2532 (N_2532,N_934,N_1613);
nor U2533 (N_2533,N_770,N_1724);
nor U2534 (N_2534,N_717,N_423);
or U2535 (N_2535,N_196,N_290);
or U2536 (N_2536,N_51,N_386);
nand U2537 (N_2537,N_37,N_1341);
nand U2538 (N_2538,N_1979,N_2283);
nor U2539 (N_2539,N_286,N_2024);
and U2540 (N_2540,N_1859,N_741);
xnor U2541 (N_2541,N_874,N_2021);
or U2542 (N_2542,N_1966,N_2170);
or U2543 (N_2543,N_831,N_421);
and U2544 (N_2544,N_681,N_2348);
nand U2545 (N_2545,N_1797,N_1533);
or U2546 (N_2546,N_802,N_1016);
and U2547 (N_2547,N_1962,N_1861);
and U2548 (N_2548,N_2217,N_851);
and U2549 (N_2549,N_2052,N_287);
and U2550 (N_2550,N_1864,N_1151);
nor U2551 (N_2551,N_464,N_1122);
nor U2552 (N_2552,N_2417,N_279);
nand U2553 (N_2553,N_1807,N_2085);
nand U2554 (N_2554,N_928,N_588);
and U2555 (N_2555,N_974,N_2412);
nand U2556 (N_2556,N_923,N_98);
and U2557 (N_2557,N_1478,N_715);
and U2558 (N_2558,N_1805,N_1135);
nand U2559 (N_2559,N_1143,N_1761);
or U2560 (N_2560,N_2211,N_1798);
or U2561 (N_2561,N_424,N_88);
or U2562 (N_2562,N_2465,N_194);
nand U2563 (N_2563,N_2034,N_243);
or U2564 (N_2564,N_2193,N_12);
and U2565 (N_2565,N_1931,N_305);
nor U2566 (N_2566,N_731,N_740);
and U2567 (N_2567,N_394,N_2084);
or U2568 (N_2568,N_1399,N_1528);
nor U2569 (N_2569,N_228,N_2261);
or U2570 (N_2570,N_111,N_110);
and U2571 (N_2571,N_9,N_1294);
or U2572 (N_2572,N_584,N_130);
or U2573 (N_2573,N_1058,N_1249);
or U2574 (N_2574,N_2364,N_651);
or U2575 (N_2575,N_2065,N_2213);
and U2576 (N_2576,N_862,N_1087);
and U2577 (N_2577,N_1474,N_238);
nand U2578 (N_2578,N_2480,N_1624);
nand U2579 (N_2579,N_1241,N_1775);
or U2580 (N_2580,N_1263,N_93);
nor U2581 (N_2581,N_1838,N_702);
or U2582 (N_2582,N_70,N_408);
nor U2583 (N_2583,N_2011,N_1148);
or U2584 (N_2584,N_1353,N_1066);
nand U2585 (N_2585,N_552,N_747);
xnor U2586 (N_2586,N_1187,N_2387);
and U2587 (N_2587,N_2461,N_507);
and U2588 (N_2588,N_1052,N_1637);
or U2589 (N_2589,N_1220,N_280);
or U2590 (N_2590,N_861,N_1776);
or U2591 (N_2591,N_160,N_1813);
nand U2592 (N_2592,N_376,N_719);
nand U2593 (N_2593,N_1914,N_2016);
nor U2594 (N_2594,N_1972,N_2308);
nor U2595 (N_2595,N_393,N_1096);
and U2596 (N_2596,N_1995,N_701);
and U2597 (N_2597,N_44,N_1197);
xnor U2598 (N_2598,N_213,N_1117);
nand U2599 (N_2599,N_1909,N_1215);
nor U2600 (N_2600,N_2228,N_100);
nor U2601 (N_2601,N_763,N_915);
nand U2602 (N_2602,N_2466,N_403);
or U2603 (N_2603,N_1827,N_546);
nor U2604 (N_2604,N_2102,N_954);
or U2605 (N_2605,N_2468,N_1941);
nor U2606 (N_2606,N_2293,N_866);
nand U2607 (N_2607,N_1547,N_840);
nand U2608 (N_2608,N_2190,N_2302);
or U2609 (N_2609,N_1401,N_344);
and U2610 (N_2610,N_1453,N_167);
and U2611 (N_2611,N_1740,N_640);
nor U2612 (N_2612,N_492,N_1127);
and U2613 (N_2613,N_1707,N_2200);
nand U2614 (N_2614,N_631,N_1206);
nand U2615 (N_2615,N_858,N_173);
xor U2616 (N_2616,N_2270,N_790);
and U2617 (N_2617,N_532,N_1120);
and U2618 (N_2618,N_1397,N_863);
nor U2619 (N_2619,N_1473,N_1810);
or U2620 (N_2620,N_1076,N_446);
nand U2621 (N_2621,N_1361,N_1934);
and U2622 (N_2622,N_1216,N_1984);
and U2623 (N_2623,N_1403,N_147);
xor U2624 (N_2624,N_199,N_759);
nand U2625 (N_2625,N_1328,N_306);
or U2626 (N_2626,N_1883,N_1088);
nor U2627 (N_2627,N_1631,N_1383);
and U2628 (N_2628,N_1849,N_4);
nor U2629 (N_2629,N_65,N_2240);
and U2630 (N_2630,N_89,N_115);
nand U2631 (N_2631,N_2029,N_2186);
or U2632 (N_2632,N_2418,N_303);
nand U2633 (N_2633,N_1794,N_8);
nand U2634 (N_2634,N_1326,N_444);
and U2635 (N_2635,N_338,N_1565);
nor U2636 (N_2636,N_1261,N_114);
and U2637 (N_2637,N_294,N_1629);
and U2638 (N_2638,N_1584,N_148);
or U2639 (N_2639,N_1105,N_1507);
and U2640 (N_2640,N_610,N_2401);
nor U2641 (N_2641,N_1213,N_1057);
or U2642 (N_2642,N_1365,N_1650);
nand U2643 (N_2643,N_1510,N_307);
nand U2644 (N_2644,N_2379,N_2122);
nand U2645 (N_2645,N_1293,N_1010);
or U2646 (N_2646,N_1375,N_471);
xor U2647 (N_2647,N_328,N_664);
or U2648 (N_2648,N_2166,N_467);
nor U2649 (N_2649,N_938,N_1374);
nand U2650 (N_2650,N_1517,N_1494);
and U2651 (N_2651,N_875,N_1428);
nor U2652 (N_2652,N_2274,N_970);
xor U2653 (N_2653,N_1072,N_34);
nor U2654 (N_2654,N_1053,N_935);
nor U2655 (N_2655,N_1758,N_289);
or U2656 (N_2656,N_169,N_485);
or U2657 (N_2657,N_636,N_1444);
or U2658 (N_2658,N_956,N_99);
and U2659 (N_2659,N_2239,N_135);
and U2660 (N_2660,N_700,N_1607);
or U2661 (N_2661,N_733,N_544);
and U2662 (N_2662,N_1929,N_1723);
nor U2663 (N_2663,N_516,N_1376);
nor U2664 (N_2664,N_2457,N_1172);
nor U2665 (N_2665,N_810,N_538);
nand U2666 (N_2666,N_1410,N_940);
or U2667 (N_2667,N_991,N_2235);
nand U2668 (N_2668,N_2316,N_1068);
and U2669 (N_2669,N_750,N_29);
and U2670 (N_2670,N_794,N_1133);
or U2671 (N_2671,N_709,N_2093);
or U2672 (N_2672,N_657,N_1304);
and U2673 (N_2673,N_2215,N_2427);
nand U2674 (N_2674,N_2244,N_1898);
nand U2675 (N_2675,N_902,N_136);
nor U2676 (N_2676,N_891,N_697);
or U2677 (N_2677,N_869,N_132);
and U2678 (N_2678,N_325,N_987);
nand U2679 (N_2679,N_563,N_1286);
or U2680 (N_2680,N_767,N_1946);
and U2681 (N_2681,N_2287,N_198);
and U2682 (N_2682,N_574,N_905);
nor U2683 (N_2683,N_1874,N_942);
or U2684 (N_2684,N_1933,N_1051);
and U2685 (N_2685,N_2403,N_1270);
nor U2686 (N_2686,N_896,N_1344);
nor U2687 (N_2687,N_1947,N_1106);
and U2688 (N_2688,N_821,N_601);
or U2689 (N_2689,N_1209,N_273);
nor U2690 (N_2690,N_1067,N_941);
nor U2691 (N_2691,N_1048,N_824);
and U2692 (N_2692,N_1884,N_803);
and U2693 (N_2693,N_1654,N_52);
and U2694 (N_2694,N_221,N_1003);
nand U2695 (N_2695,N_556,N_1039);
or U2696 (N_2696,N_1070,N_1099);
nor U2697 (N_2697,N_1784,N_855);
nor U2698 (N_2698,N_487,N_2271);
or U2699 (N_2699,N_1795,N_1082);
nand U2700 (N_2700,N_2053,N_497);
nor U2701 (N_2701,N_1773,N_798);
and U2702 (N_2702,N_834,N_479);
nand U2703 (N_2703,N_1549,N_128);
and U2704 (N_2704,N_1590,N_2091);
and U2705 (N_2705,N_877,N_2454);
or U2706 (N_2706,N_2139,N_462);
and U2707 (N_2707,N_1904,N_1566);
and U2708 (N_2708,N_220,N_2266);
nor U2709 (N_2709,N_1207,N_1621);
or U2710 (N_2710,N_1450,N_2336);
or U2711 (N_2711,N_1183,N_2298);
or U2712 (N_2712,N_1692,N_2191);
or U2713 (N_2713,N_224,N_663);
nor U2714 (N_2714,N_899,N_880);
and U2715 (N_2715,N_2320,N_2149);
nor U2716 (N_2716,N_2231,N_2407);
or U2717 (N_2717,N_451,N_1689);
or U2718 (N_2718,N_1081,N_414);
nand U2719 (N_2719,N_410,N_1644);
nand U2720 (N_2720,N_1322,N_815);
or U2721 (N_2721,N_490,N_509);
nand U2722 (N_2722,N_2214,N_704);
nor U2723 (N_2723,N_2435,N_1586);
and U2724 (N_2724,N_87,N_60);
nor U2725 (N_2725,N_2471,N_628);
and U2726 (N_2726,N_578,N_1520);
or U2727 (N_2727,N_1880,N_458);
or U2728 (N_2728,N_1219,N_748);
nor U2729 (N_2729,N_814,N_1515);
nor U2730 (N_2730,N_1466,N_972);
or U2731 (N_2731,N_1281,N_1377);
and U2732 (N_2732,N_336,N_1819);
nand U2733 (N_2733,N_1809,N_2155);
xor U2734 (N_2734,N_1182,N_1938);
and U2735 (N_2735,N_2323,N_2265);
and U2736 (N_2736,N_1338,N_2046);
or U2737 (N_2737,N_453,N_503);
nor U2738 (N_2738,N_1086,N_1953);
nor U2739 (N_2739,N_553,N_2141);
nand U2740 (N_2740,N_1866,N_714);
nor U2741 (N_2741,N_2385,N_316);
and U2742 (N_2742,N_1333,N_1845);
or U2743 (N_2743,N_1711,N_1038);
and U2744 (N_2744,N_2055,N_463);
nand U2745 (N_2745,N_1415,N_335);
and U2746 (N_2746,N_1368,N_1308);
nor U2747 (N_2747,N_784,N_301);
nor U2748 (N_2748,N_1400,N_1661);
or U2749 (N_2749,N_1824,N_1);
or U2750 (N_2750,N_2377,N_1881);
nor U2751 (N_2751,N_2444,N_1955);
nor U2752 (N_2752,N_758,N_1716);
nor U2753 (N_2753,N_2460,N_620);
nor U2754 (N_2754,N_1548,N_1901);
and U2755 (N_2755,N_241,N_982);
xnor U2756 (N_2756,N_1483,N_835);
nand U2757 (N_2757,N_1306,N_1935);
and U2758 (N_2758,N_1539,N_2491);
nand U2759 (N_2759,N_1899,N_2243);
nor U2760 (N_2760,N_127,N_297);
and U2761 (N_2761,N_1564,N_2337);
nor U2762 (N_2762,N_64,N_2382);
nand U2763 (N_2763,N_775,N_1465);
or U2764 (N_2764,N_1872,N_1063);
and U2765 (N_2765,N_2241,N_2246);
nor U2766 (N_2766,N_619,N_1289);
or U2767 (N_2767,N_427,N_1493);
nand U2768 (N_2768,N_1158,N_473);
nand U2769 (N_2769,N_641,N_2236);
nand U2770 (N_2770,N_2426,N_47);
nor U2771 (N_2771,N_2497,N_250);
and U2772 (N_2772,N_1089,N_2340);
nor U2773 (N_2773,N_1917,N_957);
and U2774 (N_2774,N_1029,N_2109);
or U2775 (N_2775,N_2356,N_859);
and U2776 (N_2776,N_669,N_2318);
nor U2777 (N_2777,N_886,N_432);
nor U2778 (N_2778,N_369,N_1451);
nand U2779 (N_2779,N_1214,N_2359);
and U2780 (N_2780,N_121,N_2115);
nor U2781 (N_2781,N_2386,N_153);
nand U2782 (N_2782,N_1169,N_1768);
xnor U2783 (N_2783,N_2317,N_2459);
nor U2784 (N_2784,N_166,N_2182);
and U2785 (N_2785,N_590,N_2448);
or U2786 (N_2786,N_183,N_1372);
or U2787 (N_2787,N_107,N_1447);
nand U2788 (N_2788,N_252,N_826);
or U2789 (N_2789,N_936,N_86);
nand U2790 (N_2790,N_1324,N_1656);
nand U2791 (N_2791,N_1567,N_1876);
and U2792 (N_2792,N_1657,N_925);
or U2793 (N_2793,N_2060,N_2446);
nand U2794 (N_2794,N_2179,N_1427);
nor U2795 (N_2795,N_1648,N_1856);
nand U2796 (N_2796,N_2409,N_841);
or U2797 (N_2797,N_1731,N_1118);
nand U2798 (N_2798,N_1942,N_543);
nor U2799 (N_2799,N_833,N_1753);
nand U2800 (N_2800,N_245,N_2372);
and U2801 (N_2801,N_392,N_1178);
nand U2802 (N_2802,N_1497,N_2090);
and U2803 (N_2803,N_124,N_901);
or U2804 (N_2804,N_1468,N_2363);
or U2805 (N_2805,N_1958,N_558);
nand U2806 (N_2806,N_260,N_2496);
and U2807 (N_2807,N_367,N_382);
or U2808 (N_2808,N_1682,N_2140);
nand U2809 (N_2809,N_248,N_1643);
nand U2810 (N_2810,N_2004,N_1339);
and U2811 (N_2811,N_1759,N_2424);
or U2812 (N_2812,N_955,N_1992);
nor U2813 (N_2813,N_1814,N_356);
nor U2814 (N_2814,N_1258,N_2487);
and U2815 (N_2815,N_1228,N_515);
nor U2816 (N_2816,N_2116,N_1006);
and U2817 (N_2817,N_140,N_1925);
nor U2818 (N_2818,N_2378,N_2260);
nor U2819 (N_2819,N_2108,N_1445);
nor U2820 (N_2820,N_616,N_623);
nand U2821 (N_2821,N_1442,N_1913);
nor U2822 (N_2822,N_2104,N_1327);
nand U2823 (N_2823,N_1005,N_1820);
and U2824 (N_2824,N_292,N_2007);
nor U2825 (N_2825,N_1464,N_692);
and U2826 (N_2826,N_712,N_1248);
nor U2827 (N_2827,N_419,N_582);
and U2828 (N_2828,N_2013,N_1893);
nand U2829 (N_2829,N_2389,N_182);
nor U2830 (N_2830,N_2063,N_1748);
and U2831 (N_2831,N_13,N_1595);
nor U2832 (N_2832,N_2258,N_1968);
and U2833 (N_2833,N_2070,N_1093);
and U2834 (N_2834,N_2032,N_926);
nand U2835 (N_2835,N_366,N_1406);
and U2836 (N_2836,N_90,N_1770);
nand U2837 (N_2837,N_375,N_1458);
and U2838 (N_2838,N_650,N_2105);
and U2839 (N_2839,N_1181,N_1491);
nand U2840 (N_2840,N_654,N_1446);
nand U2841 (N_2841,N_2118,N_117);
and U2842 (N_2842,N_2351,N_1069);
or U2843 (N_2843,N_357,N_1439);
xnor U2844 (N_2844,N_1459,N_152);
nor U2845 (N_2845,N_1936,N_1392);
nor U2846 (N_2846,N_572,N_1085);
and U2847 (N_2847,N_2451,N_1257);
or U2848 (N_2848,N_40,N_2473);
or U2849 (N_2849,N_484,N_499);
or U2850 (N_2850,N_255,N_168);
nor U2851 (N_2851,N_156,N_897);
or U2852 (N_2852,N_1479,N_1298);
and U2853 (N_2853,N_1211,N_1132);
and U2854 (N_2854,N_1134,N_2202);
or U2855 (N_2855,N_2037,N_2);
or U2856 (N_2856,N_1982,N_22);
nor U2857 (N_2857,N_1930,N_1012);
and U2858 (N_2858,N_1949,N_1223);
nand U2859 (N_2859,N_2165,N_626);
or U2860 (N_2860,N_913,N_258);
or U2861 (N_2861,N_953,N_2018);
and U2862 (N_2862,N_53,N_1389);
nand U2863 (N_2863,N_1605,N_2475);
nand U2864 (N_2864,N_512,N_486);
nand U2865 (N_2865,N_1062,N_1243);
or U2866 (N_2866,N_468,N_1275);
nor U2867 (N_2867,N_276,N_358);
nor U2868 (N_2868,N_1647,N_215);
nand U2869 (N_2869,N_1552,N_425);
nor U2870 (N_2870,N_908,N_1652);
and U2871 (N_2871,N_757,N_383);
nor U2872 (N_2872,N_137,N_402);
nor U2873 (N_2873,N_300,N_943);
nand U2874 (N_2874,N_129,N_679);
nand U2875 (N_2875,N_2410,N_2411);
and U2876 (N_2876,N_207,N_244);
nor U2877 (N_2877,N_1430,N_1190);
and U2878 (N_2878,N_1890,N_932);
and U2879 (N_2879,N_202,N_2344);
nand U2880 (N_2880,N_2429,N_2100);
or U2881 (N_2881,N_978,N_265);
or U2882 (N_2882,N_1040,N_716);
and U2883 (N_2883,N_1987,N_347);
nand U2884 (N_2884,N_109,N_673);
nand U2885 (N_2885,N_460,N_760);
nor U2886 (N_2886,N_1642,N_919);
nor U2887 (N_2887,N_1699,N_1997);
or U2888 (N_2888,N_592,N_74);
nand U2889 (N_2889,N_611,N_870);
nor U2890 (N_2890,N_2147,N_2189);
and U2891 (N_2891,N_629,N_1409);
or U2892 (N_2892,N_526,N_2173);
and U2893 (N_2893,N_1416,N_1354);
and U2894 (N_2894,N_2284,N_612);
and U2895 (N_2895,N_873,N_498);
nand U2896 (N_2896,N_1568,N_254);
xor U2897 (N_2897,N_1556,N_890);
nand U2898 (N_2898,N_964,N_165);
and U2899 (N_2899,N_263,N_2077);
or U2900 (N_2900,N_1367,N_1073);
nand U2901 (N_2901,N_1033,N_3);
and U2902 (N_2902,N_776,N_62);
nor U2903 (N_2903,N_652,N_1673);
nor U2904 (N_2904,N_635,N_1502);
nand U2905 (N_2905,N_441,N_1046);
or U2906 (N_2906,N_416,N_565);
and U2907 (N_2907,N_1840,N_38);
and U2908 (N_2908,N_240,N_1791);
and U2909 (N_2909,N_727,N_181);
and U2910 (N_2910,N_2120,N_283);
or U2911 (N_2911,N_892,N_1886);
nand U2912 (N_2912,N_1448,N_2230);
nand U2913 (N_2913,N_214,N_355);
nor U2914 (N_2914,N_541,N_1765);
or U2915 (N_2915,N_66,N_2148);
nor U2916 (N_2916,N_1690,N_1969);
or U2917 (N_2917,N_363,N_1380);
nor U2918 (N_2918,N_969,N_1176);
or U2919 (N_2919,N_726,N_1971);
nand U2920 (N_2920,N_1164,N_1269);
or U2921 (N_2921,N_365,N_1104);
nor U2922 (N_2922,N_184,N_1769);
and U2923 (N_2923,N_615,N_293);
nor U2924 (N_2924,N_744,N_1109);
nand U2925 (N_2925,N_278,N_14);
or U2926 (N_2926,N_2449,N_2368);
nand U2927 (N_2927,N_1800,N_576);
nand U2928 (N_2928,N_2488,N_881);
nand U2929 (N_2929,N_1009,N_333);
and U2930 (N_2930,N_743,N_268);
and U2931 (N_2931,N_175,N_1578);
and U2932 (N_2932,N_372,N_1574);
nor U2933 (N_2933,N_83,N_1208);
or U2934 (N_2934,N_2039,N_2499);
nor U2935 (N_2935,N_2432,N_178);
nand U2936 (N_2936,N_1267,N_966);
nor U2937 (N_2937,N_1571,N_2399);
or U2938 (N_2938,N_288,N_508);
nor U2939 (N_2939,N_75,N_1633);
nand U2940 (N_2940,N_2197,N_1885);
nand U2941 (N_2941,N_431,N_646);
and U2942 (N_2942,N_1092,N_2218);
and U2943 (N_2943,N_493,N_1264);
or U2944 (N_2944,N_1419,N_2474);
nand U2945 (N_2945,N_1577,N_2137);
nor U2946 (N_2946,N_906,N_381);
and U2947 (N_2947,N_2392,N_1390);
and U2948 (N_2948,N_1245,N_229);
and U2949 (N_2949,N_341,N_1764);
nand U2950 (N_2950,N_1725,N_2201);
nand U2951 (N_2951,N_488,N_2168);
nor U2952 (N_2952,N_1369,N_1921);
or U2953 (N_2953,N_511,N_1816);
or U2954 (N_2954,N_540,N_1527);
nand U2955 (N_2955,N_1541,N_2479);
nand U2956 (N_2956,N_1569,N_443);
or U2957 (N_2957,N_1391,N_19);
nor U2958 (N_2958,N_1659,N_879);
nand U2959 (N_2959,N_1470,N_236);
nand U2960 (N_2960,N_736,N_43);
nor U2961 (N_2961,N_2408,N_1671);
or U2962 (N_2962,N_1168,N_2415);
nor U2963 (N_2963,N_161,N_118);
nand U2964 (N_2964,N_561,N_1179);
or U2965 (N_2965,N_1115,N_1627);
or U2966 (N_2966,N_754,N_1441);
or U2967 (N_2967,N_1665,N_35);
nand U2968 (N_2968,N_568,N_1687);
nor U2969 (N_2969,N_1818,N_1894);
and U2970 (N_2970,N_2249,N_350);
or U2971 (N_2971,N_465,N_61);
and U2972 (N_2972,N_190,N_1970);
nor U2973 (N_2973,N_1858,N_537);
nor U2974 (N_2974,N_1734,N_2003);
or U2975 (N_2975,N_1329,N_1513);
or U2976 (N_2976,N_1922,N_2101);
nor U2977 (N_2977,N_1545,N_2152);
and U2978 (N_2978,N_1425,N_1149);
and U2979 (N_2979,N_688,N_330);
xor U2980 (N_2980,N_2045,N_2309);
or U2981 (N_2981,N_1514,N_143);
or U2982 (N_2982,N_2079,N_361);
or U2983 (N_2983,N_2282,N_353);
or U2984 (N_2984,N_1091,N_2089);
and U2985 (N_2985,N_1836,N_2292);
xor U2986 (N_2986,N_2047,N_420);
and U2987 (N_2987,N_436,N_822);
nor U2988 (N_2988,N_1456,N_557);
nand U2989 (N_2989,N_2125,N_266);
and U2990 (N_2990,N_1873,N_1695);
nand U2991 (N_2991,N_2489,N_1783);
nor U2992 (N_2992,N_1524,N_1782);
nand U2993 (N_2993,N_1625,N_2273);
and U2994 (N_2994,N_2113,N_2352);
nor U2995 (N_2995,N_1706,N_0);
nor U2996 (N_2996,N_1617,N_2027);
nand U2997 (N_2997,N_722,N_723);
or U2998 (N_2998,N_2028,N_1075);
or U2999 (N_2999,N_1454,N_331);
or U3000 (N_3000,N_614,N_2126);
nor U3001 (N_3001,N_1140,N_304);
nand U3002 (N_3002,N_586,N_2000);
and U3003 (N_3003,N_1582,N_2278);
and U3004 (N_3004,N_489,N_31);
nor U3005 (N_3005,N_2478,N_2291);
and U3006 (N_3006,N_608,N_162);
and U3007 (N_3007,N_1019,N_2048);
and U3008 (N_3008,N_1234,N_1229);
or U3009 (N_3009,N_1755,N_2251);
or U3010 (N_3010,N_2159,N_1926);
and U3011 (N_3011,N_1256,N_2082);
and U3012 (N_3012,N_1988,N_725);
and U3013 (N_3013,N_345,N_2406);
nor U3014 (N_3014,N_1806,N_1870);
and U3015 (N_3015,N_1312,N_1171);
nor U3016 (N_3016,N_2428,N_2438);
and U3017 (N_3017,N_1609,N_104);
xor U3018 (N_3018,N_560,N_1841);
or U3019 (N_3019,N_2188,N_1685);
nor U3020 (N_3020,N_2321,N_2367);
nand U3021 (N_3021,N_602,N_1679);
nand U3022 (N_3022,N_496,N_2440);
nand U3023 (N_3023,N_191,N_1653);
nor U3024 (N_3024,N_1945,N_1366);
nor U3025 (N_3025,N_1603,N_1743);
nor U3026 (N_3026,N_342,N_1314);
nor U3027 (N_3027,N_1200,N_2374);
nand U3028 (N_3028,N_2472,N_1260);
nand U3029 (N_3029,N_1424,N_948);
and U3030 (N_3030,N_78,N_1443);
nor U3031 (N_3031,N_352,N_604);
and U3032 (N_3032,N_1788,N_2275);
nor U3033 (N_3033,N_1337,N_2307);
and U3034 (N_3034,N_505,N_668);
and U3035 (N_3035,N_751,N_1635);
or U3036 (N_3036,N_766,N_1634);
or U3037 (N_3037,N_1518,N_1932);
nand U3038 (N_3038,N_1897,N_549);
nand U3039 (N_3039,N_1576,N_2312);
nand U3040 (N_3040,N_1056,N_749);
nor U3041 (N_3041,N_1462,N_1559);
nor U3042 (N_3042,N_1583,N_945);
and U3043 (N_3043,N_251,N_536);
nand U3044 (N_3044,N_659,N_1230);
or U3045 (N_3045,N_277,N_116);
and U3046 (N_3046,N_1268,N_2391);
nand U3047 (N_3047,N_261,N_2080);
nor U3048 (N_3048,N_1993,N_1792);
or U3049 (N_3049,N_2434,N_1646);
or U3050 (N_3050,N_2425,N_2484);
nor U3051 (N_3051,N_1512,N_554);
and U3052 (N_3052,N_1340,N_1145);
nand U3053 (N_3053,N_1944,N_947);
and U3054 (N_3054,N_1130,N_2206);
nor U3055 (N_3055,N_1839,N_2262);
or U3056 (N_3056,N_530,N_1094);
or U3057 (N_3057,N_1757,N_1318);
or U3058 (N_3058,N_1508,N_2464);
nand U3059 (N_3059,N_1131,N_2127);
nor U3060 (N_3060,N_1499,N_849);
or U3061 (N_3061,N_524,N_1486);
nand U3062 (N_3062,N_1177,N_1728);
or U3063 (N_3063,N_1173,N_1868);
or U3064 (N_3064,N_1546,N_455);
nand U3065 (N_3065,N_84,N_1618);
or U3066 (N_3066,N_742,N_373);
nor U3067 (N_3067,N_823,N_1055);
nor U3068 (N_3068,N_1021,N_1747);
and U3069 (N_3069,N_865,N_1279);
and U3070 (N_3070,N_2431,N_1786);
nand U3071 (N_3071,N_1903,N_2031);
nand U3072 (N_3072,N_728,N_518);
and U3073 (N_3073,N_618,N_359);
nand U3074 (N_3074,N_105,N_322);
or U3075 (N_3075,N_1084,N_729);
and U3076 (N_3076,N_1610,N_141);
and U3077 (N_3077,N_975,N_2267);
or U3078 (N_3078,N_2430,N_2483);
or U3079 (N_3079,N_1771,N_371);
nand U3080 (N_3080,N_477,N_1244);
nor U3081 (N_3081,N_1581,N_1498);
nor U3082 (N_3082,N_2022,N_71);
nand U3083 (N_3083,N_1004,N_598);
nand U3084 (N_3084,N_2121,N_206);
or U3085 (N_3085,N_1735,N_2494);
nor U3086 (N_3086,N_409,N_1166);
nor U3087 (N_3087,N_1271,N_694);
nand U3088 (N_3088,N_1475,N_1976);
nor U3089 (N_3089,N_893,N_2074);
or U3090 (N_3090,N_1259,N_1888);
or U3091 (N_3091,N_1817,N_470);
nand U3092 (N_3092,N_491,N_779);
nand U3093 (N_3093,N_1604,N_684);
and U3094 (N_3094,N_1772,N_2397);
nand U3095 (N_3095,N_171,N_1906);
nor U3096 (N_3096,N_2072,N_223);
and U3097 (N_3097,N_2482,N_1205);
nand U3098 (N_3098,N_2111,N_192);
or U3099 (N_3099,N_2445,N_564);
nand U3100 (N_3100,N_1703,N_1250);
nand U3101 (N_3101,N_825,N_1394);
nor U3102 (N_3102,N_1896,N_778);
nand U3103 (N_3103,N_1355,N_1273);
nand U3104 (N_3104,N_1481,N_11);
or U3105 (N_3105,N_1018,N_1460);
nor U3106 (N_3106,N_1965,N_2381);
or U3107 (N_3107,N_2059,N_2207);
nor U3108 (N_3108,N_1575,N_1908);
nor U3109 (N_3109,N_706,N_2138);
nor U3110 (N_3110,N_2061,N_1860);
nor U3111 (N_3111,N_852,N_1877);
or U3112 (N_3112,N_1385,N_950);
or U3113 (N_3113,N_1825,N_2123);
nand U3114 (N_3114,N_1821,N_2248);
and U3115 (N_3115,N_1954,N_326);
and U3116 (N_3116,N_327,N_958);
nand U3117 (N_3117,N_321,N_1655);
nor U3118 (N_3118,N_415,N_1011);
and U3119 (N_3119,N_730,N_1108);
or U3120 (N_3120,N_996,N_910);
or U3121 (N_3121,N_17,N_320);
and U3122 (N_3122,N_1323,N_1693);
nand U3123 (N_3123,N_1153,N_314);
or U3124 (N_3124,N_872,N_680);
or U3125 (N_3125,N_1887,N_1746);
and U3126 (N_3126,N_1283,N_1668);
or U3127 (N_3127,N_724,N_1680);
nor U3128 (N_3128,N_1660,N_1147);
nand U3129 (N_3129,N_1420,N_112);
and U3130 (N_3130,N_985,N_1619);
or U3131 (N_3131,N_2208,N_63);
or U3132 (N_3132,N_189,N_1697);
and U3133 (N_3133,N_1879,N_2119);
and U3134 (N_3134,N_1503,N_937);
nand U3135 (N_3135,N_2162,N_1822);
or U3136 (N_3136,N_961,N_2221);
or U3137 (N_3137,N_1429,N_459);
nor U3138 (N_3138,N_788,N_1395);
and U3139 (N_3139,N_2436,N_466);
nor U3140 (N_3140,N_603,N_1097);
nor U3141 (N_3141,N_816,N_644);
and U3142 (N_3142,N_1265,N_656);
nand U3143 (N_3143,N_411,N_514);
nand U3144 (N_3144,N_1589,N_227);
nand U3145 (N_3145,N_1347,N_1325);
nand U3146 (N_3146,N_2001,N_1918);
nand U3147 (N_3147,N_275,N_1246);
or U3148 (N_3148,N_378,N_1550);
nand U3149 (N_3149,N_1891,N_1967);
nand U3150 (N_3150,N_1119,N_203);
xor U3151 (N_3151,N_627,N_2301);
nand U3152 (N_3152,N_1756,N_1364);
nand U3153 (N_3153,N_412,N_1013);
or U3154 (N_3154,N_1952,N_2198);
nand U3155 (N_3155,N_478,N_617);
and U3156 (N_3156,N_1843,N_2212);
and U3157 (N_3157,N_808,N_800);
and U3158 (N_3158,N_1100,N_2002);
or U3159 (N_3159,N_698,N_387);
nand U3160 (N_3160,N_310,N_1334);
or U3161 (N_3161,N_1139,N_1146);
or U3162 (N_3162,N_1867,N_1781);
or U3163 (N_3163,N_1951,N_1534);
nand U3164 (N_3164,N_917,N_720);
nor U3165 (N_3165,N_2237,N_2124);
nand U3166 (N_3166,N_1438,N_149);
and U3167 (N_3167,N_2294,N_738);
nand U3168 (N_3168,N_2209,N_1254);
or U3169 (N_3169,N_1017,N_2419);
or U3170 (N_3170,N_755,N_246);
and U3171 (N_3171,N_1540,N_146);
nor U3172 (N_3172,N_1159,N_205);
and U3173 (N_3173,N_1461,N_1174);
and U3174 (N_3174,N_1752,N_2020);
or U3175 (N_3175,N_689,N_2437);
nor U3176 (N_3176,N_395,N_1760);
nand U3177 (N_3177,N_2036,N_2360);
nand U3178 (N_3178,N_1912,N_2005);
and U3179 (N_3179,N_399,N_1506);
nor U3180 (N_3180,N_1960,N_222);
nor U3181 (N_3181,N_682,N_1123);
or U3182 (N_3182,N_418,N_667);
nand U3183 (N_3183,N_1985,N_2224);
nor U3184 (N_3184,N_1688,N_1892);
and U3185 (N_3185,N_2075,N_597);
nand U3186 (N_3186,N_921,N_2299);
nand U3187 (N_3187,N_2232,N_1645);
or U3188 (N_3188,N_247,N_217);
and U3189 (N_3189,N_559,N_649);
nand U3190 (N_3190,N_535,N_2184);
or U3191 (N_3191,N_1015,N_2277);
nand U3192 (N_3192,N_2158,N_67);
xnor U3193 (N_3193,N_270,N_1495);
or U3194 (N_3194,N_2154,N_1433);
or U3195 (N_3195,N_2167,N_1767);
nor U3196 (N_3196,N_1349,N_1436);
nand U3197 (N_3197,N_2355,N_2087);
and U3198 (N_3198,N_1343,N_1226);
and U3199 (N_3199,N_1237,N_475);
and U3200 (N_3200,N_20,N_2433);
or U3201 (N_3201,N_676,N_2470);
or U3202 (N_3202,N_2328,N_2313);
nand U3203 (N_3203,N_430,N_7);
nand U3204 (N_3204,N_979,N_2143);
or U3205 (N_3205,N_2255,N_2269);
nand U3206 (N_3206,N_73,N_1192);
nor U3207 (N_3207,N_2187,N_1677);
nand U3208 (N_3208,N_317,N_2279);
nand U3209 (N_3209,N_389,N_1240);
or U3210 (N_3210,N_1608,N_1193);
nor U3211 (N_3211,N_632,N_318);
nor U3212 (N_3212,N_1718,N_1080);
and U3213 (N_3213,N_483,N_844);
nand U3214 (N_3214,N_1684,N_1332);
or U3215 (N_3215,N_2145,N_1778);
or U3216 (N_3216,N_1712,N_133);
nand U3217 (N_3217,N_1986,N_2306);
and U3218 (N_3218,N_609,N_204);
nor U3219 (N_3219,N_707,N_76);
and U3220 (N_3220,N_1407,N_2069);
nand U3221 (N_3221,N_1079,N_21);
nor U3222 (N_3222,N_1457,N_131);
or U3223 (N_3223,N_1686,N_1382);
nor U3224 (N_3224,N_594,N_703);
nor U3225 (N_3225,N_853,N_1316);
xor U3226 (N_3226,N_1227,N_1563);
nand U3227 (N_3227,N_1423,N_1045);
nor U3228 (N_3228,N_1247,N_2073);
nor U3229 (N_3229,N_1191,N_360);
or U3230 (N_3230,N_155,N_151);
nand U3231 (N_3231,N_513,N_1532);
nor U3232 (N_3232,N_139,N_1373);
nand U3233 (N_3233,N_2157,N_571);
nand U3234 (N_3234,N_1150,N_525);
nand U3235 (N_3235,N_1895,N_449);
and U3236 (N_3236,N_1698,N_428);
xnor U3237 (N_3237,N_447,N_787);
and U3238 (N_3238,N_291,N_1418);
or U3239 (N_3239,N_1666,N_119);
and U3240 (N_3240,N_1830,N_1078);
and U3241 (N_3241,N_2456,N_939);
nor U3242 (N_3242,N_469,N_2049);
or U3243 (N_3243,N_1440,N_1225);
xor U3244 (N_3244,N_1696,N_642);
and U3245 (N_3245,N_1125,N_2133);
or U3246 (N_3246,N_1504,N_1722);
nor U3247 (N_3247,N_1787,N_1194);
nand U3248 (N_3248,N_1594,N_786);
or U3249 (N_3249,N_2463,N_868);
or U3250 (N_3250,N_1683,N_569);
nand U3251 (N_3251,N_1516,N_1847);
or U3252 (N_3252,N_648,N_843);
or U3253 (N_3253,N_370,N_888);
nand U3254 (N_3254,N_918,N_272);
nor U3255 (N_3255,N_1059,N_2219);
and U3256 (N_3256,N_256,N_1710);
and U3257 (N_3257,N_142,N_660);
and U3258 (N_3258,N_2394,N_1141);
and U3259 (N_3259,N_1558,N_1032);
nor U3260 (N_3260,N_27,N_1255);
and U3261 (N_3261,N_1796,N_1157);
and U3262 (N_3262,N_2486,N_1994);
nor U3263 (N_3263,N_284,N_354);
or U3264 (N_3264,N_929,N_789);
and U3265 (N_3265,N_1739,N_138);
or U3266 (N_3266,N_1356,N_907);
nand U3267 (N_3267,N_696,N_1136);
nor U3268 (N_3268,N_2257,N_585);
and U3269 (N_3269,N_539,N_384);
nand U3270 (N_3270,N_42,N_1623);
and U3271 (N_3271,N_1165,N_323);
or U3272 (N_3272,N_2009,N_2288);
nor U3273 (N_3273,N_1562,N_1709);
nand U3274 (N_3274,N_1405,N_2442);
or U3275 (N_3275,N_157,N_2150);
nand U3276 (N_3276,N_2339,N_1763);
nand U3277 (N_3277,N_349,N_854);
nand U3278 (N_3278,N_2253,N_1602);
and U3279 (N_3279,N_2019,N_2322);
and U3280 (N_3280,N_120,N_77);
nor U3281 (N_3281,N_1235,N_1300);
nor U3282 (N_3282,N_2324,N_1572);
nand U3283 (N_3283,N_1302,N_613);
or U3284 (N_3284,N_976,N_951);
and U3285 (N_3285,N_1291,N_931);
or U3286 (N_3286,N_2066,N_2146);
and U3287 (N_3287,N_2106,N_312);
nor U3288 (N_3288,N_2014,N_977);
nand U3289 (N_3289,N_1026,N_1490);
and U3290 (N_3290,N_633,N_1212);
nor U3291 (N_3291,N_434,N_806);
xnor U3292 (N_3292,N_695,N_634);
nand U3293 (N_3293,N_102,N_2493);
or U3294 (N_3294,N_1551,N_1875);
nor U3295 (N_3295,N_2238,N_2263);
or U3296 (N_3296,N_2259,N_1606);
nand U3297 (N_3297,N_528,N_1266);
nor U3298 (N_3298,N_2362,N_573);
nand U3299 (N_3299,N_1766,N_1359);
nand U3300 (N_3300,N_1393,N_1278);
nand U3301 (N_3301,N_1203,N_1095);
or U3302 (N_3302,N_1991,N_1754);
nor U3303 (N_3303,N_1485,N_1854);
or U3304 (N_3304,N_832,N_871);
or U3305 (N_3305,N_397,N_2422);
nor U3306 (N_3306,N_828,N_1154);
and U3307 (N_3307,N_2376,N_930);
nor U3308 (N_3308,N_1292,N_180);
nor U3309 (N_3309,N_1948,N_1272);
or U3310 (N_3310,N_1370,N_1320);
and U3311 (N_3311,N_1396,N_756);
and U3312 (N_3312,N_2384,N_1037);
nor U3313 (N_3313,N_400,N_1622);
and U3314 (N_3314,N_655,N_1850);
and U3315 (N_3315,N_398,N_1388);
or U3316 (N_3316,N_1331,N_542);
and U3317 (N_3317,N_782,N_2156);
nand U3318 (N_3318,N_1455,N_599);
nor U3319 (N_3319,N_1184,N_1599);
nor U3320 (N_3320,N_2099,N_1842);
nand U3321 (N_3321,N_334,N_2095);
or U3322 (N_3322,N_687,N_2112);
xor U3323 (N_3323,N_927,N_1102);
nand U3324 (N_3324,N_495,N_764);
and U3325 (N_3325,N_113,N_26);
nand U3326 (N_3326,N_126,N_1253);
nor U3327 (N_3327,N_1167,N_2346);
and U3328 (N_3328,N_2172,N_32);
or U3329 (N_3329,N_864,N_2195);
nor U3330 (N_3330,N_2071,N_1557);
nor U3331 (N_3331,N_1330,N_2056);
nand U3332 (N_3332,N_2268,N_45);
nor U3333 (N_3333,N_1630,N_271);
nand U3334 (N_3334,N_362,N_1142);
or U3335 (N_3335,N_867,N_1708);
nand U3336 (N_3336,N_949,N_1579);
nand U3337 (N_3337,N_1526,N_1844);
nand U3338 (N_3338,N_1348,N_1831);
or U3339 (N_3339,N_2250,N_2310);
nand U3340 (N_3340,N_2083,N_878);
nand U3341 (N_3341,N_134,N_1044);
nor U3342 (N_3342,N_593,N_677);
nand U3343 (N_3343,N_2423,N_1199);
and U3344 (N_3344,N_1452,N_2256);
and U3345 (N_3345,N_1007,N_385);
and U3346 (N_3346,N_1889,N_2107);
and U3347 (N_3347,N_1705,N_2295);
nor U3348 (N_3348,N_1835,N_653);
nor U3349 (N_3349,N_445,N_811);
nand U3350 (N_3350,N_262,N_216);
or U3351 (N_3351,N_2314,N_123);
nand U3352 (N_3352,N_1990,N_1116);
nor U3353 (N_3353,N_2151,N_998);
nand U3354 (N_3354,N_59,N_1155);
and U3355 (N_3355,N_2131,N_474);
xor U3356 (N_3356,N_46,N_638);
or U3357 (N_3357,N_1750,N_188);
and U3358 (N_3358,N_596,N_2174);
nor U3359 (N_3359,N_1098,N_2025);
and U3360 (N_3360,N_997,N_2183);
and U3361 (N_3361,N_269,N_2455);
nand U3362 (N_3362,N_1694,N_2289);
or U3363 (N_3363,N_710,N_2114);
nor U3364 (N_3364,N_1449,N_2286);
nand U3365 (N_3365,N_745,N_2341);
nand U3366 (N_3366,N_197,N_299);
nand U3367 (N_3367,N_1977,N_2134);
or U3368 (N_3368,N_1296,N_993);
or U3369 (N_3369,N_647,N_2033);
nand U3370 (N_3370,N_1251,N_172);
or U3371 (N_3371,N_422,N_1384);
nor U3372 (N_3372,N_1744,N_1780);
and U3373 (N_3373,N_179,N_2040);
and U3374 (N_3374,N_1001,N_946);
and U3375 (N_3375,N_555,N_311);
nand U3376 (N_3376,N_914,N_922);
nor U3377 (N_3377,N_2220,N_1749);
nor U3378 (N_3378,N_1598,N_2110);
xnor U3379 (N_3379,N_1804,N_1138);
and U3380 (N_3380,N_2247,N_1587);
or U3381 (N_3381,N_302,N_2199);
nand U3382 (N_3382,N_718,N_95);
and U3383 (N_3383,N_1981,N_2361);
and U3384 (N_3384,N_324,N_1144);
nor U3385 (N_3385,N_1239,N_2178);
nand U3386 (N_3386,N_1980,N_2375);
or U3387 (N_3387,N_2062,N_1411);
and U3388 (N_3388,N_2136,N_771);
nand U3389 (N_3389,N_622,N_797);
nand U3390 (N_3390,N_2338,N_807);
or U3391 (N_3391,N_2050,N_607);
nand U3392 (N_3392,N_639,N_379);
or U3393 (N_3393,N_1833,N_170);
xnor U3394 (N_3394,N_2103,N_339);
or U3395 (N_3395,N_960,N_517);
nor U3396 (N_3396,N_674,N_933);
and U3397 (N_3397,N_296,N_1596);
nor U3398 (N_3398,N_1832,N_1288);
and U3399 (N_3399,N_2400,N_1871);
and U3400 (N_3400,N_2413,N_309);
nor U3401 (N_3401,N_54,N_2176);
or U3402 (N_3402,N_200,N_2160);
and U3403 (N_3403,N_2396,N_346);
nor U3404 (N_3404,N_753,N_2242);
or U3405 (N_3405,N_1531,N_440);
and U3406 (N_3406,N_675,N_735);
nand U3407 (N_3407,N_2452,N_1218);
and U3408 (N_3408,N_2371,N_1615);
nor U3409 (N_3409,N_1422,N_1789);
nor U3410 (N_3410,N_1701,N_1905);
and U3411 (N_3411,N_920,N_857);
nor U3412 (N_3412,N_2094,N_1002);
or U3413 (N_3413,N_836,N_1352);
and U3414 (N_3414,N_158,N_846);
or U3415 (N_3415,N_1726,N_1943);
and U3416 (N_3416,N_900,N_438);
and U3417 (N_3417,N_1014,N_637);
or U3418 (N_3418,N_2343,N_1204);
and U3419 (N_3419,N_2161,N_1061);
and U3420 (N_3420,N_721,N_1195);
nor U3421 (N_3421,N_2216,N_2233);
nand U3422 (N_3422,N_1907,N_1924);
nand U3423 (N_3423,N_1402,N_1628);
or U3424 (N_3424,N_2332,N_2030);
nand U3425 (N_3425,N_1161,N_1350);
nor U3426 (N_3426,N_80,N_2038);
nand U3427 (N_3427,N_212,N_1107);
nor U3428 (N_3428,N_1492,N_1593);
nand U3429 (N_3429,N_1927,N_1779);
nor U3430 (N_3430,N_1801,N_1358);
and U3431 (N_3431,N_1111,N_201);
nor U3432 (N_3432,N_1509,N_2416);
nor U3433 (N_3433,N_1224,N_1077);
and U3434 (N_3434,N_235,N_1342);
nand U3435 (N_3435,N_2333,N_2092);
and U3436 (N_3436,N_1658,N_1233);
nand U3437 (N_3437,N_1309,N_661);
and U3438 (N_3438,N_159,N_81);
and U3439 (N_3439,N_1371,N_630);
and U3440 (N_3440,N_2398,N_1505);
and U3441 (N_3441,N_1301,N_1882);
nand U3442 (N_3442,N_989,N_551);
and U3443 (N_3443,N_769,N_177);
xor U3444 (N_3444,N_898,N_1638);
nor U3445 (N_3445,N_1742,N_343);
nor U3446 (N_3446,N_1471,N_481);
nor U3447 (N_3447,N_780,N_1834);
nor U3448 (N_3448,N_1730,N_10);
and U3449 (N_3449,N_28,N_2035);
nor U3450 (N_3450,N_1902,N_2326);
and U3451 (N_3451,N_1413,N_5);
nand U3452 (N_3452,N_2347,N_259);
and U3453 (N_3453,N_1803,N_2370);
nand U3454 (N_3454,N_1500,N_522);
nand U3455 (N_3455,N_2281,N_2194);
and U3456 (N_3456,N_2315,N_1489);
nand U3457 (N_3457,N_566,N_842);
or U3458 (N_3458,N_233,N_1983);
and U3459 (N_3459,N_209,N_783);
nor U3460 (N_3460,N_959,N_1065);
and U3461 (N_3461,N_1031,N_2304);
nand U3462 (N_3462,N_1050,N_2180);
and U3463 (N_3463,N_562,N_1519);
nor U3464 (N_3464,N_884,N_1928);
nand U3465 (N_3465,N_995,N_448);
and U3466 (N_3466,N_390,N_407);
or U3467 (N_3467,N_830,N_671);
or U3468 (N_3468,N_1188,N_1315);
and U3469 (N_3469,N_2462,N_1345);
nor U3470 (N_3470,N_845,N_2383);
nand U3471 (N_3471,N_1920,N_313);
and U3472 (N_3472,N_662,N_1956);
xnor U3473 (N_3473,N_96,N_1437);
nand U3474 (N_3474,N_2420,N_2234);
nand U3475 (N_3475,N_144,N_1482);
nor U3476 (N_3476,N_2469,N_1054);
and U3477 (N_3477,N_2057,N_1636);
and U3478 (N_3478,N_882,N_1027);
nor U3479 (N_3479,N_2334,N_282);
xor U3480 (N_3480,N_2196,N_461);
and U3481 (N_3481,N_693,N_820);
nand U3482 (N_3482,N_737,N_1030);
nor U3483 (N_3483,N_1362,N_2169);
and U3484 (N_3484,N_285,N_219);
or U3485 (N_3485,N_1210,N_1651);
nand U3486 (N_3486,N_1878,N_605);
nor U3487 (N_3487,N_2226,N_550);
nand U3488 (N_3488,N_1198,N_984);
nand U3489 (N_3489,N_1851,N_818);
nand U3490 (N_3490,N_1295,N_885);
nor U3491 (N_3491,N_1114,N_2447);
xnor U3492 (N_3492,N_1232,N_973);
nor U3493 (N_3493,N_670,N_1745);
and U3494 (N_3494,N_1848,N_963);
nor U3495 (N_3495,N_1363,N_2325);
nor U3496 (N_3496,N_1614,N_812);
and U3497 (N_3497,N_581,N_547);
or U3498 (N_3498,N_1110,N_621);
nand U3499 (N_3499,N_1404,N_827);
nand U3500 (N_3500,N_2043,N_1311);
and U3501 (N_3501,N_801,N_988);
or U3502 (N_3502,N_230,N_992);
and U3503 (N_3503,N_1074,N_1580);
nand U3504 (N_3504,N_2068,N_49);
or U3505 (N_3505,N_2280,N_1542);
or U3506 (N_3506,N_1476,N_2296);
and U3507 (N_3507,N_1812,N_1674);
and U3508 (N_3508,N_1121,N_1900);
or U3509 (N_3509,N_1035,N_1414);
nand U3510 (N_3510,N_231,N_2086);
nor U3511 (N_3511,N_1616,N_2076);
or U3512 (N_3512,N_2010,N_1357);
or U3513 (N_3513,N_2458,N_1185);
or U3514 (N_3514,N_2453,N_2421);
and U3515 (N_3515,N_1714,N_1175);
nand U3516 (N_3516,N_2365,N_329);
nor U3517 (N_3517,N_1525,N_1815);
and U3518 (N_3518,N_176,N_1112);
xor U3519 (N_3519,N_795,N_924);
or U3520 (N_3520,N_1762,N_1855);
and U3521 (N_3521,N_2041,N_234);
and U3522 (N_3522,N_450,N_761);
nor U3523 (N_3523,N_504,N_1484);
nor U3524 (N_3524,N_417,N_340);
nor U3525 (N_3525,N_986,N_2203);
or U3526 (N_3526,N_773,N_1434);
or U3527 (N_3527,N_2373,N_1252);
and U3528 (N_3528,N_2319,N_405);
and U3529 (N_3529,N_1853,N_1544);
and U3530 (N_3530,N_1555,N_1336);
nor U3531 (N_3531,N_1978,N_2054);
nor U3532 (N_3532,N_1008,N_232);
and U3533 (N_3533,N_2393,N_2252);
nand U3534 (N_3534,N_887,N_18);
xor U3535 (N_3535,N_711,N_1799);
or U3536 (N_3536,N_218,N_791);
nor U3537 (N_3537,N_708,N_527);
nor U3538 (N_3538,N_591,N_237);
or U3539 (N_3539,N_437,N_690);
and U3540 (N_3540,N_1793,N_1543);
and U3541 (N_3541,N_456,N_413);
nor U3542 (N_3542,N_1663,N_1285);
and U3543 (N_3543,N_1846,N_1964);
nand U3544 (N_3544,N_48,N_968);
nand U3545 (N_3545,N_1521,N_1672);
and U3546 (N_3546,N_2369,N_257);
and U3547 (N_3547,N_817,N_426);
nor U3548 (N_3548,N_2300,N_1313);
nand U3549 (N_3549,N_1537,N_332);
and U3550 (N_3550,N_1640,N_583);
nor U3551 (N_3551,N_2395,N_683);
xor U3552 (N_3552,N_1303,N_2477);
and U3553 (N_3553,N_380,N_1592);
or U3554 (N_3554,N_502,N_1170);
and U3555 (N_3555,N_952,N_1591);
or U3556 (N_3556,N_895,N_2390);
or U3557 (N_3557,N_2495,N_1919);
or U3558 (N_3558,N_944,N_2051);
nand U3559 (N_3559,N_1319,N_1785);
or U3560 (N_3560,N_799,N_1238);
and U3561 (N_3561,N_510,N_56);
nor U3562 (N_3562,N_570,N_16);
or U3563 (N_3563,N_1620,N_2357);
nor U3564 (N_3564,N_580,N_2481);
nor U3565 (N_3565,N_665,N_624);
and U3566 (N_3566,N_186,N_1561);
nand U3567 (N_3567,N_1837,N_876);
or U3568 (N_3568,N_2229,N_2142);
nor U3569 (N_3569,N_374,N_1284);
xnor U3570 (N_3570,N_2096,N_838);
and U3571 (N_3571,N_2358,N_2192);
nor U3572 (N_3572,N_1083,N_533);
nand U3573 (N_3573,N_1998,N_2042);
nor U3574 (N_3574,N_55,N_1000);
nand U3575 (N_3575,N_781,N_1321);
nand U3576 (N_3576,N_1487,N_1536);
nor U3577 (N_3577,N_523,N_705);
and U3578 (N_3578,N_2097,N_2130);
nor U3579 (N_3579,N_1041,N_79);
or U3580 (N_3580,N_1702,N_2144);
nand U3581 (N_3581,N_1802,N_1996);
or U3582 (N_3582,N_765,N_1911);
nand U3583 (N_3583,N_2078,N_1222);
nand U3584 (N_3584,N_193,N_315);
and U3585 (N_3585,N_2329,N_531);
or U3586 (N_3586,N_2015,N_500);
or U3587 (N_3587,N_1585,N_519);
nor U3588 (N_3588,N_805,N_2175);
or U3589 (N_3589,N_1426,N_253);
and U3590 (N_3590,N_1378,N_364);
and U3591 (N_3591,N_2276,N_1217);
nor U3592 (N_3592,N_1305,N_645);
and U3593 (N_3593,N_2058,N_226);
or U3594 (N_3594,N_768,N_1047);
xnor U3595 (N_3595,N_1042,N_476);
and U3596 (N_3596,N_1412,N_472);
or U3597 (N_3597,N_1808,N_1940);
nor U3598 (N_3598,N_793,N_1573);
nor U3599 (N_3599,N_1186,N_804);
nand U3600 (N_3600,N_1863,N_122);
nor U3601 (N_3601,N_41,N_225);
and U3602 (N_3602,N_792,N_1398);
nand U3603 (N_3603,N_1287,N_2402);
or U3604 (N_3604,N_242,N_185);
nor U3605 (N_3605,N_587,N_785);
nand U3606 (N_3606,N_1915,N_1720);
nand U3607 (N_3607,N_1828,N_672);
and U3608 (N_3608,N_1282,N_2353);
or U3609 (N_3609,N_734,N_1916);
nor U3610 (N_3610,N_1060,N_1790);
nand U3611 (N_3611,N_1715,N_2311);
nand U3612 (N_3612,N_163,N_2450);
or U3613 (N_3613,N_24,N_2026);
nand U3614 (N_3614,N_2006,N_2345);
and U3615 (N_3615,N_2129,N_1501);
nand U3616 (N_3616,N_1691,N_1477);
nand U3617 (N_3617,N_1387,N_1124);
nand U3618 (N_3618,N_847,N_1432);
nand U3619 (N_3619,N_1939,N_125);
nand U3620 (N_3620,N_912,N_1522);
nor U3621 (N_3621,N_994,N_2388);
nand U3622 (N_3622,N_981,N_2064);
or U3623 (N_3623,N_625,N_839);
nand U3624 (N_3624,N_860,N_2088);
nor U3625 (N_3625,N_1360,N_2350);
or U3626 (N_3626,N_666,N_1386);
and U3627 (N_3627,N_643,N_1025);
nand U3628 (N_3628,N_2163,N_1741);
nor U3629 (N_3629,N_1923,N_101);
and U3630 (N_3630,N_1463,N_1681);
and U3631 (N_3631,N_50,N_1989);
or U3632 (N_3632,N_579,N_1727);
xnor U3633 (N_3633,N_25,N_713);
or U3634 (N_3634,N_850,N_1649);
nor U3635 (N_3635,N_368,N_1469);
and U3636 (N_3636,N_2290,N_337);
xnor U3637 (N_3637,N_1335,N_267);
and U3638 (N_3638,N_1523,N_2081);
nor U3639 (N_3639,N_746,N_678);
and U3640 (N_3640,N_1736,N_58);
nand U3641 (N_3641,N_1113,N_1910);
nor U3642 (N_3642,N_1297,N_2254);
and U3643 (N_3643,N_439,N_1535);
and U3644 (N_3644,N_600,N_2331);
and U3645 (N_3645,N_97,N_1128);
nand U3646 (N_3646,N_2490,N_1975);
nand U3647 (N_3647,N_2044,N_1732);
nand U3648 (N_3648,N_2354,N_1152);
or U3649 (N_3649,N_108,N_2067);
or U3650 (N_3650,N_1274,N_575);
nand U3651 (N_3651,N_429,N_308);
nor U3652 (N_3652,N_2181,N_883);
nand U3653 (N_3653,N_1676,N_68);
or U3654 (N_3654,N_1670,N_911);
and U3655 (N_3655,N_567,N_39);
or U3656 (N_3656,N_452,N_150);
nor U3657 (N_3657,N_1262,N_2225);
xnor U3658 (N_3658,N_1950,N_772);
or U3659 (N_3659,N_2012,N_2492);
or U3660 (N_3660,N_983,N_1307);
and U3661 (N_3661,N_494,N_999);
and U3662 (N_3662,N_1530,N_819);
or U3663 (N_3663,N_348,N_1221);
nor U3664 (N_3664,N_848,N_2128);
and U3665 (N_3665,N_520,N_1669);
and U3666 (N_3666,N_2164,N_2245);
nand U3667 (N_3667,N_1043,N_1704);
or U3668 (N_3668,N_391,N_1236);
or U3669 (N_3669,N_2467,N_69);
nor U3670 (N_3670,N_699,N_2349);
and U3671 (N_3671,N_796,N_1700);
and U3672 (N_3672,N_1553,N_1713);
nand U3673 (N_3673,N_433,N_577);
and U3674 (N_3674,N_2439,N_1588);
nor U3675 (N_3675,N_1751,N_211);
or U3676 (N_3676,N_1662,N_1597);
xnor U3677 (N_3677,N_2017,N_2285);
and U3678 (N_3678,N_2330,N_1937);
nand U3679 (N_3679,N_837,N_208);
and U3680 (N_3680,N_903,N_1467);
and U3681 (N_3681,N_2303,N_967);
or U3682 (N_3682,N_57,N_548);
or U3683 (N_3683,N_401,N_1554);
and U3684 (N_3684,N_2223,N_351);
nor U3685 (N_3685,N_457,N_94);
or U3686 (N_3686,N_962,N_1600);
nor U3687 (N_3687,N_1733,N_319);
nor U3688 (N_3688,N_1310,N_691);
nor U3689 (N_3689,N_2132,N_435);
nand U3690 (N_3690,N_264,N_1180);
xor U3691 (N_3691,N_1611,N_606);
or U3692 (N_3692,N_1999,N_2177);
nand U3693 (N_3693,N_2153,N_1641);
or U3694 (N_3694,N_210,N_1379);
nor U3695 (N_3695,N_1678,N_1529);
or U3696 (N_3696,N_658,N_809);
nor U3697 (N_3697,N_1717,N_965);
nand U3698 (N_3698,N_274,N_1729);
and U3699 (N_3699,N_2380,N_2405);
or U3700 (N_3700,N_1961,N_1959);
or U3701 (N_3701,N_752,N_534);
nand U3702 (N_3702,N_195,N_545);
nor U3703 (N_3703,N_249,N_1777);
nor U3704 (N_3704,N_298,N_239);
nor U3705 (N_3705,N_1036,N_2335);
nand U3706 (N_3706,N_762,N_454);
and U3707 (N_3707,N_1496,N_1189);
nor U3708 (N_3708,N_1826,N_1538);
or U3709 (N_3709,N_103,N_1129);
or U3710 (N_3710,N_1280,N_1675);
nand U3711 (N_3711,N_1560,N_777);
and U3712 (N_3712,N_1963,N_1290);
or U3713 (N_3713,N_2404,N_685);
nor U3714 (N_3714,N_1667,N_1022);
or U3715 (N_3715,N_1829,N_1957);
nor U3716 (N_3716,N_1408,N_1163);
xor U3717 (N_3717,N_2441,N_1721);
or U3718 (N_3718,N_909,N_1242);
nand U3719 (N_3719,N_1823,N_1511);
nor U3720 (N_3720,N_2204,N_2443);
and U3721 (N_3721,N_1351,N_686);
or U3722 (N_3722,N_1774,N_904);
nand U3723 (N_3723,N_1612,N_2205);
and U3724 (N_3724,N_732,N_1064);
nand U3725 (N_3725,N_1034,N_154);
nand U3726 (N_3726,N_1601,N_1317);
nor U3727 (N_3727,N_2227,N_1737);
nor U3728 (N_3728,N_442,N_813);
and U3729 (N_3729,N_894,N_1472);
nor U3730 (N_3730,N_1417,N_1626);
and U3731 (N_3731,N_404,N_187);
nor U3732 (N_3732,N_1639,N_1071);
or U3733 (N_3733,N_396,N_2366);
or U3734 (N_3734,N_2117,N_1101);
nand U3735 (N_3735,N_1277,N_15);
nand U3736 (N_3736,N_856,N_739);
and U3737 (N_3737,N_1570,N_916);
or U3738 (N_3738,N_174,N_595);
nand U3739 (N_3739,N_1869,N_2185);
nand U3740 (N_3740,N_1811,N_1126);
or U3741 (N_3741,N_2327,N_1973);
nand U3742 (N_3742,N_1480,N_1090);
nand U3743 (N_3743,N_1435,N_1299);
or U3744 (N_3744,N_1023,N_1231);
or U3745 (N_3745,N_406,N_2297);
nor U3746 (N_3746,N_2414,N_829);
nor U3747 (N_3747,N_1738,N_1865);
nor U3748 (N_3748,N_82,N_92);
and U3749 (N_3749,N_2023,N_1857);
nor U3750 (N_3750,N_907,N_1457);
and U3751 (N_3751,N_2073,N_1996);
or U3752 (N_3752,N_1434,N_2439);
and U3753 (N_3753,N_2435,N_173);
or U3754 (N_3754,N_1200,N_2388);
and U3755 (N_3755,N_2386,N_848);
or U3756 (N_3756,N_1594,N_1569);
and U3757 (N_3757,N_2460,N_2256);
and U3758 (N_3758,N_1872,N_588);
nor U3759 (N_3759,N_1321,N_2035);
and U3760 (N_3760,N_962,N_2262);
nor U3761 (N_3761,N_125,N_1757);
nand U3762 (N_3762,N_1618,N_1580);
and U3763 (N_3763,N_1866,N_1874);
and U3764 (N_3764,N_905,N_1159);
or U3765 (N_3765,N_1281,N_2411);
and U3766 (N_3766,N_2276,N_143);
nand U3767 (N_3767,N_2352,N_37);
and U3768 (N_3768,N_262,N_1363);
nand U3769 (N_3769,N_964,N_1984);
or U3770 (N_3770,N_2230,N_1660);
nand U3771 (N_3771,N_878,N_253);
or U3772 (N_3772,N_2410,N_120);
nand U3773 (N_3773,N_2084,N_1291);
nor U3774 (N_3774,N_560,N_2396);
nand U3775 (N_3775,N_260,N_2353);
and U3776 (N_3776,N_2045,N_514);
nor U3777 (N_3777,N_515,N_1469);
and U3778 (N_3778,N_1120,N_928);
or U3779 (N_3779,N_1162,N_751);
nand U3780 (N_3780,N_2427,N_1485);
nand U3781 (N_3781,N_1416,N_299);
or U3782 (N_3782,N_2210,N_582);
and U3783 (N_3783,N_1977,N_671);
nor U3784 (N_3784,N_2446,N_1739);
and U3785 (N_3785,N_2020,N_880);
nand U3786 (N_3786,N_911,N_685);
or U3787 (N_3787,N_2018,N_38);
nand U3788 (N_3788,N_150,N_22);
and U3789 (N_3789,N_114,N_1106);
and U3790 (N_3790,N_396,N_1909);
nor U3791 (N_3791,N_1471,N_781);
and U3792 (N_3792,N_267,N_388);
or U3793 (N_3793,N_2301,N_2079);
nand U3794 (N_3794,N_971,N_165);
nor U3795 (N_3795,N_2187,N_1538);
and U3796 (N_3796,N_553,N_787);
nand U3797 (N_3797,N_2159,N_1943);
or U3798 (N_3798,N_1426,N_670);
and U3799 (N_3799,N_151,N_1012);
or U3800 (N_3800,N_1943,N_1034);
or U3801 (N_3801,N_763,N_1337);
xor U3802 (N_3802,N_601,N_84);
or U3803 (N_3803,N_1908,N_1031);
nand U3804 (N_3804,N_196,N_1985);
nor U3805 (N_3805,N_2017,N_550);
or U3806 (N_3806,N_1008,N_2140);
or U3807 (N_3807,N_176,N_2274);
nand U3808 (N_3808,N_1658,N_2347);
nor U3809 (N_3809,N_1565,N_1908);
nand U3810 (N_3810,N_518,N_859);
nor U3811 (N_3811,N_2418,N_1048);
xor U3812 (N_3812,N_162,N_513);
nor U3813 (N_3813,N_1951,N_2136);
nand U3814 (N_3814,N_199,N_380);
xnor U3815 (N_3815,N_1003,N_645);
or U3816 (N_3816,N_2018,N_1671);
and U3817 (N_3817,N_41,N_689);
nand U3818 (N_3818,N_2077,N_758);
nand U3819 (N_3819,N_1620,N_2467);
nand U3820 (N_3820,N_1144,N_1611);
nor U3821 (N_3821,N_916,N_1648);
nor U3822 (N_3822,N_173,N_1465);
nor U3823 (N_3823,N_2285,N_748);
or U3824 (N_3824,N_2137,N_822);
or U3825 (N_3825,N_1949,N_2391);
and U3826 (N_3826,N_888,N_1275);
and U3827 (N_3827,N_842,N_1158);
or U3828 (N_3828,N_1819,N_993);
nor U3829 (N_3829,N_412,N_1313);
nor U3830 (N_3830,N_1028,N_141);
nand U3831 (N_3831,N_1455,N_421);
and U3832 (N_3832,N_1534,N_1864);
nand U3833 (N_3833,N_2121,N_180);
or U3834 (N_3834,N_725,N_124);
or U3835 (N_3835,N_1193,N_971);
nand U3836 (N_3836,N_842,N_554);
nor U3837 (N_3837,N_441,N_2000);
nand U3838 (N_3838,N_2144,N_596);
or U3839 (N_3839,N_1033,N_519);
nand U3840 (N_3840,N_1544,N_2218);
nand U3841 (N_3841,N_790,N_2176);
nand U3842 (N_3842,N_589,N_1026);
and U3843 (N_3843,N_2009,N_359);
nor U3844 (N_3844,N_2408,N_1722);
and U3845 (N_3845,N_350,N_1332);
nand U3846 (N_3846,N_122,N_1156);
and U3847 (N_3847,N_938,N_182);
nor U3848 (N_3848,N_962,N_1624);
or U3849 (N_3849,N_156,N_2225);
and U3850 (N_3850,N_599,N_1459);
or U3851 (N_3851,N_907,N_240);
nor U3852 (N_3852,N_677,N_1447);
nand U3853 (N_3853,N_873,N_1312);
and U3854 (N_3854,N_352,N_2225);
nand U3855 (N_3855,N_983,N_2219);
and U3856 (N_3856,N_1706,N_1932);
or U3857 (N_3857,N_2368,N_74);
and U3858 (N_3858,N_132,N_828);
or U3859 (N_3859,N_2488,N_2158);
nand U3860 (N_3860,N_2163,N_2202);
nand U3861 (N_3861,N_2362,N_101);
or U3862 (N_3862,N_2198,N_747);
nand U3863 (N_3863,N_1994,N_934);
or U3864 (N_3864,N_672,N_1024);
and U3865 (N_3865,N_1138,N_1174);
nand U3866 (N_3866,N_1471,N_2256);
or U3867 (N_3867,N_624,N_769);
nand U3868 (N_3868,N_767,N_509);
nor U3869 (N_3869,N_1236,N_1614);
nor U3870 (N_3870,N_232,N_1884);
and U3871 (N_3871,N_967,N_214);
or U3872 (N_3872,N_775,N_122);
nand U3873 (N_3873,N_2037,N_2032);
nor U3874 (N_3874,N_2341,N_2136);
and U3875 (N_3875,N_1267,N_2172);
or U3876 (N_3876,N_156,N_2240);
nand U3877 (N_3877,N_743,N_1681);
nand U3878 (N_3878,N_823,N_1514);
or U3879 (N_3879,N_1723,N_849);
and U3880 (N_3880,N_1158,N_364);
or U3881 (N_3881,N_27,N_569);
nand U3882 (N_3882,N_827,N_1278);
and U3883 (N_3883,N_1067,N_556);
and U3884 (N_3884,N_2407,N_235);
nand U3885 (N_3885,N_1570,N_2270);
and U3886 (N_3886,N_2088,N_2275);
nor U3887 (N_3887,N_2168,N_531);
nor U3888 (N_3888,N_473,N_2006);
nor U3889 (N_3889,N_1124,N_1279);
and U3890 (N_3890,N_146,N_1144);
nand U3891 (N_3891,N_703,N_1984);
nand U3892 (N_3892,N_1014,N_43);
nor U3893 (N_3893,N_1243,N_2090);
nand U3894 (N_3894,N_1058,N_897);
and U3895 (N_3895,N_831,N_2004);
nor U3896 (N_3896,N_198,N_284);
or U3897 (N_3897,N_211,N_139);
and U3898 (N_3898,N_1230,N_748);
and U3899 (N_3899,N_592,N_778);
and U3900 (N_3900,N_2032,N_1067);
nand U3901 (N_3901,N_1071,N_1169);
and U3902 (N_3902,N_561,N_321);
and U3903 (N_3903,N_2450,N_522);
nand U3904 (N_3904,N_2292,N_77);
nand U3905 (N_3905,N_1725,N_2378);
and U3906 (N_3906,N_1251,N_2320);
or U3907 (N_3907,N_2180,N_940);
nor U3908 (N_3908,N_1024,N_1327);
nor U3909 (N_3909,N_1704,N_980);
and U3910 (N_3910,N_1439,N_1114);
and U3911 (N_3911,N_1042,N_1928);
nand U3912 (N_3912,N_940,N_221);
and U3913 (N_3913,N_2143,N_1090);
nor U3914 (N_3914,N_474,N_1105);
or U3915 (N_3915,N_124,N_2193);
nor U3916 (N_3916,N_1978,N_2330);
or U3917 (N_3917,N_1964,N_1808);
nor U3918 (N_3918,N_446,N_1092);
and U3919 (N_3919,N_335,N_2209);
or U3920 (N_3920,N_47,N_642);
nor U3921 (N_3921,N_1347,N_2049);
or U3922 (N_3922,N_1606,N_1699);
and U3923 (N_3923,N_2479,N_292);
or U3924 (N_3924,N_598,N_876);
and U3925 (N_3925,N_1311,N_131);
or U3926 (N_3926,N_1168,N_463);
nor U3927 (N_3927,N_1550,N_1893);
nor U3928 (N_3928,N_1923,N_851);
nand U3929 (N_3929,N_267,N_1323);
xnor U3930 (N_3930,N_1632,N_1833);
or U3931 (N_3931,N_895,N_2017);
nand U3932 (N_3932,N_386,N_2490);
nand U3933 (N_3933,N_954,N_2084);
nand U3934 (N_3934,N_1256,N_296);
nand U3935 (N_3935,N_1892,N_1047);
or U3936 (N_3936,N_448,N_1366);
nor U3937 (N_3937,N_107,N_1397);
nand U3938 (N_3938,N_1105,N_2205);
nor U3939 (N_3939,N_2359,N_881);
and U3940 (N_3940,N_1634,N_1222);
and U3941 (N_3941,N_1931,N_805);
nand U3942 (N_3942,N_1130,N_1373);
nor U3943 (N_3943,N_2148,N_1728);
nand U3944 (N_3944,N_220,N_2134);
nand U3945 (N_3945,N_670,N_42);
or U3946 (N_3946,N_1824,N_879);
or U3947 (N_3947,N_1501,N_737);
nand U3948 (N_3948,N_1837,N_858);
nor U3949 (N_3949,N_1025,N_1893);
nand U3950 (N_3950,N_2347,N_1413);
and U3951 (N_3951,N_1040,N_2193);
nand U3952 (N_3952,N_2291,N_739);
and U3953 (N_3953,N_39,N_1944);
nor U3954 (N_3954,N_1310,N_542);
or U3955 (N_3955,N_354,N_2065);
xor U3956 (N_3956,N_138,N_126);
and U3957 (N_3957,N_2110,N_1191);
or U3958 (N_3958,N_719,N_2481);
xor U3959 (N_3959,N_419,N_1482);
or U3960 (N_3960,N_100,N_1910);
nand U3961 (N_3961,N_535,N_285);
nor U3962 (N_3962,N_1840,N_2399);
or U3963 (N_3963,N_1882,N_381);
and U3964 (N_3964,N_2021,N_950);
nor U3965 (N_3965,N_1473,N_1335);
and U3966 (N_3966,N_694,N_639);
nand U3967 (N_3967,N_67,N_2038);
or U3968 (N_3968,N_1194,N_1936);
nand U3969 (N_3969,N_347,N_2488);
or U3970 (N_3970,N_163,N_1475);
nor U3971 (N_3971,N_998,N_770);
nor U3972 (N_3972,N_1145,N_767);
and U3973 (N_3973,N_2145,N_951);
or U3974 (N_3974,N_1228,N_2387);
or U3975 (N_3975,N_810,N_2241);
nor U3976 (N_3976,N_2056,N_771);
and U3977 (N_3977,N_2181,N_101);
nand U3978 (N_3978,N_490,N_2326);
nor U3979 (N_3979,N_884,N_1146);
nor U3980 (N_3980,N_437,N_612);
nor U3981 (N_3981,N_774,N_423);
nand U3982 (N_3982,N_1368,N_1491);
or U3983 (N_3983,N_1810,N_266);
and U3984 (N_3984,N_2158,N_404);
nand U3985 (N_3985,N_766,N_1948);
or U3986 (N_3986,N_2256,N_2315);
and U3987 (N_3987,N_554,N_524);
or U3988 (N_3988,N_2406,N_229);
or U3989 (N_3989,N_813,N_2177);
nand U3990 (N_3990,N_904,N_837);
nand U3991 (N_3991,N_1849,N_2125);
or U3992 (N_3992,N_154,N_396);
or U3993 (N_3993,N_852,N_743);
nor U3994 (N_3994,N_1007,N_1941);
and U3995 (N_3995,N_2043,N_1137);
and U3996 (N_3996,N_1278,N_1818);
or U3997 (N_3997,N_801,N_2079);
and U3998 (N_3998,N_715,N_2379);
or U3999 (N_3999,N_941,N_230);
nor U4000 (N_4000,N_729,N_1046);
nor U4001 (N_4001,N_558,N_2381);
nor U4002 (N_4002,N_1066,N_532);
nor U4003 (N_4003,N_1,N_1586);
nor U4004 (N_4004,N_2167,N_150);
and U4005 (N_4005,N_1492,N_1854);
and U4006 (N_4006,N_1292,N_1036);
or U4007 (N_4007,N_813,N_2424);
nor U4008 (N_4008,N_1029,N_890);
nand U4009 (N_4009,N_2108,N_1454);
nor U4010 (N_4010,N_576,N_331);
nand U4011 (N_4011,N_157,N_691);
nand U4012 (N_4012,N_2482,N_476);
and U4013 (N_4013,N_71,N_481);
nand U4014 (N_4014,N_2454,N_1613);
or U4015 (N_4015,N_568,N_1473);
and U4016 (N_4016,N_1968,N_1959);
nand U4017 (N_4017,N_1539,N_1055);
and U4018 (N_4018,N_2250,N_209);
nor U4019 (N_4019,N_2361,N_800);
or U4020 (N_4020,N_774,N_1693);
or U4021 (N_4021,N_1632,N_299);
nor U4022 (N_4022,N_1159,N_7);
or U4023 (N_4023,N_2059,N_772);
nor U4024 (N_4024,N_1345,N_2039);
or U4025 (N_4025,N_2377,N_894);
nor U4026 (N_4026,N_2114,N_1983);
nand U4027 (N_4027,N_2335,N_1388);
and U4028 (N_4028,N_607,N_638);
nand U4029 (N_4029,N_1199,N_1941);
nor U4030 (N_4030,N_812,N_846);
and U4031 (N_4031,N_1014,N_824);
and U4032 (N_4032,N_513,N_540);
or U4033 (N_4033,N_1527,N_1811);
or U4034 (N_4034,N_1228,N_945);
or U4035 (N_4035,N_2219,N_659);
and U4036 (N_4036,N_1052,N_1992);
nand U4037 (N_4037,N_689,N_1831);
or U4038 (N_4038,N_262,N_1486);
nor U4039 (N_4039,N_1630,N_1348);
and U4040 (N_4040,N_162,N_461);
nand U4041 (N_4041,N_2334,N_1456);
and U4042 (N_4042,N_2353,N_2483);
and U4043 (N_4043,N_2179,N_1315);
nand U4044 (N_4044,N_1180,N_734);
and U4045 (N_4045,N_2429,N_1342);
nand U4046 (N_4046,N_735,N_1343);
nor U4047 (N_4047,N_185,N_1265);
nor U4048 (N_4048,N_900,N_1314);
nand U4049 (N_4049,N_9,N_2254);
xnor U4050 (N_4050,N_420,N_571);
nand U4051 (N_4051,N_76,N_1978);
nor U4052 (N_4052,N_1149,N_1919);
or U4053 (N_4053,N_1009,N_336);
nand U4054 (N_4054,N_1958,N_1886);
or U4055 (N_4055,N_40,N_2165);
nand U4056 (N_4056,N_1191,N_2381);
or U4057 (N_4057,N_1081,N_1914);
nor U4058 (N_4058,N_763,N_2075);
and U4059 (N_4059,N_1809,N_1186);
and U4060 (N_4060,N_2438,N_1224);
nor U4061 (N_4061,N_1848,N_891);
or U4062 (N_4062,N_1475,N_153);
nor U4063 (N_4063,N_260,N_1221);
or U4064 (N_4064,N_392,N_1104);
nor U4065 (N_4065,N_1856,N_1398);
or U4066 (N_4066,N_1768,N_1120);
nor U4067 (N_4067,N_1371,N_1642);
or U4068 (N_4068,N_2205,N_1213);
nor U4069 (N_4069,N_644,N_1912);
and U4070 (N_4070,N_333,N_1221);
and U4071 (N_4071,N_1820,N_1340);
nor U4072 (N_4072,N_2226,N_378);
nand U4073 (N_4073,N_570,N_1900);
or U4074 (N_4074,N_2475,N_741);
and U4075 (N_4075,N_1612,N_2363);
nand U4076 (N_4076,N_744,N_112);
and U4077 (N_4077,N_1363,N_2219);
nor U4078 (N_4078,N_1839,N_2311);
and U4079 (N_4079,N_1470,N_2045);
and U4080 (N_4080,N_1330,N_828);
nor U4081 (N_4081,N_822,N_1967);
and U4082 (N_4082,N_2342,N_277);
nand U4083 (N_4083,N_1724,N_1071);
and U4084 (N_4084,N_971,N_1497);
or U4085 (N_4085,N_1529,N_195);
or U4086 (N_4086,N_2243,N_1736);
xor U4087 (N_4087,N_305,N_596);
nor U4088 (N_4088,N_2173,N_1170);
or U4089 (N_4089,N_1772,N_1727);
and U4090 (N_4090,N_189,N_1531);
and U4091 (N_4091,N_576,N_1949);
nand U4092 (N_4092,N_231,N_2448);
and U4093 (N_4093,N_1152,N_589);
nand U4094 (N_4094,N_1582,N_473);
and U4095 (N_4095,N_374,N_1950);
nor U4096 (N_4096,N_2460,N_2110);
xnor U4097 (N_4097,N_1841,N_3);
nor U4098 (N_4098,N_1,N_2356);
and U4099 (N_4099,N_1021,N_925);
or U4100 (N_4100,N_859,N_2207);
nor U4101 (N_4101,N_1165,N_1103);
and U4102 (N_4102,N_1956,N_1381);
and U4103 (N_4103,N_245,N_2301);
nand U4104 (N_4104,N_2124,N_1312);
nor U4105 (N_4105,N_1215,N_2345);
or U4106 (N_4106,N_39,N_2400);
nand U4107 (N_4107,N_2086,N_968);
and U4108 (N_4108,N_1379,N_1067);
nand U4109 (N_4109,N_1232,N_1539);
and U4110 (N_4110,N_313,N_2240);
and U4111 (N_4111,N_1718,N_422);
or U4112 (N_4112,N_2139,N_1487);
and U4113 (N_4113,N_741,N_1527);
or U4114 (N_4114,N_1172,N_1241);
and U4115 (N_4115,N_441,N_1507);
and U4116 (N_4116,N_2025,N_54);
nand U4117 (N_4117,N_1438,N_512);
or U4118 (N_4118,N_2328,N_773);
nor U4119 (N_4119,N_52,N_1869);
nor U4120 (N_4120,N_86,N_1761);
and U4121 (N_4121,N_856,N_304);
or U4122 (N_4122,N_1038,N_1902);
nand U4123 (N_4123,N_741,N_1858);
xnor U4124 (N_4124,N_1999,N_1133);
and U4125 (N_4125,N_2061,N_843);
nand U4126 (N_4126,N_3,N_2250);
and U4127 (N_4127,N_773,N_2474);
or U4128 (N_4128,N_164,N_763);
and U4129 (N_4129,N_2009,N_455);
or U4130 (N_4130,N_562,N_1153);
nor U4131 (N_4131,N_218,N_1240);
and U4132 (N_4132,N_601,N_400);
and U4133 (N_4133,N_1498,N_834);
nor U4134 (N_4134,N_1857,N_2353);
nand U4135 (N_4135,N_2015,N_1229);
nor U4136 (N_4136,N_520,N_77);
nor U4137 (N_4137,N_1041,N_226);
and U4138 (N_4138,N_906,N_1410);
nor U4139 (N_4139,N_2054,N_646);
nor U4140 (N_4140,N_1416,N_981);
nor U4141 (N_4141,N_173,N_1883);
nor U4142 (N_4142,N_2187,N_506);
and U4143 (N_4143,N_2260,N_916);
nor U4144 (N_4144,N_2260,N_1155);
nand U4145 (N_4145,N_962,N_1573);
and U4146 (N_4146,N_1370,N_1471);
and U4147 (N_4147,N_1234,N_2395);
nand U4148 (N_4148,N_676,N_775);
and U4149 (N_4149,N_2163,N_289);
nand U4150 (N_4150,N_1029,N_407);
nor U4151 (N_4151,N_1179,N_2019);
nor U4152 (N_4152,N_838,N_2478);
nand U4153 (N_4153,N_1190,N_396);
nand U4154 (N_4154,N_1720,N_142);
or U4155 (N_4155,N_1649,N_518);
and U4156 (N_4156,N_2332,N_566);
nand U4157 (N_4157,N_2002,N_1498);
nor U4158 (N_4158,N_1145,N_462);
and U4159 (N_4159,N_2136,N_357);
nor U4160 (N_4160,N_1156,N_1859);
xnor U4161 (N_4161,N_710,N_1244);
nor U4162 (N_4162,N_1521,N_1575);
and U4163 (N_4163,N_900,N_2493);
or U4164 (N_4164,N_1081,N_288);
nor U4165 (N_4165,N_626,N_2035);
and U4166 (N_4166,N_1441,N_739);
or U4167 (N_4167,N_2259,N_1795);
nor U4168 (N_4168,N_1891,N_2048);
nand U4169 (N_4169,N_1054,N_1971);
nand U4170 (N_4170,N_1965,N_1978);
nand U4171 (N_4171,N_1634,N_498);
or U4172 (N_4172,N_1342,N_1397);
nor U4173 (N_4173,N_1185,N_1866);
nor U4174 (N_4174,N_2059,N_1870);
nor U4175 (N_4175,N_2475,N_2429);
or U4176 (N_4176,N_1190,N_2277);
nand U4177 (N_4177,N_1275,N_477);
nand U4178 (N_4178,N_1701,N_1652);
or U4179 (N_4179,N_1726,N_590);
and U4180 (N_4180,N_2413,N_1960);
and U4181 (N_4181,N_264,N_1039);
and U4182 (N_4182,N_1325,N_1602);
or U4183 (N_4183,N_12,N_1364);
nor U4184 (N_4184,N_312,N_1824);
nand U4185 (N_4185,N_129,N_1560);
nand U4186 (N_4186,N_1787,N_1369);
and U4187 (N_4187,N_516,N_374);
nor U4188 (N_4188,N_461,N_1330);
and U4189 (N_4189,N_2163,N_742);
nand U4190 (N_4190,N_40,N_1879);
and U4191 (N_4191,N_1885,N_2026);
nor U4192 (N_4192,N_583,N_918);
nor U4193 (N_4193,N_2086,N_416);
nor U4194 (N_4194,N_241,N_583);
and U4195 (N_4195,N_2341,N_118);
nor U4196 (N_4196,N_289,N_1974);
xor U4197 (N_4197,N_638,N_632);
xnor U4198 (N_4198,N_1649,N_969);
and U4199 (N_4199,N_2207,N_674);
nand U4200 (N_4200,N_106,N_1413);
and U4201 (N_4201,N_455,N_301);
nand U4202 (N_4202,N_1872,N_14);
or U4203 (N_4203,N_868,N_335);
nand U4204 (N_4204,N_1604,N_1765);
or U4205 (N_4205,N_1328,N_2170);
or U4206 (N_4206,N_48,N_174);
or U4207 (N_4207,N_2361,N_2303);
nand U4208 (N_4208,N_575,N_1210);
and U4209 (N_4209,N_1203,N_1552);
and U4210 (N_4210,N_1803,N_2421);
or U4211 (N_4211,N_2083,N_1396);
nor U4212 (N_4212,N_2386,N_1788);
nand U4213 (N_4213,N_418,N_212);
or U4214 (N_4214,N_556,N_2421);
nor U4215 (N_4215,N_525,N_1522);
and U4216 (N_4216,N_742,N_2261);
nand U4217 (N_4217,N_112,N_313);
nand U4218 (N_4218,N_768,N_598);
nor U4219 (N_4219,N_2,N_691);
nor U4220 (N_4220,N_793,N_1955);
xnor U4221 (N_4221,N_2252,N_2218);
and U4222 (N_4222,N_1585,N_96);
or U4223 (N_4223,N_163,N_24);
nor U4224 (N_4224,N_2309,N_438);
and U4225 (N_4225,N_468,N_1139);
nor U4226 (N_4226,N_393,N_44);
nor U4227 (N_4227,N_2134,N_787);
nand U4228 (N_4228,N_2475,N_2086);
nand U4229 (N_4229,N_1851,N_1454);
nor U4230 (N_4230,N_2436,N_1277);
nor U4231 (N_4231,N_542,N_1153);
xor U4232 (N_4232,N_502,N_1081);
nand U4233 (N_4233,N_580,N_1957);
or U4234 (N_4234,N_306,N_1740);
and U4235 (N_4235,N_1925,N_468);
or U4236 (N_4236,N_422,N_1914);
nand U4237 (N_4237,N_631,N_2204);
or U4238 (N_4238,N_1722,N_1464);
nor U4239 (N_4239,N_1013,N_1901);
nor U4240 (N_4240,N_2196,N_2188);
or U4241 (N_4241,N_210,N_401);
nor U4242 (N_4242,N_2397,N_980);
xnor U4243 (N_4243,N_586,N_729);
and U4244 (N_4244,N_2358,N_1061);
nand U4245 (N_4245,N_931,N_887);
or U4246 (N_4246,N_283,N_1791);
or U4247 (N_4247,N_2021,N_1780);
and U4248 (N_4248,N_608,N_1660);
or U4249 (N_4249,N_2425,N_1118);
and U4250 (N_4250,N_2355,N_1381);
and U4251 (N_4251,N_1269,N_1968);
and U4252 (N_4252,N_1656,N_1337);
nor U4253 (N_4253,N_1519,N_1366);
nor U4254 (N_4254,N_1376,N_1270);
nor U4255 (N_4255,N_1089,N_988);
or U4256 (N_4256,N_2176,N_1689);
or U4257 (N_4257,N_1440,N_1334);
nor U4258 (N_4258,N_2206,N_1046);
nand U4259 (N_4259,N_836,N_471);
nor U4260 (N_4260,N_1692,N_935);
nor U4261 (N_4261,N_1021,N_1037);
xnor U4262 (N_4262,N_1632,N_703);
and U4263 (N_4263,N_2065,N_1870);
and U4264 (N_4264,N_375,N_784);
nor U4265 (N_4265,N_2371,N_1137);
nand U4266 (N_4266,N_1726,N_2059);
nor U4267 (N_4267,N_149,N_337);
nor U4268 (N_4268,N_2134,N_908);
nand U4269 (N_4269,N_2165,N_1847);
nor U4270 (N_4270,N_1302,N_1666);
nor U4271 (N_4271,N_2173,N_1449);
and U4272 (N_4272,N_783,N_631);
nand U4273 (N_4273,N_535,N_1690);
and U4274 (N_4274,N_994,N_1333);
or U4275 (N_4275,N_1572,N_140);
and U4276 (N_4276,N_1623,N_1014);
and U4277 (N_4277,N_1785,N_11);
and U4278 (N_4278,N_507,N_832);
nor U4279 (N_4279,N_2186,N_80);
nand U4280 (N_4280,N_836,N_1788);
nor U4281 (N_4281,N_641,N_1462);
and U4282 (N_4282,N_1667,N_965);
nand U4283 (N_4283,N_1080,N_178);
and U4284 (N_4284,N_809,N_1383);
nor U4285 (N_4285,N_773,N_849);
nor U4286 (N_4286,N_19,N_1530);
and U4287 (N_4287,N_704,N_1872);
or U4288 (N_4288,N_170,N_280);
nor U4289 (N_4289,N_1535,N_978);
nor U4290 (N_4290,N_2345,N_2290);
nor U4291 (N_4291,N_2177,N_1249);
nor U4292 (N_4292,N_286,N_2489);
nand U4293 (N_4293,N_2136,N_938);
nor U4294 (N_4294,N_2321,N_1606);
nand U4295 (N_4295,N_2325,N_1898);
nand U4296 (N_4296,N_1110,N_1015);
or U4297 (N_4297,N_2430,N_2446);
xnor U4298 (N_4298,N_1663,N_898);
and U4299 (N_4299,N_1093,N_1773);
nand U4300 (N_4300,N_2002,N_1469);
or U4301 (N_4301,N_452,N_1491);
or U4302 (N_4302,N_1641,N_1046);
nor U4303 (N_4303,N_908,N_983);
nand U4304 (N_4304,N_1033,N_6);
or U4305 (N_4305,N_1745,N_2381);
or U4306 (N_4306,N_2061,N_1430);
nand U4307 (N_4307,N_1153,N_719);
or U4308 (N_4308,N_1239,N_287);
nor U4309 (N_4309,N_1894,N_1665);
or U4310 (N_4310,N_2416,N_215);
nand U4311 (N_4311,N_1781,N_953);
or U4312 (N_4312,N_2243,N_1045);
nand U4313 (N_4313,N_497,N_1842);
nand U4314 (N_4314,N_1038,N_230);
or U4315 (N_4315,N_2330,N_108);
nand U4316 (N_4316,N_313,N_1712);
or U4317 (N_4317,N_421,N_358);
or U4318 (N_4318,N_35,N_1724);
nor U4319 (N_4319,N_663,N_1967);
nor U4320 (N_4320,N_1351,N_544);
nand U4321 (N_4321,N_1027,N_847);
and U4322 (N_4322,N_705,N_1240);
and U4323 (N_4323,N_937,N_2022);
nand U4324 (N_4324,N_2352,N_1072);
nor U4325 (N_4325,N_553,N_2313);
nor U4326 (N_4326,N_2220,N_1958);
nor U4327 (N_4327,N_38,N_1268);
nor U4328 (N_4328,N_1103,N_2215);
or U4329 (N_4329,N_206,N_1075);
nand U4330 (N_4330,N_1418,N_547);
and U4331 (N_4331,N_585,N_882);
or U4332 (N_4332,N_1910,N_2318);
or U4333 (N_4333,N_958,N_2351);
nand U4334 (N_4334,N_1226,N_1023);
and U4335 (N_4335,N_1787,N_1537);
nor U4336 (N_4336,N_428,N_379);
nor U4337 (N_4337,N_265,N_133);
and U4338 (N_4338,N_2001,N_733);
nor U4339 (N_4339,N_386,N_822);
or U4340 (N_4340,N_490,N_1874);
and U4341 (N_4341,N_335,N_2078);
nor U4342 (N_4342,N_687,N_1525);
and U4343 (N_4343,N_1024,N_2288);
nor U4344 (N_4344,N_2057,N_325);
nor U4345 (N_4345,N_1376,N_1698);
nor U4346 (N_4346,N_342,N_136);
nand U4347 (N_4347,N_2188,N_1098);
nor U4348 (N_4348,N_64,N_765);
and U4349 (N_4349,N_560,N_953);
nor U4350 (N_4350,N_468,N_1869);
and U4351 (N_4351,N_1995,N_19);
and U4352 (N_4352,N_392,N_14);
and U4353 (N_4353,N_671,N_1691);
nand U4354 (N_4354,N_1855,N_25);
or U4355 (N_4355,N_487,N_666);
and U4356 (N_4356,N_1713,N_1158);
nand U4357 (N_4357,N_1319,N_2254);
or U4358 (N_4358,N_2487,N_2073);
nor U4359 (N_4359,N_1087,N_673);
nand U4360 (N_4360,N_243,N_1201);
nor U4361 (N_4361,N_1200,N_772);
or U4362 (N_4362,N_2031,N_2157);
and U4363 (N_4363,N_503,N_2115);
nor U4364 (N_4364,N_1876,N_587);
nand U4365 (N_4365,N_463,N_1444);
and U4366 (N_4366,N_531,N_1654);
nor U4367 (N_4367,N_2301,N_1098);
nand U4368 (N_4368,N_482,N_966);
nand U4369 (N_4369,N_1863,N_194);
and U4370 (N_4370,N_1534,N_2165);
nor U4371 (N_4371,N_1625,N_445);
nor U4372 (N_4372,N_922,N_1357);
nand U4373 (N_4373,N_839,N_2205);
and U4374 (N_4374,N_1414,N_1031);
nand U4375 (N_4375,N_1378,N_1725);
and U4376 (N_4376,N_2399,N_1627);
and U4377 (N_4377,N_1849,N_459);
or U4378 (N_4378,N_577,N_2260);
nor U4379 (N_4379,N_2355,N_1632);
nand U4380 (N_4380,N_147,N_1368);
and U4381 (N_4381,N_723,N_1121);
and U4382 (N_4382,N_2097,N_1169);
nor U4383 (N_4383,N_1459,N_865);
nand U4384 (N_4384,N_516,N_243);
or U4385 (N_4385,N_1270,N_784);
or U4386 (N_4386,N_892,N_2064);
and U4387 (N_4387,N_2030,N_1014);
nand U4388 (N_4388,N_2226,N_1909);
nor U4389 (N_4389,N_145,N_1589);
nor U4390 (N_4390,N_1517,N_1070);
nor U4391 (N_4391,N_2460,N_2085);
or U4392 (N_4392,N_1707,N_276);
nor U4393 (N_4393,N_1832,N_886);
xor U4394 (N_4394,N_2072,N_1264);
or U4395 (N_4395,N_632,N_1464);
or U4396 (N_4396,N_1407,N_1922);
nor U4397 (N_4397,N_2330,N_2020);
and U4398 (N_4398,N_1309,N_435);
nor U4399 (N_4399,N_2167,N_966);
or U4400 (N_4400,N_497,N_1423);
nor U4401 (N_4401,N_599,N_368);
nor U4402 (N_4402,N_1022,N_940);
nor U4403 (N_4403,N_2454,N_820);
or U4404 (N_4404,N_1271,N_2301);
xor U4405 (N_4405,N_1421,N_1217);
and U4406 (N_4406,N_2275,N_1465);
or U4407 (N_4407,N_1117,N_272);
or U4408 (N_4408,N_2337,N_1634);
nor U4409 (N_4409,N_2237,N_563);
nor U4410 (N_4410,N_2359,N_2449);
nor U4411 (N_4411,N_1519,N_1797);
or U4412 (N_4412,N_1974,N_1185);
nand U4413 (N_4413,N_1788,N_296);
nor U4414 (N_4414,N_150,N_1517);
or U4415 (N_4415,N_2441,N_635);
or U4416 (N_4416,N_1615,N_1228);
nand U4417 (N_4417,N_1436,N_1233);
or U4418 (N_4418,N_1893,N_1156);
nand U4419 (N_4419,N_944,N_1320);
nand U4420 (N_4420,N_354,N_1479);
or U4421 (N_4421,N_2449,N_2006);
and U4422 (N_4422,N_366,N_1734);
nor U4423 (N_4423,N_183,N_198);
nand U4424 (N_4424,N_987,N_1520);
nand U4425 (N_4425,N_2257,N_1217);
nor U4426 (N_4426,N_502,N_1208);
nand U4427 (N_4427,N_1665,N_2113);
or U4428 (N_4428,N_644,N_297);
or U4429 (N_4429,N_2061,N_1535);
nand U4430 (N_4430,N_622,N_891);
nand U4431 (N_4431,N_1175,N_1853);
or U4432 (N_4432,N_2023,N_1963);
nand U4433 (N_4433,N_1709,N_1828);
nand U4434 (N_4434,N_2338,N_520);
nor U4435 (N_4435,N_1906,N_2411);
or U4436 (N_4436,N_697,N_104);
and U4437 (N_4437,N_495,N_327);
nand U4438 (N_4438,N_2053,N_2216);
and U4439 (N_4439,N_2435,N_1724);
nor U4440 (N_4440,N_2125,N_1832);
nor U4441 (N_4441,N_980,N_2159);
and U4442 (N_4442,N_1857,N_2386);
nor U4443 (N_4443,N_1278,N_939);
nor U4444 (N_4444,N_1134,N_1975);
nand U4445 (N_4445,N_2174,N_331);
or U4446 (N_4446,N_161,N_2097);
and U4447 (N_4447,N_214,N_1426);
nand U4448 (N_4448,N_1944,N_481);
or U4449 (N_4449,N_2052,N_58);
or U4450 (N_4450,N_247,N_507);
or U4451 (N_4451,N_1450,N_646);
nor U4452 (N_4452,N_2455,N_1186);
nor U4453 (N_4453,N_1783,N_1627);
or U4454 (N_4454,N_1247,N_981);
and U4455 (N_4455,N_608,N_2094);
or U4456 (N_4456,N_1383,N_2495);
and U4457 (N_4457,N_919,N_357);
xor U4458 (N_4458,N_1134,N_309);
nor U4459 (N_4459,N_1560,N_2106);
nand U4460 (N_4460,N_891,N_1613);
and U4461 (N_4461,N_404,N_508);
and U4462 (N_4462,N_553,N_1604);
nand U4463 (N_4463,N_299,N_312);
nor U4464 (N_4464,N_706,N_1844);
and U4465 (N_4465,N_1422,N_1327);
nor U4466 (N_4466,N_841,N_1085);
nand U4467 (N_4467,N_242,N_359);
and U4468 (N_4468,N_912,N_953);
nor U4469 (N_4469,N_378,N_584);
and U4470 (N_4470,N_97,N_2207);
nand U4471 (N_4471,N_1844,N_221);
nor U4472 (N_4472,N_183,N_2114);
and U4473 (N_4473,N_2380,N_911);
and U4474 (N_4474,N_1323,N_1636);
nand U4475 (N_4475,N_1820,N_991);
or U4476 (N_4476,N_348,N_448);
or U4477 (N_4477,N_1377,N_937);
or U4478 (N_4478,N_1137,N_509);
nand U4479 (N_4479,N_21,N_466);
or U4480 (N_4480,N_601,N_336);
or U4481 (N_4481,N_286,N_1434);
nand U4482 (N_4482,N_1939,N_1185);
and U4483 (N_4483,N_432,N_2218);
and U4484 (N_4484,N_2134,N_1482);
and U4485 (N_4485,N_1390,N_1626);
nand U4486 (N_4486,N_1066,N_770);
nor U4487 (N_4487,N_2485,N_1997);
xnor U4488 (N_4488,N_599,N_1225);
nand U4489 (N_4489,N_613,N_232);
nor U4490 (N_4490,N_1568,N_2319);
nor U4491 (N_4491,N_293,N_521);
or U4492 (N_4492,N_2297,N_1363);
or U4493 (N_4493,N_455,N_113);
nand U4494 (N_4494,N_2381,N_732);
nor U4495 (N_4495,N_1228,N_1753);
and U4496 (N_4496,N_2389,N_1588);
and U4497 (N_4497,N_983,N_308);
nand U4498 (N_4498,N_13,N_545);
or U4499 (N_4499,N_1380,N_2063);
nand U4500 (N_4500,N_2380,N_1005);
nand U4501 (N_4501,N_1717,N_543);
or U4502 (N_4502,N_1071,N_995);
or U4503 (N_4503,N_333,N_953);
nor U4504 (N_4504,N_76,N_2278);
and U4505 (N_4505,N_955,N_1378);
and U4506 (N_4506,N_477,N_1709);
or U4507 (N_4507,N_901,N_2480);
nand U4508 (N_4508,N_2139,N_2336);
nand U4509 (N_4509,N_2499,N_1112);
and U4510 (N_4510,N_1240,N_954);
or U4511 (N_4511,N_2248,N_1627);
nor U4512 (N_4512,N_609,N_1187);
nor U4513 (N_4513,N_1184,N_642);
and U4514 (N_4514,N_964,N_119);
and U4515 (N_4515,N_1357,N_163);
nor U4516 (N_4516,N_1323,N_1324);
nor U4517 (N_4517,N_406,N_499);
nand U4518 (N_4518,N_829,N_1868);
nor U4519 (N_4519,N_989,N_1271);
and U4520 (N_4520,N_507,N_52);
and U4521 (N_4521,N_820,N_986);
or U4522 (N_4522,N_1865,N_5);
and U4523 (N_4523,N_122,N_1738);
nor U4524 (N_4524,N_706,N_1611);
or U4525 (N_4525,N_151,N_725);
or U4526 (N_4526,N_943,N_1561);
or U4527 (N_4527,N_1886,N_2298);
nand U4528 (N_4528,N_756,N_806);
and U4529 (N_4529,N_2350,N_912);
nand U4530 (N_4530,N_614,N_1681);
nand U4531 (N_4531,N_937,N_158);
and U4532 (N_4532,N_2332,N_1266);
or U4533 (N_4533,N_1620,N_2065);
nand U4534 (N_4534,N_23,N_594);
nor U4535 (N_4535,N_247,N_1551);
or U4536 (N_4536,N_2015,N_2243);
nand U4537 (N_4537,N_104,N_1565);
and U4538 (N_4538,N_2159,N_257);
or U4539 (N_4539,N_2241,N_2227);
nand U4540 (N_4540,N_1605,N_2450);
or U4541 (N_4541,N_2269,N_2188);
and U4542 (N_4542,N_800,N_754);
or U4543 (N_4543,N_683,N_490);
or U4544 (N_4544,N_977,N_1840);
and U4545 (N_4545,N_1185,N_1622);
nor U4546 (N_4546,N_1257,N_1919);
nor U4547 (N_4547,N_1425,N_2331);
nand U4548 (N_4548,N_2372,N_101);
or U4549 (N_4549,N_1363,N_656);
and U4550 (N_4550,N_682,N_97);
or U4551 (N_4551,N_794,N_1917);
and U4552 (N_4552,N_1323,N_1802);
nor U4553 (N_4553,N_1426,N_872);
nand U4554 (N_4554,N_1486,N_1071);
nand U4555 (N_4555,N_745,N_2302);
and U4556 (N_4556,N_1617,N_2298);
xnor U4557 (N_4557,N_1277,N_1014);
or U4558 (N_4558,N_2437,N_648);
and U4559 (N_4559,N_1082,N_1974);
and U4560 (N_4560,N_1753,N_1570);
or U4561 (N_4561,N_1157,N_1584);
or U4562 (N_4562,N_1321,N_1);
nor U4563 (N_4563,N_1294,N_2121);
and U4564 (N_4564,N_2451,N_326);
nor U4565 (N_4565,N_281,N_193);
nor U4566 (N_4566,N_1135,N_78);
and U4567 (N_4567,N_1550,N_894);
or U4568 (N_4568,N_1087,N_2330);
nand U4569 (N_4569,N_1725,N_800);
nor U4570 (N_4570,N_2313,N_1578);
and U4571 (N_4571,N_2080,N_1900);
nor U4572 (N_4572,N_506,N_2388);
or U4573 (N_4573,N_2384,N_350);
or U4574 (N_4574,N_2099,N_1576);
nand U4575 (N_4575,N_1506,N_2348);
or U4576 (N_4576,N_1485,N_1119);
xor U4577 (N_4577,N_402,N_683);
and U4578 (N_4578,N_994,N_2111);
and U4579 (N_4579,N_1540,N_1083);
or U4580 (N_4580,N_260,N_2082);
or U4581 (N_4581,N_122,N_1541);
nand U4582 (N_4582,N_1157,N_632);
nand U4583 (N_4583,N_931,N_1274);
and U4584 (N_4584,N_1112,N_721);
and U4585 (N_4585,N_82,N_718);
nand U4586 (N_4586,N_1657,N_1063);
nor U4587 (N_4587,N_2395,N_2219);
nor U4588 (N_4588,N_1990,N_2315);
and U4589 (N_4589,N_1624,N_366);
nor U4590 (N_4590,N_1868,N_808);
or U4591 (N_4591,N_893,N_2165);
and U4592 (N_4592,N_213,N_2463);
and U4593 (N_4593,N_455,N_2065);
and U4594 (N_4594,N_1851,N_2316);
nor U4595 (N_4595,N_1171,N_1385);
nor U4596 (N_4596,N_2181,N_2078);
and U4597 (N_4597,N_2442,N_1205);
nor U4598 (N_4598,N_1122,N_499);
or U4599 (N_4599,N_977,N_1530);
or U4600 (N_4600,N_59,N_1649);
and U4601 (N_4601,N_2114,N_167);
nand U4602 (N_4602,N_342,N_1415);
nand U4603 (N_4603,N_1015,N_1214);
nor U4604 (N_4604,N_331,N_387);
nand U4605 (N_4605,N_994,N_88);
or U4606 (N_4606,N_553,N_2472);
nor U4607 (N_4607,N_760,N_1368);
and U4608 (N_4608,N_1690,N_1936);
and U4609 (N_4609,N_584,N_1994);
or U4610 (N_4610,N_2398,N_418);
nor U4611 (N_4611,N_299,N_2403);
nand U4612 (N_4612,N_2243,N_944);
nor U4613 (N_4613,N_1225,N_719);
xor U4614 (N_4614,N_320,N_46);
or U4615 (N_4615,N_1317,N_881);
or U4616 (N_4616,N_2245,N_1239);
or U4617 (N_4617,N_1413,N_966);
and U4618 (N_4618,N_777,N_1290);
and U4619 (N_4619,N_1807,N_1980);
nor U4620 (N_4620,N_2204,N_1211);
or U4621 (N_4621,N_1023,N_516);
and U4622 (N_4622,N_2174,N_2007);
nand U4623 (N_4623,N_1082,N_886);
nor U4624 (N_4624,N_1870,N_2439);
and U4625 (N_4625,N_1614,N_872);
and U4626 (N_4626,N_2392,N_1213);
nor U4627 (N_4627,N_2240,N_2015);
nand U4628 (N_4628,N_1410,N_353);
nor U4629 (N_4629,N_1185,N_2397);
nor U4630 (N_4630,N_1822,N_1534);
nand U4631 (N_4631,N_2436,N_991);
or U4632 (N_4632,N_1964,N_1085);
or U4633 (N_4633,N_2288,N_1042);
nor U4634 (N_4634,N_884,N_2315);
nor U4635 (N_4635,N_1231,N_1735);
nand U4636 (N_4636,N_380,N_1088);
nand U4637 (N_4637,N_887,N_975);
nor U4638 (N_4638,N_2289,N_2337);
nor U4639 (N_4639,N_2499,N_2234);
nor U4640 (N_4640,N_2444,N_834);
nor U4641 (N_4641,N_1360,N_112);
or U4642 (N_4642,N_1668,N_861);
or U4643 (N_4643,N_1512,N_2162);
nand U4644 (N_4644,N_1105,N_213);
nand U4645 (N_4645,N_235,N_1344);
nor U4646 (N_4646,N_2367,N_1993);
nand U4647 (N_4647,N_1831,N_1148);
nand U4648 (N_4648,N_1050,N_1268);
and U4649 (N_4649,N_79,N_2490);
and U4650 (N_4650,N_1904,N_2229);
nor U4651 (N_4651,N_1110,N_762);
or U4652 (N_4652,N_2155,N_1563);
nand U4653 (N_4653,N_816,N_1316);
or U4654 (N_4654,N_1891,N_2098);
or U4655 (N_4655,N_272,N_1625);
nand U4656 (N_4656,N_1000,N_1894);
or U4657 (N_4657,N_1058,N_539);
and U4658 (N_4658,N_2439,N_268);
nor U4659 (N_4659,N_1554,N_130);
nor U4660 (N_4660,N_163,N_1448);
nor U4661 (N_4661,N_578,N_582);
nor U4662 (N_4662,N_2156,N_831);
or U4663 (N_4663,N_839,N_1776);
or U4664 (N_4664,N_1965,N_1775);
nor U4665 (N_4665,N_793,N_1245);
or U4666 (N_4666,N_111,N_2000);
or U4667 (N_4667,N_1279,N_2407);
nor U4668 (N_4668,N_1102,N_114);
nand U4669 (N_4669,N_708,N_1022);
nand U4670 (N_4670,N_744,N_1275);
and U4671 (N_4671,N_298,N_2482);
nand U4672 (N_4672,N_2120,N_1515);
and U4673 (N_4673,N_2332,N_1704);
nand U4674 (N_4674,N_2279,N_280);
nand U4675 (N_4675,N_1553,N_2297);
nand U4676 (N_4676,N_134,N_78);
nor U4677 (N_4677,N_1833,N_126);
or U4678 (N_4678,N_2072,N_1087);
nor U4679 (N_4679,N_1160,N_233);
nor U4680 (N_4680,N_853,N_956);
nor U4681 (N_4681,N_2046,N_1858);
or U4682 (N_4682,N_1875,N_1770);
nand U4683 (N_4683,N_534,N_2182);
nand U4684 (N_4684,N_1924,N_1711);
nand U4685 (N_4685,N_1573,N_1127);
nor U4686 (N_4686,N_1497,N_42);
nand U4687 (N_4687,N_1698,N_320);
xnor U4688 (N_4688,N_1018,N_2407);
nor U4689 (N_4689,N_699,N_1994);
or U4690 (N_4690,N_845,N_2102);
nand U4691 (N_4691,N_1304,N_1333);
or U4692 (N_4692,N_1464,N_678);
nor U4693 (N_4693,N_506,N_1085);
or U4694 (N_4694,N_636,N_112);
nor U4695 (N_4695,N_1724,N_885);
nand U4696 (N_4696,N_1290,N_1984);
nor U4697 (N_4697,N_1972,N_417);
or U4698 (N_4698,N_1765,N_665);
or U4699 (N_4699,N_1836,N_2307);
nor U4700 (N_4700,N_2108,N_2361);
or U4701 (N_4701,N_1644,N_972);
and U4702 (N_4702,N_2487,N_1151);
and U4703 (N_4703,N_1012,N_1546);
and U4704 (N_4704,N_1436,N_1296);
or U4705 (N_4705,N_316,N_1437);
and U4706 (N_4706,N_1615,N_1139);
nand U4707 (N_4707,N_1762,N_1220);
and U4708 (N_4708,N_1686,N_557);
nor U4709 (N_4709,N_478,N_982);
and U4710 (N_4710,N_2334,N_1604);
or U4711 (N_4711,N_1527,N_383);
nor U4712 (N_4712,N_581,N_1315);
and U4713 (N_4713,N_1260,N_2144);
nand U4714 (N_4714,N_1699,N_722);
nor U4715 (N_4715,N_761,N_623);
nor U4716 (N_4716,N_887,N_2250);
nand U4717 (N_4717,N_239,N_1391);
or U4718 (N_4718,N_1396,N_2117);
nor U4719 (N_4719,N_535,N_1433);
or U4720 (N_4720,N_2299,N_151);
or U4721 (N_4721,N_2471,N_1859);
and U4722 (N_4722,N_519,N_1726);
nor U4723 (N_4723,N_1598,N_1412);
nor U4724 (N_4724,N_2203,N_952);
nor U4725 (N_4725,N_1113,N_751);
nand U4726 (N_4726,N_349,N_1859);
or U4727 (N_4727,N_2489,N_150);
or U4728 (N_4728,N_2135,N_110);
and U4729 (N_4729,N_735,N_1554);
nor U4730 (N_4730,N_918,N_1415);
and U4731 (N_4731,N_513,N_904);
nand U4732 (N_4732,N_1922,N_1877);
nand U4733 (N_4733,N_97,N_1570);
nand U4734 (N_4734,N_2374,N_1805);
nand U4735 (N_4735,N_1616,N_2089);
or U4736 (N_4736,N_1230,N_482);
nand U4737 (N_4737,N_181,N_548);
or U4738 (N_4738,N_1873,N_898);
or U4739 (N_4739,N_639,N_1656);
nand U4740 (N_4740,N_2370,N_655);
nor U4741 (N_4741,N_248,N_782);
or U4742 (N_4742,N_1218,N_66);
xnor U4743 (N_4743,N_441,N_0);
or U4744 (N_4744,N_965,N_1217);
and U4745 (N_4745,N_1599,N_113);
or U4746 (N_4746,N_993,N_1446);
nand U4747 (N_4747,N_1660,N_2432);
and U4748 (N_4748,N_1977,N_1988);
nand U4749 (N_4749,N_738,N_86);
nor U4750 (N_4750,N_1496,N_1727);
nand U4751 (N_4751,N_1699,N_1506);
or U4752 (N_4752,N_1693,N_2246);
and U4753 (N_4753,N_1403,N_811);
nand U4754 (N_4754,N_468,N_2312);
nor U4755 (N_4755,N_695,N_2143);
or U4756 (N_4756,N_1317,N_1427);
and U4757 (N_4757,N_870,N_2284);
nand U4758 (N_4758,N_16,N_2311);
nand U4759 (N_4759,N_1242,N_1659);
nand U4760 (N_4760,N_595,N_1005);
xor U4761 (N_4761,N_1936,N_1814);
nand U4762 (N_4762,N_699,N_1064);
and U4763 (N_4763,N_2206,N_568);
or U4764 (N_4764,N_1690,N_1131);
nor U4765 (N_4765,N_1336,N_492);
nand U4766 (N_4766,N_1934,N_642);
or U4767 (N_4767,N_891,N_1275);
nand U4768 (N_4768,N_76,N_2094);
or U4769 (N_4769,N_979,N_2318);
and U4770 (N_4770,N_368,N_2448);
and U4771 (N_4771,N_2266,N_139);
xor U4772 (N_4772,N_1005,N_928);
or U4773 (N_4773,N_1258,N_664);
or U4774 (N_4774,N_1644,N_910);
nor U4775 (N_4775,N_2208,N_1447);
and U4776 (N_4776,N_3,N_706);
and U4777 (N_4777,N_1166,N_10);
or U4778 (N_4778,N_1232,N_2440);
nand U4779 (N_4779,N_1278,N_1299);
or U4780 (N_4780,N_1957,N_1732);
and U4781 (N_4781,N_1328,N_1831);
or U4782 (N_4782,N_1471,N_1691);
nor U4783 (N_4783,N_2307,N_663);
nor U4784 (N_4784,N_446,N_160);
or U4785 (N_4785,N_1057,N_2148);
and U4786 (N_4786,N_1801,N_2476);
xor U4787 (N_4787,N_691,N_2110);
and U4788 (N_4788,N_1842,N_422);
or U4789 (N_4789,N_1399,N_2151);
and U4790 (N_4790,N_1215,N_617);
and U4791 (N_4791,N_1947,N_1719);
nand U4792 (N_4792,N_1216,N_2491);
and U4793 (N_4793,N_1846,N_2192);
or U4794 (N_4794,N_1926,N_41);
and U4795 (N_4795,N_1104,N_330);
nand U4796 (N_4796,N_1782,N_1501);
or U4797 (N_4797,N_2057,N_1591);
and U4798 (N_4798,N_1200,N_2211);
and U4799 (N_4799,N_1814,N_2449);
nor U4800 (N_4800,N_1393,N_1919);
or U4801 (N_4801,N_1909,N_601);
nor U4802 (N_4802,N_1258,N_265);
nand U4803 (N_4803,N_604,N_2422);
and U4804 (N_4804,N_2268,N_2419);
and U4805 (N_4805,N_42,N_919);
or U4806 (N_4806,N_1498,N_1838);
or U4807 (N_4807,N_1252,N_2442);
and U4808 (N_4808,N_426,N_2023);
nand U4809 (N_4809,N_1444,N_2443);
or U4810 (N_4810,N_115,N_262);
xor U4811 (N_4811,N_296,N_499);
nor U4812 (N_4812,N_1557,N_694);
nand U4813 (N_4813,N_170,N_2358);
nand U4814 (N_4814,N_214,N_632);
or U4815 (N_4815,N_764,N_611);
nor U4816 (N_4816,N_347,N_2220);
nand U4817 (N_4817,N_956,N_1781);
and U4818 (N_4818,N_572,N_1496);
and U4819 (N_4819,N_927,N_1752);
nand U4820 (N_4820,N_1838,N_1943);
and U4821 (N_4821,N_1848,N_299);
or U4822 (N_4822,N_725,N_1253);
nor U4823 (N_4823,N_282,N_1533);
and U4824 (N_4824,N_605,N_981);
nand U4825 (N_4825,N_1726,N_279);
and U4826 (N_4826,N_1914,N_380);
xor U4827 (N_4827,N_107,N_513);
and U4828 (N_4828,N_1146,N_230);
and U4829 (N_4829,N_2005,N_2319);
or U4830 (N_4830,N_1245,N_867);
or U4831 (N_4831,N_2098,N_511);
and U4832 (N_4832,N_1269,N_1346);
or U4833 (N_4833,N_1542,N_1749);
and U4834 (N_4834,N_838,N_1614);
or U4835 (N_4835,N_1506,N_1598);
and U4836 (N_4836,N_1381,N_1160);
nand U4837 (N_4837,N_1735,N_1034);
nand U4838 (N_4838,N_540,N_829);
and U4839 (N_4839,N_369,N_1687);
nor U4840 (N_4840,N_2491,N_1702);
nor U4841 (N_4841,N_1729,N_1646);
and U4842 (N_4842,N_1357,N_744);
nand U4843 (N_4843,N_1827,N_1925);
nand U4844 (N_4844,N_2091,N_1146);
or U4845 (N_4845,N_200,N_703);
nand U4846 (N_4846,N_793,N_1414);
nand U4847 (N_4847,N_488,N_246);
nor U4848 (N_4848,N_1134,N_920);
nor U4849 (N_4849,N_1693,N_1163);
nor U4850 (N_4850,N_1266,N_2305);
nor U4851 (N_4851,N_2338,N_2202);
or U4852 (N_4852,N_906,N_1031);
and U4853 (N_4853,N_1203,N_2336);
nor U4854 (N_4854,N_2013,N_1020);
and U4855 (N_4855,N_1901,N_2231);
nand U4856 (N_4856,N_2229,N_2002);
and U4857 (N_4857,N_844,N_300);
or U4858 (N_4858,N_1528,N_1198);
nor U4859 (N_4859,N_907,N_1085);
nand U4860 (N_4860,N_1937,N_836);
or U4861 (N_4861,N_886,N_1546);
xor U4862 (N_4862,N_2109,N_525);
nand U4863 (N_4863,N_1015,N_262);
or U4864 (N_4864,N_852,N_1532);
nand U4865 (N_4865,N_588,N_1655);
nand U4866 (N_4866,N_1514,N_479);
nor U4867 (N_4867,N_1813,N_2057);
or U4868 (N_4868,N_1245,N_771);
nor U4869 (N_4869,N_1410,N_812);
nor U4870 (N_4870,N_1632,N_2123);
nand U4871 (N_4871,N_2253,N_1822);
and U4872 (N_4872,N_1661,N_1403);
nor U4873 (N_4873,N_1225,N_1487);
or U4874 (N_4874,N_2423,N_168);
or U4875 (N_4875,N_1029,N_148);
nand U4876 (N_4876,N_1182,N_2387);
nand U4877 (N_4877,N_629,N_1000);
and U4878 (N_4878,N_1590,N_1011);
and U4879 (N_4879,N_216,N_804);
nand U4880 (N_4880,N_879,N_1499);
nor U4881 (N_4881,N_2157,N_1937);
or U4882 (N_4882,N_1291,N_1494);
or U4883 (N_4883,N_163,N_1786);
nand U4884 (N_4884,N_1930,N_1929);
and U4885 (N_4885,N_276,N_905);
or U4886 (N_4886,N_26,N_2030);
or U4887 (N_4887,N_720,N_378);
nor U4888 (N_4888,N_926,N_1607);
nand U4889 (N_4889,N_1588,N_2412);
or U4890 (N_4890,N_2097,N_20);
nand U4891 (N_4891,N_2043,N_1979);
and U4892 (N_4892,N_2190,N_1150);
nand U4893 (N_4893,N_1201,N_1938);
nand U4894 (N_4894,N_2184,N_785);
or U4895 (N_4895,N_363,N_2390);
nand U4896 (N_4896,N_1187,N_1940);
or U4897 (N_4897,N_1094,N_1109);
nor U4898 (N_4898,N_929,N_1726);
nor U4899 (N_4899,N_711,N_2038);
or U4900 (N_4900,N_986,N_879);
and U4901 (N_4901,N_1798,N_1344);
nand U4902 (N_4902,N_1837,N_2079);
or U4903 (N_4903,N_419,N_173);
and U4904 (N_4904,N_1037,N_12);
or U4905 (N_4905,N_1736,N_257);
or U4906 (N_4906,N_1268,N_197);
nor U4907 (N_4907,N_205,N_841);
nand U4908 (N_4908,N_577,N_590);
nor U4909 (N_4909,N_921,N_1791);
nand U4910 (N_4910,N_1603,N_1692);
and U4911 (N_4911,N_460,N_510);
nor U4912 (N_4912,N_838,N_1670);
or U4913 (N_4913,N_1895,N_72);
or U4914 (N_4914,N_1916,N_2248);
and U4915 (N_4915,N_1829,N_1208);
nand U4916 (N_4916,N_784,N_1448);
nor U4917 (N_4917,N_1839,N_2316);
and U4918 (N_4918,N_1617,N_288);
or U4919 (N_4919,N_359,N_26);
nor U4920 (N_4920,N_2042,N_449);
nor U4921 (N_4921,N_673,N_1173);
nand U4922 (N_4922,N_1159,N_144);
or U4923 (N_4923,N_1494,N_802);
nor U4924 (N_4924,N_89,N_407);
nand U4925 (N_4925,N_1063,N_659);
nand U4926 (N_4926,N_1397,N_46);
or U4927 (N_4927,N_1552,N_1668);
nand U4928 (N_4928,N_1265,N_895);
or U4929 (N_4929,N_596,N_144);
nand U4930 (N_4930,N_772,N_2487);
or U4931 (N_4931,N_1824,N_1080);
and U4932 (N_4932,N_1476,N_279);
and U4933 (N_4933,N_931,N_401);
nand U4934 (N_4934,N_745,N_287);
nand U4935 (N_4935,N_801,N_2362);
or U4936 (N_4936,N_1044,N_2035);
and U4937 (N_4937,N_1225,N_289);
and U4938 (N_4938,N_2404,N_1800);
nor U4939 (N_4939,N_2292,N_553);
and U4940 (N_4940,N_725,N_969);
nand U4941 (N_4941,N_1163,N_493);
xor U4942 (N_4942,N_341,N_609);
nor U4943 (N_4943,N_771,N_2288);
or U4944 (N_4944,N_2121,N_356);
nor U4945 (N_4945,N_2423,N_1506);
and U4946 (N_4946,N_1007,N_1153);
and U4947 (N_4947,N_365,N_1647);
nor U4948 (N_4948,N_1730,N_2036);
or U4949 (N_4949,N_1216,N_1813);
nand U4950 (N_4950,N_712,N_1989);
nor U4951 (N_4951,N_276,N_2463);
nor U4952 (N_4952,N_2438,N_134);
nor U4953 (N_4953,N_640,N_16);
and U4954 (N_4954,N_1560,N_1158);
or U4955 (N_4955,N_4,N_1293);
nor U4956 (N_4956,N_968,N_1132);
xor U4957 (N_4957,N_175,N_920);
nand U4958 (N_4958,N_1915,N_1769);
or U4959 (N_4959,N_424,N_2252);
or U4960 (N_4960,N_1368,N_1211);
nand U4961 (N_4961,N_1804,N_2265);
or U4962 (N_4962,N_263,N_206);
or U4963 (N_4963,N_393,N_179);
and U4964 (N_4964,N_1007,N_1479);
or U4965 (N_4965,N_267,N_389);
and U4966 (N_4966,N_1883,N_756);
nand U4967 (N_4967,N_2099,N_2165);
or U4968 (N_4968,N_1838,N_1861);
or U4969 (N_4969,N_184,N_1763);
nor U4970 (N_4970,N_1066,N_549);
nand U4971 (N_4971,N_1557,N_1531);
and U4972 (N_4972,N_88,N_1455);
or U4973 (N_4973,N_2125,N_1340);
nand U4974 (N_4974,N_2208,N_558);
and U4975 (N_4975,N_168,N_1211);
nand U4976 (N_4976,N_2037,N_1058);
nand U4977 (N_4977,N_1695,N_2005);
and U4978 (N_4978,N_1021,N_771);
nor U4979 (N_4979,N_1491,N_2018);
and U4980 (N_4980,N_2379,N_1266);
nand U4981 (N_4981,N_869,N_694);
xor U4982 (N_4982,N_2158,N_1407);
nor U4983 (N_4983,N_597,N_1305);
nand U4984 (N_4984,N_1668,N_58);
or U4985 (N_4985,N_1475,N_1643);
and U4986 (N_4986,N_2440,N_1787);
nand U4987 (N_4987,N_105,N_262);
and U4988 (N_4988,N_2377,N_731);
or U4989 (N_4989,N_7,N_2126);
nor U4990 (N_4990,N_2460,N_2334);
and U4991 (N_4991,N_2043,N_1596);
and U4992 (N_4992,N_1541,N_1106);
and U4993 (N_4993,N_2465,N_1222);
and U4994 (N_4994,N_1574,N_1191);
xnor U4995 (N_4995,N_991,N_1142);
nor U4996 (N_4996,N_1649,N_362);
nor U4997 (N_4997,N_70,N_1746);
or U4998 (N_4998,N_2099,N_1766);
and U4999 (N_4999,N_2227,N_1495);
nand U5000 (N_5000,N_2678,N_3308);
nand U5001 (N_5001,N_2582,N_4532);
or U5002 (N_5002,N_2908,N_2619);
nor U5003 (N_5003,N_3105,N_4584);
and U5004 (N_5004,N_3736,N_2841);
nor U5005 (N_5005,N_2725,N_4766);
and U5006 (N_5006,N_3184,N_4399);
nor U5007 (N_5007,N_3616,N_3435);
nand U5008 (N_5008,N_4717,N_4329);
nor U5009 (N_5009,N_4923,N_3710);
nor U5010 (N_5010,N_4088,N_2903);
and U5011 (N_5011,N_2805,N_4758);
nor U5012 (N_5012,N_3844,N_4554);
and U5013 (N_5013,N_3699,N_4103);
nand U5014 (N_5014,N_4223,N_4209);
nand U5015 (N_5015,N_3356,N_4507);
and U5016 (N_5016,N_4574,N_4370);
or U5017 (N_5017,N_2770,N_3144);
and U5018 (N_5018,N_2694,N_3695);
and U5019 (N_5019,N_3962,N_4215);
or U5020 (N_5020,N_3499,N_4233);
nand U5021 (N_5021,N_2729,N_2552);
nor U5022 (N_5022,N_3168,N_4345);
nor U5023 (N_5023,N_4426,N_4855);
nor U5024 (N_5024,N_2917,N_3574);
nor U5025 (N_5025,N_4489,N_3653);
or U5026 (N_5026,N_3452,N_3246);
nand U5027 (N_5027,N_4889,N_4334);
xor U5028 (N_5028,N_3069,N_4149);
or U5029 (N_5029,N_4017,N_2786);
xor U5030 (N_5030,N_2751,N_4913);
nor U5031 (N_5031,N_4390,N_4304);
and U5032 (N_5032,N_4914,N_4236);
nor U5033 (N_5033,N_4364,N_3428);
nand U5034 (N_5034,N_3118,N_3276);
nand U5035 (N_5035,N_3421,N_2513);
nor U5036 (N_5036,N_3556,N_3854);
or U5037 (N_5037,N_4313,N_4521);
and U5038 (N_5038,N_4934,N_3601);
nor U5039 (N_5039,N_3117,N_4039);
or U5040 (N_5040,N_4277,N_3460);
and U5041 (N_5041,N_4371,N_2734);
nor U5042 (N_5042,N_2957,N_4721);
and U5043 (N_5043,N_4629,N_3002);
nor U5044 (N_5044,N_4533,N_4095);
nor U5045 (N_5045,N_3581,N_2809);
nand U5046 (N_5046,N_4021,N_3919);
or U5047 (N_5047,N_3289,N_4622);
nand U5048 (N_5048,N_2956,N_3973);
or U5049 (N_5049,N_3315,N_4705);
nand U5050 (N_5050,N_3891,N_4099);
nor U5051 (N_5051,N_4501,N_2715);
or U5052 (N_5052,N_2924,N_3610);
nor U5053 (N_5053,N_4094,N_4098);
and U5054 (N_5054,N_3388,N_3011);
and U5055 (N_5055,N_4443,N_2865);
nor U5056 (N_5056,N_2973,N_2521);
or U5057 (N_5057,N_2772,N_3974);
nor U5058 (N_5058,N_4548,N_2716);
xor U5059 (N_5059,N_3794,N_4949);
nand U5060 (N_5060,N_2664,N_3864);
or U5061 (N_5061,N_2667,N_3382);
nand U5062 (N_5062,N_2516,N_2897);
nand U5063 (N_5063,N_2847,N_4743);
nand U5064 (N_5064,N_3186,N_4177);
or U5065 (N_5065,N_3339,N_3155);
or U5066 (N_5066,N_4481,N_2609);
nor U5067 (N_5067,N_4248,N_4151);
or U5068 (N_5068,N_2870,N_4765);
and U5069 (N_5069,N_4627,N_4479);
and U5070 (N_5070,N_3153,N_4915);
nand U5071 (N_5071,N_4641,N_3991);
nand U5072 (N_5072,N_4247,N_3223);
nand U5073 (N_5073,N_2768,N_2835);
nand U5074 (N_5074,N_3612,N_2789);
and U5075 (N_5075,N_4956,N_2830);
xor U5076 (N_5076,N_3325,N_3907);
nor U5077 (N_5077,N_4222,N_2987);
nand U5078 (N_5078,N_3423,N_3625);
or U5079 (N_5079,N_2748,N_4587);
nor U5080 (N_5080,N_2673,N_4530);
or U5081 (N_5081,N_3116,N_4414);
nand U5082 (N_5082,N_4578,N_4971);
nand U5083 (N_5083,N_4969,N_2628);
nor U5084 (N_5084,N_3009,N_4990);
nand U5085 (N_5085,N_3783,N_2881);
nor U5086 (N_5086,N_3389,N_4272);
nor U5087 (N_5087,N_4073,N_3094);
and U5088 (N_5088,N_3501,N_4490);
nor U5089 (N_5089,N_2524,N_4219);
and U5090 (N_5090,N_3174,N_4702);
nor U5091 (N_5091,N_4729,N_4411);
nor U5092 (N_5092,N_4428,N_4275);
and U5093 (N_5093,N_2693,N_4077);
nand U5094 (N_5094,N_3990,N_4427);
and U5095 (N_5095,N_3750,N_2606);
xor U5096 (N_5096,N_2810,N_4875);
or U5097 (N_5097,N_2773,N_2629);
xnor U5098 (N_5098,N_3586,N_3860);
nor U5099 (N_5099,N_4645,N_3062);
nor U5100 (N_5100,N_2849,N_3534);
nand U5101 (N_5101,N_4857,N_4006);
and U5102 (N_5102,N_2544,N_4106);
nor U5103 (N_5103,N_3227,N_3291);
and U5104 (N_5104,N_4284,N_4071);
nand U5105 (N_5105,N_4305,N_3861);
and U5106 (N_5106,N_2802,N_4534);
or U5107 (N_5107,N_3050,N_3960);
nor U5108 (N_5108,N_3355,N_4356);
nor U5109 (N_5109,N_4461,N_4775);
or U5110 (N_5110,N_2819,N_3154);
and U5111 (N_5111,N_4323,N_4366);
nor U5112 (N_5112,N_3815,N_3141);
and U5113 (N_5113,N_4535,N_4303);
or U5114 (N_5114,N_3923,N_3606);
and U5115 (N_5115,N_3803,N_2696);
and U5116 (N_5116,N_4497,N_3835);
or U5117 (N_5117,N_4659,N_3784);
nand U5118 (N_5118,N_4415,N_3992);
or U5119 (N_5119,N_4599,N_4311);
nor U5120 (N_5120,N_4013,N_3211);
nor U5121 (N_5121,N_2576,N_2700);
xor U5122 (N_5122,N_2690,N_3497);
nor U5123 (N_5123,N_4592,N_2775);
nor U5124 (N_5124,N_2764,N_3218);
nand U5125 (N_5125,N_4817,N_3941);
nor U5126 (N_5126,N_4699,N_4435);
nand U5127 (N_5127,N_4315,N_2587);
or U5128 (N_5128,N_4877,N_2646);
nor U5129 (N_5129,N_2663,N_3214);
or U5130 (N_5130,N_4205,N_4518);
and U5131 (N_5131,N_4563,N_2867);
nand U5132 (N_5132,N_4101,N_4935);
nor U5133 (N_5133,N_2630,N_4963);
nor U5134 (N_5134,N_2602,N_4928);
or U5135 (N_5135,N_4774,N_3594);
and U5136 (N_5136,N_2793,N_3071);
nand U5137 (N_5137,N_3448,N_3839);
and U5138 (N_5138,N_4447,N_2566);
nor U5139 (N_5139,N_4450,N_3916);
and U5140 (N_5140,N_4338,N_2531);
or U5141 (N_5141,N_4035,N_3280);
nor U5142 (N_5142,N_4029,N_2861);
or U5143 (N_5143,N_4639,N_4108);
or U5144 (N_5144,N_3231,N_4133);
and U5145 (N_5145,N_2871,N_3019);
or U5146 (N_5146,N_4191,N_3819);
nand U5147 (N_5147,N_4217,N_2644);
nor U5148 (N_5148,N_2540,N_4084);
nand U5149 (N_5149,N_3731,N_4231);
nor U5150 (N_5150,N_4797,N_3171);
nand U5151 (N_5151,N_3929,N_2791);
and U5152 (N_5152,N_3544,N_3807);
or U5153 (N_5153,N_3471,N_3961);
and U5154 (N_5154,N_3446,N_3772);
nand U5155 (N_5155,N_4286,N_3309);
nor U5156 (N_5156,N_4686,N_3089);
nand U5157 (N_5157,N_2929,N_3052);
xor U5158 (N_5158,N_3818,N_4167);
nand U5159 (N_5159,N_4425,N_3351);
and U5160 (N_5160,N_4352,N_2741);
nor U5161 (N_5161,N_4328,N_3795);
nand U5162 (N_5162,N_4001,N_4912);
or U5163 (N_5163,N_3107,N_4493);
or U5164 (N_5164,N_4972,N_3102);
nand U5165 (N_5165,N_4747,N_3755);
nor U5166 (N_5166,N_4561,N_4092);
nand U5167 (N_5167,N_3965,N_3669);
nor U5168 (N_5168,N_2800,N_3734);
nor U5169 (N_5169,N_4666,N_4188);
nor U5170 (N_5170,N_2844,N_4250);
and U5171 (N_5171,N_3195,N_4351);
nor U5172 (N_5172,N_4009,N_4948);
and U5173 (N_5173,N_2633,N_4090);
nand U5174 (N_5174,N_4762,N_3593);
nand U5175 (N_5175,N_2889,N_2965);
nand U5176 (N_5176,N_2625,N_2549);
and U5177 (N_5177,N_3547,N_2899);
xnor U5178 (N_5178,N_4241,N_3233);
and U5179 (N_5179,N_4647,N_4033);
nand U5180 (N_5180,N_2616,N_4089);
nand U5181 (N_5181,N_3294,N_4121);
or U5182 (N_5182,N_3926,N_4291);
nor U5183 (N_5183,N_3337,N_4353);
nor U5184 (N_5184,N_3932,N_2698);
and U5185 (N_5185,N_4925,N_3904);
nor U5186 (N_5186,N_2780,N_4267);
and U5187 (N_5187,N_4322,N_4638);
nand U5188 (N_5188,N_3955,N_2938);
nand U5189 (N_5189,N_4945,N_3030);
or U5190 (N_5190,N_4940,N_4392);
nor U5191 (N_5191,N_3061,N_4036);
or U5192 (N_5192,N_2817,N_4342);
or U5193 (N_5193,N_2868,N_3433);
nor U5194 (N_5194,N_4330,N_3851);
nor U5195 (N_5195,N_4874,N_3346);
nor U5196 (N_5196,N_4410,N_3443);
or U5197 (N_5197,N_4871,N_3360);
nand U5198 (N_5198,N_3078,N_2506);
nand U5199 (N_5199,N_4876,N_4617);
or U5200 (N_5200,N_3559,N_3417);
and U5201 (N_5201,N_2683,N_3424);
or U5202 (N_5202,N_4238,N_3867);
or U5203 (N_5203,N_4244,N_4016);
nor U5204 (N_5204,N_4865,N_4879);
or U5205 (N_5205,N_2568,N_4448);
or U5206 (N_5206,N_3347,N_3311);
nand U5207 (N_5207,N_4727,N_4166);
and U5208 (N_5208,N_2922,N_2717);
or U5209 (N_5209,N_2508,N_4266);
nor U5210 (N_5210,N_3666,N_3158);
nor U5211 (N_5211,N_3997,N_3405);
nand U5212 (N_5212,N_4495,N_2901);
and U5213 (N_5213,N_3954,N_4680);
and U5214 (N_5214,N_2744,N_4919);
nor U5215 (N_5215,N_2788,N_3461);
nand U5216 (N_5216,N_3114,N_4572);
nand U5217 (N_5217,N_2620,N_4673);
and U5218 (N_5218,N_3512,N_4527);
and U5219 (N_5219,N_3100,N_2782);
and U5220 (N_5220,N_4846,N_2787);
nand U5221 (N_5221,N_2906,N_4294);
nand U5222 (N_5222,N_3624,N_4559);
nor U5223 (N_5223,N_4581,N_2704);
nand U5224 (N_5224,N_3528,N_4158);
nor U5225 (N_5225,N_4357,N_4640);
nand U5226 (N_5226,N_4449,N_4218);
xor U5227 (N_5227,N_3737,N_4711);
nor U5228 (N_5228,N_4258,N_2913);
or U5229 (N_5229,N_3642,N_3359);
or U5230 (N_5230,N_2910,N_2632);
or U5231 (N_5231,N_2848,N_3732);
or U5232 (N_5232,N_4786,N_4880);
and U5233 (N_5233,N_4350,N_3913);
and U5234 (N_5234,N_3542,N_2944);
or U5235 (N_5235,N_4187,N_3567);
or U5236 (N_5236,N_2911,N_3757);
nor U5237 (N_5237,N_3345,N_2950);
and U5238 (N_5238,N_2745,N_3228);
nand U5239 (N_5239,N_2977,N_3940);
and U5240 (N_5240,N_2947,N_3475);
or U5241 (N_5241,N_4653,N_3825);
nor U5242 (N_5242,N_4536,N_4769);
or U5243 (N_5243,N_2588,N_4795);
nor U5244 (N_5244,N_3777,N_3401);
and U5245 (N_5245,N_3152,N_3530);
or U5246 (N_5246,N_2798,N_2740);
nor U5247 (N_5247,N_4199,N_2797);
and U5248 (N_5248,N_3072,N_3871);
or U5249 (N_5249,N_3711,N_4684);
nor U5250 (N_5250,N_4895,N_4718);
and U5251 (N_5251,N_4979,N_3331);
nor U5252 (N_5252,N_2739,N_2671);
nor U5253 (N_5253,N_2526,N_2753);
and U5254 (N_5254,N_3580,N_3674);
and U5255 (N_5255,N_3582,N_4918);
or U5256 (N_5256,N_3853,N_3915);
and U5257 (N_5257,N_4897,N_3073);
nor U5258 (N_5258,N_3147,N_3708);
xnor U5259 (N_5259,N_3693,N_3746);
nand U5260 (N_5260,N_4204,N_4053);
nand U5261 (N_5261,N_3265,N_4591);
nor U5262 (N_5262,N_4847,N_4454);
or U5263 (N_5263,N_3077,N_4589);
xor U5264 (N_5264,N_4970,N_3447);
or U5265 (N_5265,N_2660,N_2732);
and U5266 (N_5266,N_3244,N_3070);
nor U5267 (N_5267,N_4400,N_3872);
and U5268 (N_5268,N_4982,N_2921);
xnor U5269 (N_5269,N_4469,N_4619);
or U5270 (N_5270,N_2651,N_2880);
nand U5271 (N_5271,N_4114,N_3414);
nand U5272 (N_5272,N_3368,N_3741);
or U5273 (N_5273,N_4451,N_3268);
xor U5274 (N_5274,N_4531,N_3826);
nor U5275 (N_5275,N_4045,N_4391);
or U5276 (N_5276,N_3828,N_3876);
or U5277 (N_5277,N_4379,N_4768);
and U5278 (N_5278,N_3549,N_3936);
or U5279 (N_5279,N_4626,N_4181);
and U5280 (N_5280,N_4992,N_3049);
or U5281 (N_5281,N_2680,N_4007);
nor U5282 (N_5282,N_4946,N_4525);
nor U5283 (N_5283,N_3022,N_4520);
and U5284 (N_5284,N_4180,N_3909);
nor U5285 (N_5285,N_2610,N_2733);
nand U5286 (N_5286,N_3546,N_4719);
nand U5287 (N_5287,N_2752,N_3063);
xor U5288 (N_5288,N_2648,N_3720);
nor U5289 (N_5289,N_4129,N_4930);
xnor U5290 (N_5290,N_2954,N_3979);
nor U5291 (N_5291,N_4260,N_2631);
or U5292 (N_5292,N_3245,N_2650);
nand U5293 (N_5293,N_3577,N_2529);
nand U5294 (N_5294,N_3886,N_3655);
nor U5295 (N_5295,N_3361,N_4337);
and U5296 (N_5296,N_3238,N_3620);
and U5297 (N_5297,N_2642,N_4839);
or U5298 (N_5298,N_4409,N_4920);
nor U5299 (N_5299,N_4256,N_3419);
nor U5300 (N_5300,N_3332,N_2681);
and U5301 (N_5301,N_3774,N_4343);
or U5302 (N_5302,N_2501,N_3626);
or U5303 (N_5303,N_4438,N_2946);
or U5304 (N_5304,N_2893,N_4784);
and U5305 (N_5305,N_4549,N_4821);
or U5306 (N_5306,N_3604,N_4904);
and U5307 (N_5307,N_3957,N_3834);
nor U5308 (N_5308,N_4668,N_3744);
nand U5309 (N_5309,N_4200,N_4632);
nand U5310 (N_5310,N_3455,N_3404);
nand U5311 (N_5311,N_3456,N_3910);
and U5312 (N_5312,N_3240,N_4174);
nor U5313 (N_5313,N_4703,N_3525);
or U5314 (N_5314,N_2927,N_3873);
or U5315 (N_5315,N_3562,N_3921);
or U5316 (N_5316,N_4202,N_3202);
nor U5317 (N_5317,N_4005,N_3659);
nand U5318 (N_5318,N_4615,N_3949);
nor U5319 (N_5319,N_4383,N_3589);
and U5320 (N_5320,N_3204,N_3207);
nor U5321 (N_5321,N_2873,N_4600);
nand U5322 (N_5322,N_4417,N_3875);
and U5323 (N_5323,N_3899,N_4573);
or U5324 (N_5324,N_3817,N_3827);
nor U5325 (N_5325,N_4613,N_4714);
nor U5326 (N_5326,N_4220,N_2846);
nor U5327 (N_5327,N_3432,N_2686);
nor U5328 (N_5328,N_4601,N_2543);
and U5329 (N_5329,N_3253,N_2557);
or U5330 (N_5330,N_4463,N_3751);
nand U5331 (N_5331,N_3264,N_2858);
nor U5332 (N_5332,N_3014,N_2843);
or U5333 (N_5333,N_3931,N_4326);
and U5334 (N_5334,N_3637,N_3366);
nand U5335 (N_5335,N_3120,N_3125);
nand U5336 (N_5336,N_2866,N_4843);
and U5337 (N_5337,N_3608,N_4375);
nor U5338 (N_5338,N_3928,N_4239);
and U5339 (N_5339,N_3192,N_4207);
or U5340 (N_5340,N_3307,N_4796);
and U5341 (N_5341,N_2695,N_4713);
nor U5342 (N_5342,N_3016,N_4608);
and U5343 (N_5343,N_3273,N_2823);
nor U5344 (N_5344,N_3524,N_4741);
nand U5345 (N_5345,N_3691,N_2998);
nor U5346 (N_5346,N_4069,N_2909);
and U5347 (N_5347,N_3636,N_4393);
or U5348 (N_5348,N_4254,N_3464);
xor U5349 (N_5349,N_3395,N_4881);
nand U5350 (N_5350,N_4404,N_3671);
nor U5351 (N_5351,N_4862,N_4178);
nand U5352 (N_5352,N_3801,N_4168);
and U5353 (N_5353,N_3129,N_4606);
nor U5354 (N_5354,N_2555,N_2718);
and U5355 (N_5355,N_2553,N_4269);
or U5356 (N_5356,N_4614,N_3785);
or U5357 (N_5357,N_2983,N_4942);
or U5358 (N_5358,N_2854,N_2721);
and U5359 (N_5359,N_3031,N_4810);
nand U5360 (N_5360,N_4130,N_4866);
or U5361 (N_5361,N_3765,N_4363);
or U5362 (N_5362,N_2685,N_4767);
nand U5363 (N_5363,N_3059,N_4980);
or U5364 (N_5364,N_2654,N_3866);
nand U5365 (N_5365,N_3088,N_3793);
or U5366 (N_5366,N_4938,N_3564);
nor U5367 (N_5367,N_2682,N_4683);
nor U5368 (N_5368,N_3182,N_4115);
and U5369 (N_5369,N_3937,N_3193);
nand U5370 (N_5370,N_4093,N_4354);
nor U5371 (N_5371,N_3598,N_4550);
or U5372 (N_5372,N_4757,N_3064);
or U5373 (N_5373,N_3187,N_3043);
nor U5374 (N_5374,N_3442,N_3983);
and U5375 (N_5375,N_3830,N_3602);
nor U5376 (N_5376,N_4398,N_2724);
nor U5377 (N_5377,N_3232,N_4558);
and U5378 (N_5378,N_4104,N_2503);
and U5379 (N_5379,N_3838,N_4772);
nand U5380 (N_5380,N_4709,N_3792);
nor U5381 (N_5381,N_3033,N_4864);
or U5382 (N_5382,N_3545,N_3229);
and U5383 (N_5383,N_4249,N_4395);
nor U5384 (N_5384,N_4171,N_4694);
or U5385 (N_5385,N_4655,N_2759);
and U5386 (N_5386,N_4118,N_2807);
and U5387 (N_5387,N_3648,N_2972);
nor U5388 (N_5388,N_3393,N_2853);
or U5389 (N_5389,N_3672,N_3733);
and U5390 (N_5390,N_3707,N_2592);
and U5391 (N_5391,N_4319,N_4165);
xor U5392 (N_5392,N_2643,N_2584);
nor U5393 (N_5393,N_4245,N_3380);
xnor U5394 (N_5394,N_2687,N_4771);
or U5395 (N_5395,N_3563,N_3681);
nor U5396 (N_5396,N_3329,N_3618);
nor U5397 (N_5397,N_4813,N_2862);
nor U5398 (N_5398,N_4112,N_4860);
nand U5399 (N_5399,N_4382,N_3491);
and U5400 (N_5400,N_3684,N_2522);
nand U5401 (N_5401,N_3142,N_4793);
or U5402 (N_5402,N_3771,N_4465);
and U5403 (N_5403,N_4477,N_2703);
nor U5404 (N_5404,N_3816,N_3312);
or U5405 (N_5405,N_3326,N_4022);
and U5406 (N_5406,N_3947,N_4085);
or U5407 (N_5407,N_3135,N_2514);
and U5408 (N_5408,N_3484,N_2743);
and U5409 (N_5409,N_2500,N_3013);
or U5410 (N_5410,N_3370,N_2528);
and U5411 (N_5411,N_2596,N_3647);
and U5412 (N_5412,N_4210,N_4936);
nor U5413 (N_5413,N_3474,N_3165);
or U5414 (N_5414,N_3194,N_3427);
and U5415 (N_5415,N_4373,N_4825);
nor U5416 (N_5416,N_2888,N_4442);
and U5417 (N_5417,N_2986,N_3086);
nand U5418 (N_5418,N_3948,N_3159);
nand U5419 (N_5419,N_3422,N_2608);
nand U5420 (N_5420,N_2656,N_3048);
or U5421 (N_5421,N_2623,N_3166);
and U5422 (N_5422,N_4564,N_3725);
and U5423 (N_5423,N_4902,N_3500);
nand U5424 (N_5424,N_4792,N_2808);
nor U5425 (N_5425,N_3314,N_3327);
and U5426 (N_5426,N_4063,N_4339);
nor U5427 (N_5427,N_3136,N_4137);
and U5428 (N_5428,N_4027,N_3167);
or U5429 (N_5429,N_4939,N_4716);
nand U5430 (N_5430,N_3481,N_3786);
or U5431 (N_5431,N_4041,N_3358);
nor U5432 (N_5432,N_4991,N_3927);
or U5433 (N_5433,N_2711,N_2585);
nor U5434 (N_5434,N_4812,N_3883);
nor U5435 (N_5435,N_3944,N_3344);
nor U5436 (N_5436,N_3999,N_3286);
nor U5437 (N_5437,N_3700,N_2845);
and U5438 (N_5438,N_2958,N_3548);
nor U5439 (N_5439,N_3338,N_4954);
or U5440 (N_5440,N_3112,N_3203);
nand U5441 (N_5441,N_3068,N_4586);
and U5442 (N_5442,N_3639,N_2816);
and U5443 (N_5443,N_3426,N_3300);
and U5444 (N_5444,N_3813,N_3814);
nor U5445 (N_5445,N_4408,N_3398);
or U5446 (N_5446,N_4805,N_2688);
nand U5447 (N_5447,N_4967,N_3532);
and U5448 (N_5448,N_2794,N_3946);
nand U5449 (N_5449,N_2615,N_3702);
nor U5450 (N_5450,N_4726,N_4648);
and U5451 (N_5451,N_4265,N_2532);
and U5452 (N_5452,N_3942,N_2665);
nand U5453 (N_5453,N_2869,N_4482);
xor U5454 (N_5454,N_3079,N_3560);
nand U5455 (N_5455,N_2974,N_3901);
nor U5456 (N_5456,N_3034,N_3216);
nor U5457 (N_5457,N_3995,N_4884);
nor U5458 (N_5458,N_4916,N_3865);
nand U5459 (N_5459,N_2590,N_2525);
and U5460 (N_5460,N_3713,N_2952);
and U5461 (N_5461,N_2626,N_4135);
and U5462 (N_5462,N_4751,N_3971);
nor U5463 (N_5463,N_4734,N_3980);
and U5464 (N_5464,N_2603,N_2661);
and U5465 (N_5465,N_2738,N_3958);
and U5466 (N_5466,N_4320,N_4941);
or U5467 (N_5467,N_4910,N_4025);
nand U5468 (N_5468,N_3018,N_4937);
or U5469 (N_5469,N_3256,N_4422);
nor U5470 (N_5470,N_3701,N_2919);
and U5471 (N_5471,N_3402,N_4074);
nor U5472 (N_5472,N_4075,N_4776);
nor U5473 (N_5473,N_2624,N_4252);
or U5474 (N_5474,N_4541,N_2517);
nand U5475 (N_5475,N_4457,N_2666);
and U5476 (N_5476,N_3622,N_2670);
and U5477 (N_5477,N_3824,N_4867);
or U5478 (N_5478,N_4308,N_2747);
nand U5479 (N_5479,N_4289,N_3880);
or U5480 (N_5480,N_4700,N_3161);
nor U5481 (N_5481,N_4685,N_4560);
or U5482 (N_5482,N_3150,N_3027);
nor U5483 (N_5483,N_4290,N_3799);
nand U5484 (N_5484,N_2679,N_3664);
nand U5485 (N_5485,N_3148,N_3287);
or U5486 (N_5486,N_3956,N_4540);
nand U5487 (N_5487,N_3284,N_3967);
or U5488 (N_5488,N_4605,N_3236);
and U5489 (N_5489,N_3721,N_2771);
or U5490 (N_5490,N_4724,N_4111);
nor U5491 (N_5491,N_2883,N_4459);
and U5492 (N_5492,N_2641,N_4015);
and U5493 (N_5493,N_2542,N_4898);
or U5494 (N_5494,N_2662,N_4506);
and U5495 (N_5495,N_2940,N_4385);
or U5496 (N_5496,N_4508,N_4173);
nor U5497 (N_5497,N_2502,N_4926);
nor U5498 (N_5498,N_2799,N_2948);
and U5499 (N_5499,N_4455,N_3103);
nor U5500 (N_5500,N_3668,N_3650);
nand U5501 (N_5501,N_3970,N_2923);
nand U5502 (N_5502,N_4346,N_4566);
and U5503 (N_5503,N_3551,N_4259);
nand U5504 (N_5504,N_2579,N_4983);
nor U5505 (N_5505,N_3806,N_4844);
nand U5506 (N_5506,N_4814,N_3369);
or U5507 (N_5507,N_3917,N_4280);
or U5508 (N_5508,N_4081,N_3037);
or U5509 (N_5509,N_3330,N_3180);
nand U5510 (N_5510,N_2618,N_4957);
or U5511 (N_5511,N_4389,N_3561);
nand U5512 (N_5512,N_3199,N_4512);
and U5513 (N_5513,N_4467,N_4542);
xnor U5514 (N_5514,N_3576,N_3762);
nor U5515 (N_5515,N_4546,N_3340);
or U5516 (N_5516,N_3262,N_4911);
or U5517 (N_5517,N_4838,N_3543);
nand U5518 (N_5518,N_3157,N_4958);
or U5519 (N_5519,N_2826,N_3748);
and U5520 (N_5520,N_4607,N_3270);
or U5521 (N_5521,N_4262,N_4787);
nor U5522 (N_5522,N_3015,N_2991);
nor U5523 (N_5523,N_4123,N_4431);
or U5524 (N_5524,N_4890,N_2763);
or U5525 (N_5525,N_4959,N_3087);
nand U5526 (N_5526,N_2614,N_4687);
nor U5527 (N_5527,N_4325,N_4677);
or U5528 (N_5528,N_4068,N_3663);
nand U5529 (N_5529,N_3565,N_3488);
or U5530 (N_5530,N_2563,N_3843);
nand U5531 (N_5531,N_2774,N_4761);
or U5532 (N_5532,N_3884,N_4080);
or U5533 (N_5533,N_3058,N_2635);
or U5534 (N_5534,N_3966,N_4018);
xnor U5535 (N_5535,N_3324,N_2545);
xnor U5536 (N_5536,N_4748,N_4675);
and U5537 (N_5537,N_3968,N_3178);
nand U5538 (N_5538,N_3673,N_4841);
and U5539 (N_5539,N_4460,N_2672);
nand U5540 (N_5540,N_3688,N_2801);
or U5541 (N_5541,N_3123,N_3084);
nor U5542 (N_5542,N_3343,N_2776);
nand U5543 (N_5543,N_3788,N_4961);
nor U5544 (N_5544,N_3162,N_3296);
and U5545 (N_5545,N_3924,N_2537);
or U5546 (N_5546,N_3209,N_3728);
nand U5547 (N_5547,N_2939,N_4661);
or U5548 (N_5548,N_3399,N_3466);
or U5549 (N_5549,N_3400,N_2837);
nand U5550 (N_5550,N_2904,N_3096);
nor U5551 (N_5551,N_4401,N_4062);
or U5552 (N_5552,N_2784,N_4362);
and U5553 (N_5553,N_4698,N_3657);
and U5554 (N_5554,N_3482,N_2601);
and U5555 (N_5555,N_4380,N_2885);
nand U5556 (N_5556,N_3590,N_3540);
or U5557 (N_5557,N_2890,N_3313);
nand U5558 (N_5558,N_4296,N_3093);
or U5559 (N_5559,N_4785,N_4552);
or U5560 (N_5560,N_2995,N_3996);
nand U5561 (N_5561,N_4635,N_3467);
and U5562 (N_5562,N_4585,N_3521);
and U5563 (N_5563,N_4044,N_3766);
and U5564 (N_5564,N_3489,N_4999);
or U5565 (N_5565,N_3583,N_3763);
and U5566 (N_5566,N_3823,N_4809);
and U5567 (N_5567,N_4047,N_2559);
nor U5568 (N_5568,N_3646,N_4828);
and U5569 (N_5569,N_2561,N_4150);
and U5570 (N_5570,N_2600,N_3945);
xor U5571 (N_5571,N_4396,N_3040);
nor U5572 (N_5572,N_3279,N_4544);
nand U5573 (N_5573,N_3354,N_2945);
nand U5574 (N_5574,N_4462,N_4208);
nand U5575 (N_5575,N_2551,N_3579);
and U5576 (N_5576,N_4834,N_4046);
nand U5577 (N_5577,N_4037,N_4042);
nand U5578 (N_5578,N_4660,N_3463);
or U5579 (N_5579,N_4593,N_3752);
nor U5580 (N_5580,N_2838,N_3328);
nand U5581 (N_5581,N_3535,N_4569);
nor U5582 (N_5582,N_2720,N_2898);
nand U5583 (N_5583,N_3175,N_4799);
nor U5584 (N_5584,N_3200,N_3503);
and U5585 (N_5585,N_4195,N_4050);
nor U5586 (N_5586,N_3840,N_3255);
and U5587 (N_5587,N_3889,N_2580);
nor U5588 (N_5588,N_4453,N_4800);
and U5589 (N_5589,N_4194,N_2839);
nor U5590 (N_5590,N_4054,N_3682);
and U5591 (N_5591,N_4824,N_4140);
nor U5592 (N_5592,N_3221,N_3504);
and U5593 (N_5593,N_2538,N_3082);
and U5594 (N_5594,N_2822,N_4806);
nand U5595 (N_5595,N_2951,N_4281);
nor U5596 (N_5596,N_4227,N_3696);
or U5597 (N_5597,N_4225,N_4545);
or U5598 (N_5598,N_4358,N_4206);
nor U5599 (N_5599,N_3566,N_3754);
xnor U5600 (N_5600,N_3042,N_4298);
nand U5601 (N_5601,N_4372,N_4432);
or U5602 (N_5602,N_3457,N_3384);
or U5603 (N_5603,N_3115,N_4837);
nor U5604 (N_5604,N_4226,N_2769);
nor U5605 (N_5605,N_2605,N_2964);
and U5606 (N_5606,N_4456,N_3390);
nor U5607 (N_5607,N_3578,N_2994);
nand U5608 (N_5608,N_3789,N_4061);
nand U5609 (N_5609,N_3798,N_4376);
and U5610 (N_5610,N_3894,N_3529);
nand U5611 (N_5611,N_3643,N_3781);
or U5612 (N_5612,N_3411,N_3494);
nand U5613 (N_5613,N_2785,N_3617);
or U5614 (N_5614,N_2996,N_4906);
and U5615 (N_5615,N_3208,N_4723);
and U5616 (N_5616,N_4973,N_4251);
nor U5617 (N_5617,N_4028,N_3514);
nor U5618 (N_5618,N_4882,N_2640);
nand U5619 (N_5619,N_2675,N_4583);
and U5620 (N_5620,N_3697,N_4657);
nor U5621 (N_5621,N_2878,N_2708);
or U5622 (N_5622,N_3051,N_3372);
and U5623 (N_5623,N_3434,N_3882);
nor U5624 (N_5624,N_4725,N_3878);
nand U5625 (N_5625,N_2742,N_4276);
or U5626 (N_5626,N_3341,N_4197);
or U5627 (N_5627,N_3000,N_4185);
nand U5628 (N_5628,N_3299,N_4480);
or U5629 (N_5629,N_4929,N_4498);
nand U5630 (N_5630,N_4708,N_4086);
nand U5631 (N_5631,N_4873,N_4528);
nor U5632 (N_5632,N_4139,N_4515);
and U5633 (N_5633,N_3278,N_4434);
or U5634 (N_5634,N_2746,N_3282);
nor U5635 (N_5635,N_3520,N_3764);
and U5636 (N_5636,N_3879,N_3829);
or U5637 (N_5637,N_4690,N_4756);
nand U5638 (N_5638,N_3722,N_4788);
nand U5639 (N_5639,N_3951,N_4316);
nand U5640 (N_5640,N_3383,N_3163);
and U5641 (N_5641,N_3397,N_4295);
nor U5642 (N_5642,N_4893,N_2892);
nor U5643 (N_5643,N_3729,N_3272);
and U5644 (N_5644,N_2891,N_3984);
nor U5645 (N_5645,N_2936,N_4689);
nor U5646 (N_5646,N_3248,N_4826);
nand U5647 (N_5647,N_4894,N_2701);
or U5648 (N_5648,N_3686,N_4423);
nor U5649 (N_5649,N_3905,N_3523);
nor U5650 (N_5650,N_3133,N_3656);
and U5651 (N_5651,N_3887,N_2968);
nand U5652 (N_5652,N_4492,N_4654);
or U5653 (N_5653,N_2872,N_3800);
nand U5654 (N_5654,N_3943,N_4011);
nor U5655 (N_5655,N_3685,N_4679);
or U5656 (N_5656,N_3550,N_3164);
or U5657 (N_5657,N_3258,N_4688);
nor U5658 (N_5658,N_3055,N_4968);
or U5659 (N_5659,N_2527,N_4331);
nand U5660 (N_5660,N_3060,N_4628);
nor U5661 (N_5661,N_3486,N_4976);
or U5662 (N_5662,N_4141,N_3409);
nand U5663 (N_5663,N_4539,N_4868);
nand U5664 (N_5664,N_2530,N_4856);
and U5665 (N_5665,N_4519,N_4603);
nand U5666 (N_5666,N_3742,N_2560);
xor U5667 (N_5667,N_4625,N_4440);
nor U5668 (N_5668,N_3661,N_4598);
or U5669 (N_5669,N_4537,N_4038);
or U5670 (N_5670,N_4175,N_2882);
xnor U5671 (N_5671,N_3453,N_4056);
and U5672 (N_5672,N_3334,N_4750);
nand U5673 (N_5673,N_4040,N_2857);
or U5674 (N_5674,N_3436,N_3743);
xnor U5675 (N_5675,N_4312,N_4620);
and U5676 (N_5676,N_2594,N_2980);
and U5677 (N_5677,N_4927,N_4933);
or U5678 (N_5678,N_2591,N_2966);
nor U5679 (N_5679,N_2534,N_4735);
nor U5680 (N_5680,N_3075,N_4728);
nand U5681 (N_5681,N_2879,N_3634);
or U5682 (N_5682,N_4845,N_2856);
nand U5683 (N_5683,N_4246,N_3126);
nor U5684 (N_5684,N_3495,N_3241);
or U5685 (N_5685,N_3363,N_4529);
or U5686 (N_5686,N_3054,N_3885);
nor U5687 (N_5687,N_4833,N_3281);
or U5688 (N_5688,N_4696,N_4570);
nand U5689 (N_5689,N_3437,N_3859);
nor U5690 (N_5690,N_4365,N_4349);
and U5691 (N_5691,N_3056,N_4943);
or U5692 (N_5692,N_3767,N_4547);
or U5693 (N_5693,N_3874,N_3274);
and U5694 (N_5694,N_2659,N_3895);
nor U5695 (N_5695,N_2992,N_4905);
nand U5696 (N_5696,N_2604,N_4023);
and U5697 (N_5697,N_2691,N_3985);
and U5698 (N_5698,N_2520,N_2505);
or U5699 (N_5699,N_4475,N_3251);
nor U5700 (N_5700,N_4124,N_3091);
or U5701 (N_5701,N_2935,N_3538);
nor U5702 (N_5702,N_3490,N_3502);
or U5703 (N_5703,N_3425,N_4755);
and U5704 (N_5704,N_4794,N_3558);
or U5705 (N_5705,N_3478,N_3130);
xnor U5706 (N_5706,N_3185,N_4087);
and U5707 (N_5707,N_4773,N_3808);
nand U5708 (N_5708,N_3953,N_3727);
and U5709 (N_5709,N_2655,N_3172);
and U5710 (N_5710,N_2988,N_3621);
nor U5711 (N_5711,N_3440,N_3812);
nor U5712 (N_5712,N_3554,N_4662);
or U5713 (N_5713,N_4978,N_3012);
nand U5714 (N_5714,N_4485,N_2581);
or U5715 (N_5715,N_4778,N_3645);
and U5716 (N_5716,N_3333,N_2953);
and U5717 (N_5717,N_3290,N_4163);
nand U5718 (N_5718,N_4117,N_2636);
xor U5719 (N_5719,N_3134,N_4565);
nand U5720 (N_5720,N_3320,N_2933);
or U5721 (N_5721,N_3470,N_3095);
nand U5722 (N_5722,N_2855,N_3321);
or U5723 (N_5723,N_4848,N_2969);
xnor U5724 (N_5724,N_3595,N_4962);
nor U5725 (N_5725,N_3715,N_4909);
and U5726 (N_5726,N_4858,N_4987);
nand U5727 (N_5727,N_3092,N_3024);
or U5728 (N_5728,N_3930,N_3477);
nand U5729 (N_5729,N_4851,N_3526);
or U5730 (N_5730,N_4674,N_4995);
and U5731 (N_5731,N_3510,N_2617);
nor U5732 (N_5732,N_3323,N_3127);
nand U5733 (N_5733,N_4596,N_4419);
or U5734 (N_5734,N_2825,N_3170);
xor U5735 (N_5735,N_3632,N_3704);
or U5736 (N_5736,N_2840,N_3357);
and U5737 (N_5737,N_2727,N_4198);
or U5738 (N_5738,N_4000,N_3687);
nand U5739 (N_5739,N_3065,N_2931);
nand U5740 (N_5740,N_4324,N_2999);
or U5741 (N_5741,N_3465,N_4058);
nor U5742 (N_5742,N_3881,N_3469);
nor U5743 (N_5743,N_3537,N_3938);
nand U5744 (N_5744,N_3215,N_2510);
xor U5745 (N_5745,N_3348,N_3007);
and U5746 (N_5746,N_2820,N_4588);
nor U5747 (N_5747,N_4297,N_4307);
and U5748 (N_5748,N_4861,N_4820);
or U5749 (N_5749,N_2915,N_4255);
nor U5750 (N_5750,N_2942,N_4503);
and U5751 (N_5751,N_4831,N_2962);
nor U5752 (N_5752,N_2766,N_4452);
nand U5753 (N_5753,N_4505,N_2705);
and U5754 (N_5754,N_4887,N_4908);
and U5755 (N_5755,N_4514,N_4283);
and U5756 (N_5756,N_2697,N_4517);
nand U5757 (N_5757,N_3146,N_3438);
nand U5758 (N_5758,N_4522,N_2760);
nand U5759 (N_5759,N_4815,N_4779);
nand U5760 (N_5760,N_4644,N_4649);
nand U5761 (N_5761,N_4102,N_2960);
nor U5762 (N_5762,N_2750,N_4100);
xor U5763 (N_5763,N_3444,N_4424);
nor U5764 (N_5764,N_2577,N_3585);
nor U5765 (N_5765,N_2895,N_3753);
nand U5766 (N_5766,N_4076,N_4243);
nor U5767 (N_5767,N_3613,N_3908);
nand U5768 (N_5768,N_3782,N_2886);
nand U5769 (N_5769,N_3005,N_2569);
or U5770 (N_5770,N_3035,N_4553);
nor U5771 (N_5771,N_3662,N_4891);
nor U5772 (N_5772,N_3109,N_3374);
nand U5773 (N_5773,N_3571,N_2887);
or U5774 (N_5774,N_4234,N_4224);
nor U5775 (N_5775,N_2541,N_4418);
nor U5776 (N_5776,N_2990,N_3804);
and U5777 (N_5777,N_3138,N_4557);
and U5778 (N_5778,N_4827,N_3462);
nand U5779 (N_5779,N_3877,N_2834);
and U5780 (N_5780,N_3066,N_3090);
and U5781 (N_5781,N_3021,N_3242);
or U5782 (N_5782,N_3679,N_2719);
and U5783 (N_5783,N_3310,N_4268);
and U5784 (N_5784,N_3675,N_3254);
nor U5785 (N_5785,N_2593,N_3988);
and U5786 (N_5786,N_4516,N_2976);
nor U5787 (N_5787,N_2509,N_2754);
and U5788 (N_5788,N_2971,N_4145);
nand U5789 (N_5789,N_3841,N_2836);
nor U5790 (N_5790,N_4196,N_4742);
nor U5791 (N_5791,N_2767,N_4032);
or U5792 (N_5792,N_3508,N_3615);
or U5793 (N_5793,N_2597,N_2761);
or U5794 (N_5794,N_4031,N_4739);
nand U5795 (N_5795,N_4950,N_4610);
nor U5796 (N_5796,N_2916,N_4302);
nor U5797 (N_5797,N_3692,N_2578);
nor U5798 (N_5798,N_3403,N_4836);
or U5799 (N_5799,N_4318,N_3104);
and U5800 (N_5800,N_4055,N_4502);
or U5801 (N_5801,N_3920,N_4984);
nor U5802 (N_5802,N_3796,N_3429);
or U5803 (N_5803,N_2595,N_4484);
or U5804 (N_5804,N_4623,N_3379);
or U5805 (N_5805,N_3275,N_3212);
and U5806 (N_5806,N_3833,N_3099);
nor U5807 (N_5807,N_3292,N_3317);
nor U5808 (N_5808,N_4416,N_4070);
nand U5809 (N_5809,N_4960,N_3206);
nand U5810 (N_5810,N_3717,N_2832);
nor U5811 (N_5811,N_3391,N_4261);
or U5812 (N_5812,N_4989,N_3977);
nor U5813 (N_5813,N_3151,N_4731);
or U5814 (N_5814,N_3667,N_4746);
nor U5815 (N_5815,N_4377,N_4203);
and U5816 (N_5816,N_4402,N_3969);
and U5817 (N_5817,N_4732,N_3173);
and U5818 (N_5818,N_3847,N_2981);
and U5819 (N_5819,N_3352,N_4681);
nand U5820 (N_5820,N_4361,N_4486);
and U5821 (N_5821,N_3097,N_4474);
nor U5822 (N_5822,N_4336,N_4921);
nor U5823 (N_5823,N_4072,N_4369);
nor U5824 (N_5824,N_3181,N_2943);
nand U5825 (N_5825,N_3496,N_3026);
nand U5826 (N_5826,N_3230,N_4212);
nor U5827 (N_5827,N_4996,N_4388);
nor U5828 (N_5828,N_3023,N_4693);
nand U5829 (N_5829,N_3527,N_3283);
or U5830 (N_5830,N_3981,N_3235);
nor U5831 (N_5831,N_4242,N_2706);
and U5832 (N_5832,N_3832,N_4221);
nand U5833 (N_5833,N_4125,N_4155);
and U5834 (N_5834,N_3705,N_4783);
and U5835 (N_5835,N_2613,N_3213);
and U5836 (N_5836,N_3385,N_3472);
nor U5837 (N_5837,N_3837,N_3694);
nand U5838 (N_5838,N_3644,N_3271);
or U5839 (N_5839,N_3260,N_4010);
and U5840 (N_5840,N_2611,N_3822);
or U5841 (N_5841,N_2565,N_4807);
nor U5842 (N_5842,N_3293,N_3890);
and U5843 (N_5843,N_4406,N_3020);
or U5844 (N_5844,N_4595,N_3689);
nor U5845 (N_5845,N_3719,N_4637);
nor U5846 (N_5846,N_4335,N_3266);
and U5847 (N_5847,N_4300,N_4273);
nand U5848 (N_5848,N_4715,N_3575);
nor U5849 (N_5849,N_4977,N_3776);
nor U5850 (N_5850,N_4116,N_3863);
nor U5851 (N_5851,N_4483,N_4730);
nor U5852 (N_5852,N_4816,N_3994);
and U5853 (N_5853,N_2586,N_4944);
and U5854 (N_5854,N_4830,N_3739);
xor U5855 (N_5855,N_2558,N_4279);
and U5856 (N_5856,N_3239,N_4229);
and U5857 (N_5857,N_4083,N_4159);
and U5858 (N_5858,N_4403,N_4953);
nand U5859 (N_5859,N_4965,N_4186);
or U5860 (N_5860,N_3950,N_4157);
and U5861 (N_5861,N_4682,N_3787);
nor U5862 (N_5862,N_3053,N_3038);
or U5863 (N_5863,N_4576,N_4811);
nand U5864 (N_5864,N_4643,N_4669);
or U5865 (N_5865,N_4386,N_4160);
nor U5866 (N_5866,N_4476,N_4513);
and U5867 (N_5867,N_4790,N_2932);
and U5868 (N_5868,N_4738,N_2731);
nor U5869 (N_5869,N_4314,N_4823);
and U5870 (N_5870,N_3473,N_2790);
nor U5871 (N_5871,N_2702,N_4780);
nand U5872 (N_5872,N_3407,N_4154);
or U5873 (N_5873,N_4510,N_3591);
nand U5874 (N_5874,N_4985,N_4240);
xor U5875 (N_5875,N_4310,N_4446);
and U5876 (N_5876,N_4213,N_2804);
and U5877 (N_5877,N_3531,N_4571);
nor U5878 (N_5878,N_3386,N_3375);
and U5879 (N_5879,N_4701,N_2627);
nor U5880 (N_5880,N_3364,N_3857);
and U5881 (N_5881,N_4466,N_4002);
and U5882 (N_5882,N_3935,N_4043);
nand U5883 (N_5883,N_3128,N_3252);
or U5884 (N_5884,N_3934,N_4340);
nor U5885 (N_5885,N_4109,N_3458);
and U5886 (N_5886,N_3387,N_4192);
nor U5887 (N_5887,N_3987,N_3493);
nand U5888 (N_5888,N_3964,N_3301);
and U5889 (N_5889,N_4509,N_4230);
and U5890 (N_5890,N_2713,N_4113);
or U5891 (N_5891,N_4777,N_2649);
nand U5892 (N_5892,N_4131,N_4019);
and U5893 (N_5893,N_4119,N_4804);
or U5894 (N_5894,N_2984,N_4214);
nand U5895 (N_5895,N_3113,N_3085);
and U5896 (N_5896,N_4012,N_3408);
and U5897 (N_5897,N_3810,N_3716);
nand U5898 (N_5898,N_3139,N_2905);
or U5899 (N_5899,N_4132,N_3603);
nand U5900 (N_5900,N_3449,N_3519);
or U5901 (N_5901,N_4886,N_4672);
and U5902 (N_5902,N_3111,N_4096);
or U5903 (N_5903,N_4753,N_3376);
or U5904 (N_5904,N_4859,N_3631);
nor U5905 (N_5905,N_3773,N_3665);
and U5906 (N_5906,N_2914,N_3441);
or U5907 (N_5907,N_4744,N_3553);
nand U5908 (N_5908,N_2533,N_4282);
nor U5909 (N_5909,N_3342,N_3573);
or U5910 (N_5910,N_4201,N_2722);
nor U5911 (N_5911,N_3633,N_3536);
or U5912 (N_5912,N_3160,N_3335);
nor U5913 (N_5913,N_4609,N_3852);
or U5914 (N_5914,N_2778,N_4650);
or U5915 (N_5915,N_3454,N_3098);
or U5916 (N_5916,N_4270,N_4646);
nor U5917 (N_5917,N_4764,N_3036);
nand U5918 (N_5918,N_2612,N_4458);
nor U5919 (N_5919,N_3902,N_4162);
nand U5920 (N_5920,N_3285,N_2570);
xnor U5921 (N_5921,N_2599,N_4594);
nand U5922 (N_5922,N_3505,N_4872);
and U5923 (N_5923,N_4333,N_3416);
or U5924 (N_5924,N_4412,N_3611);
or U5925 (N_5925,N_4896,N_3846);
nand U5926 (N_5926,N_4763,N_4128);
nor U5927 (N_5927,N_2884,N_4543);
or U5928 (N_5928,N_4436,N_4618);
nand U5929 (N_5929,N_3775,N_3836);
and U5930 (N_5930,N_3267,N_3394);
nor U5931 (N_5931,N_4110,N_2511);
and U5932 (N_5932,N_4078,N_3677);
or U5933 (N_5933,N_3316,N_3476);
and U5934 (N_5934,N_3745,N_3201);
nand U5935 (N_5935,N_4184,N_4378);
nor U5936 (N_5936,N_3004,N_3522);
or U5937 (N_5937,N_4253,N_3740);
and U5938 (N_5938,N_3450,N_3849);
nor U5939 (N_5939,N_2736,N_3619);
nor U5940 (N_5940,N_3651,N_4487);
and U5941 (N_5941,N_2978,N_2714);
or U5942 (N_5942,N_4892,N_4782);
or U5943 (N_5943,N_4917,N_3892);
or U5944 (N_5944,N_3820,N_3978);
nor U5945 (N_5945,N_3101,N_4228);
and U5946 (N_5946,N_4579,N_3224);
or U5947 (N_5947,N_4292,N_3976);
nand U5948 (N_5948,N_4707,N_3678);
and U5949 (N_5949,N_3205,N_3628);
or U5950 (N_5950,N_4932,N_2571);
nor U5951 (N_5951,N_2689,N_4232);
or U5952 (N_5952,N_3226,N_3143);
and U5953 (N_5953,N_4656,N_2907);
and U5954 (N_5954,N_3076,N_2926);
nand U5955 (N_5955,N_3552,N_3110);
or U5956 (N_5956,N_4791,N_3641);
nand U5957 (N_5957,N_2783,N_3698);
or U5958 (N_5958,N_3652,N_2975);
nor U5959 (N_5959,N_3237,N_2634);
nor U5960 (N_5960,N_2941,N_3047);
and U5961 (N_5961,N_4523,N_4580);
and U5962 (N_5962,N_4341,N_2589);
nand U5963 (N_5963,N_2564,N_3658);
or U5964 (N_5964,N_3431,N_2583);
nor U5965 (N_5965,N_2737,N_3080);
and U5966 (N_5966,N_3498,N_3690);
and U5967 (N_5967,N_4819,N_4500);
or U5968 (N_5968,N_4288,N_3779);
or U5969 (N_5969,N_4170,N_4468);
nor U5970 (N_5970,N_3217,N_4433);
nor U5971 (N_5971,N_2959,N_4692);
nor U5972 (N_5972,N_4556,N_4321);
nor U5973 (N_5973,N_4381,N_3912);
or U5974 (N_5974,N_3305,N_4429);
nor U5975 (N_5975,N_4789,N_4922);
nand U5976 (N_5976,N_4667,N_4752);
and U5977 (N_5977,N_3336,N_2792);
nand U5978 (N_5978,N_3196,N_2811);
or U5979 (N_5979,N_4818,N_4067);
nand U5980 (N_5980,N_3210,N_4955);
and U5981 (N_5981,N_2652,N_4008);
or U5982 (N_5982,N_4883,N_3057);
nand U5983 (N_5983,N_3156,N_3197);
and U5984 (N_5984,N_2818,N_4051);
nor U5985 (N_5985,N_4120,N_4182);
nor U5986 (N_5986,N_3190,N_3778);
nand U5987 (N_5987,N_3044,N_4624);
nand U5988 (N_5988,N_2864,N_3119);
or U5989 (N_5989,N_4499,N_3001);
nor U5990 (N_5990,N_3247,N_3288);
or U5991 (N_5991,N_4091,N_4014);
and U5992 (N_5992,N_4439,N_3029);
nor U5993 (N_5993,N_3306,N_2937);
nand U5994 (N_5994,N_3588,N_2707);
and U5995 (N_5995,N_4931,N_2827);
and U5996 (N_5996,N_4664,N_4712);
and U5997 (N_5997,N_3373,N_3858);
and U5998 (N_5998,N_2515,N_3670);
and U5999 (N_5999,N_3515,N_4172);
or U6000 (N_6000,N_4437,N_2863);
and U6001 (N_6001,N_4271,N_3277);
nor U6002 (N_6002,N_4161,N_3898);
nor U6003 (N_6003,N_3780,N_4327);
nand U6004 (N_6004,N_4759,N_3541);
and U6005 (N_6005,N_3761,N_4849);
nor U6006 (N_6006,N_3605,N_4237);
xnor U6007 (N_6007,N_2961,N_2674);
and U6008 (N_6008,N_2795,N_3017);
nand U6009 (N_6009,N_3925,N_2758);
and U6010 (N_6010,N_2852,N_2550);
nand U6011 (N_6011,N_3511,N_2985);
or U6012 (N_6012,N_3811,N_4975);
nand U6013 (N_6013,N_4526,N_4444);
or U6014 (N_6014,N_2668,N_2979);
and U6015 (N_6015,N_3010,N_4538);
and U6016 (N_6016,N_3225,N_3257);
nand U6017 (N_6017,N_3623,N_4697);
and U6018 (N_6018,N_3790,N_4840);
or U6019 (N_6019,N_2902,N_4888);
nor U6020 (N_6020,N_4974,N_3989);
nor U6021 (N_6021,N_4634,N_3074);
and U6022 (N_6022,N_4413,N_2723);
nor U6023 (N_6023,N_4754,N_3259);
nand U6024 (N_6024,N_4024,N_3914);
or U6025 (N_6025,N_3596,N_2755);
and U6026 (N_6026,N_4781,N_2710);
nor U6027 (N_6027,N_4360,N_2554);
or U6028 (N_6028,N_3365,N_3584);
and U6029 (N_6029,N_2967,N_2546);
and U6030 (N_6030,N_3614,N_4397);
and U6031 (N_6031,N_4347,N_4951);
nor U6032 (N_6032,N_2669,N_3738);
or U6033 (N_6033,N_3831,N_4720);
or U6034 (N_6034,N_4835,N_4066);
nand U6035 (N_6035,N_4870,N_3188);
nand U6036 (N_6036,N_4478,N_4832);
or U6037 (N_6037,N_4211,N_2647);
nor U6038 (N_6038,N_4445,N_4179);
or U6039 (N_6039,N_4189,N_3485);
nor U6040 (N_6040,N_4988,N_3718);
or U6041 (N_6041,N_4691,N_3507);
or U6042 (N_6042,N_2735,N_2765);
and U6043 (N_6043,N_3303,N_3108);
nor U6044 (N_6044,N_4138,N_2860);
nor U6045 (N_6045,N_3121,N_2536);
and U6046 (N_6046,N_4633,N_2877);
nor U6047 (N_6047,N_2851,N_4274);
xor U6048 (N_6048,N_2730,N_2989);
or U6049 (N_6049,N_4355,N_3509);
nand U6050 (N_6050,N_4524,N_4803);
or U6051 (N_6051,N_2657,N_3724);
nand U6052 (N_6052,N_2894,N_4706);
or U6053 (N_6053,N_3406,N_3714);
and U6054 (N_6054,N_3627,N_3802);
nor U6055 (N_6055,N_3756,N_4216);
or U6056 (N_6056,N_2918,N_4808);
nor U6057 (N_6057,N_2779,N_4368);
nor U6058 (N_6058,N_3747,N_4496);
nor U6059 (N_6059,N_2547,N_3353);
or U6060 (N_6060,N_2831,N_4344);
nand U6061 (N_6061,N_3145,N_3749);
nand U6062 (N_6062,N_3735,N_4317);
nor U6063 (N_6063,N_4602,N_3169);
nor U6064 (N_6064,N_4285,N_4670);
nand U6065 (N_6065,N_3557,N_3896);
nand U6066 (N_6066,N_3302,N_3959);
and U6067 (N_6067,N_4678,N_2567);
or U6068 (N_6068,N_4642,N_3349);
and U6069 (N_6069,N_4473,N_4869);
and U6070 (N_6070,N_4878,N_3640);
xnor U6071 (N_6071,N_2638,N_2645);
and U6072 (N_6072,N_4287,N_4127);
and U6073 (N_6073,N_2639,N_4582);
nand U6074 (N_6074,N_3791,N_4852);
nor U6075 (N_6075,N_2658,N_4146);
or U6076 (N_6076,N_2934,N_3480);
nand U6077 (N_6077,N_4562,N_4278);
and U6078 (N_6078,N_4430,N_4900);
nor U6079 (N_6079,N_4264,N_2955);
nor U6080 (N_6080,N_2548,N_4964);
or U6081 (N_6081,N_3572,N_2824);
or U6082 (N_6082,N_4994,N_4760);
or U6083 (N_6083,N_2756,N_3797);
or U6084 (N_6084,N_4193,N_2762);
nand U6085 (N_6085,N_3219,N_4394);
nand U6086 (N_6086,N_3568,N_4491);
or U6087 (N_6087,N_3993,N_3533);
or U6088 (N_6088,N_3845,N_2796);
and U6089 (N_6089,N_4064,N_4636);
or U6090 (N_6090,N_3518,N_3998);
nand U6091 (N_6091,N_4567,N_4577);
nor U6092 (N_6092,N_3234,N_2709);
nor U6093 (N_6093,N_3868,N_2749);
or U6094 (N_6094,N_3140,N_3177);
nand U6095 (N_6095,N_4494,N_4332);
nor U6096 (N_6096,N_3587,N_2813);
nand U6097 (N_6097,N_3420,N_3410);
or U6098 (N_6098,N_4555,N_4144);
nand U6099 (N_6099,N_3842,N_4901);
or U6100 (N_6100,N_3760,N_4652);
and U6101 (N_6101,N_3805,N_2828);
or U6102 (N_6102,N_4770,N_3081);
nor U6103 (N_6103,N_4169,N_3041);
and U6104 (N_6104,N_4190,N_2573);
and U6105 (N_6105,N_2963,N_4885);
or U6106 (N_6106,N_4616,N_3862);
nand U6107 (N_6107,N_2728,N_4293);
nand U6108 (N_6108,N_3712,N_3418);
or U6109 (N_6109,N_4136,N_4049);
nand U6110 (N_6110,N_2815,N_3367);
nand U6111 (N_6111,N_4152,N_2875);
or U6112 (N_6112,N_4299,N_4348);
and U6113 (N_6113,N_4740,N_3592);
or U6114 (N_6114,N_4176,N_2806);
nand U6115 (N_6115,N_3972,N_4464);
nand U6116 (N_6116,N_3350,N_3703);
nand U6117 (N_6117,N_4057,N_3952);
nand U6118 (N_6118,N_4059,N_2677);
and U6119 (N_6119,N_2726,N_3377);
nor U6120 (N_6120,N_3683,N_4903);
and U6121 (N_6121,N_3975,N_4026);
nand U6122 (N_6122,N_2757,N_3222);
nand U6123 (N_6123,N_2574,N_4143);
or U6124 (N_6124,N_3319,N_3680);
nor U6125 (N_6125,N_3003,N_4952);
nor U6126 (N_6126,N_4105,N_3630);
nor U6127 (N_6127,N_3304,N_3045);
or U6128 (N_6128,N_2535,N_3479);
nor U6129 (N_6129,N_3517,N_3706);
nor U6130 (N_6130,N_3132,N_3638);
and U6131 (N_6131,N_2842,N_4993);
and U6132 (N_6132,N_2970,N_3451);
nor U6133 (N_6133,N_4148,N_3821);
nand U6134 (N_6134,N_3249,N_3025);
or U6135 (N_6135,N_4030,N_4107);
or U6136 (N_6136,N_2812,N_2653);
nand U6137 (N_6137,N_4822,N_3122);
or U6138 (N_6138,N_2821,N_4387);
nand U6139 (N_6139,N_3032,N_3893);
and U6140 (N_6140,N_4367,N_4612);
or U6141 (N_6141,N_3600,N_3850);
or U6142 (N_6142,N_4802,N_2781);
or U6143 (N_6143,N_4004,N_3046);
nand U6144 (N_6144,N_2637,N_4421);
or U6145 (N_6145,N_2712,N_4359);
nand U6146 (N_6146,N_2993,N_4997);
and U6147 (N_6147,N_3220,N_2507);
nand U6148 (N_6148,N_3413,N_3986);
nor U6149 (N_6149,N_4003,N_3709);
or U6150 (N_6150,N_4551,N_4309);
nand U6151 (N_6151,N_3261,N_3597);
or U6152 (N_6152,N_4853,N_4147);
nand U6153 (N_6153,N_4704,N_4801);
nand U6154 (N_6154,N_3911,N_3855);
nand U6155 (N_6155,N_4597,N_4733);
and U6156 (N_6156,N_3635,N_4060);
or U6157 (N_6157,N_4850,N_4235);
and U6158 (N_6158,N_4651,N_3318);
and U6159 (N_6159,N_3539,N_2982);
nand U6160 (N_6160,N_4631,N_3297);
and U6161 (N_6161,N_2833,N_4863);
nor U6162 (N_6162,N_4156,N_2523);
or U6163 (N_6163,N_4749,N_3903);
nand U6164 (N_6164,N_4671,N_3870);
nor U6165 (N_6165,N_3263,N_3106);
nor U6166 (N_6166,N_3439,N_3906);
and U6167 (N_6167,N_4504,N_2997);
nor U6168 (N_6168,N_3191,N_2874);
or U6169 (N_6169,N_4981,N_3131);
or U6170 (N_6170,N_3900,N_4488);
nand U6171 (N_6171,N_3918,N_3555);
nor U6172 (N_6172,N_2607,N_4829);
nand U6173 (N_6173,N_3809,N_2598);
and U6174 (N_6174,N_3322,N_3445);
nand U6175 (N_6175,N_4568,N_3770);
nor U6176 (N_6176,N_3362,N_3295);
and U6177 (N_6177,N_4695,N_3654);
nor U6178 (N_6178,N_4384,N_3067);
or U6179 (N_6179,N_3415,N_4034);
nor U6180 (N_6180,N_4048,N_3137);
or U6181 (N_6181,N_2699,N_3758);
or U6182 (N_6182,N_2900,N_3897);
or U6183 (N_6183,N_4907,N_3028);
or U6184 (N_6184,N_4745,N_3396);
nor U6185 (N_6185,N_4899,N_3649);
nand U6186 (N_6186,N_3856,N_2539);
or U6187 (N_6187,N_3008,N_3570);
and U6188 (N_6188,N_4153,N_4420);
nor U6189 (N_6189,N_3459,N_3506);
and U6190 (N_6190,N_4621,N_4590);
or U6191 (N_6191,N_3183,N_4134);
or U6192 (N_6192,N_3513,N_4710);
nor U6193 (N_6193,N_3607,N_3198);
and U6194 (N_6194,N_2575,N_4966);
or U6195 (N_6195,N_4142,N_4405);
and U6196 (N_6196,N_3176,N_2896);
and U6197 (N_6197,N_3179,N_4924);
or U6198 (N_6198,N_3039,N_4986);
and U6199 (N_6199,N_3769,N_2512);
and U6200 (N_6200,N_3149,N_3939);
or U6201 (N_6201,N_3468,N_2928);
or U6202 (N_6202,N_4183,N_2562);
or U6203 (N_6203,N_4842,N_4470);
and U6204 (N_6204,N_4658,N_2692);
and U6205 (N_6205,N_3243,N_4306);
nor U6206 (N_6206,N_3378,N_3250);
nand U6207 (N_6207,N_4947,N_3492);
nand U6208 (N_6208,N_3599,N_3269);
and U6209 (N_6209,N_3483,N_3922);
nand U6210 (N_6210,N_3933,N_2676);
and U6211 (N_6211,N_4079,N_4126);
and U6212 (N_6212,N_2504,N_4164);
nor U6213 (N_6213,N_2814,N_2556);
nor U6214 (N_6214,N_4472,N_4736);
nor U6215 (N_6215,N_3006,N_3848);
nor U6216 (N_6216,N_3430,N_2925);
nor U6217 (N_6217,N_3963,N_3723);
nor U6218 (N_6218,N_4511,N_3768);
or U6219 (N_6219,N_4737,N_4676);
nor U6220 (N_6220,N_4854,N_2803);
nor U6221 (N_6221,N_4082,N_2949);
and U6222 (N_6222,N_3660,N_2920);
and U6223 (N_6223,N_4052,N_4798);
nor U6224 (N_6224,N_3381,N_4263);
or U6225 (N_6225,N_4065,N_4604);
nor U6226 (N_6226,N_2912,N_4097);
nor U6227 (N_6227,N_4257,N_2777);
or U6228 (N_6228,N_4663,N_4998);
nor U6229 (N_6229,N_3124,N_4722);
nor U6230 (N_6230,N_3569,N_2572);
or U6231 (N_6231,N_3982,N_3392);
nand U6232 (N_6232,N_4407,N_3298);
or U6233 (N_6233,N_2621,N_4122);
or U6234 (N_6234,N_4020,N_3676);
nor U6235 (N_6235,N_2519,N_4471);
nand U6236 (N_6236,N_4301,N_4575);
nor U6237 (N_6237,N_2518,N_3412);
and U6238 (N_6238,N_3516,N_2829);
nor U6239 (N_6239,N_3726,N_4665);
or U6240 (N_6240,N_3759,N_4611);
nand U6241 (N_6241,N_3888,N_2930);
and U6242 (N_6242,N_3609,N_4630);
or U6243 (N_6243,N_4374,N_3083);
or U6244 (N_6244,N_3371,N_2859);
and U6245 (N_6245,N_2876,N_3869);
nor U6246 (N_6246,N_3730,N_4441);
or U6247 (N_6247,N_3487,N_3189);
or U6248 (N_6248,N_2684,N_2622);
and U6249 (N_6249,N_3629,N_2850);
or U6250 (N_6250,N_2642,N_4313);
and U6251 (N_6251,N_3679,N_4356);
xnor U6252 (N_6252,N_4063,N_4985);
and U6253 (N_6253,N_2525,N_4307);
nand U6254 (N_6254,N_3266,N_3825);
nand U6255 (N_6255,N_3183,N_3503);
and U6256 (N_6256,N_4439,N_4592);
or U6257 (N_6257,N_2957,N_2859);
and U6258 (N_6258,N_4838,N_3647);
nand U6259 (N_6259,N_3622,N_3215);
nand U6260 (N_6260,N_2920,N_3819);
xor U6261 (N_6261,N_2944,N_3666);
nand U6262 (N_6262,N_3123,N_4713);
and U6263 (N_6263,N_3129,N_3367);
nor U6264 (N_6264,N_2935,N_3434);
nand U6265 (N_6265,N_4368,N_3973);
xnor U6266 (N_6266,N_2881,N_2771);
nor U6267 (N_6267,N_3097,N_4342);
or U6268 (N_6268,N_3231,N_3945);
or U6269 (N_6269,N_2989,N_4932);
nand U6270 (N_6270,N_4086,N_3708);
nor U6271 (N_6271,N_3565,N_4113);
nand U6272 (N_6272,N_3789,N_3464);
nor U6273 (N_6273,N_2752,N_2754);
and U6274 (N_6274,N_2852,N_4984);
nor U6275 (N_6275,N_3859,N_3710);
nand U6276 (N_6276,N_2625,N_3340);
nand U6277 (N_6277,N_3114,N_4069);
or U6278 (N_6278,N_4196,N_2673);
and U6279 (N_6279,N_3065,N_4164);
nor U6280 (N_6280,N_3688,N_2732);
and U6281 (N_6281,N_4124,N_3109);
or U6282 (N_6282,N_2753,N_4252);
or U6283 (N_6283,N_2742,N_3056);
xor U6284 (N_6284,N_2887,N_3743);
or U6285 (N_6285,N_4244,N_2552);
or U6286 (N_6286,N_4148,N_3962);
nand U6287 (N_6287,N_4549,N_3911);
nor U6288 (N_6288,N_3477,N_4939);
nor U6289 (N_6289,N_3890,N_3782);
or U6290 (N_6290,N_2575,N_3083);
and U6291 (N_6291,N_3633,N_3263);
and U6292 (N_6292,N_4736,N_3359);
xor U6293 (N_6293,N_4496,N_3554);
or U6294 (N_6294,N_4522,N_4757);
or U6295 (N_6295,N_4248,N_3981);
or U6296 (N_6296,N_2990,N_2962);
or U6297 (N_6297,N_2599,N_4261);
or U6298 (N_6298,N_2979,N_3319);
nor U6299 (N_6299,N_3737,N_4271);
nand U6300 (N_6300,N_4519,N_3800);
nor U6301 (N_6301,N_4829,N_2798);
and U6302 (N_6302,N_2897,N_2762);
and U6303 (N_6303,N_4651,N_3629);
or U6304 (N_6304,N_3583,N_2902);
or U6305 (N_6305,N_3027,N_2885);
nand U6306 (N_6306,N_3477,N_2853);
or U6307 (N_6307,N_3542,N_2595);
and U6308 (N_6308,N_4869,N_4435);
nor U6309 (N_6309,N_4540,N_3924);
and U6310 (N_6310,N_4785,N_4639);
nand U6311 (N_6311,N_2512,N_4324);
or U6312 (N_6312,N_2956,N_3212);
or U6313 (N_6313,N_3142,N_4566);
or U6314 (N_6314,N_4283,N_3062);
or U6315 (N_6315,N_4885,N_3069);
and U6316 (N_6316,N_4443,N_4359);
and U6317 (N_6317,N_3124,N_2606);
or U6318 (N_6318,N_3864,N_3070);
nor U6319 (N_6319,N_2963,N_4878);
nand U6320 (N_6320,N_3710,N_2792);
and U6321 (N_6321,N_2684,N_3658);
nand U6322 (N_6322,N_3702,N_3834);
nor U6323 (N_6323,N_3050,N_4267);
or U6324 (N_6324,N_4999,N_3117);
nand U6325 (N_6325,N_2750,N_2869);
and U6326 (N_6326,N_4007,N_4189);
nor U6327 (N_6327,N_3331,N_2632);
nand U6328 (N_6328,N_4209,N_4245);
nor U6329 (N_6329,N_4120,N_4952);
nor U6330 (N_6330,N_4551,N_4508);
and U6331 (N_6331,N_3268,N_4688);
or U6332 (N_6332,N_2879,N_3461);
or U6333 (N_6333,N_3639,N_3203);
or U6334 (N_6334,N_3445,N_4136);
and U6335 (N_6335,N_3889,N_2859);
or U6336 (N_6336,N_2694,N_3367);
nor U6337 (N_6337,N_2977,N_4303);
and U6338 (N_6338,N_3174,N_3996);
nor U6339 (N_6339,N_4350,N_4689);
or U6340 (N_6340,N_4592,N_4232);
and U6341 (N_6341,N_3058,N_4076);
and U6342 (N_6342,N_3099,N_3601);
and U6343 (N_6343,N_2676,N_4906);
nor U6344 (N_6344,N_4877,N_4376);
or U6345 (N_6345,N_3791,N_4243);
nor U6346 (N_6346,N_3237,N_4098);
or U6347 (N_6347,N_2504,N_3661);
or U6348 (N_6348,N_4400,N_3634);
nor U6349 (N_6349,N_3493,N_3288);
nand U6350 (N_6350,N_2731,N_4375);
nand U6351 (N_6351,N_2898,N_4348);
nor U6352 (N_6352,N_4250,N_3102);
or U6353 (N_6353,N_2852,N_2605);
nor U6354 (N_6354,N_4625,N_2927);
nor U6355 (N_6355,N_4466,N_3231);
nor U6356 (N_6356,N_3270,N_4666);
or U6357 (N_6357,N_4296,N_4167);
nor U6358 (N_6358,N_3693,N_4969);
nor U6359 (N_6359,N_3770,N_4079);
or U6360 (N_6360,N_4338,N_4740);
nand U6361 (N_6361,N_3191,N_3259);
or U6362 (N_6362,N_4110,N_4336);
or U6363 (N_6363,N_2541,N_2746);
and U6364 (N_6364,N_3622,N_3104);
and U6365 (N_6365,N_4969,N_4814);
and U6366 (N_6366,N_4418,N_3487);
nand U6367 (N_6367,N_3710,N_4340);
nor U6368 (N_6368,N_4753,N_4951);
nor U6369 (N_6369,N_3445,N_4007);
nor U6370 (N_6370,N_4512,N_3152);
nor U6371 (N_6371,N_2922,N_4085);
nand U6372 (N_6372,N_3803,N_3229);
and U6373 (N_6373,N_3422,N_2545);
or U6374 (N_6374,N_3162,N_4014);
or U6375 (N_6375,N_2999,N_4122);
or U6376 (N_6376,N_3585,N_4327);
nand U6377 (N_6377,N_4849,N_3437);
or U6378 (N_6378,N_3697,N_2644);
nand U6379 (N_6379,N_2789,N_4917);
xor U6380 (N_6380,N_4225,N_3918);
or U6381 (N_6381,N_3657,N_3660);
nand U6382 (N_6382,N_3627,N_4566);
nor U6383 (N_6383,N_3152,N_4994);
nor U6384 (N_6384,N_3038,N_4598);
or U6385 (N_6385,N_3668,N_4046);
nor U6386 (N_6386,N_2976,N_3744);
or U6387 (N_6387,N_4469,N_3201);
nor U6388 (N_6388,N_3886,N_4628);
and U6389 (N_6389,N_2804,N_3596);
or U6390 (N_6390,N_4768,N_3176);
nor U6391 (N_6391,N_3395,N_2849);
nand U6392 (N_6392,N_3938,N_4079);
nor U6393 (N_6393,N_3568,N_2830);
nor U6394 (N_6394,N_3019,N_3881);
and U6395 (N_6395,N_4750,N_3540);
and U6396 (N_6396,N_4624,N_4050);
nand U6397 (N_6397,N_3535,N_4856);
and U6398 (N_6398,N_2515,N_2875);
or U6399 (N_6399,N_3249,N_3007);
nor U6400 (N_6400,N_3823,N_3013);
nor U6401 (N_6401,N_4621,N_4644);
or U6402 (N_6402,N_2754,N_2617);
and U6403 (N_6403,N_2759,N_4772);
or U6404 (N_6404,N_2935,N_3178);
or U6405 (N_6405,N_3357,N_4357);
or U6406 (N_6406,N_3332,N_4972);
nor U6407 (N_6407,N_3750,N_3023);
or U6408 (N_6408,N_3106,N_2724);
nand U6409 (N_6409,N_4874,N_3660);
and U6410 (N_6410,N_2676,N_3151);
nand U6411 (N_6411,N_4577,N_4007);
or U6412 (N_6412,N_2749,N_4918);
nor U6413 (N_6413,N_3477,N_3003);
nor U6414 (N_6414,N_4532,N_4088);
xnor U6415 (N_6415,N_4372,N_4899);
nand U6416 (N_6416,N_3570,N_4933);
or U6417 (N_6417,N_3779,N_3346);
nor U6418 (N_6418,N_3458,N_4784);
nand U6419 (N_6419,N_3397,N_4661);
and U6420 (N_6420,N_4562,N_4869);
nand U6421 (N_6421,N_3161,N_3999);
nor U6422 (N_6422,N_3617,N_3633);
or U6423 (N_6423,N_2536,N_2769);
nor U6424 (N_6424,N_4451,N_3361);
nor U6425 (N_6425,N_4329,N_2815);
or U6426 (N_6426,N_4294,N_4401);
or U6427 (N_6427,N_4203,N_4849);
and U6428 (N_6428,N_3847,N_3933);
nand U6429 (N_6429,N_4802,N_4312);
nor U6430 (N_6430,N_3117,N_4401);
and U6431 (N_6431,N_4112,N_3847);
nand U6432 (N_6432,N_4025,N_3248);
or U6433 (N_6433,N_2974,N_3961);
or U6434 (N_6434,N_4602,N_4072);
or U6435 (N_6435,N_4345,N_4308);
or U6436 (N_6436,N_4336,N_4905);
nand U6437 (N_6437,N_3158,N_3810);
nor U6438 (N_6438,N_3941,N_3286);
nand U6439 (N_6439,N_3113,N_4862);
and U6440 (N_6440,N_3245,N_3432);
and U6441 (N_6441,N_4334,N_4617);
or U6442 (N_6442,N_4571,N_2563);
nor U6443 (N_6443,N_3066,N_3484);
nor U6444 (N_6444,N_3721,N_3291);
and U6445 (N_6445,N_4200,N_4760);
nand U6446 (N_6446,N_4534,N_4510);
and U6447 (N_6447,N_3636,N_3819);
nand U6448 (N_6448,N_4466,N_3614);
nor U6449 (N_6449,N_3340,N_4539);
nand U6450 (N_6450,N_4421,N_4700);
or U6451 (N_6451,N_4789,N_3447);
or U6452 (N_6452,N_4736,N_3827);
nand U6453 (N_6453,N_4600,N_3903);
nor U6454 (N_6454,N_4692,N_2914);
and U6455 (N_6455,N_3253,N_2667);
or U6456 (N_6456,N_3804,N_2632);
or U6457 (N_6457,N_2768,N_2619);
nand U6458 (N_6458,N_4992,N_4013);
nor U6459 (N_6459,N_3337,N_4619);
nor U6460 (N_6460,N_3156,N_4520);
nor U6461 (N_6461,N_3004,N_3824);
nor U6462 (N_6462,N_4485,N_3068);
or U6463 (N_6463,N_4380,N_2985);
nand U6464 (N_6464,N_3980,N_4660);
and U6465 (N_6465,N_3155,N_2531);
nor U6466 (N_6466,N_3185,N_4034);
and U6467 (N_6467,N_2564,N_3383);
nor U6468 (N_6468,N_3912,N_4780);
nand U6469 (N_6469,N_3816,N_4515);
nand U6470 (N_6470,N_3040,N_4255);
nand U6471 (N_6471,N_3422,N_4938);
nand U6472 (N_6472,N_2882,N_3936);
nand U6473 (N_6473,N_3017,N_4170);
nand U6474 (N_6474,N_4477,N_3690);
or U6475 (N_6475,N_3588,N_4984);
nand U6476 (N_6476,N_2706,N_4868);
or U6477 (N_6477,N_3533,N_4513);
or U6478 (N_6478,N_3861,N_3855);
nor U6479 (N_6479,N_4533,N_4238);
or U6480 (N_6480,N_4439,N_2633);
nand U6481 (N_6481,N_2576,N_3706);
nor U6482 (N_6482,N_3459,N_4858);
nand U6483 (N_6483,N_4116,N_4636);
nand U6484 (N_6484,N_4923,N_3435);
nand U6485 (N_6485,N_3402,N_3482);
and U6486 (N_6486,N_3735,N_2587);
nor U6487 (N_6487,N_4427,N_2941);
and U6488 (N_6488,N_3723,N_2647);
or U6489 (N_6489,N_4398,N_3246);
and U6490 (N_6490,N_3455,N_3422);
nand U6491 (N_6491,N_3708,N_3695);
and U6492 (N_6492,N_2971,N_4389);
nand U6493 (N_6493,N_4671,N_3383);
or U6494 (N_6494,N_4133,N_4481);
or U6495 (N_6495,N_3150,N_2802);
nand U6496 (N_6496,N_4395,N_3262);
or U6497 (N_6497,N_4562,N_2956);
nor U6498 (N_6498,N_2547,N_4078);
nor U6499 (N_6499,N_3262,N_2700);
nor U6500 (N_6500,N_3702,N_2850);
and U6501 (N_6501,N_4545,N_2504);
or U6502 (N_6502,N_3046,N_3302);
nor U6503 (N_6503,N_4412,N_4116);
nor U6504 (N_6504,N_4605,N_4256);
nand U6505 (N_6505,N_4989,N_4675);
or U6506 (N_6506,N_4359,N_3544);
and U6507 (N_6507,N_4007,N_3113);
or U6508 (N_6508,N_4061,N_3588);
or U6509 (N_6509,N_4884,N_3165);
nand U6510 (N_6510,N_2846,N_3941);
nand U6511 (N_6511,N_3854,N_3931);
and U6512 (N_6512,N_2636,N_4774);
nand U6513 (N_6513,N_2654,N_3083);
and U6514 (N_6514,N_3216,N_2921);
nor U6515 (N_6515,N_4111,N_3109);
nor U6516 (N_6516,N_2599,N_4580);
and U6517 (N_6517,N_4818,N_3281);
nor U6518 (N_6518,N_3886,N_3852);
nand U6519 (N_6519,N_2693,N_4477);
nor U6520 (N_6520,N_2850,N_2863);
and U6521 (N_6521,N_4635,N_4165);
and U6522 (N_6522,N_2633,N_2567);
nand U6523 (N_6523,N_3417,N_4734);
or U6524 (N_6524,N_4885,N_4167);
or U6525 (N_6525,N_4599,N_2806);
and U6526 (N_6526,N_2694,N_3709);
and U6527 (N_6527,N_4245,N_4057);
xnor U6528 (N_6528,N_4919,N_3486);
nand U6529 (N_6529,N_3774,N_3141);
or U6530 (N_6530,N_3150,N_3830);
xnor U6531 (N_6531,N_4937,N_2683);
nor U6532 (N_6532,N_3540,N_4066);
or U6533 (N_6533,N_2658,N_3386);
nand U6534 (N_6534,N_4360,N_4150);
and U6535 (N_6535,N_2715,N_2672);
nand U6536 (N_6536,N_3305,N_3890);
and U6537 (N_6537,N_4806,N_4431);
nor U6538 (N_6538,N_3005,N_4095);
nor U6539 (N_6539,N_3549,N_4842);
nor U6540 (N_6540,N_4559,N_3996);
nand U6541 (N_6541,N_3433,N_3116);
nor U6542 (N_6542,N_4889,N_3905);
or U6543 (N_6543,N_3878,N_3469);
nand U6544 (N_6544,N_4970,N_4900);
nor U6545 (N_6545,N_4231,N_3945);
nand U6546 (N_6546,N_3021,N_3465);
nor U6547 (N_6547,N_3820,N_2677);
nand U6548 (N_6548,N_3797,N_2522);
and U6549 (N_6549,N_3670,N_4178);
nor U6550 (N_6550,N_4262,N_4546);
and U6551 (N_6551,N_4409,N_3804);
nand U6552 (N_6552,N_4841,N_4329);
or U6553 (N_6553,N_3380,N_3007);
nand U6554 (N_6554,N_3132,N_3818);
and U6555 (N_6555,N_2900,N_4922);
and U6556 (N_6556,N_4255,N_4462);
or U6557 (N_6557,N_3184,N_4154);
and U6558 (N_6558,N_3604,N_4508);
nor U6559 (N_6559,N_3886,N_3296);
or U6560 (N_6560,N_4423,N_3331);
nor U6561 (N_6561,N_3138,N_3216);
nand U6562 (N_6562,N_3458,N_3569);
nand U6563 (N_6563,N_4622,N_3514);
nor U6564 (N_6564,N_2767,N_2983);
nand U6565 (N_6565,N_3191,N_4816);
and U6566 (N_6566,N_4565,N_4122);
xor U6567 (N_6567,N_4358,N_2883);
and U6568 (N_6568,N_3416,N_4789);
nor U6569 (N_6569,N_3091,N_3684);
nand U6570 (N_6570,N_4916,N_3353);
nand U6571 (N_6571,N_3026,N_3070);
nand U6572 (N_6572,N_4498,N_3030);
and U6573 (N_6573,N_3187,N_3722);
and U6574 (N_6574,N_3453,N_4901);
or U6575 (N_6575,N_3306,N_4628);
and U6576 (N_6576,N_4078,N_3021);
and U6577 (N_6577,N_3118,N_4527);
nand U6578 (N_6578,N_3669,N_2910);
and U6579 (N_6579,N_4886,N_4967);
xor U6580 (N_6580,N_2926,N_4690);
nand U6581 (N_6581,N_4420,N_3414);
or U6582 (N_6582,N_3580,N_4080);
nand U6583 (N_6583,N_2920,N_4191);
nor U6584 (N_6584,N_2598,N_4044);
nand U6585 (N_6585,N_4904,N_3765);
and U6586 (N_6586,N_2641,N_2606);
nor U6587 (N_6587,N_4208,N_4223);
nand U6588 (N_6588,N_4067,N_3271);
and U6589 (N_6589,N_4540,N_2783);
and U6590 (N_6590,N_2657,N_4859);
nor U6591 (N_6591,N_4076,N_4902);
nand U6592 (N_6592,N_3987,N_2636);
or U6593 (N_6593,N_3258,N_3690);
or U6594 (N_6594,N_2626,N_4977);
or U6595 (N_6595,N_3512,N_3228);
and U6596 (N_6596,N_4547,N_4484);
and U6597 (N_6597,N_4544,N_4666);
or U6598 (N_6598,N_4462,N_4782);
nor U6599 (N_6599,N_4172,N_2872);
nor U6600 (N_6600,N_3364,N_3150);
nand U6601 (N_6601,N_3555,N_3314);
nor U6602 (N_6602,N_3586,N_3990);
nor U6603 (N_6603,N_4319,N_4075);
or U6604 (N_6604,N_3823,N_3716);
and U6605 (N_6605,N_4352,N_3271);
nor U6606 (N_6606,N_4574,N_3528);
nor U6607 (N_6607,N_2944,N_4244);
nor U6608 (N_6608,N_3451,N_3152);
nor U6609 (N_6609,N_3157,N_4007);
nor U6610 (N_6610,N_3150,N_2533);
and U6611 (N_6611,N_4056,N_3828);
nor U6612 (N_6612,N_2763,N_3629);
or U6613 (N_6613,N_4650,N_3144);
or U6614 (N_6614,N_3638,N_2967);
xnor U6615 (N_6615,N_3223,N_4777);
or U6616 (N_6616,N_4662,N_4285);
nand U6617 (N_6617,N_4960,N_4540);
nand U6618 (N_6618,N_3535,N_2805);
nor U6619 (N_6619,N_3840,N_4356);
and U6620 (N_6620,N_4378,N_4256);
nand U6621 (N_6621,N_4018,N_4979);
nor U6622 (N_6622,N_4269,N_4536);
nor U6623 (N_6623,N_2660,N_3294);
nand U6624 (N_6624,N_3424,N_4006);
and U6625 (N_6625,N_4410,N_2731);
or U6626 (N_6626,N_3271,N_2830);
and U6627 (N_6627,N_4547,N_2743);
or U6628 (N_6628,N_3940,N_3490);
or U6629 (N_6629,N_4997,N_2896);
and U6630 (N_6630,N_3220,N_3444);
and U6631 (N_6631,N_2975,N_3089);
or U6632 (N_6632,N_3207,N_4807);
nor U6633 (N_6633,N_3501,N_3790);
nor U6634 (N_6634,N_2850,N_4324);
nor U6635 (N_6635,N_3171,N_3121);
and U6636 (N_6636,N_3744,N_4526);
nand U6637 (N_6637,N_4011,N_4077);
nor U6638 (N_6638,N_3164,N_4332);
nor U6639 (N_6639,N_2729,N_2547);
or U6640 (N_6640,N_3098,N_4141);
and U6641 (N_6641,N_4280,N_4553);
nor U6642 (N_6642,N_3217,N_2717);
or U6643 (N_6643,N_4895,N_3145);
nand U6644 (N_6644,N_3026,N_4934);
and U6645 (N_6645,N_4137,N_4887);
nand U6646 (N_6646,N_2735,N_2693);
or U6647 (N_6647,N_3935,N_4118);
nand U6648 (N_6648,N_4074,N_3645);
nor U6649 (N_6649,N_3323,N_4510);
nor U6650 (N_6650,N_3640,N_3412);
and U6651 (N_6651,N_4782,N_3680);
or U6652 (N_6652,N_4070,N_3172);
nor U6653 (N_6653,N_3773,N_3500);
nand U6654 (N_6654,N_2928,N_4534);
or U6655 (N_6655,N_3064,N_4249);
nor U6656 (N_6656,N_4593,N_3462);
nand U6657 (N_6657,N_3539,N_4389);
and U6658 (N_6658,N_3946,N_4443);
nand U6659 (N_6659,N_2676,N_3993);
and U6660 (N_6660,N_3440,N_4308);
or U6661 (N_6661,N_4238,N_4022);
nor U6662 (N_6662,N_3733,N_4587);
nand U6663 (N_6663,N_3916,N_2805);
nor U6664 (N_6664,N_4035,N_3236);
and U6665 (N_6665,N_4047,N_4275);
and U6666 (N_6666,N_4722,N_2737);
nand U6667 (N_6667,N_4775,N_3294);
or U6668 (N_6668,N_3410,N_4519);
nand U6669 (N_6669,N_2957,N_4959);
or U6670 (N_6670,N_3898,N_4046);
or U6671 (N_6671,N_3781,N_4832);
and U6672 (N_6672,N_3874,N_3064);
and U6673 (N_6673,N_4477,N_2758);
nand U6674 (N_6674,N_4447,N_3989);
nand U6675 (N_6675,N_3659,N_2563);
nand U6676 (N_6676,N_2858,N_4192);
nand U6677 (N_6677,N_3526,N_4372);
or U6678 (N_6678,N_2991,N_2899);
nand U6679 (N_6679,N_4707,N_3116);
nor U6680 (N_6680,N_2861,N_4356);
nor U6681 (N_6681,N_3940,N_4966);
and U6682 (N_6682,N_3421,N_2772);
and U6683 (N_6683,N_3448,N_4154);
or U6684 (N_6684,N_3267,N_4413);
and U6685 (N_6685,N_4014,N_4397);
nor U6686 (N_6686,N_3530,N_3031);
nand U6687 (N_6687,N_3589,N_2857);
nand U6688 (N_6688,N_3009,N_4508);
or U6689 (N_6689,N_3981,N_4106);
or U6690 (N_6690,N_4008,N_3025);
and U6691 (N_6691,N_3025,N_4490);
nor U6692 (N_6692,N_4762,N_4288);
or U6693 (N_6693,N_3944,N_4575);
and U6694 (N_6694,N_4627,N_3556);
nor U6695 (N_6695,N_4728,N_4053);
and U6696 (N_6696,N_3260,N_4557);
and U6697 (N_6697,N_4577,N_2834);
nor U6698 (N_6698,N_4042,N_2523);
nor U6699 (N_6699,N_3821,N_3603);
nor U6700 (N_6700,N_4457,N_3607);
and U6701 (N_6701,N_2911,N_4022);
nand U6702 (N_6702,N_2571,N_2671);
nor U6703 (N_6703,N_3367,N_3071);
nand U6704 (N_6704,N_3581,N_4649);
or U6705 (N_6705,N_3853,N_4576);
nand U6706 (N_6706,N_4680,N_3108);
xor U6707 (N_6707,N_3757,N_2660);
or U6708 (N_6708,N_4769,N_3579);
xnor U6709 (N_6709,N_4796,N_2641);
nor U6710 (N_6710,N_3211,N_3320);
nor U6711 (N_6711,N_4579,N_3372);
nand U6712 (N_6712,N_3548,N_4726);
nand U6713 (N_6713,N_2906,N_4377);
or U6714 (N_6714,N_4154,N_4224);
nor U6715 (N_6715,N_4822,N_3501);
and U6716 (N_6716,N_4605,N_4040);
or U6717 (N_6717,N_4010,N_3983);
nor U6718 (N_6718,N_3044,N_2880);
or U6719 (N_6719,N_3188,N_2978);
or U6720 (N_6720,N_3054,N_4507);
and U6721 (N_6721,N_4003,N_4721);
or U6722 (N_6722,N_4978,N_4350);
nor U6723 (N_6723,N_3571,N_3467);
or U6724 (N_6724,N_3889,N_3546);
or U6725 (N_6725,N_2653,N_4332);
nor U6726 (N_6726,N_3227,N_4893);
or U6727 (N_6727,N_3012,N_2822);
nor U6728 (N_6728,N_2940,N_3852);
nand U6729 (N_6729,N_2765,N_2881);
or U6730 (N_6730,N_3883,N_4577);
and U6731 (N_6731,N_2578,N_4320);
nand U6732 (N_6732,N_4989,N_3677);
and U6733 (N_6733,N_4620,N_2939);
or U6734 (N_6734,N_4649,N_2714);
nand U6735 (N_6735,N_4342,N_4481);
or U6736 (N_6736,N_3714,N_3371);
and U6737 (N_6737,N_3664,N_4082);
and U6738 (N_6738,N_3315,N_2571);
nor U6739 (N_6739,N_4685,N_3584);
nor U6740 (N_6740,N_3486,N_4283);
and U6741 (N_6741,N_2648,N_3792);
or U6742 (N_6742,N_2735,N_3294);
and U6743 (N_6743,N_4007,N_4667);
nor U6744 (N_6744,N_2776,N_3731);
and U6745 (N_6745,N_3981,N_3369);
xor U6746 (N_6746,N_3267,N_4674);
and U6747 (N_6747,N_2546,N_2896);
and U6748 (N_6748,N_4489,N_2840);
nor U6749 (N_6749,N_3250,N_3814);
and U6750 (N_6750,N_4126,N_2940);
nand U6751 (N_6751,N_4313,N_4723);
and U6752 (N_6752,N_3241,N_3130);
xnor U6753 (N_6753,N_4044,N_2773);
or U6754 (N_6754,N_3476,N_4034);
nor U6755 (N_6755,N_3278,N_4846);
and U6756 (N_6756,N_2547,N_2541);
and U6757 (N_6757,N_3691,N_4115);
or U6758 (N_6758,N_3696,N_4727);
nor U6759 (N_6759,N_4627,N_2906);
and U6760 (N_6760,N_3599,N_2837);
or U6761 (N_6761,N_2683,N_3754);
nor U6762 (N_6762,N_2926,N_3363);
nor U6763 (N_6763,N_4198,N_4872);
nand U6764 (N_6764,N_4799,N_4772);
nor U6765 (N_6765,N_4129,N_4978);
and U6766 (N_6766,N_4402,N_3157);
nor U6767 (N_6767,N_3575,N_3132);
and U6768 (N_6768,N_4232,N_4901);
nor U6769 (N_6769,N_3148,N_2870);
nor U6770 (N_6770,N_2685,N_3396);
nor U6771 (N_6771,N_3728,N_4445);
or U6772 (N_6772,N_2951,N_3945);
nand U6773 (N_6773,N_3298,N_4031);
nor U6774 (N_6774,N_3907,N_3359);
nand U6775 (N_6775,N_4234,N_4896);
or U6776 (N_6776,N_3494,N_3162);
nor U6777 (N_6777,N_3390,N_3504);
or U6778 (N_6778,N_4356,N_3040);
nand U6779 (N_6779,N_4056,N_4963);
or U6780 (N_6780,N_4095,N_3077);
or U6781 (N_6781,N_3064,N_3633);
or U6782 (N_6782,N_4445,N_2649);
or U6783 (N_6783,N_4573,N_4342);
and U6784 (N_6784,N_4992,N_3945);
nand U6785 (N_6785,N_4326,N_3586);
or U6786 (N_6786,N_4954,N_3514);
nor U6787 (N_6787,N_2863,N_3332);
nand U6788 (N_6788,N_4030,N_3625);
or U6789 (N_6789,N_4604,N_3540);
or U6790 (N_6790,N_4207,N_4422);
nand U6791 (N_6791,N_4817,N_3667);
and U6792 (N_6792,N_3762,N_3724);
and U6793 (N_6793,N_4944,N_4621);
or U6794 (N_6794,N_3267,N_3077);
and U6795 (N_6795,N_4464,N_2729);
and U6796 (N_6796,N_4754,N_4979);
nor U6797 (N_6797,N_4940,N_2511);
nand U6798 (N_6798,N_3616,N_3159);
or U6799 (N_6799,N_3037,N_4738);
nor U6800 (N_6800,N_4468,N_2954);
and U6801 (N_6801,N_2535,N_4725);
nor U6802 (N_6802,N_3228,N_4947);
nand U6803 (N_6803,N_3812,N_2568);
or U6804 (N_6804,N_4515,N_3783);
or U6805 (N_6805,N_4590,N_4456);
and U6806 (N_6806,N_4265,N_2674);
nor U6807 (N_6807,N_3461,N_3397);
nand U6808 (N_6808,N_3089,N_3259);
and U6809 (N_6809,N_2893,N_3531);
nor U6810 (N_6810,N_4591,N_3338);
and U6811 (N_6811,N_4509,N_4417);
nor U6812 (N_6812,N_3202,N_3826);
or U6813 (N_6813,N_3940,N_2937);
or U6814 (N_6814,N_4157,N_3436);
nor U6815 (N_6815,N_4030,N_4093);
nor U6816 (N_6816,N_4669,N_3581);
nand U6817 (N_6817,N_4077,N_3601);
or U6818 (N_6818,N_4210,N_3688);
nor U6819 (N_6819,N_4944,N_2853);
xor U6820 (N_6820,N_4167,N_2825);
and U6821 (N_6821,N_2742,N_4034);
and U6822 (N_6822,N_3722,N_4831);
or U6823 (N_6823,N_4557,N_3917);
nor U6824 (N_6824,N_3255,N_4589);
nor U6825 (N_6825,N_4358,N_3896);
nor U6826 (N_6826,N_3972,N_3952);
nand U6827 (N_6827,N_4829,N_2809);
nand U6828 (N_6828,N_2962,N_2903);
or U6829 (N_6829,N_4199,N_2991);
nand U6830 (N_6830,N_4361,N_2979);
nand U6831 (N_6831,N_4166,N_3316);
nand U6832 (N_6832,N_3599,N_4797);
nor U6833 (N_6833,N_4018,N_3283);
or U6834 (N_6834,N_2555,N_4048);
nand U6835 (N_6835,N_3605,N_2666);
or U6836 (N_6836,N_3899,N_4759);
or U6837 (N_6837,N_2918,N_4777);
or U6838 (N_6838,N_3294,N_4405);
or U6839 (N_6839,N_4509,N_3493);
nand U6840 (N_6840,N_3164,N_3875);
nand U6841 (N_6841,N_4645,N_4408);
and U6842 (N_6842,N_4107,N_3715);
nand U6843 (N_6843,N_3836,N_4263);
nand U6844 (N_6844,N_3794,N_3104);
nor U6845 (N_6845,N_4569,N_3376);
nand U6846 (N_6846,N_3398,N_4874);
and U6847 (N_6847,N_3868,N_2763);
and U6848 (N_6848,N_3141,N_4189);
nor U6849 (N_6849,N_3611,N_4880);
or U6850 (N_6850,N_3003,N_3008);
or U6851 (N_6851,N_4232,N_4745);
nor U6852 (N_6852,N_4308,N_4342);
nor U6853 (N_6853,N_4707,N_4176);
or U6854 (N_6854,N_4651,N_4105);
and U6855 (N_6855,N_3676,N_4003);
xor U6856 (N_6856,N_4834,N_3323);
or U6857 (N_6857,N_4433,N_3003);
and U6858 (N_6858,N_2724,N_3079);
nand U6859 (N_6859,N_2583,N_4534);
xor U6860 (N_6860,N_4296,N_4102);
nand U6861 (N_6861,N_4378,N_3835);
nand U6862 (N_6862,N_3614,N_3144);
or U6863 (N_6863,N_2825,N_3699);
nand U6864 (N_6864,N_2762,N_2562);
or U6865 (N_6865,N_4178,N_4045);
nand U6866 (N_6866,N_2639,N_3222);
nor U6867 (N_6867,N_2910,N_3797);
nand U6868 (N_6868,N_4712,N_4307);
nor U6869 (N_6869,N_4947,N_2883);
or U6870 (N_6870,N_2737,N_2899);
nor U6871 (N_6871,N_3519,N_4268);
or U6872 (N_6872,N_4146,N_2551);
nor U6873 (N_6873,N_2670,N_4772);
and U6874 (N_6874,N_3552,N_3575);
or U6875 (N_6875,N_2675,N_3652);
nor U6876 (N_6876,N_3701,N_3987);
or U6877 (N_6877,N_4228,N_3077);
nor U6878 (N_6878,N_3863,N_3634);
nand U6879 (N_6879,N_4226,N_3684);
nor U6880 (N_6880,N_4927,N_3419);
or U6881 (N_6881,N_4679,N_4745);
nand U6882 (N_6882,N_4618,N_3563);
or U6883 (N_6883,N_4585,N_4796);
nor U6884 (N_6884,N_3566,N_4102);
nor U6885 (N_6885,N_3017,N_3692);
nand U6886 (N_6886,N_4175,N_3714);
nand U6887 (N_6887,N_2615,N_2981);
xor U6888 (N_6888,N_2695,N_4529);
or U6889 (N_6889,N_3695,N_4093);
nand U6890 (N_6890,N_2758,N_3315);
nor U6891 (N_6891,N_4935,N_4927);
and U6892 (N_6892,N_4077,N_4146);
nor U6893 (N_6893,N_3870,N_2919);
nor U6894 (N_6894,N_3685,N_3444);
or U6895 (N_6895,N_3596,N_4652);
or U6896 (N_6896,N_2547,N_3002);
nor U6897 (N_6897,N_3022,N_4150);
nor U6898 (N_6898,N_3979,N_2969);
nand U6899 (N_6899,N_4017,N_4475);
nor U6900 (N_6900,N_3947,N_3518);
nand U6901 (N_6901,N_3844,N_4296);
and U6902 (N_6902,N_4464,N_3314);
nand U6903 (N_6903,N_4292,N_4045);
nand U6904 (N_6904,N_3916,N_3688);
and U6905 (N_6905,N_4484,N_3626);
nor U6906 (N_6906,N_3645,N_3987);
and U6907 (N_6907,N_2991,N_4404);
nand U6908 (N_6908,N_4429,N_3237);
nor U6909 (N_6909,N_4968,N_4240);
or U6910 (N_6910,N_3136,N_4140);
nor U6911 (N_6911,N_3205,N_3468);
or U6912 (N_6912,N_4342,N_3435);
nor U6913 (N_6913,N_3022,N_4326);
or U6914 (N_6914,N_3417,N_4706);
nand U6915 (N_6915,N_3949,N_3062);
and U6916 (N_6916,N_4243,N_3151);
or U6917 (N_6917,N_2529,N_4947);
nor U6918 (N_6918,N_3301,N_2600);
nand U6919 (N_6919,N_4213,N_2688);
nand U6920 (N_6920,N_4929,N_2597);
and U6921 (N_6921,N_3692,N_4614);
nor U6922 (N_6922,N_4617,N_2835);
xor U6923 (N_6923,N_3405,N_3939);
nor U6924 (N_6924,N_3066,N_2981);
nor U6925 (N_6925,N_2889,N_4269);
nand U6926 (N_6926,N_3647,N_3277);
and U6927 (N_6927,N_3283,N_2529);
and U6928 (N_6928,N_2645,N_2644);
or U6929 (N_6929,N_3054,N_2649);
nand U6930 (N_6930,N_4111,N_3641);
or U6931 (N_6931,N_3784,N_3480);
nand U6932 (N_6932,N_4117,N_4933);
nand U6933 (N_6933,N_4098,N_4953);
and U6934 (N_6934,N_3702,N_4140);
nand U6935 (N_6935,N_2833,N_4178);
and U6936 (N_6936,N_2912,N_2512);
or U6937 (N_6937,N_4958,N_4378);
nor U6938 (N_6938,N_3820,N_3285);
nor U6939 (N_6939,N_3468,N_3214);
and U6940 (N_6940,N_3134,N_2933);
and U6941 (N_6941,N_4687,N_2704);
or U6942 (N_6942,N_3676,N_3084);
or U6943 (N_6943,N_3963,N_3748);
and U6944 (N_6944,N_3631,N_4424);
nor U6945 (N_6945,N_4370,N_2948);
or U6946 (N_6946,N_3517,N_4344);
nand U6947 (N_6947,N_4854,N_2911);
nand U6948 (N_6948,N_3038,N_4022);
or U6949 (N_6949,N_4948,N_4674);
nor U6950 (N_6950,N_4704,N_4173);
and U6951 (N_6951,N_3441,N_4856);
nand U6952 (N_6952,N_4910,N_2516);
nor U6953 (N_6953,N_3786,N_4737);
nand U6954 (N_6954,N_4635,N_4861);
nor U6955 (N_6955,N_4920,N_3785);
or U6956 (N_6956,N_2888,N_2571);
or U6957 (N_6957,N_3631,N_3376);
or U6958 (N_6958,N_3096,N_3543);
nand U6959 (N_6959,N_3964,N_3258);
nor U6960 (N_6960,N_2856,N_4250);
or U6961 (N_6961,N_4485,N_4100);
and U6962 (N_6962,N_3028,N_2737);
nor U6963 (N_6963,N_3499,N_3539);
nand U6964 (N_6964,N_3547,N_2780);
xor U6965 (N_6965,N_2589,N_3245);
nand U6966 (N_6966,N_4273,N_4800);
nor U6967 (N_6967,N_2570,N_4265);
nor U6968 (N_6968,N_4982,N_4643);
and U6969 (N_6969,N_2713,N_4640);
and U6970 (N_6970,N_3003,N_3838);
and U6971 (N_6971,N_3735,N_4191);
nor U6972 (N_6972,N_2515,N_2724);
nand U6973 (N_6973,N_2731,N_4196);
or U6974 (N_6974,N_4300,N_3203);
nand U6975 (N_6975,N_4085,N_4989);
nand U6976 (N_6976,N_2609,N_2810);
nand U6977 (N_6977,N_2598,N_4786);
or U6978 (N_6978,N_3946,N_3683);
nor U6979 (N_6979,N_2874,N_4936);
nor U6980 (N_6980,N_4127,N_3605);
xnor U6981 (N_6981,N_4567,N_2744);
or U6982 (N_6982,N_3945,N_3311);
and U6983 (N_6983,N_4743,N_2623);
and U6984 (N_6984,N_3682,N_3199);
and U6985 (N_6985,N_2921,N_2858);
nor U6986 (N_6986,N_4089,N_2768);
or U6987 (N_6987,N_4351,N_2783);
or U6988 (N_6988,N_2768,N_2525);
nor U6989 (N_6989,N_2957,N_3946);
nand U6990 (N_6990,N_3565,N_3806);
or U6991 (N_6991,N_4813,N_3991);
nor U6992 (N_6992,N_2829,N_3911);
nor U6993 (N_6993,N_3589,N_4635);
nand U6994 (N_6994,N_4033,N_2937);
xor U6995 (N_6995,N_4073,N_4507);
or U6996 (N_6996,N_3422,N_4860);
or U6997 (N_6997,N_4793,N_3655);
nor U6998 (N_6998,N_4569,N_3079);
and U6999 (N_6999,N_4081,N_4374);
and U7000 (N_7000,N_2802,N_3073);
or U7001 (N_7001,N_2760,N_4762);
and U7002 (N_7002,N_3075,N_4117);
nand U7003 (N_7003,N_3668,N_3899);
nor U7004 (N_7004,N_4010,N_4152);
or U7005 (N_7005,N_4703,N_4615);
and U7006 (N_7006,N_2825,N_4449);
or U7007 (N_7007,N_3650,N_4518);
and U7008 (N_7008,N_4545,N_3135);
nor U7009 (N_7009,N_2865,N_4105);
or U7010 (N_7010,N_4438,N_2769);
nand U7011 (N_7011,N_3954,N_4676);
or U7012 (N_7012,N_4425,N_2842);
nor U7013 (N_7013,N_3021,N_3295);
nor U7014 (N_7014,N_2742,N_2765);
and U7015 (N_7015,N_4496,N_4592);
nor U7016 (N_7016,N_4854,N_4237);
nand U7017 (N_7017,N_4760,N_4495);
nor U7018 (N_7018,N_3950,N_3178);
nor U7019 (N_7019,N_3815,N_4685);
nand U7020 (N_7020,N_4056,N_3014);
nand U7021 (N_7021,N_4262,N_3681);
nor U7022 (N_7022,N_3437,N_4290);
and U7023 (N_7023,N_3683,N_3100);
nand U7024 (N_7024,N_2836,N_2535);
and U7025 (N_7025,N_2627,N_4015);
and U7026 (N_7026,N_2734,N_4288);
nor U7027 (N_7027,N_4607,N_2826);
nand U7028 (N_7028,N_2517,N_4427);
or U7029 (N_7029,N_4338,N_4480);
or U7030 (N_7030,N_4328,N_3468);
and U7031 (N_7031,N_3940,N_3829);
nand U7032 (N_7032,N_2602,N_3213);
nor U7033 (N_7033,N_4091,N_4694);
or U7034 (N_7034,N_4346,N_4752);
nand U7035 (N_7035,N_4045,N_4495);
nor U7036 (N_7036,N_2685,N_2649);
nor U7037 (N_7037,N_4505,N_2791);
or U7038 (N_7038,N_4184,N_3097);
or U7039 (N_7039,N_2897,N_4655);
xor U7040 (N_7040,N_4192,N_4745);
or U7041 (N_7041,N_2812,N_3583);
nor U7042 (N_7042,N_4185,N_4397);
nand U7043 (N_7043,N_4369,N_4898);
and U7044 (N_7044,N_3449,N_4463);
and U7045 (N_7045,N_3791,N_4170);
or U7046 (N_7046,N_3881,N_2725);
and U7047 (N_7047,N_3936,N_2648);
nand U7048 (N_7048,N_2525,N_4554);
and U7049 (N_7049,N_3902,N_3252);
nor U7050 (N_7050,N_3696,N_3720);
or U7051 (N_7051,N_2513,N_3775);
or U7052 (N_7052,N_4659,N_3589);
or U7053 (N_7053,N_4674,N_4169);
xor U7054 (N_7054,N_2565,N_2659);
nor U7055 (N_7055,N_4559,N_2988);
and U7056 (N_7056,N_4210,N_3804);
nor U7057 (N_7057,N_4213,N_3700);
nand U7058 (N_7058,N_4487,N_4514);
nor U7059 (N_7059,N_4234,N_3347);
and U7060 (N_7060,N_3230,N_3879);
nor U7061 (N_7061,N_3719,N_3339);
or U7062 (N_7062,N_3144,N_4877);
and U7063 (N_7063,N_3095,N_3988);
and U7064 (N_7064,N_3374,N_2946);
and U7065 (N_7065,N_4190,N_4224);
nand U7066 (N_7066,N_4853,N_4588);
or U7067 (N_7067,N_2637,N_3302);
or U7068 (N_7068,N_4250,N_3896);
nand U7069 (N_7069,N_3547,N_2969);
nor U7070 (N_7070,N_3505,N_3230);
and U7071 (N_7071,N_3124,N_2855);
nand U7072 (N_7072,N_2702,N_3008);
or U7073 (N_7073,N_4126,N_3077);
or U7074 (N_7074,N_4217,N_2811);
nor U7075 (N_7075,N_2691,N_3024);
nor U7076 (N_7076,N_3460,N_4314);
nand U7077 (N_7077,N_2641,N_4845);
or U7078 (N_7078,N_3261,N_3686);
and U7079 (N_7079,N_2861,N_3571);
or U7080 (N_7080,N_4038,N_4789);
nor U7081 (N_7081,N_4542,N_3164);
and U7082 (N_7082,N_3379,N_4148);
or U7083 (N_7083,N_3404,N_2881);
nor U7084 (N_7084,N_2828,N_4538);
and U7085 (N_7085,N_3237,N_4818);
nand U7086 (N_7086,N_4277,N_2671);
nor U7087 (N_7087,N_4780,N_2732);
nor U7088 (N_7088,N_2596,N_4206);
xor U7089 (N_7089,N_4298,N_3803);
nand U7090 (N_7090,N_2908,N_4503);
nand U7091 (N_7091,N_2858,N_2501);
xnor U7092 (N_7092,N_3418,N_4497);
nor U7093 (N_7093,N_3093,N_4682);
and U7094 (N_7094,N_3779,N_3172);
or U7095 (N_7095,N_4222,N_4053);
nor U7096 (N_7096,N_4426,N_4440);
nor U7097 (N_7097,N_3431,N_3124);
nand U7098 (N_7098,N_3306,N_4007);
nand U7099 (N_7099,N_2664,N_2616);
nand U7100 (N_7100,N_4509,N_4004);
nand U7101 (N_7101,N_3062,N_4372);
or U7102 (N_7102,N_3917,N_2769);
or U7103 (N_7103,N_3041,N_4763);
nor U7104 (N_7104,N_4604,N_2997);
nor U7105 (N_7105,N_3151,N_2808);
or U7106 (N_7106,N_4915,N_2524);
nor U7107 (N_7107,N_3961,N_2829);
nor U7108 (N_7108,N_2605,N_2877);
and U7109 (N_7109,N_4579,N_4134);
nand U7110 (N_7110,N_3372,N_4143);
nand U7111 (N_7111,N_4436,N_3855);
or U7112 (N_7112,N_4520,N_4985);
and U7113 (N_7113,N_2871,N_2642);
nor U7114 (N_7114,N_3620,N_3542);
nor U7115 (N_7115,N_4819,N_2870);
nor U7116 (N_7116,N_4486,N_4278);
nand U7117 (N_7117,N_3417,N_2835);
or U7118 (N_7118,N_2850,N_4957);
or U7119 (N_7119,N_2805,N_2879);
nand U7120 (N_7120,N_4743,N_3059);
and U7121 (N_7121,N_3638,N_4958);
nor U7122 (N_7122,N_3376,N_4194);
nand U7123 (N_7123,N_4397,N_3802);
or U7124 (N_7124,N_3653,N_3389);
or U7125 (N_7125,N_3228,N_4942);
or U7126 (N_7126,N_3483,N_4762);
or U7127 (N_7127,N_3664,N_4417);
or U7128 (N_7128,N_3680,N_2584);
and U7129 (N_7129,N_2807,N_4585);
and U7130 (N_7130,N_4282,N_3993);
nand U7131 (N_7131,N_2862,N_3329);
and U7132 (N_7132,N_4292,N_3950);
nor U7133 (N_7133,N_4963,N_3725);
or U7134 (N_7134,N_3694,N_2929);
xor U7135 (N_7135,N_3117,N_3422);
nor U7136 (N_7136,N_4046,N_4954);
nor U7137 (N_7137,N_3865,N_4325);
nand U7138 (N_7138,N_2766,N_3779);
or U7139 (N_7139,N_3681,N_3378);
nand U7140 (N_7140,N_4130,N_4014);
or U7141 (N_7141,N_3168,N_2688);
and U7142 (N_7142,N_4926,N_4218);
and U7143 (N_7143,N_3461,N_2824);
or U7144 (N_7144,N_3714,N_3438);
and U7145 (N_7145,N_4319,N_3473);
and U7146 (N_7146,N_3310,N_3691);
or U7147 (N_7147,N_3782,N_3203);
and U7148 (N_7148,N_2760,N_3055);
and U7149 (N_7149,N_3653,N_2793);
nand U7150 (N_7150,N_4675,N_4950);
or U7151 (N_7151,N_4305,N_3370);
or U7152 (N_7152,N_4390,N_3126);
nand U7153 (N_7153,N_3980,N_3419);
and U7154 (N_7154,N_3648,N_4976);
nor U7155 (N_7155,N_2664,N_4401);
nand U7156 (N_7156,N_3412,N_3731);
or U7157 (N_7157,N_3186,N_4702);
and U7158 (N_7158,N_3707,N_4267);
and U7159 (N_7159,N_4195,N_2983);
or U7160 (N_7160,N_2544,N_4627);
or U7161 (N_7161,N_4196,N_3921);
and U7162 (N_7162,N_2658,N_2685);
nor U7163 (N_7163,N_4805,N_4095);
nor U7164 (N_7164,N_2589,N_4858);
nor U7165 (N_7165,N_4201,N_4572);
and U7166 (N_7166,N_2856,N_2746);
or U7167 (N_7167,N_4903,N_3346);
nor U7168 (N_7168,N_3155,N_3069);
or U7169 (N_7169,N_3257,N_4052);
and U7170 (N_7170,N_3868,N_3464);
or U7171 (N_7171,N_3095,N_3766);
nor U7172 (N_7172,N_4090,N_3638);
or U7173 (N_7173,N_2873,N_4485);
nor U7174 (N_7174,N_4904,N_3576);
and U7175 (N_7175,N_3388,N_4563);
and U7176 (N_7176,N_3139,N_3507);
and U7177 (N_7177,N_4573,N_3907);
and U7178 (N_7178,N_4477,N_4221);
nor U7179 (N_7179,N_4242,N_4646);
and U7180 (N_7180,N_4212,N_3545);
nand U7181 (N_7181,N_3373,N_3952);
nand U7182 (N_7182,N_3440,N_4584);
nand U7183 (N_7183,N_3967,N_4908);
or U7184 (N_7184,N_2958,N_4253);
and U7185 (N_7185,N_4617,N_3310);
or U7186 (N_7186,N_4858,N_3647);
nor U7187 (N_7187,N_4071,N_3515);
nor U7188 (N_7188,N_4128,N_4923);
or U7189 (N_7189,N_2822,N_4684);
or U7190 (N_7190,N_3477,N_3989);
nand U7191 (N_7191,N_2568,N_4548);
nor U7192 (N_7192,N_4768,N_3398);
and U7193 (N_7193,N_4855,N_2518);
and U7194 (N_7194,N_4678,N_4404);
nor U7195 (N_7195,N_3710,N_2803);
or U7196 (N_7196,N_4784,N_4638);
nand U7197 (N_7197,N_3309,N_2613);
nand U7198 (N_7198,N_4857,N_2740);
and U7199 (N_7199,N_4031,N_3641);
nand U7200 (N_7200,N_3317,N_3694);
nand U7201 (N_7201,N_2712,N_4192);
nor U7202 (N_7202,N_4144,N_2676);
nand U7203 (N_7203,N_4343,N_2892);
xor U7204 (N_7204,N_4961,N_3617);
or U7205 (N_7205,N_3205,N_3066);
or U7206 (N_7206,N_3897,N_4146);
nor U7207 (N_7207,N_4921,N_3309);
nor U7208 (N_7208,N_4139,N_3667);
and U7209 (N_7209,N_3187,N_4644);
xnor U7210 (N_7210,N_4685,N_2703);
nor U7211 (N_7211,N_4297,N_4248);
nor U7212 (N_7212,N_3752,N_2566);
nor U7213 (N_7213,N_4723,N_4179);
nand U7214 (N_7214,N_4341,N_4806);
or U7215 (N_7215,N_3064,N_4352);
and U7216 (N_7216,N_4610,N_3073);
nor U7217 (N_7217,N_2712,N_2825);
nand U7218 (N_7218,N_4148,N_4397);
or U7219 (N_7219,N_4979,N_3957);
nor U7220 (N_7220,N_4724,N_3672);
nor U7221 (N_7221,N_2571,N_2515);
or U7222 (N_7222,N_3603,N_4596);
and U7223 (N_7223,N_2872,N_4124);
nor U7224 (N_7224,N_2719,N_4935);
xor U7225 (N_7225,N_2852,N_3886);
and U7226 (N_7226,N_2640,N_3277);
nand U7227 (N_7227,N_3067,N_3126);
nand U7228 (N_7228,N_3506,N_3797);
nand U7229 (N_7229,N_3597,N_2645);
or U7230 (N_7230,N_4258,N_4112);
nor U7231 (N_7231,N_3206,N_4994);
xor U7232 (N_7232,N_4517,N_2748);
and U7233 (N_7233,N_4970,N_3971);
or U7234 (N_7234,N_4592,N_2937);
nor U7235 (N_7235,N_4282,N_4341);
nor U7236 (N_7236,N_4392,N_3014);
nand U7237 (N_7237,N_3353,N_3069);
and U7238 (N_7238,N_2569,N_3845);
and U7239 (N_7239,N_3643,N_3491);
and U7240 (N_7240,N_3961,N_2633);
nor U7241 (N_7241,N_4136,N_3515);
nand U7242 (N_7242,N_3432,N_3499);
and U7243 (N_7243,N_3315,N_4388);
nand U7244 (N_7244,N_3216,N_3967);
nor U7245 (N_7245,N_3130,N_3127);
nor U7246 (N_7246,N_2612,N_3252);
and U7247 (N_7247,N_3149,N_4434);
nor U7248 (N_7248,N_2782,N_3020);
and U7249 (N_7249,N_3111,N_4996);
and U7250 (N_7250,N_3693,N_3441);
nand U7251 (N_7251,N_2705,N_4851);
or U7252 (N_7252,N_4434,N_4404);
nand U7253 (N_7253,N_4754,N_3170);
xnor U7254 (N_7254,N_2527,N_2520);
or U7255 (N_7255,N_4158,N_4195);
nor U7256 (N_7256,N_3517,N_4588);
and U7257 (N_7257,N_2800,N_2552);
and U7258 (N_7258,N_3464,N_4845);
nor U7259 (N_7259,N_3365,N_3991);
and U7260 (N_7260,N_3871,N_2969);
or U7261 (N_7261,N_3858,N_2601);
nand U7262 (N_7262,N_2897,N_3155);
nand U7263 (N_7263,N_2853,N_4687);
or U7264 (N_7264,N_3990,N_3428);
nor U7265 (N_7265,N_4057,N_2859);
or U7266 (N_7266,N_4408,N_3411);
or U7267 (N_7267,N_4110,N_3874);
nor U7268 (N_7268,N_3887,N_4699);
and U7269 (N_7269,N_4406,N_2774);
nor U7270 (N_7270,N_2542,N_2570);
nor U7271 (N_7271,N_3406,N_3730);
and U7272 (N_7272,N_3729,N_4574);
or U7273 (N_7273,N_4922,N_3451);
nand U7274 (N_7274,N_4584,N_3744);
nor U7275 (N_7275,N_2896,N_4186);
and U7276 (N_7276,N_3103,N_4325);
and U7277 (N_7277,N_4933,N_2726);
or U7278 (N_7278,N_3501,N_4584);
nor U7279 (N_7279,N_4296,N_2575);
or U7280 (N_7280,N_3620,N_4876);
and U7281 (N_7281,N_3658,N_4234);
nand U7282 (N_7282,N_3628,N_4217);
and U7283 (N_7283,N_4167,N_4836);
and U7284 (N_7284,N_3235,N_3614);
or U7285 (N_7285,N_4399,N_2666);
nand U7286 (N_7286,N_4315,N_4565);
or U7287 (N_7287,N_3274,N_3100);
and U7288 (N_7288,N_3746,N_3058);
and U7289 (N_7289,N_3290,N_4266);
nand U7290 (N_7290,N_4932,N_4594);
nor U7291 (N_7291,N_3322,N_3344);
nor U7292 (N_7292,N_4587,N_3070);
and U7293 (N_7293,N_2622,N_2936);
nor U7294 (N_7294,N_2916,N_2747);
nand U7295 (N_7295,N_2867,N_3445);
nor U7296 (N_7296,N_4956,N_3580);
or U7297 (N_7297,N_4173,N_2509);
and U7298 (N_7298,N_4914,N_4970);
nand U7299 (N_7299,N_3247,N_4608);
or U7300 (N_7300,N_2897,N_4249);
xnor U7301 (N_7301,N_4707,N_2554);
and U7302 (N_7302,N_3534,N_4976);
nor U7303 (N_7303,N_4017,N_3023);
nand U7304 (N_7304,N_3189,N_4077);
and U7305 (N_7305,N_3202,N_4756);
or U7306 (N_7306,N_4964,N_4589);
and U7307 (N_7307,N_3609,N_3470);
and U7308 (N_7308,N_4170,N_3612);
and U7309 (N_7309,N_2632,N_3450);
and U7310 (N_7310,N_4401,N_4295);
nor U7311 (N_7311,N_4302,N_4777);
or U7312 (N_7312,N_3682,N_3224);
or U7313 (N_7313,N_2911,N_4416);
and U7314 (N_7314,N_4689,N_3316);
and U7315 (N_7315,N_3409,N_4606);
or U7316 (N_7316,N_3695,N_3164);
nor U7317 (N_7317,N_2879,N_4029);
nor U7318 (N_7318,N_4281,N_3237);
nand U7319 (N_7319,N_2949,N_2826);
and U7320 (N_7320,N_3279,N_3729);
nor U7321 (N_7321,N_2934,N_3361);
nand U7322 (N_7322,N_3196,N_2829);
nor U7323 (N_7323,N_2639,N_3202);
nor U7324 (N_7324,N_2908,N_3279);
nor U7325 (N_7325,N_4508,N_3677);
nor U7326 (N_7326,N_2760,N_4370);
and U7327 (N_7327,N_2992,N_3911);
nand U7328 (N_7328,N_4118,N_3912);
or U7329 (N_7329,N_3569,N_4335);
and U7330 (N_7330,N_4739,N_2503);
nor U7331 (N_7331,N_4993,N_2750);
nand U7332 (N_7332,N_2646,N_4622);
or U7333 (N_7333,N_4401,N_4221);
nand U7334 (N_7334,N_4600,N_3246);
nor U7335 (N_7335,N_3225,N_4039);
or U7336 (N_7336,N_3820,N_3099);
or U7337 (N_7337,N_2670,N_3071);
and U7338 (N_7338,N_3819,N_4319);
nor U7339 (N_7339,N_4279,N_4891);
or U7340 (N_7340,N_4180,N_4140);
or U7341 (N_7341,N_2792,N_3000);
nand U7342 (N_7342,N_3729,N_3359);
and U7343 (N_7343,N_3911,N_2983);
nand U7344 (N_7344,N_3405,N_2666);
nor U7345 (N_7345,N_3064,N_3718);
nand U7346 (N_7346,N_2722,N_3002);
or U7347 (N_7347,N_2522,N_3003);
or U7348 (N_7348,N_2924,N_3427);
xnor U7349 (N_7349,N_4970,N_3796);
and U7350 (N_7350,N_3695,N_3947);
nand U7351 (N_7351,N_3792,N_4667);
or U7352 (N_7352,N_3168,N_2956);
or U7353 (N_7353,N_2935,N_4047);
nor U7354 (N_7354,N_4029,N_2983);
nand U7355 (N_7355,N_3500,N_4043);
nand U7356 (N_7356,N_4166,N_4398);
or U7357 (N_7357,N_2500,N_4074);
and U7358 (N_7358,N_4624,N_2657);
or U7359 (N_7359,N_3125,N_4326);
nor U7360 (N_7360,N_4581,N_4315);
and U7361 (N_7361,N_3726,N_4389);
nand U7362 (N_7362,N_4319,N_4613);
nand U7363 (N_7363,N_3951,N_2580);
and U7364 (N_7364,N_3867,N_4688);
nand U7365 (N_7365,N_2678,N_3949);
nand U7366 (N_7366,N_4204,N_3063);
nand U7367 (N_7367,N_2588,N_2901);
or U7368 (N_7368,N_4357,N_2902);
and U7369 (N_7369,N_4267,N_3508);
and U7370 (N_7370,N_4975,N_3485);
or U7371 (N_7371,N_4909,N_2644);
or U7372 (N_7372,N_4164,N_3142);
nor U7373 (N_7373,N_4032,N_4881);
nand U7374 (N_7374,N_3905,N_4694);
nand U7375 (N_7375,N_3163,N_3927);
and U7376 (N_7376,N_4018,N_2678);
nand U7377 (N_7377,N_4315,N_2524);
or U7378 (N_7378,N_3997,N_2667);
nor U7379 (N_7379,N_2655,N_2850);
nor U7380 (N_7380,N_3137,N_3086);
nor U7381 (N_7381,N_4411,N_2875);
nor U7382 (N_7382,N_3101,N_3365);
or U7383 (N_7383,N_3446,N_4298);
nand U7384 (N_7384,N_3221,N_3208);
and U7385 (N_7385,N_4474,N_2693);
and U7386 (N_7386,N_3054,N_3461);
nand U7387 (N_7387,N_2899,N_3495);
or U7388 (N_7388,N_4371,N_3728);
nand U7389 (N_7389,N_3375,N_3472);
nor U7390 (N_7390,N_2644,N_4407);
or U7391 (N_7391,N_3867,N_3664);
nand U7392 (N_7392,N_3243,N_3535);
nor U7393 (N_7393,N_3480,N_2795);
nor U7394 (N_7394,N_4858,N_4336);
or U7395 (N_7395,N_4340,N_4095);
nor U7396 (N_7396,N_2582,N_3131);
or U7397 (N_7397,N_3333,N_3478);
nor U7398 (N_7398,N_3090,N_3759);
nand U7399 (N_7399,N_3403,N_3135);
nor U7400 (N_7400,N_3208,N_4062);
and U7401 (N_7401,N_4911,N_3549);
nor U7402 (N_7402,N_3722,N_2941);
or U7403 (N_7403,N_3486,N_2623);
and U7404 (N_7404,N_4653,N_2689);
and U7405 (N_7405,N_3103,N_3650);
nor U7406 (N_7406,N_4627,N_3499);
nor U7407 (N_7407,N_4646,N_2794);
and U7408 (N_7408,N_4775,N_4850);
nor U7409 (N_7409,N_3257,N_3343);
nor U7410 (N_7410,N_4013,N_3509);
or U7411 (N_7411,N_4268,N_2823);
nand U7412 (N_7412,N_4266,N_2666);
and U7413 (N_7413,N_4750,N_2761);
nand U7414 (N_7414,N_4230,N_2520);
or U7415 (N_7415,N_4725,N_4594);
and U7416 (N_7416,N_3181,N_4003);
and U7417 (N_7417,N_3314,N_2785);
or U7418 (N_7418,N_3355,N_3705);
nor U7419 (N_7419,N_3891,N_4115);
nor U7420 (N_7420,N_4069,N_3733);
xnor U7421 (N_7421,N_3227,N_4528);
nand U7422 (N_7422,N_2967,N_4747);
or U7423 (N_7423,N_4626,N_4826);
or U7424 (N_7424,N_3280,N_3235);
nor U7425 (N_7425,N_2867,N_2787);
nand U7426 (N_7426,N_4387,N_3611);
nand U7427 (N_7427,N_4988,N_4913);
and U7428 (N_7428,N_3296,N_2810);
or U7429 (N_7429,N_3862,N_2830);
nor U7430 (N_7430,N_3671,N_4664);
nor U7431 (N_7431,N_4266,N_4354);
or U7432 (N_7432,N_3914,N_3494);
and U7433 (N_7433,N_4274,N_4784);
or U7434 (N_7434,N_2749,N_4033);
xnor U7435 (N_7435,N_4196,N_3332);
or U7436 (N_7436,N_3785,N_3625);
nor U7437 (N_7437,N_4388,N_3401);
and U7438 (N_7438,N_3331,N_2932);
or U7439 (N_7439,N_3968,N_4360);
and U7440 (N_7440,N_3997,N_3738);
or U7441 (N_7441,N_3106,N_2685);
or U7442 (N_7442,N_2615,N_3562);
or U7443 (N_7443,N_3567,N_3674);
and U7444 (N_7444,N_4950,N_3989);
or U7445 (N_7445,N_2631,N_4920);
nor U7446 (N_7446,N_2830,N_4332);
nand U7447 (N_7447,N_4650,N_2668);
and U7448 (N_7448,N_4477,N_4824);
nor U7449 (N_7449,N_2567,N_2559);
or U7450 (N_7450,N_4847,N_4646);
and U7451 (N_7451,N_3751,N_3342);
nand U7452 (N_7452,N_3187,N_3517);
or U7453 (N_7453,N_3870,N_2968);
nor U7454 (N_7454,N_3675,N_3434);
and U7455 (N_7455,N_4402,N_3671);
nor U7456 (N_7456,N_3516,N_4101);
nand U7457 (N_7457,N_4027,N_3696);
nor U7458 (N_7458,N_4727,N_4284);
or U7459 (N_7459,N_2580,N_4938);
and U7460 (N_7460,N_3749,N_3921);
nor U7461 (N_7461,N_3404,N_2829);
or U7462 (N_7462,N_3072,N_2810);
nand U7463 (N_7463,N_4360,N_4875);
and U7464 (N_7464,N_2947,N_3281);
or U7465 (N_7465,N_3401,N_3851);
and U7466 (N_7466,N_3360,N_3536);
nand U7467 (N_7467,N_3416,N_4509);
nand U7468 (N_7468,N_4423,N_3841);
and U7469 (N_7469,N_4680,N_3236);
or U7470 (N_7470,N_2607,N_4533);
or U7471 (N_7471,N_4684,N_4334);
or U7472 (N_7472,N_4976,N_3692);
and U7473 (N_7473,N_3872,N_4742);
nand U7474 (N_7474,N_4140,N_4606);
nand U7475 (N_7475,N_3041,N_4099);
nand U7476 (N_7476,N_3042,N_4063);
nand U7477 (N_7477,N_4761,N_3559);
nand U7478 (N_7478,N_2519,N_2607);
nand U7479 (N_7479,N_4542,N_3917);
and U7480 (N_7480,N_4042,N_2879);
or U7481 (N_7481,N_3716,N_4424);
xnor U7482 (N_7482,N_3462,N_3838);
nor U7483 (N_7483,N_3464,N_4962);
or U7484 (N_7484,N_3232,N_2913);
xnor U7485 (N_7485,N_3863,N_2678);
nor U7486 (N_7486,N_4831,N_4873);
nor U7487 (N_7487,N_2591,N_4263);
xor U7488 (N_7488,N_2855,N_4309);
nor U7489 (N_7489,N_4609,N_3567);
or U7490 (N_7490,N_4085,N_4977);
nor U7491 (N_7491,N_4722,N_4449);
nor U7492 (N_7492,N_3747,N_3934);
and U7493 (N_7493,N_4310,N_2552);
nor U7494 (N_7494,N_3202,N_3678);
nand U7495 (N_7495,N_4524,N_3824);
nand U7496 (N_7496,N_3477,N_4378);
nand U7497 (N_7497,N_3455,N_4783);
nand U7498 (N_7498,N_4315,N_4844);
nand U7499 (N_7499,N_3365,N_3050);
and U7500 (N_7500,N_6781,N_5423);
or U7501 (N_7501,N_6711,N_7256);
nand U7502 (N_7502,N_5893,N_5536);
and U7503 (N_7503,N_6935,N_5636);
or U7504 (N_7504,N_5164,N_5931);
nand U7505 (N_7505,N_5960,N_7221);
and U7506 (N_7506,N_5713,N_5583);
or U7507 (N_7507,N_6103,N_6651);
nand U7508 (N_7508,N_6078,N_6617);
nor U7509 (N_7509,N_6331,N_6934);
or U7510 (N_7510,N_7405,N_5548);
nand U7511 (N_7511,N_6429,N_7022);
and U7512 (N_7512,N_5836,N_6374);
or U7513 (N_7513,N_6569,N_6663);
nand U7514 (N_7514,N_7245,N_6948);
and U7515 (N_7515,N_6991,N_7003);
or U7516 (N_7516,N_6978,N_6485);
xnor U7517 (N_7517,N_5947,N_6951);
and U7518 (N_7518,N_5890,N_6507);
or U7519 (N_7519,N_7372,N_5675);
nor U7520 (N_7520,N_5585,N_5072);
and U7521 (N_7521,N_5137,N_7373);
nor U7522 (N_7522,N_7420,N_6520);
xor U7523 (N_7523,N_6529,N_6113);
nand U7524 (N_7524,N_7271,N_6330);
and U7525 (N_7525,N_5527,N_5922);
nor U7526 (N_7526,N_5278,N_5083);
or U7527 (N_7527,N_6905,N_5531);
and U7528 (N_7528,N_6051,N_6001);
and U7529 (N_7529,N_7430,N_7314);
nand U7530 (N_7530,N_6707,N_6914);
nand U7531 (N_7531,N_5982,N_5584);
or U7532 (N_7532,N_6325,N_5436);
xnor U7533 (N_7533,N_5253,N_5441);
or U7534 (N_7534,N_6973,N_5188);
nand U7535 (N_7535,N_7422,N_5352);
nand U7536 (N_7536,N_5267,N_6696);
nor U7537 (N_7537,N_6567,N_5353);
nor U7538 (N_7538,N_6438,N_5217);
or U7539 (N_7539,N_7121,N_6558);
or U7540 (N_7540,N_7016,N_6010);
nand U7541 (N_7541,N_5777,N_6445);
and U7542 (N_7542,N_5538,N_6189);
and U7543 (N_7543,N_5582,N_7493);
or U7544 (N_7544,N_6441,N_5132);
or U7545 (N_7545,N_7228,N_7268);
or U7546 (N_7546,N_5943,N_7112);
nor U7547 (N_7547,N_6662,N_5081);
nand U7548 (N_7548,N_6106,N_5738);
nand U7549 (N_7549,N_6862,N_5948);
or U7550 (N_7550,N_7125,N_5274);
and U7551 (N_7551,N_5884,N_7429);
nand U7552 (N_7552,N_6299,N_5104);
nand U7553 (N_7553,N_5649,N_5528);
nor U7554 (N_7554,N_6022,N_6112);
nand U7555 (N_7555,N_7053,N_7357);
or U7556 (N_7556,N_5568,N_6263);
or U7557 (N_7557,N_6518,N_5085);
nor U7558 (N_7558,N_6576,N_5248);
and U7559 (N_7559,N_6913,N_7036);
nor U7560 (N_7560,N_5607,N_7288);
or U7561 (N_7561,N_5163,N_6882);
nor U7562 (N_7562,N_6767,N_7129);
nand U7563 (N_7563,N_5741,N_5261);
and U7564 (N_7564,N_6346,N_7331);
nor U7565 (N_7565,N_7078,N_5417);
xor U7566 (N_7566,N_6093,N_5219);
and U7567 (N_7567,N_5485,N_6535);
nand U7568 (N_7568,N_7048,N_5869);
nand U7569 (N_7569,N_5464,N_5133);
and U7570 (N_7570,N_6494,N_5972);
nor U7571 (N_7571,N_5341,N_5720);
nand U7572 (N_7572,N_6750,N_5399);
nand U7573 (N_7573,N_6616,N_7047);
nor U7574 (N_7574,N_6413,N_5180);
nor U7575 (N_7575,N_6497,N_5546);
nor U7576 (N_7576,N_5109,N_5829);
and U7577 (N_7577,N_5116,N_6721);
nand U7578 (N_7578,N_6650,N_5867);
nand U7579 (N_7579,N_6185,N_6876);
nand U7580 (N_7580,N_6820,N_7486);
and U7581 (N_7581,N_6077,N_6594);
or U7582 (N_7582,N_5051,N_6436);
xnor U7583 (N_7583,N_5925,N_7365);
and U7584 (N_7584,N_5186,N_7173);
or U7585 (N_7585,N_5511,N_6958);
xnor U7586 (N_7586,N_5593,N_5413);
nor U7587 (N_7587,N_7386,N_5858);
or U7588 (N_7588,N_5192,N_6336);
or U7589 (N_7589,N_5973,N_6961);
xnor U7590 (N_7590,N_5037,N_6015);
and U7591 (N_7591,N_7251,N_6194);
and U7592 (N_7592,N_5386,N_6603);
nor U7593 (N_7593,N_7382,N_5087);
nand U7594 (N_7594,N_6805,N_5375);
nor U7595 (N_7595,N_7073,N_6684);
or U7596 (N_7596,N_6005,N_6070);
nand U7597 (N_7597,N_6170,N_5339);
or U7598 (N_7598,N_6853,N_6916);
nor U7599 (N_7599,N_7227,N_6851);
and U7600 (N_7600,N_5385,N_7324);
nand U7601 (N_7601,N_5648,N_6240);
xnor U7602 (N_7602,N_5052,N_6858);
nand U7603 (N_7603,N_6364,N_6703);
or U7604 (N_7604,N_5055,N_6908);
and U7605 (N_7605,N_5557,N_6579);
xnor U7606 (N_7606,N_7274,N_7187);
xnor U7607 (N_7607,N_7403,N_6954);
and U7608 (N_7608,N_5840,N_6704);
nor U7609 (N_7609,N_6880,N_7341);
or U7610 (N_7610,N_5610,N_7337);
nor U7611 (N_7611,N_7072,N_6729);
nand U7612 (N_7612,N_5977,N_6047);
nand U7613 (N_7613,N_6584,N_6503);
nor U7614 (N_7614,N_7316,N_5018);
nor U7615 (N_7615,N_6629,N_5785);
nand U7616 (N_7616,N_7496,N_7024);
nor U7617 (N_7617,N_6502,N_5886);
and U7618 (N_7618,N_5329,N_5150);
or U7619 (N_7619,N_5257,N_6139);
xor U7620 (N_7620,N_7332,N_6116);
nand U7621 (N_7621,N_7298,N_5558);
or U7622 (N_7622,N_6418,N_6555);
and U7623 (N_7623,N_5733,N_7065);
and U7624 (N_7624,N_6164,N_7211);
or U7625 (N_7625,N_5690,N_6631);
nor U7626 (N_7626,N_5949,N_5486);
nor U7627 (N_7627,N_6832,N_6526);
xor U7628 (N_7628,N_5287,N_7296);
and U7629 (N_7629,N_7077,N_6447);
nand U7630 (N_7630,N_6976,N_6821);
nand U7631 (N_7631,N_6673,N_7344);
nand U7632 (N_7632,N_6014,N_6621);
nand U7633 (N_7633,N_5643,N_5476);
and U7634 (N_7634,N_5455,N_5667);
nand U7635 (N_7635,N_6151,N_6100);
nor U7636 (N_7636,N_7363,N_7094);
and U7637 (N_7637,N_7278,N_5942);
nand U7638 (N_7638,N_6203,N_7292);
or U7639 (N_7639,N_5612,N_6333);
or U7640 (N_7640,N_7428,N_7285);
and U7641 (N_7641,N_5303,N_6233);
nand U7642 (N_7642,N_7495,N_6216);
nand U7643 (N_7643,N_5903,N_5623);
nand U7644 (N_7644,N_5915,N_5802);
and U7645 (N_7645,N_5856,N_7389);
and U7646 (N_7646,N_5337,N_7179);
nor U7647 (N_7647,N_6857,N_7297);
xnor U7648 (N_7648,N_5497,N_5026);
nand U7649 (N_7649,N_5070,N_5280);
nand U7650 (N_7650,N_6126,N_6319);
and U7651 (N_7651,N_7335,N_5433);
and U7652 (N_7652,N_7485,N_6271);
nor U7653 (N_7653,N_5999,N_7433);
nand U7654 (N_7654,N_6306,N_5173);
nand U7655 (N_7655,N_5149,N_5182);
nor U7656 (N_7656,N_5294,N_5388);
nand U7657 (N_7657,N_7273,N_6053);
and U7658 (N_7658,N_5556,N_7074);
or U7659 (N_7659,N_6893,N_6562);
nand U7660 (N_7660,N_7404,N_7415);
nor U7661 (N_7661,N_7396,N_5064);
and U7662 (N_7662,N_5595,N_5065);
or U7663 (N_7663,N_5160,N_5233);
nor U7664 (N_7664,N_7455,N_6697);
and U7665 (N_7665,N_5514,N_5803);
and U7666 (N_7666,N_6796,N_7066);
nand U7667 (N_7667,N_6264,N_5053);
nand U7668 (N_7668,N_6700,N_5758);
and U7669 (N_7669,N_7425,N_7023);
nand U7670 (N_7670,N_6570,N_5314);
nor U7671 (N_7671,N_5806,N_6534);
and U7672 (N_7672,N_5014,N_7416);
nor U7673 (N_7673,N_5835,N_5794);
and U7674 (N_7674,N_6049,N_7131);
nor U7675 (N_7675,N_6204,N_7358);
or U7676 (N_7676,N_5826,N_6907);
and U7677 (N_7677,N_6727,N_6826);
nand U7678 (N_7678,N_6715,N_7242);
and U7679 (N_7679,N_6597,N_5761);
or U7680 (N_7680,N_5379,N_7265);
and U7681 (N_7681,N_5390,N_5533);
nand U7682 (N_7682,N_7175,N_6870);
nor U7683 (N_7683,N_6746,N_5542);
xnor U7684 (N_7684,N_7069,N_6165);
and U7685 (N_7685,N_7472,N_6394);
or U7686 (N_7686,N_6722,N_7134);
and U7687 (N_7687,N_7307,N_5962);
xnor U7688 (N_7688,N_5708,N_6708);
nor U7689 (N_7689,N_6743,N_7200);
nor U7690 (N_7690,N_6459,N_5235);
nand U7691 (N_7691,N_7317,N_5193);
and U7692 (N_7692,N_6361,N_5916);
and U7693 (N_7693,N_7064,N_6278);
and U7694 (N_7694,N_5488,N_7427);
or U7695 (N_7695,N_5504,N_6176);
nor U7696 (N_7696,N_6309,N_6351);
and U7697 (N_7697,N_5951,N_5953);
nor U7698 (N_7698,N_5816,N_5776);
nor U7699 (N_7699,N_7349,N_5577);
nor U7700 (N_7700,N_6775,N_6301);
nand U7701 (N_7701,N_6793,N_5786);
nor U7702 (N_7702,N_6774,N_5174);
nor U7703 (N_7703,N_5753,N_7398);
nor U7704 (N_7704,N_6467,N_5586);
or U7705 (N_7705,N_6384,N_6777);
nand U7706 (N_7706,N_5209,N_6886);
nor U7707 (N_7707,N_5566,N_5978);
nor U7708 (N_7708,N_6699,N_7436);
or U7709 (N_7709,N_5112,N_6895);
nand U7710 (N_7710,N_6039,N_7026);
and U7711 (N_7711,N_7119,N_5468);
or U7712 (N_7712,N_5660,N_6448);
or U7713 (N_7713,N_6052,N_6736);
nor U7714 (N_7714,N_5853,N_7007);
nand U7715 (N_7715,N_5359,N_5172);
and U7716 (N_7716,N_5707,N_6768);
nand U7717 (N_7717,N_6614,N_7124);
or U7718 (N_7718,N_5218,N_7088);
and U7719 (N_7719,N_5606,N_6063);
nand U7720 (N_7720,N_5622,N_7244);
or U7721 (N_7721,N_5282,N_6933);
or U7722 (N_7722,N_7194,N_6242);
and U7723 (N_7723,N_6510,N_5271);
xnor U7724 (N_7724,N_7402,N_6407);
nand U7725 (N_7725,N_5317,N_5935);
nand U7726 (N_7726,N_6387,N_5555);
or U7727 (N_7727,N_6249,N_6468);
nand U7728 (N_7728,N_6382,N_7340);
nor U7729 (N_7729,N_7474,N_7231);
nor U7730 (N_7730,N_5700,N_6313);
or U7731 (N_7731,N_6745,N_6486);
nor U7732 (N_7732,N_6643,N_5693);
or U7733 (N_7733,N_5318,N_5493);
nand U7734 (N_7734,N_7159,N_5797);
or U7735 (N_7735,N_6298,N_7034);
or U7736 (N_7736,N_6237,N_5967);
nand U7737 (N_7737,N_5449,N_5213);
nand U7738 (N_7738,N_5872,N_6446);
or U7739 (N_7739,N_7042,N_5347);
nand U7740 (N_7740,N_6927,N_6683);
nand U7741 (N_7741,N_5429,N_6653);
and U7742 (N_7742,N_5238,N_6002);
or U7743 (N_7743,N_5461,N_5196);
nor U7744 (N_7744,N_5703,N_6023);
and U7745 (N_7745,N_6910,N_7126);
nand U7746 (N_7746,N_6060,N_5204);
or U7747 (N_7747,N_7356,N_6389);
nand U7748 (N_7748,N_5025,N_6265);
or U7749 (N_7749,N_5078,N_5283);
or U7750 (N_7750,N_5778,N_5161);
or U7751 (N_7751,N_6232,N_6037);
or U7752 (N_7752,N_5073,N_7446);
and U7753 (N_7753,N_5006,N_7461);
nand U7754 (N_7754,N_6094,N_5565);
and U7755 (N_7755,N_6284,N_5575);
nand U7756 (N_7756,N_6142,N_6071);
and U7757 (N_7757,N_6637,N_7199);
and U7758 (N_7758,N_5602,N_5743);
nor U7759 (N_7759,N_5631,N_5831);
nand U7760 (N_7760,N_6644,N_5661);
nand U7761 (N_7761,N_6321,N_6557);
or U7762 (N_7762,N_6957,N_5941);
nand U7763 (N_7763,N_5662,N_7190);
or U7764 (N_7764,N_5044,N_6524);
nor U7765 (N_7765,N_5765,N_6725);
or U7766 (N_7766,N_6160,N_5599);
nor U7767 (N_7767,N_6551,N_5594);
nor U7768 (N_7768,N_6871,N_6897);
xnor U7769 (N_7769,N_5928,N_5001);
or U7770 (N_7770,N_5270,N_5677);
or U7771 (N_7771,N_5721,N_6169);
and U7772 (N_7772,N_6463,N_5343);
or U7773 (N_7773,N_6422,N_5820);
nor U7774 (N_7774,N_5189,N_7246);
or U7775 (N_7775,N_7452,N_6028);
nor U7776 (N_7776,N_6152,N_7106);
nand U7777 (N_7777,N_5907,N_5264);
and U7778 (N_7778,N_6251,N_6872);
and U7779 (N_7779,N_5710,N_6068);
and U7780 (N_7780,N_6695,N_5428);
or U7781 (N_7781,N_7409,N_6952);
and U7782 (N_7782,N_5443,N_5042);
and U7783 (N_7783,N_5888,N_6716);
or U7784 (N_7784,N_7417,N_7305);
nand U7785 (N_7785,N_6754,N_6399);
and U7786 (N_7786,N_6492,N_6188);
and U7787 (N_7787,N_6756,N_6223);
nor U7788 (N_7788,N_7489,N_5800);
nor U7789 (N_7789,N_7424,N_5279);
nor U7790 (N_7790,N_5405,N_7328);
and U7791 (N_7791,N_6148,N_6785);
xor U7792 (N_7792,N_6818,N_5860);
nand U7793 (N_7793,N_5492,N_5277);
and U7794 (N_7794,N_6092,N_5658);
and U7795 (N_7795,N_6274,N_7054);
and U7796 (N_7796,N_5458,N_7043);
or U7797 (N_7797,N_6838,N_6064);
nand U7798 (N_7798,N_6811,N_5451);
and U7799 (N_7799,N_5746,N_5234);
nor U7800 (N_7800,N_5847,N_7321);
nand U7801 (N_7801,N_6450,N_5121);
nor U7802 (N_7802,N_6055,N_6356);
or U7803 (N_7803,N_6589,N_5704);
nand U7804 (N_7804,N_5141,N_5273);
and U7805 (N_7805,N_6168,N_6211);
or U7806 (N_7806,N_5683,N_6987);
xor U7807 (N_7807,N_7157,N_6606);
nor U7808 (N_7808,N_6867,N_6545);
nand U7809 (N_7809,N_5203,N_6848);
or U7810 (N_7810,N_7249,N_5139);
and U7811 (N_7811,N_5790,N_5987);
nor U7812 (N_7812,N_5370,N_6806);
nor U7813 (N_7813,N_5611,N_5914);
and U7814 (N_7814,N_6656,N_5571);
and U7815 (N_7815,N_5205,N_6532);
nand U7816 (N_7816,N_6975,N_7250);
and U7817 (N_7817,N_6084,N_7395);
nor U7818 (N_7818,N_7336,N_7174);
nor U7819 (N_7819,N_5047,N_6780);
and U7820 (N_7820,N_5288,N_5002);
or U7821 (N_7821,N_5851,N_5041);
nand U7822 (N_7822,N_6638,N_5515);
nor U7823 (N_7823,N_7475,N_5102);
and U7824 (N_7824,N_5090,N_5828);
nor U7825 (N_7825,N_5082,N_5088);
nand U7826 (N_7826,N_7439,N_5854);
nor U7827 (N_7827,N_5115,N_6276);
and U7828 (N_7828,N_5739,N_7441);
nand U7829 (N_7829,N_6288,N_5010);
or U7830 (N_7830,N_5861,N_6726);
nand U7831 (N_7831,N_6326,N_6732);
and U7832 (N_7832,N_7302,N_5201);
xor U7833 (N_7833,N_6046,N_5769);
nand U7834 (N_7834,N_5034,N_6904);
and U7835 (N_7835,N_7276,N_6040);
or U7836 (N_7836,N_5430,N_5499);
nor U7837 (N_7837,N_5258,N_6409);
and U7838 (N_7838,N_6006,N_6235);
nand U7839 (N_7839,N_5153,N_6665);
or U7840 (N_7840,N_5197,N_6802);
nand U7841 (N_7841,N_5123,N_7193);
nand U7842 (N_7842,N_5130,N_5729);
nor U7843 (N_7843,N_5437,N_6936);
nor U7844 (N_7844,N_7361,N_5605);
nand U7845 (N_7845,N_5742,N_6931);
and U7846 (N_7846,N_6191,N_7044);
and U7847 (N_7847,N_5609,N_6672);
and U7848 (N_7848,N_7029,N_6482);
and U7849 (N_7849,N_5899,N_5954);
or U7850 (N_7850,N_5841,N_7240);
nor U7851 (N_7851,N_5313,N_5269);
nor U7852 (N_7852,N_6842,N_6034);
nor U7853 (N_7853,N_6342,N_7095);
nor U7854 (N_7854,N_6115,N_7368);
nand U7855 (N_7855,N_6813,N_6398);
nor U7856 (N_7856,N_6733,N_7442);
nand U7857 (N_7857,N_7058,N_6368);
or U7858 (N_7858,N_6369,N_7261);
nand U7859 (N_7859,N_5466,N_6314);
or U7860 (N_7860,N_5712,N_6628);
or U7861 (N_7861,N_6065,N_7153);
or U7862 (N_7862,N_5927,N_6088);
and U7863 (N_7863,N_6324,N_7380);
nor U7864 (N_7864,N_7113,N_5208);
or U7865 (N_7865,N_5517,N_5618);
nor U7866 (N_7866,N_5652,N_5415);
or U7867 (N_7867,N_5224,N_6588);
nand U7868 (N_7868,N_6879,N_6619);
nor U7869 (N_7869,N_5509,N_7394);
nor U7870 (N_7870,N_7338,N_6636);
nand U7871 (N_7871,N_6270,N_6391);
and U7872 (N_7872,N_6779,N_6512);
nand U7873 (N_7873,N_6041,N_5796);
or U7874 (N_7874,N_5645,N_5381);
nand U7875 (N_7875,N_7306,N_6220);
or U7876 (N_7876,N_6903,N_7289);
nor U7877 (N_7877,N_5033,N_5118);
nor U7878 (N_7878,N_6412,N_7186);
or U7879 (N_7879,N_6568,N_5988);
nor U7880 (N_7880,N_6846,N_5679);
and U7881 (N_7881,N_5852,N_5236);
nor U7882 (N_7882,N_5748,N_5136);
or U7883 (N_7883,N_5633,N_5603);
nand U7884 (N_7884,N_5911,N_5022);
nor U7885 (N_7885,N_7046,N_5276);
nand U7886 (N_7886,N_7201,N_5537);
or U7887 (N_7887,N_6114,N_6547);
or U7888 (N_7888,N_5470,N_6222);
nand U7889 (N_7889,N_5545,N_7255);
or U7890 (N_7890,N_5501,N_5245);
and U7891 (N_7891,N_5570,N_7217);
and U7892 (N_7892,N_5870,N_7258);
xor U7893 (N_7893,N_5810,N_6787);
and U7894 (N_7894,N_6839,N_6538);
and U7895 (N_7895,N_6424,N_5342);
and U7896 (N_7896,N_7342,N_5754);
nand U7897 (N_7897,N_6283,N_5457);
or U7898 (N_7898,N_6860,N_6076);
nand U7899 (N_7899,N_5069,N_6472);
and U7900 (N_7900,N_7421,N_6375);
or U7901 (N_7901,N_6601,N_7115);
nand U7902 (N_7902,N_5335,N_7165);
xnor U7903 (N_7903,N_6670,N_5165);
nand U7904 (N_7904,N_5963,N_7435);
or U7905 (N_7905,N_5183,N_6523);
or U7906 (N_7906,N_5589,N_7020);
nor U7907 (N_7907,N_5480,N_6640);
nand U7908 (N_7908,N_5009,N_5292);
xnor U7909 (N_7909,N_5334,N_6344);
nand U7910 (N_7910,N_5706,N_7359);
xnor U7911 (N_7911,N_5992,N_5642);
nor U7912 (N_7912,N_6290,N_6335);
nand U7913 (N_7913,N_6930,N_6849);
nand U7914 (N_7914,N_7414,N_6671);
and U7915 (N_7915,N_5863,N_5502);
nor U7916 (N_7916,N_7346,N_6997);
nor U7917 (N_7917,N_5285,N_5672);
nand U7918 (N_7918,N_5075,N_5946);
nand U7919 (N_7919,N_6845,N_6003);
or U7920 (N_7920,N_5289,N_7408);
and U7921 (N_7921,N_6807,N_6117);
or U7922 (N_7922,N_7032,N_5979);
nor U7923 (N_7923,N_5663,N_6552);
nand U7924 (N_7924,N_6789,N_5145);
or U7925 (N_7925,N_5788,N_5625);
or U7926 (N_7926,N_7039,N_5553);
and U7927 (N_7927,N_7313,N_5795);
and U7928 (N_7928,N_6676,N_5510);
nand U7929 (N_7929,N_6835,N_7028);
and U7930 (N_7930,N_6723,N_7438);
nand U7931 (N_7931,N_5926,N_6172);
or U7932 (N_7932,N_5834,N_6912);
or U7933 (N_7933,N_7293,N_6373);
nand U7934 (N_7934,N_6564,N_5837);
or U7935 (N_7935,N_5873,N_6207);
and U7936 (N_7936,N_5275,N_6949);
or U7937 (N_7937,N_5237,N_6067);
nand U7938 (N_7938,N_5808,N_5923);
and U7939 (N_7939,N_6371,N_6423);
and U7940 (N_7940,N_6761,N_6253);
or U7941 (N_7941,N_5671,N_6928);
and U7942 (N_7942,N_5030,N_6004);
or U7943 (N_7943,N_6759,N_7009);
or U7944 (N_7944,N_5822,N_5627);
nor U7945 (N_7945,N_6804,N_6501);
nor U7946 (N_7946,N_5930,N_5398);
or U7947 (N_7947,N_6219,N_5411);
nor U7948 (N_7948,N_5507,N_6110);
and U7949 (N_7949,N_7146,N_6577);
nor U7950 (N_7950,N_6701,N_7225);
or U7951 (N_7951,N_6019,N_5590);
nand U7952 (N_7952,N_6527,N_6362);
or U7953 (N_7953,N_6944,N_7456);
nand U7954 (N_7954,N_5737,N_6747);
or U7955 (N_7955,N_7238,N_5408);
or U7956 (N_7956,N_5881,N_5908);
or U7957 (N_7957,N_7312,N_5143);
and U7958 (N_7958,N_6825,N_5877);
or U7959 (N_7959,N_5906,N_6575);
xnor U7960 (N_7960,N_7303,N_6924);
nand U7961 (N_7961,N_6593,N_5670);
or U7962 (N_7962,N_6377,N_5995);
nand U7963 (N_7963,N_7379,N_5198);
nand U7964 (N_7964,N_7236,N_6144);
or U7965 (N_7965,N_6660,N_5815);
nand U7966 (N_7966,N_6082,N_5079);
or U7967 (N_7967,N_5843,N_6347);
or U7968 (N_7968,N_7458,N_5020);
and U7969 (N_7969,N_7291,N_7052);
and U7970 (N_7970,N_5581,N_5924);
nand U7971 (N_7971,N_5715,N_5695);
nand U7972 (N_7972,N_5940,N_6668);
nor U7973 (N_7973,N_7170,N_5354);
nand U7974 (N_7974,N_6909,N_6795);
or U7975 (N_7975,N_7377,N_6231);
nand U7976 (N_7976,N_6059,N_7197);
or U7977 (N_7977,N_5503,N_7070);
nor U7978 (N_7978,N_6247,N_6718);
nand U7979 (N_7979,N_5396,N_5789);
or U7980 (N_7980,N_5215,N_6018);
and U7981 (N_7981,N_5159,N_6964);
nand U7982 (N_7982,N_7041,N_6517);
nand U7983 (N_7983,N_5475,N_6658);
and U7984 (N_7984,N_5444,N_7209);
nor U7985 (N_7985,N_6618,N_5422);
nor U7986 (N_7986,N_7309,N_7378);
or U7987 (N_7987,N_6980,N_5360);
and U7988 (N_7988,N_5157,N_6828);
nand U7989 (N_7989,N_5832,N_6647);
and U7990 (N_7990,N_6180,N_5284);
nor U7991 (N_7991,N_5015,N_7375);
xor U7992 (N_7992,N_5574,N_5063);
nand U7993 (N_7993,N_7447,N_5176);
and U7994 (N_7994,N_7055,N_5067);
xnor U7995 (N_7995,N_6427,N_6841);
nor U7996 (N_7996,N_5784,N_5855);
xor U7997 (N_7997,N_7253,N_5358);
nand U7998 (N_7998,N_5956,N_7451);
nor U7999 (N_7999,N_6762,N_6045);
or U8000 (N_8000,N_5591,N_7391);
nor U8001 (N_8001,N_5554,N_7329);
nand U8002 (N_8002,N_6221,N_7367);
nand U8003 (N_8003,N_6434,N_5698);
nand U8004 (N_8004,N_7037,N_5680);
xor U8005 (N_8005,N_6228,N_7166);
or U8006 (N_8006,N_6030,N_5036);
nor U8007 (N_8007,N_6955,N_5697);
and U8008 (N_8008,N_6519,N_7318);
nor U8009 (N_8009,N_5750,N_5120);
and U8010 (N_8010,N_5702,N_6452);
or U8011 (N_8011,N_5369,N_5098);
or U8012 (N_8012,N_6227,N_6224);
nor U8013 (N_8013,N_6989,N_7116);
xor U8014 (N_8014,N_6887,N_7364);
xor U8015 (N_8015,N_6977,N_5857);
or U8016 (N_8016,N_6465,N_6343);
or U8017 (N_8017,N_6317,N_6884);
xor U8018 (N_8018,N_5541,N_6932);
nand U8019 (N_8019,N_6072,N_5617);
nand U8020 (N_8020,N_5896,N_5228);
nor U8021 (N_8021,N_5027,N_7400);
nand U8022 (N_8022,N_6633,N_7011);
nor U8023 (N_8023,N_6121,N_6033);
or U8024 (N_8024,N_6359,N_6021);
nand U8025 (N_8025,N_6738,N_6354);
and U8026 (N_8026,N_7185,N_6856);
or U8027 (N_8027,N_5561,N_7347);
or U8028 (N_8028,N_7334,N_6246);
or U8029 (N_8029,N_5225,N_5902);
and U8030 (N_8030,N_6200,N_7013);
and U8031 (N_8031,N_5489,N_7206);
xor U8032 (N_8032,N_5821,N_6544);
and U8033 (N_8033,N_6020,N_6815);
and U8034 (N_8034,N_6130,N_5391);
or U8035 (N_8035,N_5268,N_7345);
and U8036 (N_8036,N_5547,N_7093);
or U8037 (N_8037,N_6560,N_7330);
nand U8038 (N_8038,N_6769,N_5409);
nor U8039 (N_8039,N_5040,N_5779);
nor U8040 (N_8040,N_7243,N_6784);
and U8041 (N_8041,N_5990,N_5673);
and U8042 (N_8042,N_6590,N_7056);
nand U8043 (N_8043,N_6748,N_6918);
or U8044 (N_8044,N_7478,N_5387);
nand U8045 (N_8045,N_6902,N_6259);
nor U8046 (N_8046,N_5952,N_5412);
nand U8047 (N_8047,N_7381,N_5074);
or U8048 (N_8048,N_6016,N_6837);
and U8049 (N_8049,N_6066,N_7263);
nor U8050 (N_8050,N_5106,N_7141);
and U8051 (N_8051,N_5263,N_6624);
nand U8052 (N_8052,N_6256,N_6735);
or U8053 (N_8053,N_5024,N_6044);
and U8054 (N_8054,N_6613,N_5879);
nor U8055 (N_8055,N_5937,N_5050);
and U8056 (N_8056,N_6488,N_5366);
nor U8057 (N_8057,N_5687,N_5424);
or U8058 (N_8058,N_6822,N_5874);
nand U8059 (N_8059,N_6153,N_7287);
and U8060 (N_8060,N_5876,N_6268);
nand U8061 (N_8061,N_7497,N_5402);
nor U8062 (N_8062,N_7230,N_7254);
or U8063 (N_8063,N_6899,N_6303);
nor U8064 (N_8064,N_5534,N_5897);
nand U8065 (N_8065,N_6599,N_7448);
nor U8066 (N_8066,N_6109,N_5901);
or U8067 (N_8067,N_7492,N_5168);
or U8068 (N_8068,N_6766,N_5580);
nand U8069 (N_8069,N_7311,N_5699);
nand U8070 (N_8070,N_7155,N_6571);
and U8071 (N_8071,N_5077,N_7387);
nand U8072 (N_8072,N_7150,N_6854);
xnor U8073 (N_8073,N_7136,N_6102);
or U8074 (N_8074,N_6505,N_5587);
or U8075 (N_8075,N_5383,N_5440);
and U8076 (N_8076,N_5560,N_6740);
and U8077 (N_8077,N_7140,N_5483);
nor U8078 (N_8078,N_6241,N_6600);
and U8079 (N_8079,N_6426,N_6753);
nor U8080 (N_8080,N_6120,N_7130);
xor U8081 (N_8081,N_5850,N_6824);
nor U8082 (N_8082,N_5921,N_5066);
and U8083 (N_8083,N_7101,N_5151);
and U8084 (N_8084,N_6458,N_5046);
or U8085 (N_8085,N_5985,N_7120);
nand U8086 (N_8086,N_6892,N_6686);
nand U8087 (N_8087,N_6181,N_6710);
nand U8088 (N_8088,N_6864,N_5421);
nand U8089 (N_8089,N_6607,N_7067);
nor U8090 (N_8090,N_6277,N_7484);
or U8091 (N_8091,N_7160,N_5374);
or U8092 (N_8092,N_7222,N_6511);
nor U8093 (N_8093,N_5416,N_5350);
nor U8094 (N_8094,N_6993,N_6294);
nand U8095 (N_8095,N_5838,N_5752);
nor U8096 (N_8096,N_5304,N_5525);
nand U8097 (N_8097,N_5105,N_5844);
nand U8098 (N_8098,N_7117,N_5969);
nor U8099 (N_8099,N_5091,N_5434);
nand U8100 (N_8100,N_5054,N_5717);
or U8101 (N_8101,N_7223,N_5559);
and U8102 (N_8102,N_7152,N_6122);
or U8103 (N_8103,N_7213,N_6236);
or U8104 (N_8104,N_6580,N_5508);
or U8105 (N_8105,N_5848,N_6027);
nand U8106 (N_8106,N_6554,N_5068);
nor U8107 (N_8107,N_5035,N_6585);
nand U8108 (N_8108,N_7308,N_6129);
and U8109 (N_8109,N_7370,N_6500);
nand U8110 (N_8110,N_6042,N_6455);
nor U8111 (N_8111,N_5327,N_6755);
and U8112 (N_8112,N_6210,N_6057);
or U8113 (N_8113,N_5813,N_6490);
nor U8114 (N_8114,N_7315,N_6548);
or U8115 (N_8115,N_7488,N_6891);
nand U8116 (N_8116,N_7085,N_5320);
and U8117 (N_8117,N_7195,N_6182);
nor U8118 (N_8118,N_7283,N_7105);
nand U8119 (N_8119,N_7004,N_6792);
nor U8120 (N_8120,N_6058,N_5539);
nor U8121 (N_8121,N_5306,N_5725);
nor U8122 (N_8122,N_6128,N_7108);
nand U8123 (N_8123,N_6026,N_5563);
nand U8124 (N_8124,N_6782,N_5669);
or U8125 (N_8125,N_7167,N_7279);
nor U8126 (N_8126,N_6681,N_7235);
nor U8127 (N_8127,N_6469,N_6454);
nor U8128 (N_8128,N_6996,N_6208);
or U8129 (N_8129,N_7272,N_6192);
nor U8130 (N_8130,N_5825,N_6230);
or U8131 (N_8131,N_7169,N_5056);
nor U8132 (N_8132,N_7010,N_5771);
nand U8133 (N_8133,N_6473,N_5138);
or U8134 (N_8134,N_6788,N_5099);
or U8135 (N_8135,N_6542,N_5128);
nor U8136 (N_8136,N_5716,N_5281);
and U8137 (N_8137,N_5195,N_6392);
or U8138 (N_8138,N_6719,N_5601);
and U8139 (N_8139,N_5604,N_5997);
and U8140 (N_8140,N_5471,N_5249);
nand U8141 (N_8141,N_6062,N_6541);
or U8142 (N_8142,N_6741,N_5728);
and U8143 (N_8143,N_5005,N_5216);
and U8144 (N_8144,N_5103,N_5058);
nand U8145 (N_8145,N_7183,N_5092);
and U8146 (N_8146,N_7203,N_6285);
and U8147 (N_8147,N_5919,N_6400);
and U8148 (N_8148,N_7470,N_6690);
and U8149 (N_8149,N_5062,N_7295);
and U8150 (N_8150,N_5071,N_7202);
nand U8151 (N_8151,N_7025,N_6456);
nand U8152 (N_8152,N_5096,N_7142);
nor U8153 (N_8153,N_6937,N_5016);
nand U8154 (N_8154,N_6183,N_7100);
nor U8155 (N_8155,N_7476,N_5659);
xor U8156 (N_8156,N_6383,N_7033);
and U8157 (N_8157,N_5640,N_7431);
and U8158 (N_8158,N_5406,N_6669);
or U8159 (N_8159,N_6451,N_6850);
or U8160 (N_8160,N_6682,N_5763);
nor U8161 (N_8161,N_6565,N_5759);
and U8162 (N_8162,N_6460,N_6147);
nor U8163 (N_8163,N_5781,N_5597);
and U8164 (N_8164,N_6430,N_6213);
or U8165 (N_8165,N_5125,N_5191);
and U8166 (N_8166,N_5722,N_6595);
and U8167 (N_8167,N_6917,N_5004);
nor U8168 (N_8168,N_7339,N_6202);
or U8169 (N_8169,N_7463,N_6950);
or U8170 (N_8170,N_7366,N_7216);
nand U8171 (N_8171,N_6218,N_6525);
or U8172 (N_8172,N_6372,N_5447);
nand U8173 (N_8173,N_6974,N_5827);
or U8174 (N_8174,N_5167,N_6272);
nand U8175 (N_8175,N_7212,N_6808);
nand U8176 (N_8176,N_6437,N_7107);
and U8177 (N_8177,N_6877,N_7079);
or U8178 (N_8178,N_7499,N_5108);
and U8179 (N_8179,N_7284,N_5262);
nand U8180 (N_8180,N_7397,N_6763);
and U8181 (N_8181,N_5770,N_5964);
and U8182 (N_8182,N_5222,N_5348);
nor U8183 (N_8183,N_5839,N_5849);
nand U8184 (N_8184,N_6641,N_6573);
and U8185 (N_8185,N_6646,N_6664);
nand U8186 (N_8186,N_5003,N_7333);
nand U8187 (N_8187,N_7133,N_7494);
nor U8188 (N_8188,N_5450,N_6966);
or U8189 (N_8189,N_5747,N_5368);
nand U8190 (N_8190,N_5818,N_6135);
or U8191 (N_8191,N_5472,N_6098);
nand U8192 (N_8192,N_5199,N_5309);
nand U8193 (N_8193,N_5126,N_6744);
nor U8194 (N_8194,N_7423,N_5635);
or U8195 (N_8195,N_5255,N_7266);
and U8196 (N_8196,N_6289,N_6124);
nor U8197 (N_8197,N_5400,N_6801);
nand U8198 (N_8198,N_5202,N_5340);
nand U8199 (N_8199,N_6890,N_5305);
and U8200 (N_8200,N_7269,N_5637);
nand U8201 (N_8201,N_7127,N_5315);
nor U8202 (N_8202,N_6765,N_6156);
nor U8203 (N_8203,N_6731,N_5319);
nor U8204 (N_8204,N_7362,N_5393);
nor U8205 (N_8205,N_6985,N_7144);
nor U8206 (N_8206,N_6118,N_7371);
xnor U8207 (N_8207,N_7111,N_5266);
or U8208 (N_8208,N_6480,N_6328);
and U8209 (N_8209,N_7189,N_6474);
nor U8210 (N_8210,N_5719,N_5324);
nand U8211 (N_8211,N_5535,N_7450);
nor U8212 (N_8212,N_7454,N_7017);
or U8213 (N_8213,N_6275,N_6691);
nor U8214 (N_8214,N_5694,N_6435);
nor U8215 (N_8215,N_6069,N_7498);
nor U8216 (N_8216,N_6481,N_6096);
and U8217 (N_8217,N_5600,N_6171);
and U8218 (N_8218,N_5970,N_6591);
nand U8219 (N_8219,N_5377,N_6645);
or U8220 (N_8220,N_5975,N_6419);
or U8221 (N_8221,N_7280,N_5043);
nand U8222 (N_8222,N_7090,N_6868);
and U8223 (N_8223,N_5380,N_7360);
or U8224 (N_8224,N_5709,N_5917);
or U8225 (N_8225,N_6988,N_6803);
nor U8226 (N_8226,N_6678,N_7449);
or U8227 (N_8227,N_5404,N_6406);
and U8228 (N_8228,N_6730,N_5127);
nor U8229 (N_8229,N_6863,N_6883);
nand U8230 (N_8230,N_5653,N_5119);
nor U8231 (N_8231,N_5107,N_6679);
nor U8232 (N_8232,N_7286,N_6137);
nor U8233 (N_8233,N_7132,N_6657);
and U8234 (N_8234,N_5361,N_6967);
nand U8235 (N_8235,N_5812,N_7172);
nor U8236 (N_8236,N_5792,N_6615);
nand U8237 (N_8237,N_6357,N_5060);
and U8238 (N_8238,N_5316,N_7156);
or U8239 (N_8239,N_7021,N_5310);
and U8240 (N_8240,N_7353,N_6471);
nor U8241 (N_8241,N_6659,N_5664);
nor U8242 (N_8242,N_5376,N_6245);
or U8243 (N_8243,N_7412,N_5651);
nand U8244 (N_8244,N_7040,N_6091);
and U8245 (N_8245,N_5243,N_5291);
nor U8246 (N_8246,N_5993,N_5665);
nor U8247 (N_8247,N_5093,N_6428);
xnor U8248 (N_8248,N_6866,N_6556);
nand U8249 (N_8249,N_7392,N_6184);
and U8250 (N_8250,N_5868,N_6693);
nor U8251 (N_8251,N_5338,N_5454);
or U8252 (N_8252,N_7218,N_5783);
and U8253 (N_8253,N_6339,N_5668);
or U8254 (N_8254,N_5101,N_6385);
or U8255 (N_8255,N_7076,N_6844);
nand U8256 (N_8256,N_7204,N_5619);
nor U8257 (N_8257,N_5212,N_7399);
and U8258 (N_8258,N_6894,N_5564);
xor U8259 (N_8259,N_5629,N_7143);
xor U8260 (N_8260,N_5804,N_5626);
nand U8261 (N_8261,N_6734,N_6865);
nor U8262 (N_8262,N_6773,N_6386);
and U8263 (N_8263,N_5705,N_5023);
nor U8264 (N_8264,N_5805,N_6986);
nand U8265 (N_8265,N_6861,N_5456);
or U8266 (N_8266,N_5971,N_7210);
xor U8267 (N_8267,N_6111,N_5206);
or U8268 (N_8268,N_7014,N_6244);
nor U8269 (N_8269,N_5181,N_7158);
nand U8270 (N_8270,N_5551,N_5000);
and U8271 (N_8271,N_7406,N_7182);
nor U8272 (N_8272,N_7445,N_5462);
or U8273 (N_8273,N_6366,N_5365);
or U8274 (N_8274,N_5147,N_5297);
nor U8275 (N_8275,N_6179,N_5723);
nand U8276 (N_8276,N_5596,N_6900);
nand U8277 (N_8277,N_6982,N_5944);
nor U8278 (N_8278,N_5148,N_5029);
or U8279 (N_8279,N_5344,N_6712);
nand U8280 (N_8280,N_5809,N_7473);
xnor U8281 (N_8281,N_6827,N_5482);
and U8282 (N_8282,N_5166,N_5220);
and U8283 (N_8283,N_5487,N_5491);
nor U8284 (N_8284,N_5934,N_5567);
or U8285 (N_8285,N_7479,N_6167);
nor U8286 (N_8286,N_6315,N_6770);
nor U8287 (N_8287,N_6087,N_7299);
or U8288 (N_8288,N_5308,N_7031);
xnor U8289 (N_8289,N_5474,N_5012);
nor U8290 (N_8290,N_6915,N_5124);
and U8291 (N_8291,N_7000,N_6345);
and U8292 (N_8292,N_5184,N_7012);
nor U8293 (N_8293,N_5371,N_6654);
and U8294 (N_8294,N_6190,N_6390);
and U8295 (N_8295,N_5986,N_5656);
and U8296 (N_8296,N_5549,N_5755);
nor U8297 (N_8297,N_6296,N_6496);
and U8298 (N_8298,N_6360,N_5395);
nand U8299 (N_8299,N_5048,N_5576);
or U8300 (N_8300,N_6206,N_5500);
or U8301 (N_8301,N_5431,N_5293);
or U8302 (N_8302,N_5918,N_6859);
or U8303 (N_8303,N_6292,N_6367);
or U8304 (N_8304,N_5239,N_6363);
nand U8305 (N_8305,N_5936,N_5397);
or U8306 (N_8306,N_7301,N_5364);
and U8307 (N_8307,N_5562,N_6476);
nor U8308 (N_8308,N_5957,N_6720);
nor U8309 (N_8309,N_6261,N_5976);
and U8310 (N_8310,N_6622,N_5345);
or U8311 (N_8311,N_5039,N_7139);
nand U8312 (N_8312,N_6572,N_5823);
nand U8313 (N_8313,N_6310,N_6239);
nand U8314 (N_8314,N_7383,N_6349);
and U8315 (N_8315,N_6634,N_5286);
nand U8316 (N_8316,N_7219,N_6509);
and U8317 (N_8317,N_5866,N_5933);
or U8318 (N_8318,N_7413,N_7063);
nor U8319 (N_8319,N_5432,N_6608);
and U8320 (N_8320,N_7393,N_5242);
or U8321 (N_8321,N_6348,N_5736);
xnor U8322 (N_8322,N_6178,N_5331);
and U8323 (N_8323,N_5959,N_6376);
and U8324 (N_8324,N_7468,N_6834);
nand U8325 (N_8325,N_6706,N_7320);
or U8326 (N_8326,N_6959,N_5259);
and U8327 (N_8327,N_7466,N_6702);
nand U8328 (N_8328,N_5152,N_5814);
and U8329 (N_8329,N_7128,N_6404);
nand U8330 (N_8330,N_5241,N_6140);
nor U8331 (N_8331,N_5330,N_5628);
nor U8332 (N_8332,N_6054,N_5889);
and U8333 (N_8333,N_5732,N_5057);
and U8334 (N_8334,N_5760,N_7161);
and U8335 (N_8335,N_6453,N_5410);
or U8336 (N_8336,N_6995,N_5974);
nor U8337 (N_8337,N_6604,N_6107);
nor U8338 (N_8338,N_6799,N_7050);
or U8339 (N_8339,N_5453,N_5211);
nor U8340 (N_8340,N_6941,N_5989);
nand U8341 (N_8341,N_5830,N_5529);
and U8342 (N_8342,N_5333,N_5938);
or U8343 (N_8343,N_5882,N_6388);
nor U8344 (N_8344,N_5214,N_5674);
xnor U8345 (N_8345,N_7233,N_6186);
nor U8346 (N_8346,N_5438,N_5641);
nand U8347 (N_8347,N_5490,N_7482);
nor U8348 (N_8348,N_7401,N_6025);
nand U8349 (N_8349,N_5146,N_6174);
nor U8350 (N_8350,N_5639,N_5256);
nor U8351 (N_8351,N_5654,N_7322);
nand U8352 (N_8352,N_6393,N_6709);
nor U8353 (N_8353,N_6953,N_7385);
and U8354 (N_8354,N_7005,N_5394);
and U8355 (N_8355,N_6442,N_5414);
or U8356 (N_8356,N_5389,N_6352);
or U8357 (N_8357,N_5177,N_6625);
and U8358 (N_8358,N_5170,N_5407);
and U8359 (N_8359,N_5021,N_6605);
and U8360 (N_8360,N_5425,N_6035);
nand U8361 (N_8361,N_5251,N_6104);
or U8362 (N_8362,N_5095,N_6757);
nand U8363 (N_8363,N_6829,N_5505);
or U8364 (N_8364,N_5221,N_7062);
nor U8365 (N_8365,N_6992,N_7135);
nor U8366 (N_8366,N_6305,N_7092);
and U8367 (N_8367,N_6611,N_5312);
and U8368 (N_8368,N_6878,N_5230);
and U8369 (N_8369,N_7138,N_6483);
nand U8370 (N_8370,N_5129,N_7188);
or U8371 (N_8371,N_5540,N_7091);
nor U8372 (N_8372,N_7462,N_7464);
nand U8373 (N_8373,N_6358,N_5349);
nand U8374 (N_8374,N_5356,N_6163);
and U8375 (N_8375,N_5135,N_5961);
and U8376 (N_8376,N_6714,N_7081);
and U8377 (N_8377,N_6417,N_6635);
nor U8378 (N_8378,N_6798,N_5382);
and U8379 (N_8379,N_7049,N_7234);
or U8380 (N_8380,N_7351,N_7418);
or U8381 (N_8381,N_7205,N_6300);
xor U8382 (N_8382,N_5965,N_5378);
and U8383 (N_8383,N_5302,N_7098);
nor U8384 (N_8384,N_6282,N_5007);
xor U8385 (N_8385,N_6008,N_6999);
nor U8386 (N_8386,N_7467,N_5764);
and U8387 (N_8387,N_5929,N_6692);
or U8388 (N_8388,N_7149,N_6685);
nor U8389 (N_8389,N_5401,N_6561);
and U8390 (N_8390,N_6431,N_6158);
or U8391 (N_8391,N_5782,N_7087);
and U8392 (N_8392,N_7083,N_5448);
or U8393 (N_8393,N_6281,N_7481);
nand U8394 (N_8394,N_6537,N_6758);
or U8395 (N_8395,N_6405,N_7057);
nor U8396 (N_8396,N_5955,N_5169);
and U8397 (N_8397,N_7260,N_6790);
nand U8398 (N_8398,N_7300,N_6786);
nor U8399 (N_8399,N_5724,N_5445);
and U8400 (N_8400,N_5880,N_6433);
or U8401 (N_8401,N_7198,N_6772);
and U8402 (N_8402,N_5701,N_6508);
nor U8403 (N_8403,N_5403,N_5384);
or U8404 (N_8404,N_6083,N_5496);
or U8405 (N_8405,N_6279,N_7281);
nor U8406 (N_8406,N_5573,N_6150);
and U8407 (N_8407,N_7035,N_5484);
nor U8408 (N_8408,N_6403,N_5311);
and U8409 (N_8409,N_7262,N_6800);
nand U8410 (N_8410,N_6771,N_5871);
nand U8411 (N_8411,N_6248,N_5467);
or U8412 (N_8412,N_5530,N_6133);
nor U8413 (N_8413,N_6814,N_6267);
nand U8414 (N_8414,N_5252,N_5891);
nor U8415 (N_8415,N_7232,N_5446);
nor U8416 (N_8416,N_6108,N_5086);
nor U8417 (N_8417,N_5113,N_6085);
nor U8418 (N_8418,N_5846,N_6370);
nor U8419 (N_8419,N_5247,N_5774);
nand U8420 (N_8420,N_5920,N_6612);
or U8421 (N_8421,N_6925,N_7038);
and U8422 (N_8422,N_5740,N_6979);
nand U8423 (N_8423,N_5756,N_5076);
and U8424 (N_8424,N_7018,N_7180);
nand U8425 (N_8425,N_6688,N_6778);
or U8426 (N_8426,N_6029,N_5520);
xor U8427 (N_8427,N_6449,N_6079);
nor U8428 (N_8428,N_7259,N_5892);
nor U8429 (N_8429,N_5495,N_6559);
or U8430 (N_8430,N_5059,N_6764);
or U8431 (N_8431,N_7410,N_5061);
nand U8432 (N_8432,N_5226,N_6632);
nor U8433 (N_8433,N_5684,N_5775);
or U8434 (N_8434,N_5142,N_5592);
and U8435 (N_8435,N_6843,N_5644);
nand U8436 (N_8436,N_6255,N_6969);
nor U8437 (N_8437,N_6320,N_5817);
or U8438 (N_8438,N_5171,N_5735);
and U8439 (N_8439,N_7348,N_5745);
or U8440 (N_8440,N_6293,N_5154);
and U8441 (N_8441,N_5655,N_6630);
and U8442 (N_8442,N_6627,N_5357);
nand U8443 (N_8443,N_7027,N_6238);
or U8444 (N_8444,N_6498,N_7352);
or U8445 (N_8445,N_5097,N_5932);
nor U8446 (N_8446,N_7118,N_7453);
nor U8447 (N_8447,N_7109,N_5013);
and U8448 (N_8448,N_7168,N_6705);
and U8449 (N_8449,N_6408,N_7068);
or U8450 (N_8450,N_6395,N_6295);
or U8451 (N_8451,N_6549,N_7325);
or U8452 (N_8452,N_6048,N_6197);
nor U8453 (N_8453,N_7355,N_6831);
nand U8454 (N_8454,N_5569,N_5824);
nand U8455 (N_8455,N_5865,N_5094);
nand U8456 (N_8456,N_7440,N_6751);
or U8457 (N_8457,N_7237,N_7407);
or U8458 (N_8458,N_6540,N_5634);
nand U8459 (N_8459,N_7252,N_6487);
nor U8460 (N_8460,N_5473,N_6254);
or U8461 (N_8461,N_7323,N_5532);
nand U8462 (N_8462,N_7327,N_5994);
nand U8463 (N_8463,N_5045,N_5945);
or U8464 (N_8464,N_5833,N_6262);
nor U8465 (N_8465,N_7163,N_6243);
nand U8466 (N_8466,N_7019,N_7241);
nand U8467 (N_8467,N_6302,N_6043);
nand U8468 (N_8468,N_7114,N_6582);
and U8469 (N_8469,N_7229,N_6136);
and U8470 (N_8470,N_5260,N_6410);
xnor U8471 (N_8471,N_7104,N_7215);
or U8472 (N_8472,N_6794,N_7419);
and U8473 (N_8473,N_5650,N_7491);
and U8474 (N_8474,N_6984,N_6141);
or U8475 (N_8475,N_5028,N_5494);
or U8476 (N_8476,N_7103,N_6687);
nand U8477 (N_8477,N_5966,N_5223);
nand U8478 (N_8478,N_7294,N_6099);
or U8479 (N_8479,N_6215,N_7207);
or U8480 (N_8480,N_6353,N_6970);
or U8481 (N_8481,N_5598,N_6214);
nand U8482 (N_8482,N_6286,N_6489);
nor U8483 (N_8483,N_6642,N_5883);
nor U8484 (N_8484,N_6173,N_6873);
nand U8485 (N_8485,N_5793,N_7145);
or U8486 (N_8486,N_7154,N_7178);
nor U8487 (N_8487,N_6816,N_5621);
nand U8488 (N_8488,N_5608,N_7171);
and U8489 (N_8489,N_6226,N_5322);
xor U8490 (N_8490,N_5647,N_6378);
and U8491 (N_8491,N_7267,N_6416);
nor U8492 (N_8492,N_6817,N_6516);
and U8493 (N_8493,N_6131,N_5200);
nor U8494 (N_8494,N_7465,N_6050);
and U8495 (N_8495,N_5272,N_7214);
nand U8496 (N_8496,N_6209,N_6443);
and U8497 (N_8497,N_5910,N_5900);
nand U8498 (N_8498,N_7443,N_5615);
or U8499 (N_8499,N_6543,N_5730);
nand U8500 (N_8500,N_5950,N_6484);
nand U8501 (N_8501,N_6420,N_6513);
nand U8502 (N_8502,N_5646,N_5996);
xor U8503 (N_8503,N_6947,N_5162);
nand U8504 (N_8504,N_6439,N_6260);
or U8505 (N_8505,N_5254,N_5210);
nand U8506 (N_8506,N_5114,N_6875);
nand U8507 (N_8507,N_6493,N_5666);
nor U8508 (N_8508,N_5772,N_6031);
and U8509 (N_8509,N_6157,N_5419);
or U8510 (N_8510,N_7147,N_7411);
nor U8511 (N_8511,N_7226,N_6648);
nand U8512 (N_8512,N_6724,N_6365);
nand U8513 (N_8513,N_6906,N_6024);
nor U8514 (N_8514,N_6332,N_6316);
and U8515 (N_8515,N_7151,N_5158);
or U8516 (N_8516,N_6649,N_6012);
nand U8517 (N_8517,N_6514,N_6578);
and U8518 (N_8518,N_6962,N_6921);
or U8519 (N_8519,N_6531,N_6089);
xor U8520 (N_8520,N_6713,N_7390);
nor U8521 (N_8521,N_6998,N_7480);
or U8522 (N_8522,N_6195,N_6457);
nor U8523 (N_8523,N_6478,N_5749);
and U8524 (N_8524,N_5898,N_7045);
and U8525 (N_8525,N_6553,N_6161);
nor U8526 (N_8526,N_6833,N_6504);
or U8527 (N_8527,N_7459,N_5726);
and U8528 (N_8528,N_7086,N_5519);
nand U8529 (N_8529,N_6444,N_6154);
or U8530 (N_8530,N_6061,N_6329);
nand U8531 (N_8531,N_7264,N_6341);
or U8532 (N_8532,N_6198,N_7247);
and U8533 (N_8533,N_6193,N_6689);
nor U8534 (N_8534,N_6090,N_5862);
and U8535 (N_8535,N_5801,N_5469);
nand U8536 (N_8536,N_5689,N_6229);
nand U8537 (N_8537,N_5613,N_6304);
and U8538 (N_8538,N_6466,N_6602);
nor U8539 (N_8539,N_6983,N_5681);
nand U8540 (N_8540,N_7137,N_5657);
nor U8541 (N_8541,N_6205,N_6666);
and U8542 (N_8542,N_6566,N_6940);
nor U8543 (N_8543,N_5232,N_6960);
and U8544 (N_8544,N_6586,N_6923);
or U8545 (N_8545,N_7122,N_7376);
nand U8546 (N_8546,N_5110,N_5744);
and U8547 (N_8547,N_6546,N_5894);
or U8548 (N_8548,N_7471,N_6652);
nand U8549 (N_8549,N_7304,N_5346);
nor U8550 (N_8550,N_7162,N_5676);
nand U8551 (N_8551,N_6675,N_5465);
or U8552 (N_8552,N_6522,N_6381);
nand U8553 (N_8553,N_6972,N_7164);
and U8554 (N_8554,N_6926,N_5578);
xor U8555 (N_8555,N_7001,N_5155);
nand U8556 (N_8556,N_5632,N_5768);
or U8557 (N_8557,N_6105,N_5682);
and U8558 (N_8558,N_5523,N_6919);
and U8559 (N_8559,N_6312,N_6212);
nand U8560 (N_8560,N_5766,N_6965);
nor U8561 (N_8561,N_5731,N_5442);
and U8562 (N_8562,N_5620,N_6337);
nand U8563 (N_8563,N_5301,N_6783);
nand U8564 (N_8564,N_6250,N_7099);
nor U8565 (N_8565,N_6269,N_7434);
nor U8566 (N_8566,N_5131,N_6574);
or U8567 (N_8567,N_6506,N_5864);
or U8568 (N_8568,N_6280,N_6836);
nor U8569 (N_8569,N_5875,N_6809);
nand U8570 (N_8570,N_6609,N_5799);
nand U8571 (N_8571,N_6920,N_5185);
or U8572 (N_8572,N_7148,N_6086);
or U8573 (N_8573,N_6938,N_6739);
and U8574 (N_8574,N_5762,N_5011);
and U8575 (N_8575,N_6728,N_7257);
nand U8576 (N_8576,N_5991,N_6199);
nor U8577 (N_8577,N_5905,N_5904);
nand U8578 (N_8578,N_6797,N_5481);
nand U8579 (N_8579,N_5506,N_6823);
nand U8580 (N_8580,N_5798,N_5552);
or U8581 (N_8581,N_7059,N_6159);
nand U8582 (N_8582,N_5895,N_5332);
and U8583 (N_8583,N_6123,N_6258);
and U8584 (N_8584,N_7290,N_6162);
nand U8585 (N_8585,N_6307,N_6166);
or U8586 (N_8586,N_7426,N_7469);
nand U8587 (N_8587,N_5080,N_5522);
or U8588 (N_8588,N_5227,N_5246);
nor U8589 (N_8589,N_7354,N_5460);
nand U8590 (N_8590,N_5518,N_5134);
nor U8591 (N_8591,N_6425,N_6411);
or U8592 (N_8592,N_6149,N_7444);
nor U8593 (N_8593,N_6737,N_5328);
and U8594 (N_8594,N_5692,N_6297);
or U8595 (N_8595,N_5909,N_6217);
nand U8596 (N_8596,N_6874,N_6922);
nand U8597 (N_8597,N_6234,N_6596);
nor U8598 (N_8598,N_7369,N_5265);
or U8599 (N_8599,N_6655,N_6074);
nand U8600 (N_8600,N_5807,N_6011);
nand U8601 (N_8601,N_5156,N_5787);
and U8602 (N_8602,N_5714,N_6530);
and U8603 (N_8603,N_7075,N_6073);
nand U8604 (N_8604,N_6462,N_6901);
nand U8605 (N_8605,N_5913,N_7184);
nor U8606 (N_8606,N_5049,N_6929);
nor U8607 (N_8607,N_5968,N_6994);
nand U8608 (N_8608,N_7437,N_5757);
and U8609 (N_8609,N_6840,N_6810);
nor U8610 (N_8610,N_6847,N_6495);
or U8611 (N_8611,N_6397,N_6499);
nand U8612 (N_8612,N_6539,N_5887);
nand U8613 (N_8613,N_5439,N_5300);
nand U8614 (N_8614,N_6266,N_6667);
nand U8615 (N_8615,N_7110,N_6717);
nand U8616 (N_8616,N_6491,N_5017);
and U8617 (N_8617,N_5355,N_5624);
nor U8618 (N_8618,N_6414,N_6132);
nand U8619 (N_8619,N_7002,N_7196);
or U8620 (N_8620,N_5842,N_5122);
and U8621 (N_8621,N_5190,N_6639);
nand U8622 (N_8622,N_6533,N_6963);
nor U8623 (N_8623,N_7102,N_6583);
nor U8624 (N_8624,N_6943,N_5290);
nand U8625 (N_8625,N_6038,N_5250);
and U8626 (N_8626,N_7326,N_5718);
and U8627 (N_8627,N_6095,N_6355);
and U8628 (N_8628,N_7096,N_5939);
and U8629 (N_8629,N_6968,N_5435);
and U8630 (N_8630,N_5298,N_6036);
and U8631 (N_8631,N_6855,N_5325);
nand U8632 (N_8632,N_6945,N_7008);
or U8633 (N_8633,N_6592,N_6812);
nand U8634 (N_8634,N_5773,N_6475);
or U8635 (N_8635,N_5767,N_7282);
nand U8636 (N_8636,N_6550,N_5478);
nor U8637 (N_8637,N_6971,N_6032);
and U8638 (N_8638,N_5543,N_6563);
or U8639 (N_8639,N_7239,N_6379);
or U8640 (N_8640,N_5179,N_6101);
or U8641 (N_8641,N_5513,N_6477);
and U8642 (N_8642,N_6990,N_6273);
nor U8643 (N_8643,N_6852,N_7220);
nand U8644 (N_8644,N_6528,N_5175);
and U8645 (N_8645,N_5678,N_5427);
and U8646 (N_8646,N_5516,N_5187);
or U8647 (N_8647,N_6338,N_6536);
or U8648 (N_8648,N_6201,N_5984);
nand U8649 (N_8649,N_7457,N_6017);
and U8650 (N_8650,N_7191,N_7176);
or U8651 (N_8651,N_7061,N_7181);
or U8652 (N_8652,N_6007,N_6127);
or U8653 (N_8653,N_7006,N_6401);
or U8654 (N_8654,N_5336,N_6881);
nand U8655 (N_8655,N_7097,N_5117);
nand U8656 (N_8656,N_6322,N_7248);
xor U8657 (N_8657,N_6885,N_5550);
nand U8658 (N_8658,N_6464,N_5459);
nor U8659 (N_8659,N_6080,N_7483);
or U8660 (N_8660,N_5845,N_6752);
and U8661 (N_8661,N_5084,N_6134);
nand U8662 (N_8662,N_6056,N_7460);
and U8663 (N_8663,N_5392,N_6898);
nor U8664 (N_8664,N_7051,N_6581);
or U8665 (N_8665,N_6402,N_6911);
and U8666 (N_8666,N_5008,N_6075);
and U8667 (N_8667,N_6340,N_5426);
xor U8668 (N_8668,N_5463,N_6350);
or U8669 (N_8669,N_5912,N_6942);
or U8670 (N_8670,N_5019,N_5512);
nand U8671 (N_8671,N_5420,N_5111);
or U8672 (N_8672,N_5811,N_5372);
xnor U8673 (N_8673,N_6175,N_5630);
nand U8674 (N_8674,N_5526,N_6869);
and U8675 (N_8675,N_6521,N_6009);
nand U8676 (N_8676,N_6461,N_5998);
or U8677 (N_8677,N_6318,N_7343);
nand U8678 (N_8678,N_7208,N_7310);
and U8679 (N_8679,N_7270,N_6939);
or U8680 (N_8680,N_5791,N_5326);
nor U8681 (N_8681,N_7432,N_5144);
and U8682 (N_8682,N_6415,N_5296);
nor U8683 (N_8683,N_6291,N_5859);
and U8684 (N_8684,N_5240,N_5231);
nor U8685 (N_8685,N_5321,N_6097);
nand U8686 (N_8686,N_6396,N_6674);
and U8687 (N_8687,N_5479,N_6143);
nand U8688 (N_8688,N_5373,N_6680);
nor U8689 (N_8689,N_7277,N_5878);
nand U8690 (N_8690,N_5685,N_5363);
nor U8691 (N_8691,N_6470,N_7084);
nand U8692 (N_8692,N_6440,N_6196);
or U8693 (N_8693,N_5958,N_6421);
nor U8694 (N_8694,N_7060,N_6119);
and U8695 (N_8695,N_5983,N_6138);
nand U8696 (N_8696,N_7388,N_7319);
nand U8697 (N_8697,N_6225,N_6432);
and U8698 (N_8698,N_6323,N_6749);
or U8699 (N_8699,N_5031,N_6146);
and U8700 (N_8700,N_5885,N_6694);
nand U8701 (N_8701,N_7030,N_6791);
nor U8702 (N_8702,N_5734,N_5367);
and U8703 (N_8703,N_5418,N_5498);
nand U8704 (N_8704,N_6981,N_6308);
and U8705 (N_8705,N_5780,N_5638);
or U8706 (N_8706,N_5544,N_6177);
and U8707 (N_8707,N_5727,N_6776);
nand U8708 (N_8708,N_5980,N_6698);
nor U8709 (N_8709,N_7487,N_6760);
nor U8710 (N_8710,N_6888,N_6610);
or U8711 (N_8711,N_6145,N_5691);
nand U8712 (N_8712,N_6252,N_5362);
nand U8713 (N_8713,N_5524,N_5299);
nor U8714 (N_8714,N_7490,N_6661);
nand U8715 (N_8715,N_5140,N_5323);
nand U8716 (N_8716,N_5819,N_5178);
nor U8717 (N_8717,N_7080,N_5614);
and U8718 (N_8718,N_5616,N_6380);
or U8719 (N_8719,N_5711,N_7082);
nand U8720 (N_8720,N_6626,N_7089);
nand U8721 (N_8721,N_7177,N_6000);
or U8722 (N_8722,N_6334,N_6896);
nand U8723 (N_8723,N_7275,N_6587);
or U8724 (N_8724,N_5229,N_6677);
and U8725 (N_8725,N_6620,N_5207);
nor U8726 (N_8726,N_7123,N_6125);
nand U8727 (N_8727,N_5572,N_5688);
and U8728 (N_8728,N_5100,N_5751);
or U8729 (N_8729,N_5452,N_5981);
and U8730 (N_8730,N_5038,N_6742);
and U8731 (N_8731,N_6598,N_6956);
or U8732 (N_8732,N_6311,N_6889);
and U8733 (N_8733,N_7477,N_7015);
nand U8734 (N_8734,N_5244,N_5194);
nand U8735 (N_8735,N_5295,N_5089);
nand U8736 (N_8736,N_5032,N_5351);
nand U8737 (N_8737,N_7224,N_7350);
and U8738 (N_8738,N_7374,N_6013);
nor U8739 (N_8739,N_5686,N_7192);
nor U8740 (N_8740,N_5588,N_5696);
and U8741 (N_8741,N_6155,N_5307);
nor U8742 (N_8742,N_6819,N_6081);
nand U8743 (N_8743,N_5477,N_7384);
nor U8744 (N_8744,N_6287,N_6946);
or U8745 (N_8745,N_6257,N_5521);
nor U8746 (N_8746,N_6830,N_7071);
or U8747 (N_8747,N_6623,N_6187);
or U8748 (N_8748,N_6479,N_6515);
or U8749 (N_8749,N_5579,N_6327);
and U8750 (N_8750,N_6375,N_7444);
or U8751 (N_8751,N_6192,N_6466);
or U8752 (N_8752,N_7240,N_7289);
and U8753 (N_8753,N_5138,N_7262);
and U8754 (N_8754,N_5626,N_6661);
or U8755 (N_8755,N_6578,N_7133);
and U8756 (N_8756,N_7064,N_5430);
nand U8757 (N_8757,N_7365,N_6829);
nand U8758 (N_8758,N_6330,N_5901);
or U8759 (N_8759,N_5275,N_7066);
nand U8760 (N_8760,N_5028,N_7413);
nor U8761 (N_8761,N_6390,N_6815);
nor U8762 (N_8762,N_7463,N_7159);
or U8763 (N_8763,N_5619,N_5049);
nand U8764 (N_8764,N_5373,N_5791);
and U8765 (N_8765,N_6362,N_5363);
or U8766 (N_8766,N_7256,N_6641);
nand U8767 (N_8767,N_6133,N_5693);
nand U8768 (N_8768,N_6388,N_7300);
nand U8769 (N_8769,N_5182,N_5366);
nor U8770 (N_8770,N_7316,N_6248);
or U8771 (N_8771,N_6589,N_5515);
or U8772 (N_8772,N_6897,N_7454);
nand U8773 (N_8773,N_7011,N_6938);
xnor U8774 (N_8774,N_5438,N_5227);
nand U8775 (N_8775,N_7058,N_5523);
and U8776 (N_8776,N_6039,N_6286);
and U8777 (N_8777,N_5800,N_6938);
and U8778 (N_8778,N_6000,N_6472);
and U8779 (N_8779,N_7343,N_5815);
xor U8780 (N_8780,N_7262,N_6202);
nand U8781 (N_8781,N_6616,N_5006);
and U8782 (N_8782,N_6510,N_6647);
nor U8783 (N_8783,N_6914,N_5203);
nand U8784 (N_8784,N_6530,N_6333);
or U8785 (N_8785,N_6063,N_7087);
or U8786 (N_8786,N_5226,N_5019);
or U8787 (N_8787,N_5975,N_5910);
nand U8788 (N_8788,N_6950,N_7103);
nor U8789 (N_8789,N_6307,N_6421);
and U8790 (N_8790,N_5215,N_5974);
or U8791 (N_8791,N_7171,N_5431);
nor U8792 (N_8792,N_7317,N_6126);
and U8793 (N_8793,N_7164,N_6200);
nand U8794 (N_8794,N_6887,N_6370);
or U8795 (N_8795,N_5589,N_5214);
nor U8796 (N_8796,N_7242,N_6776);
or U8797 (N_8797,N_7191,N_6260);
or U8798 (N_8798,N_5336,N_6454);
nor U8799 (N_8799,N_6646,N_7257);
nand U8800 (N_8800,N_6908,N_5497);
or U8801 (N_8801,N_5830,N_5642);
nor U8802 (N_8802,N_5527,N_7077);
nand U8803 (N_8803,N_6640,N_5237);
xnor U8804 (N_8804,N_6388,N_7179);
and U8805 (N_8805,N_7134,N_5823);
nor U8806 (N_8806,N_7328,N_7326);
and U8807 (N_8807,N_6140,N_5718);
and U8808 (N_8808,N_7428,N_6265);
nor U8809 (N_8809,N_7270,N_6853);
nor U8810 (N_8810,N_7404,N_5947);
or U8811 (N_8811,N_6004,N_6824);
nor U8812 (N_8812,N_5654,N_6760);
xor U8813 (N_8813,N_5100,N_5624);
or U8814 (N_8814,N_7322,N_7363);
and U8815 (N_8815,N_6611,N_7471);
nor U8816 (N_8816,N_6774,N_6921);
and U8817 (N_8817,N_7104,N_7241);
nand U8818 (N_8818,N_5297,N_5870);
nor U8819 (N_8819,N_5911,N_7369);
or U8820 (N_8820,N_6679,N_6787);
nand U8821 (N_8821,N_5893,N_7390);
nor U8822 (N_8822,N_5155,N_6861);
nand U8823 (N_8823,N_6582,N_6840);
or U8824 (N_8824,N_6290,N_6371);
nor U8825 (N_8825,N_7427,N_6408);
or U8826 (N_8826,N_7003,N_6588);
nand U8827 (N_8827,N_6406,N_7070);
nor U8828 (N_8828,N_7380,N_5042);
nor U8829 (N_8829,N_6524,N_5104);
nor U8830 (N_8830,N_6004,N_7012);
nand U8831 (N_8831,N_6238,N_5627);
nand U8832 (N_8832,N_7328,N_6291);
or U8833 (N_8833,N_7372,N_7304);
nor U8834 (N_8834,N_6814,N_7293);
nor U8835 (N_8835,N_5960,N_6172);
nor U8836 (N_8836,N_7253,N_5186);
and U8837 (N_8837,N_6039,N_7319);
or U8838 (N_8838,N_5584,N_6126);
nand U8839 (N_8839,N_6999,N_6179);
and U8840 (N_8840,N_6598,N_6020);
nand U8841 (N_8841,N_6040,N_5461);
or U8842 (N_8842,N_5051,N_6413);
and U8843 (N_8843,N_6479,N_6119);
or U8844 (N_8844,N_6411,N_5895);
nand U8845 (N_8845,N_6323,N_5674);
and U8846 (N_8846,N_6790,N_7099);
and U8847 (N_8847,N_6097,N_6428);
or U8848 (N_8848,N_5482,N_7329);
or U8849 (N_8849,N_5024,N_6015);
nand U8850 (N_8850,N_7200,N_6161);
nand U8851 (N_8851,N_6090,N_5029);
nand U8852 (N_8852,N_5556,N_5593);
and U8853 (N_8853,N_5268,N_6154);
or U8854 (N_8854,N_6597,N_6116);
and U8855 (N_8855,N_7133,N_5370);
and U8856 (N_8856,N_6753,N_5162);
nor U8857 (N_8857,N_5267,N_6407);
nor U8858 (N_8858,N_6401,N_6054);
nand U8859 (N_8859,N_6748,N_6549);
nand U8860 (N_8860,N_6496,N_6554);
nand U8861 (N_8861,N_5709,N_5139);
or U8862 (N_8862,N_7417,N_5053);
nor U8863 (N_8863,N_5946,N_6479);
and U8864 (N_8864,N_7391,N_6157);
and U8865 (N_8865,N_6410,N_7132);
nor U8866 (N_8866,N_6848,N_5961);
and U8867 (N_8867,N_5689,N_6731);
nor U8868 (N_8868,N_7317,N_7112);
nand U8869 (N_8869,N_5950,N_5193);
and U8870 (N_8870,N_6215,N_6212);
nand U8871 (N_8871,N_6916,N_6047);
nand U8872 (N_8872,N_6950,N_6482);
xor U8873 (N_8873,N_5028,N_6198);
or U8874 (N_8874,N_5454,N_6592);
and U8875 (N_8875,N_5503,N_5907);
and U8876 (N_8876,N_7487,N_5335);
nor U8877 (N_8877,N_7274,N_7057);
or U8878 (N_8878,N_6487,N_5696);
xnor U8879 (N_8879,N_6321,N_6179);
nor U8880 (N_8880,N_7023,N_6956);
and U8881 (N_8881,N_5010,N_6852);
and U8882 (N_8882,N_7090,N_5917);
or U8883 (N_8883,N_5118,N_6951);
and U8884 (N_8884,N_6336,N_5496);
nand U8885 (N_8885,N_6100,N_7270);
nand U8886 (N_8886,N_6325,N_5066);
or U8887 (N_8887,N_6649,N_6751);
and U8888 (N_8888,N_6843,N_5370);
nand U8889 (N_8889,N_6685,N_5641);
nor U8890 (N_8890,N_6721,N_7426);
and U8891 (N_8891,N_5205,N_6966);
and U8892 (N_8892,N_6455,N_6779);
and U8893 (N_8893,N_7065,N_6537);
or U8894 (N_8894,N_5312,N_6617);
nand U8895 (N_8895,N_7321,N_6480);
and U8896 (N_8896,N_6817,N_6814);
and U8897 (N_8897,N_6342,N_5007);
or U8898 (N_8898,N_5198,N_6523);
xnor U8899 (N_8899,N_7155,N_5589);
and U8900 (N_8900,N_5930,N_6412);
and U8901 (N_8901,N_7255,N_5564);
or U8902 (N_8902,N_5549,N_7003);
and U8903 (N_8903,N_5554,N_5479);
or U8904 (N_8904,N_5624,N_7479);
nand U8905 (N_8905,N_6238,N_5502);
or U8906 (N_8906,N_7211,N_6858);
nand U8907 (N_8907,N_6424,N_7064);
and U8908 (N_8908,N_6985,N_6994);
and U8909 (N_8909,N_6014,N_6122);
nand U8910 (N_8910,N_5245,N_7260);
or U8911 (N_8911,N_5740,N_6539);
nand U8912 (N_8912,N_6624,N_5924);
and U8913 (N_8913,N_7427,N_7210);
nor U8914 (N_8914,N_5110,N_6775);
and U8915 (N_8915,N_7359,N_5665);
xnor U8916 (N_8916,N_6488,N_6664);
nor U8917 (N_8917,N_6960,N_5772);
nor U8918 (N_8918,N_7425,N_6165);
nor U8919 (N_8919,N_5341,N_6750);
and U8920 (N_8920,N_6476,N_5366);
or U8921 (N_8921,N_5652,N_6432);
and U8922 (N_8922,N_5439,N_5869);
nand U8923 (N_8923,N_5087,N_7145);
nor U8924 (N_8924,N_6215,N_6499);
and U8925 (N_8925,N_7017,N_5592);
or U8926 (N_8926,N_5532,N_6415);
or U8927 (N_8927,N_7177,N_5419);
and U8928 (N_8928,N_5438,N_5600);
or U8929 (N_8929,N_7296,N_5433);
nor U8930 (N_8930,N_5631,N_5495);
or U8931 (N_8931,N_6247,N_5822);
or U8932 (N_8932,N_5452,N_6836);
or U8933 (N_8933,N_6411,N_5651);
nand U8934 (N_8934,N_5176,N_5086);
and U8935 (N_8935,N_5499,N_7397);
or U8936 (N_8936,N_6630,N_6195);
and U8937 (N_8937,N_6478,N_7359);
nor U8938 (N_8938,N_5387,N_6757);
nand U8939 (N_8939,N_5794,N_6795);
nor U8940 (N_8940,N_7248,N_6943);
and U8941 (N_8941,N_6561,N_6374);
and U8942 (N_8942,N_6017,N_6030);
nand U8943 (N_8943,N_6706,N_5070);
or U8944 (N_8944,N_6906,N_6293);
nor U8945 (N_8945,N_6232,N_5034);
nor U8946 (N_8946,N_5855,N_6690);
or U8947 (N_8947,N_5781,N_7320);
nor U8948 (N_8948,N_5155,N_6508);
or U8949 (N_8949,N_6431,N_6240);
xor U8950 (N_8950,N_5919,N_5544);
nor U8951 (N_8951,N_5747,N_7086);
nor U8952 (N_8952,N_7162,N_6872);
and U8953 (N_8953,N_5063,N_5509);
or U8954 (N_8954,N_6151,N_6905);
xnor U8955 (N_8955,N_6848,N_6490);
and U8956 (N_8956,N_5688,N_7159);
and U8957 (N_8957,N_5098,N_6247);
nor U8958 (N_8958,N_5525,N_6201);
nor U8959 (N_8959,N_5697,N_5169);
nand U8960 (N_8960,N_6570,N_5490);
and U8961 (N_8961,N_6076,N_7464);
nor U8962 (N_8962,N_5041,N_6569);
nor U8963 (N_8963,N_7016,N_6136);
and U8964 (N_8964,N_6289,N_7327);
nor U8965 (N_8965,N_6102,N_6472);
nor U8966 (N_8966,N_6573,N_5214);
nand U8967 (N_8967,N_7385,N_7429);
xor U8968 (N_8968,N_7322,N_5066);
xor U8969 (N_8969,N_6214,N_5542);
and U8970 (N_8970,N_6040,N_6392);
nor U8971 (N_8971,N_5073,N_7216);
and U8972 (N_8972,N_5225,N_5376);
xor U8973 (N_8973,N_5150,N_5060);
or U8974 (N_8974,N_5121,N_6764);
nand U8975 (N_8975,N_5877,N_7382);
and U8976 (N_8976,N_5750,N_6768);
and U8977 (N_8977,N_6208,N_7138);
nand U8978 (N_8978,N_5133,N_5801);
or U8979 (N_8979,N_6087,N_6196);
and U8980 (N_8980,N_6629,N_6437);
xor U8981 (N_8981,N_5968,N_6599);
or U8982 (N_8982,N_5017,N_6114);
or U8983 (N_8983,N_6742,N_5963);
nand U8984 (N_8984,N_6895,N_5535);
or U8985 (N_8985,N_6783,N_5433);
and U8986 (N_8986,N_6509,N_6208);
nand U8987 (N_8987,N_5999,N_6895);
or U8988 (N_8988,N_6037,N_6653);
nand U8989 (N_8989,N_6372,N_7355);
or U8990 (N_8990,N_6793,N_6086);
and U8991 (N_8991,N_5345,N_5261);
nand U8992 (N_8992,N_7109,N_5475);
xnor U8993 (N_8993,N_5129,N_7272);
or U8994 (N_8994,N_6771,N_7419);
nand U8995 (N_8995,N_7460,N_7298);
and U8996 (N_8996,N_6297,N_6779);
nor U8997 (N_8997,N_5848,N_5512);
or U8998 (N_8998,N_5059,N_7405);
and U8999 (N_8999,N_6113,N_6043);
nor U9000 (N_9000,N_5008,N_5395);
or U9001 (N_9001,N_5720,N_5345);
and U9002 (N_9002,N_6972,N_5775);
or U9003 (N_9003,N_5078,N_5111);
and U9004 (N_9004,N_7008,N_6905);
nor U9005 (N_9005,N_7391,N_7062);
xor U9006 (N_9006,N_7079,N_6765);
or U9007 (N_9007,N_6474,N_6957);
and U9008 (N_9008,N_7208,N_5208);
or U9009 (N_9009,N_5539,N_5079);
or U9010 (N_9010,N_6389,N_5103);
nand U9011 (N_9011,N_5993,N_7041);
nor U9012 (N_9012,N_7446,N_6662);
or U9013 (N_9013,N_6974,N_6440);
or U9014 (N_9014,N_7266,N_5879);
nor U9015 (N_9015,N_5403,N_6198);
nand U9016 (N_9016,N_5803,N_5356);
and U9017 (N_9017,N_5637,N_5957);
xor U9018 (N_9018,N_5959,N_6249);
and U9019 (N_9019,N_6938,N_6707);
and U9020 (N_9020,N_5237,N_5372);
and U9021 (N_9021,N_6838,N_5679);
nor U9022 (N_9022,N_6327,N_7217);
and U9023 (N_9023,N_6813,N_5105);
nor U9024 (N_9024,N_5469,N_6140);
and U9025 (N_9025,N_5366,N_5463);
nor U9026 (N_9026,N_6400,N_5391);
nor U9027 (N_9027,N_6271,N_6744);
or U9028 (N_9028,N_6499,N_7029);
and U9029 (N_9029,N_6231,N_5433);
and U9030 (N_9030,N_5310,N_6888);
nor U9031 (N_9031,N_6683,N_6769);
and U9032 (N_9032,N_6662,N_6383);
or U9033 (N_9033,N_7051,N_7090);
and U9034 (N_9034,N_6665,N_6243);
xor U9035 (N_9035,N_5941,N_5157);
nand U9036 (N_9036,N_6441,N_6661);
and U9037 (N_9037,N_7260,N_6570);
nand U9038 (N_9038,N_5787,N_6814);
and U9039 (N_9039,N_6681,N_5778);
nand U9040 (N_9040,N_5184,N_6760);
or U9041 (N_9041,N_6318,N_7292);
and U9042 (N_9042,N_5804,N_6287);
and U9043 (N_9043,N_7246,N_6424);
nor U9044 (N_9044,N_7151,N_7250);
nor U9045 (N_9045,N_5640,N_7078);
nor U9046 (N_9046,N_5930,N_7287);
nor U9047 (N_9047,N_6690,N_5306);
and U9048 (N_9048,N_6907,N_6285);
or U9049 (N_9049,N_7218,N_6268);
nand U9050 (N_9050,N_6144,N_6311);
and U9051 (N_9051,N_6830,N_7202);
nand U9052 (N_9052,N_6581,N_7146);
or U9053 (N_9053,N_5667,N_5754);
and U9054 (N_9054,N_6286,N_6938);
or U9055 (N_9055,N_6516,N_7013);
nand U9056 (N_9056,N_6176,N_5418);
nand U9057 (N_9057,N_6679,N_6559);
nand U9058 (N_9058,N_6079,N_5808);
or U9059 (N_9059,N_6639,N_6931);
or U9060 (N_9060,N_6044,N_7255);
nor U9061 (N_9061,N_5943,N_6393);
or U9062 (N_9062,N_5305,N_6349);
and U9063 (N_9063,N_7107,N_5130);
or U9064 (N_9064,N_6035,N_7088);
and U9065 (N_9065,N_6164,N_6036);
or U9066 (N_9066,N_5585,N_5054);
nor U9067 (N_9067,N_5783,N_7495);
or U9068 (N_9068,N_5147,N_6334);
and U9069 (N_9069,N_6579,N_5178);
and U9070 (N_9070,N_5110,N_7322);
nor U9071 (N_9071,N_6660,N_7309);
nor U9072 (N_9072,N_5744,N_5784);
nor U9073 (N_9073,N_5295,N_7376);
nand U9074 (N_9074,N_5963,N_7292);
or U9075 (N_9075,N_5025,N_5079);
or U9076 (N_9076,N_5224,N_5114);
nand U9077 (N_9077,N_6969,N_5734);
and U9078 (N_9078,N_5037,N_7184);
nand U9079 (N_9079,N_6075,N_6457);
or U9080 (N_9080,N_6990,N_5592);
nand U9081 (N_9081,N_5243,N_6131);
and U9082 (N_9082,N_5063,N_5534);
nor U9083 (N_9083,N_6937,N_6047);
and U9084 (N_9084,N_5317,N_6077);
xor U9085 (N_9085,N_7356,N_5819);
or U9086 (N_9086,N_6984,N_6589);
and U9087 (N_9087,N_6957,N_7056);
or U9088 (N_9088,N_6820,N_5216);
and U9089 (N_9089,N_5133,N_7072);
and U9090 (N_9090,N_6823,N_6437);
and U9091 (N_9091,N_5948,N_6503);
nand U9092 (N_9092,N_7201,N_5818);
nand U9093 (N_9093,N_6306,N_6898);
nor U9094 (N_9094,N_6473,N_6796);
or U9095 (N_9095,N_7282,N_5428);
nor U9096 (N_9096,N_6708,N_5680);
nor U9097 (N_9097,N_6928,N_6981);
nor U9098 (N_9098,N_5172,N_5029);
or U9099 (N_9099,N_5296,N_5790);
nand U9100 (N_9100,N_7248,N_5693);
nand U9101 (N_9101,N_5616,N_6300);
or U9102 (N_9102,N_6083,N_7102);
or U9103 (N_9103,N_5996,N_7233);
nor U9104 (N_9104,N_6797,N_6875);
or U9105 (N_9105,N_7086,N_6356);
nor U9106 (N_9106,N_7001,N_5034);
nand U9107 (N_9107,N_5849,N_6636);
nand U9108 (N_9108,N_7493,N_6569);
or U9109 (N_9109,N_5200,N_7394);
nor U9110 (N_9110,N_6729,N_6399);
nor U9111 (N_9111,N_6722,N_5008);
nor U9112 (N_9112,N_6647,N_6567);
nand U9113 (N_9113,N_6033,N_5850);
nor U9114 (N_9114,N_7192,N_5444);
nor U9115 (N_9115,N_6453,N_7173);
or U9116 (N_9116,N_6764,N_5399);
nand U9117 (N_9117,N_6314,N_5948);
xnor U9118 (N_9118,N_6377,N_5708);
and U9119 (N_9119,N_6831,N_5382);
and U9120 (N_9120,N_6725,N_6004);
or U9121 (N_9121,N_6054,N_5863);
and U9122 (N_9122,N_5315,N_6671);
or U9123 (N_9123,N_7425,N_6887);
and U9124 (N_9124,N_5604,N_5044);
nand U9125 (N_9125,N_5081,N_7149);
nor U9126 (N_9126,N_5868,N_7262);
and U9127 (N_9127,N_7021,N_5228);
nand U9128 (N_9128,N_7209,N_6803);
nor U9129 (N_9129,N_6971,N_6364);
nand U9130 (N_9130,N_5596,N_6372);
nor U9131 (N_9131,N_6548,N_6710);
nor U9132 (N_9132,N_6003,N_6800);
nor U9133 (N_9133,N_6416,N_7293);
nand U9134 (N_9134,N_5517,N_6065);
nor U9135 (N_9135,N_7014,N_5049);
and U9136 (N_9136,N_6097,N_7397);
or U9137 (N_9137,N_5438,N_5234);
nor U9138 (N_9138,N_5773,N_6912);
nand U9139 (N_9139,N_6264,N_5434);
and U9140 (N_9140,N_6040,N_5833);
and U9141 (N_9141,N_5180,N_5048);
nor U9142 (N_9142,N_7100,N_6277);
nand U9143 (N_9143,N_6376,N_7443);
nand U9144 (N_9144,N_5153,N_5188);
or U9145 (N_9145,N_6286,N_7252);
nor U9146 (N_9146,N_6786,N_5307);
and U9147 (N_9147,N_7391,N_6638);
and U9148 (N_9148,N_6655,N_6707);
nor U9149 (N_9149,N_7184,N_7409);
or U9150 (N_9150,N_6225,N_6596);
nor U9151 (N_9151,N_5137,N_7260);
nor U9152 (N_9152,N_6413,N_6914);
nand U9153 (N_9153,N_6631,N_5517);
or U9154 (N_9154,N_5950,N_6984);
nor U9155 (N_9155,N_5504,N_5722);
nor U9156 (N_9156,N_7055,N_5716);
nand U9157 (N_9157,N_7355,N_7098);
xor U9158 (N_9158,N_6125,N_6731);
nand U9159 (N_9159,N_6514,N_6376);
and U9160 (N_9160,N_5250,N_5088);
nor U9161 (N_9161,N_5143,N_6257);
nand U9162 (N_9162,N_5910,N_5509);
and U9163 (N_9163,N_5480,N_5819);
and U9164 (N_9164,N_6279,N_6520);
nand U9165 (N_9165,N_5844,N_6726);
and U9166 (N_9166,N_6428,N_7254);
nand U9167 (N_9167,N_6274,N_5101);
nand U9168 (N_9168,N_5899,N_7005);
or U9169 (N_9169,N_5431,N_7056);
or U9170 (N_9170,N_5599,N_5885);
nand U9171 (N_9171,N_7412,N_6890);
nor U9172 (N_9172,N_6306,N_5271);
or U9173 (N_9173,N_5532,N_6758);
and U9174 (N_9174,N_7090,N_6534);
and U9175 (N_9175,N_6601,N_6353);
nor U9176 (N_9176,N_5405,N_6286);
and U9177 (N_9177,N_5721,N_6562);
and U9178 (N_9178,N_5900,N_6958);
or U9179 (N_9179,N_6312,N_5432);
nand U9180 (N_9180,N_6770,N_6732);
nor U9181 (N_9181,N_6113,N_5965);
nor U9182 (N_9182,N_7358,N_6904);
nand U9183 (N_9183,N_7246,N_5352);
nor U9184 (N_9184,N_7440,N_6116);
nor U9185 (N_9185,N_5011,N_6822);
nor U9186 (N_9186,N_6365,N_6031);
nand U9187 (N_9187,N_5394,N_6199);
nand U9188 (N_9188,N_7223,N_6657);
and U9189 (N_9189,N_5936,N_7418);
and U9190 (N_9190,N_6474,N_5154);
or U9191 (N_9191,N_7389,N_7484);
and U9192 (N_9192,N_5582,N_5940);
and U9193 (N_9193,N_7384,N_6266);
nand U9194 (N_9194,N_5166,N_6786);
nor U9195 (N_9195,N_6045,N_5494);
xor U9196 (N_9196,N_5791,N_6049);
and U9197 (N_9197,N_5942,N_5646);
and U9198 (N_9198,N_7376,N_6996);
xnor U9199 (N_9199,N_6017,N_7403);
or U9200 (N_9200,N_6586,N_6709);
and U9201 (N_9201,N_7139,N_5092);
or U9202 (N_9202,N_6377,N_5562);
and U9203 (N_9203,N_6997,N_6535);
nor U9204 (N_9204,N_6774,N_6038);
nor U9205 (N_9205,N_6970,N_6883);
nor U9206 (N_9206,N_6940,N_5747);
nand U9207 (N_9207,N_5819,N_6198);
or U9208 (N_9208,N_6689,N_6931);
or U9209 (N_9209,N_7308,N_5341);
nor U9210 (N_9210,N_6099,N_5007);
nor U9211 (N_9211,N_5198,N_5979);
or U9212 (N_9212,N_7471,N_6946);
nor U9213 (N_9213,N_5200,N_6396);
and U9214 (N_9214,N_6356,N_7347);
or U9215 (N_9215,N_5519,N_5749);
and U9216 (N_9216,N_7244,N_6636);
nor U9217 (N_9217,N_6751,N_5550);
and U9218 (N_9218,N_5707,N_6748);
nand U9219 (N_9219,N_5520,N_6661);
and U9220 (N_9220,N_6414,N_5190);
and U9221 (N_9221,N_5469,N_6839);
and U9222 (N_9222,N_5140,N_6422);
and U9223 (N_9223,N_6399,N_5262);
nand U9224 (N_9224,N_7292,N_6019);
or U9225 (N_9225,N_6002,N_5669);
or U9226 (N_9226,N_5799,N_7065);
or U9227 (N_9227,N_5482,N_6530);
nor U9228 (N_9228,N_5850,N_6316);
or U9229 (N_9229,N_6650,N_6761);
nand U9230 (N_9230,N_6674,N_6068);
and U9231 (N_9231,N_6606,N_7068);
nor U9232 (N_9232,N_5655,N_6153);
and U9233 (N_9233,N_6609,N_6940);
nor U9234 (N_9234,N_7223,N_6831);
nand U9235 (N_9235,N_6657,N_7213);
nor U9236 (N_9236,N_6240,N_5592);
or U9237 (N_9237,N_6731,N_5301);
nand U9238 (N_9238,N_5048,N_7375);
nand U9239 (N_9239,N_6170,N_7493);
or U9240 (N_9240,N_5446,N_5384);
nand U9241 (N_9241,N_7020,N_5082);
nor U9242 (N_9242,N_5535,N_5451);
or U9243 (N_9243,N_7404,N_6353);
and U9244 (N_9244,N_5966,N_5196);
nand U9245 (N_9245,N_6707,N_7359);
or U9246 (N_9246,N_5987,N_5250);
or U9247 (N_9247,N_6861,N_6518);
or U9248 (N_9248,N_6631,N_5259);
and U9249 (N_9249,N_6002,N_6108);
and U9250 (N_9250,N_6479,N_6105);
or U9251 (N_9251,N_5644,N_5454);
or U9252 (N_9252,N_5802,N_5603);
or U9253 (N_9253,N_7172,N_6567);
and U9254 (N_9254,N_6466,N_6188);
nor U9255 (N_9255,N_7168,N_6613);
nand U9256 (N_9256,N_6902,N_5883);
and U9257 (N_9257,N_5692,N_5656);
xnor U9258 (N_9258,N_5441,N_5164);
and U9259 (N_9259,N_6785,N_6160);
nor U9260 (N_9260,N_7179,N_5538);
nor U9261 (N_9261,N_6541,N_6219);
and U9262 (N_9262,N_7113,N_6983);
nand U9263 (N_9263,N_6567,N_7386);
and U9264 (N_9264,N_6271,N_5376);
nand U9265 (N_9265,N_5774,N_5440);
and U9266 (N_9266,N_5762,N_6005);
or U9267 (N_9267,N_5023,N_5932);
and U9268 (N_9268,N_5521,N_7086);
nor U9269 (N_9269,N_6631,N_5333);
xnor U9270 (N_9270,N_7274,N_6977);
nand U9271 (N_9271,N_6057,N_7389);
nor U9272 (N_9272,N_7204,N_6370);
and U9273 (N_9273,N_7175,N_5699);
xnor U9274 (N_9274,N_7006,N_7340);
nand U9275 (N_9275,N_5370,N_6294);
and U9276 (N_9276,N_7183,N_5941);
nor U9277 (N_9277,N_7102,N_7152);
or U9278 (N_9278,N_5755,N_6072);
nor U9279 (N_9279,N_5250,N_7308);
nand U9280 (N_9280,N_6791,N_7304);
nor U9281 (N_9281,N_5695,N_6696);
nand U9282 (N_9282,N_5226,N_6012);
nor U9283 (N_9283,N_5136,N_6272);
nand U9284 (N_9284,N_6363,N_6515);
or U9285 (N_9285,N_7336,N_7207);
nand U9286 (N_9286,N_7418,N_7136);
and U9287 (N_9287,N_5298,N_5944);
and U9288 (N_9288,N_6619,N_5937);
xnor U9289 (N_9289,N_6661,N_7352);
nand U9290 (N_9290,N_7107,N_6195);
nor U9291 (N_9291,N_5759,N_5501);
nor U9292 (N_9292,N_7201,N_6807);
nor U9293 (N_9293,N_7040,N_5708);
nor U9294 (N_9294,N_7260,N_6254);
or U9295 (N_9295,N_5232,N_7415);
or U9296 (N_9296,N_7187,N_5396);
or U9297 (N_9297,N_6422,N_5995);
and U9298 (N_9298,N_5219,N_5300);
nor U9299 (N_9299,N_5854,N_6398);
and U9300 (N_9300,N_5753,N_5965);
nand U9301 (N_9301,N_6113,N_5087);
nor U9302 (N_9302,N_7383,N_7126);
nand U9303 (N_9303,N_6718,N_5169);
and U9304 (N_9304,N_7273,N_5288);
nand U9305 (N_9305,N_5002,N_6518);
or U9306 (N_9306,N_5001,N_5618);
or U9307 (N_9307,N_5918,N_7086);
nor U9308 (N_9308,N_7094,N_7026);
and U9309 (N_9309,N_5348,N_5535);
or U9310 (N_9310,N_5394,N_5234);
and U9311 (N_9311,N_6760,N_7003);
and U9312 (N_9312,N_5917,N_6581);
nor U9313 (N_9313,N_7309,N_5395);
and U9314 (N_9314,N_7031,N_6010);
nor U9315 (N_9315,N_5939,N_6935);
xnor U9316 (N_9316,N_6234,N_7408);
or U9317 (N_9317,N_5988,N_6407);
nand U9318 (N_9318,N_6635,N_7192);
and U9319 (N_9319,N_5390,N_5738);
and U9320 (N_9320,N_6952,N_6342);
and U9321 (N_9321,N_7186,N_5713);
nor U9322 (N_9322,N_5034,N_5203);
nand U9323 (N_9323,N_7429,N_6926);
or U9324 (N_9324,N_6610,N_6822);
and U9325 (N_9325,N_5488,N_5018);
nand U9326 (N_9326,N_7152,N_5571);
nor U9327 (N_9327,N_6709,N_5296);
and U9328 (N_9328,N_5383,N_5945);
and U9329 (N_9329,N_5926,N_6830);
and U9330 (N_9330,N_6643,N_5888);
or U9331 (N_9331,N_5868,N_6675);
nand U9332 (N_9332,N_6015,N_6238);
nor U9333 (N_9333,N_5531,N_7104);
nand U9334 (N_9334,N_6026,N_7119);
nor U9335 (N_9335,N_5592,N_6331);
nor U9336 (N_9336,N_6513,N_7295);
nor U9337 (N_9337,N_5516,N_6778);
xnor U9338 (N_9338,N_6569,N_7219);
nand U9339 (N_9339,N_5192,N_5785);
nand U9340 (N_9340,N_5276,N_5185);
nand U9341 (N_9341,N_6461,N_5485);
nand U9342 (N_9342,N_6410,N_6101);
nor U9343 (N_9343,N_6481,N_6705);
nor U9344 (N_9344,N_6016,N_7058);
and U9345 (N_9345,N_7394,N_6859);
nor U9346 (N_9346,N_5839,N_6720);
nand U9347 (N_9347,N_7088,N_7205);
and U9348 (N_9348,N_6672,N_5285);
or U9349 (N_9349,N_5579,N_5333);
nand U9350 (N_9350,N_5376,N_7480);
nand U9351 (N_9351,N_6375,N_6152);
nor U9352 (N_9352,N_7111,N_7444);
nand U9353 (N_9353,N_6546,N_6658);
and U9354 (N_9354,N_6359,N_7282);
nand U9355 (N_9355,N_5892,N_6657);
nor U9356 (N_9356,N_6072,N_6356);
and U9357 (N_9357,N_5884,N_5622);
or U9358 (N_9358,N_5091,N_7493);
and U9359 (N_9359,N_5014,N_6634);
nand U9360 (N_9360,N_5796,N_7082);
nand U9361 (N_9361,N_5369,N_6524);
and U9362 (N_9362,N_5505,N_5223);
or U9363 (N_9363,N_7364,N_5872);
and U9364 (N_9364,N_6548,N_6274);
nor U9365 (N_9365,N_5001,N_5858);
nor U9366 (N_9366,N_6686,N_7224);
or U9367 (N_9367,N_5346,N_7243);
xor U9368 (N_9368,N_6944,N_6919);
and U9369 (N_9369,N_5638,N_6805);
or U9370 (N_9370,N_6147,N_6026);
nor U9371 (N_9371,N_7004,N_5012);
nand U9372 (N_9372,N_6821,N_7120);
and U9373 (N_9373,N_7207,N_6046);
nor U9374 (N_9374,N_5905,N_5549);
and U9375 (N_9375,N_5129,N_6105);
nand U9376 (N_9376,N_7277,N_6682);
nand U9377 (N_9377,N_6023,N_7240);
and U9378 (N_9378,N_6730,N_6807);
or U9379 (N_9379,N_6887,N_5359);
and U9380 (N_9380,N_6607,N_6572);
or U9381 (N_9381,N_5292,N_6648);
nor U9382 (N_9382,N_6259,N_6345);
nand U9383 (N_9383,N_6320,N_6207);
nor U9384 (N_9384,N_6717,N_5364);
xnor U9385 (N_9385,N_6013,N_6837);
nor U9386 (N_9386,N_5211,N_7342);
nand U9387 (N_9387,N_6900,N_6101);
and U9388 (N_9388,N_7121,N_5611);
and U9389 (N_9389,N_6299,N_6417);
and U9390 (N_9390,N_6041,N_6551);
or U9391 (N_9391,N_6018,N_6761);
or U9392 (N_9392,N_6185,N_7373);
or U9393 (N_9393,N_7062,N_5870);
nand U9394 (N_9394,N_6927,N_5244);
or U9395 (N_9395,N_6513,N_6937);
nand U9396 (N_9396,N_6671,N_6308);
and U9397 (N_9397,N_6036,N_5712);
or U9398 (N_9398,N_6653,N_5480);
and U9399 (N_9399,N_6531,N_5695);
and U9400 (N_9400,N_6769,N_7436);
nand U9401 (N_9401,N_5948,N_5849);
and U9402 (N_9402,N_7026,N_6590);
xnor U9403 (N_9403,N_5172,N_6796);
and U9404 (N_9404,N_6791,N_6748);
and U9405 (N_9405,N_5788,N_7477);
or U9406 (N_9406,N_7089,N_7247);
nor U9407 (N_9407,N_6515,N_6144);
or U9408 (N_9408,N_5695,N_6981);
or U9409 (N_9409,N_7310,N_6109);
nor U9410 (N_9410,N_5104,N_5517);
and U9411 (N_9411,N_6488,N_5321);
or U9412 (N_9412,N_7087,N_7263);
or U9413 (N_9413,N_6395,N_6914);
nor U9414 (N_9414,N_5797,N_6417);
nor U9415 (N_9415,N_5973,N_6454);
and U9416 (N_9416,N_7022,N_7349);
nand U9417 (N_9417,N_5719,N_7408);
and U9418 (N_9418,N_5576,N_5420);
and U9419 (N_9419,N_7247,N_5776);
xor U9420 (N_9420,N_5793,N_5392);
or U9421 (N_9421,N_6613,N_5759);
nand U9422 (N_9422,N_6393,N_6978);
nor U9423 (N_9423,N_6889,N_6325);
nor U9424 (N_9424,N_6102,N_6017);
nand U9425 (N_9425,N_5473,N_6635);
or U9426 (N_9426,N_6832,N_6189);
or U9427 (N_9427,N_7219,N_7114);
or U9428 (N_9428,N_7276,N_5008);
nor U9429 (N_9429,N_7388,N_6754);
nand U9430 (N_9430,N_6461,N_5707);
or U9431 (N_9431,N_5831,N_7435);
nor U9432 (N_9432,N_5110,N_6862);
nor U9433 (N_9433,N_5333,N_7276);
and U9434 (N_9434,N_7085,N_6962);
and U9435 (N_9435,N_6564,N_5627);
or U9436 (N_9436,N_6947,N_7484);
and U9437 (N_9437,N_5366,N_6596);
nor U9438 (N_9438,N_5733,N_6249);
nand U9439 (N_9439,N_5435,N_5214);
and U9440 (N_9440,N_5583,N_6935);
or U9441 (N_9441,N_6790,N_5711);
nand U9442 (N_9442,N_7489,N_6297);
nor U9443 (N_9443,N_5184,N_5538);
and U9444 (N_9444,N_5568,N_6643);
and U9445 (N_9445,N_6799,N_6116);
or U9446 (N_9446,N_6706,N_6634);
and U9447 (N_9447,N_6236,N_5248);
nand U9448 (N_9448,N_5113,N_6026);
nor U9449 (N_9449,N_6151,N_5098);
nand U9450 (N_9450,N_7009,N_6401);
nand U9451 (N_9451,N_7443,N_5985);
or U9452 (N_9452,N_6822,N_7236);
nor U9453 (N_9453,N_6751,N_5130);
nor U9454 (N_9454,N_6576,N_5484);
nand U9455 (N_9455,N_6670,N_5084);
and U9456 (N_9456,N_6400,N_5935);
or U9457 (N_9457,N_6093,N_5052);
nand U9458 (N_9458,N_6441,N_6724);
nand U9459 (N_9459,N_6277,N_5495);
or U9460 (N_9460,N_5733,N_7173);
nand U9461 (N_9461,N_5067,N_6049);
or U9462 (N_9462,N_6900,N_6490);
xor U9463 (N_9463,N_5395,N_5233);
and U9464 (N_9464,N_5228,N_5253);
or U9465 (N_9465,N_7303,N_5972);
nand U9466 (N_9466,N_6441,N_5608);
or U9467 (N_9467,N_5899,N_5812);
or U9468 (N_9468,N_7243,N_6111);
or U9469 (N_9469,N_5005,N_7415);
and U9470 (N_9470,N_6584,N_6269);
xnor U9471 (N_9471,N_7126,N_5076);
or U9472 (N_9472,N_7214,N_6256);
or U9473 (N_9473,N_6689,N_5718);
nor U9474 (N_9474,N_5086,N_6913);
nand U9475 (N_9475,N_7275,N_5960);
nor U9476 (N_9476,N_6199,N_6870);
and U9477 (N_9477,N_6163,N_7365);
nor U9478 (N_9478,N_5182,N_5197);
nand U9479 (N_9479,N_6791,N_6599);
or U9480 (N_9480,N_5197,N_6652);
and U9481 (N_9481,N_5876,N_6802);
nor U9482 (N_9482,N_5132,N_6981);
and U9483 (N_9483,N_7170,N_5797);
nor U9484 (N_9484,N_5235,N_5829);
nor U9485 (N_9485,N_7495,N_5170);
and U9486 (N_9486,N_7023,N_6703);
and U9487 (N_9487,N_7064,N_5465);
and U9488 (N_9488,N_5379,N_7234);
xnor U9489 (N_9489,N_6344,N_6412);
nor U9490 (N_9490,N_6481,N_5583);
nor U9491 (N_9491,N_6824,N_5678);
nand U9492 (N_9492,N_6824,N_5087);
nand U9493 (N_9493,N_5951,N_6009);
or U9494 (N_9494,N_7269,N_7447);
or U9495 (N_9495,N_6819,N_5860);
and U9496 (N_9496,N_6544,N_7028);
and U9497 (N_9497,N_6500,N_5086);
and U9498 (N_9498,N_6562,N_7147);
xnor U9499 (N_9499,N_5546,N_5076);
nand U9500 (N_9500,N_6760,N_5358);
xnor U9501 (N_9501,N_5339,N_6557);
or U9502 (N_9502,N_7377,N_5169);
nor U9503 (N_9503,N_5039,N_7042);
and U9504 (N_9504,N_7422,N_6560);
nor U9505 (N_9505,N_7186,N_5662);
nand U9506 (N_9506,N_7165,N_6320);
or U9507 (N_9507,N_5832,N_6026);
nor U9508 (N_9508,N_5925,N_6490);
nand U9509 (N_9509,N_6767,N_5760);
nand U9510 (N_9510,N_7363,N_6753);
nor U9511 (N_9511,N_5449,N_5282);
xor U9512 (N_9512,N_5529,N_5286);
or U9513 (N_9513,N_6109,N_6037);
or U9514 (N_9514,N_6524,N_6584);
and U9515 (N_9515,N_7093,N_6454);
nand U9516 (N_9516,N_6364,N_7498);
nor U9517 (N_9517,N_6598,N_7377);
nor U9518 (N_9518,N_6478,N_6261);
or U9519 (N_9519,N_7176,N_5144);
nor U9520 (N_9520,N_6245,N_7202);
nand U9521 (N_9521,N_6266,N_6695);
or U9522 (N_9522,N_6817,N_7343);
and U9523 (N_9523,N_5250,N_5207);
nor U9524 (N_9524,N_7198,N_5048);
or U9525 (N_9525,N_6562,N_6612);
nand U9526 (N_9526,N_6891,N_5790);
or U9527 (N_9527,N_5979,N_7365);
and U9528 (N_9528,N_5775,N_5876);
nor U9529 (N_9529,N_5300,N_5087);
nor U9530 (N_9530,N_5684,N_6710);
xnor U9531 (N_9531,N_6354,N_5716);
or U9532 (N_9532,N_5275,N_5982);
or U9533 (N_9533,N_5596,N_5300);
or U9534 (N_9534,N_5184,N_7347);
nor U9535 (N_9535,N_6994,N_5711);
nor U9536 (N_9536,N_5120,N_6671);
or U9537 (N_9537,N_5956,N_5362);
and U9538 (N_9538,N_6395,N_5479);
and U9539 (N_9539,N_5046,N_6572);
and U9540 (N_9540,N_6516,N_6022);
or U9541 (N_9541,N_6134,N_6834);
nand U9542 (N_9542,N_6322,N_5723);
or U9543 (N_9543,N_5992,N_7321);
nor U9544 (N_9544,N_5084,N_5277);
and U9545 (N_9545,N_6237,N_5167);
or U9546 (N_9546,N_6691,N_6510);
or U9547 (N_9547,N_6244,N_5988);
or U9548 (N_9548,N_6187,N_5265);
or U9549 (N_9549,N_5935,N_5536);
nor U9550 (N_9550,N_6555,N_6944);
nor U9551 (N_9551,N_5662,N_6683);
and U9552 (N_9552,N_5594,N_5900);
and U9553 (N_9553,N_7078,N_7194);
nand U9554 (N_9554,N_6885,N_5118);
and U9555 (N_9555,N_5992,N_6304);
and U9556 (N_9556,N_5082,N_6969);
nand U9557 (N_9557,N_6893,N_5028);
or U9558 (N_9558,N_5133,N_5354);
nand U9559 (N_9559,N_7418,N_6261);
or U9560 (N_9560,N_5713,N_6278);
and U9561 (N_9561,N_6512,N_6170);
and U9562 (N_9562,N_6505,N_6425);
nand U9563 (N_9563,N_7156,N_7422);
and U9564 (N_9564,N_7469,N_7042);
nand U9565 (N_9565,N_7314,N_5773);
nand U9566 (N_9566,N_6919,N_6022);
and U9567 (N_9567,N_5117,N_5333);
and U9568 (N_9568,N_6141,N_6409);
nand U9569 (N_9569,N_5557,N_5783);
or U9570 (N_9570,N_6431,N_6150);
or U9571 (N_9571,N_7319,N_6111);
nor U9572 (N_9572,N_7373,N_6270);
and U9573 (N_9573,N_6674,N_5419);
xnor U9574 (N_9574,N_5096,N_7447);
or U9575 (N_9575,N_6584,N_5277);
nor U9576 (N_9576,N_6110,N_7253);
or U9577 (N_9577,N_7313,N_7056);
nand U9578 (N_9578,N_6045,N_6378);
or U9579 (N_9579,N_6080,N_7409);
and U9580 (N_9580,N_5250,N_7365);
and U9581 (N_9581,N_5273,N_7206);
or U9582 (N_9582,N_6703,N_5333);
or U9583 (N_9583,N_6734,N_5677);
xnor U9584 (N_9584,N_5924,N_6286);
nor U9585 (N_9585,N_5060,N_7125);
or U9586 (N_9586,N_6471,N_6843);
and U9587 (N_9587,N_5025,N_6133);
or U9588 (N_9588,N_7485,N_7141);
and U9589 (N_9589,N_7309,N_5907);
nand U9590 (N_9590,N_6547,N_6662);
nand U9591 (N_9591,N_6520,N_6663);
and U9592 (N_9592,N_5189,N_6071);
nand U9593 (N_9593,N_5247,N_6076);
and U9594 (N_9594,N_5246,N_6367);
nand U9595 (N_9595,N_6270,N_6631);
xor U9596 (N_9596,N_5711,N_6928);
nand U9597 (N_9597,N_5534,N_6166);
and U9598 (N_9598,N_6633,N_7086);
or U9599 (N_9599,N_6961,N_7349);
nand U9600 (N_9600,N_6542,N_7365);
or U9601 (N_9601,N_6895,N_7025);
and U9602 (N_9602,N_6487,N_5672);
nor U9603 (N_9603,N_6390,N_7340);
and U9604 (N_9604,N_5276,N_5223);
and U9605 (N_9605,N_6567,N_6867);
nor U9606 (N_9606,N_5257,N_6791);
nor U9607 (N_9607,N_5063,N_5704);
xor U9608 (N_9608,N_6845,N_5716);
nand U9609 (N_9609,N_5079,N_5542);
or U9610 (N_9610,N_5162,N_6240);
or U9611 (N_9611,N_6905,N_5295);
and U9612 (N_9612,N_7060,N_5917);
nor U9613 (N_9613,N_6647,N_6087);
and U9614 (N_9614,N_5859,N_7228);
nand U9615 (N_9615,N_6368,N_5680);
nand U9616 (N_9616,N_7115,N_6178);
and U9617 (N_9617,N_5402,N_5604);
nand U9618 (N_9618,N_6602,N_6503);
nand U9619 (N_9619,N_6863,N_5591);
xnor U9620 (N_9620,N_6228,N_6441);
nor U9621 (N_9621,N_7286,N_5438);
nand U9622 (N_9622,N_5366,N_6583);
nand U9623 (N_9623,N_5527,N_6384);
and U9624 (N_9624,N_5966,N_7181);
nand U9625 (N_9625,N_5505,N_7246);
nand U9626 (N_9626,N_5230,N_6856);
or U9627 (N_9627,N_6471,N_6052);
or U9628 (N_9628,N_6042,N_5526);
nand U9629 (N_9629,N_7098,N_6215);
nand U9630 (N_9630,N_7002,N_6355);
or U9631 (N_9631,N_6445,N_6352);
xor U9632 (N_9632,N_6901,N_6167);
and U9633 (N_9633,N_7471,N_7130);
or U9634 (N_9634,N_6480,N_5140);
nor U9635 (N_9635,N_6602,N_5183);
nor U9636 (N_9636,N_5301,N_5002);
nor U9637 (N_9637,N_6452,N_5290);
nor U9638 (N_9638,N_5711,N_5954);
nand U9639 (N_9639,N_6431,N_6678);
nand U9640 (N_9640,N_6675,N_6737);
nand U9641 (N_9641,N_5487,N_6861);
or U9642 (N_9642,N_6794,N_5669);
nand U9643 (N_9643,N_6839,N_6694);
nand U9644 (N_9644,N_6709,N_6568);
or U9645 (N_9645,N_6682,N_6201);
nand U9646 (N_9646,N_5573,N_6545);
xor U9647 (N_9647,N_5887,N_7241);
and U9648 (N_9648,N_6866,N_5569);
nand U9649 (N_9649,N_5577,N_7149);
nand U9650 (N_9650,N_6804,N_6315);
nand U9651 (N_9651,N_6407,N_5370);
nand U9652 (N_9652,N_5445,N_6502);
nand U9653 (N_9653,N_6631,N_5017);
and U9654 (N_9654,N_6053,N_5290);
nand U9655 (N_9655,N_5756,N_7330);
nor U9656 (N_9656,N_7176,N_5338);
and U9657 (N_9657,N_6170,N_5002);
or U9658 (N_9658,N_6496,N_6053);
nand U9659 (N_9659,N_5187,N_6182);
nand U9660 (N_9660,N_5204,N_5668);
or U9661 (N_9661,N_6569,N_5956);
and U9662 (N_9662,N_5292,N_7229);
or U9663 (N_9663,N_5283,N_6593);
nand U9664 (N_9664,N_7149,N_6498);
and U9665 (N_9665,N_5449,N_5522);
or U9666 (N_9666,N_5835,N_5014);
or U9667 (N_9667,N_7273,N_5798);
and U9668 (N_9668,N_6136,N_6082);
nor U9669 (N_9669,N_5313,N_5582);
nand U9670 (N_9670,N_6580,N_5383);
and U9671 (N_9671,N_6867,N_5779);
nand U9672 (N_9672,N_5133,N_6424);
and U9673 (N_9673,N_7052,N_6984);
nor U9674 (N_9674,N_6332,N_5770);
and U9675 (N_9675,N_5895,N_6522);
nor U9676 (N_9676,N_5066,N_6461);
nand U9677 (N_9677,N_6972,N_6656);
and U9678 (N_9678,N_6378,N_5334);
or U9679 (N_9679,N_6271,N_7378);
nor U9680 (N_9680,N_5548,N_6525);
nand U9681 (N_9681,N_5731,N_6914);
nor U9682 (N_9682,N_6326,N_6372);
nor U9683 (N_9683,N_6584,N_7386);
nand U9684 (N_9684,N_6552,N_5395);
and U9685 (N_9685,N_5460,N_6531);
and U9686 (N_9686,N_7127,N_5268);
nor U9687 (N_9687,N_6618,N_6876);
nand U9688 (N_9688,N_5308,N_6148);
or U9689 (N_9689,N_6540,N_7119);
nor U9690 (N_9690,N_5033,N_5373);
nand U9691 (N_9691,N_7454,N_6938);
nand U9692 (N_9692,N_6644,N_5255);
and U9693 (N_9693,N_6186,N_5707);
nor U9694 (N_9694,N_5647,N_6656);
nand U9695 (N_9695,N_6508,N_6226);
and U9696 (N_9696,N_5492,N_5493);
nand U9697 (N_9697,N_5136,N_5013);
and U9698 (N_9698,N_6969,N_6876);
xnor U9699 (N_9699,N_5389,N_7140);
and U9700 (N_9700,N_7303,N_7266);
or U9701 (N_9701,N_7332,N_6476);
or U9702 (N_9702,N_5945,N_6215);
nor U9703 (N_9703,N_6993,N_6614);
nor U9704 (N_9704,N_6244,N_5889);
and U9705 (N_9705,N_6684,N_6606);
nand U9706 (N_9706,N_6231,N_6132);
xnor U9707 (N_9707,N_6402,N_6020);
nand U9708 (N_9708,N_5484,N_7398);
and U9709 (N_9709,N_5318,N_6389);
xor U9710 (N_9710,N_6805,N_6210);
nand U9711 (N_9711,N_5477,N_6259);
nand U9712 (N_9712,N_6024,N_6529);
or U9713 (N_9713,N_5770,N_5460);
nand U9714 (N_9714,N_7458,N_5200);
nand U9715 (N_9715,N_5601,N_5934);
nand U9716 (N_9716,N_5668,N_5771);
nand U9717 (N_9717,N_5885,N_5816);
and U9718 (N_9718,N_6580,N_5940);
nor U9719 (N_9719,N_7330,N_6953);
nor U9720 (N_9720,N_5044,N_7468);
nor U9721 (N_9721,N_5419,N_6940);
nor U9722 (N_9722,N_5942,N_7342);
nor U9723 (N_9723,N_6187,N_7329);
nor U9724 (N_9724,N_7115,N_6865);
and U9725 (N_9725,N_5600,N_7257);
nor U9726 (N_9726,N_6842,N_7353);
nand U9727 (N_9727,N_6648,N_5608);
nand U9728 (N_9728,N_6117,N_7163);
nor U9729 (N_9729,N_6448,N_5475);
and U9730 (N_9730,N_6571,N_5528);
or U9731 (N_9731,N_5341,N_6520);
nand U9732 (N_9732,N_6239,N_7102);
or U9733 (N_9733,N_7364,N_5851);
xor U9734 (N_9734,N_7259,N_5590);
and U9735 (N_9735,N_5410,N_5820);
nor U9736 (N_9736,N_5497,N_7249);
nand U9737 (N_9737,N_7437,N_6554);
or U9738 (N_9738,N_5336,N_5023);
and U9739 (N_9739,N_7341,N_5722);
and U9740 (N_9740,N_5030,N_6457);
nor U9741 (N_9741,N_6228,N_5654);
nand U9742 (N_9742,N_5039,N_5877);
nor U9743 (N_9743,N_6539,N_6226);
and U9744 (N_9744,N_5231,N_6103);
nor U9745 (N_9745,N_6485,N_6351);
nand U9746 (N_9746,N_5410,N_6800);
nor U9747 (N_9747,N_7085,N_6621);
and U9748 (N_9748,N_7021,N_6669);
nor U9749 (N_9749,N_5297,N_5638);
nor U9750 (N_9750,N_6378,N_6882);
or U9751 (N_9751,N_7281,N_5210);
nand U9752 (N_9752,N_6638,N_5690);
or U9753 (N_9753,N_5697,N_5720);
nand U9754 (N_9754,N_6918,N_7486);
nand U9755 (N_9755,N_6747,N_6097);
nor U9756 (N_9756,N_5193,N_5425);
or U9757 (N_9757,N_6321,N_6066);
or U9758 (N_9758,N_6546,N_6007);
nor U9759 (N_9759,N_5220,N_6152);
or U9760 (N_9760,N_5237,N_5774);
and U9761 (N_9761,N_6905,N_5233);
nor U9762 (N_9762,N_6289,N_5160);
nor U9763 (N_9763,N_5902,N_5735);
nor U9764 (N_9764,N_6955,N_7346);
nor U9765 (N_9765,N_5890,N_5571);
and U9766 (N_9766,N_6547,N_5259);
nor U9767 (N_9767,N_5401,N_6395);
nand U9768 (N_9768,N_7396,N_6344);
or U9769 (N_9769,N_7169,N_7144);
nor U9770 (N_9770,N_6208,N_6270);
nand U9771 (N_9771,N_6370,N_5589);
nor U9772 (N_9772,N_7154,N_7391);
nor U9773 (N_9773,N_6996,N_6976);
and U9774 (N_9774,N_5010,N_5690);
nor U9775 (N_9775,N_5289,N_5774);
and U9776 (N_9776,N_5256,N_6291);
nor U9777 (N_9777,N_5698,N_7190);
nand U9778 (N_9778,N_6040,N_6820);
nor U9779 (N_9779,N_7062,N_5480);
or U9780 (N_9780,N_6793,N_6110);
nor U9781 (N_9781,N_5773,N_6878);
nor U9782 (N_9782,N_5108,N_7163);
nand U9783 (N_9783,N_6413,N_7175);
or U9784 (N_9784,N_6553,N_6632);
nor U9785 (N_9785,N_6279,N_7246);
nand U9786 (N_9786,N_5582,N_6483);
or U9787 (N_9787,N_5442,N_5322);
and U9788 (N_9788,N_5558,N_5789);
and U9789 (N_9789,N_5613,N_6481);
nand U9790 (N_9790,N_5649,N_5634);
nor U9791 (N_9791,N_5411,N_6397);
nor U9792 (N_9792,N_5411,N_7096);
nand U9793 (N_9793,N_7431,N_6946);
nand U9794 (N_9794,N_7475,N_5190);
nor U9795 (N_9795,N_5879,N_6169);
or U9796 (N_9796,N_5053,N_7374);
xnor U9797 (N_9797,N_7413,N_5023);
or U9798 (N_9798,N_6404,N_5510);
and U9799 (N_9799,N_7034,N_6295);
and U9800 (N_9800,N_7080,N_7276);
and U9801 (N_9801,N_7167,N_5727);
nand U9802 (N_9802,N_6480,N_5117);
nor U9803 (N_9803,N_7270,N_5146);
and U9804 (N_9804,N_5429,N_6817);
or U9805 (N_9805,N_5716,N_6757);
nand U9806 (N_9806,N_7040,N_5521);
nor U9807 (N_9807,N_5696,N_7420);
nor U9808 (N_9808,N_6431,N_5415);
nand U9809 (N_9809,N_6632,N_6167);
nand U9810 (N_9810,N_5761,N_5505);
and U9811 (N_9811,N_6721,N_7335);
or U9812 (N_9812,N_6344,N_5661);
nor U9813 (N_9813,N_6252,N_6001);
or U9814 (N_9814,N_6873,N_5508);
xnor U9815 (N_9815,N_6295,N_6737);
nand U9816 (N_9816,N_7214,N_6643);
and U9817 (N_9817,N_5311,N_5855);
nand U9818 (N_9818,N_7421,N_7074);
and U9819 (N_9819,N_7398,N_5210);
and U9820 (N_9820,N_6793,N_5323);
and U9821 (N_9821,N_6324,N_5543);
or U9822 (N_9822,N_5828,N_7025);
nor U9823 (N_9823,N_5802,N_6899);
xnor U9824 (N_9824,N_5944,N_5504);
or U9825 (N_9825,N_6423,N_6526);
and U9826 (N_9826,N_6086,N_5440);
nor U9827 (N_9827,N_5041,N_6410);
nor U9828 (N_9828,N_6690,N_5737);
nor U9829 (N_9829,N_5217,N_5771);
nand U9830 (N_9830,N_6620,N_5490);
or U9831 (N_9831,N_7031,N_6894);
or U9832 (N_9832,N_7270,N_6593);
or U9833 (N_9833,N_5074,N_6621);
or U9834 (N_9834,N_7111,N_6436);
nand U9835 (N_9835,N_6929,N_5125);
and U9836 (N_9836,N_6782,N_6231);
nand U9837 (N_9837,N_6524,N_6579);
and U9838 (N_9838,N_6183,N_5748);
and U9839 (N_9839,N_5541,N_6237);
nor U9840 (N_9840,N_6132,N_6074);
nand U9841 (N_9841,N_6090,N_6285);
nand U9842 (N_9842,N_6292,N_5560);
nor U9843 (N_9843,N_5024,N_5872);
nand U9844 (N_9844,N_6545,N_5837);
nor U9845 (N_9845,N_6639,N_6618);
nor U9846 (N_9846,N_6210,N_6697);
nor U9847 (N_9847,N_6180,N_6717);
and U9848 (N_9848,N_5620,N_6385);
or U9849 (N_9849,N_7254,N_7378);
or U9850 (N_9850,N_7003,N_7360);
nand U9851 (N_9851,N_5429,N_6619);
nor U9852 (N_9852,N_7190,N_5740);
or U9853 (N_9853,N_6971,N_5694);
and U9854 (N_9854,N_7082,N_6140);
nand U9855 (N_9855,N_6795,N_5989);
and U9856 (N_9856,N_7190,N_5573);
nor U9857 (N_9857,N_7022,N_6662);
nor U9858 (N_9858,N_5185,N_6153);
nor U9859 (N_9859,N_6098,N_5648);
or U9860 (N_9860,N_6654,N_7107);
or U9861 (N_9861,N_5719,N_6938);
xnor U9862 (N_9862,N_6866,N_7005);
and U9863 (N_9863,N_6026,N_5493);
and U9864 (N_9864,N_5593,N_6699);
xor U9865 (N_9865,N_7453,N_7159);
and U9866 (N_9866,N_7413,N_6989);
or U9867 (N_9867,N_6124,N_5969);
and U9868 (N_9868,N_6767,N_6317);
or U9869 (N_9869,N_5726,N_6517);
nand U9870 (N_9870,N_6174,N_6693);
nand U9871 (N_9871,N_6011,N_6929);
and U9872 (N_9872,N_5850,N_6589);
or U9873 (N_9873,N_6149,N_5861);
nor U9874 (N_9874,N_6685,N_5088);
and U9875 (N_9875,N_5953,N_7328);
and U9876 (N_9876,N_5925,N_7119);
xnor U9877 (N_9877,N_5007,N_5517);
and U9878 (N_9878,N_7153,N_5700);
nor U9879 (N_9879,N_5353,N_6594);
nand U9880 (N_9880,N_6866,N_7043);
and U9881 (N_9881,N_5945,N_6991);
or U9882 (N_9882,N_5521,N_6524);
or U9883 (N_9883,N_5595,N_6693);
or U9884 (N_9884,N_6202,N_7457);
and U9885 (N_9885,N_5780,N_5180);
nor U9886 (N_9886,N_5232,N_5886);
nand U9887 (N_9887,N_6334,N_6615);
nand U9888 (N_9888,N_6409,N_7153);
and U9889 (N_9889,N_7305,N_6803);
nor U9890 (N_9890,N_6290,N_7329);
or U9891 (N_9891,N_5392,N_6244);
and U9892 (N_9892,N_6193,N_5475);
and U9893 (N_9893,N_5648,N_7445);
nor U9894 (N_9894,N_5375,N_6121);
and U9895 (N_9895,N_6522,N_7302);
nand U9896 (N_9896,N_6970,N_6557);
nand U9897 (N_9897,N_7120,N_5917);
nor U9898 (N_9898,N_7120,N_6304);
nand U9899 (N_9899,N_6202,N_6526);
or U9900 (N_9900,N_5237,N_5150);
or U9901 (N_9901,N_5208,N_5091);
nand U9902 (N_9902,N_5533,N_5727);
or U9903 (N_9903,N_6186,N_7467);
xnor U9904 (N_9904,N_7254,N_5789);
nand U9905 (N_9905,N_6739,N_5175);
nand U9906 (N_9906,N_6859,N_5178);
and U9907 (N_9907,N_5104,N_7333);
or U9908 (N_9908,N_6599,N_5568);
or U9909 (N_9909,N_5942,N_5098);
or U9910 (N_9910,N_5206,N_7083);
nor U9911 (N_9911,N_5718,N_6334);
or U9912 (N_9912,N_7302,N_5323);
nand U9913 (N_9913,N_7271,N_7215);
nor U9914 (N_9914,N_6939,N_6693);
nand U9915 (N_9915,N_6308,N_6828);
nor U9916 (N_9916,N_6284,N_6635);
xor U9917 (N_9917,N_6889,N_6871);
or U9918 (N_9918,N_5728,N_5967);
and U9919 (N_9919,N_6462,N_6376);
nand U9920 (N_9920,N_5897,N_6712);
nand U9921 (N_9921,N_6698,N_6169);
or U9922 (N_9922,N_5239,N_5764);
or U9923 (N_9923,N_5100,N_6594);
nor U9924 (N_9924,N_5210,N_6571);
nor U9925 (N_9925,N_5076,N_5911);
and U9926 (N_9926,N_7187,N_5691);
nand U9927 (N_9927,N_6138,N_5493);
or U9928 (N_9928,N_5747,N_5388);
nand U9929 (N_9929,N_5621,N_5033);
nor U9930 (N_9930,N_5164,N_6778);
or U9931 (N_9931,N_5401,N_6579);
and U9932 (N_9932,N_7141,N_6591);
nand U9933 (N_9933,N_7148,N_6266);
and U9934 (N_9934,N_5972,N_5497);
and U9935 (N_9935,N_5024,N_7087);
nand U9936 (N_9936,N_6767,N_5651);
nand U9937 (N_9937,N_6000,N_5106);
nand U9938 (N_9938,N_7158,N_5381);
nand U9939 (N_9939,N_5472,N_5567);
nor U9940 (N_9940,N_5459,N_7014);
or U9941 (N_9941,N_5861,N_6108);
nor U9942 (N_9942,N_6094,N_7243);
nand U9943 (N_9943,N_5948,N_5155);
nand U9944 (N_9944,N_7183,N_7120);
nor U9945 (N_9945,N_5055,N_6830);
nand U9946 (N_9946,N_6842,N_5627);
nand U9947 (N_9947,N_6984,N_7371);
or U9948 (N_9948,N_6257,N_5455);
nor U9949 (N_9949,N_5678,N_7482);
or U9950 (N_9950,N_7254,N_6599);
nor U9951 (N_9951,N_6607,N_5338);
or U9952 (N_9952,N_7271,N_5054);
and U9953 (N_9953,N_5380,N_5265);
nand U9954 (N_9954,N_5626,N_6210);
and U9955 (N_9955,N_7178,N_6876);
nand U9956 (N_9956,N_7286,N_7029);
nand U9957 (N_9957,N_5630,N_5349);
or U9958 (N_9958,N_5635,N_5727);
nor U9959 (N_9959,N_5537,N_5448);
nand U9960 (N_9960,N_7226,N_5698);
nor U9961 (N_9961,N_7350,N_6138);
or U9962 (N_9962,N_5383,N_6144);
nor U9963 (N_9963,N_5680,N_7350);
and U9964 (N_9964,N_7299,N_5701);
nand U9965 (N_9965,N_6314,N_6247);
nor U9966 (N_9966,N_5501,N_6150);
xnor U9967 (N_9967,N_5591,N_7193);
and U9968 (N_9968,N_6883,N_7252);
nand U9969 (N_9969,N_7025,N_5345);
nand U9970 (N_9970,N_6264,N_6055);
nor U9971 (N_9971,N_6397,N_6822);
or U9972 (N_9972,N_5592,N_5594);
and U9973 (N_9973,N_5315,N_6747);
or U9974 (N_9974,N_6652,N_6973);
nor U9975 (N_9975,N_5965,N_6463);
and U9976 (N_9976,N_5285,N_5943);
or U9977 (N_9977,N_6676,N_5612);
xnor U9978 (N_9978,N_6088,N_6992);
nor U9979 (N_9979,N_6465,N_6733);
nor U9980 (N_9980,N_5605,N_5582);
or U9981 (N_9981,N_5325,N_7439);
nor U9982 (N_9982,N_6647,N_5487);
or U9983 (N_9983,N_5502,N_6790);
nand U9984 (N_9984,N_6599,N_5937);
and U9985 (N_9985,N_6533,N_5823);
or U9986 (N_9986,N_5527,N_6954);
nand U9987 (N_9987,N_7449,N_6413);
nand U9988 (N_9988,N_6768,N_7008);
nand U9989 (N_9989,N_5535,N_6558);
or U9990 (N_9990,N_5858,N_6753);
and U9991 (N_9991,N_5129,N_5808);
nand U9992 (N_9992,N_5062,N_7179);
or U9993 (N_9993,N_6118,N_6316);
nand U9994 (N_9994,N_7288,N_6940);
or U9995 (N_9995,N_6133,N_7410);
nor U9996 (N_9996,N_7122,N_7487);
or U9997 (N_9997,N_5056,N_6592);
and U9998 (N_9998,N_7058,N_5724);
and U9999 (N_9999,N_5997,N_5231);
nor UO_0 (O_0,N_8995,N_7786);
and UO_1 (O_1,N_8923,N_8239);
and UO_2 (O_2,N_9777,N_9944);
and UO_3 (O_3,N_8513,N_9984);
nor UO_4 (O_4,N_8050,N_9327);
and UO_5 (O_5,N_9381,N_9189);
nand UO_6 (O_6,N_9823,N_8293);
nand UO_7 (O_7,N_8784,N_9828);
nand UO_8 (O_8,N_8730,N_8336);
and UO_9 (O_9,N_8181,N_9998);
nor UO_10 (O_10,N_9871,N_9743);
and UO_11 (O_11,N_7754,N_8176);
nor UO_12 (O_12,N_7915,N_8347);
nand UO_13 (O_13,N_9168,N_9304);
or UO_14 (O_14,N_8426,N_9046);
nor UO_15 (O_15,N_9987,N_8165);
nor UO_16 (O_16,N_9230,N_7942);
or UO_17 (O_17,N_8779,N_9044);
xor UO_18 (O_18,N_9425,N_8331);
or UO_19 (O_19,N_7838,N_8467);
nand UO_20 (O_20,N_9771,N_9147);
nor UO_21 (O_21,N_8414,N_9899);
nor UO_22 (O_22,N_8459,N_9047);
or UO_23 (O_23,N_7825,N_8968);
nand UO_24 (O_24,N_9224,N_8522);
nand UO_25 (O_25,N_7662,N_9036);
or UO_26 (O_26,N_7553,N_9174);
nor UO_27 (O_27,N_7758,N_8411);
nand UO_28 (O_28,N_9589,N_8096);
and UO_29 (O_29,N_8281,N_7990);
and UO_30 (O_30,N_9506,N_7850);
and UO_31 (O_31,N_8958,N_9467);
nor UO_32 (O_32,N_9225,N_8728);
nand UO_33 (O_33,N_9878,N_8041);
nand UO_34 (O_34,N_8270,N_8847);
and UO_35 (O_35,N_7775,N_8277);
and UO_36 (O_36,N_8353,N_9517);
nand UO_37 (O_37,N_8228,N_9384);
nor UO_38 (O_38,N_8882,N_7853);
and UO_39 (O_39,N_9336,N_8648);
nor UO_40 (O_40,N_9027,N_9917);
nor UO_41 (O_41,N_7813,N_8564);
and UO_42 (O_42,N_9612,N_9827);
or UO_43 (O_43,N_8567,N_8764);
and UO_44 (O_44,N_9710,N_8514);
or UO_45 (O_45,N_9145,N_8042);
or UO_46 (O_46,N_7847,N_8694);
or UO_47 (O_47,N_7628,N_8590);
or UO_48 (O_48,N_7556,N_7968);
nand UO_49 (O_49,N_9974,N_8273);
and UO_50 (O_50,N_9958,N_9964);
nand UO_51 (O_51,N_8319,N_9433);
nand UO_52 (O_52,N_7760,N_8120);
xnor UO_53 (O_53,N_8868,N_8424);
and UO_54 (O_54,N_8404,N_7576);
or UO_55 (O_55,N_7660,N_8260);
or UO_56 (O_56,N_7964,N_7987);
and UO_57 (O_57,N_8951,N_8945);
nor UO_58 (O_58,N_8295,N_9696);
and UO_59 (O_59,N_9086,N_9947);
and UO_60 (O_60,N_9200,N_7574);
nor UO_61 (O_61,N_8160,N_8828);
nand UO_62 (O_62,N_8544,N_9795);
nand UO_63 (O_63,N_9724,N_7588);
nor UO_64 (O_64,N_9244,N_8027);
nor UO_65 (O_65,N_8210,N_8299);
nor UO_66 (O_66,N_8431,N_8103);
nand UO_67 (O_67,N_9892,N_8225);
nand UO_68 (O_68,N_7560,N_9955);
nand UO_69 (O_69,N_8139,N_9687);
or UO_70 (O_70,N_8509,N_8778);
and UO_71 (O_71,N_9383,N_9308);
or UO_72 (O_72,N_8562,N_9848);
nor UO_73 (O_73,N_8623,N_9786);
nand UO_74 (O_74,N_7674,N_7913);
xnor UO_75 (O_75,N_7642,N_9034);
nor UO_76 (O_76,N_8141,N_9029);
and UO_77 (O_77,N_8804,N_8048);
or UO_78 (O_78,N_9177,N_9317);
nor UO_79 (O_79,N_9246,N_8019);
or UO_80 (O_80,N_7746,N_8841);
and UO_81 (O_81,N_9785,N_9581);
and UO_82 (O_82,N_9202,N_8724);
or UO_83 (O_83,N_8300,N_8925);
nand UO_84 (O_84,N_8512,N_8002);
or UO_85 (O_85,N_8954,N_7870);
nand UO_86 (O_86,N_9812,N_7601);
or UO_87 (O_87,N_9717,N_9411);
or UO_88 (O_88,N_7637,N_8960);
nor UO_89 (O_89,N_8856,N_9942);
or UO_90 (O_90,N_9709,N_9925);
or UO_91 (O_91,N_8739,N_9928);
or UO_92 (O_92,N_7720,N_9948);
or UO_93 (O_93,N_9720,N_9111);
and UO_94 (O_94,N_8261,N_8116);
nand UO_95 (O_95,N_9302,N_9500);
and UO_96 (O_96,N_9719,N_9161);
nand UO_97 (O_97,N_9443,N_9166);
or UO_98 (O_98,N_9770,N_8162);
nor UO_99 (O_99,N_9836,N_7879);
or UO_100 (O_100,N_8574,N_8114);
and UO_101 (O_101,N_9496,N_9728);
and UO_102 (O_102,N_9756,N_8851);
nor UO_103 (O_103,N_8859,N_7741);
nand UO_104 (O_104,N_8576,N_9560);
nor UO_105 (O_105,N_8021,N_9755);
or UO_106 (O_106,N_8504,N_9085);
nand UO_107 (O_107,N_9653,N_8583);
or UO_108 (O_108,N_8036,N_8057);
nor UO_109 (O_109,N_7757,N_8146);
nand UO_110 (O_110,N_8571,N_8267);
and UO_111 (O_111,N_8642,N_9761);
or UO_112 (O_112,N_8731,N_7520);
nand UO_113 (O_113,N_7785,N_8364);
and UO_114 (O_114,N_7876,N_9254);
and UO_115 (O_115,N_8090,N_7614);
and UO_116 (O_116,N_8494,N_8844);
nand UO_117 (O_117,N_8624,N_7695);
or UO_118 (O_118,N_8896,N_7510);
or UO_119 (O_119,N_8385,N_8199);
and UO_120 (O_120,N_9454,N_8020);
or UO_121 (O_121,N_8689,N_8743);
and UO_122 (O_122,N_8713,N_9397);
or UO_123 (O_123,N_9193,N_9949);
or UO_124 (O_124,N_7536,N_9704);
xnor UO_125 (O_125,N_9956,N_9543);
nand UO_126 (O_126,N_9257,N_9701);
and UO_127 (O_127,N_8285,N_7833);
nand UO_128 (O_128,N_9576,N_9766);
and UO_129 (O_129,N_7708,N_8810);
nor UO_130 (O_130,N_8985,N_9686);
nor UO_131 (O_131,N_8323,N_9595);
nor UO_132 (O_132,N_7690,N_7533);
or UO_133 (O_133,N_9982,N_7511);
or UO_134 (O_134,N_9850,N_9160);
nor UO_135 (O_135,N_7594,N_9556);
and UO_136 (O_136,N_9866,N_9421);
and UO_137 (O_137,N_9416,N_9076);
nand UO_138 (O_138,N_7527,N_8388);
and UO_139 (O_139,N_9460,N_7515);
and UO_140 (O_140,N_8678,N_9475);
nor UO_141 (O_141,N_9860,N_7592);
or UO_142 (O_142,N_8102,N_7729);
and UO_143 (O_143,N_8733,N_9830);
nor UO_144 (O_144,N_8455,N_8534);
and UO_145 (O_145,N_7989,N_8537);
nor UO_146 (O_146,N_9452,N_8524);
nand UO_147 (O_147,N_9937,N_8366);
or UO_148 (O_148,N_9343,N_9342);
or UO_149 (O_149,N_8831,N_8227);
and UO_150 (O_150,N_7514,N_9374);
and UO_151 (O_151,N_8203,N_7617);
nor UO_152 (O_152,N_9057,N_8776);
nor UO_153 (O_153,N_9398,N_8445);
nor UO_154 (O_154,N_8437,N_7716);
xnor UO_155 (O_155,N_8486,N_9285);
nand UO_156 (O_156,N_8344,N_8127);
nor UO_157 (O_157,N_9075,N_8992);
nor UO_158 (O_158,N_8461,N_7559);
nand UO_159 (O_159,N_7792,N_8064);
and UO_160 (O_160,N_8205,N_9021);
and UO_161 (O_161,N_8518,N_9705);
nor UO_162 (O_162,N_9572,N_9468);
nor UO_163 (O_163,N_9915,N_7562);
or UO_164 (O_164,N_7540,N_7569);
or UO_165 (O_165,N_9172,N_8785);
or UO_166 (O_166,N_7784,N_7701);
and UO_167 (O_167,N_9370,N_8664);
nand UO_168 (O_168,N_7797,N_9056);
nor UO_169 (O_169,N_9877,N_9862);
nand UO_170 (O_170,N_9415,N_7826);
nand UO_171 (O_171,N_8348,N_8044);
nor UO_172 (O_172,N_8091,N_8873);
nor UO_173 (O_173,N_9791,N_9000);
nand UO_174 (O_174,N_9992,N_7781);
nor UO_175 (O_175,N_8558,N_7806);
and UO_176 (O_176,N_8125,N_9681);
and UO_177 (O_177,N_9391,N_9657);
nor UO_178 (O_178,N_8809,N_9497);
or UO_179 (O_179,N_9676,N_8378);
or UO_180 (O_180,N_9980,N_9015);
nand UO_181 (O_181,N_9215,N_8993);
nor UO_182 (O_182,N_8183,N_7904);
or UO_183 (O_183,N_7609,N_9447);
and UO_184 (O_184,N_9604,N_8208);
or UO_185 (O_185,N_8994,N_9226);
or UO_186 (O_186,N_8981,N_9249);
nand UO_187 (O_187,N_7945,N_8812);
or UO_188 (O_188,N_9074,N_9292);
and UO_189 (O_189,N_8088,N_9555);
and UO_190 (O_190,N_9377,N_8974);
nor UO_191 (O_191,N_9598,N_7507);
and UO_192 (O_192,N_9584,N_7868);
nand UO_193 (O_193,N_9049,N_8175);
nor UO_194 (O_194,N_7591,N_7763);
and UO_195 (O_195,N_7564,N_8098);
nor UO_196 (O_196,N_8858,N_8843);
or UO_197 (O_197,N_8238,N_7636);
and UO_198 (O_198,N_7842,N_9819);
and UO_199 (O_199,N_8072,N_8454);
or UO_200 (O_200,N_8618,N_9300);
or UO_201 (O_201,N_8189,N_8074);
or UO_202 (O_202,N_8516,N_8961);
or UO_203 (O_203,N_8909,N_7856);
and UO_204 (O_204,N_9176,N_9538);
or UO_205 (O_205,N_8190,N_9624);
nor UO_206 (O_206,N_8458,N_7871);
nor UO_207 (O_207,N_8085,N_9644);
and UO_208 (O_208,N_8649,N_8555);
nand UO_209 (O_209,N_8005,N_8258);
and UO_210 (O_210,N_9312,N_7956);
or UO_211 (O_211,N_8839,N_8794);
and UO_212 (O_212,N_7726,N_9339);
and UO_213 (O_213,N_8172,N_9376);
and UO_214 (O_214,N_8708,N_9059);
nor UO_215 (O_215,N_8895,N_7638);
nand UO_216 (O_216,N_9675,N_8886);
and UO_217 (O_217,N_9325,N_9641);
nor UO_218 (O_218,N_8263,N_8322);
nor UO_219 (O_219,N_8440,N_7656);
nand UO_220 (O_220,N_8766,N_7652);
or UO_221 (O_221,N_8406,N_9531);
and UO_222 (O_222,N_8602,N_7770);
nand UO_223 (O_223,N_8241,N_9006);
nor UO_224 (O_224,N_9872,N_8410);
nor UO_225 (O_225,N_9549,N_7725);
and UO_226 (O_226,N_8750,N_9801);
nor UO_227 (O_227,N_8919,N_8453);
and UO_228 (O_228,N_7975,N_8640);
and UO_229 (O_229,N_8680,N_7789);
nand UO_230 (O_230,N_7903,N_9981);
nand UO_231 (O_231,N_8675,N_8326);
nor UO_232 (O_232,N_7762,N_9155);
and UO_233 (O_233,N_8852,N_7571);
nand UO_234 (O_234,N_8656,N_7737);
nor UO_235 (O_235,N_9236,N_8927);
nor UO_236 (O_236,N_9119,N_7764);
nand UO_237 (O_237,N_8177,N_9600);
nand UO_238 (O_238,N_8421,N_8620);
or UO_239 (O_239,N_9678,N_8673);
nand UO_240 (O_240,N_7509,N_9844);
and UO_241 (O_241,N_9185,N_9393);
nor UO_242 (O_242,N_9286,N_8483);
nand UO_243 (O_243,N_8413,N_9586);
and UO_244 (O_244,N_9101,N_9267);
nor UO_245 (O_245,N_9229,N_8290);
nor UO_246 (O_246,N_8752,N_8798);
and UO_247 (O_247,N_9703,N_9472);
nand UO_248 (O_248,N_7889,N_9727);
nand UO_249 (O_249,N_8755,N_9404);
or UO_250 (O_250,N_9627,N_9431);
and UO_251 (O_251,N_8032,N_9718);
and UO_252 (O_252,N_8737,N_9638);
nor UO_253 (O_253,N_7552,N_8899);
nand UO_254 (O_254,N_7530,N_7654);
nor UO_255 (O_255,N_8906,N_7772);
xnor UO_256 (O_256,N_9395,N_7687);
or UO_257 (O_257,N_8200,N_9889);
nand UO_258 (O_258,N_7955,N_7863);
and UO_259 (O_259,N_9401,N_9930);
nand UO_260 (O_260,N_8825,N_8612);
or UO_261 (O_261,N_9732,N_7947);
nor UO_262 (O_262,N_8606,N_9923);
and UO_263 (O_263,N_9869,N_8118);
nand UO_264 (O_264,N_7615,N_8861);
or UO_265 (O_265,N_9833,N_7901);
xnor UO_266 (O_266,N_9248,N_8706);
or UO_267 (O_267,N_9534,N_9438);
and UO_268 (O_268,N_9127,N_9941);
or UO_269 (O_269,N_9505,N_7969);
nor UO_270 (O_270,N_8670,N_9297);
or UO_271 (O_271,N_9037,N_8417);
nand UO_272 (O_272,N_9615,N_9216);
nand UO_273 (O_273,N_8119,N_8374);
nand UO_274 (O_274,N_9861,N_7860);
nor UO_275 (O_275,N_8536,N_7818);
or UO_276 (O_276,N_7765,N_9323);
and UO_277 (O_277,N_8188,N_9313);
or UO_278 (O_278,N_8449,N_8399);
and UO_279 (O_279,N_8986,N_8511);
or UO_280 (O_280,N_9977,N_9768);
nand UO_281 (O_281,N_9250,N_7517);
nand UO_282 (O_282,N_9753,N_9737);
or UO_283 (O_283,N_7547,N_8481);
and UO_284 (O_284,N_9330,N_9184);
nor UO_285 (O_285,N_9135,N_9541);
or UO_286 (O_286,N_9150,N_7886);
and UO_287 (O_287,N_8936,N_8055);
or UO_288 (O_288,N_9334,N_8529);
or UO_289 (O_289,N_8464,N_8818);
and UO_290 (O_290,N_7516,N_9252);
and UO_291 (O_291,N_8444,N_9445);
or UO_292 (O_292,N_7551,N_7704);
or UO_293 (O_293,N_9396,N_8419);
nor UO_294 (O_294,N_9986,N_8506);
nor UO_295 (O_295,N_9702,N_8206);
nand UO_296 (O_296,N_7963,N_8924);
and UO_297 (O_297,N_9060,N_9010);
nor UO_298 (O_298,N_8677,N_9769);
nor UO_299 (O_299,N_9243,N_9341);
or UO_300 (O_300,N_7976,N_8218);
and UO_301 (O_301,N_7997,N_8488);
nand UO_302 (O_302,N_9792,N_7914);
and UO_303 (O_303,N_8645,N_8835);
nor UO_304 (O_304,N_9364,N_9960);
nand UO_305 (O_305,N_7897,N_8772);
nand UO_306 (O_306,N_9389,N_9289);
nor UO_307 (O_307,N_9845,N_9832);
and UO_308 (O_308,N_9876,N_9122);
and UO_309 (O_309,N_7561,N_7633);
and UO_310 (O_310,N_9590,N_8060);
nor UO_311 (O_311,N_9750,N_8638);
and UO_312 (O_312,N_8530,N_8446);
or UO_313 (O_313,N_8546,N_7805);
and UO_314 (O_314,N_8156,N_9052);
nor UO_315 (O_315,N_8774,N_8871);
nor UO_316 (O_316,N_9841,N_9504);
or UO_317 (O_317,N_7523,N_9118);
and UO_318 (O_318,N_8807,N_9896);
or UO_319 (O_319,N_9731,N_8948);
or UO_320 (O_320,N_9146,N_9032);
or UO_321 (O_321,N_9817,N_8519);
and UO_322 (O_322,N_8163,N_8138);
nand UO_323 (O_323,N_7873,N_9684);
and UO_324 (O_324,N_9479,N_8051);
or UO_325 (O_325,N_8790,N_8617);
and UO_326 (O_326,N_7844,N_8422);
nand UO_327 (O_327,N_8997,N_9359);
or UO_328 (O_328,N_9901,N_8140);
nor UO_329 (O_329,N_8869,N_8716);
or UO_330 (O_330,N_8174,N_7621);
or UO_331 (O_331,N_7902,N_9124);
nand UO_332 (O_332,N_7965,N_9592);
or UO_333 (O_333,N_9815,N_7927);
nor UO_334 (O_334,N_8879,N_8877);
nor UO_335 (O_335,N_9091,N_9485);
or UO_336 (O_336,N_8220,N_8372);
nor UO_337 (O_337,N_9634,N_7796);
nand UO_338 (O_338,N_8226,N_8217);
and UO_339 (O_339,N_7512,N_7550);
nand UO_340 (O_340,N_8480,N_7835);
nand UO_341 (O_341,N_9978,N_7557);
and UO_342 (O_342,N_7735,N_8685);
or UO_343 (O_343,N_9256,N_9126);
or UO_344 (O_344,N_7974,N_9671);
nor UO_345 (O_345,N_9163,N_8040);
nand UO_346 (O_346,N_7728,N_9729);
nand UO_347 (O_347,N_8129,N_8984);
and UO_348 (O_348,N_9423,N_9587);
and UO_349 (O_349,N_9080,N_9407);
and UO_350 (O_350,N_8012,N_8365);
and UO_351 (O_351,N_7984,N_9322);
nand UO_352 (O_352,N_9533,N_8307);
xor UO_353 (O_353,N_7608,N_8965);
nand UO_354 (O_354,N_7727,N_8736);
or UO_355 (O_355,N_7867,N_8478);
or UO_356 (O_356,N_9898,N_8697);
nor UO_357 (O_357,N_9142,N_8988);
xor UO_358 (O_358,N_8663,N_8266);
and UO_359 (O_359,N_7898,N_8479);
or UO_360 (O_360,N_8605,N_7973);
nor UO_361 (O_361,N_7712,N_7837);
xnor UO_362 (O_362,N_9363,N_8379);
nand UO_363 (O_363,N_9561,N_8741);
nand UO_364 (O_364,N_9408,N_8709);
nand UO_365 (O_365,N_8732,N_7875);
nor UO_366 (O_366,N_9886,N_8324);
or UO_367 (O_367,N_9255,N_7679);
and UO_368 (O_368,N_8104,N_9692);
and UO_369 (O_369,N_9204,N_7791);
and UO_370 (O_370,N_7694,N_9979);
and UO_371 (O_371,N_9968,N_8133);
nor UO_372 (O_372,N_7800,N_8943);
nand UO_373 (O_373,N_7703,N_8355);
nor UO_374 (O_374,N_8161,N_9940);
nor UO_375 (O_375,N_7713,N_9270);
nor UO_376 (O_376,N_8944,N_7851);
nor UO_377 (O_377,N_9603,N_8275);
nor UO_378 (O_378,N_9430,N_7983);
nor UO_379 (O_379,N_7864,N_8117);
nor UO_380 (O_380,N_9571,N_9864);
nor UO_381 (O_381,N_9806,N_9579);
or UO_382 (O_382,N_9945,N_9347);
and UO_383 (O_383,N_8317,N_9242);
nand UO_384 (O_384,N_8823,N_8236);
and UO_385 (O_385,N_7597,N_9999);
and UO_386 (O_386,N_9477,N_7709);
nand UO_387 (O_387,N_9321,N_8942);
and UO_388 (O_388,N_8803,N_8634);
and UO_389 (O_389,N_9783,N_9706);
or UO_390 (O_390,N_9435,N_9131);
and UO_391 (O_391,N_7506,N_8552);
nor UO_392 (O_392,N_8912,N_7865);
and UO_393 (O_393,N_8628,N_8539);
nand UO_394 (O_394,N_8854,N_8933);
or UO_395 (O_395,N_8510,N_9854);
nand UO_396 (O_396,N_8598,N_9623);
or UO_397 (O_397,N_8561,N_8435);
or UO_398 (O_398,N_7528,N_9963);
and UO_399 (O_399,N_9629,N_8124);
nor UO_400 (O_400,N_9759,N_9959);
nand UO_401 (O_401,N_9662,N_9640);
nand UO_402 (O_402,N_7659,N_9690);
nand UO_403 (O_403,N_7535,N_9446);
or UO_404 (O_404,N_9482,N_9716);
nor UO_405 (O_405,N_8891,N_8863);
nand UO_406 (O_406,N_8354,N_8065);
and UO_407 (O_407,N_8073,N_7878);
nand UO_408 (O_408,N_9933,N_8375);
or UO_409 (O_409,N_8523,N_8526);
and UO_410 (O_410,N_9361,N_8097);
or UO_411 (O_411,N_8682,N_9412);
xor UO_412 (O_412,N_9069,N_8022);
nor UO_413 (O_413,N_9642,N_8830);
or UO_414 (O_414,N_8157,N_8145);
nand UO_415 (O_415,N_8672,N_8350);
nor UO_416 (O_416,N_8373,N_8765);
or UO_417 (O_417,N_8463,N_9782);
nor UO_418 (O_418,N_9156,N_8250);
nand UO_419 (O_419,N_7666,N_9680);
or UO_420 (O_420,N_8693,N_9611);
nand UO_421 (O_421,N_8262,N_8788);
and UO_422 (O_422,N_9462,N_7639);
nand UO_423 (O_423,N_9171,N_8213);
nor UO_424 (O_424,N_7620,N_7830);
and UO_425 (O_425,N_7732,N_8497);
or UO_426 (O_426,N_8184,N_9097);
or UO_427 (O_427,N_9526,N_9647);
and UO_428 (O_428,N_9668,N_9622);
nand UO_429 (O_429,N_8885,N_8007);
and UO_430 (O_430,N_9221,N_9351);
nor UO_431 (O_431,N_8930,N_7986);
and UO_432 (O_432,N_9666,N_8237);
nor UO_433 (O_433,N_9108,N_9050);
or UO_434 (O_434,N_8452,N_7584);
nand UO_435 (O_435,N_7573,N_8089);
and UO_436 (O_436,N_8609,N_9700);
or UO_437 (O_437,N_8934,N_9259);
and UO_438 (O_438,N_9673,N_8581);
or UO_439 (O_439,N_8112,N_8596);
nand UO_440 (O_440,N_8575,N_9328);
nor UO_441 (O_441,N_8989,N_8130);
and UO_442 (O_442,N_9989,N_9400);
or UO_443 (O_443,N_9318,N_9616);
nor UO_444 (O_444,N_7630,N_7959);
or UO_445 (O_445,N_8159,N_9633);
and UO_446 (O_446,N_9455,N_7750);
nand UO_447 (O_447,N_9023,N_7663);
nor UO_448 (O_448,N_7521,N_9851);
and UO_449 (O_449,N_9907,N_7738);
nand UO_450 (O_450,N_7954,N_7960);
or UO_451 (O_451,N_9188,N_9508);
nand UO_452 (O_452,N_9601,N_8178);
nand UO_453 (O_453,N_9975,N_7539);
or UO_454 (O_454,N_9966,N_9846);
or UO_455 (O_455,N_8698,N_9880);
or UO_456 (O_456,N_9664,N_7855);
nand UO_457 (O_457,N_8259,N_9209);
nor UO_458 (O_458,N_9382,N_7948);
and UO_459 (O_459,N_7650,N_8137);
and UO_460 (O_460,N_8004,N_8749);
nand UO_461 (O_461,N_8676,N_9222);
nor UO_462 (O_462,N_8330,N_9314);
or UO_463 (O_463,N_9818,N_8126);
or UO_464 (O_464,N_8441,N_8541);
nand UO_465 (O_465,N_8806,N_8474);
and UO_466 (O_466,N_7549,N_9488);
nand UO_467 (O_467,N_9619,N_8791);
nor UO_468 (O_468,N_9733,N_8362);
xnor UO_469 (O_469,N_8469,N_8268);
or UO_470 (O_470,N_9137,N_9491);
or UO_471 (O_471,N_9487,N_7631);
or UO_472 (O_472,N_9138,N_8627);
and UO_473 (O_473,N_8517,N_8231);
and UO_474 (O_474,N_8855,N_9625);
and UO_475 (O_475,N_9042,N_9970);
nor UO_476 (O_476,N_8180,N_8626);
or UO_477 (O_477,N_7783,N_9262);
nand UO_478 (O_478,N_8179,N_8381);
and UO_479 (O_479,N_8745,N_7680);
or UO_480 (O_480,N_9182,N_9495);
or UO_481 (O_481,N_8363,N_9070);
or UO_482 (O_482,N_9211,N_8607);
or UO_483 (O_483,N_8701,N_8235);
nand UO_484 (O_484,N_8786,N_8893);
and UO_485 (O_485,N_8636,N_7700);
nand UO_486 (O_486,N_8515,N_8801);
nand UO_487 (O_487,N_9307,N_9760);
nor UO_488 (O_488,N_9708,N_8695);
nor UO_489 (O_489,N_8466,N_7866);
and UO_490 (O_490,N_8193,N_8377);
nand UO_491 (O_491,N_9208,N_9829);
or UO_492 (O_492,N_8889,N_8535);
nand UO_493 (O_493,N_7607,N_9002);
and UO_494 (O_494,N_9797,N_8341);
or UO_495 (O_495,N_7793,N_7756);
or UO_496 (O_496,N_9626,N_9583);
xnor UO_497 (O_497,N_7888,N_8099);
nor UO_498 (O_498,N_9077,N_8062);
nor UO_499 (O_499,N_8904,N_8545);
and UO_500 (O_500,N_9026,N_9996);
and UO_501 (O_501,N_9319,N_8361);
and UO_502 (O_502,N_8692,N_9449);
xnor UO_503 (O_503,N_9711,N_8144);
nor UO_504 (O_504,N_9367,N_8507);
and UO_505 (O_505,N_7721,N_7755);
xor UO_506 (O_506,N_8473,N_7739);
nor UO_507 (O_507,N_7843,N_9082);
nand UO_508 (O_508,N_8611,N_8430);
nand UO_509 (O_509,N_9481,N_9528);
and UO_510 (O_510,N_9929,N_8318);
nand UO_511 (O_511,N_9373,N_8719);
and UO_512 (O_512,N_7524,N_8274);
or UO_513 (O_513,N_9258,N_9016);
or UO_514 (O_514,N_8991,N_8723);
or UO_515 (O_515,N_7596,N_8325);
nand UO_516 (O_516,N_9240,N_8123);
nand UO_517 (O_517,N_7988,N_9570);
or UO_518 (O_518,N_8757,N_9178);
nor UO_519 (O_519,N_8397,N_9061);
nor UO_520 (O_520,N_8940,N_9276);
nor UO_521 (O_521,N_7773,N_9133);
or UO_522 (O_522,N_7894,N_8848);
and UO_523 (O_523,N_9542,N_8908);
nor UO_524 (O_524,N_9284,N_8554);
or UO_525 (O_525,N_9924,N_7967);
and UO_526 (O_526,N_8782,N_9350);
nand UO_527 (O_527,N_9946,N_8409);
or UO_528 (O_528,N_8067,N_7920);
or UO_529 (O_529,N_7613,N_8914);
nor UO_530 (O_530,N_8836,N_7619);
and UO_531 (O_531,N_8291,N_8900);
and UO_532 (O_532,N_8921,N_8195);
nor UO_533 (O_533,N_8760,N_9811);
and UO_534 (O_534,N_9175,N_7603);
nand UO_535 (O_535,N_7678,N_8661);
nor UO_536 (O_536,N_8376,N_9802);
or UO_537 (O_537,N_9651,N_9148);
and UO_538 (O_538,N_7885,N_8465);
or UO_539 (O_539,N_9162,N_8838);
and UO_540 (O_540,N_8857,N_9913);
nand UO_541 (O_541,N_7599,N_7808);
or UO_542 (O_542,N_7926,N_9656);
and UO_543 (O_543,N_7731,N_9269);
or UO_544 (O_544,N_9345,N_7541);
xor UO_545 (O_545,N_8310,N_8725);
nand UO_546 (O_546,N_8505,N_8240);
nor UO_547 (O_547,N_9762,N_9024);
nor UO_548 (O_548,N_8427,N_8996);
or UO_549 (O_549,N_8527,N_7958);
nor UO_550 (O_550,N_8025,N_9458);
nor UO_551 (O_551,N_9129,N_9509);
or UO_552 (O_552,N_8312,N_8297);
nor UO_553 (O_553,N_7640,N_8563);
or UO_554 (O_554,N_7909,N_9220);
and UO_555 (O_555,N_8443,N_9905);
nand UO_556 (O_556,N_9331,N_8920);
and UO_557 (O_557,N_7604,N_9501);
nand UO_558 (O_558,N_7612,N_9067);
and UO_559 (O_559,N_9235,N_9738);
or UO_560 (O_560,N_8052,N_8122);
nand UO_561 (O_561,N_8686,N_8603);
or UO_562 (O_562,N_7919,N_9985);
nor UO_563 (O_563,N_8086,N_8013);
xor UO_564 (O_564,N_7743,N_9428);
and UO_565 (O_565,N_9170,N_9020);
and UO_566 (O_566,N_8559,N_9265);
or UO_567 (O_567,N_7623,N_9853);
and UO_568 (O_568,N_8644,N_8938);
or UO_569 (O_569,N_8548,N_8704);
xor UO_570 (O_570,N_9816,N_7538);
or UO_571 (O_571,N_8169,N_8614);
and UO_572 (O_572,N_8586,N_9456);
or UO_573 (O_573,N_8219,N_8647);
nand UO_574 (O_574,N_8797,N_9223);
nor UO_575 (O_575,N_9281,N_8566);
or UO_576 (O_576,N_9195,N_9593);
and UO_577 (O_577,N_7717,N_7625);
nor UO_578 (O_578,N_9839,N_7935);
nand UO_579 (O_579,N_7982,N_8173);
and UO_580 (O_580,N_9419,N_8009);
nor UO_581 (O_581,N_7992,N_9808);
nand UO_582 (O_582,N_8671,N_8202);
or UO_583 (O_583,N_8211,N_8721);
and UO_584 (O_584,N_9144,N_7747);
nand UO_585 (O_585,N_8436,N_9048);
and UO_586 (O_586,N_8633,N_7896);
nor UO_587 (O_587,N_9887,N_7624);
and UO_588 (O_588,N_9008,N_8304);
nand UO_589 (O_589,N_7724,N_9707);
nor UO_590 (O_590,N_8342,N_7719);
and UO_591 (O_591,N_9062,N_9809);
nand UO_592 (O_592,N_9311,N_9282);
nor UO_593 (O_593,N_7544,N_7675);
or UO_594 (O_594,N_7665,N_8305);
and UO_595 (O_595,N_7714,N_7626);
nor UO_596 (O_596,N_9369,N_8538);
nor UO_597 (O_597,N_8014,N_7653);
or UO_598 (O_598,N_9745,N_8589);
nand UO_599 (O_599,N_9834,N_9721);
or UO_600 (O_600,N_8393,N_8963);
or UO_601 (O_601,N_8712,N_9368);
nand UO_602 (O_602,N_9186,N_9521);
nor UO_603 (O_603,N_8977,N_8814);
or UO_604 (O_604,N_8294,N_9253);
nand UO_605 (O_605,N_9514,N_8043);
xnor UO_606 (O_606,N_8271,N_7972);
and UO_607 (O_607,N_9512,N_8328);
and UO_608 (O_608,N_9112,N_9677);
nand UO_609 (O_609,N_9165,N_9470);
nand UO_610 (O_610,N_9659,N_8499);
nor UO_611 (O_611,N_8451,N_7985);
nand UO_612 (O_612,N_9066,N_9306);
nor UO_613 (O_613,N_9551,N_8018);
nand UO_614 (O_614,N_7908,N_9781);
nor UO_615 (O_615,N_7682,N_9754);
and UO_616 (O_616,N_9606,N_8982);
nand UO_617 (O_617,N_9459,N_9012);
nor UO_618 (O_618,N_9713,N_8321);
and UO_619 (O_619,N_7565,N_9565);
and UO_620 (O_620,N_8101,N_8148);
or UO_621 (O_621,N_7705,N_9483);
nor UO_622 (O_622,N_8593,N_9780);
nand UO_623 (O_623,N_9375,N_9128);
and UO_624 (O_624,N_8389,N_8008);
or UO_625 (O_625,N_9261,N_9346);
and UO_626 (O_626,N_9294,N_8557);
and UO_627 (O_627,N_7883,N_7568);
xor UO_628 (O_628,N_9420,N_8151);
and UO_629 (O_629,N_8931,N_7513);
and UO_630 (O_630,N_8902,N_9746);
and UO_631 (O_631,N_9654,N_9151);
nand UO_632 (O_632,N_9380,N_8000);
nor UO_633 (O_633,N_7500,N_7782);
nand UO_634 (O_634,N_8705,N_8619);
nor UO_635 (O_635,N_9413,N_7907);
and UO_636 (O_636,N_9893,N_8734);
xor UO_637 (O_637,N_7598,N_8484);
nand UO_638 (O_638,N_9305,N_7670);
nor UO_639 (O_639,N_7912,N_9752);
nor UO_640 (O_640,N_9498,N_7869);
nand UO_641 (O_641,N_8916,N_8476);
or UO_642 (O_642,N_7616,N_8864);
and UO_643 (O_643,N_9440,N_9406);
nand UO_644 (O_644,N_8953,N_9763);
and UO_645 (O_645,N_9663,N_7602);
and UO_646 (O_646,N_8356,N_9793);
nand UO_647 (O_647,N_7811,N_8058);
or UO_648 (O_648,N_8070,N_8460);
and UO_649 (O_649,N_9670,N_8521);
nand UO_650 (O_650,N_9278,N_8482);
or UO_651 (O_651,N_8939,N_9742);
nor UO_652 (O_652,N_7941,N_9238);
nand UO_653 (O_653,N_9798,N_9807);
or UO_654 (O_654,N_7683,N_8001);
xnor UO_655 (O_655,N_9296,N_9453);
or UO_656 (O_656,N_8246,N_7854);
and UO_657 (O_657,N_9814,N_8998);
and UO_658 (O_658,N_8433,N_9765);
nand UO_659 (O_659,N_8815,N_7676);
nand UO_660 (O_660,N_8746,N_9194);
and UO_661 (O_661,N_9045,N_7829);
nand UO_662 (O_662,N_8442,N_9859);
and UO_663 (O_663,N_9824,N_9568);
and UO_664 (O_664,N_8629,N_7768);
or UO_665 (O_665,N_7657,N_8111);
or UO_666 (O_666,N_8171,N_9231);
or UO_667 (O_667,N_8212,N_8550);
and UO_668 (O_668,N_9885,N_7803);
and UO_669 (O_669,N_8585,N_8252);
nor UO_670 (O_670,N_7991,N_8683);
or UO_671 (O_671,N_7939,N_9614);
nor UO_672 (O_672,N_9139,N_8061);
and UO_673 (O_673,N_8880,N_9599);
nand UO_674 (O_674,N_8800,N_7643);
or UO_675 (O_675,N_9125,N_9884);
nand UO_676 (O_676,N_9532,N_9320);
nor UO_677 (O_677,N_9852,N_8301);
nand UO_678 (O_678,N_9493,N_7861);
nor UO_679 (O_679,N_9329,N_9530);
nor UO_680 (O_680,N_9507,N_7970);
nand UO_681 (O_681,N_8747,N_7925);
and UO_682 (O_682,N_9104,N_8870);
or UO_683 (O_683,N_9471,N_9993);
and UO_684 (O_684,N_9699,N_8471);
nor UO_685 (O_685,N_9983,N_8349);
nand UO_686 (O_686,N_9199,N_8248);
xor UO_687 (O_687,N_7828,N_9007);
xnor UO_688 (O_688,N_8472,N_9212);
and UO_689 (O_689,N_9667,N_9569);
or UO_690 (O_690,N_8487,N_8296);
or UO_691 (O_691,N_9973,N_7748);
nor UO_692 (O_692,N_8412,N_8781);
nand UO_693 (O_693,N_7734,N_8547);
nand UO_694 (O_694,N_9058,N_7501);
nor UO_695 (O_695,N_9725,N_9372);
nor UO_696 (O_696,N_8758,N_9805);
nor UO_697 (O_697,N_9356,N_9197);
nand UO_698 (O_698,N_7580,N_9405);
and UO_699 (O_699,N_9510,N_8082);
and UO_700 (O_700,N_7943,N_9715);
nor UO_701 (O_701,N_9410,N_8853);
and UO_702 (O_702,N_9432,N_9120);
nand UO_703 (O_703,N_9218,N_9228);
nor UO_704 (O_704,N_7706,N_8371);
nand UO_705 (O_705,N_8046,N_9926);
or UO_706 (O_706,N_7502,N_9113);
nand UO_707 (O_707,N_8315,N_8158);
and UO_708 (O_708,N_8795,N_7848);
nor UO_709 (O_709,N_8134,N_9922);
nor UO_710 (O_710,N_8540,N_9337);
nor UO_711 (O_711,N_9879,N_8865);
or UO_712 (O_712,N_9610,N_8155);
nor UO_713 (O_713,N_7644,N_8339);
or UO_714 (O_714,N_7600,N_7641);
nor UO_715 (O_715,N_7744,N_8255);
and UO_716 (O_716,N_8850,N_9299);
nand UO_717 (O_717,N_8884,N_8495);
nor UO_718 (O_718,N_7966,N_8491);
nand UO_719 (O_719,N_9904,N_9545);
or UO_720 (O_720,N_8875,N_9298);
and UO_721 (O_721,N_9378,N_8937);
or UO_722 (O_722,N_7794,N_9213);
and UO_723 (O_723,N_8078,N_9390);
and UO_724 (O_724,N_7749,N_9630);
or UO_725 (O_725,N_9473,N_9494);
nand UO_726 (O_726,N_9883,N_8395);
and UO_727 (O_727,N_7548,N_9478);
and UO_728 (O_728,N_9293,N_8687);
and UO_729 (O_729,N_8653,N_7777);
or UO_730 (O_730,N_8946,N_8773);
nand UO_731 (O_731,N_8679,N_8681);
nor UO_732 (O_732,N_9053,N_8654);
nor UO_733 (O_733,N_9643,N_8556);
nor UO_734 (O_734,N_8599,N_9207);
or UO_735 (O_735,N_9909,N_8744);
and UO_736 (O_736,N_9529,N_9863);
or UO_737 (O_737,N_9617,N_8971);
or UO_738 (O_738,N_9691,N_7578);
xor UO_739 (O_739,N_8358,N_9063);
nand UO_740 (O_740,N_8717,N_7618);
or UO_741 (O_741,N_9272,N_9800);
nand UO_742 (O_742,N_8722,N_9838);
nand UO_743 (O_743,N_8657,N_9219);
nand UO_744 (O_744,N_8592,N_9547);
xor UO_745 (O_745,N_9559,N_7834);
nand UO_746 (O_746,N_8063,N_8655);
and UO_747 (O_747,N_8878,N_8026);
nor UO_748 (O_748,N_8384,N_9758);
nand UO_749 (O_749,N_8957,N_8659);
nor UO_750 (O_750,N_7769,N_9562);
and UO_751 (O_751,N_9098,N_8768);
or UO_752 (O_752,N_7880,N_9679);
nand UO_753 (O_753,N_8136,N_9490);
nor UO_754 (O_754,N_9001,N_8793);
or UO_755 (O_755,N_7846,N_9078);
or UO_756 (O_756,N_8087,N_7911);
or UO_757 (O_757,N_7815,N_8477);
nor UO_758 (O_758,N_9003,N_9712);
or UO_759 (O_759,N_8287,N_9789);
xor UO_760 (O_760,N_7605,N_8980);
or UO_761 (O_761,N_8876,N_9943);
or UO_762 (O_762,N_9039,N_7978);
or UO_763 (O_763,N_9566,N_9698);
or UO_764 (O_764,N_9988,N_9489);
nor UO_765 (O_765,N_9264,N_9748);
nand UO_766 (O_766,N_7693,N_9333);
or UO_767 (O_767,N_9972,N_8799);
nor UO_768 (O_768,N_7778,N_8660);
nand UO_769 (O_769,N_8820,N_7821);
nand UO_770 (O_770,N_8767,N_8143);
or UO_771 (O_771,N_8955,N_7733);
and UO_772 (O_772,N_8282,N_8470);
and UO_773 (O_773,N_9646,N_9523);
nand UO_774 (O_774,N_9167,N_8827);
nand UO_775 (O_775,N_9295,N_8894);
and UO_776 (O_776,N_8334,N_8720);
nand UO_777 (O_777,N_8630,N_7771);
nor UO_778 (O_778,N_9234,N_9102);
or UO_779 (O_779,N_9273,N_9110);
or UO_780 (O_780,N_9628,N_8508);
nand UO_781 (O_781,N_8973,N_7918);
nor UO_782 (O_782,N_8771,N_8068);
or UO_783 (O_783,N_7661,N_7537);
or UO_784 (O_784,N_7816,N_8573);
and UO_785 (O_785,N_8352,N_9919);
and UO_786 (O_786,N_8662,N_8327);
and UO_787 (O_787,N_7809,N_8003);
or UO_788 (O_788,N_8279,N_8432);
or UO_789 (O_789,N_9842,N_8832);
nor UO_790 (O_790,N_8276,N_9655);
or UO_791 (O_791,N_9203,N_9072);
or UO_792 (O_792,N_8715,N_7722);
or UO_793 (O_793,N_7882,N_7788);
nor UO_794 (O_794,N_9025,N_9198);
and UO_795 (O_795,N_9558,N_9348);
and UO_796 (O_796,N_8926,N_9525);
and UO_797 (O_797,N_8551,N_8950);
and UO_798 (O_798,N_9461,N_9088);
nand UO_799 (O_799,N_7845,N_8641);
and UO_800 (O_800,N_8254,N_8813);
nor UO_801 (O_801,N_7577,N_8710);
nand UO_802 (O_802,N_8192,N_9804);
nand UO_803 (O_803,N_8502,N_9040);
and UO_804 (O_804,N_8718,N_9548);
nor UO_805 (O_805,N_7715,N_7923);
xor UO_806 (O_806,N_9279,N_9856);
nand UO_807 (O_807,N_8168,N_8872);
xnor UO_808 (O_808,N_8108,N_8822);
or UO_809 (O_809,N_8867,N_7900);
nand UO_810 (O_810,N_7944,N_8525);
or UO_811 (O_811,N_8897,N_9038);
xor UO_812 (O_812,N_8346,N_9041);
nand UO_813 (O_813,N_8223,N_8845);
and UO_814 (O_814,N_9847,N_8320);
xor UO_815 (O_815,N_8631,N_8761);
and UO_816 (O_816,N_8135,N_9868);
and UO_817 (O_817,N_7795,N_9123);
and UO_818 (O_818,N_8438,N_9744);
or UO_819 (O_819,N_8170,N_9444);
xnor UO_820 (O_820,N_9775,N_7852);
nor UO_821 (O_821,N_8083,N_7723);
and UO_822 (O_822,N_8756,N_9894);
and UO_823 (O_823,N_8601,N_8343);
or UO_824 (O_824,N_9825,N_9577);
nor UO_825 (O_825,N_8054,N_8269);
nor UO_826 (O_826,N_9439,N_7971);
nor UO_827 (O_827,N_8500,N_9739);
and UO_828 (O_828,N_9196,N_9043);
nand UO_829 (O_829,N_8383,N_8216);
nor UO_830 (O_830,N_8329,N_9697);
nor UO_831 (O_831,N_7593,N_8039);
nand UO_832 (O_832,N_8149,N_9263);
xor UO_833 (O_833,N_8214,N_9179);
nand UO_834 (O_834,N_7691,N_8245);
and UO_835 (O_835,N_7979,N_7799);
xor UO_836 (O_836,N_9914,N_9991);
or UO_837 (O_837,N_9735,N_7622);
nand UO_838 (O_838,N_8588,N_9513);
nor UO_839 (O_839,N_7585,N_8748);
nand UO_840 (O_840,N_7892,N_9858);
or UO_841 (O_841,N_9106,N_9429);
nor UO_842 (O_842,N_9326,N_8615);
or UO_843 (O_843,N_7822,N_8674);
and UO_844 (O_844,N_8234,N_8265);
xnor UO_845 (O_845,N_9092,N_7698);
and UO_846 (O_846,N_9418,N_7840);
or UO_847 (O_847,N_7936,N_8742);
nor UO_848 (O_848,N_8735,N_9967);
nor UO_849 (O_849,N_8837,N_7582);
and UO_850 (O_850,N_8956,N_7859);
nor UO_851 (O_851,N_9803,N_8577);
nand UO_852 (O_852,N_7994,N_7877);
or UO_853 (O_853,N_8688,N_8910);
or UO_854 (O_854,N_8367,N_7570);
nand UO_855 (O_855,N_9134,N_9740);
xnor UO_856 (O_856,N_9465,N_8475);
or UO_857 (O_857,N_8668,N_9187);
nor UO_858 (O_858,N_8796,N_8898);
nand UO_859 (O_859,N_7586,N_9773);
nand UO_860 (O_860,N_8394,N_9054);
and UO_861 (O_861,N_8714,N_8351);
nor UO_862 (O_862,N_9903,N_9068);
nor UO_863 (O_863,N_9511,N_9386);
and UO_864 (O_864,N_9751,N_8967);
and UO_865 (O_865,N_9426,N_9141);
or UO_866 (O_866,N_8100,N_9157);
and UO_867 (O_867,N_7922,N_9457);
and UO_868 (O_868,N_7718,N_8622);
and UO_869 (O_869,N_7938,N_8229);
nand UO_870 (O_870,N_7503,N_8883);
and UO_871 (O_871,N_8696,N_8769);
or UO_872 (O_872,N_8501,N_8826);
nor UO_873 (O_873,N_9580,N_8531);
or UO_874 (O_874,N_7993,N_8121);
nand UO_875 (O_875,N_7647,N_8932);
or UO_876 (O_876,N_8415,N_8579);
and UO_877 (O_877,N_7581,N_8498);
nand UO_878 (O_878,N_8283,N_9882);
or UO_879 (O_879,N_8303,N_8684);
and UO_880 (O_880,N_9011,N_9649);
nor UO_881 (O_881,N_8221,N_8264);
nor UO_882 (O_882,N_9422,N_9388);
nand UO_883 (O_883,N_8700,N_7692);
xor UO_884 (O_884,N_9014,N_8191);
nand UO_885 (O_885,N_8726,N_9484);
or UO_886 (O_886,N_8075,N_7632);
nand UO_887 (O_887,N_7921,N_9103);
nor UO_888 (O_888,N_7519,N_8401);
and UO_889 (O_889,N_9159,N_7887);
nand UO_890 (O_890,N_7646,N_9233);
or UO_891 (O_891,N_9206,N_9362);
or UO_892 (O_892,N_8528,N_7862);
or UO_893 (O_893,N_8418,N_8613);
and UO_894 (O_894,N_7505,N_8979);
nor UO_895 (O_895,N_9214,N_7555);
or UO_896 (O_896,N_9976,N_9180);
or UO_897 (O_897,N_9031,N_9371);
or UO_898 (O_898,N_9140,N_8224);
nor UO_899 (O_899,N_9957,N_7858);
and UO_900 (O_900,N_7526,N_7891);
and UO_901 (O_901,N_9620,N_7962);
or UO_902 (O_902,N_9965,N_8106);
nand UO_903 (O_903,N_9778,N_8272);
or UO_904 (O_904,N_7884,N_7518);
nand UO_905 (O_905,N_7977,N_8632);
nand UO_906 (O_906,N_8915,N_9519);
nand UO_907 (O_907,N_7583,N_9121);
nand UO_908 (O_908,N_9087,N_7831);
and UO_909 (O_909,N_9096,N_9005);
nor UO_910 (O_910,N_9631,N_9650);
nor UO_911 (O_911,N_7917,N_9567);
nand UO_912 (O_912,N_7686,N_9837);
nand UO_913 (O_913,N_9424,N_8901);
nor UO_914 (O_914,N_7629,N_7787);
nand UO_915 (O_915,N_7688,N_8147);
nor UO_916 (O_916,N_8059,N_8016);
nand UO_917 (O_917,N_8416,N_7766);
and UO_918 (O_918,N_8569,N_9268);
nor UO_919 (O_919,N_9492,N_9100);
and UO_920 (O_920,N_8187,N_7677);
or UO_921 (O_921,N_9205,N_7801);
nor UO_922 (O_922,N_8196,N_9636);
nor UO_923 (O_923,N_7648,N_7981);
nand UO_924 (O_924,N_8142,N_7910);
nand UO_925 (O_925,N_7933,N_9990);
or UO_926 (O_926,N_9515,N_9332);
and UO_927 (O_927,N_9881,N_7872);
nor UO_928 (O_928,N_9409,N_9682);
nand UO_929 (O_929,N_8922,N_7710);
nand UO_930 (O_930,N_8045,N_9360);
and UO_931 (O_931,N_9303,N_9190);
nor UO_932 (O_932,N_9910,N_9952);
or UO_933 (O_933,N_8094,N_8759);
or UO_934 (O_934,N_8153,N_9897);
nor UO_935 (O_935,N_9183,N_7881);
nor UO_936 (O_936,N_8959,N_7684);
or UO_937 (O_937,N_7671,N_8978);
or UO_938 (O_938,N_9607,N_9064);
or UO_939 (O_939,N_8360,N_9694);
nand UO_940 (O_940,N_8249,N_8763);
nand UO_941 (O_941,N_8468,N_8233);
and UO_942 (O_942,N_9486,N_7767);
and UO_943 (O_943,N_8860,N_8903);
or UO_944 (O_944,N_8711,N_9239);
or UO_945 (O_945,N_9578,N_8817);
nor UO_946 (O_946,N_9030,N_9779);
or UO_947 (O_947,N_8400,N_8802);
and UO_948 (O_948,N_9546,N_9961);
nand UO_949 (O_949,N_8284,N_9660);
nand UO_950 (O_950,N_9290,N_9605);
and UO_951 (O_951,N_9747,N_7874);
or UO_952 (O_952,N_7946,N_9813);
and UO_953 (O_953,N_7610,N_7836);
nand UO_954 (O_954,N_8382,N_9635);
or UO_955 (O_955,N_7668,N_9004);
xor UO_956 (O_956,N_9315,N_8990);
or UO_957 (O_957,N_8703,N_8194);
or UO_958 (O_958,N_9994,N_8034);
and UO_959 (O_959,N_8913,N_8639);
or UO_960 (O_960,N_7893,N_9033);
and UO_961 (O_961,N_9810,N_9843);
nor UO_962 (O_962,N_9237,N_9639);
or UO_963 (O_963,N_9051,N_8947);
nor UO_964 (O_964,N_7649,N_8150);
and UO_965 (O_965,N_8311,N_7841);
nor UO_966 (O_966,N_9764,N_7673);
nor UO_967 (O_967,N_9117,N_7534);
nor UO_968 (O_968,N_8787,N_8069);
and UO_969 (O_969,N_9217,N_9757);
nand UO_970 (O_970,N_8077,N_8053);
nand UO_971 (O_971,N_8811,N_8298);
nor UO_972 (O_972,N_8568,N_9683);
nor UO_973 (O_973,N_8243,N_9895);
or UO_974 (O_974,N_9414,N_8842);
nand UO_975 (O_975,N_9536,N_9908);
and UO_976 (O_976,N_7804,N_9164);
nor UO_977 (O_977,N_7849,N_9522);
nand UO_978 (O_978,N_8109,N_9951);
nor UO_979 (O_979,N_8423,N_7832);
nor UO_980 (O_980,N_8888,N_7751);
nor UO_981 (O_981,N_8316,N_7931);
nand UO_982 (O_982,N_9274,N_8313);
and UO_983 (O_983,N_9537,N_9469);
or UO_984 (O_984,N_9266,N_8390);
and UO_985 (O_985,N_8429,N_9158);
nor UO_986 (O_986,N_8833,N_7776);
or UO_987 (O_987,N_9535,N_8197);
nor UO_988 (O_988,N_8584,N_9550);
and UO_989 (O_989,N_7780,N_8222);
or UO_990 (O_990,N_8028,N_7522);
and UO_991 (O_991,N_8829,N_7957);
nor UO_992 (O_992,N_8565,N_9090);
or UO_993 (O_993,N_9734,N_9109);
nor UO_994 (O_994,N_8941,N_8637);
nor UO_995 (O_995,N_8819,N_8892);
or UO_996 (O_996,N_8572,N_7508);
nor UO_997 (O_997,N_8047,N_9609);
or UO_998 (O_998,N_7940,N_8669);
and UO_999 (O_999,N_8338,N_9114);
or UO_1000 (O_1000,N_8907,N_9873);
nand UO_1001 (O_1001,N_9169,N_8727);
or UO_1002 (O_1002,N_7759,N_9366);
and UO_1003 (O_1003,N_8594,N_8570);
nand UO_1004 (O_1004,N_8076,N_8071);
nand UO_1005 (O_1005,N_9767,N_7611);
and UO_1006 (O_1006,N_8251,N_7566);
nor UO_1007 (O_1007,N_9271,N_8056);
or UO_1008 (O_1008,N_9324,N_9632);
and UO_1009 (O_1009,N_7579,N_8420);
nor UO_1010 (O_1010,N_8917,N_9918);
nand UO_1011 (O_1011,N_8666,N_9669);
or UO_1012 (O_1012,N_9695,N_8667);
nand UO_1013 (O_1013,N_7587,N_8232);
nor UO_1014 (O_1014,N_9065,N_9192);
or UO_1015 (O_1015,N_7681,N_8131);
or UO_1016 (O_1016,N_9115,N_7572);
nor UO_1017 (O_1017,N_8646,N_8408);
nand UO_1018 (O_1018,N_9354,N_9291);
or UO_1019 (O_1019,N_8975,N_7953);
or UO_1020 (O_1020,N_9890,N_8306);
nor UO_1021 (O_1021,N_8387,N_9575);
and UO_1022 (O_1022,N_9136,N_9417);
and UO_1023 (O_1023,N_8066,N_8402);
or UO_1024 (O_1024,N_7689,N_8780);
or UO_1025 (O_1025,N_7817,N_7819);
nor UO_1026 (O_1026,N_7664,N_9277);
or UO_1027 (O_1027,N_9083,N_9826);
or UO_1028 (O_1028,N_8775,N_8770);
or UO_1029 (O_1029,N_8359,N_8049);
or UO_1030 (O_1030,N_8132,N_7590);
nor UO_1031 (O_1031,N_9645,N_8092);
nand UO_1032 (O_1032,N_7928,N_9130);
and UO_1033 (O_1033,N_9073,N_7814);
nor UO_1034 (O_1034,N_9621,N_7905);
nor UO_1035 (O_1035,N_9107,N_9340);
and UO_1036 (O_1036,N_8010,N_8380);
xor UO_1037 (O_1037,N_9953,N_8532);
or UO_1038 (O_1038,N_8115,N_8215);
or UO_1039 (O_1039,N_8849,N_9776);
and UO_1040 (O_1040,N_7807,N_8198);
nor UO_1041 (O_1041,N_9152,N_7824);
or UO_1042 (O_1042,N_8970,N_8866);
or UO_1043 (O_1043,N_7934,N_8166);
nor UO_1044 (O_1044,N_9714,N_8386);
nor UO_1045 (O_1045,N_8824,N_9927);
nand UO_1046 (O_1046,N_8015,N_9585);
or UO_1047 (O_1047,N_9352,N_8369);
nor UO_1048 (O_1048,N_9939,N_9516);
nand UO_1049 (O_1049,N_9099,N_9685);
nand UO_1050 (O_1050,N_8370,N_7742);
nor UO_1051 (O_1051,N_8201,N_9402);
nor UO_1052 (O_1052,N_9870,N_9035);
and UO_1053 (O_1053,N_9950,N_9434);
or UO_1054 (O_1054,N_8887,N_9855);
and UO_1055 (O_1055,N_9749,N_9524);
nor UO_1056 (O_1056,N_7790,N_8107);
or UO_1057 (O_1057,N_9387,N_9232);
nor UO_1058 (O_1058,N_9009,N_8278);
or UO_1059 (O_1059,N_8578,N_9287);
and UO_1060 (O_1060,N_8999,N_9790);
nand UO_1061 (O_1061,N_9392,N_7525);
nor UO_1062 (O_1062,N_7730,N_9900);
nand UO_1063 (O_1063,N_9730,N_9245);
nand UO_1064 (O_1064,N_7531,N_8520);
nor UO_1065 (O_1065,N_9867,N_9210);
or UO_1066 (O_1066,N_7995,N_8553);
or UO_1067 (O_1067,N_9280,N_9466);
or UO_1068 (O_1068,N_8890,N_8635);
nand UO_1069 (O_1069,N_8690,N_9722);
nor UO_1070 (O_1070,N_9723,N_8079);
and UO_1071 (O_1071,N_8911,N_9385);
nand UO_1072 (O_1072,N_8840,N_8337);
or UO_1073 (O_1073,N_8595,N_9143);
and UO_1074 (O_1074,N_7736,N_8983);
nor UO_1075 (O_1075,N_9574,N_9902);
and UO_1076 (O_1076,N_8600,N_9316);
nand UO_1077 (O_1077,N_8105,N_8543);
or UO_1078 (O_1078,N_7916,N_8729);
nor UO_1079 (O_1079,N_8333,N_8207);
nor UO_1080 (O_1080,N_8456,N_9554);
or UO_1081 (O_1081,N_8625,N_8964);
nor UO_1082 (O_1082,N_9594,N_9931);
and UO_1083 (O_1083,N_8345,N_8335);
nand UO_1084 (O_1084,N_9149,N_9442);
nor UO_1085 (O_1085,N_8616,N_7627);
nand UO_1086 (O_1086,N_8702,N_8496);
or UO_1087 (O_1087,N_7949,N_7827);
nor UO_1088 (O_1088,N_9181,N_9573);
nor UO_1089 (O_1089,N_9338,N_9693);
or UO_1090 (O_1090,N_9028,N_9474);
or UO_1091 (O_1091,N_9934,N_7890);
nand UO_1092 (O_1092,N_8230,N_9932);
or UO_1093 (O_1093,N_8292,N_9018);
or UO_1094 (O_1094,N_9596,N_9355);
or UO_1095 (O_1095,N_9672,N_9597);
and UO_1096 (O_1096,N_7529,N_9540);
nand UO_1097 (O_1097,N_8972,N_8011);
nor UO_1098 (O_1098,N_8874,N_9962);
and UO_1099 (O_1099,N_8580,N_8405);
nand UO_1100 (O_1100,N_7950,N_7980);
and UO_1101 (O_1101,N_8391,N_9427);
nor UO_1102 (O_1102,N_7711,N_9480);
or UO_1103 (O_1103,N_9799,N_9095);
or UO_1104 (O_1104,N_7932,N_9283);
and UO_1105 (O_1105,N_9971,N_7635);
or UO_1106 (O_1106,N_7996,N_8006);
or UO_1107 (O_1107,N_9344,N_8549);
or UO_1108 (O_1108,N_9995,N_7542);
and UO_1109 (O_1109,N_8533,N_7685);
or UO_1110 (O_1110,N_9831,N_9539);
nor UO_1111 (O_1111,N_7651,N_9288);
nand UO_1112 (O_1112,N_8396,N_9784);
or UO_1113 (O_1113,N_9774,N_7999);
nand UO_1114 (O_1114,N_9938,N_9618);
and UO_1115 (O_1115,N_9661,N_7839);
nor UO_1116 (O_1116,N_9935,N_9451);
or UO_1117 (O_1117,N_9518,N_9019);
nor UO_1118 (O_1118,N_8095,N_9921);
and UO_1119 (O_1119,N_9464,N_9652);
nor UO_1120 (O_1120,N_9017,N_8256);
nand UO_1121 (O_1121,N_7545,N_8392);
and UO_1122 (O_1122,N_7810,N_8665);
or UO_1123 (O_1123,N_9788,N_7672);
nor UO_1124 (O_1124,N_9349,N_8244);
xnor UO_1125 (O_1125,N_9463,N_9201);
and UO_1126 (O_1126,N_9013,N_8439);
or UO_1127 (O_1127,N_8164,N_8738);
and UO_1128 (O_1128,N_8434,N_9602);
nand UO_1129 (O_1129,N_9502,N_8398);
and UO_1130 (O_1130,N_8242,N_8777);
and UO_1131 (O_1131,N_9450,N_8652);
or UO_1132 (O_1132,N_8038,N_8037);
or UO_1133 (O_1133,N_8033,N_8542);
nor UO_1134 (O_1134,N_9954,N_8302);
or UO_1135 (O_1135,N_9055,N_8167);
nand UO_1136 (O_1136,N_8332,N_9637);
and UO_1137 (O_1137,N_7543,N_9888);
xor UO_1138 (O_1138,N_8966,N_9241);
nor UO_1139 (O_1139,N_7667,N_9403);
nor UO_1140 (O_1140,N_7812,N_8186);
or UO_1141 (O_1141,N_7697,N_9726);
and UO_1142 (O_1142,N_8110,N_9436);
and UO_1143 (O_1143,N_8182,N_9379);
nor UO_1144 (O_1144,N_8952,N_8080);
and UO_1145 (O_1145,N_7567,N_7554);
nor UO_1146 (O_1146,N_9476,N_9582);
nand UO_1147 (O_1147,N_8357,N_8309);
nor UO_1148 (O_1148,N_8031,N_7961);
or UO_1149 (O_1149,N_8023,N_8608);
nand UO_1150 (O_1150,N_8816,N_9089);
and UO_1151 (O_1151,N_9553,N_9665);
or UO_1152 (O_1152,N_8591,N_7634);
nand UO_1153 (O_1153,N_8610,N_9448);
nand UO_1154 (O_1154,N_7645,N_9613);
nor UO_1155 (O_1155,N_7899,N_8582);
nor UO_1156 (O_1156,N_9499,N_8834);
nand UO_1157 (O_1157,N_7798,N_9527);
nand UO_1158 (O_1158,N_8257,N_9772);
nor UO_1159 (O_1159,N_9688,N_9247);
nand UO_1160 (O_1160,N_7930,N_9796);
or UO_1161 (O_1161,N_9564,N_8017);
nand UO_1162 (O_1162,N_8691,N_9365);
or UO_1163 (O_1163,N_9648,N_8846);
nand UO_1164 (O_1164,N_8450,N_8407);
and UO_1165 (O_1165,N_9437,N_9310);
nand UO_1166 (O_1166,N_8288,N_8651);
nand UO_1167 (O_1167,N_9094,N_8862);
or UO_1168 (O_1168,N_8792,N_7696);
nor UO_1169 (O_1169,N_8969,N_7563);
nor UO_1170 (O_1170,N_7745,N_8247);
and UO_1171 (O_1171,N_8918,N_8560);
nor UO_1172 (O_1172,N_9275,N_7779);
and UO_1173 (O_1173,N_7532,N_8308);
nand UO_1174 (O_1174,N_7740,N_8081);
nor UO_1175 (O_1175,N_8929,N_9689);
nor UO_1176 (O_1176,N_7753,N_9920);
nor UO_1177 (O_1177,N_7655,N_9116);
nor UO_1178 (O_1178,N_9260,N_7774);
nor UO_1179 (O_1179,N_7699,N_7702);
nand UO_1180 (O_1180,N_9857,N_8489);
or UO_1181 (O_1181,N_8403,N_8492);
nor UO_1182 (O_1182,N_9588,N_8084);
nand UO_1183 (O_1183,N_9357,N_8808);
nor UO_1184 (O_1184,N_9835,N_8740);
nor UO_1185 (O_1185,N_9227,N_9358);
nor UO_1186 (O_1186,N_9820,N_8340);
nor UO_1187 (O_1187,N_9301,N_8805);
or UO_1188 (O_1188,N_8881,N_8024);
and UO_1189 (O_1189,N_8368,N_9153);
nand UO_1190 (O_1190,N_9503,N_9674);
nor UO_1191 (O_1191,N_9309,N_9912);
or UO_1192 (O_1192,N_9022,N_8650);
or UO_1193 (O_1193,N_8604,N_9335);
nand UO_1194 (O_1194,N_8493,N_9658);
and UO_1195 (O_1195,N_8658,N_8485);
nor UO_1196 (O_1196,N_9132,N_8289);
nand UO_1197 (O_1197,N_9741,N_8128);
and UO_1198 (O_1198,N_9563,N_9840);
nor UO_1199 (O_1199,N_9081,N_7761);
nor UO_1200 (O_1200,N_8905,N_8789);
nand UO_1201 (O_1201,N_9079,N_8935);
nor UO_1202 (O_1202,N_7820,N_9105);
nor UO_1203 (O_1203,N_8093,N_7606);
or UO_1204 (O_1204,N_7857,N_8597);
and UO_1205 (O_1205,N_9865,N_7558);
or UO_1206 (O_1206,N_8314,N_8987);
nor UO_1207 (O_1207,N_8448,N_7906);
nor UO_1208 (O_1208,N_8503,N_8113);
nand UO_1209 (O_1209,N_9936,N_9916);
or UO_1210 (O_1210,N_9394,N_8962);
nand UO_1211 (O_1211,N_7929,N_8462);
or UO_1212 (O_1212,N_9557,N_8280);
nand UO_1213 (O_1213,N_9191,N_9441);
or UO_1214 (O_1214,N_8753,N_8425);
and UO_1215 (O_1215,N_8035,N_9093);
nand UO_1216 (O_1216,N_9821,N_8587);
and UO_1217 (O_1217,N_9071,N_8490);
nand UO_1218 (O_1218,N_7802,N_9875);
and UO_1219 (O_1219,N_8457,N_9544);
nand UO_1220 (O_1220,N_8643,N_8152);
or UO_1221 (O_1221,N_7504,N_8253);
or UO_1222 (O_1222,N_8707,N_8428);
xor UO_1223 (O_1223,N_8976,N_8699);
nor UO_1224 (O_1224,N_9822,N_7951);
or UO_1225 (O_1225,N_8185,N_9787);
and UO_1226 (O_1226,N_7752,N_9608);
or UO_1227 (O_1227,N_9969,N_8751);
and UO_1228 (O_1228,N_9849,N_9552);
and UO_1229 (O_1229,N_7895,N_9736);
nand UO_1230 (O_1230,N_9874,N_7823);
nor UO_1231 (O_1231,N_8821,N_7924);
and UO_1232 (O_1232,N_9906,N_7658);
or UO_1233 (O_1233,N_9251,N_8030);
or UO_1234 (O_1234,N_8029,N_8209);
nand UO_1235 (O_1235,N_9794,N_7589);
or UO_1236 (O_1236,N_9154,N_8621);
or UO_1237 (O_1237,N_7575,N_8286);
nor UO_1238 (O_1238,N_9084,N_9173);
nor UO_1239 (O_1239,N_8154,N_9891);
and UO_1240 (O_1240,N_9997,N_9353);
and UO_1241 (O_1241,N_7595,N_7669);
and UO_1242 (O_1242,N_7937,N_9399);
and UO_1243 (O_1243,N_8949,N_8204);
nor UO_1244 (O_1244,N_7546,N_7998);
nor UO_1245 (O_1245,N_9520,N_8447);
and UO_1246 (O_1246,N_7707,N_8754);
or UO_1247 (O_1247,N_9911,N_8762);
or UO_1248 (O_1248,N_9591,N_8783);
or UO_1249 (O_1249,N_8928,N_7952);
or UO_1250 (O_1250,N_8615,N_9906);
nor UO_1251 (O_1251,N_8390,N_8488);
or UO_1252 (O_1252,N_9806,N_9226);
or UO_1253 (O_1253,N_7886,N_9407);
or UO_1254 (O_1254,N_9999,N_9611);
nand UO_1255 (O_1255,N_8896,N_8214);
xnor UO_1256 (O_1256,N_7872,N_8192);
or UO_1257 (O_1257,N_7651,N_7662);
or UO_1258 (O_1258,N_7584,N_8955);
and UO_1259 (O_1259,N_9020,N_7529);
or UO_1260 (O_1260,N_9494,N_8222);
nand UO_1261 (O_1261,N_9124,N_8237);
nor UO_1262 (O_1262,N_9113,N_8806);
nor UO_1263 (O_1263,N_9106,N_9681);
or UO_1264 (O_1264,N_8794,N_8072);
or UO_1265 (O_1265,N_9949,N_8231);
or UO_1266 (O_1266,N_8720,N_8987);
and UO_1267 (O_1267,N_7925,N_7689);
nor UO_1268 (O_1268,N_9819,N_8361);
nor UO_1269 (O_1269,N_7881,N_7565);
and UO_1270 (O_1270,N_9389,N_8098);
nand UO_1271 (O_1271,N_9054,N_7910);
nand UO_1272 (O_1272,N_7803,N_9497);
nor UO_1273 (O_1273,N_9803,N_9833);
and UO_1274 (O_1274,N_8950,N_9323);
or UO_1275 (O_1275,N_7979,N_9441);
and UO_1276 (O_1276,N_7804,N_8078);
or UO_1277 (O_1277,N_9091,N_9315);
nor UO_1278 (O_1278,N_9320,N_8135);
and UO_1279 (O_1279,N_8072,N_8879);
and UO_1280 (O_1280,N_8608,N_8860);
nand UO_1281 (O_1281,N_9303,N_9311);
and UO_1282 (O_1282,N_8104,N_7772);
nor UO_1283 (O_1283,N_9649,N_8740);
nor UO_1284 (O_1284,N_9691,N_9690);
and UO_1285 (O_1285,N_9653,N_9347);
and UO_1286 (O_1286,N_7957,N_8296);
and UO_1287 (O_1287,N_9234,N_9233);
nor UO_1288 (O_1288,N_9690,N_9649);
nand UO_1289 (O_1289,N_9983,N_9322);
and UO_1290 (O_1290,N_7825,N_9920);
nor UO_1291 (O_1291,N_9839,N_8275);
nand UO_1292 (O_1292,N_9319,N_9771);
nor UO_1293 (O_1293,N_8848,N_7982);
nor UO_1294 (O_1294,N_8132,N_7525);
nand UO_1295 (O_1295,N_8901,N_8543);
and UO_1296 (O_1296,N_8930,N_8545);
and UO_1297 (O_1297,N_9268,N_8939);
nor UO_1298 (O_1298,N_9079,N_9367);
and UO_1299 (O_1299,N_7772,N_7681);
nand UO_1300 (O_1300,N_9953,N_9046);
nor UO_1301 (O_1301,N_8393,N_8560);
and UO_1302 (O_1302,N_7762,N_9823);
nor UO_1303 (O_1303,N_7682,N_9324);
nand UO_1304 (O_1304,N_9874,N_9138);
and UO_1305 (O_1305,N_9944,N_9675);
and UO_1306 (O_1306,N_9722,N_9092);
or UO_1307 (O_1307,N_9919,N_8079);
or UO_1308 (O_1308,N_7512,N_9482);
or UO_1309 (O_1309,N_8676,N_9010);
and UO_1310 (O_1310,N_8593,N_9608);
or UO_1311 (O_1311,N_9960,N_9306);
and UO_1312 (O_1312,N_8646,N_8591);
and UO_1313 (O_1313,N_8734,N_7958);
and UO_1314 (O_1314,N_9980,N_8331);
and UO_1315 (O_1315,N_9527,N_8486);
and UO_1316 (O_1316,N_8720,N_9916);
nand UO_1317 (O_1317,N_9833,N_8668);
or UO_1318 (O_1318,N_9401,N_8870);
nor UO_1319 (O_1319,N_8844,N_8127);
and UO_1320 (O_1320,N_8522,N_9714);
and UO_1321 (O_1321,N_9025,N_8420);
and UO_1322 (O_1322,N_9720,N_9134);
nor UO_1323 (O_1323,N_9011,N_7653);
nor UO_1324 (O_1324,N_8820,N_7942);
xor UO_1325 (O_1325,N_8706,N_9686);
nand UO_1326 (O_1326,N_8004,N_9523);
nand UO_1327 (O_1327,N_9624,N_9274);
and UO_1328 (O_1328,N_7580,N_8076);
xor UO_1329 (O_1329,N_9431,N_9260);
nand UO_1330 (O_1330,N_8205,N_8446);
and UO_1331 (O_1331,N_8421,N_8612);
and UO_1332 (O_1332,N_9692,N_9382);
nor UO_1333 (O_1333,N_9997,N_8598);
and UO_1334 (O_1334,N_9576,N_9221);
nor UO_1335 (O_1335,N_8266,N_9995);
nor UO_1336 (O_1336,N_8051,N_8045);
nor UO_1337 (O_1337,N_9962,N_9907);
nand UO_1338 (O_1338,N_7640,N_9519);
or UO_1339 (O_1339,N_9939,N_8902);
or UO_1340 (O_1340,N_8567,N_8475);
nor UO_1341 (O_1341,N_7652,N_9113);
nand UO_1342 (O_1342,N_9355,N_8094);
nor UO_1343 (O_1343,N_8547,N_9995);
and UO_1344 (O_1344,N_9998,N_8279);
nand UO_1345 (O_1345,N_8669,N_7989);
and UO_1346 (O_1346,N_7547,N_8296);
and UO_1347 (O_1347,N_7898,N_9335);
nor UO_1348 (O_1348,N_8050,N_8966);
and UO_1349 (O_1349,N_8660,N_9046);
nand UO_1350 (O_1350,N_8347,N_9298);
nand UO_1351 (O_1351,N_8103,N_8867);
nor UO_1352 (O_1352,N_9169,N_7888);
and UO_1353 (O_1353,N_8361,N_9168);
nor UO_1354 (O_1354,N_9610,N_8259);
xnor UO_1355 (O_1355,N_8587,N_9091);
and UO_1356 (O_1356,N_9164,N_7567);
nor UO_1357 (O_1357,N_8759,N_8542);
nand UO_1358 (O_1358,N_8970,N_8376);
and UO_1359 (O_1359,N_9954,N_8952);
nand UO_1360 (O_1360,N_9977,N_8116);
nand UO_1361 (O_1361,N_7818,N_9800);
nor UO_1362 (O_1362,N_9457,N_9073);
and UO_1363 (O_1363,N_8404,N_7918);
nor UO_1364 (O_1364,N_9062,N_9303);
or UO_1365 (O_1365,N_8204,N_9962);
or UO_1366 (O_1366,N_9985,N_7719);
nor UO_1367 (O_1367,N_8672,N_8102);
nor UO_1368 (O_1368,N_9508,N_8597);
or UO_1369 (O_1369,N_9801,N_9548);
nor UO_1370 (O_1370,N_9883,N_8621);
and UO_1371 (O_1371,N_9135,N_8904);
nand UO_1372 (O_1372,N_8533,N_8829);
nand UO_1373 (O_1373,N_8155,N_9414);
and UO_1374 (O_1374,N_8152,N_8179);
and UO_1375 (O_1375,N_8276,N_8851);
or UO_1376 (O_1376,N_9481,N_7571);
nor UO_1377 (O_1377,N_9367,N_8192);
nor UO_1378 (O_1378,N_8155,N_9890);
or UO_1379 (O_1379,N_8773,N_8520);
and UO_1380 (O_1380,N_8012,N_7648);
and UO_1381 (O_1381,N_8305,N_9967);
nor UO_1382 (O_1382,N_9423,N_8997);
or UO_1383 (O_1383,N_8619,N_8615);
and UO_1384 (O_1384,N_9301,N_9448);
nor UO_1385 (O_1385,N_9692,N_8824);
and UO_1386 (O_1386,N_8999,N_7506);
or UO_1387 (O_1387,N_9967,N_9840);
nor UO_1388 (O_1388,N_9239,N_9883);
or UO_1389 (O_1389,N_9384,N_9416);
or UO_1390 (O_1390,N_8883,N_8756);
nor UO_1391 (O_1391,N_9030,N_8998);
or UO_1392 (O_1392,N_8470,N_9668);
or UO_1393 (O_1393,N_7619,N_8899);
and UO_1394 (O_1394,N_7599,N_8576);
nor UO_1395 (O_1395,N_8350,N_7712);
nand UO_1396 (O_1396,N_8441,N_9540);
or UO_1397 (O_1397,N_9662,N_8870);
or UO_1398 (O_1398,N_9473,N_9250);
nor UO_1399 (O_1399,N_8704,N_8253);
or UO_1400 (O_1400,N_9225,N_9274);
nor UO_1401 (O_1401,N_7512,N_8966);
xor UO_1402 (O_1402,N_8175,N_9229);
and UO_1403 (O_1403,N_7675,N_9675);
nand UO_1404 (O_1404,N_8088,N_9688);
xnor UO_1405 (O_1405,N_9689,N_8857);
or UO_1406 (O_1406,N_7524,N_7784);
and UO_1407 (O_1407,N_8709,N_9377);
nand UO_1408 (O_1408,N_7577,N_7862);
nand UO_1409 (O_1409,N_7619,N_8347);
nor UO_1410 (O_1410,N_9121,N_7865);
and UO_1411 (O_1411,N_7840,N_8367);
nand UO_1412 (O_1412,N_7951,N_9157);
and UO_1413 (O_1413,N_8331,N_9602);
and UO_1414 (O_1414,N_9173,N_9202);
nand UO_1415 (O_1415,N_9766,N_7776);
or UO_1416 (O_1416,N_7793,N_9420);
nand UO_1417 (O_1417,N_9959,N_7580);
nand UO_1418 (O_1418,N_9059,N_7555);
nand UO_1419 (O_1419,N_8869,N_8806);
and UO_1420 (O_1420,N_7988,N_8361);
and UO_1421 (O_1421,N_8838,N_7957);
nor UO_1422 (O_1422,N_8815,N_9333);
or UO_1423 (O_1423,N_8086,N_9877);
and UO_1424 (O_1424,N_8480,N_9238);
nor UO_1425 (O_1425,N_9591,N_9502);
nand UO_1426 (O_1426,N_7770,N_8259);
nor UO_1427 (O_1427,N_9275,N_9041);
and UO_1428 (O_1428,N_8573,N_9248);
nor UO_1429 (O_1429,N_8472,N_9120);
or UO_1430 (O_1430,N_8812,N_9487);
or UO_1431 (O_1431,N_8449,N_7796);
or UO_1432 (O_1432,N_7529,N_9781);
xnor UO_1433 (O_1433,N_9426,N_9260);
and UO_1434 (O_1434,N_8201,N_9403);
nor UO_1435 (O_1435,N_9451,N_9099);
or UO_1436 (O_1436,N_8620,N_7985);
nor UO_1437 (O_1437,N_7897,N_8920);
or UO_1438 (O_1438,N_9880,N_8543);
or UO_1439 (O_1439,N_8472,N_8855);
and UO_1440 (O_1440,N_8357,N_8945);
or UO_1441 (O_1441,N_8815,N_7796);
and UO_1442 (O_1442,N_8920,N_8295);
and UO_1443 (O_1443,N_9951,N_7813);
nand UO_1444 (O_1444,N_7880,N_8018);
or UO_1445 (O_1445,N_8200,N_7964);
or UO_1446 (O_1446,N_9823,N_8945);
and UO_1447 (O_1447,N_8049,N_8548);
nand UO_1448 (O_1448,N_9845,N_7511);
nor UO_1449 (O_1449,N_8737,N_7642);
and UO_1450 (O_1450,N_7910,N_9759);
nand UO_1451 (O_1451,N_9650,N_8655);
nand UO_1452 (O_1452,N_8037,N_9237);
and UO_1453 (O_1453,N_7777,N_7875);
nand UO_1454 (O_1454,N_8565,N_7891);
nor UO_1455 (O_1455,N_9453,N_9276);
nor UO_1456 (O_1456,N_9483,N_8157);
nor UO_1457 (O_1457,N_9449,N_8262);
nand UO_1458 (O_1458,N_8980,N_9221);
nand UO_1459 (O_1459,N_9964,N_9931);
nor UO_1460 (O_1460,N_7791,N_9649);
nand UO_1461 (O_1461,N_8880,N_9324);
or UO_1462 (O_1462,N_9996,N_8899);
and UO_1463 (O_1463,N_8081,N_9787);
nand UO_1464 (O_1464,N_8716,N_7685);
nand UO_1465 (O_1465,N_9683,N_9877);
nor UO_1466 (O_1466,N_9656,N_7706);
or UO_1467 (O_1467,N_9766,N_8725);
xor UO_1468 (O_1468,N_8108,N_8138);
nand UO_1469 (O_1469,N_8257,N_8839);
or UO_1470 (O_1470,N_7922,N_8974);
and UO_1471 (O_1471,N_9488,N_9503);
nor UO_1472 (O_1472,N_9047,N_8259);
or UO_1473 (O_1473,N_8879,N_8327);
and UO_1474 (O_1474,N_9785,N_8515);
and UO_1475 (O_1475,N_8404,N_8070);
xnor UO_1476 (O_1476,N_7987,N_8128);
nor UO_1477 (O_1477,N_8838,N_7501);
or UO_1478 (O_1478,N_7929,N_8285);
or UO_1479 (O_1479,N_9645,N_8950);
nand UO_1480 (O_1480,N_9273,N_9681);
nor UO_1481 (O_1481,N_8720,N_9841);
nor UO_1482 (O_1482,N_9076,N_8343);
or UO_1483 (O_1483,N_8417,N_7742);
and UO_1484 (O_1484,N_8133,N_7941);
and UO_1485 (O_1485,N_8418,N_8147);
nor UO_1486 (O_1486,N_9922,N_8486);
nand UO_1487 (O_1487,N_8550,N_9279);
or UO_1488 (O_1488,N_9270,N_9261);
nand UO_1489 (O_1489,N_7732,N_7968);
and UO_1490 (O_1490,N_8236,N_8084);
nor UO_1491 (O_1491,N_9674,N_7963);
and UO_1492 (O_1492,N_7578,N_8978);
and UO_1493 (O_1493,N_9414,N_8929);
nand UO_1494 (O_1494,N_9106,N_9585);
and UO_1495 (O_1495,N_8377,N_9591);
and UO_1496 (O_1496,N_9615,N_8705);
nand UO_1497 (O_1497,N_8372,N_8027);
nor UO_1498 (O_1498,N_7636,N_8351);
and UO_1499 (O_1499,N_8008,N_7773);
endmodule