module basic_1000_10000_1500_4_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_709,In_120);
nor U1 (N_1,In_876,In_721);
nor U2 (N_2,In_112,In_40);
and U3 (N_3,In_740,In_691);
nand U4 (N_4,In_355,In_164);
nand U5 (N_5,In_555,In_698);
and U6 (N_6,In_574,In_313);
or U7 (N_7,In_783,In_339);
xnor U8 (N_8,In_485,In_602);
nor U9 (N_9,In_174,In_294);
nand U10 (N_10,In_639,In_128);
nand U11 (N_11,In_391,In_357);
nand U12 (N_12,In_542,In_860);
nor U13 (N_13,In_205,In_605);
or U14 (N_14,In_63,In_118);
or U15 (N_15,In_182,In_848);
or U16 (N_16,In_929,In_233);
nor U17 (N_17,In_133,In_809);
and U18 (N_18,In_351,In_912);
nor U19 (N_19,In_749,In_955);
nand U20 (N_20,In_445,In_841);
nor U21 (N_21,In_27,In_416);
or U22 (N_22,In_972,In_75);
nor U23 (N_23,In_96,In_773);
xnor U24 (N_24,In_79,In_948);
and U25 (N_25,In_41,In_380);
xnor U26 (N_26,In_735,In_633);
or U27 (N_27,In_431,In_314);
xnor U28 (N_28,In_386,In_882);
xnor U29 (N_29,In_76,In_219);
nor U30 (N_30,In_812,In_757);
nor U31 (N_31,In_413,In_614);
nor U32 (N_32,In_80,In_449);
or U33 (N_33,In_301,In_251);
nand U34 (N_34,In_651,In_402);
and U35 (N_35,In_708,In_221);
or U36 (N_36,In_341,In_212);
nor U37 (N_37,In_702,In_608);
and U38 (N_38,In_305,In_694);
or U39 (N_39,In_423,In_31);
and U40 (N_40,In_454,In_42);
xor U41 (N_41,In_477,In_778);
and U42 (N_42,In_218,In_310);
nor U43 (N_43,In_422,In_887);
or U44 (N_44,In_201,In_412);
or U45 (N_45,In_178,In_784);
and U46 (N_46,In_629,In_269);
and U47 (N_47,In_25,In_901);
xor U48 (N_48,In_279,In_909);
nor U49 (N_49,In_267,In_469);
and U50 (N_50,In_820,In_532);
nor U51 (N_51,In_681,In_607);
or U52 (N_52,In_932,In_177);
nand U53 (N_53,In_468,In_870);
nor U54 (N_54,In_747,In_951);
and U55 (N_55,In_987,In_793);
xnor U56 (N_56,In_985,In_452);
or U57 (N_57,In_828,In_894);
and U58 (N_58,In_840,In_395);
nand U59 (N_59,In_968,In_459);
nor U60 (N_60,In_624,In_154);
or U61 (N_61,In_22,In_800);
and U62 (N_62,In_97,In_687);
and U63 (N_63,In_915,In_361);
nand U64 (N_64,In_601,In_831);
nor U65 (N_65,In_609,In_216);
or U66 (N_66,In_737,In_879);
xnor U67 (N_67,In_679,In_705);
nor U68 (N_68,In_969,In_772);
nor U69 (N_69,In_561,In_530);
and U70 (N_70,In_883,In_817);
or U71 (N_71,In_913,In_648);
nor U72 (N_72,In_170,In_275);
nand U73 (N_73,In_329,In_388);
nor U74 (N_74,In_807,In_898);
nand U75 (N_75,In_464,In_796);
nand U76 (N_76,In_842,In_242);
nor U77 (N_77,In_563,In_964);
nor U78 (N_78,In_718,In_751);
or U79 (N_79,In_936,In_787);
nor U80 (N_80,In_662,In_891);
nor U81 (N_81,In_845,In_488);
nand U82 (N_82,In_917,In_153);
nor U83 (N_83,In_239,In_546);
nand U84 (N_84,In_768,In_222);
or U85 (N_85,In_824,In_761);
nand U86 (N_86,In_653,In_760);
xnor U87 (N_87,In_973,In_382);
and U88 (N_88,In_764,In_295);
nand U89 (N_89,In_179,In_387);
or U90 (N_90,In_461,In_880);
nand U91 (N_91,In_712,In_259);
nor U92 (N_92,In_20,In_957);
nor U93 (N_93,In_213,In_754);
xor U94 (N_94,In_980,In_701);
nor U95 (N_95,In_52,In_849);
nand U96 (N_96,In_881,In_660);
nor U97 (N_97,In_515,In_941);
and U98 (N_98,In_473,In_258);
or U99 (N_99,In_87,In_302);
nor U100 (N_100,In_244,In_846);
and U101 (N_101,In_372,In_874);
and U102 (N_102,In_720,In_405);
and U103 (N_103,In_224,In_308);
and U104 (N_104,In_204,In_30);
xnor U105 (N_105,In_726,In_229);
and U106 (N_106,In_743,In_871);
and U107 (N_107,In_211,In_11);
nor U108 (N_108,In_537,In_695);
nand U109 (N_109,In_186,In_151);
nor U110 (N_110,In_113,In_180);
nor U111 (N_111,In_441,In_270);
nor U112 (N_112,In_952,In_136);
or U113 (N_113,In_669,In_167);
or U114 (N_114,In_495,In_419);
xor U115 (N_115,In_283,In_524);
and U116 (N_116,In_160,In_13);
nor U117 (N_117,In_374,In_114);
nor U118 (N_118,In_19,In_700);
and U119 (N_119,In_24,In_309);
and U120 (N_120,In_611,In_489);
nor U121 (N_121,In_794,In_818);
nor U122 (N_122,In_480,In_577);
nand U123 (N_123,In_869,In_215);
or U124 (N_124,In_710,In_939);
nand U125 (N_125,In_398,In_82);
nor U126 (N_126,In_2,In_644);
nand U127 (N_127,In_396,In_837);
or U128 (N_128,In_707,In_947);
nand U129 (N_129,In_665,In_248);
nand U130 (N_130,In_714,In_271);
nand U131 (N_131,In_364,In_130);
nand U132 (N_132,In_4,In_910);
or U133 (N_133,In_435,In_976);
nand U134 (N_134,In_919,In_203);
nand U135 (N_135,In_826,In_630);
nor U136 (N_136,In_35,In_392);
nor U137 (N_137,In_241,In_632);
or U138 (N_138,In_425,In_847);
and U139 (N_139,In_297,In_795);
or U140 (N_140,In_496,In_432);
nor U141 (N_141,In_78,In_621);
xor U142 (N_142,In_394,In_750);
nand U143 (N_143,In_210,In_942);
or U144 (N_144,In_744,In_690);
nor U145 (N_145,In_979,In_507);
or U146 (N_146,In_428,In_474);
nand U147 (N_147,In_767,In_81);
nand U148 (N_148,In_706,In_988);
nor U149 (N_149,In_326,In_805);
nor U150 (N_150,In_619,In_777);
nor U151 (N_151,In_821,In_86);
or U152 (N_152,In_554,In_265);
and U153 (N_153,In_672,In_786);
or U154 (N_154,In_885,In_646);
or U155 (N_155,In_978,In_526);
nand U156 (N_156,In_616,In_360);
and U157 (N_157,In_453,In_763);
nand U158 (N_158,In_873,In_29);
or U159 (N_159,In_322,In_333);
nor U160 (N_160,In_12,In_667);
nor U161 (N_161,In_791,In_755);
nor U162 (N_162,In_933,In_200);
xor U163 (N_163,In_433,In_728);
or U164 (N_164,In_59,In_567);
nor U165 (N_165,In_816,In_799);
nand U166 (N_166,In_383,In_491);
and U167 (N_167,In_552,In_553);
or U168 (N_168,In_520,In_102);
and U169 (N_169,In_770,In_187);
and U170 (N_170,In_243,In_264);
nor U171 (N_171,In_73,In_946);
nand U172 (N_172,In_358,In_106);
nor U173 (N_173,In_534,In_850);
xor U174 (N_174,In_490,In_483);
nor U175 (N_175,In_995,In_634);
nor U176 (N_176,In_45,In_176);
and U177 (N_177,In_253,In_370);
nand U178 (N_178,In_17,In_580);
nor U179 (N_179,In_977,In_606);
nand U180 (N_180,In_37,In_103);
nor U181 (N_181,In_467,In_911);
and U182 (N_182,In_108,In_74);
or U183 (N_183,In_658,In_522);
nand U184 (N_184,In_782,In_171);
and U185 (N_185,In_509,In_195);
or U186 (N_186,In_974,In_654);
nor U187 (N_187,In_332,In_337);
or U188 (N_188,In_47,In_642);
or U189 (N_189,In_217,In_647);
nor U190 (N_190,In_6,In_323);
xnor U191 (N_191,In_199,In_833);
or U192 (N_192,In_442,In_236);
and U193 (N_193,In_115,In_902);
nor U194 (N_194,In_207,In_157);
xnor U195 (N_195,In_727,In_142);
and U196 (N_196,In_588,In_385);
or U197 (N_197,In_722,In_330);
nor U198 (N_198,In_231,In_125);
nand U199 (N_199,In_937,In_684);
and U200 (N_200,In_126,In_196);
nand U201 (N_201,In_247,In_797);
nand U202 (N_202,In_677,In_328);
or U203 (N_203,In_839,In_280);
nor U204 (N_204,In_688,In_255);
nand U205 (N_205,In_521,In_340);
xnor U206 (N_206,In_462,In_792);
nor U207 (N_207,In_299,In_94);
and U208 (N_208,In_140,In_100);
xor U209 (N_209,In_945,In_890);
or U210 (N_210,In_905,In_149);
nor U211 (N_211,In_692,In_685);
or U212 (N_212,In_771,In_225);
nand U213 (N_213,In_220,In_877);
nand U214 (N_214,In_502,In_935);
and U215 (N_215,In_717,In_752);
nand U216 (N_216,In_581,In_626);
or U217 (N_217,In_723,In_146);
nor U218 (N_218,In_830,In_859);
and U219 (N_219,In_316,In_408);
or U220 (N_220,In_209,In_730);
and U221 (N_221,In_900,In_535);
nor U222 (N_222,In_926,In_732);
and U223 (N_223,In_371,In_557);
nand U224 (N_224,In_482,In_921);
or U225 (N_225,In_739,In_513);
nand U226 (N_226,In_741,In_774);
xor U227 (N_227,In_888,In_536);
or U228 (N_228,In_158,In_368);
nor U229 (N_229,In_77,In_682);
nor U230 (N_230,In_811,In_612);
xor U231 (N_231,In_815,In_121);
xor U232 (N_232,In_983,In_861);
nor U233 (N_233,In_625,In_344);
or U234 (N_234,In_237,In_298);
nand U235 (N_235,In_585,In_352);
or U236 (N_236,In_202,In_623);
nand U237 (N_237,In_208,In_291);
nand U238 (N_238,In_367,In_517);
nor U239 (N_239,In_188,In_533);
xnor U240 (N_240,In_998,In_345);
and U241 (N_241,In_172,In_938);
nor U242 (N_242,In_856,In_960);
and U243 (N_243,In_834,In_285);
nand U244 (N_244,In_397,In_430);
nor U245 (N_245,In_904,In_274);
or U246 (N_246,In_595,In_953);
nand U247 (N_247,In_853,In_33);
or U248 (N_248,In_982,In_70);
nand U249 (N_249,In_348,In_814);
and U250 (N_250,In_362,In_753);
nor U251 (N_251,In_956,In_16);
and U252 (N_252,In_117,In_583);
and U253 (N_253,In_928,In_104);
nand U254 (N_254,In_862,In_0);
nor U255 (N_255,In_363,In_227);
and U256 (N_256,In_756,In_666);
and U257 (N_257,In_966,In_373);
xnor U258 (N_258,In_599,In_852);
or U259 (N_259,In_779,In_250);
nor U260 (N_260,In_661,In_197);
xor U261 (N_261,In_384,In_131);
nor U262 (N_262,In_994,In_23);
nand U263 (N_263,In_393,In_48);
nand U264 (N_264,In_159,In_109);
or U265 (N_265,In_970,In_541);
xor U266 (N_266,In_50,In_716);
or U267 (N_267,In_127,In_389);
and U268 (N_268,In_66,In_965);
nor U269 (N_269,In_864,In_465);
nand U270 (N_270,In_822,In_895);
nor U271 (N_271,In_353,In_311);
nand U272 (N_272,In_290,In_906);
nand U273 (N_273,In_137,In_404);
or U274 (N_274,In_827,In_317);
and U275 (N_275,In_668,In_663);
and U276 (N_276,In_451,In_84);
nand U277 (N_277,In_868,In_808);
or U278 (N_278,In_282,In_892);
nand U279 (N_279,In_576,In_284);
and U280 (N_280,In_855,In_235);
or U281 (N_281,In_578,In_414);
nand U282 (N_282,In_922,In_107);
nand U283 (N_283,In_379,In_95);
nor U284 (N_284,In_443,In_369);
or U285 (N_285,In_503,In_803);
nand U286 (N_286,In_518,In_736);
xnor U287 (N_287,In_145,In_494);
nand U288 (N_288,In_155,In_99);
nand U289 (N_289,In_303,In_993);
nand U290 (N_290,In_68,In_587);
nand U291 (N_291,In_657,In_189);
nor U292 (N_292,In_636,In_631);
or U293 (N_293,In_234,In_460);
nor U294 (N_294,In_168,In_276);
and U295 (N_295,In_996,In_409);
or U296 (N_296,In_55,In_49);
nor U297 (N_297,In_643,In_613);
or U298 (N_298,In_69,In_628);
or U299 (N_299,In_439,In_65);
and U300 (N_300,In_548,In_867);
nand U301 (N_301,In_598,In_637);
nor U302 (N_302,In_296,In_32);
and U303 (N_303,In_72,In_139);
and U304 (N_304,In_46,In_872);
or U305 (N_305,In_927,In_600);
and U306 (N_306,In_266,In_181);
nor U307 (N_307,In_105,In_418);
or U308 (N_308,In_999,In_547);
or U309 (N_309,In_427,In_544);
and U310 (N_310,In_278,In_954);
and U311 (N_311,In_659,In_436);
nor U312 (N_312,In_450,In_590);
xnor U313 (N_313,In_725,In_897);
nor U314 (N_314,In_246,In_748);
xnor U315 (N_315,In_514,In_759);
nor U316 (N_316,In_958,In_406);
or U317 (N_317,In_731,In_620);
or U318 (N_318,In_62,In_949);
xnor U319 (N_319,In_689,In_531);
or U320 (N_320,In_375,In_110);
nor U321 (N_321,In_7,In_60);
and U322 (N_322,In_479,In_655);
and U323 (N_323,In_836,In_124);
and U324 (N_324,In_724,In_400);
or U325 (N_325,In_504,In_981);
or U326 (N_326,In_615,In_734);
or U327 (N_327,In_914,In_429);
nor U328 (N_328,In_318,In_597);
xnor U329 (N_329,In_641,In_390);
xor U330 (N_330,In_696,In_550);
nor U331 (N_331,In_132,In_43);
or U332 (N_332,In_505,In_604);
nor U333 (N_333,In_893,In_147);
nor U334 (N_334,In_71,In_683);
nand U335 (N_335,In_312,In_699);
nand U336 (N_336,In_523,In_338);
xor U337 (N_337,In_463,In_471);
nor U338 (N_338,In_572,In_582);
nand U339 (N_339,In_539,In_458);
and U340 (N_340,In_889,In_93);
nand U341 (N_341,In_420,In_674);
nor U342 (N_342,In_569,In_512);
and U343 (N_343,In_769,In_790);
nand U344 (N_344,In_519,In_798);
nor U345 (N_345,In_67,In_448);
nand U346 (N_346,In_802,In_959);
and U347 (N_347,In_378,In_281);
nor U348 (N_348,In_963,In_528);
nand U349 (N_349,In_780,In_697);
or U350 (N_350,In_226,In_693);
or U351 (N_351,In_650,In_950);
nand U352 (N_352,In_486,In_971);
nor U353 (N_353,In_766,In_56);
xnor U354 (N_354,In_729,In_719);
and U355 (N_355,In_781,In_670);
and U356 (N_356,In_162,In_560);
or U357 (N_357,In_549,In_975);
and U358 (N_358,In_635,In_884);
or U359 (N_359,In_543,In_123);
nor U360 (N_360,In_262,In_315);
and U361 (N_361,In_129,In_343);
or U362 (N_362,In_711,In_51);
or U363 (N_363,In_579,In_410);
or U364 (N_364,In_596,In_161);
nor U365 (N_365,In_472,In_516);
and U366 (N_366,In_350,In_58);
or U367 (N_367,In_556,In_14);
xor U368 (N_368,In_943,In_335);
and U369 (N_369,In_381,In_64);
nand U370 (N_370,In_788,In_306);
nor U371 (N_371,In_497,In_854);
and U372 (N_372,In_640,In_589);
nor U373 (N_373,In_18,In_26);
and U374 (N_374,In_875,In_810);
and U375 (N_375,In_704,In_1);
nand U376 (N_376,In_575,In_678);
and U377 (N_377,In_785,In_789);
nor U378 (N_378,In_365,In_499);
and U379 (N_379,In_85,In_342);
nand U380 (N_380,In_347,In_143);
xor U381 (N_381,In_832,In_961);
and U382 (N_382,In_627,In_475);
and U383 (N_383,In_254,In_823);
nor U384 (N_384,In_622,In_566);
nor U385 (N_385,In_907,In_36);
nand U386 (N_386,In_9,In_366);
xnor U387 (N_387,In_508,In_715);
and U388 (N_388,In_111,In_134);
nor U389 (N_389,In_593,In_119);
or U390 (N_390,In_165,In_421);
nand U391 (N_391,In_256,In_903);
xor U392 (N_392,In_562,In_991);
and U393 (N_393,In_440,In_289);
and U394 (N_394,In_183,In_745);
and U395 (N_395,In_878,In_138);
and U396 (N_396,In_481,In_173);
nor U397 (N_397,In_407,In_263);
nor U398 (N_398,In_122,In_559);
nand U399 (N_399,In_38,In_565);
or U400 (N_400,In_804,In_493);
or U401 (N_401,In_232,In_500);
nor U402 (N_402,In_934,In_962);
nor U403 (N_403,In_260,In_967);
nand U404 (N_404,In_349,In_101);
nand U405 (N_405,In_510,In_238);
nor U406 (N_406,In_286,In_838);
nand U407 (N_407,In_617,In_277);
nand U408 (N_408,In_775,In_156);
and U409 (N_409,In_190,In_835);
xor U410 (N_410,In_652,In_300);
and U411 (N_411,In_758,In_98);
and U412 (N_412,In_571,In_568);
nand U413 (N_413,In_192,In_272);
nor U414 (N_414,In_34,In_455);
or U415 (N_415,In_252,In_478);
or U416 (N_416,In_415,In_813);
and U417 (N_417,In_135,In_899);
nor U418 (N_418,In_851,In_664);
xor U419 (N_419,In_551,In_470);
and U420 (N_420,In_83,In_527);
nand U421 (N_421,In_584,In_399);
and U422 (N_422,In_829,In_148);
or U423 (N_423,In_356,In_986);
and U424 (N_424,In_920,In_90);
nand U425 (N_425,In_206,In_924);
nand U426 (N_426,In_377,In_434);
or U427 (N_427,In_564,In_733);
nand U428 (N_428,In_586,In_857);
or U429 (N_429,In_484,In_39);
nor U430 (N_430,In_908,In_447);
or U431 (N_431,In_525,In_287);
and U432 (N_432,In_765,In_538);
xnor U433 (N_433,In_886,In_594);
or U434 (N_434,In_511,In_91);
and U435 (N_435,In_673,In_931);
nand U436 (N_436,In_191,In_558);
nor U437 (N_437,In_150,In_417);
nor U438 (N_438,In_675,In_742);
nor U439 (N_439,In_3,In_603);
nor U440 (N_440,In_334,In_863);
nand U441 (N_441,In_175,In_918);
or U442 (N_442,In_437,In_680);
or U443 (N_443,In_61,In_166);
or U444 (N_444,In_319,In_257);
or U445 (N_445,In_249,In_293);
xor U446 (N_446,In_656,In_610);
or U447 (N_447,In_529,In_498);
and U448 (N_448,In_476,In_738);
and U449 (N_449,In_354,In_424);
nor U450 (N_450,In_843,In_426);
nand U451 (N_451,In_865,In_776);
nor U452 (N_452,In_268,In_806);
xor U453 (N_453,In_292,In_185);
nor U454 (N_454,In_866,In_230);
or U455 (N_455,In_506,In_746);
nor U456 (N_456,In_618,In_573);
and U457 (N_457,In_858,In_261);
or U458 (N_458,In_703,In_194);
nand U459 (N_459,In_403,In_944);
nand U460 (N_460,In_336,In_8);
or U461 (N_461,In_327,In_819);
nand U462 (N_462,In_193,In_44);
xnor U463 (N_463,In_15,In_116);
xnor U464 (N_464,In_5,In_671);
nor U465 (N_465,In_169,In_545);
or U466 (N_466,In_916,In_92);
xnor U467 (N_467,In_456,In_321);
and U468 (N_468,In_89,In_989);
nand U469 (N_469,In_638,In_141);
nand U470 (N_470,In_346,In_88);
and U471 (N_471,In_649,In_446);
and U472 (N_472,In_940,In_28);
or U473 (N_473,In_240,In_487);
or U474 (N_474,In_645,In_54);
nor U475 (N_475,In_307,In_444);
nand U476 (N_476,In_144,In_457);
xnor U477 (N_477,In_925,In_896);
nand U478 (N_478,In_501,In_492);
and U479 (N_479,In_990,In_401);
xnor U480 (N_480,In_801,In_184);
or U481 (N_481,In_570,In_10);
nand U482 (N_482,In_825,In_288);
nor U483 (N_483,In_228,In_466);
and U484 (N_484,In_676,In_214);
nand U485 (N_485,In_320,In_844);
or U486 (N_486,In_762,In_163);
or U487 (N_487,In_592,In_53);
or U488 (N_488,In_325,In_930);
nand U489 (N_489,In_359,In_331);
nor U490 (N_490,In_997,In_57);
and U491 (N_491,In_540,In_152);
xor U492 (N_492,In_273,In_223);
and U493 (N_493,In_923,In_21);
nand U494 (N_494,In_376,In_984);
and U495 (N_495,In_324,In_713);
nor U496 (N_496,In_438,In_591);
and U497 (N_497,In_992,In_304);
nand U498 (N_498,In_686,In_198);
and U499 (N_499,In_245,In_411);
and U500 (N_500,In_543,In_669);
or U501 (N_501,In_77,In_499);
nor U502 (N_502,In_448,In_733);
and U503 (N_503,In_316,In_361);
or U504 (N_504,In_446,In_70);
xor U505 (N_505,In_743,In_694);
or U506 (N_506,In_275,In_898);
or U507 (N_507,In_606,In_813);
xor U508 (N_508,In_44,In_676);
nor U509 (N_509,In_903,In_948);
and U510 (N_510,In_92,In_176);
nor U511 (N_511,In_424,In_945);
or U512 (N_512,In_888,In_794);
xnor U513 (N_513,In_354,In_289);
nor U514 (N_514,In_930,In_168);
and U515 (N_515,In_810,In_462);
nor U516 (N_516,In_204,In_450);
and U517 (N_517,In_222,In_576);
or U518 (N_518,In_324,In_311);
or U519 (N_519,In_440,In_877);
or U520 (N_520,In_795,In_590);
and U521 (N_521,In_242,In_734);
nor U522 (N_522,In_293,In_170);
nor U523 (N_523,In_645,In_843);
nand U524 (N_524,In_563,In_305);
xnor U525 (N_525,In_175,In_683);
xor U526 (N_526,In_394,In_731);
nand U527 (N_527,In_784,In_760);
or U528 (N_528,In_152,In_143);
nand U529 (N_529,In_600,In_755);
and U530 (N_530,In_866,In_632);
and U531 (N_531,In_620,In_257);
xnor U532 (N_532,In_95,In_247);
nand U533 (N_533,In_563,In_25);
or U534 (N_534,In_308,In_460);
and U535 (N_535,In_147,In_771);
nor U536 (N_536,In_765,In_951);
nor U537 (N_537,In_186,In_831);
or U538 (N_538,In_816,In_672);
nand U539 (N_539,In_965,In_557);
nor U540 (N_540,In_139,In_636);
and U541 (N_541,In_552,In_757);
nand U542 (N_542,In_120,In_953);
nor U543 (N_543,In_530,In_899);
nor U544 (N_544,In_390,In_158);
nand U545 (N_545,In_490,In_12);
nor U546 (N_546,In_556,In_853);
nor U547 (N_547,In_574,In_116);
or U548 (N_548,In_802,In_82);
nand U549 (N_549,In_468,In_905);
or U550 (N_550,In_399,In_632);
or U551 (N_551,In_919,In_552);
and U552 (N_552,In_193,In_890);
nor U553 (N_553,In_21,In_196);
and U554 (N_554,In_288,In_293);
nand U555 (N_555,In_52,In_67);
and U556 (N_556,In_863,In_933);
nor U557 (N_557,In_224,In_718);
nor U558 (N_558,In_684,In_310);
or U559 (N_559,In_864,In_296);
xor U560 (N_560,In_581,In_848);
or U561 (N_561,In_620,In_853);
nor U562 (N_562,In_982,In_906);
xor U563 (N_563,In_773,In_64);
nand U564 (N_564,In_992,In_702);
xor U565 (N_565,In_953,In_629);
or U566 (N_566,In_920,In_485);
or U567 (N_567,In_780,In_289);
nor U568 (N_568,In_249,In_318);
nor U569 (N_569,In_752,In_36);
nand U570 (N_570,In_293,In_552);
xor U571 (N_571,In_306,In_964);
nor U572 (N_572,In_549,In_302);
and U573 (N_573,In_466,In_134);
nand U574 (N_574,In_380,In_831);
xnor U575 (N_575,In_221,In_414);
or U576 (N_576,In_20,In_721);
nor U577 (N_577,In_843,In_477);
nand U578 (N_578,In_923,In_809);
or U579 (N_579,In_492,In_203);
nand U580 (N_580,In_954,In_86);
xor U581 (N_581,In_99,In_83);
or U582 (N_582,In_112,In_287);
or U583 (N_583,In_360,In_335);
and U584 (N_584,In_751,In_120);
nand U585 (N_585,In_936,In_418);
nor U586 (N_586,In_7,In_45);
or U587 (N_587,In_587,In_598);
nor U588 (N_588,In_858,In_180);
or U589 (N_589,In_327,In_655);
or U590 (N_590,In_153,In_660);
nor U591 (N_591,In_586,In_906);
nor U592 (N_592,In_713,In_480);
xnor U593 (N_593,In_924,In_328);
nand U594 (N_594,In_951,In_637);
and U595 (N_595,In_378,In_519);
and U596 (N_596,In_405,In_986);
nand U597 (N_597,In_83,In_260);
or U598 (N_598,In_570,In_187);
and U599 (N_599,In_710,In_706);
nor U600 (N_600,In_436,In_913);
or U601 (N_601,In_31,In_825);
or U602 (N_602,In_620,In_135);
nand U603 (N_603,In_764,In_824);
and U604 (N_604,In_902,In_425);
nor U605 (N_605,In_581,In_304);
nand U606 (N_606,In_113,In_576);
nor U607 (N_607,In_196,In_606);
nor U608 (N_608,In_914,In_312);
xnor U609 (N_609,In_347,In_634);
nand U610 (N_610,In_632,In_747);
or U611 (N_611,In_292,In_49);
nand U612 (N_612,In_515,In_63);
nand U613 (N_613,In_513,In_393);
nor U614 (N_614,In_313,In_227);
xor U615 (N_615,In_317,In_669);
or U616 (N_616,In_715,In_491);
and U617 (N_617,In_807,In_746);
or U618 (N_618,In_993,In_72);
or U619 (N_619,In_668,In_300);
and U620 (N_620,In_482,In_802);
nand U621 (N_621,In_909,In_33);
xor U622 (N_622,In_755,In_458);
nor U623 (N_623,In_258,In_247);
and U624 (N_624,In_738,In_426);
or U625 (N_625,In_861,In_995);
nand U626 (N_626,In_856,In_240);
xor U627 (N_627,In_946,In_277);
nor U628 (N_628,In_176,In_26);
nand U629 (N_629,In_838,In_3);
nor U630 (N_630,In_459,In_756);
nand U631 (N_631,In_519,In_413);
nand U632 (N_632,In_674,In_783);
and U633 (N_633,In_346,In_216);
and U634 (N_634,In_138,In_200);
nor U635 (N_635,In_275,In_991);
nand U636 (N_636,In_814,In_126);
or U637 (N_637,In_32,In_587);
and U638 (N_638,In_9,In_343);
or U639 (N_639,In_527,In_376);
and U640 (N_640,In_558,In_982);
nor U641 (N_641,In_74,In_197);
and U642 (N_642,In_649,In_215);
or U643 (N_643,In_127,In_508);
xor U644 (N_644,In_934,In_856);
and U645 (N_645,In_140,In_447);
and U646 (N_646,In_526,In_869);
or U647 (N_647,In_413,In_491);
or U648 (N_648,In_650,In_680);
or U649 (N_649,In_163,In_546);
or U650 (N_650,In_685,In_856);
or U651 (N_651,In_611,In_931);
or U652 (N_652,In_567,In_299);
nand U653 (N_653,In_609,In_932);
nor U654 (N_654,In_792,In_922);
and U655 (N_655,In_127,In_992);
nor U656 (N_656,In_97,In_53);
or U657 (N_657,In_538,In_7);
nand U658 (N_658,In_202,In_203);
and U659 (N_659,In_187,In_243);
and U660 (N_660,In_428,In_110);
and U661 (N_661,In_533,In_114);
or U662 (N_662,In_832,In_881);
nor U663 (N_663,In_683,In_350);
nand U664 (N_664,In_408,In_389);
or U665 (N_665,In_193,In_34);
or U666 (N_666,In_469,In_43);
or U667 (N_667,In_856,In_492);
or U668 (N_668,In_584,In_122);
nor U669 (N_669,In_408,In_262);
nand U670 (N_670,In_653,In_413);
nand U671 (N_671,In_870,In_196);
nor U672 (N_672,In_284,In_39);
nand U673 (N_673,In_172,In_48);
and U674 (N_674,In_71,In_630);
nor U675 (N_675,In_727,In_390);
nor U676 (N_676,In_774,In_552);
nand U677 (N_677,In_906,In_214);
xor U678 (N_678,In_100,In_959);
nor U679 (N_679,In_114,In_717);
nand U680 (N_680,In_276,In_948);
and U681 (N_681,In_739,In_726);
nand U682 (N_682,In_638,In_852);
nand U683 (N_683,In_832,In_19);
and U684 (N_684,In_335,In_307);
or U685 (N_685,In_433,In_335);
or U686 (N_686,In_587,In_858);
nor U687 (N_687,In_502,In_91);
xnor U688 (N_688,In_888,In_582);
or U689 (N_689,In_126,In_110);
nand U690 (N_690,In_793,In_245);
or U691 (N_691,In_414,In_499);
nand U692 (N_692,In_783,In_190);
and U693 (N_693,In_951,In_532);
nor U694 (N_694,In_985,In_560);
nor U695 (N_695,In_943,In_796);
or U696 (N_696,In_289,In_742);
nand U697 (N_697,In_871,In_829);
or U698 (N_698,In_247,In_266);
nor U699 (N_699,In_59,In_164);
and U700 (N_700,In_124,In_20);
nor U701 (N_701,In_636,In_490);
nand U702 (N_702,In_465,In_582);
nand U703 (N_703,In_88,In_701);
or U704 (N_704,In_702,In_323);
and U705 (N_705,In_991,In_70);
or U706 (N_706,In_60,In_171);
or U707 (N_707,In_455,In_77);
and U708 (N_708,In_436,In_679);
or U709 (N_709,In_325,In_343);
nand U710 (N_710,In_706,In_908);
nor U711 (N_711,In_748,In_312);
and U712 (N_712,In_912,In_470);
nor U713 (N_713,In_135,In_709);
nor U714 (N_714,In_144,In_320);
nor U715 (N_715,In_404,In_739);
or U716 (N_716,In_453,In_846);
and U717 (N_717,In_423,In_854);
or U718 (N_718,In_420,In_226);
nand U719 (N_719,In_969,In_114);
nand U720 (N_720,In_925,In_241);
nor U721 (N_721,In_690,In_863);
nor U722 (N_722,In_115,In_180);
and U723 (N_723,In_631,In_448);
xnor U724 (N_724,In_242,In_968);
or U725 (N_725,In_256,In_538);
nor U726 (N_726,In_303,In_179);
and U727 (N_727,In_880,In_329);
and U728 (N_728,In_730,In_329);
and U729 (N_729,In_565,In_935);
or U730 (N_730,In_701,In_441);
and U731 (N_731,In_393,In_653);
nor U732 (N_732,In_365,In_427);
nor U733 (N_733,In_707,In_343);
nand U734 (N_734,In_73,In_834);
nand U735 (N_735,In_786,In_146);
nand U736 (N_736,In_796,In_470);
xnor U737 (N_737,In_554,In_673);
xnor U738 (N_738,In_740,In_151);
and U739 (N_739,In_700,In_272);
or U740 (N_740,In_19,In_907);
nor U741 (N_741,In_963,In_150);
and U742 (N_742,In_720,In_880);
nand U743 (N_743,In_316,In_533);
nor U744 (N_744,In_373,In_892);
nor U745 (N_745,In_50,In_668);
nor U746 (N_746,In_122,In_735);
xnor U747 (N_747,In_583,In_398);
xor U748 (N_748,In_311,In_601);
nor U749 (N_749,In_338,In_529);
nand U750 (N_750,In_593,In_976);
and U751 (N_751,In_957,In_151);
nand U752 (N_752,In_719,In_504);
and U753 (N_753,In_27,In_949);
nor U754 (N_754,In_200,In_116);
and U755 (N_755,In_829,In_118);
or U756 (N_756,In_647,In_613);
or U757 (N_757,In_816,In_198);
nor U758 (N_758,In_73,In_829);
nand U759 (N_759,In_890,In_473);
nand U760 (N_760,In_19,In_360);
and U761 (N_761,In_509,In_975);
xnor U762 (N_762,In_41,In_364);
xor U763 (N_763,In_850,In_727);
or U764 (N_764,In_531,In_167);
and U765 (N_765,In_74,In_802);
nand U766 (N_766,In_522,In_15);
nor U767 (N_767,In_552,In_792);
and U768 (N_768,In_845,In_180);
and U769 (N_769,In_106,In_948);
and U770 (N_770,In_20,In_269);
nand U771 (N_771,In_167,In_134);
or U772 (N_772,In_55,In_915);
and U773 (N_773,In_349,In_194);
nand U774 (N_774,In_924,In_795);
and U775 (N_775,In_54,In_777);
nand U776 (N_776,In_309,In_348);
and U777 (N_777,In_515,In_364);
xor U778 (N_778,In_68,In_723);
nand U779 (N_779,In_956,In_544);
nand U780 (N_780,In_493,In_953);
xnor U781 (N_781,In_100,In_900);
nand U782 (N_782,In_757,In_497);
or U783 (N_783,In_101,In_355);
nand U784 (N_784,In_85,In_364);
and U785 (N_785,In_413,In_155);
nor U786 (N_786,In_916,In_96);
nor U787 (N_787,In_962,In_6);
and U788 (N_788,In_46,In_409);
nand U789 (N_789,In_791,In_955);
or U790 (N_790,In_121,In_875);
and U791 (N_791,In_350,In_793);
nand U792 (N_792,In_201,In_982);
nor U793 (N_793,In_834,In_438);
and U794 (N_794,In_109,In_170);
nor U795 (N_795,In_666,In_361);
nor U796 (N_796,In_125,In_312);
and U797 (N_797,In_592,In_910);
nand U798 (N_798,In_444,In_361);
and U799 (N_799,In_573,In_643);
and U800 (N_800,In_414,In_451);
xnor U801 (N_801,In_696,In_688);
nand U802 (N_802,In_804,In_875);
nor U803 (N_803,In_187,In_634);
and U804 (N_804,In_348,In_810);
and U805 (N_805,In_751,In_666);
and U806 (N_806,In_421,In_792);
nor U807 (N_807,In_116,In_13);
nand U808 (N_808,In_66,In_582);
nor U809 (N_809,In_303,In_185);
nor U810 (N_810,In_660,In_411);
and U811 (N_811,In_739,In_758);
nand U812 (N_812,In_905,In_449);
nand U813 (N_813,In_589,In_59);
and U814 (N_814,In_819,In_178);
or U815 (N_815,In_103,In_118);
and U816 (N_816,In_518,In_981);
xor U817 (N_817,In_559,In_931);
or U818 (N_818,In_282,In_383);
and U819 (N_819,In_12,In_124);
nand U820 (N_820,In_696,In_597);
and U821 (N_821,In_49,In_363);
or U822 (N_822,In_150,In_304);
nand U823 (N_823,In_561,In_364);
nand U824 (N_824,In_884,In_986);
or U825 (N_825,In_208,In_262);
or U826 (N_826,In_758,In_28);
nand U827 (N_827,In_383,In_567);
and U828 (N_828,In_667,In_608);
nand U829 (N_829,In_177,In_955);
or U830 (N_830,In_871,In_519);
or U831 (N_831,In_532,In_356);
nand U832 (N_832,In_814,In_941);
nand U833 (N_833,In_343,In_190);
nand U834 (N_834,In_822,In_801);
nand U835 (N_835,In_478,In_434);
nand U836 (N_836,In_443,In_573);
nor U837 (N_837,In_908,In_766);
or U838 (N_838,In_625,In_174);
and U839 (N_839,In_460,In_267);
nor U840 (N_840,In_512,In_845);
and U841 (N_841,In_813,In_217);
xor U842 (N_842,In_410,In_497);
nand U843 (N_843,In_611,In_596);
nor U844 (N_844,In_304,In_26);
nor U845 (N_845,In_530,In_203);
or U846 (N_846,In_537,In_196);
and U847 (N_847,In_93,In_764);
or U848 (N_848,In_199,In_670);
nand U849 (N_849,In_444,In_127);
or U850 (N_850,In_801,In_29);
nor U851 (N_851,In_745,In_7);
nor U852 (N_852,In_701,In_629);
nand U853 (N_853,In_345,In_413);
or U854 (N_854,In_911,In_613);
nor U855 (N_855,In_125,In_126);
nor U856 (N_856,In_389,In_406);
nor U857 (N_857,In_185,In_342);
and U858 (N_858,In_313,In_499);
nand U859 (N_859,In_746,In_869);
nand U860 (N_860,In_224,In_90);
or U861 (N_861,In_564,In_574);
and U862 (N_862,In_328,In_983);
nand U863 (N_863,In_71,In_515);
or U864 (N_864,In_836,In_620);
and U865 (N_865,In_734,In_452);
nand U866 (N_866,In_90,In_499);
nand U867 (N_867,In_650,In_463);
nor U868 (N_868,In_132,In_141);
nor U869 (N_869,In_90,In_275);
or U870 (N_870,In_396,In_766);
nor U871 (N_871,In_992,In_980);
or U872 (N_872,In_718,In_1);
and U873 (N_873,In_198,In_733);
nor U874 (N_874,In_959,In_86);
or U875 (N_875,In_811,In_10);
nand U876 (N_876,In_615,In_159);
nor U877 (N_877,In_596,In_533);
or U878 (N_878,In_964,In_20);
and U879 (N_879,In_163,In_895);
and U880 (N_880,In_418,In_248);
and U881 (N_881,In_242,In_100);
nor U882 (N_882,In_639,In_922);
and U883 (N_883,In_646,In_596);
nor U884 (N_884,In_402,In_652);
nor U885 (N_885,In_938,In_866);
or U886 (N_886,In_198,In_807);
nor U887 (N_887,In_887,In_162);
nor U888 (N_888,In_15,In_311);
nand U889 (N_889,In_672,In_279);
nor U890 (N_890,In_146,In_13);
nor U891 (N_891,In_848,In_828);
xor U892 (N_892,In_623,In_920);
nor U893 (N_893,In_28,In_329);
and U894 (N_894,In_275,In_971);
and U895 (N_895,In_510,In_583);
or U896 (N_896,In_284,In_213);
nor U897 (N_897,In_474,In_398);
xor U898 (N_898,In_545,In_672);
or U899 (N_899,In_306,In_674);
and U900 (N_900,In_538,In_847);
xnor U901 (N_901,In_440,In_249);
nand U902 (N_902,In_893,In_499);
or U903 (N_903,In_648,In_748);
or U904 (N_904,In_958,In_117);
and U905 (N_905,In_760,In_151);
nand U906 (N_906,In_264,In_9);
or U907 (N_907,In_587,In_235);
nand U908 (N_908,In_231,In_67);
nand U909 (N_909,In_374,In_633);
or U910 (N_910,In_602,In_904);
and U911 (N_911,In_137,In_39);
nand U912 (N_912,In_183,In_288);
or U913 (N_913,In_48,In_326);
or U914 (N_914,In_303,In_175);
and U915 (N_915,In_319,In_18);
or U916 (N_916,In_578,In_217);
xnor U917 (N_917,In_887,In_333);
nor U918 (N_918,In_309,In_92);
nand U919 (N_919,In_404,In_978);
and U920 (N_920,In_640,In_506);
and U921 (N_921,In_476,In_73);
nor U922 (N_922,In_664,In_267);
and U923 (N_923,In_13,In_947);
or U924 (N_924,In_483,In_856);
nand U925 (N_925,In_622,In_375);
and U926 (N_926,In_285,In_242);
or U927 (N_927,In_457,In_757);
nand U928 (N_928,In_567,In_843);
or U929 (N_929,In_296,In_748);
nor U930 (N_930,In_194,In_718);
xor U931 (N_931,In_969,In_363);
and U932 (N_932,In_283,In_335);
or U933 (N_933,In_754,In_182);
nor U934 (N_934,In_818,In_609);
and U935 (N_935,In_670,In_447);
nor U936 (N_936,In_628,In_242);
and U937 (N_937,In_784,In_103);
or U938 (N_938,In_476,In_23);
nand U939 (N_939,In_230,In_737);
nor U940 (N_940,In_917,In_40);
and U941 (N_941,In_610,In_568);
nor U942 (N_942,In_686,In_195);
xnor U943 (N_943,In_8,In_402);
and U944 (N_944,In_170,In_188);
or U945 (N_945,In_227,In_420);
and U946 (N_946,In_778,In_269);
nand U947 (N_947,In_993,In_171);
or U948 (N_948,In_230,In_550);
xnor U949 (N_949,In_626,In_750);
and U950 (N_950,In_819,In_336);
nor U951 (N_951,In_563,In_699);
nor U952 (N_952,In_925,In_809);
and U953 (N_953,In_22,In_102);
nand U954 (N_954,In_564,In_306);
or U955 (N_955,In_66,In_869);
or U956 (N_956,In_397,In_194);
and U957 (N_957,In_525,In_500);
or U958 (N_958,In_351,In_52);
xnor U959 (N_959,In_486,In_704);
and U960 (N_960,In_921,In_376);
nor U961 (N_961,In_782,In_61);
nor U962 (N_962,In_541,In_566);
nor U963 (N_963,In_602,In_52);
and U964 (N_964,In_467,In_593);
xor U965 (N_965,In_773,In_537);
nand U966 (N_966,In_17,In_138);
nand U967 (N_967,In_452,In_713);
or U968 (N_968,In_601,In_898);
and U969 (N_969,In_195,In_894);
or U970 (N_970,In_219,In_228);
and U971 (N_971,In_176,In_524);
nor U972 (N_972,In_157,In_995);
and U973 (N_973,In_323,In_449);
or U974 (N_974,In_168,In_116);
or U975 (N_975,In_381,In_202);
and U976 (N_976,In_648,In_907);
nor U977 (N_977,In_621,In_200);
or U978 (N_978,In_922,In_365);
nand U979 (N_979,In_221,In_93);
nand U980 (N_980,In_143,In_198);
nor U981 (N_981,In_816,In_943);
nor U982 (N_982,In_206,In_744);
nand U983 (N_983,In_114,In_434);
nor U984 (N_984,In_514,In_116);
and U985 (N_985,In_599,In_395);
or U986 (N_986,In_886,In_45);
and U987 (N_987,In_296,In_256);
xnor U988 (N_988,In_71,In_944);
and U989 (N_989,In_315,In_539);
nor U990 (N_990,In_532,In_145);
or U991 (N_991,In_130,In_528);
nand U992 (N_992,In_975,In_581);
or U993 (N_993,In_33,In_246);
nand U994 (N_994,In_546,In_23);
nor U995 (N_995,In_78,In_842);
or U996 (N_996,In_431,In_285);
and U997 (N_997,In_900,In_422);
or U998 (N_998,In_679,In_480);
and U999 (N_999,In_466,In_483);
and U1000 (N_1000,In_222,In_216);
nor U1001 (N_1001,In_488,In_122);
nand U1002 (N_1002,In_461,In_835);
or U1003 (N_1003,In_881,In_188);
nor U1004 (N_1004,In_494,In_492);
and U1005 (N_1005,In_872,In_550);
nand U1006 (N_1006,In_764,In_708);
and U1007 (N_1007,In_124,In_269);
and U1008 (N_1008,In_129,In_554);
nor U1009 (N_1009,In_975,In_914);
nand U1010 (N_1010,In_325,In_320);
nand U1011 (N_1011,In_748,In_377);
or U1012 (N_1012,In_111,In_188);
and U1013 (N_1013,In_16,In_968);
nor U1014 (N_1014,In_432,In_301);
nor U1015 (N_1015,In_57,In_61);
or U1016 (N_1016,In_630,In_573);
nor U1017 (N_1017,In_642,In_163);
xor U1018 (N_1018,In_787,In_473);
and U1019 (N_1019,In_980,In_70);
nand U1020 (N_1020,In_397,In_358);
nand U1021 (N_1021,In_637,In_876);
nor U1022 (N_1022,In_506,In_976);
or U1023 (N_1023,In_384,In_625);
xor U1024 (N_1024,In_944,In_765);
nor U1025 (N_1025,In_68,In_942);
nor U1026 (N_1026,In_142,In_204);
nor U1027 (N_1027,In_208,In_553);
nand U1028 (N_1028,In_190,In_372);
or U1029 (N_1029,In_858,In_407);
xnor U1030 (N_1030,In_511,In_244);
nand U1031 (N_1031,In_821,In_962);
or U1032 (N_1032,In_169,In_146);
nor U1033 (N_1033,In_230,In_155);
nand U1034 (N_1034,In_510,In_528);
nand U1035 (N_1035,In_226,In_272);
or U1036 (N_1036,In_888,In_85);
or U1037 (N_1037,In_578,In_692);
or U1038 (N_1038,In_921,In_380);
nand U1039 (N_1039,In_257,In_445);
xnor U1040 (N_1040,In_684,In_780);
xnor U1041 (N_1041,In_294,In_689);
and U1042 (N_1042,In_493,In_475);
and U1043 (N_1043,In_573,In_117);
xnor U1044 (N_1044,In_109,In_154);
and U1045 (N_1045,In_33,In_235);
nor U1046 (N_1046,In_923,In_214);
or U1047 (N_1047,In_835,In_464);
xnor U1048 (N_1048,In_12,In_616);
nor U1049 (N_1049,In_389,In_854);
nor U1050 (N_1050,In_368,In_831);
nand U1051 (N_1051,In_834,In_712);
and U1052 (N_1052,In_432,In_624);
nand U1053 (N_1053,In_598,In_887);
and U1054 (N_1054,In_607,In_279);
nor U1055 (N_1055,In_943,In_452);
and U1056 (N_1056,In_857,In_861);
or U1057 (N_1057,In_256,In_716);
xnor U1058 (N_1058,In_73,In_999);
nor U1059 (N_1059,In_339,In_558);
nor U1060 (N_1060,In_769,In_491);
xnor U1061 (N_1061,In_622,In_667);
and U1062 (N_1062,In_340,In_406);
or U1063 (N_1063,In_246,In_963);
nand U1064 (N_1064,In_96,In_186);
nor U1065 (N_1065,In_476,In_343);
or U1066 (N_1066,In_611,In_818);
nand U1067 (N_1067,In_807,In_893);
or U1068 (N_1068,In_238,In_724);
or U1069 (N_1069,In_802,In_485);
nor U1070 (N_1070,In_220,In_687);
xnor U1071 (N_1071,In_6,In_500);
and U1072 (N_1072,In_141,In_293);
nor U1073 (N_1073,In_49,In_980);
or U1074 (N_1074,In_34,In_945);
or U1075 (N_1075,In_565,In_791);
nand U1076 (N_1076,In_103,In_284);
or U1077 (N_1077,In_273,In_293);
or U1078 (N_1078,In_276,In_40);
xor U1079 (N_1079,In_308,In_985);
and U1080 (N_1080,In_403,In_186);
and U1081 (N_1081,In_559,In_940);
and U1082 (N_1082,In_556,In_547);
or U1083 (N_1083,In_502,In_992);
and U1084 (N_1084,In_75,In_728);
and U1085 (N_1085,In_404,In_38);
or U1086 (N_1086,In_207,In_927);
or U1087 (N_1087,In_188,In_689);
or U1088 (N_1088,In_647,In_641);
nor U1089 (N_1089,In_329,In_591);
or U1090 (N_1090,In_644,In_354);
nand U1091 (N_1091,In_120,In_115);
xnor U1092 (N_1092,In_469,In_393);
and U1093 (N_1093,In_161,In_120);
or U1094 (N_1094,In_690,In_376);
nor U1095 (N_1095,In_124,In_31);
nand U1096 (N_1096,In_872,In_762);
nand U1097 (N_1097,In_550,In_573);
nor U1098 (N_1098,In_619,In_740);
and U1099 (N_1099,In_418,In_674);
nand U1100 (N_1100,In_488,In_595);
nor U1101 (N_1101,In_484,In_938);
nor U1102 (N_1102,In_926,In_583);
or U1103 (N_1103,In_599,In_87);
nor U1104 (N_1104,In_261,In_661);
nor U1105 (N_1105,In_68,In_349);
nor U1106 (N_1106,In_650,In_767);
nand U1107 (N_1107,In_329,In_515);
and U1108 (N_1108,In_104,In_169);
and U1109 (N_1109,In_418,In_800);
or U1110 (N_1110,In_2,In_825);
nor U1111 (N_1111,In_611,In_843);
and U1112 (N_1112,In_32,In_670);
nand U1113 (N_1113,In_149,In_301);
and U1114 (N_1114,In_446,In_787);
nand U1115 (N_1115,In_480,In_377);
or U1116 (N_1116,In_123,In_833);
nor U1117 (N_1117,In_643,In_754);
or U1118 (N_1118,In_837,In_237);
nor U1119 (N_1119,In_950,In_274);
and U1120 (N_1120,In_724,In_1);
or U1121 (N_1121,In_587,In_528);
and U1122 (N_1122,In_864,In_13);
nand U1123 (N_1123,In_511,In_330);
nand U1124 (N_1124,In_844,In_110);
or U1125 (N_1125,In_876,In_164);
xor U1126 (N_1126,In_293,In_280);
or U1127 (N_1127,In_929,In_331);
nand U1128 (N_1128,In_66,In_603);
nor U1129 (N_1129,In_136,In_976);
nor U1130 (N_1130,In_291,In_256);
or U1131 (N_1131,In_922,In_375);
nand U1132 (N_1132,In_371,In_185);
or U1133 (N_1133,In_942,In_885);
or U1134 (N_1134,In_978,In_53);
nand U1135 (N_1135,In_854,In_350);
or U1136 (N_1136,In_237,In_92);
or U1137 (N_1137,In_785,In_337);
xnor U1138 (N_1138,In_158,In_146);
or U1139 (N_1139,In_465,In_295);
and U1140 (N_1140,In_302,In_326);
or U1141 (N_1141,In_117,In_401);
or U1142 (N_1142,In_78,In_865);
and U1143 (N_1143,In_744,In_780);
or U1144 (N_1144,In_345,In_132);
nor U1145 (N_1145,In_880,In_202);
and U1146 (N_1146,In_505,In_37);
nor U1147 (N_1147,In_168,In_664);
and U1148 (N_1148,In_481,In_864);
xor U1149 (N_1149,In_331,In_722);
nand U1150 (N_1150,In_79,In_657);
nand U1151 (N_1151,In_603,In_72);
nor U1152 (N_1152,In_923,In_602);
or U1153 (N_1153,In_800,In_906);
nand U1154 (N_1154,In_817,In_545);
and U1155 (N_1155,In_898,In_535);
or U1156 (N_1156,In_382,In_907);
or U1157 (N_1157,In_661,In_504);
nand U1158 (N_1158,In_994,In_13);
nand U1159 (N_1159,In_76,In_622);
and U1160 (N_1160,In_592,In_386);
xnor U1161 (N_1161,In_121,In_184);
nor U1162 (N_1162,In_347,In_902);
xnor U1163 (N_1163,In_557,In_254);
nor U1164 (N_1164,In_841,In_23);
nand U1165 (N_1165,In_680,In_166);
nand U1166 (N_1166,In_614,In_849);
or U1167 (N_1167,In_310,In_973);
nor U1168 (N_1168,In_755,In_540);
and U1169 (N_1169,In_462,In_90);
nand U1170 (N_1170,In_957,In_107);
nand U1171 (N_1171,In_471,In_811);
nand U1172 (N_1172,In_706,In_870);
and U1173 (N_1173,In_985,In_144);
nand U1174 (N_1174,In_359,In_709);
nor U1175 (N_1175,In_215,In_625);
or U1176 (N_1176,In_632,In_913);
and U1177 (N_1177,In_426,In_203);
nand U1178 (N_1178,In_690,In_708);
nor U1179 (N_1179,In_460,In_516);
nor U1180 (N_1180,In_930,In_699);
and U1181 (N_1181,In_963,In_197);
nor U1182 (N_1182,In_914,In_330);
and U1183 (N_1183,In_137,In_257);
nand U1184 (N_1184,In_621,In_397);
xnor U1185 (N_1185,In_145,In_226);
or U1186 (N_1186,In_773,In_855);
nand U1187 (N_1187,In_851,In_707);
nand U1188 (N_1188,In_976,In_914);
xor U1189 (N_1189,In_703,In_830);
nor U1190 (N_1190,In_482,In_259);
nand U1191 (N_1191,In_735,In_806);
nand U1192 (N_1192,In_532,In_821);
and U1193 (N_1193,In_527,In_872);
and U1194 (N_1194,In_202,In_821);
nand U1195 (N_1195,In_700,In_843);
and U1196 (N_1196,In_722,In_425);
xor U1197 (N_1197,In_132,In_825);
and U1198 (N_1198,In_355,In_617);
and U1199 (N_1199,In_974,In_838);
nor U1200 (N_1200,In_977,In_232);
nor U1201 (N_1201,In_206,In_570);
nand U1202 (N_1202,In_865,In_986);
and U1203 (N_1203,In_312,In_236);
or U1204 (N_1204,In_680,In_73);
or U1205 (N_1205,In_891,In_359);
nand U1206 (N_1206,In_363,In_663);
or U1207 (N_1207,In_336,In_602);
nand U1208 (N_1208,In_65,In_434);
or U1209 (N_1209,In_704,In_613);
nor U1210 (N_1210,In_238,In_112);
or U1211 (N_1211,In_360,In_220);
xnor U1212 (N_1212,In_677,In_576);
and U1213 (N_1213,In_248,In_607);
nand U1214 (N_1214,In_171,In_147);
nor U1215 (N_1215,In_866,In_507);
and U1216 (N_1216,In_196,In_548);
or U1217 (N_1217,In_52,In_790);
or U1218 (N_1218,In_278,In_994);
or U1219 (N_1219,In_650,In_407);
xnor U1220 (N_1220,In_410,In_724);
nor U1221 (N_1221,In_234,In_749);
nand U1222 (N_1222,In_459,In_166);
and U1223 (N_1223,In_135,In_148);
nor U1224 (N_1224,In_358,In_900);
and U1225 (N_1225,In_502,In_722);
or U1226 (N_1226,In_860,In_872);
nand U1227 (N_1227,In_746,In_73);
nor U1228 (N_1228,In_310,In_990);
and U1229 (N_1229,In_924,In_2);
and U1230 (N_1230,In_329,In_249);
or U1231 (N_1231,In_267,In_136);
nand U1232 (N_1232,In_523,In_422);
nor U1233 (N_1233,In_263,In_576);
and U1234 (N_1234,In_549,In_836);
xor U1235 (N_1235,In_804,In_444);
nand U1236 (N_1236,In_436,In_902);
nand U1237 (N_1237,In_409,In_611);
and U1238 (N_1238,In_511,In_4);
and U1239 (N_1239,In_117,In_539);
and U1240 (N_1240,In_973,In_963);
xnor U1241 (N_1241,In_379,In_490);
nand U1242 (N_1242,In_126,In_578);
xor U1243 (N_1243,In_207,In_729);
or U1244 (N_1244,In_132,In_309);
and U1245 (N_1245,In_474,In_533);
nand U1246 (N_1246,In_255,In_974);
nand U1247 (N_1247,In_542,In_620);
nand U1248 (N_1248,In_554,In_536);
nor U1249 (N_1249,In_204,In_724);
or U1250 (N_1250,In_433,In_984);
nor U1251 (N_1251,In_589,In_359);
nor U1252 (N_1252,In_844,In_249);
nand U1253 (N_1253,In_647,In_649);
nand U1254 (N_1254,In_160,In_192);
nand U1255 (N_1255,In_751,In_447);
and U1256 (N_1256,In_593,In_157);
xnor U1257 (N_1257,In_833,In_247);
or U1258 (N_1258,In_869,In_476);
and U1259 (N_1259,In_393,In_720);
nor U1260 (N_1260,In_924,In_769);
nor U1261 (N_1261,In_352,In_612);
and U1262 (N_1262,In_879,In_381);
or U1263 (N_1263,In_772,In_271);
or U1264 (N_1264,In_324,In_949);
and U1265 (N_1265,In_358,In_552);
nor U1266 (N_1266,In_326,In_349);
nor U1267 (N_1267,In_966,In_337);
nand U1268 (N_1268,In_303,In_46);
or U1269 (N_1269,In_623,In_705);
or U1270 (N_1270,In_701,In_787);
nand U1271 (N_1271,In_96,In_431);
nand U1272 (N_1272,In_208,In_971);
xor U1273 (N_1273,In_957,In_569);
nor U1274 (N_1274,In_17,In_771);
and U1275 (N_1275,In_982,In_364);
and U1276 (N_1276,In_488,In_91);
or U1277 (N_1277,In_928,In_260);
xor U1278 (N_1278,In_664,In_511);
nand U1279 (N_1279,In_296,In_705);
nor U1280 (N_1280,In_889,In_736);
nor U1281 (N_1281,In_561,In_524);
nand U1282 (N_1282,In_158,In_40);
and U1283 (N_1283,In_860,In_305);
nand U1284 (N_1284,In_495,In_935);
xnor U1285 (N_1285,In_655,In_888);
xnor U1286 (N_1286,In_823,In_792);
nor U1287 (N_1287,In_912,In_81);
or U1288 (N_1288,In_736,In_782);
nor U1289 (N_1289,In_790,In_794);
or U1290 (N_1290,In_786,In_199);
and U1291 (N_1291,In_324,In_993);
or U1292 (N_1292,In_615,In_774);
nand U1293 (N_1293,In_147,In_833);
or U1294 (N_1294,In_225,In_919);
nor U1295 (N_1295,In_361,In_335);
or U1296 (N_1296,In_910,In_434);
nand U1297 (N_1297,In_560,In_493);
nand U1298 (N_1298,In_353,In_953);
nor U1299 (N_1299,In_463,In_154);
nand U1300 (N_1300,In_241,In_983);
nor U1301 (N_1301,In_182,In_453);
nand U1302 (N_1302,In_175,In_624);
nand U1303 (N_1303,In_0,In_421);
nand U1304 (N_1304,In_491,In_242);
nand U1305 (N_1305,In_292,In_670);
and U1306 (N_1306,In_647,In_852);
nor U1307 (N_1307,In_543,In_228);
xor U1308 (N_1308,In_13,In_277);
and U1309 (N_1309,In_783,In_852);
or U1310 (N_1310,In_247,In_821);
and U1311 (N_1311,In_764,In_679);
nor U1312 (N_1312,In_390,In_613);
nor U1313 (N_1313,In_540,In_171);
or U1314 (N_1314,In_251,In_214);
nand U1315 (N_1315,In_376,In_959);
xor U1316 (N_1316,In_142,In_279);
xnor U1317 (N_1317,In_585,In_300);
and U1318 (N_1318,In_822,In_850);
nand U1319 (N_1319,In_227,In_998);
and U1320 (N_1320,In_244,In_101);
nand U1321 (N_1321,In_360,In_124);
nand U1322 (N_1322,In_426,In_185);
and U1323 (N_1323,In_806,In_470);
nor U1324 (N_1324,In_176,In_420);
nand U1325 (N_1325,In_836,In_304);
or U1326 (N_1326,In_297,In_716);
or U1327 (N_1327,In_466,In_162);
and U1328 (N_1328,In_117,In_281);
or U1329 (N_1329,In_312,In_987);
nand U1330 (N_1330,In_231,In_875);
nor U1331 (N_1331,In_115,In_233);
and U1332 (N_1332,In_578,In_832);
xnor U1333 (N_1333,In_79,In_624);
nor U1334 (N_1334,In_963,In_636);
nand U1335 (N_1335,In_791,In_314);
nor U1336 (N_1336,In_13,In_102);
xnor U1337 (N_1337,In_299,In_561);
nor U1338 (N_1338,In_221,In_223);
xnor U1339 (N_1339,In_590,In_484);
xor U1340 (N_1340,In_368,In_706);
and U1341 (N_1341,In_345,In_651);
nand U1342 (N_1342,In_973,In_119);
and U1343 (N_1343,In_575,In_535);
and U1344 (N_1344,In_88,In_972);
nor U1345 (N_1345,In_509,In_697);
nor U1346 (N_1346,In_448,In_960);
and U1347 (N_1347,In_171,In_674);
xor U1348 (N_1348,In_496,In_60);
nor U1349 (N_1349,In_79,In_64);
xnor U1350 (N_1350,In_981,In_416);
and U1351 (N_1351,In_269,In_967);
xor U1352 (N_1352,In_782,In_134);
nor U1353 (N_1353,In_726,In_961);
nand U1354 (N_1354,In_598,In_829);
and U1355 (N_1355,In_7,In_522);
nand U1356 (N_1356,In_124,In_54);
or U1357 (N_1357,In_412,In_437);
nand U1358 (N_1358,In_482,In_342);
and U1359 (N_1359,In_692,In_160);
and U1360 (N_1360,In_136,In_211);
nand U1361 (N_1361,In_855,In_910);
nand U1362 (N_1362,In_866,In_65);
nor U1363 (N_1363,In_899,In_168);
or U1364 (N_1364,In_191,In_433);
or U1365 (N_1365,In_369,In_484);
nand U1366 (N_1366,In_826,In_760);
nand U1367 (N_1367,In_788,In_745);
or U1368 (N_1368,In_694,In_986);
or U1369 (N_1369,In_629,In_548);
xor U1370 (N_1370,In_154,In_852);
nor U1371 (N_1371,In_855,In_284);
and U1372 (N_1372,In_744,In_106);
nand U1373 (N_1373,In_406,In_951);
nand U1374 (N_1374,In_923,In_443);
xor U1375 (N_1375,In_359,In_358);
and U1376 (N_1376,In_804,In_255);
or U1377 (N_1377,In_617,In_605);
or U1378 (N_1378,In_48,In_275);
or U1379 (N_1379,In_689,In_316);
nand U1380 (N_1380,In_973,In_83);
nand U1381 (N_1381,In_254,In_260);
and U1382 (N_1382,In_415,In_612);
and U1383 (N_1383,In_680,In_776);
and U1384 (N_1384,In_871,In_312);
or U1385 (N_1385,In_358,In_221);
nor U1386 (N_1386,In_164,In_82);
or U1387 (N_1387,In_434,In_239);
nor U1388 (N_1388,In_880,In_661);
nor U1389 (N_1389,In_288,In_850);
and U1390 (N_1390,In_141,In_625);
nand U1391 (N_1391,In_931,In_837);
nand U1392 (N_1392,In_897,In_310);
or U1393 (N_1393,In_149,In_293);
and U1394 (N_1394,In_141,In_317);
xnor U1395 (N_1395,In_902,In_17);
nor U1396 (N_1396,In_924,In_324);
and U1397 (N_1397,In_843,In_580);
nor U1398 (N_1398,In_42,In_72);
nor U1399 (N_1399,In_120,In_942);
nand U1400 (N_1400,In_290,In_904);
nor U1401 (N_1401,In_71,In_109);
nand U1402 (N_1402,In_396,In_539);
nand U1403 (N_1403,In_143,In_879);
or U1404 (N_1404,In_673,In_20);
or U1405 (N_1405,In_781,In_75);
or U1406 (N_1406,In_232,In_100);
nor U1407 (N_1407,In_869,In_724);
or U1408 (N_1408,In_654,In_106);
nor U1409 (N_1409,In_55,In_248);
nand U1410 (N_1410,In_664,In_181);
and U1411 (N_1411,In_403,In_202);
nor U1412 (N_1412,In_158,In_669);
or U1413 (N_1413,In_357,In_545);
and U1414 (N_1414,In_627,In_194);
nand U1415 (N_1415,In_291,In_616);
nor U1416 (N_1416,In_391,In_800);
or U1417 (N_1417,In_702,In_723);
nor U1418 (N_1418,In_73,In_298);
nor U1419 (N_1419,In_117,In_813);
nand U1420 (N_1420,In_721,In_626);
nor U1421 (N_1421,In_60,In_27);
nor U1422 (N_1422,In_145,In_306);
and U1423 (N_1423,In_25,In_88);
or U1424 (N_1424,In_812,In_996);
nor U1425 (N_1425,In_768,In_631);
nor U1426 (N_1426,In_43,In_564);
xnor U1427 (N_1427,In_287,In_10);
or U1428 (N_1428,In_586,In_737);
nand U1429 (N_1429,In_292,In_729);
nor U1430 (N_1430,In_926,In_568);
or U1431 (N_1431,In_408,In_585);
nor U1432 (N_1432,In_698,In_842);
and U1433 (N_1433,In_484,In_116);
and U1434 (N_1434,In_974,In_869);
nand U1435 (N_1435,In_945,In_504);
nand U1436 (N_1436,In_89,In_890);
nand U1437 (N_1437,In_951,In_217);
nor U1438 (N_1438,In_551,In_776);
or U1439 (N_1439,In_706,In_85);
and U1440 (N_1440,In_808,In_759);
or U1441 (N_1441,In_671,In_10);
or U1442 (N_1442,In_328,In_614);
xnor U1443 (N_1443,In_792,In_75);
nand U1444 (N_1444,In_348,In_209);
xnor U1445 (N_1445,In_206,In_652);
or U1446 (N_1446,In_794,In_464);
nor U1447 (N_1447,In_307,In_399);
nor U1448 (N_1448,In_368,In_766);
nand U1449 (N_1449,In_519,In_209);
or U1450 (N_1450,In_676,In_839);
nand U1451 (N_1451,In_898,In_569);
nor U1452 (N_1452,In_422,In_950);
or U1453 (N_1453,In_420,In_389);
nand U1454 (N_1454,In_431,In_640);
nor U1455 (N_1455,In_925,In_486);
nor U1456 (N_1456,In_701,In_51);
or U1457 (N_1457,In_805,In_856);
nand U1458 (N_1458,In_33,In_622);
or U1459 (N_1459,In_640,In_777);
or U1460 (N_1460,In_644,In_714);
or U1461 (N_1461,In_220,In_490);
nand U1462 (N_1462,In_570,In_910);
and U1463 (N_1463,In_964,In_93);
xor U1464 (N_1464,In_237,In_365);
nor U1465 (N_1465,In_973,In_622);
nor U1466 (N_1466,In_458,In_746);
or U1467 (N_1467,In_304,In_615);
nor U1468 (N_1468,In_330,In_509);
and U1469 (N_1469,In_359,In_110);
and U1470 (N_1470,In_703,In_425);
xor U1471 (N_1471,In_596,In_288);
and U1472 (N_1472,In_825,In_389);
and U1473 (N_1473,In_737,In_263);
nand U1474 (N_1474,In_942,In_74);
or U1475 (N_1475,In_146,In_767);
or U1476 (N_1476,In_536,In_747);
nand U1477 (N_1477,In_554,In_782);
or U1478 (N_1478,In_980,In_480);
or U1479 (N_1479,In_908,In_626);
nor U1480 (N_1480,In_313,In_739);
nand U1481 (N_1481,In_261,In_343);
and U1482 (N_1482,In_215,In_696);
nor U1483 (N_1483,In_890,In_824);
xnor U1484 (N_1484,In_738,In_14);
nor U1485 (N_1485,In_978,In_12);
and U1486 (N_1486,In_889,In_730);
and U1487 (N_1487,In_494,In_15);
nand U1488 (N_1488,In_352,In_106);
and U1489 (N_1489,In_131,In_152);
xnor U1490 (N_1490,In_571,In_855);
xor U1491 (N_1491,In_901,In_260);
or U1492 (N_1492,In_207,In_815);
nand U1493 (N_1493,In_417,In_649);
nand U1494 (N_1494,In_79,In_441);
and U1495 (N_1495,In_913,In_287);
nand U1496 (N_1496,In_390,In_421);
and U1497 (N_1497,In_369,In_342);
or U1498 (N_1498,In_459,In_687);
nor U1499 (N_1499,In_795,In_545);
nor U1500 (N_1500,In_809,In_491);
or U1501 (N_1501,In_145,In_283);
nand U1502 (N_1502,In_156,In_750);
nor U1503 (N_1503,In_353,In_477);
or U1504 (N_1504,In_641,In_91);
nand U1505 (N_1505,In_360,In_539);
and U1506 (N_1506,In_144,In_614);
and U1507 (N_1507,In_557,In_838);
or U1508 (N_1508,In_131,In_620);
nand U1509 (N_1509,In_846,In_760);
xor U1510 (N_1510,In_281,In_245);
nand U1511 (N_1511,In_943,In_912);
nor U1512 (N_1512,In_949,In_101);
nor U1513 (N_1513,In_887,In_492);
nor U1514 (N_1514,In_53,In_139);
or U1515 (N_1515,In_92,In_197);
nor U1516 (N_1516,In_34,In_199);
xnor U1517 (N_1517,In_74,In_875);
nand U1518 (N_1518,In_187,In_501);
nor U1519 (N_1519,In_695,In_405);
and U1520 (N_1520,In_890,In_810);
nor U1521 (N_1521,In_376,In_105);
nor U1522 (N_1522,In_420,In_750);
nand U1523 (N_1523,In_549,In_698);
or U1524 (N_1524,In_760,In_970);
and U1525 (N_1525,In_845,In_647);
xor U1526 (N_1526,In_88,In_161);
or U1527 (N_1527,In_621,In_450);
or U1528 (N_1528,In_642,In_519);
nand U1529 (N_1529,In_318,In_527);
nand U1530 (N_1530,In_282,In_816);
or U1531 (N_1531,In_570,In_28);
nand U1532 (N_1532,In_851,In_458);
xor U1533 (N_1533,In_217,In_378);
and U1534 (N_1534,In_435,In_932);
nor U1535 (N_1535,In_708,In_621);
and U1536 (N_1536,In_862,In_863);
nand U1537 (N_1537,In_962,In_460);
xnor U1538 (N_1538,In_249,In_206);
nand U1539 (N_1539,In_58,In_240);
and U1540 (N_1540,In_38,In_187);
nor U1541 (N_1541,In_597,In_929);
or U1542 (N_1542,In_175,In_496);
xor U1543 (N_1543,In_489,In_770);
nand U1544 (N_1544,In_335,In_258);
nand U1545 (N_1545,In_955,In_423);
or U1546 (N_1546,In_940,In_976);
and U1547 (N_1547,In_615,In_850);
nor U1548 (N_1548,In_534,In_323);
xor U1549 (N_1549,In_786,In_279);
and U1550 (N_1550,In_237,In_965);
nand U1551 (N_1551,In_21,In_985);
or U1552 (N_1552,In_296,In_246);
xnor U1553 (N_1553,In_465,In_956);
nor U1554 (N_1554,In_201,In_72);
or U1555 (N_1555,In_352,In_516);
nor U1556 (N_1556,In_345,In_56);
or U1557 (N_1557,In_981,In_263);
and U1558 (N_1558,In_233,In_286);
and U1559 (N_1559,In_419,In_77);
nand U1560 (N_1560,In_343,In_512);
and U1561 (N_1561,In_316,In_565);
and U1562 (N_1562,In_670,In_918);
nand U1563 (N_1563,In_762,In_996);
nor U1564 (N_1564,In_837,In_894);
nand U1565 (N_1565,In_559,In_612);
xnor U1566 (N_1566,In_268,In_763);
nor U1567 (N_1567,In_73,In_147);
xnor U1568 (N_1568,In_852,In_689);
nor U1569 (N_1569,In_599,In_849);
and U1570 (N_1570,In_38,In_699);
and U1571 (N_1571,In_919,In_523);
and U1572 (N_1572,In_550,In_320);
and U1573 (N_1573,In_338,In_98);
nand U1574 (N_1574,In_173,In_572);
nor U1575 (N_1575,In_704,In_739);
and U1576 (N_1576,In_479,In_733);
or U1577 (N_1577,In_285,In_421);
nor U1578 (N_1578,In_201,In_157);
or U1579 (N_1579,In_80,In_56);
and U1580 (N_1580,In_881,In_640);
nand U1581 (N_1581,In_512,In_685);
and U1582 (N_1582,In_865,In_664);
nor U1583 (N_1583,In_422,In_406);
nand U1584 (N_1584,In_900,In_703);
or U1585 (N_1585,In_765,In_742);
or U1586 (N_1586,In_136,In_770);
nor U1587 (N_1587,In_394,In_934);
nand U1588 (N_1588,In_881,In_409);
nor U1589 (N_1589,In_651,In_114);
or U1590 (N_1590,In_580,In_643);
or U1591 (N_1591,In_581,In_522);
xnor U1592 (N_1592,In_8,In_217);
and U1593 (N_1593,In_888,In_213);
nand U1594 (N_1594,In_617,In_148);
xnor U1595 (N_1595,In_0,In_15);
or U1596 (N_1596,In_557,In_648);
nand U1597 (N_1597,In_850,In_738);
nor U1598 (N_1598,In_776,In_882);
nand U1599 (N_1599,In_807,In_955);
nand U1600 (N_1600,In_348,In_692);
and U1601 (N_1601,In_839,In_326);
and U1602 (N_1602,In_510,In_795);
xor U1603 (N_1603,In_6,In_169);
and U1604 (N_1604,In_477,In_174);
nor U1605 (N_1605,In_479,In_478);
and U1606 (N_1606,In_604,In_478);
nor U1607 (N_1607,In_436,In_452);
nor U1608 (N_1608,In_945,In_508);
nand U1609 (N_1609,In_554,In_547);
or U1610 (N_1610,In_215,In_26);
nand U1611 (N_1611,In_307,In_358);
xnor U1612 (N_1612,In_13,In_477);
nor U1613 (N_1613,In_42,In_837);
and U1614 (N_1614,In_43,In_368);
and U1615 (N_1615,In_360,In_392);
or U1616 (N_1616,In_290,In_402);
and U1617 (N_1617,In_280,In_268);
xor U1618 (N_1618,In_578,In_398);
and U1619 (N_1619,In_90,In_48);
nor U1620 (N_1620,In_670,In_408);
xor U1621 (N_1621,In_224,In_342);
nor U1622 (N_1622,In_528,In_459);
nor U1623 (N_1623,In_454,In_39);
or U1624 (N_1624,In_357,In_392);
nand U1625 (N_1625,In_61,In_766);
and U1626 (N_1626,In_162,In_279);
and U1627 (N_1627,In_713,In_21);
or U1628 (N_1628,In_833,In_285);
nor U1629 (N_1629,In_30,In_43);
nand U1630 (N_1630,In_104,In_612);
nand U1631 (N_1631,In_677,In_24);
nand U1632 (N_1632,In_152,In_975);
or U1633 (N_1633,In_866,In_93);
or U1634 (N_1634,In_995,In_510);
nand U1635 (N_1635,In_912,In_575);
or U1636 (N_1636,In_247,In_697);
nand U1637 (N_1637,In_475,In_325);
nand U1638 (N_1638,In_626,In_14);
nand U1639 (N_1639,In_394,In_206);
and U1640 (N_1640,In_732,In_317);
nand U1641 (N_1641,In_39,In_402);
and U1642 (N_1642,In_205,In_57);
or U1643 (N_1643,In_743,In_748);
nor U1644 (N_1644,In_84,In_553);
nand U1645 (N_1645,In_162,In_771);
and U1646 (N_1646,In_808,In_154);
and U1647 (N_1647,In_296,In_782);
xnor U1648 (N_1648,In_630,In_165);
nor U1649 (N_1649,In_358,In_602);
and U1650 (N_1650,In_637,In_916);
nor U1651 (N_1651,In_105,In_636);
or U1652 (N_1652,In_390,In_643);
nand U1653 (N_1653,In_570,In_774);
nand U1654 (N_1654,In_881,In_710);
xnor U1655 (N_1655,In_511,In_451);
and U1656 (N_1656,In_630,In_476);
and U1657 (N_1657,In_832,In_791);
or U1658 (N_1658,In_237,In_782);
nand U1659 (N_1659,In_164,In_19);
or U1660 (N_1660,In_778,In_910);
and U1661 (N_1661,In_364,In_490);
and U1662 (N_1662,In_289,In_91);
nor U1663 (N_1663,In_425,In_220);
and U1664 (N_1664,In_14,In_878);
or U1665 (N_1665,In_607,In_722);
nand U1666 (N_1666,In_213,In_2);
or U1667 (N_1667,In_145,In_291);
nor U1668 (N_1668,In_743,In_367);
nor U1669 (N_1669,In_908,In_256);
and U1670 (N_1670,In_255,In_616);
or U1671 (N_1671,In_805,In_377);
nor U1672 (N_1672,In_354,In_265);
nand U1673 (N_1673,In_516,In_780);
nand U1674 (N_1674,In_27,In_323);
and U1675 (N_1675,In_563,In_942);
nor U1676 (N_1676,In_381,In_408);
xnor U1677 (N_1677,In_359,In_336);
and U1678 (N_1678,In_203,In_352);
or U1679 (N_1679,In_594,In_767);
or U1680 (N_1680,In_568,In_763);
nor U1681 (N_1681,In_719,In_181);
nand U1682 (N_1682,In_829,In_523);
nor U1683 (N_1683,In_625,In_895);
nor U1684 (N_1684,In_466,In_449);
nor U1685 (N_1685,In_517,In_943);
nor U1686 (N_1686,In_168,In_724);
nand U1687 (N_1687,In_563,In_526);
and U1688 (N_1688,In_883,In_813);
nand U1689 (N_1689,In_218,In_626);
nand U1690 (N_1690,In_400,In_784);
xnor U1691 (N_1691,In_540,In_163);
xnor U1692 (N_1692,In_694,In_617);
nor U1693 (N_1693,In_625,In_958);
and U1694 (N_1694,In_992,In_261);
nor U1695 (N_1695,In_393,In_541);
nor U1696 (N_1696,In_790,In_422);
nand U1697 (N_1697,In_536,In_75);
nand U1698 (N_1698,In_293,In_930);
nor U1699 (N_1699,In_872,In_757);
and U1700 (N_1700,In_356,In_263);
nand U1701 (N_1701,In_823,In_455);
and U1702 (N_1702,In_713,In_868);
xnor U1703 (N_1703,In_172,In_719);
and U1704 (N_1704,In_95,In_911);
nand U1705 (N_1705,In_816,In_544);
nand U1706 (N_1706,In_551,In_856);
or U1707 (N_1707,In_297,In_439);
nor U1708 (N_1708,In_84,In_25);
nand U1709 (N_1709,In_485,In_9);
nor U1710 (N_1710,In_391,In_978);
or U1711 (N_1711,In_254,In_796);
or U1712 (N_1712,In_399,In_234);
xor U1713 (N_1713,In_792,In_469);
nor U1714 (N_1714,In_449,In_502);
xnor U1715 (N_1715,In_842,In_163);
and U1716 (N_1716,In_251,In_125);
and U1717 (N_1717,In_835,In_745);
or U1718 (N_1718,In_61,In_813);
nand U1719 (N_1719,In_220,In_981);
nand U1720 (N_1720,In_885,In_441);
or U1721 (N_1721,In_622,In_577);
and U1722 (N_1722,In_888,In_251);
or U1723 (N_1723,In_590,In_182);
or U1724 (N_1724,In_333,In_253);
or U1725 (N_1725,In_568,In_429);
or U1726 (N_1726,In_457,In_193);
or U1727 (N_1727,In_450,In_420);
and U1728 (N_1728,In_808,In_964);
nand U1729 (N_1729,In_231,In_954);
nand U1730 (N_1730,In_786,In_905);
and U1731 (N_1731,In_604,In_280);
or U1732 (N_1732,In_978,In_792);
nand U1733 (N_1733,In_771,In_837);
nand U1734 (N_1734,In_428,In_260);
xnor U1735 (N_1735,In_417,In_82);
nand U1736 (N_1736,In_370,In_102);
and U1737 (N_1737,In_183,In_355);
and U1738 (N_1738,In_959,In_445);
or U1739 (N_1739,In_376,In_393);
or U1740 (N_1740,In_413,In_486);
nand U1741 (N_1741,In_138,In_715);
nand U1742 (N_1742,In_137,In_618);
nand U1743 (N_1743,In_955,In_28);
and U1744 (N_1744,In_69,In_597);
and U1745 (N_1745,In_679,In_962);
and U1746 (N_1746,In_915,In_690);
and U1747 (N_1747,In_869,In_462);
nand U1748 (N_1748,In_374,In_995);
nand U1749 (N_1749,In_261,In_471);
and U1750 (N_1750,In_466,In_114);
nand U1751 (N_1751,In_550,In_580);
or U1752 (N_1752,In_922,In_134);
xor U1753 (N_1753,In_623,In_425);
nor U1754 (N_1754,In_391,In_804);
and U1755 (N_1755,In_253,In_635);
nand U1756 (N_1756,In_539,In_705);
or U1757 (N_1757,In_647,In_484);
and U1758 (N_1758,In_803,In_708);
and U1759 (N_1759,In_176,In_706);
or U1760 (N_1760,In_251,In_658);
nor U1761 (N_1761,In_590,In_142);
nor U1762 (N_1762,In_815,In_763);
nor U1763 (N_1763,In_621,In_829);
or U1764 (N_1764,In_960,In_357);
or U1765 (N_1765,In_72,In_149);
xor U1766 (N_1766,In_768,In_712);
nand U1767 (N_1767,In_313,In_419);
nor U1768 (N_1768,In_998,In_295);
nor U1769 (N_1769,In_518,In_152);
or U1770 (N_1770,In_636,In_388);
or U1771 (N_1771,In_181,In_593);
or U1772 (N_1772,In_375,In_73);
or U1773 (N_1773,In_174,In_884);
nor U1774 (N_1774,In_36,In_262);
nor U1775 (N_1775,In_902,In_659);
and U1776 (N_1776,In_655,In_507);
xor U1777 (N_1777,In_601,In_649);
xnor U1778 (N_1778,In_482,In_105);
or U1779 (N_1779,In_337,In_823);
and U1780 (N_1780,In_759,In_973);
nor U1781 (N_1781,In_408,In_855);
or U1782 (N_1782,In_274,In_283);
nand U1783 (N_1783,In_147,In_635);
nor U1784 (N_1784,In_376,In_581);
nor U1785 (N_1785,In_776,In_27);
nand U1786 (N_1786,In_382,In_379);
or U1787 (N_1787,In_171,In_866);
xor U1788 (N_1788,In_765,In_843);
nor U1789 (N_1789,In_86,In_628);
and U1790 (N_1790,In_937,In_601);
or U1791 (N_1791,In_129,In_328);
nor U1792 (N_1792,In_147,In_953);
and U1793 (N_1793,In_35,In_690);
nor U1794 (N_1794,In_405,In_676);
and U1795 (N_1795,In_59,In_772);
nor U1796 (N_1796,In_602,In_107);
nand U1797 (N_1797,In_95,In_388);
xor U1798 (N_1798,In_110,In_818);
nor U1799 (N_1799,In_229,In_533);
nand U1800 (N_1800,In_965,In_907);
or U1801 (N_1801,In_518,In_176);
or U1802 (N_1802,In_201,In_497);
nor U1803 (N_1803,In_81,In_196);
or U1804 (N_1804,In_264,In_153);
xor U1805 (N_1805,In_417,In_148);
nor U1806 (N_1806,In_462,In_334);
and U1807 (N_1807,In_401,In_221);
nand U1808 (N_1808,In_506,In_291);
or U1809 (N_1809,In_212,In_997);
or U1810 (N_1810,In_623,In_813);
and U1811 (N_1811,In_865,In_962);
nand U1812 (N_1812,In_547,In_187);
and U1813 (N_1813,In_14,In_310);
nand U1814 (N_1814,In_364,In_395);
or U1815 (N_1815,In_50,In_934);
or U1816 (N_1816,In_688,In_8);
and U1817 (N_1817,In_322,In_902);
xor U1818 (N_1818,In_675,In_504);
and U1819 (N_1819,In_896,In_368);
and U1820 (N_1820,In_405,In_536);
nand U1821 (N_1821,In_387,In_928);
and U1822 (N_1822,In_153,In_704);
nand U1823 (N_1823,In_462,In_557);
nor U1824 (N_1824,In_274,In_611);
nand U1825 (N_1825,In_767,In_856);
and U1826 (N_1826,In_446,In_170);
nand U1827 (N_1827,In_156,In_963);
nand U1828 (N_1828,In_997,In_316);
and U1829 (N_1829,In_907,In_560);
or U1830 (N_1830,In_126,In_631);
nand U1831 (N_1831,In_533,In_785);
xnor U1832 (N_1832,In_162,In_394);
or U1833 (N_1833,In_478,In_467);
or U1834 (N_1834,In_831,In_79);
and U1835 (N_1835,In_135,In_915);
or U1836 (N_1836,In_572,In_237);
and U1837 (N_1837,In_291,In_50);
nand U1838 (N_1838,In_592,In_226);
and U1839 (N_1839,In_934,In_812);
or U1840 (N_1840,In_286,In_603);
or U1841 (N_1841,In_638,In_337);
nand U1842 (N_1842,In_884,In_401);
or U1843 (N_1843,In_372,In_883);
nor U1844 (N_1844,In_687,In_88);
nor U1845 (N_1845,In_771,In_134);
or U1846 (N_1846,In_180,In_473);
nand U1847 (N_1847,In_983,In_411);
xor U1848 (N_1848,In_425,In_381);
and U1849 (N_1849,In_302,In_316);
or U1850 (N_1850,In_52,In_141);
nand U1851 (N_1851,In_71,In_503);
nor U1852 (N_1852,In_185,In_301);
and U1853 (N_1853,In_790,In_667);
nor U1854 (N_1854,In_730,In_54);
or U1855 (N_1855,In_75,In_486);
and U1856 (N_1856,In_394,In_539);
xnor U1857 (N_1857,In_440,In_464);
xnor U1858 (N_1858,In_249,In_838);
nor U1859 (N_1859,In_27,In_694);
or U1860 (N_1860,In_412,In_354);
nor U1861 (N_1861,In_970,In_79);
and U1862 (N_1862,In_248,In_511);
and U1863 (N_1863,In_985,In_369);
nand U1864 (N_1864,In_899,In_801);
nor U1865 (N_1865,In_880,In_691);
and U1866 (N_1866,In_612,In_390);
nor U1867 (N_1867,In_466,In_779);
and U1868 (N_1868,In_512,In_69);
or U1869 (N_1869,In_163,In_853);
nand U1870 (N_1870,In_702,In_772);
xor U1871 (N_1871,In_715,In_354);
or U1872 (N_1872,In_543,In_96);
or U1873 (N_1873,In_233,In_303);
nand U1874 (N_1874,In_127,In_93);
xnor U1875 (N_1875,In_431,In_83);
nor U1876 (N_1876,In_458,In_818);
or U1877 (N_1877,In_546,In_298);
xnor U1878 (N_1878,In_633,In_615);
nor U1879 (N_1879,In_608,In_931);
and U1880 (N_1880,In_964,In_488);
and U1881 (N_1881,In_383,In_756);
nand U1882 (N_1882,In_318,In_880);
nand U1883 (N_1883,In_79,In_57);
nand U1884 (N_1884,In_681,In_718);
and U1885 (N_1885,In_422,In_118);
nand U1886 (N_1886,In_736,In_588);
and U1887 (N_1887,In_376,In_107);
xor U1888 (N_1888,In_134,In_450);
nand U1889 (N_1889,In_679,In_642);
and U1890 (N_1890,In_477,In_248);
or U1891 (N_1891,In_729,In_865);
or U1892 (N_1892,In_173,In_912);
xor U1893 (N_1893,In_333,In_699);
nor U1894 (N_1894,In_93,In_773);
nor U1895 (N_1895,In_536,In_278);
and U1896 (N_1896,In_143,In_40);
nand U1897 (N_1897,In_571,In_707);
and U1898 (N_1898,In_117,In_660);
nor U1899 (N_1899,In_520,In_538);
and U1900 (N_1900,In_570,In_551);
or U1901 (N_1901,In_724,In_826);
and U1902 (N_1902,In_173,In_37);
or U1903 (N_1903,In_867,In_669);
xnor U1904 (N_1904,In_330,In_313);
nor U1905 (N_1905,In_989,In_474);
nand U1906 (N_1906,In_403,In_120);
and U1907 (N_1907,In_794,In_245);
nor U1908 (N_1908,In_894,In_986);
xnor U1909 (N_1909,In_746,In_834);
xnor U1910 (N_1910,In_680,In_459);
or U1911 (N_1911,In_455,In_284);
nand U1912 (N_1912,In_674,In_97);
nor U1913 (N_1913,In_254,In_765);
xor U1914 (N_1914,In_610,In_996);
or U1915 (N_1915,In_499,In_952);
nand U1916 (N_1916,In_335,In_288);
or U1917 (N_1917,In_96,In_240);
nor U1918 (N_1918,In_388,In_626);
and U1919 (N_1919,In_212,In_296);
and U1920 (N_1920,In_592,In_607);
or U1921 (N_1921,In_503,In_81);
or U1922 (N_1922,In_253,In_776);
xor U1923 (N_1923,In_990,In_635);
and U1924 (N_1924,In_584,In_425);
and U1925 (N_1925,In_283,In_930);
nand U1926 (N_1926,In_357,In_14);
xnor U1927 (N_1927,In_107,In_38);
and U1928 (N_1928,In_608,In_176);
nand U1929 (N_1929,In_188,In_544);
or U1930 (N_1930,In_499,In_647);
xnor U1931 (N_1931,In_908,In_792);
xor U1932 (N_1932,In_273,In_549);
nor U1933 (N_1933,In_23,In_596);
nor U1934 (N_1934,In_189,In_364);
and U1935 (N_1935,In_431,In_615);
and U1936 (N_1936,In_470,In_745);
or U1937 (N_1937,In_963,In_851);
nand U1938 (N_1938,In_110,In_668);
nand U1939 (N_1939,In_806,In_170);
nand U1940 (N_1940,In_205,In_788);
or U1941 (N_1941,In_304,In_929);
or U1942 (N_1942,In_930,In_914);
and U1943 (N_1943,In_868,In_995);
or U1944 (N_1944,In_99,In_958);
and U1945 (N_1945,In_783,In_543);
nand U1946 (N_1946,In_620,In_464);
nand U1947 (N_1947,In_71,In_156);
and U1948 (N_1948,In_184,In_401);
xnor U1949 (N_1949,In_394,In_985);
and U1950 (N_1950,In_486,In_174);
nor U1951 (N_1951,In_956,In_299);
nand U1952 (N_1952,In_33,In_912);
and U1953 (N_1953,In_336,In_235);
nand U1954 (N_1954,In_546,In_888);
and U1955 (N_1955,In_493,In_957);
and U1956 (N_1956,In_581,In_437);
nand U1957 (N_1957,In_284,In_183);
nor U1958 (N_1958,In_42,In_760);
nor U1959 (N_1959,In_181,In_683);
and U1960 (N_1960,In_471,In_387);
or U1961 (N_1961,In_592,In_942);
nor U1962 (N_1962,In_691,In_186);
and U1963 (N_1963,In_801,In_986);
nor U1964 (N_1964,In_327,In_114);
nand U1965 (N_1965,In_759,In_694);
nand U1966 (N_1966,In_437,In_565);
xnor U1967 (N_1967,In_494,In_819);
nor U1968 (N_1968,In_182,In_110);
or U1969 (N_1969,In_982,In_959);
and U1970 (N_1970,In_887,In_487);
xnor U1971 (N_1971,In_87,In_340);
and U1972 (N_1972,In_762,In_334);
or U1973 (N_1973,In_452,In_183);
and U1974 (N_1974,In_779,In_521);
nand U1975 (N_1975,In_983,In_929);
nor U1976 (N_1976,In_286,In_491);
and U1977 (N_1977,In_280,In_528);
nand U1978 (N_1978,In_322,In_94);
xnor U1979 (N_1979,In_666,In_239);
or U1980 (N_1980,In_352,In_957);
nor U1981 (N_1981,In_630,In_322);
or U1982 (N_1982,In_228,In_610);
nand U1983 (N_1983,In_623,In_943);
or U1984 (N_1984,In_556,In_356);
nand U1985 (N_1985,In_824,In_713);
xnor U1986 (N_1986,In_676,In_973);
nor U1987 (N_1987,In_549,In_834);
xor U1988 (N_1988,In_666,In_729);
or U1989 (N_1989,In_368,In_948);
and U1990 (N_1990,In_118,In_815);
or U1991 (N_1991,In_796,In_760);
nor U1992 (N_1992,In_143,In_836);
or U1993 (N_1993,In_129,In_297);
nand U1994 (N_1994,In_775,In_173);
or U1995 (N_1995,In_981,In_385);
nand U1996 (N_1996,In_814,In_7);
and U1997 (N_1997,In_95,In_714);
or U1998 (N_1998,In_81,In_263);
or U1999 (N_1999,In_668,In_543);
and U2000 (N_2000,In_910,In_696);
and U2001 (N_2001,In_462,In_584);
xor U2002 (N_2002,In_44,In_26);
nor U2003 (N_2003,In_146,In_997);
xnor U2004 (N_2004,In_803,In_546);
nand U2005 (N_2005,In_534,In_935);
and U2006 (N_2006,In_458,In_142);
and U2007 (N_2007,In_194,In_806);
and U2008 (N_2008,In_254,In_634);
nor U2009 (N_2009,In_843,In_464);
nand U2010 (N_2010,In_657,In_816);
nand U2011 (N_2011,In_874,In_428);
nand U2012 (N_2012,In_348,In_211);
nor U2013 (N_2013,In_138,In_189);
or U2014 (N_2014,In_673,In_487);
nand U2015 (N_2015,In_184,In_535);
nand U2016 (N_2016,In_883,In_700);
or U2017 (N_2017,In_757,In_29);
nand U2018 (N_2018,In_709,In_903);
xnor U2019 (N_2019,In_286,In_657);
or U2020 (N_2020,In_26,In_49);
or U2021 (N_2021,In_781,In_138);
nor U2022 (N_2022,In_656,In_853);
and U2023 (N_2023,In_321,In_575);
or U2024 (N_2024,In_351,In_151);
and U2025 (N_2025,In_235,In_437);
xor U2026 (N_2026,In_293,In_427);
or U2027 (N_2027,In_470,In_256);
nand U2028 (N_2028,In_278,In_193);
and U2029 (N_2029,In_571,In_756);
nor U2030 (N_2030,In_705,In_775);
and U2031 (N_2031,In_469,In_471);
and U2032 (N_2032,In_906,In_58);
nor U2033 (N_2033,In_455,In_992);
and U2034 (N_2034,In_638,In_102);
nor U2035 (N_2035,In_557,In_981);
xnor U2036 (N_2036,In_392,In_135);
and U2037 (N_2037,In_711,In_216);
or U2038 (N_2038,In_150,In_121);
nor U2039 (N_2039,In_962,In_669);
and U2040 (N_2040,In_804,In_979);
nor U2041 (N_2041,In_226,In_593);
and U2042 (N_2042,In_768,In_119);
or U2043 (N_2043,In_249,In_900);
or U2044 (N_2044,In_497,In_511);
and U2045 (N_2045,In_810,In_563);
or U2046 (N_2046,In_590,In_165);
nor U2047 (N_2047,In_833,In_795);
nor U2048 (N_2048,In_641,In_438);
nor U2049 (N_2049,In_247,In_190);
nand U2050 (N_2050,In_518,In_952);
nor U2051 (N_2051,In_716,In_489);
nand U2052 (N_2052,In_895,In_894);
or U2053 (N_2053,In_223,In_347);
or U2054 (N_2054,In_890,In_905);
and U2055 (N_2055,In_840,In_938);
or U2056 (N_2056,In_60,In_599);
and U2057 (N_2057,In_890,In_5);
nor U2058 (N_2058,In_750,In_199);
or U2059 (N_2059,In_40,In_134);
nand U2060 (N_2060,In_974,In_459);
or U2061 (N_2061,In_984,In_884);
nor U2062 (N_2062,In_366,In_434);
and U2063 (N_2063,In_101,In_229);
and U2064 (N_2064,In_379,In_104);
nand U2065 (N_2065,In_632,In_329);
nor U2066 (N_2066,In_590,In_130);
nand U2067 (N_2067,In_708,In_807);
or U2068 (N_2068,In_547,In_71);
nand U2069 (N_2069,In_84,In_77);
and U2070 (N_2070,In_310,In_16);
or U2071 (N_2071,In_77,In_196);
nand U2072 (N_2072,In_347,In_887);
and U2073 (N_2073,In_477,In_180);
nor U2074 (N_2074,In_151,In_643);
and U2075 (N_2075,In_117,In_988);
or U2076 (N_2076,In_77,In_97);
and U2077 (N_2077,In_839,In_777);
nand U2078 (N_2078,In_10,In_872);
xor U2079 (N_2079,In_975,In_202);
xor U2080 (N_2080,In_889,In_527);
nand U2081 (N_2081,In_798,In_429);
nor U2082 (N_2082,In_922,In_174);
or U2083 (N_2083,In_42,In_84);
and U2084 (N_2084,In_233,In_674);
xnor U2085 (N_2085,In_50,In_456);
xnor U2086 (N_2086,In_432,In_772);
nand U2087 (N_2087,In_285,In_452);
or U2088 (N_2088,In_461,In_508);
nor U2089 (N_2089,In_503,In_319);
xor U2090 (N_2090,In_722,In_129);
nor U2091 (N_2091,In_716,In_5);
and U2092 (N_2092,In_800,In_863);
xor U2093 (N_2093,In_436,In_774);
nor U2094 (N_2094,In_343,In_459);
and U2095 (N_2095,In_645,In_495);
nor U2096 (N_2096,In_553,In_887);
nor U2097 (N_2097,In_338,In_646);
nand U2098 (N_2098,In_899,In_74);
and U2099 (N_2099,In_94,In_35);
nor U2100 (N_2100,In_911,In_445);
nand U2101 (N_2101,In_625,In_111);
or U2102 (N_2102,In_870,In_581);
and U2103 (N_2103,In_701,In_906);
nand U2104 (N_2104,In_730,In_196);
or U2105 (N_2105,In_717,In_670);
or U2106 (N_2106,In_864,In_155);
nand U2107 (N_2107,In_774,In_713);
or U2108 (N_2108,In_59,In_11);
xnor U2109 (N_2109,In_703,In_540);
xnor U2110 (N_2110,In_176,In_596);
nor U2111 (N_2111,In_445,In_776);
nor U2112 (N_2112,In_69,In_666);
or U2113 (N_2113,In_689,In_487);
nand U2114 (N_2114,In_507,In_796);
or U2115 (N_2115,In_294,In_906);
nand U2116 (N_2116,In_795,In_387);
nand U2117 (N_2117,In_4,In_537);
nand U2118 (N_2118,In_264,In_100);
nand U2119 (N_2119,In_812,In_278);
nand U2120 (N_2120,In_930,In_99);
nor U2121 (N_2121,In_651,In_518);
nand U2122 (N_2122,In_1,In_678);
and U2123 (N_2123,In_584,In_109);
or U2124 (N_2124,In_584,In_695);
nand U2125 (N_2125,In_491,In_99);
nand U2126 (N_2126,In_843,In_976);
or U2127 (N_2127,In_185,In_949);
or U2128 (N_2128,In_839,In_358);
and U2129 (N_2129,In_698,In_186);
nand U2130 (N_2130,In_4,In_354);
and U2131 (N_2131,In_83,In_781);
or U2132 (N_2132,In_810,In_492);
or U2133 (N_2133,In_830,In_565);
nor U2134 (N_2134,In_609,In_232);
or U2135 (N_2135,In_758,In_458);
nand U2136 (N_2136,In_801,In_31);
nor U2137 (N_2137,In_611,In_400);
and U2138 (N_2138,In_640,In_582);
nand U2139 (N_2139,In_414,In_758);
nor U2140 (N_2140,In_748,In_678);
xnor U2141 (N_2141,In_11,In_927);
and U2142 (N_2142,In_319,In_986);
nor U2143 (N_2143,In_107,In_375);
nor U2144 (N_2144,In_969,In_715);
and U2145 (N_2145,In_711,In_640);
and U2146 (N_2146,In_654,In_872);
and U2147 (N_2147,In_831,In_27);
nor U2148 (N_2148,In_171,In_909);
nor U2149 (N_2149,In_783,In_330);
nor U2150 (N_2150,In_974,In_195);
and U2151 (N_2151,In_330,In_325);
and U2152 (N_2152,In_388,In_630);
nor U2153 (N_2153,In_707,In_681);
nor U2154 (N_2154,In_818,In_568);
or U2155 (N_2155,In_485,In_799);
nor U2156 (N_2156,In_110,In_613);
xor U2157 (N_2157,In_494,In_384);
nand U2158 (N_2158,In_496,In_868);
nand U2159 (N_2159,In_567,In_263);
nor U2160 (N_2160,In_247,In_166);
and U2161 (N_2161,In_756,In_494);
nor U2162 (N_2162,In_91,In_146);
xnor U2163 (N_2163,In_470,In_614);
nor U2164 (N_2164,In_754,In_38);
and U2165 (N_2165,In_691,In_532);
or U2166 (N_2166,In_622,In_389);
and U2167 (N_2167,In_523,In_328);
nand U2168 (N_2168,In_739,In_526);
nor U2169 (N_2169,In_913,In_196);
nor U2170 (N_2170,In_512,In_280);
and U2171 (N_2171,In_816,In_138);
or U2172 (N_2172,In_27,In_678);
xor U2173 (N_2173,In_863,In_598);
or U2174 (N_2174,In_560,In_557);
and U2175 (N_2175,In_123,In_239);
or U2176 (N_2176,In_974,In_309);
or U2177 (N_2177,In_710,In_810);
nand U2178 (N_2178,In_259,In_934);
nand U2179 (N_2179,In_842,In_956);
nand U2180 (N_2180,In_549,In_360);
nand U2181 (N_2181,In_223,In_768);
xnor U2182 (N_2182,In_434,In_13);
nor U2183 (N_2183,In_377,In_11);
nor U2184 (N_2184,In_885,In_616);
and U2185 (N_2185,In_472,In_342);
nand U2186 (N_2186,In_145,In_247);
nor U2187 (N_2187,In_130,In_765);
and U2188 (N_2188,In_651,In_840);
or U2189 (N_2189,In_602,In_689);
nand U2190 (N_2190,In_36,In_268);
and U2191 (N_2191,In_494,In_690);
nor U2192 (N_2192,In_719,In_194);
nor U2193 (N_2193,In_694,In_885);
or U2194 (N_2194,In_88,In_333);
xnor U2195 (N_2195,In_12,In_271);
nand U2196 (N_2196,In_4,In_754);
nor U2197 (N_2197,In_578,In_409);
nand U2198 (N_2198,In_13,In_855);
xor U2199 (N_2199,In_456,In_487);
and U2200 (N_2200,In_89,In_207);
and U2201 (N_2201,In_34,In_195);
nor U2202 (N_2202,In_332,In_322);
nand U2203 (N_2203,In_437,In_746);
or U2204 (N_2204,In_338,In_774);
or U2205 (N_2205,In_766,In_993);
or U2206 (N_2206,In_449,In_585);
nor U2207 (N_2207,In_640,In_919);
and U2208 (N_2208,In_448,In_602);
and U2209 (N_2209,In_127,In_559);
nor U2210 (N_2210,In_779,In_670);
or U2211 (N_2211,In_582,In_401);
nor U2212 (N_2212,In_799,In_214);
nor U2213 (N_2213,In_727,In_133);
and U2214 (N_2214,In_979,In_593);
or U2215 (N_2215,In_501,In_319);
or U2216 (N_2216,In_122,In_207);
and U2217 (N_2217,In_552,In_897);
nor U2218 (N_2218,In_966,In_619);
nor U2219 (N_2219,In_145,In_262);
and U2220 (N_2220,In_883,In_156);
nand U2221 (N_2221,In_233,In_343);
nor U2222 (N_2222,In_980,In_208);
and U2223 (N_2223,In_170,In_749);
or U2224 (N_2224,In_482,In_232);
nor U2225 (N_2225,In_823,In_227);
nor U2226 (N_2226,In_579,In_577);
nand U2227 (N_2227,In_815,In_357);
xnor U2228 (N_2228,In_59,In_204);
and U2229 (N_2229,In_462,In_133);
and U2230 (N_2230,In_287,In_635);
nand U2231 (N_2231,In_583,In_22);
nor U2232 (N_2232,In_171,In_119);
and U2233 (N_2233,In_799,In_838);
nor U2234 (N_2234,In_921,In_785);
nand U2235 (N_2235,In_396,In_973);
nor U2236 (N_2236,In_16,In_82);
nor U2237 (N_2237,In_985,In_427);
nand U2238 (N_2238,In_59,In_735);
nand U2239 (N_2239,In_552,In_45);
or U2240 (N_2240,In_909,In_203);
nor U2241 (N_2241,In_113,In_941);
and U2242 (N_2242,In_77,In_762);
nand U2243 (N_2243,In_740,In_35);
or U2244 (N_2244,In_32,In_276);
nor U2245 (N_2245,In_306,In_863);
nor U2246 (N_2246,In_523,In_503);
and U2247 (N_2247,In_143,In_564);
and U2248 (N_2248,In_17,In_987);
xnor U2249 (N_2249,In_340,In_254);
nor U2250 (N_2250,In_772,In_312);
and U2251 (N_2251,In_684,In_823);
nand U2252 (N_2252,In_555,In_785);
nor U2253 (N_2253,In_884,In_763);
and U2254 (N_2254,In_303,In_174);
or U2255 (N_2255,In_215,In_870);
or U2256 (N_2256,In_720,In_245);
nand U2257 (N_2257,In_359,In_479);
and U2258 (N_2258,In_120,In_307);
nand U2259 (N_2259,In_262,In_674);
or U2260 (N_2260,In_789,In_778);
nand U2261 (N_2261,In_344,In_695);
nand U2262 (N_2262,In_427,In_831);
nor U2263 (N_2263,In_691,In_674);
or U2264 (N_2264,In_185,In_552);
or U2265 (N_2265,In_570,In_382);
nand U2266 (N_2266,In_364,In_287);
nand U2267 (N_2267,In_390,In_573);
nand U2268 (N_2268,In_560,In_401);
nor U2269 (N_2269,In_499,In_327);
or U2270 (N_2270,In_453,In_547);
nand U2271 (N_2271,In_757,In_545);
xor U2272 (N_2272,In_662,In_596);
nand U2273 (N_2273,In_195,In_304);
and U2274 (N_2274,In_528,In_620);
or U2275 (N_2275,In_213,In_875);
xnor U2276 (N_2276,In_965,In_437);
and U2277 (N_2277,In_187,In_797);
nor U2278 (N_2278,In_45,In_879);
and U2279 (N_2279,In_530,In_350);
or U2280 (N_2280,In_368,In_293);
or U2281 (N_2281,In_131,In_683);
nand U2282 (N_2282,In_661,In_625);
nand U2283 (N_2283,In_603,In_702);
and U2284 (N_2284,In_119,In_451);
nand U2285 (N_2285,In_639,In_476);
nor U2286 (N_2286,In_270,In_429);
xor U2287 (N_2287,In_313,In_23);
nor U2288 (N_2288,In_412,In_278);
and U2289 (N_2289,In_149,In_967);
or U2290 (N_2290,In_762,In_51);
nor U2291 (N_2291,In_394,In_470);
nand U2292 (N_2292,In_565,In_646);
or U2293 (N_2293,In_970,In_425);
nor U2294 (N_2294,In_513,In_329);
and U2295 (N_2295,In_353,In_641);
nand U2296 (N_2296,In_105,In_237);
nor U2297 (N_2297,In_163,In_919);
nand U2298 (N_2298,In_969,In_516);
nor U2299 (N_2299,In_315,In_562);
nor U2300 (N_2300,In_890,In_341);
nand U2301 (N_2301,In_848,In_538);
and U2302 (N_2302,In_209,In_321);
nor U2303 (N_2303,In_646,In_85);
and U2304 (N_2304,In_654,In_621);
or U2305 (N_2305,In_608,In_290);
and U2306 (N_2306,In_212,In_418);
xor U2307 (N_2307,In_831,In_801);
and U2308 (N_2308,In_695,In_574);
or U2309 (N_2309,In_952,In_460);
or U2310 (N_2310,In_655,In_704);
and U2311 (N_2311,In_680,In_345);
nand U2312 (N_2312,In_840,In_989);
nor U2313 (N_2313,In_606,In_333);
nand U2314 (N_2314,In_661,In_275);
nand U2315 (N_2315,In_391,In_476);
nand U2316 (N_2316,In_197,In_290);
nand U2317 (N_2317,In_756,In_882);
nand U2318 (N_2318,In_452,In_346);
or U2319 (N_2319,In_98,In_125);
nand U2320 (N_2320,In_796,In_39);
or U2321 (N_2321,In_953,In_124);
or U2322 (N_2322,In_653,In_525);
xnor U2323 (N_2323,In_398,In_745);
or U2324 (N_2324,In_978,In_899);
nand U2325 (N_2325,In_653,In_304);
nand U2326 (N_2326,In_556,In_87);
nand U2327 (N_2327,In_992,In_187);
or U2328 (N_2328,In_854,In_748);
and U2329 (N_2329,In_200,In_675);
and U2330 (N_2330,In_972,In_457);
or U2331 (N_2331,In_537,In_288);
xnor U2332 (N_2332,In_703,In_192);
and U2333 (N_2333,In_721,In_334);
or U2334 (N_2334,In_422,In_522);
nand U2335 (N_2335,In_623,In_499);
nand U2336 (N_2336,In_734,In_861);
nor U2337 (N_2337,In_145,In_591);
xor U2338 (N_2338,In_754,In_324);
nand U2339 (N_2339,In_79,In_631);
nor U2340 (N_2340,In_100,In_426);
nand U2341 (N_2341,In_402,In_746);
xor U2342 (N_2342,In_335,In_249);
and U2343 (N_2343,In_113,In_388);
or U2344 (N_2344,In_581,In_902);
nand U2345 (N_2345,In_379,In_539);
nand U2346 (N_2346,In_15,In_118);
nand U2347 (N_2347,In_880,In_379);
nand U2348 (N_2348,In_64,In_463);
nand U2349 (N_2349,In_147,In_491);
nor U2350 (N_2350,In_767,In_154);
nor U2351 (N_2351,In_934,In_402);
and U2352 (N_2352,In_223,In_406);
nor U2353 (N_2353,In_991,In_160);
or U2354 (N_2354,In_305,In_206);
and U2355 (N_2355,In_322,In_109);
nand U2356 (N_2356,In_889,In_457);
nand U2357 (N_2357,In_950,In_931);
xnor U2358 (N_2358,In_940,In_691);
or U2359 (N_2359,In_194,In_166);
nor U2360 (N_2360,In_223,In_327);
nand U2361 (N_2361,In_701,In_370);
or U2362 (N_2362,In_171,In_323);
xor U2363 (N_2363,In_429,In_281);
and U2364 (N_2364,In_703,In_683);
nor U2365 (N_2365,In_478,In_65);
and U2366 (N_2366,In_123,In_599);
nand U2367 (N_2367,In_260,In_422);
nor U2368 (N_2368,In_189,In_311);
and U2369 (N_2369,In_364,In_294);
or U2370 (N_2370,In_122,In_365);
xnor U2371 (N_2371,In_809,In_815);
xnor U2372 (N_2372,In_336,In_20);
or U2373 (N_2373,In_84,In_912);
or U2374 (N_2374,In_537,In_888);
and U2375 (N_2375,In_650,In_396);
or U2376 (N_2376,In_390,In_222);
and U2377 (N_2377,In_357,In_228);
or U2378 (N_2378,In_229,In_872);
or U2379 (N_2379,In_967,In_609);
nor U2380 (N_2380,In_433,In_378);
nand U2381 (N_2381,In_985,In_193);
or U2382 (N_2382,In_35,In_403);
nand U2383 (N_2383,In_361,In_258);
and U2384 (N_2384,In_593,In_320);
and U2385 (N_2385,In_297,In_649);
nor U2386 (N_2386,In_199,In_120);
and U2387 (N_2387,In_391,In_291);
nor U2388 (N_2388,In_432,In_607);
and U2389 (N_2389,In_939,In_856);
nand U2390 (N_2390,In_371,In_88);
nor U2391 (N_2391,In_404,In_22);
or U2392 (N_2392,In_302,In_775);
nand U2393 (N_2393,In_314,In_711);
nand U2394 (N_2394,In_778,In_408);
nor U2395 (N_2395,In_762,In_227);
or U2396 (N_2396,In_881,In_490);
and U2397 (N_2397,In_811,In_427);
and U2398 (N_2398,In_910,In_876);
and U2399 (N_2399,In_928,In_627);
xor U2400 (N_2400,In_845,In_774);
and U2401 (N_2401,In_926,In_570);
nand U2402 (N_2402,In_279,In_229);
nand U2403 (N_2403,In_298,In_335);
nand U2404 (N_2404,In_260,In_506);
or U2405 (N_2405,In_657,In_548);
nand U2406 (N_2406,In_15,In_127);
xnor U2407 (N_2407,In_488,In_432);
nand U2408 (N_2408,In_794,In_254);
and U2409 (N_2409,In_374,In_962);
and U2410 (N_2410,In_931,In_948);
and U2411 (N_2411,In_335,In_233);
nor U2412 (N_2412,In_474,In_707);
nand U2413 (N_2413,In_694,In_985);
nor U2414 (N_2414,In_918,In_24);
and U2415 (N_2415,In_734,In_217);
or U2416 (N_2416,In_299,In_738);
or U2417 (N_2417,In_911,In_522);
or U2418 (N_2418,In_550,In_902);
or U2419 (N_2419,In_236,In_250);
xor U2420 (N_2420,In_21,In_53);
nor U2421 (N_2421,In_184,In_333);
and U2422 (N_2422,In_256,In_226);
nand U2423 (N_2423,In_1,In_183);
nor U2424 (N_2424,In_618,In_894);
and U2425 (N_2425,In_131,In_572);
nor U2426 (N_2426,In_895,In_398);
nand U2427 (N_2427,In_10,In_51);
nand U2428 (N_2428,In_264,In_523);
or U2429 (N_2429,In_546,In_924);
or U2430 (N_2430,In_106,In_740);
or U2431 (N_2431,In_414,In_510);
or U2432 (N_2432,In_314,In_510);
and U2433 (N_2433,In_137,In_298);
and U2434 (N_2434,In_473,In_226);
nor U2435 (N_2435,In_529,In_370);
xor U2436 (N_2436,In_371,In_867);
xnor U2437 (N_2437,In_4,In_321);
xor U2438 (N_2438,In_680,In_951);
nor U2439 (N_2439,In_607,In_899);
nor U2440 (N_2440,In_454,In_591);
or U2441 (N_2441,In_59,In_738);
and U2442 (N_2442,In_825,In_959);
nand U2443 (N_2443,In_28,In_706);
or U2444 (N_2444,In_404,In_220);
xor U2445 (N_2445,In_331,In_210);
and U2446 (N_2446,In_849,In_800);
or U2447 (N_2447,In_828,In_943);
nor U2448 (N_2448,In_840,In_669);
nand U2449 (N_2449,In_495,In_540);
xor U2450 (N_2450,In_239,In_808);
or U2451 (N_2451,In_479,In_499);
and U2452 (N_2452,In_467,In_604);
nor U2453 (N_2453,In_442,In_428);
and U2454 (N_2454,In_121,In_36);
or U2455 (N_2455,In_179,In_759);
nor U2456 (N_2456,In_970,In_755);
and U2457 (N_2457,In_672,In_133);
and U2458 (N_2458,In_971,In_756);
nor U2459 (N_2459,In_230,In_728);
nor U2460 (N_2460,In_60,In_843);
or U2461 (N_2461,In_20,In_27);
nor U2462 (N_2462,In_346,In_721);
or U2463 (N_2463,In_303,In_716);
and U2464 (N_2464,In_694,In_280);
nand U2465 (N_2465,In_335,In_39);
nand U2466 (N_2466,In_841,In_198);
xnor U2467 (N_2467,In_910,In_425);
and U2468 (N_2468,In_575,In_828);
or U2469 (N_2469,In_930,In_591);
nand U2470 (N_2470,In_127,In_973);
nand U2471 (N_2471,In_595,In_489);
nand U2472 (N_2472,In_694,In_222);
or U2473 (N_2473,In_115,In_762);
and U2474 (N_2474,In_883,In_261);
or U2475 (N_2475,In_721,In_367);
xor U2476 (N_2476,In_920,In_740);
and U2477 (N_2477,In_651,In_598);
or U2478 (N_2478,In_870,In_803);
nand U2479 (N_2479,In_199,In_584);
nand U2480 (N_2480,In_785,In_66);
xor U2481 (N_2481,In_629,In_503);
and U2482 (N_2482,In_685,In_324);
nor U2483 (N_2483,In_389,In_336);
and U2484 (N_2484,In_817,In_925);
or U2485 (N_2485,In_698,In_55);
nand U2486 (N_2486,In_682,In_769);
or U2487 (N_2487,In_729,In_57);
or U2488 (N_2488,In_510,In_738);
or U2489 (N_2489,In_104,In_280);
and U2490 (N_2490,In_950,In_594);
and U2491 (N_2491,In_138,In_951);
or U2492 (N_2492,In_997,In_726);
nand U2493 (N_2493,In_869,In_757);
or U2494 (N_2494,In_684,In_548);
and U2495 (N_2495,In_487,In_77);
or U2496 (N_2496,In_705,In_942);
nor U2497 (N_2497,In_28,In_552);
and U2498 (N_2498,In_841,In_318);
nand U2499 (N_2499,In_102,In_513);
or U2500 (N_2500,N_1396,N_2219);
xnor U2501 (N_2501,N_841,N_166);
nand U2502 (N_2502,N_908,N_2388);
or U2503 (N_2503,N_1828,N_2231);
nor U2504 (N_2504,N_1203,N_2435);
and U2505 (N_2505,N_1504,N_1322);
nand U2506 (N_2506,N_92,N_950);
nor U2507 (N_2507,N_832,N_84);
xor U2508 (N_2508,N_1569,N_207);
and U2509 (N_2509,N_102,N_1669);
xnor U2510 (N_2510,N_1318,N_251);
nor U2511 (N_2511,N_2122,N_419);
and U2512 (N_2512,N_1999,N_461);
and U2513 (N_2513,N_354,N_75);
nor U2514 (N_2514,N_107,N_663);
nor U2515 (N_2515,N_564,N_399);
nand U2516 (N_2516,N_239,N_934);
and U2517 (N_2517,N_662,N_1502);
and U2518 (N_2518,N_1503,N_516);
or U2519 (N_2519,N_1297,N_2112);
nor U2520 (N_2520,N_1264,N_2434);
nand U2521 (N_2521,N_1973,N_2205);
or U2522 (N_2522,N_121,N_1236);
xnor U2523 (N_2523,N_1710,N_1283);
and U2524 (N_2524,N_1085,N_1523);
and U2525 (N_2525,N_1323,N_1935);
nor U2526 (N_2526,N_2255,N_275);
nand U2527 (N_2527,N_1694,N_476);
nand U2528 (N_2528,N_1703,N_729);
and U2529 (N_2529,N_2496,N_1276);
or U2530 (N_2530,N_271,N_1905);
nand U2531 (N_2531,N_1632,N_1863);
or U2532 (N_2532,N_1348,N_2004);
or U2533 (N_2533,N_890,N_1723);
nand U2534 (N_2534,N_1631,N_1361);
and U2535 (N_2535,N_1280,N_2428);
or U2536 (N_2536,N_465,N_714);
nor U2537 (N_2537,N_853,N_792);
or U2538 (N_2538,N_1540,N_2287);
nor U2539 (N_2539,N_1803,N_546);
nor U2540 (N_2540,N_835,N_308);
xnor U2541 (N_2541,N_1653,N_816);
xnor U2542 (N_2542,N_2081,N_1417);
and U2543 (N_2543,N_2348,N_535);
or U2544 (N_2544,N_919,N_109);
nor U2545 (N_2545,N_1613,N_2313);
nand U2546 (N_2546,N_2281,N_254);
and U2547 (N_2547,N_1445,N_1518);
or U2548 (N_2548,N_1759,N_2245);
or U2549 (N_2549,N_263,N_2354);
or U2550 (N_2550,N_1096,N_2389);
nand U2551 (N_2551,N_1375,N_805);
and U2552 (N_2552,N_1994,N_2054);
nand U2553 (N_2553,N_1598,N_1215);
or U2554 (N_2554,N_2183,N_397);
nor U2555 (N_2555,N_1897,N_1146);
or U2556 (N_2556,N_101,N_2096);
nor U2557 (N_2557,N_1906,N_650);
nor U2558 (N_2558,N_1367,N_1350);
xnor U2559 (N_2559,N_1550,N_660);
or U2560 (N_2560,N_15,N_1861);
nor U2561 (N_2561,N_1692,N_133);
nand U2562 (N_2562,N_2184,N_1953);
nor U2563 (N_2563,N_1910,N_2468);
and U2564 (N_2564,N_1822,N_1337);
nand U2565 (N_2565,N_2003,N_2429);
xnor U2566 (N_2566,N_1381,N_1729);
nor U2567 (N_2567,N_1516,N_1624);
nand U2568 (N_2568,N_2252,N_621);
or U2569 (N_2569,N_356,N_2253);
and U2570 (N_2570,N_1791,N_149);
and U2571 (N_2571,N_2375,N_61);
nor U2572 (N_2572,N_2346,N_603);
and U2573 (N_2573,N_1011,N_2393);
nand U2574 (N_2574,N_1434,N_1988);
and U2575 (N_2575,N_1244,N_1036);
nor U2576 (N_2576,N_1886,N_1545);
nand U2577 (N_2577,N_2075,N_1431);
and U2578 (N_2578,N_1577,N_768);
nand U2579 (N_2579,N_763,N_144);
or U2580 (N_2580,N_1878,N_1940);
nor U2581 (N_2581,N_2339,N_407);
nand U2582 (N_2582,N_2444,N_1553);
nor U2583 (N_2583,N_2022,N_1104);
or U2584 (N_2584,N_1709,N_1533);
or U2585 (N_2585,N_1529,N_180);
nand U2586 (N_2586,N_2335,N_2325);
xor U2587 (N_2587,N_1904,N_2203);
nand U2588 (N_2588,N_1730,N_846);
nand U2589 (N_2589,N_1854,N_754);
nor U2590 (N_2590,N_2316,N_1450);
nor U2591 (N_2591,N_2030,N_917);
or U2592 (N_2592,N_920,N_57);
nor U2593 (N_2593,N_2074,N_173);
nor U2594 (N_2594,N_1483,N_1301);
nand U2595 (N_2595,N_1734,N_624);
xnor U2596 (N_2596,N_1595,N_2297);
xor U2597 (N_2597,N_800,N_795);
nor U2598 (N_2598,N_30,N_1981);
nor U2599 (N_2599,N_775,N_866);
and U2600 (N_2600,N_2083,N_2194);
nand U2601 (N_2601,N_1138,N_1415);
and U2602 (N_2602,N_2362,N_376);
and U2603 (N_2603,N_1900,N_319);
nor U2604 (N_2604,N_563,N_1118);
or U2605 (N_2605,N_616,N_1616);
or U2606 (N_2606,N_2187,N_1333);
xnor U2607 (N_2607,N_1064,N_304);
or U2608 (N_2608,N_979,N_830);
nand U2609 (N_2609,N_2498,N_11);
or U2610 (N_2610,N_2251,N_484);
nand U2611 (N_2611,N_1461,N_868);
nor U2612 (N_2612,N_18,N_683);
and U2613 (N_2613,N_371,N_478);
and U2614 (N_2614,N_2300,N_470);
nor U2615 (N_2615,N_2410,N_987);
nor U2616 (N_2616,N_1050,N_786);
nand U2617 (N_2617,N_1401,N_1979);
xnor U2618 (N_2618,N_163,N_1630);
and U2619 (N_2619,N_1660,N_2403);
nand U2620 (N_2620,N_441,N_76);
or U2621 (N_2621,N_241,N_274);
nor U2622 (N_2622,N_1066,N_2053);
nand U2623 (N_2623,N_1095,N_691);
nand U2624 (N_2624,N_1419,N_2177);
and U2625 (N_2625,N_1026,N_1629);
nand U2626 (N_2626,N_2132,N_580);
nand U2627 (N_2627,N_1558,N_448);
or U2628 (N_2628,N_2180,N_871);
nor U2629 (N_2629,N_1058,N_1365);
or U2630 (N_2630,N_1115,N_436);
nand U2631 (N_2631,N_1342,N_1758);
nor U2632 (N_2632,N_588,N_1737);
and U2633 (N_2633,N_248,N_2036);
nand U2634 (N_2634,N_1037,N_153);
nor U2635 (N_2635,N_688,N_31);
and U2636 (N_2636,N_1738,N_556);
and U2637 (N_2637,N_2282,N_433);
xnor U2638 (N_2638,N_424,N_422);
and U2639 (N_2639,N_384,N_1527);
nand U2640 (N_2640,N_1475,N_1054);
or U2641 (N_2641,N_391,N_992);
nand U2642 (N_2642,N_1801,N_730);
or U2643 (N_2643,N_492,N_1986);
xor U2644 (N_2644,N_396,N_209);
or U2645 (N_2645,N_472,N_678);
and U2646 (N_2646,N_825,N_1284);
nand U2647 (N_2647,N_996,N_342);
nand U2648 (N_2648,N_1290,N_2499);
xnor U2649 (N_2649,N_286,N_625);
xnor U2650 (N_2650,N_454,N_1373);
xnor U2651 (N_2651,N_1573,N_1427);
nand U2652 (N_2652,N_1741,N_2414);
nor U2653 (N_2653,N_669,N_2303);
nor U2654 (N_2654,N_1884,N_1772);
xnor U2655 (N_2655,N_1046,N_2064);
nor U2656 (N_2656,N_734,N_1153);
nor U2657 (N_2657,N_45,N_639);
xnor U2658 (N_2658,N_400,N_1038);
or U2659 (N_2659,N_1536,N_883);
nand U2660 (N_2660,N_2484,N_2065);
xor U2661 (N_2661,N_157,N_1622);
and U2662 (N_2662,N_976,N_970);
nor U2663 (N_2663,N_609,N_781);
nand U2664 (N_2664,N_867,N_1699);
or U2665 (N_2665,N_1198,N_2280);
nor U2666 (N_2666,N_1499,N_1877);
or U2667 (N_2667,N_2438,N_674);
or U2668 (N_2668,N_44,N_591);
nand U2669 (N_2669,N_320,N_2350);
or U2670 (N_2670,N_115,N_412);
nand U2671 (N_2671,N_1921,N_1248);
xnor U2672 (N_2672,N_265,N_1552);
nand U2673 (N_2673,N_2246,N_1874);
and U2674 (N_2674,N_764,N_2491);
and U2675 (N_2675,N_2012,N_221);
nand U2676 (N_2676,N_2050,N_2174);
xnor U2677 (N_2677,N_904,N_1336);
and U2678 (N_2678,N_2480,N_42);
and U2679 (N_2679,N_925,N_205);
nor U2680 (N_2680,N_2199,N_2033);
or U2681 (N_2681,N_1689,N_2411);
or U2682 (N_2682,N_502,N_2150);
and U2683 (N_2683,N_935,N_1390);
or U2684 (N_2684,N_2148,N_1209);
nor U2685 (N_2685,N_287,N_949);
xor U2686 (N_2686,N_1469,N_1343);
nand U2687 (N_2687,N_1376,N_1834);
and U2688 (N_2688,N_2059,N_1857);
nand U2689 (N_2689,N_607,N_1785);
nand U2690 (N_2690,N_2018,N_242);
nor U2691 (N_2691,N_833,N_1128);
or U2692 (N_2692,N_962,N_2138);
and U2693 (N_2693,N_1915,N_716);
nand U2694 (N_2694,N_713,N_573);
nand U2695 (N_2695,N_2320,N_2170);
and U2696 (N_2696,N_2493,N_2417);
or U2697 (N_2697,N_2242,N_2326);
and U2698 (N_2698,N_208,N_493);
xnor U2699 (N_2699,N_743,N_1426);
nand U2700 (N_2700,N_684,N_26);
or U2701 (N_2701,N_1459,N_848);
nand U2702 (N_2702,N_1964,N_2043);
nand U2703 (N_2703,N_40,N_1161);
and U2704 (N_2704,N_105,N_1141);
nand U2705 (N_2705,N_77,N_175);
nand U2706 (N_2706,N_374,N_1812);
nor U2707 (N_2707,N_1928,N_24);
and U2708 (N_2708,N_1938,N_1195);
xnor U2709 (N_2709,N_330,N_2309);
or U2710 (N_2710,N_485,N_1982);
or U2711 (N_2711,N_145,N_395);
nor U2712 (N_2712,N_2135,N_51);
and U2713 (N_2713,N_757,N_328);
nor U2714 (N_2714,N_587,N_1090);
nand U2715 (N_2715,N_537,N_1142);
and U2716 (N_2716,N_554,N_916);
xor U2717 (N_2717,N_1420,N_341);
nand U2718 (N_2718,N_1867,N_827);
and U2719 (N_2719,N_652,N_2475);
nor U2720 (N_2720,N_2085,N_893);
or U2721 (N_2721,N_682,N_295);
xor U2722 (N_2722,N_1230,N_1509);
nor U2723 (N_2723,N_106,N_2229);
and U2724 (N_2724,N_1654,N_1351);
nand U2725 (N_2725,N_2164,N_948);
or U2726 (N_2726,N_1512,N_23);
and U2727 (N_2727,N_2159,N_467);
nand U2728 (N_2728,N_566,N_1073);
nor U2729 (N_2729,N_323,N_2178);
nor U2730 (N_2730,N_2204,N_301);
and U2731 (N_2731,N_820,N_194);
and U2732 (N_2732,N_1313,N_2146);
nand U2733 (N_2733,N_110,N_1658);
or U2734 (N_2734,N_708,N_788);
or U2735 (N_2735,N_2017,N_428);
nand U2736 (N_2736,N_94,N_2477);
nor U2737 (N_2737,N_1392,N_1926);
and U2738 (N_2738,N_791,N_2042);
xnor U2739 (N_2739,N_528,N_93);
or U2740 (N_2740,N_629,N_95);
and U2741 (N_2741,N_1505,N_1978);
or U2742 (N_2742,N_363,N_936);
or U2743 (N_2743,N_2295,N_722);
and U2744 (N_2744,N_1476,N_1651);
and U2745 (N_2745,N_601,N_469);
nor U2746 (N_2746,N_1133,N_1934);
nand U2747 (N_2747,N_879,N_2118);
or U2748 (N_2748,N_1646,N_338);
and U2749 (N_2749,N_1438,N_2176);
nand U2750 (N_2750,N_872,N_47);
and U2751 (N_2751,N_1633,N_2386);
and U2752 (N_2752,N_331,N_1384);
and U2753 (N_2753,N_2436,N_1970);
and U2754 (N_2754,N_733,N_1186);
or U2755 (N_2755,N_1676,N_2190);
nand U2756 (N_2756,N_1102,N_2091);
nor U2757 (N_2757,N_1300,N_1454);
nor U2758 (N_2758,N_1468,N_168);
and U2759 (N_2759,N_269,N_728);
and U2760 (N_2760,N_1247,N_303);
or U2761 (N_2761,N_1876,N_1017);
nor U2762 (N_2762,N_1131,N_553);
or U2763 (N_2763,N_522,N_531);
and U2764 (N_2764,N_1293,N_1241);
and U2765 (N_2765,N_316,N_513);
nand U2766 (N_2766,N_515,N_1566);
nor U2767 (N_2767,N_2472,N_1164);
or U2768 (N_2768,N_353,N_1991);
nor U2769 (N_2769,N_690,N_1787);
nor U2770 (N_2770,N_1289,N_1793);
or U2771 (N_2771,N_1072,N_1391);
or U2772 (N_2772,N_246,N_1757);
and U2773 (N_2773,N_711,N_809);
nor U2774 (N_2774,N_2430,N_545);
nand U2775 (N_2775,N_1299,N_1189);
nand U2776 (N_2776,N_1647,N_1845);
xor U2777 (N_2777,N_1923,N_1020);
nand U2778 (N_2778,N_235,N_2358);
nor U2779 (N_2779,N_2328,N_794);
nor U2780 (N_2780,N_912,N_847);
or U2781 (N_2781,N_1196,N_1081);
and U2782 (N_2782,N_514,N_1794);
or U2783 (N_2783,N_1188,N_1178);
or U2784 (N_2784,N_1500,N_642);
nor U2785 (N_2785,N_2378,N_2031);
nand U2786 (N_2786,N_1025,N_1267);
and U2787 (N_2787,N_1868,N_372);
or U2788 (N_2788,N_1029,N_118);
and U2789 (N_2789,N_410,N_2001);
nand U2790 (N_2790,N_1539,N_48);
nor U2791 (N_2791,N_2024,N_785);
xor U2792 (N_2792,N_1948,N_406);
nor U2793 (N_2793,N_79,N_1548);
and U2794 (N_2794,N_2084,N_946);
or U2795 (N_2795,N_1399,N_704);
and U2796 (N_2796,N_900,N_598);
or U2797 (N_2797,N_736,N_1958);
and U2798 (N_2798,N_193,N_1374);
nand U2799 (N_2799,N_1329,N_2243);
or U2800 (N_2800,N_1274,N_2010);
nor U2801 (N_2801,N_905,N_1060);
nor U2802 (N_2802,N_124,N_2175);
or U2803 (N_2803,N_2158,N_2342);
and U2804 (N_2804,N_631,N_1407);
and U2805 (N_2805,N_2363,N_1259);
and U2806 (N_2806,N_2140,N_1465);
or U2807 (N_2807,N_2236,N_1722);
nand U2808 (N_2808,N_2171,N_2329);
nor U2809 (N_2809,N_1895,N_1298);
nor U2810 (N_2810,N_653,N_2123);
xnor U2811 (N_2811,N_2109,N_1514);
nor U2812 (N_2812,N_1767,N_901);
nor U2813 (N_2813,N_2056,N_252);
or U2814 (N_2814,N_599,N_725);
nor U2815 (N_2815,N_2294,N_1177);
nand U2816 (N_2816,N_2323,N_1311);
nand U2817 (N_2817,N_1588,N_2361);
nor U2818 (N_2818,N_80,N_783);
xnor U2819 (N_2819,N_2424,N_726);
xnor U2820 (N_2820,N_855,N_2293);
xor U2821 (N_2821,N_1668,N_1009);
and U2822 (N_2822,N_96,N_1602);
nor U2823 (N_2823,N_765,N_1466);
nor U2824 (N_2824,N_20,N_709);
or U2825 (N_2825,N_226,N_2374);
xor U2826 (N_2826,N_140,N_2037);
nor U2827 (N_2827,N_444,N_244);
and U2828 (N_2828,N_1262,N_2366);
nand U2829 (N_2829,N_2088,N_2100);
and U2830 (N_2830,N_471,N_1605);
nor U2831 (N_2831,N_2395,N_2008);
or U2832 (N_2832,N_1010,N_1253);
and U2833 (N_2833,N_1510,N_2306);
or U2834 (N_2834,N_1478,N_1043);
nor U2835 (N_2835,N_561,N_322);
or U2836 (N_2836,N_1252,N_750);
and U2837 (N_2837,N_1261,N_1082);
nor U2838 (N_2838,N_658,N_62);
or U2839 (N_2839,N_388,N_1725);
nand U2840 (N_2840,N_2057,N_499);
and U2841 (N_2841,N_1429,N_1447);
or U2842 (N_2842,N_926,N_1652);
or U2843 (N_2843,N_1893,N_2299);
or U2844 (N_2844,N_686,N_8);
nand U2845 (N_2845,N_2239,N_612);
xor U2846 (N_2846,N_1184,N_1482);
xnor U2847 (N_2847,N_2283,N_1600);
nand U2848 (N_2848,N_2248,N_1670);
and U2849 (N_2849,N_2097,N_280);
and U2850 (N_2850,N_993,N_1966);
nor U2851 (N_2851,N_2298,N_706);
nor U2852 (N_2852,N_865,N_21);
nand U2853 (N_2853,N_318,N_1170);
or U2854 (N_2854,N_745,N_2029);
and U2855 (N_2855,N_2355,N_2360);
nor U2856 (N_2856,N_1719,N_1712);
and U2857 (N_2857,N_258,N_2278);
xor U2858 (N_2858,N_1976,N_1077);
and U2859 (N_2859,N_954,N_2167);
xor U2860 (N_2860,N_1818,N_1040);
or U2861 (N_2861,N_132,N_1349);
and U2862 (N_2862,N_52,N_270);
xnor U2863 (N_2863,N_1380,N_1798);
and U2864 (N_2864,N_789,N_1062);
nand U2865 (N_2865,N_2021,N_468);
nand U2866 (N_2866,N_877,N_243);
xor U2867 (N_2867,N_1696,N_1368);
and U2868 (N_2868,N_426,N_2489);
or U2869 (N_2869,N_2381,N_1557);
nor U2870 (N_2870,N_2291,N_411);
xor U2871 (N_2871,N_125,N_146);
nor U2872 (N_2872,N_2090,N_2071);
or U2873 (N_2873,N_771,N_2086);
and U2874 (N_2874,N_1693,N_2347);
nor U2875 (N_2875,N_2222,N_1603);
nand U2876 (N_2876,N_198,N_1615);
nand U2877 (N_2877,N_481,N_869);
nor U2878 (N_2878,N_628,N_532);
nand U2879 (N_2879,N_2206,N_2353);
or U2880 (N_2880,N_1339,N_136);
or U2881 (N_2881,N_2212,N_1372);
xor U2882 (N_2882,N_2377,N_2332);
xnor U2883 (N_2883,N_1113,N_332);
nand U2884 (N_2884,N_863,N_790);
and U2885 (N_2885,N_1789,N_681);
nand U2886 (N_2886,N_483,N_1835);
xnor U2887 (N_2887,N_1051,N_1152);
nor U2888 (N_2888,N_2481,N_336);
nor U2889 (N_2889,N_358,N_1258);
or U2890 (N_2890,N_654,N_55);
and U2891 (N_2891,N_1614,N_1139);
nor U2892 (N_2892,N_2139,N_1012);
or U2893 (N_2893,N_1838,N_1007);
and U2894 (N_2894,N_1357,N_1508);
nand U2895 (N_2895,N_517,N_1853);
nor U2896 (N_2896,N_2216,N_891);
nor U2897 (N_2897,N_1858,N_261);
nand U2898 (N_2898,N_1494,N_28);
or U2899 (N_2899,N_309,N_112);
or U2900 (N_2900,N_637,N_2023);
or U2901 (N_2901,N_1150,N_1724);
nand U2902 (N_2902,N_1525,N_2465);
and U2903 (N_2903,N_1872,N_819);
or U2904 (N_2904,N_2483,N_1875);
nand U2905 (N_2905,N_417,N_1987);
nand U2906 (N_2906,N_159,N_1578);
or U2907 (N_2907,N_1059,N_842);
and U2908 (N_2908,N_1522,N_199);
nor U2909 (N_2909,N_590,N_2113);
nor U2910 (N_2910,N_673,N_273);
and U2911 (N_2911,N_447,N_2220);
and U2912 (N_2912,N_1920,N_836);
nand U2913 (N_2913,N_2127,N_2032);
or U2914 (N_2914,N_99,N_521);
nor U2915 (N_2915,N_850,N_355);
xor U2916 (N_2916,N_431,N_558);
and U2917 (N_2917,N_1462,N_928);
xor U2918 (N_2918,N_1456,N_1980);
nor U2919 (N_2919,N_1176,N_1572);
or U2920 (N_2920,N_82,N_456);
nand U2921 (N_2921,N_2224,N_2191);
and U2922 (N_2922,N_782,N_1918);
and U2923 (N_2923,N_60,N_2416);
or U2924 (N_2924,N_2128,N_2440);
nor U2925 (N_2925,N_1996,N_1972);
xor U2926 (N_2926,N_2192,N_1366);
nor U2927 (N_2927,N_873,N_2093);
and U2928 (N_2928,N_984,N_1484);
or U2929 (N_2929,N_2268,N_473);
or U2930 (N_2930,N_364,N_2349);
and U2931 (N_2931,N_2103,N_941);
and U2932 (N_2932,N_1648,N_2455);
nor U2933 (N_2933,N_2409,N_1601);
or U2934 (N_2934,N_1831,N_1288);
and U2935 (N_2935,N_600,N_2060);
and U2936 (N_2936,N_423,N_1044);
nor U2937 (N_2937,N_969,N_1846);
and U2938 (N_2938,N_2382,N_672);
nand U2939 (N_2939,N_1507,N_1852);
nand U2940 (N_2940,N_2145,N_297);
nand U2941 (N_2941,N_2232,N_1753);
nand U2942 (N_2942,N_929,N_1561);
and U2943 (N_2943,N_2413,N_2277);
or U2944 (N_2944,N_1887,N_2172);
nand U2945 (N_2945,N_1477,N_1894);
nor U2946 (N_2946,N_1022,N_1974);
xor U2947 (N_2947,N_347,N_651);
xor U2948 (N_2948,N_1451,N_512);
xnor U2949 (N_2949,N_1400,N_1439);
nor U2950 (N_2950,N_975,N_1591);
nor U2951 (N_2951,N_1819,N_1441);
and U2952 (N_2952,N_2116,N_898);
nor U2953 (N_2953,N_1989,N_1213);
nor U2954 (N_2954,N_307,N_169);
or U2955 (N_2955,N_887,N_740);
or U2956 (N_2956,N_1312,N_1984);
nand U2957 (N_2957,N_2196,N_1049);
nand U2958 (N_2958,N_315,N_488);
xnor U2959 (N_2959,N_416,N_2262);
and U2960 (N_2960,N_1903,N_1830);
nor U2961 (N_2961,N_46,N_1467);
or U2962 (N_2962,N_2379,N_126);
nor U2963 (N_2963,N_365,N_2336);
nor U2964 (N_2964,N_647,N_760);
nor U2965 (N_2965,N_1379,N_302);
nand U2966 (N_2966,N_2331,N_875);
or U2967 (N_2967,N_1815,N_1119);
nor U2968 (N_2968,N_1493,N_1021);
nand U2969 (N_2969,N_870,N_851);
xnor U2970 (N_2970,N_1406,N_1242);
xnor U2971 (N_2971,N_2257,N_340);
or U2972 (N_2972,N_635,N_1107);
nor U2973 (N_2973,N_519,N_755);
and U2974 (N_2974,N_188,N_965);
nand U2975 (N_2975,N_627,N_1216);
and U2976 (N_2976,N_1807,N_2259);
and U2977 (N_2977,N_2406,N_68);
nand U2978 (N_2978,N_747,N_615);
xor U2979 (N_2979,N_1358,N_909);
nand U2980 (N_2980,N_1486,N_1266);
or U2981 (N_2981,N_1316,N_982);
or U2982 (N_2982,N_0,N_1674);
or U2983 (N_2983,N_961,N_1287);
nor U2984 (N_2984,N_1565,N_1187);
nor U2985 (N_2985,N_278,N_695);
and U2986 (N_2986,N_1950,N_1664);
and U2987 (N_2987,N_2476,N_2284);
nand U2988 (N_2988,N_577,N_1464);
nand U2989 (N_2989,N_2225,N_22);
nor U2990 (N_2990,N_1899,N_1820);
and U2991 (N_2991,N_2230,N_1701);
or U2992 (N_2992,N_1394,N_1779);
nand U2993 (N_2993,N_1233,N_1089);
nor U2994 (N_2994,N_2420,N_2423);
and U2995 (N_2995,N_2020,N_606);
nand U2996 (N_2996,N_1795,N_202);
nand U2997 (N_2997,N_2,N_487);
xor U2998 (N_2998,N_1364,N_496);
nor U2999 (N_2999,N_14,N_1555);
or U3000 (N_3000,N_176,N_510);
and U3001 (N_3001,N_390,N_117);
nand U3002 (N_3002,N_834,N_712);
nor U3003 (N_3003,N_1409,N_1382);
nand U3004 (N_3004,N_2398,N_1158);
nor U3005 (N_3005,N_2110,N_1599);
nand U3006 (N_3006,N_1488,N_636);
nand U3007 (N_3007,N_1250,N_4);
xnor U3008 (N_3008,N_1446,N_951);
or U3009 (N_3009,N_325,N_1506);
nor U3010 (N_3010,N_649,N_2399);
and U3011 (N_3011,N_1008,N_379);
or U3012 (N_3012,N_748,N_111);
or U3013 (N_3013,N_277,N_1255);
nand U3014 (N_3014,N_1123,N_958);
or U3015 (N_3015,N_1697,N_583);
nand U3016 (N_3016,N_1960,N_876);
nand U3017 (N_3017,N_2376,N_228);
nor U3018 (N_3018,N_389,N_361);
nand U3019 (N_3019,N_2387,N_2474);
and U3020 (N_3020,N_2357,N_368);
xnor U3021 (N_3021,N_2119,N_229);
nand U3022 (N_3022,N_2047,N_458);
nor U3023 (N_3023,N_2288,N_445);
and U3024 (N_3024,N_2025,N_1797);
nor U3025 (N_3025,N_2391,N_1659);
and U3026 (N_3026,N_1360,N_1519);
or U3027 (N_3027,N_503,N_1747);
nor U3028 (N_3028,N_230,N_858);
and U3029 (N_3029,N_2422,N_120);
or U3030 (N_3030,N_1945,N_1678);
and U3031 (N_3031,N_1781,N_977);
or U3032 (N_3032,N_565,N_1929);
or U3033 (N_3033,N_787,N_1806);
nor U3034 (N_3034,N_1850,N_1035);
nand U3035 (N_3035,N_1571,N_1657);
and U3036 (N_3036,N_482,N_1889);
nor U3037 (N_3037,N_1760,N_2005);
nor U3038 (N_3038,N_1408,N_1776);
nor U3039 (N_3039,N_696,N_86);
and U3040 (N_3040,N_1279,N_25);
nor U3041 (N_3041,N_326,N_1109);
xor U3042 (N_3042,N_2314,N_1080);
or U3043 (N_3043,N_6,N_610);
nand U3044 (N_3044,N_2106,N_2153);
and U3045 (N_3045,N_1637,N_1907);
nor U3046 (N_3046,N_2317,N_2486);
xor U3047 (N_3047,N_2111,N_2421);
nor U3048 (N_3048,N_569,N_418);
nor U3049 (N_3049,N_1922,N_1744);
nand U3050 (N_3050,N_1067,N_1892);
and U3051 (N_3051,N_122,N_192);
and U3052 (N_3052,N_1879,N_2181);
or U3053 (N_3053,N_632,N_1680);
and U3054 (N_3054,N_1901,N_1969);
or U3055 (N_3055,N_386,N_1204);
nor U3056 (N_3056,N_437,N_1655);
nand U3057 (N_3057,N_1695,N_2371);
or U3058 (N_3058,N_414,N_2394);
and U3059 (N_3059,N_1520,N_1665);
and U3060 (N_3060,N_1702,N_2302);
nor U3061 (N_3061,N_387,N_2473);
or U3062 (N_3062,N_1121,N_2142);
or U3063 (N_3063,N_2301,N_1556);
xor U3064 (N_3064,N_1112,N_1028);
nor U3065 (N_3065,N_1265,N_837);
or U3066 (N_3066,N_944,N_643);
nor U3067 (N_3067,N_97,N_1698);
or U3068 (N_3068,N_375,N_1816);
nand U3069 (N_3069,N_679,N_619);
and U3070 (N_3070,N_139,N_1720);
xnor U3071 (N_3071,N_2445,N_1226);
nand U3072 (N_3072,N_1127,N_1933);
nand U3073 (N_3073,N_408,N_1403);
and U3074 (N_3074,N_2055,N_1732);
nand U3075 (N_3075,N_1526,N_994);
nand U3076 (N_3076,N_2451,N_2009);
or U3077 (N_3077,N_81,N_1913);
nor U3078 (N_3078,N_2460,N_2104);
nand U3079 (N_3079,N_1428,N_542);
nor U3080 (N_3080,N_413,N_1814);
nand U3081 (N_3081,N_2208,N_568);
or U3082 (N_3082,N_1786,N_1310);
nand U3083 (N_3083,N_839,N_200);
or U3084 (N_3084,N_2341,N_1625);
xnor U3085 (N_3085,N_2045,N_896);
nand U3086 (N_3086,N_551,N_2210);
or U3087 (N_3087,N_1748,N_1847);
xnor U3088 (N_3088,N_2385,N_2337);
and U3089 (N_3089,N_2099,N_1083);
nor U3090 (N_3090,N_543,N_366);
and U3091 (N_3091,N_699,N_1681);
nand U3092 (N_3092,N_104,N_440);
nor U3093 (N_3093,N_843,N_1015);
nor U3094 (N_3094,N_1930,N_2221);
nor U3095 (N_3095,N_902,N_702);
nor U3096 (N_3096,N_776,N_2040);
xor U3097 (N_3097,N_1157,N_1129);
nand U3098 (N_3098,N_1227,N_1871);
nor U3099 (N_3099,N_710,N_1257);
xor U3100 (N_3100,N_147,N_504);
or U3101 (N_3101,N_1649,N_1330);
or U3102 (N_3102,N_881,N_1335);
nor U3103 (N_3103,N_2497,N_559);
nor U3104 (N_3104,N_214,N_2426);
xor U3105 (N_3105,N_1743,N_2453);
nor U3106 (N_3106,N_780,N_38);
nor U3107 (N_3107,N_1727,N_486);
and U3108 (N_3108,N_623,N_752);
nand U3109 (N_3109,N_58,N_1205);
nor U3110 (N_3110,N_1075,N_1370);
nor U3111 (N_3111,N_256,N_2079);
xnor U3112 (N_3112,N_2443,N_2107);
or U3113 (N_3113,N_818,N_523);
and U3114 (N_3114,N_675,N_2344);
nand U3115 (N_3115,N_224,N_13);
nand U3116 (N_3116,N_1735,N_2163);
or U3117 (N_3117,N_995,N_1355);
nand U3118 (N_3118,N_253,N_1042);
nor U3119 (N_3119,N_1823,N_490);
and U3120 (N_3120,N_885,N_220);
and U3121 (N_3121,N_1345,N_910);
and U3122 (N_3122,N_1517,N_1057);
and U3123 (N_3123,N_1004,N_2405);
or U3124 (N_3124,N_605,N_2401);
xnor U3125 (N_3125,N_1563,N_751);
or U3126 (N_3126,N_1808,N_16);
or U3127 (N_3127,N_43,N_2343);
or U3128 (N_3128,N_1718,N_227);
nor U3129 (N_3129,N_1378,N_2365);
or U3130 (N_3130,N_2141,N_1777);
and U3131 (N_3131,N_327,N_774);
nor U3132 (N_3132,N_940,N_1587);
and U3133 (N_3133,N_291,N_2265);
nor U3134 (N_3134,N_317,N_134);
nor U3135 (N_3135,N_74,N_1841);
or U3136 (N_3136,N_1473,N_1160);
nor U3137 (N_3137,N_1627,N_29);
and U3138 (N_3138,N_2402,N_1685);
nand U3139 (N_3139,N_1746,N_283);
nand U3140 (N_3140,N_1888,N_1386);
and U3141 (N_3141,N_1584,N_9);
nand U3142 (N_3142,N_2241,N_1024);
and U3143 (N_3143,N_184,N_296);
or U3144 (N_3144,N_1640,N_2407);
or U3145 (N_3145,N_1272,N_351);
nand U3146 (N_3146,N_1421,N_945);
nor U3147 (N_3147,N_141,N_172);
xnor U3148 (N_3148,N_1005,N_1639);
or U3149 (N_3149,N_2179,N_1586);
xnor U3150 (N_3150,N_453,N_130);
nor U3151 (N_3151,N_1749,N_2494);
xnor U3152 (N_3152,N_838,N_2272);
and U3153 (N_3153,N_1604,N_533);
or U3154 (N_3154,N_1581,N_1448);
nor U3155 (N_3155,N_335,N_2026);
nor U3156 (N_3156,N_1644,N_50);
nand U3157 (N_3157,N_1489,N_2345);
and U3158 (N_3158,N_1319,N_218);
or U3159 (N_3159,N_1495,N_2067);
nand U3160 (N_3160,N_700,N_1898);
nand U3161 (N_3161,N_1433,N_761);
nand U3162 (N_3162,N_821,N_394);
and U3163 (N_3163,N_592,N_439);
or U3164 (N_3164,N_262,N_2215);
nand U3165 (N_3165,N_1402,N_1137);
nand U3166 (N_3166,N_1078,N_2157);
xor U3167 (N_3167,N_1320,N_1324);
or U3168 (N_3168,N_2290,N_2442);
and U3169 (N_3169,N_2450,N_1544);
xor U3170 (N_3170,N_2396,N_534);
and U3171 (N_3171,N_784,N_1728);
xnor U3172 (N_3172,N_2062,N_1087);
nand U3173 (N_3173,N_2186,N_1034);
or U3174 (N_3174,N_549,N_856);
nor U3175 (N_3175,N_796,N_1105);
nand U3176 (N_3176,N_907,N_1091);
and U3177 (N_3177,N_1612,N_1916);
xnor U3178 (N_3178,N_87,N_802);
xnor U3179 (N_3179,N_1416,N_1890);
or U3180 (N_3180,N_2105,N_2404);
or U3181 (N_3181,N_2425,N_1687);
nor U3182 (N_3182,N_1114,N_1220);
or U3183 (N_3183,N_281,N_849);
and U3184 (N_3184,N_1765,N_2066);
or U3185 (N_3185,N_53,N_1377);
nand U3186 (N_3186,N_2271,N_1610);
and U3187 (N_3187,N_1179,N_1268);
or U3188 (N_3188,N_803,N_756);
nand U3189 (N_3189,N_2319,N_1458);
and U3190 (N_3190,N_1191,N_245);
and U3191 (N_3191,N_1027,N_1745);
and U3192 (N_3192,N_988,N_103);
or U3193 (N_3193,N_334,N_701);
nor U3194 (N_3194,N_1334,N_1848);
or U3195 (N_3195,N_491,N_2495);
nand U3196 (N_3196,N_2213,N_429);
or U3197 (N_3197,N_1155,N_2144);
or U3198 (N_3198,N_1271,N_998);
xor U3199 (N_3199,N_442,N_617);
nor U3200 (N_3200,N_2408,N_581);
and U3201 (N_3201,N_1936,N_1092);
or U3202 (N_3202,N_352,N_1194);
or U3203 (N_3203,N_2463,N_1424);
nand U3204 (N_3204,N_1132,N_1773);
and U3205 (N_3205,N_113,N_718);
nand U3206 (N_3206,N_1688,N_778);
nor U3207 (N_3207,N_1885,N_2035);
nand U3208 (N_3208,N_1623,N_806);
or U3209 (N_3209,N_1766,N_1990);
or U3210 (N_3210,N_446,N_2228);
and U3211 (N_3211,N_2439,N_1711);
xnor U3212 (N_3212,N_2296,N_1663);
nand U3213 (N_3213,N_593,N_1452);
or U3214 (N_3214,N_798,N_255);
and U3215 (N_3215,N_1638,N_1110);
and U3216 (N_3216,N_1911,N_2197);
nand U3217 (N_3217,N_247,N_1750);
or U3218 (N_3218,N_2114,N_947);
nor U3219 (N_3219,N_1097,N_1763);
xnor U3220 (N_3220,N_520,N_586);
nand U3221 (N_3221,N_1873,N_2092);
or U3222 (N_3222,N_2169,N_595);
or U3223 (N_3223,N_644,N_2072);
and U3224 (N_3224,N_161,N_480);
nand U3225 (N_3225,N_1515,N_2256);
and U3226 (N_3226,N_1881,N_1387);
or U3227 (N_3227,N_1956,N_2095);
nor U3228 (N_3228,N_1398,N_1733);
and U3229 (N_3229,N_562,N_2264);
nand U3230 (N_3230,N_2101,N_2115);
or U3231 (N_3231,N_1346,N_434);
or U3232 (N_3232,N_2461,N_801);
and U3233 (N_3233,N_1582,N_1941);
nor U3234 (N_3234,N_1997,N_129);
or U3235 (N_3235,N_614,N_817);
nor U3236 (N_3236,N_2261,N_544);
and U3237 (N_3237,N_1344,N_1325);
nand U3238 (N_3238,N_185,N_420);
nand U3239 (N_3239,N_236,N_1321);
or U3240 (N_3240,N_1173,N_2156);
nand U3241 (N_3241,N_1413,N_1912);
and U3242 (N_3242,N_203,N_88);
nor U3243 (N_3243,N_213,N_813);
or U3244 (N_3244,N_2415,N_311);
xnor U3245 (N_3245,N_739,N_799);
or U3246 (N_3246,N_1751,N_1144);
or U3247 (N_3247,N_217,N_972);
and U3248 (N_3248,N_1388,N_2244);
and U3249 (N_3249,N_73,N_459);
nand U3250 (N_3250,N_234,N_611);
nor U3251 (N_3251,N_1116,N_1780);
nor U3252 (N_3252,N_807,N_1190);
or U3253 (N_3253,N_1641,N_65);
nand U3254 (N_3254,N_1455,N_1611);
nand U3255 (N_3255,N_779,N_2352);
nor U3256 (N_3256,N_1959,N_2087);
and U3257 (N_3257,N_634,N_2143);
or U3258 (N_3258,N_1263,N_1100);
or U3259 (N_3259,N_1645,N_2063);
nand U3260 (N_3260,N_2250,N_222);
or U3261 (N_3261,N_1955,N_1802);
nor U3262 (N_3262,N_811,N_530);
xnor U3263 (N_3263,N_862,N_233);
nand U3264 (N_3264,N_1993,N_143);
and U3265 (N_3265,N_989,N_1410);
nand U3266 (N_3266,N_201,N_676);
nand U3267 (N_3267,N_276,N_829);
nand U3268 (N_3268,N_638,N_2202);
or U3269 (N_3269,N_895,N_1395);
nand U3270 (N_3270,N_742,N_2471);
nor U3271 (N_3271,N_324,N_2125);
and U3272 (N_3272,N_1606,N_845);
nand U3273 (N_3273,N_2351,N_2419);
and U3274 (N_3274,N_1414,N_312);
nor U3275 (N_3275,N_2292,N_475);
nand U3276 (N_3276,N_1285,N_769);
nand U3277 (N_3277,N_938,N_823);
nor U3278 (N_3278,N_2195,N_1909);
and U3279 (N_3279,N_508,N_1353);
nor U3280 (N_3280,N_430,N_1341);
nand U3281 (N_3281,N_1869,N_727);
nor U3282 (N_3282,N_500,N_1371);
and U3283 (N_3283,N_1307,N_574);
or U3284 (N_3284,N_69,N_2469);
nor U3285 (N_3285,N_955,N_1423);
or U3286 (N_3286,N_2058,N_2002);
nor U3287 (N_3287,N_293,N_345);
nand U3288 (N_3288,N_812,N_1222);
nand U3289 (N_3289,N_1783,N_2446);
and U3290 (N_3290,N_524,N_1317);
nand U3291 (N_3291,N_914,N_1174);
nand U3292 (N_3292,N_179,N_1229);
or U3293 (N_3293,N_1891,N_1961);
or U3294 (N_3294,N_1824,N_991);
nor U3295 (N_3295,N_1590,N_63);
and U3296 (N_3296,N_1821,N_1221);
nand U3297 (N_3297,N_7,N_1844);
nand U3298 (N_3298,N_1575,N_1542);
and U3299 (N_3299,N_489,N_1609);
or U3300 (N_3300,N_884,N_1405);
and U3301 (N_3301,N_548,N_421);
and U3302 (N_3302,N_1422,N_2485);
nor U3303 (N_3303,N_1675,N_1944);
and U3304 (N_3304,N_463,N_381);
or U3305 (N_3305,N_804,N_1594);
and U3306 (N_3306,N_1120,N_1620);
and U3307 (N_3307,N_620,N_1440);
xnor U3308 (N_3308,N_1576,N_1716);
nor U3309 (N_3309,N_560,N_1608);
nor U3310 (N_3310,N_464,N_2076);
or U3311 (N_3311,N_1056,N_927);
nand U3312 (N_3312,N_2226,N_1971);
and U3313 (N_3313,N_1094,N_2458);
nor U3314 (N_3314,N_1169,N_2318);
or U3315 (N_3315,N_2285,N_1634);
or U3316 (N_3316,N_2046,N_2340);
or U3317 (N_3317,N_717,N_409);
nand U3318 (N_3318,N_2233,N_1618);
and U3319 (N_3319,N_957,N_35);
nand U3320 (N_3320,N_131,N_655);
or U3321 (N_3321,N_2028,N_174);
xor U3322 (N_3322,N_1185,N_687);
xnor U3323 (N_3323,N_2082,N_1234);
nor U3324 (N_3324,N_2370,N_1583);
nand U3325 (N_3325,N_1792,N_770);
nor U3326 (N_3326,N_479,N_579);
nor U3327 (N_3327,N_1117,N_321);
xor U3328 (N_3328,N_1145,N_648);
nand U3329 (N_3329,N_550,N_2173);
nor U3330 (N_3330,N_720,N_1055);
nor U3331 (N_3331,N_34,N_2151);
nor U3332 (N_3332,N_2137,N_1332);
nor U3333 (N_3333,N_155,N_1471);
and U3334 (N_3334,N_2249,N_1975);
or U3335 (N_3335,N_369,N_1151);
or U3336 (N_3336,N_2223,N_2124);
and U3337 (N_3337,N_1404,N_692);
nor U3338 (N_3338,N_2166,N_657);
nand U3339 (N_3339,N_1013,N_943);
nor U3340 (N_3340,N_567,N_1045);
or U3341 (N_3341,N_859,N_735);
and U3342 (N_3342,N_1235,N_1532);
or U3343 (N_3343,N_219,N_589);
and U3344 (N_3344,N_186,N_2247);
nand U3345 (N_3345,N_1065,N_1686);
or U3346 (N_3346,N_2207,N_981);
and U3347 (N_3347,N_1296,N_1162);
nand U3348 (N_3348,N_1679,N_854);
and U3349 (N_3349,N_2267,N_1383);
xor U3350 (N_3350,N_2089,N_613);
xnor U3351 (N_3351,N_1328,N_697);
nor U3352 (N_3352,N_1327,N_1061);
nor U3353 (N_3353,N_626,N_1954);
or U3354 (N_3354,N_2098,N_999);
nor U3355 (N_3355,N_892,N_1245);
and U3356 (N_3356,N_1214,N_1992);
xor U3357 (N_3357,N_2312,N_1016);
and U3358 (N_3358,N_2117,N_238);
nor U3359 (N_3359,N_1521,N_939);
or U3360 (N_3360,N_392,N_259);
and U3361 (N_3361,N_158,N_216);
nor U3362 (N_3362,N_667,N_1962);
nor U3363 (N_3363,N_633,N_344);
and U3364 (N_3364,N_937,N_1947);
and U3365 (N_3365,N_1666,N_1496);
and U3366 (N_3366,N_1430,N_432);
nand U3367 (N_3367,N_2467,N_2427);
or U3368 (N_3368,N_507,N_1106);
or U3369 (N_3369,N_474,N_2338);
or U3370 (N_3370,N_135,N_54);
nand U3371 (N_3371,N_2147,N_378);
xor U3372 (N_3372,N_1356,N_1130);
nor U3373 (N_3373,N_305,N_127);
nor U3374 (N_3374,N_2492,N_963);
nor U3375 (N_3375,N_960,N_1002);
nor U3376 (N_3376,N_1347,N_455);
nor U3377 (N_3377,N_738,N_2305);
nand U3378 (N_3378,N_913,N_1487);
nor U3379 (N_3379,N_2077,N_272);
nor U3380 (N_3380,N_2322,N_2070);
or U3381 (N_3381,N_1628,N_1708);
and U3382 (N_3382,N_1707,N_195);
or U3383 (N_3383,N_1700,N_1635);
and U3384 (N_3384,N_2240,N_2487);
nor U3385 (N_3385,N_33,N_119);
xnor U3386 (N_3386,N_1736,N_1030);
or U3387 (N_3387,N_1560,N_1472);
and U3388 (N_3388,N_1559,N_495);
and U3389 (N_3389,N_1256,N_1172);
and U3390 (N_3390,N_108,N_2027);
nand U3391 (N_3391,N_1006,N_2266);
xnor U3392 (N_3392,N_933,N_2327);
nand U3393 (N_3393,N_918,N_266);
nand U3394 (N_3394,N_450,N_1126);
or U3395 (N_3395,N_2490,N_1023);
xnor U3396 (N_3396,N_732,N_1053);
and U3397 (N_3397,N_1228,N_2380);
nand U3398 (N_3398,N_19,N_526);
and U3399 (N_3399,N_2182,N_1159);
or U3400 (N_3400,N_401,N_231);
or U3401 (N_3401,N_915,N_886);
nor U3402 (N_3402,N_983,N_425);
and U3403 (N_3403,N_570,N_17);
nor U3404 (N_3404,N_1168,N_932);
and U3405 (N_3405,N_861,N_282);
and U3406 (N_3406,N_2160,N_931);
and U3407 (N_3407,N_1951,N_2227);
and U3408 (N_3408,N_1309,N_880);
and U3409 (N_3409,N_497,N_903);
or U3410 (N_3410,N_2279,N_1165);
nand U3411 (N_3411,N_1249,N_990);
and U3412 (N_3412,N_346,N_1661);
nor U3413 (N_3413,N_1756,N_156);
nand U3414 (N_3414,N_1442,N_694);
nor U3415 (N_3415,N_1225,N_715);
xor U3416 (N_3416,N_1574,N_1393);
and U3417 (N_3417,N_2437,N_71);
and U3418 (N_3418,N_329,N_12);
nand U3419 (N_3419,N_1554,N_864);
and U3420 (N_3420,N_279,N_555);
and U3421 (N_3421,N_2310,N_1774);
nor U3422 (N_3422,N_2038,N_1154);
and U3423 (N_3423,N_2136,N_826);
nor U3424 (N_3424,N_2121,N_1840);
xor U3425 (N_3425,N_1385,N_2185);
nor U3426 (N_3426,N_1770,N_1134);
nand U3427 (N_3427,N_2330,N_138);
nand U3428 (N_3428,N_314,N_36);
xor U3429 (N_3429,N_582,N_2049);
or U3430 (N_3430,N_2013,N_1580);
and U3431 (N_3431,N_1148,N_1534);
nor U3432 (N_3432,N_1485,N_527);
and U3433 (N_3433,N_1269,N_1217);
nand U3434 (N_3434,N_671,N_1436);
nand U3435 (N_3435,N_370,N_1788);
or U3436 (N_3436,N_878,N_828);
nor U3437 (N_3437,N_98,N_814);
nor U3438 (N_3438,N_1704,N_852);
and U3439 (N_3439,N_698,N_1231);
nand U3440 (N_3440,N_707,N_2189);
nand U3441 (N_3441,N_1597,N_759);
nand U3442 (N_3442,N_897,N_196);
xor U3443 (N_3443,N_1528,N_964);
or U3444 (N_3444,N_477,N_2126);
nand U3445 (N_3445,N_536,N_2165);
nor U3446 (N_3446,N_2007,N_2130);
and U3447 (N_3447,N_1667,N_415);
nor U3448 (N_3448,N_1201,N_1031);
xor U3449 (N_3449,N_1880,N_974);
and U3450 (N_3450,N_1782,N_1418);
or U3451 (N_3451,N_438,N_452);
nor U3452 (N_3452,N_985,N_1531);
and U3453 (N_3453,N_656,N_1731);
and U3454 (N_3454,N_1048,N_1470);
nand U3455 (N_3455,N_1768,N_167);
and U3456 (N_3456,N_187,N_1827);
or U3457 (N_3457,N_2200,N_2260);
or U3458 (N_3458,N_2304,N_2270);
nor U3459 (N_3459,N_1607,N_2120);
or U3460 (N_3460,N_2039,N_494);
nor U3461 (N_3461,N_840,N_2154);
and U3462 (N_3462,N_290,N_597);
nor U3463 (N_3463,N_668,N_1479);
nand U3464 (N_3464,N_59,N_1952);
or U3465 (N_3465,N_894,N_2052);
or U3466 (N_3466,N_260,N_1246);
nor U3467 (N_3467,N_1481,N_2321);
nor U3468 (N_3468,N_171,N_1800);
or U3469 (N_3469,N_1524,N_1642);
nor U3470 (N_3470,N_1326,N_1742);
nor U3471 (N_3471,N_1453,N_1931);
and U3472 (N_3472,N_1942,N_1412);
nand U3473 (N_3473,N_1171,N_1836);
nor U3474 (N_3474,N_956,N_1968);
nor U3475 (N_3475,N_2011,N_1826);
or U3476 (N_3476,N_724,N_2061);
and U3477 (N_3477,N_177,N_289);
or U3478 (N_3478,N_1919,N_349);
nor U3479 (N_3479,N_1672,N_1619);
nor U3480 (N_3480,N_1167,N_1917);
nand U3481 (N_3481,N_2308,N_758);
xor U3482 (N_3482,N_1784,N_2134);
or U3483 (N_3483,N_2201,N_1762);
nand U3484 (N_3484,N_197,N_292);
nand U3485 (N_3485,N_1,N_646);
or U3486 (N_3486,N_2161,N_2048);
and U3487 (N_3487,N_899,N_2334);
or U3488 (N_3488,N_2356,N_1714);
and U3489 (N_3489,N_1315,N_1796);
nor U3490 (N_3490,N_1810,N_1411);
or U3491 (N_3491,N_1713,N_1206);
xor U3492 (N_3492,N_1937,N_1865);
nor U3493 (N_3493,N_3,N_538);
xor U3494 (N_3494,N_749,N_2041);
nor U3495 (N_3495,N_1927,N_1136);
and U3496 (N_3496,N_1108,N_1240);
or U3497 (N_3497,N_1457,N_882);
and U3498 (N_3498,N_1535,N_1985);
or U3499 (N_3499,N_2449,N_2235);
nor U3500 (N_3500,N_1851,N_1001);
and U3501 (N_3501,N_380,N_1143);
xnor U3502 (N_3502,N_2412,N_741);
nand U3503 (N_3503,N_1896,N_1207);
and U3504 (N_3504,N_576,N_640);
nand U3505 (N_3505,N_2069,N_1754);
nor U3506 (N_3506,N_1705,N_1538);
and U3507 (N_3507,N_1860,N_547);
nand U3508 (N_3508,N_2482,N_1908);
nand U3509 (N_3509,N_1673,N_986);
nor U3510 (N_3510,N_1932,N_1579);
and U3511 (N_3511,N_1864,N_306);
nor U3512 (N_3512,N_1308,N_288);
or U3513 (N_3513,N_1182,N_1238);
nand U3514 (N_3514,N_1303,N_2448);
nor U3515 (N_3515,N_2193,N_1636);
nand U3516 (N_3516,N_1354,N_2258);
and U3517 (N_3517,N_164,N_313);
and U3518 (N_3518,N_1019,N_1626);
nand U3519 (N_3519,N_571,N_1076);
and U3520 (N_3520,N_1726,N_1883);
or U3521 (N_3521,N_2068,N_1084);
xnor U3522 (N_3522,N_1643,N_1775);
or U3523 (N_3523,N_2263,N_1682);
xnor U3524 (N_3524,N_762,N_466);
nor U3525 (N_3525,N_2454,N_1546);
and U3526 (N_3526,N_525,N_552);
xor U3527 (N_3527,N_211,N_2324);
and U3528 (N_3528,N_1183,N_2217);
and U3529 (N_3529,N_1855,N_67);
and U3530 (N_3530,N_737,N_498);
nor U3531 (N_3531,N_1069,N_1063);
and U3532 (N_3532,N_753,N_1983);
nor U3533 (N_3533,N_703,N_511);
and U3534 (N_3534,N_1965,N_2333);
or U3535 (N_3535,N_343,N_1511);
or U3536 (N_3536,N_2289,N_1088);
or U3537 (N_3537,N_357,N_1243);
nor U3538 (N_3538,N_1568,N_2372);
nor U3539 (N_3539,N_39,N_142);
and U3540 (N_3540,N_249,N_1306);
nand U3541 (N_3541,N_1541,N_810);
and U3542 (N_3542,N_1125,N_299);
nor U3543 (N_3543,N_2478,N_268);
nor U3544 (N_3544,N_2462,N_793);
or U3545 (N_3545,N_383,N_190);
nor U3546 (N_3546,N_1432,N_443);
and U3547 (N_3547,N_2211,N_359);
nor U3548 (N_3548,N_596,N_1859);
or U3549 (N_3549,N_2108,N_181);
nand U3550 (N_3550,N_966,N_2162);
or U3551 (N_3551,N_670,N_602);
xor U3552 (N_3552,N_1202,N_1498);
and U3553 (N_3553,N_719,N_1463);
xnor U3554 (N_3554,N_189,N_1166);
and U3555 (N_3555,N_1047,N_1977);
nand U3556 (N_3556,N_1799,N_460);
nand U3557 (N_3557,N_1101,N_1425);
or U3558 (N_3558,N_665,N_382);
nor U3559 (N_3559,N_505,N_1842);
and U3560 (N_3560,N_2459,N_2188);
or U3561 (N_3561,N_150,N_404);
nor U3562 (N_3562,N_2149,N_1352);
nand U3563 (N_3563,N_362,N_128);
or U3564 (N_3564,N_911,N_1052);
xnor U3565 (N_3565,N_1389,N_240);
and U3566 (N_3566,N_348,N_1585);
xor U3567 (N_3567,N_2019,N_1282);
and U3568 (N_3568,N_1181,N_1939);
nor U3569 (N_3569,N_604,N_1740);
nand U3570 (N_3570,N_1014,N_831);
or U3571 (N_3571,N_2016,N_1180);
nand U3572 (N_3572,N_539,N_402);
nor U3573 (N_3573,N_2155,N_1690);
or U3574 (N_3574,N_844,N_1677);
nor U3575 (N_3575,N_1140,N_1870);
or U3576 (N_3576,N_1998,N_1070);
nor U3577 (N_3577,N_889,N_2274);
or U3578 (N_3578,N_2198,N_1995);
xnor U3579 (N_3579,N_1547,N_1837);
nand U3580 (N_3580,N_41,N_1340);
nand U3581 (N_3581,N_2034,N_1567);
and U3582 (N_3582,N_137,N_183);
or U3583 (N_3583,N_66,N_1251);
nor U3584 (N_3584,N_541,N_1570);
xor U3585 (N_3585,N_2275,N_435);
and U3586 (N_3586,N_1208,N_250);
or U3587 (N_3587,N_952,N_1593);
and U3588 (N_3588,N_973,N_1314);
and U3589 (N_3589,N_1862,N_1491);
nor U3590 (N_3590,N_2102,N_2006);
or U3591 (N_3591,N_705,N_1362);
or U3592 (N_3592,N_151,N_1444);
or U3593 (N_3593,N_1833,N_1210);
or U3594 (N_3594,N_191,N_2168);
nand U3595 (N_3595,N_1943,N_2000);
nand U3596 (N_3596,N_360,N_225);
or U3597 (N_3597,N_264,N_1260);
and U3598 (N_3598,N_1721,N_1617);
nor U3599 (N_3599,N_1501,N_2447);
or U3600 (N_3600,N_1957,N_405);
nor U3601 (N_3601,N_501,N_310);
nand U3602 (N_3602,N_1237,N_212);
or U3603 (N_3603,N_575,N_1111);
nand U3604 (N_3604,N_959,N_666);
nor U3605 (N_3605,N_2418,N_1761);
nand U3606 (N_3606,N_953,N_2129);
and U3607 (N_3607,N_1589,N_746);
nor U3608 (N_3608,N_2209,N_1219);
or U3609 (N_3609,N_78,N_2044);
xor U3610 (N_3610,N_1490,N_971);
nor U3611 (N_3611,N_1706,N_1771);
nor U3612 (N_3612,N_2131,N_2315);
nor U3613 (N_3613,N_659,N_1018);
or U3614 (N_3614,N_540,N_2488);
nand U3615 (N_3615,N_1223,N_585);
or U3616 (N_3616,N_2273,N_509);
xor U3617 (N_3617,N_1039,N_1135);
nand U3618 (N_3618,N_1099,N_1147);
nand U3619 (N_3619,N_860,N_154);
nand U3620 (N_3620,N_1497,N_2094);
and U3621 (N_3621,N_1778,N_72);
and U3622 (N_3622,N_1592,N_1656);
nand U3623 (N_3623,N_377,N_857);
nand U3624 (N_3624,N_1946,N_618);
and U3625 (N_3625,N_37,N_1304);
nor U3626 (N_3626,N_1755,N_2479);
nor U3627 (N_3627,N_1068,N_2431);
or U3628 (N_3628,N_1278,N_1963);
nor U3629 (N_3629,N_2359,N_2456);
nor U3630 (N_3630,N_744,N_350);
nand U3631 (N_3631,N_2014,N_664);
and U3632 (N_3632,N_1295,N_661);
or U3633 (N_3633,N_1086,N_808);
nor U3634 (N_3634,N_1902,N_2392);
and U3635 (N_3635,N_906,N_1967);
nor U3636 (N_3636,N_2276,N_2383);
nor U3637 (N_3637,N_2452,N_1924);
and U3638 (N_3638,N_923,N_393);
or U3639 (N_3639,N_182,N_1925);
or U3640 (N_3640,N_1273,N_1093);
nor U3641 (N_3641,N_2307,N_518);
xor U3642 (N_3642,N_529,N_114);
or U3643 (N_3643,N_300,N_1369);
or U3644 (N_3644,N_1715,N_339);
or U3645 (N_3645,N_1562,N_1564);
and U3646 (N_3646,N_2269,N_2397);
or U3647 (N_3647,N_630,N_1291);
nand U3648 (N_3648,N_1537,N_1650);
nand U3649 (N_3649,N_1199,N_1103);
nor U3650 (N_3650,N_373,N_116);
xnor U3651 (N_3651,N_874,N_1193);
nand U3652 (N_3652,N_1832,N_1809);
or U3653 (N_3653,N_1098,N_267);
and U3654 (N_3654,N_2432,N_824);
and U3655 (N_3655,N_997,N_1239);
nor U3656 (N_3656,N_403,N_2433);
or U3657 (N_3657,N_2254,N_967);
or U3658 (N_3658,N_1829,N_2218);
xnor U3659 (N_3659,N_1825,N_822);
and U3660 (N_3660,N_162,N_451);
or U3661 (N_3661,N_1032,N_731);
or U3662 (N_3662,N_1270,N_584);
nand U3663 (N_3663,N_1359,N_223);
or U3664 (N_3664,N_772,N_1232);
and U3665 (N_3665,N_2373,N_2080);
nor U3666 (N_3666,N_1175,N_723);
and U3667 (N_3667,N_89,N_1882);
xor U3668 (N_3668,N_2286,N_206);
or U3669 (N_3669,N_1596,N_10);
and U3670 (N_3670,N_1492,N_1717);
or U3671 (N_3671,N_1149,N_930);
nand U3672 (N_3672,N_2078,N_1437);
or U3673 (N_3673,N_1003,N_2457);
nor U3674 (N_3674,N_91,N_385);
nand U3675 (N_3675,N_2369,N_204);
and U3676 (N_3676,N_693,N_27);
and U3677 (N_3677,N_2073,N_677);
nor U3678 (N_3678,N_1156,N_49);
and U3679 (N_3679,N_2441,N_1122);
nor U3680 (N_3680,N_148,N_777);
or U3681 (N_3681,N_942,N_1275);
or U3682 (N_3682,N_767,N_1804);
or U3683 (N_3683,N_170,N_2238);
or U3684 (N_3684,N_237,N_1683);
xor U3685 (N_3685,N_1684,N_506);
nand U3686 (N_3686,N_1764,N_5);
and U3687 (N_3687,N_85,N_100);
nand U3688 (N_3688,N_924,N_685);
nor U3689 (N_3689,N_888,N_1543);
nor U3690 (N_3690,N_968,N_462);
or U3691 (N_3691,N_449,N_2390);
nand U3692 (N_3692,N_160,N_1449);
and U3693 (N_3693,N_1549,N_622);
and U3694 (N_3694,N_1843,N_680);
and U3695 (N_3695,N_1277,N_257);
or U3696 (N_3696,N_232,N_1691);
xor U3697 (N_3697,N_578,N_83);
nor U3698 (N_3698,N_298,N_1739);
and U3699 (N_3699,N_922,N_1200);
nor U3700 (N_3700,N_1197,N_1331);
or U3701 (N_3701,N_1224,N_1805);
xnor U3702 (N_3702,N_1460,N_773);
nand U3703 (N_3703,N_1212,N_2400);
nand U3704 (N_3704,N_1662,N_815);
and U3705 (N_3705,N_1218,N_1074);
or U3706 (N_3706,N_294,N_427);
and U3707 (N_3707,N_2466,N_572);
or U3708 (N_3708,N_1752,N_210);
nor U3709 (N_3709,N_152,N_1551);
nand U3710 (N_3710,N_1866,N_721);
or U3711 (N_3711,N_1071,N_123);
or U3712 (N_3712,N_64,N_457);
nor U3713 (N_3713,N_1671,N_90);
nand U3714 (N_3714,N_2367,N_2234);
or U3715 (N_3715,N_2368,N_70);
nand U3716 (N_3716,N_980,N_594);
nand U3717 (N_3717,N_2015,N_1813);
nand U3718 (N_3718,N_2152,N_1302);
nand U3719 (N_3719,N_689,N_1286);
nor U3720 (N_3720,N_333,N_1294);
nand U3721 (N_3721,N_1292,N_978);
nand U3722 (N_3722,N_641,N_1769);
or U3723 (N_3723,N_1435,N_921);
xnor U3724 (N_3724,N_1474,N_1000);
nor U3725 (N_3725,N_2464,N_398);
or U3726 (N_3726,N_2470,N_1079);
or U3727 (N_3727,N_215,N_1856);
nand U3728 (N_3728,N_1849,N_797);
and U3729 (N_3729,N_1443,N_1811);
nand U3730 (N_3730,N_165,N_1211);
or U3731 (N_3731,N_56,N_178);
and U3732 (N_3732,N_1281,N_1621);
xnor U3733 (N_3733,N_1163,N_1949);
or U3734 (N_3734,N_766,N_1914);
and U3735 (N_3735,N_1033,N_1338);
and U3736 (N_3736,N_1363,N_2237);
nand U3737 (N_3737,N_1041,N_1513);
nor U3738 (N_3738,N_2051,N_645);
or U3739 (N_3739,N_2133,N_367);
nand U3740 (N_3740,N_1530,N_2364);
xnor U3741 (N_3741,N_608,N_1254);
nand U3742 (N_3742,N_32,N_1480);
nor U3743 (N_3743,N_1817,N_557);
nand U3744 (N_3744,N_285,N_1305);
nor U3745 (N_3745,N_1397,N_1192);
nor U3746 (N_3746,N_2214,N_337);
and U3747 (N_3747,N_2311,N_1790);
and U3748 (N_3748,N_1124,N_284);
or U3749 (N_3749,N_2384,N_1839);
or U3750 (N_3750,N_2215,N_469);
nand U3751 (N_3751,N_30,N_212);
nand U3752 (N_3752,N_1275,N_946);
or U3753 (N_3753,N_1698,N_1315);
nand U3754 (N_3754,N_2075,N_173);
nand U3755 (N_3755,N_1972,N_32);
nand U3756 (N_3756,N_1258,N_1600);
nand U3757 (N_3757,N_1637,N_378);
and U3758 (N_3758,N_2447,N_1757);
and U3759 (N_3759,N_1447,N_2042);
nand U3760 (N_3760,N_794,N_1680);
and U3761 (N_3761,N_786,N_1007);
and U3762 (N_3762,N_695,N_657);
nand U3763 (N_3763,N_1069,N_755);
or U3764 (N_3764,N_464,N_899);
or U3765 (N_3765,N_2446,N_1076);
or U3766 (N_3766,N_598,N_2219);
nand U3767 (N_3767,N_2255,N_2171);
and U3768 (N_3768,N_91,N_534);
nor U3769 (N_3769,N_2247,N_1353);
nand U3770 (N_3770,N_392,N_247);
nand U3771 (N_3771,N_978,N_2200);
nor U3772 (N_3772,N_121,N_516);
and U3773 (N_3773,N_1522,N_743);
or U3774 (N_3774,N_507,N_273);
xor U3775 (N_3775,N_725,N_2098);
xor U3776 (N_3776,N_514,N_1285);
nand U3777 (N_3777,N_348,N_1145);
or U3778 (N_3778,N_1513,N_998);
and U3779 (N_3779,N_403,N_295);
and U3780 (N_3780,N_2261,N_1650);
or U3781 (N_3781,N_710,N_404);
nor U3782 (N_3782,N_99,N_973);
nand U3783 (N_3783,N_255,N_1330);
and U3784 (N_3784,N_333,N_827);
nor U3785 (N_3785,N_927,N_627);
and U3786 (N_3786,N_1675,N_143);
nor U3787 (N_3787,N_2476,N_891);
nor U3788 (N_3788,N_733,N_790);
nand U3789 (N_3789,N_958,N_388);
nand U3790 (N_3790,N_365,N_1373);
nor U3791 (N_3791,N_503,N_1583);
and U3792 (N_3792,N_547,N_1155);
and U3793 (N_3793,N_2386,N_1784);
nor U3794 (N_3794,N_1754,N_2323);
xnor U3795 (N_3795,N_1403,N_830);
and U3796 (N_3796,N_2057,N_371);
xor U3797 (N_3797,N_1128,N_250);
nor U3798 (N_3798,N_1605,N_1880);
nor U3799 (N_3799,N_364,N_1317);
or U3800 (N_3800,N_1006,N_637);
nand U3801 (N_3801,N_2413,N_1730);
nand U3802 (N_3802,N_2433,N_888);
nand U3803 (N_3803,N_842,N_1366);
or U3804 (N_3804,N_2483,N_1643);
nand U3805 (N_3805,N_511,N_1214);
and U3806 (N_3806,N_1629,N_908);
nor U3807 (N_3807,N_1733,N_2375);
nand U3808 (N_3808,N_195,N_1091);
nor U3809 (N_3809,N_268,N_1832);
nand U3810 (N_3810,N_1706,N_1364);
nor U3811 (N_3811,N_804,N_641);
nor U3812 (N_3812,N_1451,N_1881);
and U3813 (N_3813,N_772,N_708);
nand U3814 (N_3814,N_1068,N_2249);
nor U3815 (N_3815,N_1589,N_1584);
and U3816 (N_3816,N_1831,N_1489);
nor U3817 (N_3817,N_2400,N_1940);
or U3818 (N_3818,N_2259,N_449);
nor U3819 (N_3819,N_1735,N_1291);
or U3820 (N_3820,N_2265,N_310);
or U3821 (N_3821,N_2325,N_584);
and U3822 (N_3822,N_1594,N_5);
and U3823 (N_3823,N_2267,N_898);
or U3824 (N_3824,N_53,N_1060);
and U3825 (N_3825,N_2408,N_1941);
and U3826 (N_3826,N_1924,N_424);
or U3827 (N_3827,N_1844,N_683);
nand U3828 (N_3828,N_2042,N_2429);
or U3829 (N_3829,N_2407,N_1201);
xor U3830 (N_3830,N_1207,N_2289);
nand U3831 (N_3831,N_59,N_2327);
xor U3832 (N_3832,N_1797,N_362);
and U3833 (N_3833,N_1234,N_893);
nand U3834 (N_3834,N_206,N_1915);
and U3835 (N_3835,N_2128,N_27);
or U3836 (N_3836,N_1360,N_393);
nor U3837 (N_3837,N_868,N_1560);
nor U3838 (N_3838,N_782,N_1600);
nand U3839 (N_3839,N_28,N_365);
nand U3840 (N_3840,N_1317,N_629);
or U3841 (N_3841,N_2467,N_544);
or U3842 (N_3842,N_6,N_2307);
nor U3843 (N_3843,N_487,N_2283);
nor U3844 (N_3844,N_1384,N_1402);
nand U3845 (N_3845,N_351,N_2372);
nand U3846 (N_3846,N_2285,N_520);
and U3847 (N_3847,N_1718,N_1926);
nand U3848 (N_3848,N_633,N_335);
and U3849 (N_3849,N_360,N_108);
or U3850 (N_3850,N_151,N_1740);
or U3851 (N_3851,N_1429,N_501);
and U3852 (N_3852,N_2240,N_1975);
or U3853 (N_3853,N_2179,N_160);
nand U3854 (N_3854,N_1974,N_163);
and U3855 (N_3855,N_1472,N_337);
nand U3856 (N_3856,N_1389,N_243);
nand U3857 (N_3857,N_1016,N_1126);
and U3858 (N_3858,N_724,N_1937);
nand U3859 (N_3859,N_648,N_1992);
nor U3860 (N_3860,N_1399,N_950);
or U3861 (N_3861,N_1510,N_1912);
nand U3862 (N_3862,N_1769,N_905);
or U3863 (N_3863,N_108,N_1042);
nand U3864 (N_3864,N_1270,N_554);
nor U3865 (N_3865,N_730,N_418);
or U3866 (N_3866,N_102,N_547);
and U3867 (N_3867,N_1678,N_1137);
or U3868 (N_3868,N_1949,N_1783);
and U3869 (N_3869,N_563,N_1655);
and U3870 (N_3870,N_1967,N_1781);
nor U3871 (N_3871,N_1375,N_1177);
xnor U3872 (N_3872,N_628,N_765);
or U3873 (N_3873,N_553,N_56);
nand U3874 (N_3874,N_1886,N_898);
nor U3875 (N_3875,N_2069,N_1479);
nor U3876 (N_3876,N_1872,N_1740);
nor U3877 (N_3877,N_1010,N_1847);
nand U3878 (N_3878,N_85,N_416);
and U3879 (N_3879,N_360,N_631);
xnor U3880 (N_3880,N_16,N_1209);
nand U3881 (N_3881,N_562,N_261);
or U3882 (N_3882,N_1897,N_554);
or U3883 (N_3883,N_1788,N_1357);
nor U3884 (N_3884,N_377,N_459);
or U3885 (N_3885,N_1291,N_525);
nor U3886 (N_3886,N_2303,N_1862);
nand U3887 (N_3887,N_1018,N_974);
nand U3888 (N_3888,N_1153,N_1759);
nand U3889 (N_3889,N_1561,N_2148);
or U3890 (N_3890,N_28,N_1386);
and U3891 (N_3891,N_781,N_1128);
xor U3892 (N_3892,N_1671,N_1790);
and U3893 (N_3893,N_219,N_534);
xor U3894 (N_3894,N_46,N_837);
nand U3895 (N_3895,N_1661,N_2104);
and U3896 (N_3896,N_397,N_835);
nand U3897 (N_3897,N_2028,N_682);
or U3898 (N_3898,N_1306,N_642);
nand U3899 (N_3899,N_107,N_2342);
xnor U3900 (N_3900,N_1879,N_726);
xor U3901 (N_3901,N_175,N_1787);
nand U3902 (N_3902,N_2188,N_563);
nand U3903 (N_3903,N_1798,N_323);
or U3904 (N_3904,N_2025,N_2404);
and U3905 (N_3905,N_1377,N_1256);
nand U3906 (N_3906,N_2370,N_1568);
or U3907 (N_3907,N_468,N_1721);
nor U3908 (N_3908,N_2135,N_1695);
and U3909 (N_3909,N_854,N_1128);
or U3910 (N_3910,N_1500,N_2166);
or U3911 (N_3911,N_1739,N_1006);
nand U3912 (N_3912,N_2394,N_1618);
and U3913 (N_3913,N_2220,N_1370);
nand U3914 (N_3914,N_496,N_1122);
or U3915 (N_3915,N_2004,N_323);
and U3916 (N_3916,N_2437,N_1600);
xnor U3917 (N_3917,N_57,N_2017);
nor U3918 (N_3918,N_1582,N_475);
nand U3919 (N_3919,N_2330,N_1380);
or U3920 (N_3920,N_2022,N_1447);
or U3921 (N_3921,N_1791,N_413);
nor U3922 (N_3922,N_836,N_672);
or U3923 (N_3923,N_532,N_956);
xor U3924 (N_3924,N_1809,N_14);
and U3925 (N_3925,N_1860,N_1703);
nor U3926 (N_3926,N_1429,N_377);
or U3927 (N_3927,N_1368,N_2022);
nand U3928 (N_3928,N_1187,N_1347);
xnor U3929 (N_3929,N_1832,N_1034);
or U3930 (N_3930,N_1527,N_1314);
and U3931 (N_3931,N_1491,N_1729);
and U3932 (N_3932,N_1105,N_278);
and U3933 (N_3933,N_2251,N_945);
and U3934 (N_3934,N_1486,N_2120);
or U3935 (N_3935,N_286,N_1570);
and U3936 (N_3936,N_212,N_1608);
or U3937 (N_3937,N_2277,N_1116);
xnor U3938 (N_3938,N_2012,N_2144);
or U3939 (N_3939,N_2149,N_1664);
and U3940 (N_3940,N_854,N_2238);
and U3941 (N_3941,N_1980,N_554);
and U3942 (N_3942,N_670,N_85);
nor U3943 (N_3943,N_25,N_548);
or U3944 (N_3944,N_1631,N_650);
and U3945 (N_3945,N_1420,N_1460);
nand U3946 (N_3946,N_850,N_521);
and U3947 (N_3947,N_1648,N_1082);
xor U3948 (N_3948,N_1937,N_400);
nand U3949 (N_3949,N_1265,N_1598);
nand U3950 (N_3950,N_190,N_2214);
and U3951 (N_3951,N_2296,N_945);
or U3952 (N_3952,N_620,N_972);
nor U3953 (N_3953,N_1918,N_2327);
xnor U3954 (N_3954,N_568,N_1567);
and U3955 (N_3955,N_2328,N_2027);
nand U3956 (N_3956,N_511,N_171);
nor U3957 (N_3957,N_618,N_1534);
and U3958 (N_3958,N_1817,N_1240);
xor U3959 (N_3959,N_2361,N_825);
nor U3960 (N_3960,N_2070,N_2304);
or U3961 (N_3961,N_1217,N_733);
nor U3962 (N_3962,N_2460,N_2463);
nor U3963 (N_3963,N_469,N_68);
nor U3964 (N_3964,N_2380,N_1446);
nor U3965 (N_3965,N_419,N_1079);
nand U3966 (N_3966,N_67,N_2388);
nand U3967 (N_3967,N_1226,N_2127);
nand U3968 (N_3968,N_2111,N_1914);
or U3969 (N_3969,N_162,N_1797);
or U3970 (N_3970,N_1550,N_2424);
nand U3971 (N_3971,N_468,N_591);
nor U3972 (N_3972,N_1709,N_1588);
nand U3973 (N_3973,N_1491,N_798);
nor U3974 (N_3974,N_68,N_1091);
or U3975 (N_3975,N_1180,N_2103);
and U3976 (N_3976,N_1945,N_2109);
or U3977 (N_3977,N_1245,N_1720);
and U3978 (N_3978,N_913,N_924);
nand U3979 (N_3979,N_540,N_1836);
and U3980 (N_3980,N_1552,N_2270);
nor U3981 (N_3981,N_985,N_2175);
nor U3982 (N_3982,N_635,N_1943);
nor U3983 (N_3983,N_1524,N_2444);
or U3984 (N_3984,N_1102,N_659);
xor U3985 (N_3985,N_841,N_1326);
nand U3986 (N_3986,N_1751,N_1126);
nor U3987 (N_3987,N_2302,N_256);
nand U3988 (N_3988,N_468,N_2181);
nor U3989 (N_3989,N_1071,N_966);
or U3990 (N_3990,N_295,N_2477);
nand U3991 (N_3991,N_2321,N_1197);
nand U3992 (N_3992,N_1858,N_1353);
and U3993 (N_3993,N_1805,N_1369);
nand U3994 (N_3994,N_748,N_662);
nor U3995 (N_3995,N_1755,N_43);
and U3996 (N_3996,N_1685,N_185);
nand U3997 (N_3997,N_2253,N_2457);
nor U3998 (N_3998,N_518,N_929);
nand U3999 (N_3999,N_2396,N_2224);
xnor U4000 (N_4000,N_1978,N_1762);
and U4001 (N_4001,N_1339,N_1043);
nand U4002 (N_4002,N_1000,N_663);
and U4003 (N_4003,N_1387,N_1086);
xor U4004 (N_4004,N_2483,N_441);
and U4005 (N_4005,N_2379,N_1697);
and U4006 (N_4006,N_1964,N_1450);
or U4007 (N_4007,N_746,N_2479);
and U4008 (N_4008,N_190,N_941);
nor U4009 (N_4009,N_1395,N_426);
and U4010 (N_4010,N_1662,N_761);
or U4011 (N_4011,N_1082,N_728);
and U4012 (N_4012,N_1695,N_2204);
and U4013 (N_4013,N_178,N_1694);
or U4014 (N_4014,N_1343,N_1099);
nand U4015 (N_4015,N_916,N_1865);
or U4016 (N_4016,N_2189,N_2104);
nand U4017 (N_4017,N_1125,N_2101);
and U4018 (N_4018,N_343,N_2291);
or U4019 (N_4019,N_817,N_1633);
nand U4020 (N_4020,N_946,N_925);
and U4021 (N_4021,N_2306,N_1014);
and U4022 (N_4022,N_1812,N_70);
and U4023 (N_4023,N_719,N_1680);
nor U4024 (N_4024,N_2079,N_2413);
nand U4025 (N_4025,N_779,N_155);
and U4026 (N_4026,N_654,N_1556);
or U4027 (N_4027,N_2407,N_1616);
xor U4028 (N_4028,N_869,N_432);
xnor U4029 (N_4029,N_641,N_809);
nor U4030 (N_4030,N_1743,N_1055);
and U4031 (N_4031,N_292,N_1606);
nand U4032 (N_4032,N_578,N_1673);
and U4033 (N_4033,N_467,N_1278);
xnor U4034 (N_4034,N_1798,N_253);
or U4035 (N_4035,N_1991,N_2466);
xor U4036 (N_4036,N_2376,N_1669);
and U4037 (N_4037,N_1533,N_1275);
and U4038 (N_4038,N_1280,N_1276);
or U4039 (N_4039,N_351,N_147);
xnor U4040 (N_4040,N_1051,N_546);
nand U4041 (N_4041,N_420,N_235);
and U4042 (N_4042,N_2368,N_198);
nor U4043 (N_4043,N_740,N_612);
and U4044 (N_4044,N_336,N_547);
and U4045 (N_4045,N_1615,N_676);
and U4046 (N_4046,N_1550,N_1705);
xor U4047 (N_4047,N_215,N_771);
nor U4048 (N_4048,N_1289,N_1338);
nor U4049 (N_4049,N_647,N_481);
and U4050 (N_4050,N_305,N_1118);
nand U4051 (N_4051,N_250,N_2060);
and U4052 (N_4052,N_1680,N_2242);
nor U4053 (N_4053,N_1484,N_1552);
nor U4054 (N_4054,N_2153,N_1117);
xor U4055 (N_4055,N_1948,N_1477);
or U4056 (N_4056,N_275,N_2129);
and U4057 (N_4057,N_1583,N_338);
nand U4058 (N_4058,N_32,N_1681);
nand U4059 (N_4059,N_2439,N_2412);
or U4060 (N_4060,N_2334,N_1447);
or U4061 (N_4061,N_126,N_1251);
and U4062 (N_4062,N_1123,N_802);
xnor U4063 (N_4063,N_1662,N_585);
nand U4064 (N_4064,N_830,N_1567);
nand U4065 (N_4065,N_2306,N_727);
and U4066 (N_4066,N_970,N_1261);
or U4067 (N_4067,N_2438,N_1842);
and U4068 (N_4068,N_1126,N_1389);
nand U4069 (N_4069,N_2361,N_477);
nand U4070 (N_4070,N_2407,N_712);
or U4071 (N_4071,N_380,N_495);
nand U4072 (N_4072,N_967,N_1709);
xnor U4073 (N_4073,N_380,N_950);
and U4074 (N_4074,N_433,N_210);
or U4075 (N_4075,N_808,N_871);
xnor U4076 (N_4076,N_602,N_366);
and U4077 (N_4077,N_1600,N_2062);
nand U4078 (N_4078,N_2245,N_2179);
or U4079 (N_4079,N_527,N_1121);
nand U4080 (N_4080,N_2013,N_1518);
nor U4081 (N_4081,N_1197,N_1204);
or U4082 (N_4082,N_383,N_1773);
or U4083 (N_4083,N_477,N_851);
xnor U4084 (N_4084,N_763,N_756);
nor U4085 (N_4085,N_593,N_1143);
and U4086 (N_4086,N_385,N_257);
and U4087 (N_4087,N_1882,N_1931);
nor U4088 (N_4088,N_2048,N_899);
and U4089 (N_4089,N_2111,N_512);
or U4090 (N_4090,N_161,N_2441);
nor U4091 (N_4091,N_1382,N_2358);
and U4092 (N_4092,N_321,N_1271);
nor U4093 (N_4093,N_1148,N_1855);
nand U4094 (N_4094,N_2135,N_636);
and U4095 (N_4095,N_989,N_1343);
or U4096 (N_4096,N_1570,N_1767);
and U4097 (N_4097,N_2466,N_2143);
nand U4098 (N_4098,N_1792,N_1858);
and U4099 (N_4099,N_11,N_1819);
xor U4100 (N_4100,N_402,N_1030);
or U4101 (N_4101,N_236,N_1329);
or U4102 (N_4102,N_2048,N_546);
nand U4103 (N_4103,N_2222,N_2162);
nand U4104 (N_4104,N_1460,N_2079);
xnor U4105 (N_4105,N_2295,N_2060);
or U4106 (N_4106,N_620,N_1112);
or U4107 (N_4107,N_708,N_1805);
nand U4108 (N_4108,N_1048,N_142);
or U4109 (N_4109,N_1680,N_835);
and U4110 (N_4110,N_844,N_1769);
or U4111 (N_4111,N_1490,N_2431);
and U4112 (N_4112,N_1057,N_1046);
nor U4113 (N_4113,N_1301,N_184);
nand U4114 (N_4114,N_929,N_2245);
and U4115 (N_4115,N_1913,N_454);
and U4116 (N_4116,N_55,N_1470);
and U4117 (N_4117,N_1966,N_839);
xor U4118 (N_4118,N_887,N_2178);
nand U4119 (N_4119,N_2418,N_774);
and U4120 (N_4120,N_1565,N_2369);
and U4121 (N_4121,N_716,N_2219);
xor U4122 (N_4122,N_1023,N_422);
and U4123 (N_4123,N_2365,N_660);
and U4124 (N_4124,N_41,N_616);
nor U4125 (N_4125,N_853,N_1343);
xor U4126 (N_4126,N_139,N_295);
nand U4127 (N_4127,N_1326,N_1392);
or U4128 (N_4128,N_1213,N_2275);
nand U4129 (N_4129,N_494,N_1008);
and U4130 (N_4130,N_1224,N_1110);
or U4131 (N_4131,N_2056,N_369);
nor U4132 (N_4132,N_31,N_1217);
nor U4133 (N_4133,N_2465,N_938);
and U4134 (N_4134,N_690,N_822);
nand U4135 (N_4135,N_77,N_177);
nand U4136 (N_4136,N_2241,N_293);
nor U4137 (N_4137,N_1166,N_126);
nand U4138 (N_4138,N_2279,N_816);
nand U4139 (N_4139,N_377,N_2476);
nand U4140 (N_4140,N_1201,N_1898);
and U4141 (N_4141,N_1536,N_588);
and U4142 (N_4142,N_1531,N_1774);
nor U4143 (N_4143,N_1885,N_1370);
or U4144 (N_4144,N_1287,N_1734);
nand U4145 (N_4145,N_1909,N_84);
nor U4146 (N_4146,N_201,N_2048);
nand U4147 (N_4147,N_1755,N_976);
nand U4148 (N_4148,N_172,N_323);
or U4149 (N_4149,N_25,N_1090);
nor U4150 (N_4150,N_146,N_1921);
nand U4151 (N_4151,N_1009,N_1654);
or U4152 (N_4152,N_708,N_2311);
nand U4153 (N_4153,N_754,N_178);
or U4154 (N_4154,N_2385,N_1167);
nand U4155 (N_4155,N_550,N_144);
nand U4156 (N_4156,N_1096,N_1260);
or U4157 (N_4157,N_1409,N_1564);
nor U4158 (N_4158,N_1903,N_1591);
and U4159 (N_4159,N_1274,N_2114);
nor U4160 (N_4160,N_696,N_1093);
or U4161 (N_4161,N_614,N_1207);
or U4162 (N_4162,N_1162,N_941);
or U4163 (N_4163,N_168,N_549);
nor U4164 (N_4164,N_706,N_1484);
xnor U4165 (N_4165,N_523,N_1995);
or U4166 (N_4166,N_1601,N_1520);
and U4167 (N_4167,N_2146,N_515);
or U4168 (N_4168,N_785,N_274);
and U4169 (N_4169,N_1561,N_1517);
nor U4170 (N_4170,N_252,N_722);
nand U4171 (N_4171,N_890,N_1042);
xor U4172 (N_4172,N_372,N_4);
nor U4173 (N_4173,N_886,N_182);
and U4174 (N_4174,N_1350,N_777);
or U4175 (N_4175,N_1581,N_1637);
nor U4176 (N_4176,N_1703,N_1730);
xor U4177 (N_4177,N_1353,N_2123);
nor U4178 (N_4178,N_711,N_363);
nor U4179 (N_4179,N_2198,N_796);
and U4180 (N_4180,N_1188,N_2317);
or U4181 (N_4181,N_2007,N_215);
and U4182 (N_4182,N_941,N_1215);
or U4183 (N_4183,N_2372,N_281);
nand U4184 (N_4184,N_223,N_385);
nand U4185 (N_4185,N_1387,N_170);
and U4186 (N_4186,N_2175,N_2449);
and U4187 (N_4187,N_1360,N_2392);
or U4188 (N_4188,N_528,N_663);
or U4189 (N_4189,N_2359,N_1543);
nor U4190 (N_4190,N_998,N_901);
nand U4191 (N_4191,N_370,N_2117);
nand U4192 (N_4192,N_1209,N_667);
and U4193 (N_4193,N_1153,N_1173);
or U4194 (N_4194,N_1825,N_1397);
and U4195 (N_4195,N_1849,N_1104);
nor U4196 (N_4196,N_1967,N_1211);
or U4197 (N_4197,N_659,N_21);
nor U4198 (N_4198,N_1252,N_2164);
nor U4199 (N_4199,N_1685,N_565);
nor U4200 (N_4200,N_1061,N_199);
nor U4201 (N_4201,N_1610,N_1802);
nor U4202 (N_4202,N_1127,N_526);
nand U4203 (N_4203,N_299,N_2212);
and U4204 (N_4204,N_337,N_2058);
and U4205 (N_4205,N_1259,N_651);
and U4206 (N_4206,N_518,N_1159);
nand U4207 (N_4207,N_1279,N_1617);
or U4208 (N_4208,N_1274,N_1757);
and U4209 (N_4209,N_2171,N_1316);
and U4210 (N_4210,N_23,N_1639);
or U4211 (N_4211,N_902,N_1180);
nor U4212 (N_4212,N_1353,N_2113);
and U4213 (N_4213,N_591,N_1195);
xor U4214 (N_4214,N_1755,N_200);
nor U4215 (N_4215,N_594,N_79);
nand U4216 (N_4216,N_707,N_338);
nor U4217 (N_4217,N_279,N_2330);
or U4218 (N_4218,N_843,N_47);
nand U4219 (N_4219,N_2185,N_31);
nand U4220 (N_4220,N_623,N_807);
and U4221 (N_4221,N_136,N_1223);
xnor U4222 (N_4222,N_2009,N_346);
nor U4223 (N_4223,N_891,N_2180);
or U4224 (N_4224,N_1859,N_102);
nor U4225 (N_4225,N_226,N_1102);
nor U4226 (N_4226,N_1439,N_1383);
and U4227 (N_4227,N_1105,N_1688);
nand U4228 (N_4228,N_2296,N_2174);
nor U4229 (N_4229,N_2147,N_1499);
and U4230 (N_4230,N_1367,N_2123);
or U4231 (N_4231,N_194,N_394);
nor U4232 (N_4232,N_408,N_1314);
or U4233 (N_4233,N_1917,N_2032);
and U4234 (N_4234,N_1470,N_1660);
and U4235 (N_4235,N_1018,N_458);
xor U4236 (N_4236,N_931,N_1572);
nand U4237 (N_4237,N_1965,N_344);
xor U4238 (N_4238,N_1236,N_2361);
nor U4239 (N_4239,N_1361,N_706);
or U4240 (N_4240,N_19,N_580);
nor U4241 (N_4241,N_788,N_793);
or U4242 (N_4242,N_1644,N_332);
or U4243 (N_4243,N_1034,N_1379);
or U4244 (N_4244,N_1914,N_2200);
nor U4245 (N_4245,N_1557,N_411);
nor U4246 (N_4246,N_1216,N_405);
xnor U4247 (N_4247,N_2032,N_439);
nand U4248 (N_4248,N_1849,N_182);
and U4249 (N_4249,N_2069,N_855);
and U4250 (N_4250,N_1265,N_2308);
and U4251 (N_4251,N_1406,N_741);
nor U4252 (N_4252,N_1302,N_545);
or U4253 (N_4253,N_1645,N_1159);
or U4254 (N_4254,N_1139,N_784);
nor U4255 (N_4255,N_29,N_1995);
nand U4256 (N_4256,N_900,N_367);
xor U4257 (N_4257,N_905,N_1289);
or U4258 (N_4258,N_1370,N_26);
xnor U4259 (N_4259,N_1350,N_2458);
and U4260 (N_4260,N_449,N_175);
or U4261 (N_4261,N_1814,N_776);
and U4262 (N_4262,N_269,N_956);
and U4263 (N_4263,N_276,N_709);
xor U4264 (N_4264,N_736,N_1073);
xnor U4265 (N_4265,N_493,N_578);
or U4266 (N_4266,N_2474,N_850);
xnor U4267 (N_4267,N_2355,N_1348);
or U4268 (N_4268,N_1831,N_2328);
nand U4269 (N_4269,N_1486,N_1223);
nor U4270 (N_4270,N_2093,N_2436);
nand U4271 (N_4271,N_1544,N_2394);
and U4272 (N_4272,N_2320,N_181);
and U4273 (N_4273,N_23,N_134);
nor U4274 (N_4274,N_2445,N_1610);
nor U4275 (N_4275,N_422,N_2061);
nand U4276 (N_4276,N_182,N_1639);
or U4277 (N_4277,N_827,N_1667);
xnor U4278 (N_4278,N_410,N_2291);
xor U4279 (N_4279,N_469,N_618);
xnor U4280 (N_4280,N_2379,N_800);
or U4281 (N_4281,N_220,N_1826);
and U4282 (N_4282,N_7,N_639);
and U4283 (N_4283,N_2068,N_568);
xor U4284 (N_4284,N_328,N_617);
xor U4285 (N_4285,N_1254,N_643);
and U4286 (N_4286,N_380,N_1713);
xnor U4287 (N_4287,N_1575,N_897);
and U4288 (N_4288,N_234,N_424);
and U4289 (N_4289,N_1948,N_606);
nand U4290 (N_4290,N_2322,N_255);
xor U4291 (N_4291,N_1550,N_808);
nand U4292 (N_4292,N_1953,N_1037);
or U4293 (N_4293,N_1529,N_1611);
nand U4294 (N_4294,N_628,N_1117);
nand U4295 (N_4295,N_2235,N_227);
nor U4296 (N_4296,N_872,N_2028);
and U4297 (N_4297,N_1948,N_519);
nor U4298 (N_4298,N_712,N_2006);
xnor U4299 (N_4299,N_26,N_2208);
or U4300 (N_4300,N_92,N_2077);
nor U4301 (N_4301,N_1821,N_202);
nand U4302 (N_4302,N_1169,N_2358);
or U4303 (N_4303,N_2343,N_978);
and U4304 (N_4304,N_139,N_1859);
and U4305 (N_4305,N_1256,N_591);
nand U4306 (N_4306,N_2053,N_1775);
nor U4307 (N_4307,N_368,N_1716);
or U4308 (N_4308,N_2155,N_327);
nand U4309 (N_4309,N_448,N_1436);
nand U4310 (N_4310,N_24,N_942);
xor U4311 (N_4311,N_1627,N_2196);
xnor U4312 (N_4312,N_918,N_1223);
xnor U4313 (N_4313,N_548,N_1883);
xor U4314 (N_4314,N_1799,N_2248);
and U4315 (N_4315,N_1384,N_1868);
nand U4316 (N_4316,N_1001,N_1474);
or U4317 (N_4317,N_2308,N_2029);
nand U4318 (N_4318,N_910,N_2151);
or U4319 (N_4319,N_389,N_417);
and U4320 (N_4320,N_228,N_348);
xor U4321 (N_4321,N_20,N_197);
nand U4322 (N_4322,N_475,N_769);
or U4323 (N_4323,N_28,N_123);
or U4324 (N_4324,N_2305,N_638);
nor U4325 (N_4325,N_2052,N_1043);
nor U4326 (N_4326,N_1245,N_2451);
nor U4327 (N_4327,N_785,N_1657);
and U4328 (N_4328,N_1923,N_1466);
and U4329 (N_4329,N_2148,N_759);
nand U4330 (N_4330,N_2058,N_1413);
nand U4331 (N_4331,N_450,N_1851);
nor U4332 (N_4332,N_657,N_2358);
and U4333 (N_4333,N_1023,N_648);
nor U4334 (N_4334,N_244,N_462);
xnor U4335 (N_4335,N_2091,N_1580);
nand U4336 (N_4336,N_1742,N_1965);
nor U4337 (N_4337,N_1255,N_932);
xnor U4338 (N_4338,N_237,N_443);
or U4339 (N_4339,N_1131,N_268);
nand U4340 (N_4340,N_2108,N_1550);
or U4341 (N_4341,N_808,N_2314);
xnor U4342 (N_4342,N_2220,N_899);
nor U4343 (N_4343,N_311,N_928);
nand U4344 (N_4344,N_1513,N_615);
nand U4345 (N_4345,N_1598,N_2097);
nor U4346 (N_4346,N_427,N_2110);
xor U4347 (N_4347,N_2454,N_1126);
and U4348 (N_4348,N_860,N_2389);
and U4349 (N_4349,N_34,N_1973);
or U4350 (N_4350,N_1323,N_1271);
or U4351 (N_4351,N_98,N_1986);
or U4352 (N_4352,N_1080,N_1822);
xor U4353 (N_4353,N_993,N_1090);
and U4354 (N_4354,N_1476,N_2388);
or U4355 (N_4355,N_1198,N_1599);
nand U4356 (N_4356,N_79,N_901);
nand U4357 (N_4357,N_1939,N_1213);
or U4358 (N_4358,N_92,N_674);
nand U4359 (N_4359,N_226,N_1885);
xnor U4360 (N_4360,N_2311,N_2222);
xor U4361 (N_4361,N_1251,N_1440);
nand U4362 (N_4362,N_408,N_923);
nand U4363 (N_4363,N_1363,N_74);
nor U4364 (N_4364,N_2437,N_436);
and U4365 (N_4365,N_2227,N_1132);
and U4366 (N_4366,N_2207,N_925);
nor U4367 (N_4367,N_1582,N_1181);
nand U4368 (N_4368,N_479,N_2331);
and U4369 (N_4369,N_1632,N_2272);
nor U4370 (N_4370,N_1450,N_277);
and U4371 (N_4371,N_2373,N_434);
or U4372 (N_4372,N_153,N_1940);
and U4373 (N_4373,N_613,N_1035);
nand U4374 (N_4374,N_1270,N_62);
xnor U4375 (N_4375,N_2197,N_1178);
or U4376 (N_4376,N_1640,N_2197);
nor U4377 (N_4377,N_1210,N_2090);
nand U4378 (N_4378,N_440,N_517);
nor U4379 (N_4379,N_385,N_141);
nand U4380 (N_4380,N_47,N_1400);
nor U4381 (N_4381,N_1906,N_572);
nor U4382 (N_4382,N_1519,N_1658);
or U4383 (N_4383,N_2420,N_577);
nor U4384 (N_4384,N_1611,N_2478);
or U4385 (N_4385,N_2036,N_1863);
xnor U4386 (N_4386,N_1758,N_2450);
or U4387 (N_4387,N_2185,N_1368);
and U4388 (N_4388,N_1329,N_1776);
or U4389 (N_4389,N_440,N_2279);
and U4390 (N_4390,N_913,N_1931);
or U4391 (N_4391,N_676,N_429);
or U4392 (N_4392,N_731,N_826);
or U4393 (N_4393,N_385,N_2347);
nand U4394 (N_4394,N_1309,N_536);
or U4395 (N_4395,N_1163,N_255);
or U4396 (N_4396,N_1834,N_362);
nor U4397 (N_4397,N_1489,N_501);
and U4398 (N_4398,N_1195,N_2101);
or U4399 (N_4399,N_1607,N_2140);
nand U4400 (N_4400,N_2493,N_2174);
and U4401 (N_4401,N_1652,N_725);
nand U4402 (N_4402,N_1603,N_2457);
nor U4403 (N_4403,N_1472,N_1077);
and U4404 (N_4404,N_249,N_52);
or U4405 (N_4405,N_508,N_958);
nor U4406 (N_4406,N_1063,N_1013);
xnor U4407 (N_4407,N_1983,N_137);
and U4408 (N_4408,N_117,N_497);
and U4409 (N_4409,N_1073,N_1831);
or U4410 (N_4410,N_2007,N_1850);
nand U4411 (N_4411,N_941,N_1414);
or U4412 (N_4412,N_311,N_90);
xnor U4413 (N_4413,N_2315,N_1126);
xor U4414 (N_4414,N_0,N_722);
nor U4415 (N_4415,N_1938,N_767);
nand U4416 (N_4416,N_1400,N_538);
nor U4417 (N_4417,N_1669,N_1104);
nor U4418 (N_4418,N_514,N_412);
nor U4419 (N_4419,N_2046,N_566);
xnor U4420 (N_4420,N_442,N_348);
and U4421 (N_4421,N_434,N_2332);
nor U4422 (N_4422,N_83,N_773);
and U4423 (N_4423,N_1932,N_2005);
nor U4424 (N_4424,N_337,N_1640);
and U4425 (N_4425,N_2215,N_2246);
and U4426 (N_4426,N_2428,N_132);
and U4427 (N_4427,N_1139,N_2309);
nor U4428 (N_4428,N_384,N_1576);
or U4429 (N_4429,N_1884,N_1069);
and U4430 (N_4430,N_1795,N_1785);
nor U4431 (N_4431,N_2124,N_1462);
nor U4432 (N_4432,N_1564,N_663);
xnor U4433 (N_4433,N_671,N_654);
nand U4434 (N_4434,N_1548,N_167);
xnor U4435 (N_4435,N_844,N_772);
nor U4436 (N_4436,N_2203,N_936);
and U4437 (N_4437,N_2150,N_1809);
xor U4438 (N_4438,N_2391,N_1469);
or U4439 (N_4439,N_1734,N_1259);
nand U4440 (N_4440,N_1208,N_1381);
or U4441 (N_4441,N_2095,N_385);
and U4442 (N_4442,N_2027,N_642);
nor U4443 (N_4443,N_229,N_2174);
nand U4444 (N_4444,N_1714,N_1087);
xor U4445 (N_4445,N_1720,N_783);
or U4446 (N_4446,N_2353,N_670);
or U4447 (N_4447,N_1600,N_1317);
nor U4448 (N_4448,N_848,N_16);
nand U4449 (N_4449,N_1326,N_265);
xor U4450 (N_4450,N_1824,N_2026);
or U4451 (N_4451,N_1938,N_1719);
or U4452 (N_4452,N_2036,N_2181);
nor U4453 (N_4453,N_1514,N_1040);
and U4454 (N_4454,N_2422,N_1718);
or U4455 (N_4455,N_545,N_188);
xnor U4456 (N_4456,N_2389,N_1441);
nor U4457 (N_4457,N_1069,N_2433);
or U4458 (N_4458,N_631,N_1589);
or U4459 (N_4459,N_2417,N_1527);
and U4460 (N_4460,N_1746,N_465);
xnor U4461 (N_4461,N_2157,N_1707);
xor U4462 (N_4462,N_1497,N_2405);
nand U4463 (N_4463,N_1109,N_1646);
and U4464 (N_4464,N_1321,N_2449);
or U4465 (N_4465,N_370,N_2279);
nand U4466 (N_4466,N_1716,N_1129);
nor U4467 (N_4467,N_2063,N_685);
xnor U4468 (N_4468,N_1341,N_157);
nand U4469 (N_4469,N_322,N_1751);
nor U4470 (N_4470,N_1968,N_1908);
nand U4471 (N_4471,N_2041,N_1006);
nand U4472 (N_4472,N_2155,N_57);
nand U4473 (N_4473,N_1006,N_1642);
and U4474 (N_4474,N_1402,N_2330);
and U4475 (N_4475,N_1014,N_1175);
or U4476 (N_4476,N_985,N_990);
and U4477 (N_4477,N_1050,N_923);
and U4478 (N_4478,N_269,N_2409);
or U4479 (N_4479,N_2328,N_1178);
or U4480 (N_4480,N_2148,N_2328);
and U4481 (N_4481,N_408,N_1195);
xor U4482 (N_4482,N_2156,N_277);
nor U4483 (N_4483,N_1737,N_1341);
and U4484 (N_4484,N_690,N_534);
nand U4485 (N_4485,N_2142,N_543);
or U4486 (N_4486,N_1178,N_1352);
nand U4487 (N_4487,N_1150,N_417);
or U4488 (N_4488,N_192,N_655);
nand U4489 (N_4489,N_1481,N_817);
nor U4490 (N_4490,N_976,N_43);
and U4491 (N_4491,N_394,N_176);
nand U4492 (N_4492,N_2300,N_1376);
and U4493 (N_4493,N_406,N_950);
and U4494 (N_4494,N_221,N_2039);
nor U4495 (N_4495,N_1534,N_1505);
xnor U4496 (N_4496,N_1123,N_487);
nor U4497 (N_4497,N_1218,N_2428);
and U4498 (N_4498,N_2334,N_1597);
and U4499 (N_4499,N_906,N_288);
or U4500 (N_4500,N_2130,N_1271);
nand U4501 (N_4501,N_1625,N_623);
xor U4502 (N_4502,N_10,N_20);
or U4503 (N_4503,N_511,N_293);
and U4504 (N_4504,N_2184,N_2078);
nand U4505 (N_4505,N_224,N_1506);
or U4506 (N_4506,N_919,N_703);
nand U4507 (N_4507,N_1543,N_858);
and U4508 (N_4508,N_1210,N_1906);
or U4509 (N_4509,N_1877,N_1727);
and U4510 (N_4510,N_1747,N_1345);
nor U4511 (N_4511,N_450,N_2151);
and U4512 (N_4512,N_158,N_673);
nor U4513 (N_4513,N_2300,N_2018);
and U4514 (N_4514,N_1645,N_1190);
nand U4515 (N_4515,N_1169,N_1201);
and U4516 (N_4516,N_221,N_2230);
and U4517 (N_4517,N_2443,N_1108);
xor U4518 (N_4518,N_2240,N_873);
nand U4519 (N_4519,N_549,N_104);
nand U4520 (N_4520,N_516,N_2282);
or U4521 (N_4521,N_1820,N_234);
xnor U4522 (N_4522,N_1156,N_1131);
nand U4523 (N_4523,N_895,N_662);
and U4524 (N_4524,N_1141,N_776);
or U4525 (N_4525,N_2195,N_968);
or U4526 (N_4526,N_66,N_2251);
and U4527 (N_4527,N_1295,N_1512);
nand U4528 (N_4528,N_2327,N_1041);
and U4529 (N_4529,N_2092,N_126);
nand U4530 (N_4530,N_1224,N_468);
and U4531 (N_4531,N_1818,N_1223);
xnor U4532 (N_4532,N_913,N_817);
xor U4533 (N_4533,N_366,N_1434);
nand U4534 (N_4534,N_131,N_343);
and U4535 (N_4535,N_514,N_2308);
and U4536 (N_4536,N_2424,N_2143);
nor U4537 (N_4537,N_2163,N_1261);
and U4538 (N_4538,N_856,N_638);
and U4539 (N_4539,N_68,N_501);
nand U4540 (N_4540,N_1407,N_2103);
xnor U4541 (N_4541,N_18,N_1445);
nor U4542 (N_4542,N_758,N_523);
nor U4543 (N_4543,N_887,N_2477);
nor U4544 (N_4544,N_1301,N_720);
or U4545 (N_4545,N_1713,N_741);
xnor U4546 (N_4546,N_2425,N_1926);
nor U4547 (N_4547,N_2114,N_2467);
nor U4548 (N_4548,N_647,N_1328);
and U4549 (N_4549,N_1509,N_399);
and U4550 (N_4550,N_2162,N_239);
nand U4551 (N_4551,N_337,N_1712);
xnor U4552 (N_4552,N_1730,N_643);
nand U4553 (N_4553,N_1858,N_451);
nand U4554 (N_4554,N_2402,N_615);
nand U4555 (N_4555,N_2435,N_414);
and U4556 (N_4556,N_433,N_636);
or U4557 (N_4557,N_1616,N_1337);
and U4558 (N_4558,N_1062,N_1993);
nand U4559 (N_4559,N_1747,N_185);
or U4560 (N_4560,N_2202,N_1393);
and U4561 (N_4561,N_1096,N_2418);
nor U4562 (N_4562,N_2159,N_1071);
nand U4563 (N_4563,N_466,N_2396);
nor U4564 (N_4564,N_104,N_894);
nor U4565 (N_4565,N_1905,N_1796);
nand U4566 (N_4566,N_2296,N_89);
nand U4567 (N_4567,N_922,N_1278);
or U4568 (N_4568,N_397,N_1029);
or U4569 (N_4569,N_1725,N_1669);
and U4570 (N_4570,N_311,N_166);
nand U4571 (N_4571,N_534,N_2329);
and U4572 (N_4572,N_1141,N_1222);
nor U4573 (N_4573,N_870,N_877);
or U4574 (N_4574,N_491,N_1777);
or U4575 (N_4575,N_912,N_1639);
and U4576 (N_4576,N_542,N_2460);
or U4577 (N_4577,N_2402,N_2179);
and U4578 (N_4578,N_1616,N_2368);
nor U4579 (N_4579,N_2160,N_1288);
nand U4580 (N_4580,N_609,N_394);
and U4581 (N_4581,N_216,N_2136);
and U4582 (N_4582,N_2296,N_526);
and U4583 (N_4583,N_658,N_1425);
nand U4584 (N_4584,N_1367,N_784);
and U4585 (N_4585,N_411,N_988);
nor U4586 (N_4586,N_2309,N_796);
nand U4587 (N_4587,N_1492,N_2004);
nand U4588 (N_4588,N_715,N_448);
and U4589 (N_4589,N_2134,N_2084);
or U4590 (N_4590,N_92,N_566);
or U4591 (N_4591,N_1855,N_2179);
and U4592 (N_4592,N_1636,N_1504);
nand U4593 (N_4593,N_266,N_668);
nand U4594 (N_4594,N_1475,N_2373);
nor U4595 (N_4595,N_1234,N_37);
or U4596 (N_4596,N_413,N_657);
nand U4597 (N_4597,N_2340,N_1450);
and U4598 (N_4598,N_1945,N_1070);
or U4599 (N_4599,N_1125,N_920);
or U4600 (N_4600,N_1144,N_2482);
or U4601 (N_4601,N_2267,N_2066);
or U4602 (N_4602,N_92,N_357);
nor U4603 (N_4603,N_2267,N_1582);
and U4604 (N_4604,N_2455,N_1840);
and U4605 (N_4605,N_1964,N_1280);
and U4606 (N_4606,N_604,N_459);
or U4607 (N_4607,N_1365,N_1320);
and U4608 (N_4608,N_745,N_1684);
nor U4609 (N_4609,N_2188,N_2491);
and U4610 (N_4610,N_487,N_1831);
nor U4611 (N_4611,N_1880,N_894);
nand U4612 (N_4612,N_2459,N_259);
or U4613 (N_4613,N_151,N_26);
or U4614 (N_4614,N_1719,N_1457);
nor U4615 (N_4615,N_962,N_121);
or U4616 (N_4616,N_1724,N_324);
xor U4617 (N_4617,N_2427,N_750);
and U4618 (N_4618,N_507,N_2440);
and U4619 (N_4619,N_1403,N_1519);
nor U4620 (N_4620,N_242,N_1283);
and U4621 (N_4621,N_843,N_446);
xor U4622 (N_4622,N_1030,N_1283);
nor U4623 (N_4623,N_297,N_1874);
nor U4624 (N_4624,N_1715,N_2292);
or U4625 (N_4625,N_2132,N_1007);
and U4626 (N_4626,N_2323,N_456);
and U4627 (N_4627,N_3,N_1502);
and U4628 (N_4628,N_40,N_2315);
nand U4629 (N_4629,N_125,N_1174);
or U4630 (N_4630,N_2313,N_2478);
xor U4631 (N_4631,N_2074,N_60);
nor U4632 (N_4632,N_342,N_1324);
or U4633 (N_4633,N_682,N_2225);
nor U4634 (N_4634,N_2352,N_2102);
and U4635 (N_4635,N_2438,N_1224);
or U4636 (N_4636,N_640,N_2023);
or U4637 (N_4637,N_2063,N_178);
nor U4638 (N_4638,N_480,N_777);
or U4639 (N_4639,N_1564,N_1421);
nand U4640 (N_4640,N_480,N_641);
nand U4641 (N_4641,N_1682,N_2295);
and U4642 (N_4642,N_2229,N_1761);
nand U4643 (N_4643,N_937,N_595);
or U4644 (N_4644,N_448,N_71);
xnor U4645 (N_4645,N_1600,N_722);
or U4646 (N_4646,N_1474,N_982);
nor U4647 (N_4647,N_1671,N_1388);
and U4648 (N_4648,N_344,N_1475);
or U4649 (N_4649,N_1316,N_2435);
nand U4650 (N_4650,N_2393,N_1672);
xor U4651 (N_4651,N_19,N_1649);
and U4652 (N_4652,N_1016,N_1547);
nand U4653 (N_4653,N_267,N_618);
nand U4654 (N_4654,N_34,N_1661);
or U4655 (N_4655,N_290,N_1043);
nand U4656 (N_4656,N_1533,N_2080);
and U4657 (N_4657,N_881,N_1426);
nor U4658 (N_4658,N_297,N_1384);
and U4659 (N_4659,N_634,N_1156);
nand U4660 (N_4660,N_2166,N_292);
nand U4661 (N_4661,N_130,N_241);
nor U4662 (N_4662,N_744,N_797);
or U4663 (N_4663,N_2431,N_231);
nor U4664 (N_4664,N_787,N_887);
or U4665 (N_4665,N_1961,N_1373);
xor U4666 (N_4666,N_1247,N_1184);
and U4667 (N_4667,N_965,N_1335);
and U4668 (N_4668,N_476,N_1271);
nor U4669 (N_4669,N_640,N_75);
nor U4670 (N_4670,N_1755,N_1503);
and U4671 (N_4671,N_1294,N_2300);
or U4672 (N_4672,N_1368,N_1075);
nand U4673 (N_4673,N_1089,N_1842);
nand U4674 (N_4674,N_1218,N_484);
xor U4675 (N_4675,N_1920,N_101);
nor U4676 (N_4676,N_1670,N_444);
xnor U4677 (N_4677,N_1551,N_82);
nand U4678 (N_4678,N_1121,N_1153);
nand U4679 (N_4679,N_952,N_329);
and U4680 (N_4680,N_1686,N_4);
nor U4681 (N_4681,N_2137,N_1597);
nand U4682 (N_4682,N_2194,N_1964);
nor U4683 (N_4683,N_266,N_1740);
and U4684 (N_4684,N_1634,N_672);
or U4685 (N_4685,N_1160,N_1695);
xnor U4686 (N_4686,N_592,N_1770);
nor U4687 (N_4687,N_543,N_1585);
or U4688 (N_4688,N_2480,N_2415);
and U4689 (N_4689,N_327,N_2451);
nand U4690 (N_4690,N_323,N_153);
nand U4691 (N_4691,N_326,N_2237);
nand U4692 (N_4692,N_2222,N_288);
and U4693 (N_4693,N_1283,N_983);
or U4694 (N_4694,N_1206,N_1835);
or U4695 (N_4695,N_925,N_1180);
nand U4696 (N_4696,N_119,N_2249);
or U4697 (N_4697,N_2191,N_2090);
xnor U4698 (N_4698,N_1183,N_380);
and U4699 (N_4699,N_2261,N_1304);
or U4700 (N_4700,N_395,N_2004);
nor U4701 (N_4701,N_816,N_1404);
nor U4702 (N_4702,N_1790,N_332);
nor U4703 (N_4703,N_1236,N_767);
nor U4704 (N_4704,N_2259,N_1688);
and U4705 (N_4705,N_242,N_2183);
xnor U4706 (N_4706,N_1381,N_211);
nor U4707 (N_4707,N_491,N_2110);
or U4708 (N_4708,N_1898,N_1978);
nor U4709 (N_4709,N_206,N_1697);
nor U4710 (N_4710,N_1555,N_736);
and U4711 (N_4711,N_1110,N_1200);
nor U4712 (N_4712,N_879,N_1523);
nand U4713 (N_4713,N_1810,N_311);
and U4714 (N_4714,N_533,N_481);
and U4715 (N_4715,N_1450,N_1198);
and U4716 (N_4716,N_1380,N_1801);
nor U4717 (N_4717,N_332,N_428);
nand U4718 (N_4718,N_62,N_2072);
and U4719 (N_4719,N_1910,N_1742);
nor U4720 (N_4720,N_900,N_341);
nor U4721 (N_4721,N_1845,N_673);
and U4722 (N_4722,N_447,N_2480);
xor U4723 (N_4723,N_409,N_272);
and U4724 (N_4724,N_1545,N_510);
nor U4725 (N_4725,N_1913,N_2129);
nor U4726 (N_4726,N_897,N_2163);
or U4727 (N_4727,N_1447,N_702);
nand U4728 (N_4728,N_397,N_2307);
nor U4729 (N_4729,N_1767,N_2366);
nand U4730 (N_4730,N_51,N_560);
and U4731 (N_4731,N_1008,N_1365);
or U4732 (N_4732,N_1756,N_2430);
nand U4733 (N_4733,N_666,N_1650);
nor U4734 (N_4734,N_1739,N_1061);
or U4735 (N_4735,N_736,N_1954);
nor U4736 (N_4736,N_2237,N_2072);
or U4737 (N_4737,N_2164,N_833);
nor U4738 (N_4738,N_1793,N_1736);
nand U4739 (N_4739,N_822,N_1513);
nand U4740 (N_4740,N_2289,N_787);
and U4741 (N_4741,N_773,N_1105);
nor U4742 (N_4742,N_330,N_2234);
or U4743 (N_4743,N_1896,N_2018);
and U4744 (N_4744,N_838,N_693);
xor U4745 (N_4745,N_2473,N_2102);
nand U4746 (N_4746,N_557,N_454);
nand U4747 (N_4747,N_1519,N_1791);
xor U4748 (N_4748,N_2057,N_351);
nand U4749 (N_4749,N_131,N_207);
nand U4750 (N_4750,N_556,N_752);
and U4751 (N_4751,N_958,N_95);
nor U4752 (N_4752,N_764,N_1616);
and U4753 (N_4753,N_1719,N_425);
and U4754 (N_4754,N_251,N_2345);
or U4755 (N_4755,N_1910,N_1316);
and U4756 (N_4756,N_1261,N_2285);
or U4757 (N_4757,N_292,N_1270);
nand U4758 (N_4758,N_279,N_1504);
or U4759 (N_4759,N_535,N_1483);
nor U4760 (N_4760,N_627,N_1705);
and U4761 (N_4761,N_80,N_115);
or U4762 (N_4762,N_1050,N_1408);
and U4763 (N_4763,N_428,N_551);
nor U4764 (N_4764,N_353,N_2389);
or U4765 (N_4765,N_450,N_1979);
nor U4766 (N_4766,N_664,N_123);
xnor U4767 (N_4767,N_518,N_392);
nand U4768 (N_4768,N_1792,N_1642);
and U4769 (N_4769,N_806,N_2215);
nand U4770 (N_4770,N_1246,N_1458);
and U4771 (N_4771,N_2430,N_2099);
and U4772 (N_4772,N_1424,N_873);
and U4773 (N_4773,N_228,N_91);
and U4774 (N_4774,N_601,N_1156);
nor U4775 (N_4775,N_764,N_374);
nand U4776 (N_4776,N_1358,N_2485);
or U4777 (N_4777,N_935,N_727);
and U4778 (N_4778,N_609,N_1362);
and U4779 (N_4779,N_556,N_2214);
and U4780 (N_4780,N_1996,N_1554);
nand U4781 (N_4781,N_336,N_2252);
or U4782 (N_4782,N_1827,N_507);
and U4783 (N_4783,N_1406,N_690);
nor U4784 (N_4784,N_388,N_1709);
nor U4785 (N_4785,N_3,N_1111);
nor U4786 (N_4786,N_178,N_2116);
and U4787 (N_4787,N_1339,N_1508);
or U4788 (N_4788,N_1115,N_1252);
or U4789 (N_4789,N_696,N_2122);
or U4790 (N_4790,N_2221,N_66);
nor U4791 (N_4791,N_1759,N_1150);
or U4792 (N_4792,N_1766,N_486);
nand U4793 (N_4793,N_1158,N_625);
and U4794 (N_4794,N_1698,N_1780);
nand U4795 (N_4795,N_957,N_5);
and U4796 (N_4796,N_2153,N_947);
and U4797 (N_4797,N_318,N_1343);
and U4798 (N_4798,N_882,N_1092);
or U4799 (N_4799,N_298,N_2249);
or U4800 (N_4800,N_2364,N_522);
or U4801 (N_4801,N_2417,N_2446);
and U4802 (N_4802,N_870,N_1228);
or U4803 (N_4803,N_2416,N_96);
and U4804 (N_4804,N_936,N_49);
nor U4805 (N_4805,N_1228,N_1940);
nor U4806 (N_4806,N_2294,N_1127);
nor U4807 (N_4807,N_1663,N_1012);
and U4808 (N_4808,N_2116,N_991);
nand U4809 (N_4809,N_232,N_492);
nand U4810 (N_4810,N_1013,N_265);
or U4811 (N_4811,N_1658,N_63);
nand U4812 (N_4812,N_369,N_2497);
nand U4813 (N_4813,N_166,N_467);
or U4814 (N_4814,N_1889,N_915);
and U4815 (N_4815,N_51,N_293);
xnor U4816 (N_4816,N_62,N_1001);
and U4817 (N_4817,N_2239,N_380);
nor U4818 (N_4818,N_315,N_332);
nand U4819 (N_4819,N_849,N_1614);
nor U4820 (N_4820,N_2421,N_2217);
or U4821 (N_4821,N_486,N_724);
nor U4822 (N_4822,N_849,N_1211);
nor U4823 (N_4823,N_1446,N_2430);
or U4824 (N_4824,N_2025,N_383);
or U4825 (N_4825,N_2306,N_252);
nand U4826 (N_4826,N_2493,N_1617);
and U4827 (N_4827,N_11,N_1752);
nand U4828 (N_4828,N_1743,N_1213);
nand U4829 (N_4829,N_1333,N_966);
or U4830 (N_4830,N_2046,N_2137);
xor U4831 (N_4831,N_2206,N_38);
nor U4832 (N_4832,N_75,N_1475);
and U4833 (N_4833,N_1605,N_2491);
or U4834 (N_4834,N_1837,N_569);
or U4835 (N_4835,N_269,N_1478);
and U4836 (N_4836,N_2485,N_1006);
xor U4837 (N_4837,N_1358,N_1697);
or U4838 (N_4838,N_2246,N_617);
nand U4839 (N_4839,N_1009,N_819);
and U4840 (N_4840,N_1488,N_1943);
xnor U4841 (N_4841,N_2087,N_904);
or U4842 (N_4842,N_453,N_174);
or U4843 (N_4843,N_18,N_195);
and U4844 (N_4844,N_1371,N_668);
and U4845 (N_4845,N_2124,N_1134);
and U4846 (N_4846,N_1490,N_2124);
or U4847 (N_4847,N_448,N_1896);
or U4848 (N_4848,N_1777,N_954);
and U4849 (N_4849,N_1374,N_1065);
nor U4850 (N_4850,N_29,N_2220);
nand U4851 (N_4851,N_1357,N_1598);
and U4852 (N_4852,N_882,N_1785);
nor U4853 (N_4853,N_886,N_2061);
nor U4854 (N_4854,N_930,N_1075);
or U4855 (N_4855,N_2448,N_989);
nand U4856 (N_4856,N_353,N_1883);
and U4857 (N_4857,N_607,N_911);
or U4858 (N_4858,N_1675,N_243);
and U4859 (N_4859,N_61,N_192);
nand U4860 (N_4860,N_2479,N_70);
and U4861 (N_4861,N_1037,N_2263);
nand U4862 (N_4862,N_468,N_1175);
nor U4863 (N_4863,N_1772,N_793);
xor U4864 (N_4864,N_2291,N_44);
xnor U4865 (N_4865,N_774,N_1984);
or U4866 (N_4866,N_1170,N_351);
nor U4867 (N_4867,N_1327,N_346);
nor U4868 (N_4868,N_2016,N_734);
nand U4869 (N_4869,N_2409,N_1097);
or U4870 (N_4870,N_1310,N_418);
or U4871 (N_4871,N_2107,N_2060);
or U4872 (N_4872,N_2047,N_1530);
nand U4873 (N_4873,N_745,N_517);
or U4874 (N_4874,N_916,N_202);
and U4875 (N_4875,N_2150,N_351);
nor U4876 (N_4876,N_621,N_485);
and U4877 (N_4877,N_1472,N_1931);
xor U4878 (N_4878,N_2196,N_932);
nand U4879 (N_4879,N_1931,N_2375);
nand U4880 (N_4880,N_609,N_2433);
nor U4881 (N_4881,N_2357,N_1065);
nor U4882 (N_4882,N_2311,N_185);
and U4883 (N_4883,N_2201,N_2188);
or U4884 (N_4884,N_817,N_1932);
and U4885 (N_4885,N_1888,N_259);
or U4886 (N_4886,N_919,N_2381);
nor U4887 (N_4887,N_317,N_2281);
nor U4888 (N_4888,N_1177,N_962);
nor U4889 (N_4889,N_20,N_1978);
or U4890 (N_4890,N_1143,N_678);
nor U4891 (N_4891,N_8,N_1517);
nand U4892 (N_4892,N_506,N_723);
nor U4893 (N_4893,N_1362,N_1176);
nor U4894 (N_4894,N_2083,N_150);
and U4895 (N_4895,N_651,N_1464);
nand U4896 (N_4896,N_2083,N_1395);
nor U4897 (N_4897,N_2129,N_2056);
nor U4898 (N_4898,N_829,N_1789);
and U4899 (N_4899,N_1649,N_2151);
or U4900 (N_4900,N_2078,N_1056);
and U4901 (N_4901,N_109,N_331);
and U4902 (N_4902,N_906,N_140);
and U4903 (N_4903,N_1049,N_648);
xor U4904 (N_4904,N_872,N_997);
nand U4905 (N_4905,N_1713,N_1649);
nor U4906 (N_4906,N_380,N_1347);
and U4907 (N_4907,N_585,N_1603);
or U4908 (N_4908,N_899,N_1664);
nand U4909 (N_4909,N_2093,N_2198);
or U4910 (N_4910,N_1640,N_2291);
or U4911 (N_4911,N_299,N_1835);
and U4912 (N_4912,N_875,N_804);
or U4913 (N_4913,N_305,N_2070);
or U4914 (N_4914,N_164,N_2397);
nor U4915 (N_4915,N_1723,N_187);
or U4916 (N_4916,N_698,N_2438);
or U4917 (N_4917,N_140,N_631);
nand U4918 (N_4918,N_715,N_845);
or U4919 (N_4919,N_1470,N_382);
nor U4920 (N_4920,N_539,N_1549);
or U4921 (N_4921,N_2034,N_1605);
nand U4922 (N_4922,N_635,N_1480);
xor U4923 (N_4923,N_390,N_991);
and U4924 (N_4924,N_2158,N_736);
and U4925 (N_4925,N_1531,N_1517);
and U4926 (N_4926,N_2193,N_1561);
nor U4927 (N_4927,N_1271,N_606);
xor U4928 (N_4928,N_538,N_1690);
or U4929 (N_4929,N_1059,N_498);
nor U4930 (N_4930,N_1740,N_1471);
or U4931 (N_4931,N_563,N_715);
xnor U4932 (N_4932,N_741,N_259);
and U4933 (N_4933,N_2121,N_1139);
nand U4934 (N_4934,N_2228,N_1849);
or U4935 (N_4935,N_353,N_98);
nand U4936 (N_4936,N_204,N_1605);
nor U4937 (N_4937,N_879,N_1750);
and U4938 (N_4938,N_1402,N_9);
nand U4939 (N_4939,N_261,N_463);
and U4940 (N_4940,N_877,N_2432);
nand U4941 (N_4941,N_1793,N_2481);
nor U4942 (N_4942,N_647,N_2040);
xnor U4943 (N_4943,N_2155,N_1074);
and U4944 (N_4944,N_778,N_600);
nor U4945 (N_4945,N_1475,N_1610);
nand U4946 (N_4946,N_1540,N_2278);
nand U4947 (N_4947,N_1347,N_1877);
nand U4948 (N_4948,N_176,N_1954);
or U4949 (N_4949,N_1771,N_1782);
nor U4950 (N_4950,N_1019,N_736);
and U4951 (N_4951,N_1774,N_729);
and U4952 (N_4952,N_496,N_847);
or U4953 (N_4953,N_2452,N_90);
and U4954 (N_4954,N_1436,N_1803);
xor U4955 (N_4955,N_1748,N_1418);
or U4956 (N_4956,N_1336,N_352);
nor U4957 (N_4957,N_1561,N_1620);
nor U4958 (N_4958,N_557,N_57);
xnor U4959 (N_4959,N_2433,N_1238);
xnor U4960 (N_4960,N_1773,N_920);
or U4961 (N_4961,N_2401,N_1713);
or U4962 (N_4962,N_1785,N_1012);
or U4963 (N_4963,N_2392,N_417);
nor U4964 (N_4964,N_1323,N_1013);
or U4965 (N_4965,N_2252,N_1823);
and U4966 (N_4966,N_981,N_2439);
nand U4967 (N_4967,N_174,N_1054);
nand U4968 (N_4968,N_1578,N_789);
nand U4969 (N_4969,N_1061,N_1685);
nand U4970 (N_4970,N_36,N_2005);
nand U4971 (N_4971,N_2305,N_809);
nand U4972 (N_4972,N_251,N_1338);
and U4973 (N_4973,N_129,N_2403);
and U4974 (N_4974,N_719,N_855);
nor U4975 (N_4975,N_607,N_342);
and U4976 (N_4976,N_1877,N_294);
nor U4977 (N_4977,N_138,N_118);
nor U4978 (N_4978,N_2085,N_442);
xnor U4979 (N_4979,N_1278,N_2004);
nor U4980 (N_4980,N_1571,N_376);
nor U4981 (N_4981,N_1869,N_2303);
nor U4982 (N_4982,N_2280,N_1238);
nand U4983 (N_4983,N_235,N_1477);
nor U4984 (N_4984,N_2235,N_1063);
xnor U4985 (N_4985,N_2105,N_871);
and U4986 (N_4986,N_1170,N_1079);
or U4987 (N_4987,N_44,N_1615);
nand U4988 (N_4988,N_2087,N_2262);
and U4989 (N_4989,N_1961,N_1385);
or U4990 (N_4990,N_378,N_1222);
and U4991 (N_4991,N_438,N_1004);
or U4992 (N_4992,N_1723,N_396);
and U4993 (N_4993,N_315,N_615);
nand U4994 (N_4994,N_1011,N_574);
nor U4995 (N_4995,N_1963,N_1701);
xor U4996 (N_4996,N_553,N_1037);
nand U4997 (N_4997,N_1871,N_1475);
nor U4998 (N_4998,N_1347,N_1550);
and U4999 (N_4999,N_173,N_1974);
nor U5000 (N_5000,N_2901,N_3920);
and U5001 (N_5001,N_4762,N_4529);
and U5002 (N_5002,N_4483,N_3691);
nor U5003 (N_5003,N_4871,N_2632);
nor U5004 (N_5004,N_4447,N_3972);
or U5005 (N_5005,N_4864,N_4884);
or U5006 (N_5006,N_2765,N_3708);
xor U5007 (N_5007,N_2665,N_4364);
nand U5008 (N_5008,N_3176,N_4831);
and U5009 (N_5009,N_4528,N_4564);
nor U5010 (N_5010,N_3990,N_4050);
nand U5011 (N_5011,N_2899,N_2880);
nor U5012 (N_5012,N_3051,N_3649);
nor U5013 (N_5013,N_2997,N_3588);
nor U5014 (N_5014,N_4499,N_4627);
nor U5015 (N_5015,N_3574,N_3712);
nand U5016 (N_5016,N_2885,N_4332);
nand U5017 (N_5017,N_3799,N_3215);
nor U5018 (N_5018,N_3887,N_3983);
and U5019 (N_5019,N_2683,N_3981);
xnor U5020 (N_5020,N_4934,N_4127);
nor U5021 (N_5021,N_2930,N_4786);
nand U5022 (N_5022,N_3303,N_4570);
and U5023 (N_5023,N_4362,N_4738);
or U5024 (N_5024,N_3808,N_4316);
and U5025 (N_5025,N_4698,N_2769);
xnor U5026 (N_5026,N_4343,N_4084);
and U5027 (N_5027,N_4446,N_4741);
nand U5028 (N_5028,N_3723,N_4173);
and U5029 (N_5029,N_3170,N_4792);
nor U5030 (N_5030,N_4730,N_4417);
or U5031 (N_5031,N_3495,N_3470);
nor U5032 (N_5032,N_4633,N_2840);
nor U5033 (N_5033,N_2964,N_3444);
or U5034 (N_5034,N_3336,N_3753);
nor U5035 (N_5035,N_3914,N_3738);
nor U5036 (N_5036,N_4830,N_3288);
or U5037 (N_5037,N_3224,N_4977);
xor U5038 (N_5038,N_2920,N_4097);
nor U5039 (N_5039,N_3474,N_3988);
and U5040 (N_5040,N_2659,N_4733);
nor U5041 (N_5041,N_4183,N_4628);
nor U5042 (N_5042,N_4102,N_3366);
xnor U5043 (N_5043,N_2688,N_4828);
or U5044 (N_5044,N_4927,N_4898);
nand U5045 (N_5045,N_4163,N_2762);
and U5046 (N_5046,N_4162,N_4487);
and U5047 (N_5047,N_2503,N_4651);
or U5048 (N_5048,N_4011,N_3824);
nand U5049 (N_5049,N_4081,N_3012);
nand U5050 (N_5050,N_4583,N_3609);
nor U5051 (N_5051,N_3938,N_3802);
nand U5052 (N_5052,N_3544,N_2676);
nor U5053 (N_5053,N_3504,N_2722);
or U5054 (N_5054,N_3459,N_4506);
or U5055 (N_5055,N_2785,N_4206);
nor U5056 (N_5056,N_2544,N_3745);
nor U5057 (N_5057,N_3950,N_2981);
nor U5058 (N_5058,N_2599,N_3897);
or U5059 (N_5059,N_2783,N_3764);
xor U5060 (N_5060,N_2628,N_2772);
or U5061 (N_5061,N_2979,N_3271);
nand U5062 (N_5062,N_3228,N_2693);
nor U5063 (N_5063,N_4375,N_3558);
xor U5064 (N_5064,N_4571,N_4134);
xor U5065 (N_5065,N_2998,N_2802);
or U5066 (N_5066,N_4582,N_3446);
nand U5067 (N_5067,N_4153,N_4405);
and U5068 (N_5068,N_2633,N_3326);
xor U5069 (N_5069,N_4608,N_2790);
and U5070 (N_5070,N_4580,N_4983);
or U5071 (N_5071,N_4881,N_3883);
nor U5072 (N_5072,N_2839,N_4131);
and U5073 (N_5073,N_3557,N_4002);
or U5074 (N_5074,N_2916,N_2625);
nor U5075 (N_5075,N_3255,N_4363);
nand U5076 (N_5076,N_3334,N_4620);
and U5077 (N_5077,N_4240,N_2572);
and U5078 (N_5078,N_4460,N_4559);
or U5079 (N_5079,N_4524,N_3299);
nand U5080 (N_5080,N_2699,N_4222);
nand U5081 (N_5081,N_3651,N_3715);
and U5082 (N_5082,N_3554,N_3596);
nand U5083 (N_5083,N_3128,N_4114);
or U5084 (N_5084,N_4243,N_3243);
nand U5085 (N_5085,N_4176,N_4412);
nand U5086 (N_5086,N_2908,N_4951);
nand U5087 (N_5087,N_4797,N_2536);
or U5088 (N_5088,N_4817,N_4381);
nand U5089 (N_5089,N_2520,N_4691);
nand U5090 (N_5090,N_4937,N_4833);
nand U5091 (N_5091,N_2977,N_3076);
or U5092 (N_5092,N_3491,N_4954);
nor U5093 (N_5093,N_3941,N_3142);
nand U5094 (N_5094,N_2975,N_3355);
and U5095 (N_5095,N_4140,N_4949);
nand U5096 (N_5096,N_4754,N_4160);
nand U5097 (N_5097,N_3817,N_3820);
and U5098 (N_5098,N_2939,N_3185);
and U5099 (N_5099,N_2960,N_3534);
and U5100 (N_5100,N_2959,N_2866);
and U5101 (N_5101,N_4029,N_4471);
or U5102 (N_5102,N_3093,N_4040);
or U5103 (N_5103,N_3907,N_3891);
or U5104 (N_5104,N_3116,N_3767);
nor U5105 (N_5105,N_3452,N_2587);
nor U5106 (N_5106,N_4530,N_4398);
xnor U5107 (N_5107,N_4109,N_4148);
or U5108 (N_5108,N_4648,N_3810);
nand U5109 (N_5109,N_2940,N_2630);
nand U5110 (N_5110,N_2661,N_3540);
and U5111 (N_5111,N_2622,N_4070);
nor U5112 (N_5112,N_3893,N_4527);
and U5113 (N_5113,N_4455,N_2867);
nor U5114 (N_5114,N_3594,N_3484);
nor U5115 (N_5115,N_4875,N_2576);
nand U5116 (N_5116,N_4277,N_3351);
and U5117 (N_5117,N_3209,N_3026);
nand U5118 (N_5118,N_2923,N_2974);
and U5119 (N_5119,N_3912,N_4517);
nor U5120 (N_5120,N_4345,N_4264);
and U5121 (N_5121,N_2517,N_3790);
nor U5122 (N_5122,N_3377,N_2623);
or U5123 (N_5123,N_4461,N_4861);
or U5124 (N_5124,N_3092,N_4731);
and U5125 (N_5125,N_3348,N_4000);
or U5126 (N_5126,N_2619,N_4966);
or U5127 (N_5127,N_4834,N_3823);
and U5128 (N_5128,N_3875,N_4950);
nor U5129 (N_5129,N_2985,N_3521);
or U5130 (N_5130,N_2640,N_2594);
nand U5131 (N_5131,N_4079,N_4210);
nor U5132 (N_5132,N_4809,N_3561);
xnor U5133 (N_5133,N_3863,N_2600);
or U5134 (N_5134,N_3350,N_3761);
or U5135 (N_5135,N_2680,N_4810);
nand U5136 (N_5136,N_4063,N_4013);
nor U5137 (N_5137,N_3239,N_4172);
or U5138 (N_5138,N_2642,N_2955);
and U5139 (N_5139,N_4065,N_4847);
nand U5140 (N_5140,N_2674,N_3547);
nor U5141 (N_5141,N_3939,N_4435);
xnor U5142 (N_5142,N_4870,N_3368);
nor U5143 (N_5143,N_4494,N_3034);
nor U5144 (N_5144,N_3434,N_4600);
xnor U5145 (N_5145,N_3187,N_4701);
or U5146 (N_5146,N_3214,N_4392);
and U5147 (N_5147,N_3282,N_2716);
and U5148 (N_5148,N_3450,N_4910);
nor U5149 (N_5149,N_4760,N_4464);
xor U5150 (N_5150,N_2730,N_4010);
nor U5151 (N_5151,N_4567,N_4561);
nor U5152 (N_5152,N_4028,N_2666);
xnor U5153 (N_5153,N_4214,N_4819);
or U5154 (N_5154,N_4226,N_2822);
or U5155 (N_5155,N_3843,N_3155);
nor U5156 (N_5156,N_4548,N_2580);
nor U5157 (N_5157,N_4024,N_3086);
nand U5158 (N_5158,N_4250,N_4837);
xnor U5159 (N_5159,N_4051,N_3762);
or U5160 (N_5160,N_4686,N_4033);
and U5161 (N_5161,N_3236,N_2675);
nor U5162 (N_5162,N_2538,N_4019);
nand U5163 (N_5163,N_4771,N_2582);
nor U5164 (N_5164,N_3993,N_2637);
and U5165 (N_5165,N_4476,N_4192);
nand U5166 (N_5166,N_3453,N_2669);
and U5167 (N_5167,N_4502,N_3970);
nor U5168 (N_5168,N_3017,N_4263);
or U5169 (N_5169,N_4511,N_2747);
or U5170 (N_5170,N_3831,N_2592);
or U5171 (N_5171,N_3905,N_4431);
nor U5172 (N_5172,N_4979,N_3841);
xnor U5173 (N_5173,N_3462,N_4616);
and U5174 (N_5174,N_2558,N_4572);
nand U5175 (N_5175,N_3065,N_4672);
nand U5176 (N_5176,N_4936,N_4347);
or U5177 (N_5177,N_3849,N_3727);
or U5178 (N_5178,N_3565,N_3295);
or U5179 (N_5179,N_4193,N_2821);
xor U5180 (N_5180,N_4613,N_3951);
and U5181 (N_5181,N_4938,N_4371);
and U5182 (N_5182,N_3418,N_4256);
and U5183 (N_5183,N_4198,N_3048);
or U5184 (N_5184,N_2505,N_2968);
or U5185 (N_5185,N_4536,N_4642);
nand U5186 (N_5186,N_3513,N_3158);
nor U5187 (N_5187,N_3748,N_4368);
and U5188 (N_5188,N_2573,N_4787);
and U5189 (N_5189,N_3073,N_3694);
nand U5190 (N_5190,N_4391,N_4619);
or U5191 (N_5191,N_4117,N_4718);
nand U5192 (N_5192,N_3263,N_3156);
nand U5193 (N_5193,N_4926,N_3948);
and U5194 (N_5194,N_3505,N_4166);
nand U5195 (N_5195,N_4423,N_4822);
or U5196 (N_5196,N_3693,N_4301);
nor U5197 (N_5197,N_3947,N_3498);
and U5198 (N_5198,N_2898,N_4728);
xnor U5199 (N_5199,N_4761,N_4299);
nor U5200 (N_5200,N_4129,N_4694);
and U5201 (N_5201,N_3848,N_2915);
and U5202 (N_5202,N_2825,N_4159);
or U5203 (N_5203,N_4308,N_3269);
or U5204 (N_5204,N_2548,N_3408);
or U5205 (N_5205,N_3333,N_3660);
and U5206 (N_5206,N_2712,N_4315);
xnor U5207 (N_5207,N_3909,N_2591);
or U5208 (N_5208,N_3690,N_3743);
and U5209 (N_5209,N_2746,N_3435);
nor U5210 (N_5210,N_2984,N_2937);
and U5211 (N_5211,N_3857,N_3900);
nor U5212 (N_5212,N_2918,N_3159);
or U5213 (N_5213,N_3946,N_3050);
or U5214 (N_5214,N_3667,N_3096);
nand U5215 (N_5215,N_4353,N_3398);
nor U5216 (N_5216,N_3670,N_3283);
nand U5217 (N_5217,N_4071,N_3620);
nand U5218 (N_5218,N_3375,N_3562);
and U5219 (N_5219,N_3056,N_3772);
nor U5220 (N_5220,N_2598,N_3494);
nand U5221 (N_5221,N_3792,N_2635);
nand U5222 (N_5222,N_2956,N_3613);
nand U5223 (N_5223,N_4851,N_4321);
nand U5224 (N_5224,N_4973,N_4604);
or U5225 (N_5225,N_2739,N_4743);
or U5226 (N_5226,N_2863,N_4451);
xor U5227 (N_5227,N_4440,N_4729);
or U5228 (N_5228,N_2673,N_3021);
and U5229 (N_5229,N_4638,N_3161);
and U5230 (N_5230,N_3526,N_4473);
or U5231 (N_5231,N_4366,N_3359);
or U5232 (N_5232,N_3140,N_3260);
nand U5233 (N_5233,N_3605,N_3612);
nor U5234 (N_5234,N_4352,N_3890);
or U5235 (N_5235,N_3686,N_4424);
and U5236 (N_5236,N_3414,N_3070);
nor U5237 (N_5237,N_3525,N_2832);
nor U5238 (N_5238,N_2828,N_3490);
and U5239 (N_5239,N_3705,N_3943);
or U5240 (N_5240,N_3742,N_4947);
xnor U5241 (N_5241,N_3785,N_3617);
or U5242 (N_5242,N_3380,N_4766);
and U5243 (N_5243,N_4626,N_3265);
and U5244 (N_5244,N_4067,N_2604);
nand U5245 (N_5245,N_4860,N_4962);
and U5246 (N_5246,N_4317,N_3137);
or U5247 (N_5247,N_2932,N_3492);
nor U5248 (N_5248,N_3741,N_3576);
or U5249 (N_5249,N_3218,N_3512);
nor U5250 (N_5250,N_4337,N_3200);
and U5251 (N_5251,N_3002,N_3147);
and U5252 (N_5252,N_4155,N_2777);
and U5253 (N_5253,N_3603,N_3461);
and U5254 (N_5254,N_3674,N_4194);
or U5255 (N_5255,N_2823,N_4048);
nand U5256 (N_5256,N_3199,N_2523);
nor U5257 (N_5257,N_2546,N_3997);
and U5258 (N_5258,N_3292,N_2824);
nand U5259 (N_5259,N_3818,N_3815);
nand U5260 (N_5260,N_4340,N_3044);
and U5261 (N_5261,N_2539,N_2578);
nor U5262 (N_5262,N_3644,N_4798);
or U5263 (N_5263,N_3212,N_2818);
or U5264 (N_5264,N_3160,N_3828);
or U5265 (N_5265,N_4699,N_3071);
xnor U5266 (N_5266,N_3248,N_4859);
or U5267 (N_5267,N_4216,N_3078);
or U5268 (N_5268,N_3211,N_2857);
or U5269 (N_5269,N_3189,N_4656);
nand U5270 (N_5270,N_3682,N_4924);
nor U5271 (N_5271,N_3967,N_2557);
nor U5272 (N_5272,N_2922,N_3033);
nor U5273 (N_5273,N_2910,N_4664);
nor U5274 (N_5274,N_4107,N_4180);
nand U5275 (N_5275,N_4096,N_2784);
xnor U5276 (N_5276,N_2826,N_4082);
and U5277 (N_5277,N_3894,N_3275);
and U5278 (N_5278,N_4684,N_4690);
or U5279 (N_5279,N_3416,N_3871);
and U5280 (N_5280,N_4960,N_3420);
nor U5281 (N_5281,N_2815,N_4657);
and U5282 (N_5282,N_3966,N_4257);
nand U5283 (N_5283,N_3892,N_3968);
nand U5284 (N_5284,N_3111,N_3971);
nor U5285 (N_5285,N_4265,N_3709);
nor U5286 (N_5286,N_4687,N_4565);
nor U5287 (N_5287,N_4212,N_4115);
or U5288 (N_5288,N_2919,N_3419);
or U5289 (N_5289,N_4985,N_3872);
nor U5290 (N_5290,N_3537,N_4827);
nor U5291 (N_5291,N_3483,N_3122);
xor U5292 (N_5292,N_3331,N_3812);
xnor U5293 (N_5293,N_2749,N_3726);
nor U5294 (N_5294,N_3870,N_3927);
and U5295 (N_5295,N_3438,N_2808);
and U5296 (N_5296,N_4453,N_3382);
or U5297 (N_5297,N_3264,N_3481);
and U5298 (N_5298,N_4201,N_2603);
nand U5299 (N_5299,N_4467,N_4280);
nand U5300 (N_5300,N_3840,N_4826);
nor U5301 (N_5301,N_3009,N_3816);
nor U5302 (N_5302,N_2629,N_3797);
and U5303 (N_5303,N_3659,N_4945);
and U5304 (N_5304,N_3110,N_2664);
and U5305 (N_5305,N_4793,N_4739);
nand U5306 (N_5306,N_4853,N_4598);
nand U5307 (N_5307,N_3245,N_2540);
nor U5308 (N_5308,N_4149,N_3364);
and U5309 (N_5309,N_3995,N_3038);
nor U5310 (N_5310,N_3782,N_3204);
or U5311 (N_5311,N_2819,N_4272);
nand U5312 (N_5312,N_2750,N_4156);
xnor U5313 (N_5313,N_4639,N_4824);
nor U5314 (N_5314,N_4596,N_3752);
or U5315 (N_5315,N_3937,N_2694);
nor U5316 (N_5316,N_4327,N_2951);
xnor U5317 (N_5317,N_4974,N_4334);
or U5318 (N_5318,N_3423,N_4085);
xor U5319 (N_5319,N_4895,N_4449);
and U5320 (N_5320,N_4229,N_3637);
or U5321 (N_5321,N_2848,N_3433);
and U5322 (N_5322,N_3706,N_4421);
nor U5323 (N_5323,N_2697,N_3737);
nand U5324 (N_5324,N_4631,N_2914);
nor U5325 (N_5325,N_3805,N_2927);
and U5326 (N_5326,N_2648,N_3787);
or U5327 (N_5327,N_3440,N_4892);
xnor U5328 (N_5328,N_4073,N_4745);
xnor U5329 (N_5329,N_4736,N_3858);
or U5330 (N_5330,N_2532,N_3475);
or U5331 (N_5331,N_3541,N_3169);
nand U5332 (N_5332,N_3680,N_2670);
nor U5333 (N_5333,N_3387,N_2967);
xnor U5334 (N_5334,N_3102,N_3079);
and U5335 (N_5335,N_3332,N_2892);
nor U5336 (N_5336,N_3567,N_3234);
nor U5337 (N_5337,N_4649,N_2983);
and U5338 (N_5338,N_3157,N_3530);
and U5339 (N_5339,N_3773,N_3354);
or U5340 (N_5340,N_3468,N_3675);
nand U5341 (N_5341,N_3961,N_3143);
nor U5342 (N_5342,N_4014,N_4181);
or U5343 (N_5343,N_3697,N_3750);
or U5344 (N_5344,N_3361,N_4746);
and U5345 (N_5345,N_3621,N_2811);
nand U5346 (N_5346,N_4535,N_4601);
nand U5347 (N_5347,N_3080,N_3172);
or U5348 (N_5348,N_3546,N_3150);
nand U5349 (N_5349,N_4843,N_4643);
and U5350 (N_5350,N_4808,N_2947);
nor U5351 (N_5351,N_3467,N_2657);
and U5352 (N_5352,N_3573,N_4144);
nand U5353 (N_5353,N_2589,N_4384);
or U5354 (N_5354,N_4965,N_3443);
or U5355 (N_5355,N_3960,N_3298);
nand U5356 (N_5356,N_2846,N_4994);
nor U5357 (N_5357,N_3488,N_3650);
nor U5358 (N_5358,N_3854,N_3619);
or U5359 (N_5359,N_4237,N_3321);
nand U5360 (N_5360,N_2537,N_4066);
nor U5361 (N_5361,N_2993,N_3986);
and U5362 (N_5362,N_2615,N_3542);
nor U5363 (N_5363,N_3087,N_4469);
or U5364 (N_5364,N_4130,N_4439);
and U5365 (N_5365,N_4080,N_2690);
nand U5366 (N_5366,N_4083,N_4143);
xnor U5367 (N_5367,N_2903,N_3486);
nand U5368 (N_5368,N_2668,N_4963);
and U5369 (N_5369,N_3869,N_3424);
or U5370 (N_5370,N_3388,N_3781);
and U5371 (N_5371,N_2634,N_3722);
and U5372 (N_5372,N_4801,N_4573);
nor U5373 (N_5373,N_3261,N_2541);
nor U5374 (N_5374,N_4360,N_2986);
nor U5375 (N_5375,N_3519,N_3149);
or U5376 (N_5376,N_4609,N_4589);
or U5377 (N_5377,N_2996,N_4268);
and U5378 (N_5378,N_3793,N_4556);
nor U5379 (N_5379,N_4800,N_3656);
xnor U5380 (N_5380,N_4658,N_4946);
nand U5381 (N_5381,N_3130,N_2510);
and U5382 (N_5382,N_3744,N_3310);
nand U5383 (N_5383,N_3877,N_3556);
or U5384 (N_5384,N_2734,N_2838);
nor U5385 (N_5385,N_3746,N_3196);
nor U5386 (N_5386,N_4549,N_3963);
or U5387 (N_5387,N_3664,N_3445);
nor U5388 (N_5388,N_4576,N_4693);
or U5389 (N_5389,N_4190,N_2677);
or U5390 (N_5390,N_2728,N_4575);
and U5391 (N_5391,N_4177,N_2731);
or U5392 (N_5392,N_2567,N_4996);
nor U5393 (N_5393,N_4984,N_2806);
and U5394 (N_5394,N_3957,N_4355);
and U5395 (N_5395,N_3208,N_3861);
nor U5396 (N_5396,N_3401,N_3482);
nor U5397 (N_5397,N_4357,N_2575);
or U5398 (N_5398,N_4395,N_2715);
nand U5399 (N_5399,N_4674,N_4901);
nand U5400 (N_5400,N_3457,N_2616);
or U5401 (N_5401,N_3578,N_4486);
nand U5402 (N_5402,N_4329,N_2949);
xor U5403 (N_5403,N_4894,N_3606);
nand U5404 (N_5404,N_4863,N_2735);
xnor U5405 (N_5405,N_4479,N_4647);
xor U5406 (N_5406,N_3778,N_4283);
or U5407 (N_5407,N_3777,N_4594);
nand U5408 (N_5408,N_2702,N_4445);
nor U5409 (N_5409,N_3655,N_4519);
nor U5410 (N_5410,N_2991,N_4169);
and U5411 (N_5411,N_2726,N_3383);
nor U5412 (N_5412,N_4661,N_2570);
and U5413 (N_5413,N_3118,N_3814);
nor U5414 (N_5414,N_3415,N_3929);
nand U5415 (N_5415,N_3590,N_4404);
or U5416 (N_5416,N_3884,N_4780);
nor U5417 (N_5417,N_4197,N_2636);
and U5418 (N_5418,N_4009,N_4992);
nor U5419 (N_5419,N_4209,N_2571);
nor U5420 (N_5420,N_4660,N_4982);
xor U5421 (N_5421,N_3795,N_3119);
nand U5422 (N_5422,N_4324,N_2876);
nor U5423 (N_5423,N_3225,N_2717);
and U5424 (N_5424,N_2654,N_4282);
nor U5425 (N_5425,N_2789,N_2556);
or U5426 (N_5426,N_3316,N_4228);
and U5427 (N_5427,N_2609,N_4630);
nor U5428 (N_5428,N_2771,N_2507);
and U5429 (N_5429,N_4734,N_4916);
nand U5430 (N_5430,N_2646,N_4059);
nor U5431 (N_5431,N_4291,N_4957);
or U5432 (N_5432,N_2687,N_2588);
xor U5433 (N_5433,N_2652,N_2549);
xnor U5434 (N_5434,N_3233,N_4818);
nor U5435 (N_5435,N_4832,N_2831);
or U5436 (N_5436,N_3284,N_3141);
xor U5437 (N_5437,N_3393,N_2973);
or U5438 (N_5438,N_2692,N_3701);
or U5439 (N_5439,N_4551,N_4058);
or U5440 (N_5440,N_4456,N_4688);
nor U5441 (N_5441,N_4663,N_4278);
nand U5442 (N_5442,N_4532,N_4390);
or U5443 (N_5443,N_3720,N_2865);
nor U5444 (N_5444,N_4060,N_3915);
nand U5445 (N_5445,N_4558,N_4425);
and U5446 (N_5446,N_3776,N_4290);
nand U5447 (N_5447,N_4704,N_4579);
and U5448 (N_5448,N_2710,N_4047);
nand U5449 (N_5449,N_2626,N_4666);
or U5450 (N_5450,N_3152,N_3400);
nor U5451 (N_5451,N_3669,N_4253);
nand U5452 (N_5452,N_3327,N_3791);
nor U5453 (N_5453,N_4659,N_3555);
nor U5454 (N_5454,N_2660,N_4933);
nand U5455 (N_5455,N_3136,N_3765);
or U5456 (N_5456,N_3129,N_4939);
nand U5457 (N_5457,N_4719,N_3936);
and U5458 (N_5458,N_4223,N_2602);
nor U5459 (N_5459,N_4932,N_3340);
xor U5460 (N_5460,N_4037,N_4422);
nand U5461 (N_5461,N_3456,N_4665);
or U5462 (N_5462,N_3135,N_3198);
xnor U5463 (N_5463,N_4720,N_2963);
nor U5464 (N_5464,N_4857,N_3365);
or U5465 (N_5465,N_3973,N_4427);
nand U5466 (N_5466,N_3273,N_3739);
nor U5467 (N_5467,N_4995,N_4577);
nand U5468 (N_5468,N_2565,N_3025);
and U5469 (N_5469,N_3297,N_3962);
xor U5470 (N_5470,N_2525,N_3725);
and U5471 (N_5471,N_4319,N_4419);
and U5472 (N_5472,N_4560,N_3511);
nor U5473 (N_5473,N_3367,N_3721);
nor U5474 (N_5474,N_3319,N_4854);
and U5475 (N_5475,N_4313,N_4935);
or U5476 (N_5476,N_3801,N_2741);
xor U5477 (N_5477,N_4091,N_4953);
or U5478 (N_5478,N_4764,N_4513);
nor U5479 (N_5479,N_3077,N_2725);
nand U5480 (N_5480,N_2764,N_4998);
and U5481 (N_5481,N_4031,N_3751);
nand U5482 (N_5482,N_4839,N_4196);
and U5483 (N_5483,N_4187,N_4510);
nor U5484 (N_5484,N_4816,N_4458);
nand U5485 (N_5485,N_3595,N_4377);
nor U5486 (N_5486,N_4813,N_4426);
and U5487 (N_5487,N_2748,N_4448);
or U5488 (N_5488,N_3213,N_2605);
and U5489 (N_5489,N_2522,N_2562);
xnor U5490 (N_5490,N_3572,N_3838);
and U5491 (N_5491,N_4872,N_4118);
nor U5492 (N_5492,N_4396,N_3487);
nor U5493 (N_5493,N_4333,N_4986);
and U5494 (N_5494,N_3272,N_3373);
nor U5495 (N_5495,N_3372,N_3984);
or U5496 (N_5496,N_3108,N_4008);
nor U5497 (N_5497,N_3789,N_3277);
nand U5498 (N_5498,N_4251,N_4230);
or U5499 (N_5499,N_3653,N_3677);
nand U5500 (N_5500,N_3935,N_2617);
or U5501 (N_5501,N_3197,N_2530);
or U5502 (N_5502,N_3252,N_4679);
nor U5503 (N_5503,N_4015,N_3632);
or U5504 (N_5504,N_4821,N_4269);
nand U5505 (N_5505,N_4068,N_4683);
xnor U5506 (N_5506,N_4611,N_3719);
nor U5507 (N_5507,N_3714,N_4629);
nand U5508 (N_5508,N_4266,N_3625);
nor U5509 (N_5509,N_3114,N_3432);
or U5510 (N_5510,N_3657,N_4751);
nand U5511 (N_5511,N_4478,N_3258);
nor U5512 (N_5512,N_4470,N_3518);
xor U5513 (N_5513,N_4023,N_4781);
or U5514 (N_5514,N_4891,N_4805);
or U5515 (N_5515,N_2946,N_3704);
nand U5516 (N_5516,N_3464,N_4538);
nand U5517 (N_5517,N_4868,N_4948);
or U5518 (N_5518,N_3507,N_3700);
nand U5519 (N_5519,N_3859,N_4902);
nand U5520 (N_5520,N_3022,N_3001);
or U5521 (N_5521,N_3850,N_4285);
nor U5522 (N_5522,N_3476,N_3192);
and U5523 (N_5523,N_2542,N_4186);
nor U5524 (N_5524,N_4918,N_3254);
nor U5525 (N_5525,N_2803,N_4005);
and U5526 (N_5526,N_4624,N_4920);
nor U5527 (N_5527,N_2655,N_3203);
nor U5528 (N_5528,N_4737,N_4389);
nor U5529 (N_5529,N_4523,N_3724);
nor U5530 (N_5530,N_4543,N_3853);
xor U5531 (N_5531,N_4711,N_3153);
or U5532 (N_5532,N_2796,N_3030);
nand U5533 (N_5533,N_3830,N_2759);
nand U5534 (N_5534,N_3626,N_3992);
nor U5535 (N_5535,N_3267,N_2577);
nor U5536 (N_5536,N_3786,N_4539);
xnor U5537 (N_5537,N_2948,N_3707);
nand U5538 (N_5538,N_4323,N_4135);
nand U5539 (N_5539,N_4325,N_3164);
nor U5540 (N_5540,N_2593,N_3113);
or U5541 (N_5541,N_4179,N_4921);
nor U5542 (N_5542,N_4367,N_4914);
xnor U5543 (N_5543,N_2529,N_3371);
or U5544 (N_5544,N_4913,N_3635);
and U5545 (N_5545,N_4597,N_3821);
and U5546 (N_5546,N_4713,N_4820);
nor U5547 (N_5547,N_4696,N_3047);
or U5548 (N_5548,N_2827,N_3409);
nor U5549 (N_5549,N_2782,N_3502);
xor U5550 (N_5550,N_3568,N_4077);
or U5551 (N_5551,N_3783,N_3522);
and U5552 (N_5552,N_3352,N_4199);
nor U5553 (N_5553,N_4929,N_4284);
or U5554 (N_5554,N_4928,N_3145);
or U5555 (N_5555,N_4605,N_3031);
and U5556 (N_5556,N_2744,N_3647);
nor U5557 (N_5557,N_4896,N_4488);
nand U5558 (N_5558,N_3134,N_4418);
nor U5559 (N_5559,N_4727,N_4776);
and U5560 (N_5560,N_3042,N_3591);
xnor U5561 (N_5561,N_4248,N_4785);
nand U5562 (N_5562,N_4931,N_3202);
and U5563 (N_5563,N_3736,N_3454);
nand U5564 (N_5564,N_4087,N_3665);
xor U5565 (N_5565,N_3049,N_4942);
nor U5566 (N_5566,N_3779,N_4707);
and U5567 (N_5567,N_4244,N_4584);
and U5568 (N_5568,N_2620,N_3085);
or U5569 (N_5569,N_4202,N_4757);
xnor U5570 (N_5570,N_3294,N_4969);
xor U5571 (N_5571,N_3583,N_3473);
and U5572 (N_5572,N_3426,N_4748);
or U5573 (N_5573,N_2791,N_3104);
nor U5574 (N_5574,N_3585,N_4838);
nor U5575 (N_5575,N_4772,N_4259);
nand U5576 (N_5576,N_3880,N_2871);
or U5577 (N_5577,N_4231,N_4182);
xnor U5578 (N_5578,N_4344,N_3923);
xnor U5579 (N_5579,N_2971,N_3592);
nand U5580 (N_5580,N_2639,N_3813);
and U5581 (N_5581,N_4123,N_3955);
and U5582 (N_5582,N_3965,N_4312);
nor U5583 (N_5583,N_3063,N_3913);
and U5584 (N_5584,N_2509,N_2774);
nand U5585 (N_5585,N_4184,N_3698);
nand U5586 (N_5586,N_2805,N_3754);
or U5587 (N_5587,N_3061,N_3345);
or U5588 (N_5588,N_4279,N_3163);
nand U5589 (N_5589,N_3796,N_4586);
or U5590 (N_5590,N_4829,N_3112);
and U5591 (N_5591,N_3337,N_4303);
and U5592 (N_5592,N_2860,N_3217);
nor U5593 (N_5593,N_2566,N_3058);
nor U5594 (N_5594,N_2767,N_2989);
or U5595 (N_5595,N_4802,N_4428);
nor U5596 (N_5596,N_3931,N_4930);
nor U5597 (N_5597,N_3188,N_4356);
nor U5598 (N_5598,N_4026,N_4883);
and U5599 (N_5599,N_4241,N_3399);
nand U5600 (N_5600,N_2995,N_2888);
and U5601 (N_5601,N_2706,N_4410);
nand U5602 (N_5602,N_3428,N_2656);
or U5603 (N_5603,N_3274,N_3095);
and U5604 (N_5604,N_4238,N_3803);
nand U5605 (N_5605,N_3449,N_4342);
or U5606 (N_5606,N_3749,N_4790);
or U5607 (N_5607,N_4915,N_3054);
and U5608 (N_5608,N_3138,N_4964);
or U5609 (N_5609,N_3126,N_3043);
xor U5610 (N_5610,N_3396,N_2928);
and U5611 (N_5611,N_4379,N_3847);
nand U5612 (N_5612,N_4443,N_3024);
and U5613 (N_5613,N_3758,N_4750);
nand U5614 (N_5614,N_4858,N_3627);
or U5615 (N_5615,N_2513,N_4141);
nand U5616 (N_5616,N_3183,N_4566);
nor U5617 (N_5617,N_2778,N_3703);
nor U5618 (N_5618,N_2607,N_3389);
or U5619 (N_5619,N_3543,N_2614);
or U5620 (N_5620,N_4940,N_3253);
nor U5621 (N_5621,N_3441,N_3903);
xor U5622 (N_5622,N_3057,N_3165);
and U5623 (N_5623,N_4689,N_4862);
or U5624 (N_5624,N_3148,N_3551);
nand U5625 (N_5625,N_4249,N_4599);
nor U5626 (N_5626,N_4374,N_4348);
nor U5627 (N_5627,N_2902,N_3788);
and U5628 (N_5628,N_4286,N_2862);
nor U5629 (N_5629,N_3671,N_3681);
nand U5630 (N_5630,N_2855,N_4952);
nor U5631 (N_5631,N_3646,N_3422);
nand U5632 (N_5632,N_4849,N_4540);
nand U5633 (N_5633,N_3683,N_4124);
and U5634 (N_5634,N_4900,N_3560);
and U5635 (N_5635,N_4120,N_4670);
or U5636 (N_5636,N_3827,N_4022);
or U5637 (N_5637,N_4438,N_2962);
nor U5638 (N_5638,N_2800,N_4703);
or U5639 (N_5639,N_3139,N_3478);
and U5640 (N_5640,N_2681,N_2696);
or U5641 (N_5641,N_3663,N_3210);
nor U5642 (N_5642,N_2816,N_4545);
xnor U5643 (N_5643,N_3771,N_3385);
or U5644 (N_5644,N_4518,N_3942);
nor U5645 (N_5645,N_2859,N_2601);
nand U5646 (N_5646,N_3571,N_2904);
nor U5647 (N_5647,N_4255,N_3531);
nor U5648 (N_5648,N_2911,N_2945);
nor U5649 (N_5649,N_4351,N_4667);
nor U5650 (N_5650,N_2727,N_3881);
and U5651 (N_5651,N_2858,N_3908);
and U5652 (N_5652,N_3959,N_2810);
and U5653 (N_5653,N_4732,N_4386);
and U5654 (N_5654,N_2740,N_3845);
and U5655 (N_5655,N_4121,N_4815);
and U5656 (N_5656,N_4814,N_4975);
and U5657 (N_5657,N_3216,N_3549);
xnor U5658 (N_5658,N_4092,N_3103);
and U5659 (N_5659,N_4569,N_2524);
nand U5660 (N_5660,N_2533,N_4922);
and U5661 (N_5661,N_2758,N_3598);
or U5662 (N_5662,N_2527,N_4840);
nand U5663 (N_5663,N_3346,N_3846);
nand U5664 (N_5664,N_4682,N_3552);
nor U5665 (N_5665,N_3013,N_3125);
and U5666 (N_5666,N_3717,N_3447);
or U5667 (N_5667,N_3489,N_3330);
nand U5668 (N_5668,N_4722,N_3286);
or U5669 (N_5669,N_3320,N_2606);
or U5670 (N_5670,N_4897,N_4799);
or U5671 (N_5671,N_4261,N_3611);
nor U5672 (N_5672,N_4046,N_2583);
and U5673 (N_5673,N_2891,N_2929);
nand U5674 (N_5674,N_4723,N_2792);
or U5675 (N_5675,N_2936,N_4306);
and U5676 (N_5676,N_4708,N_3833);
and U5677 (N_5677,N_4041,N_4526);
and U5678 (N_5678,N_2970,N_4454);
nand U5679 (N_5679,N_4382,N_2844);
nor U5680 (N_5680,N_2886,N_4311);
nor U5681 (N_5681,N_4018,N_4967);
and U5682 (N_5682,N_4715,N_4380);
and U5683 (N_5683,N_4027,N_4142);
nand U5684 (N_5684,N_4254,N_3780);
and U5685 (N_5685,N_3485,N_2686);
nor U5686 (N_5686,N_2579,N_3538);
nor U5687 (N_5687,N_3325,N_2776);
and U5688 (N_5688,N_3760,N_4553);
xor U5689 (N_5689,N_3564,N_3889);
or U5690 (N_5690,N_4758,N_4495);
nand U5691 (N_5691,N_3174,N_4170);
or U5692 (N_5692,N_3266,N_4784);
nand U5693 (N_5693,N_3645,N_4061);
and U5694 (N_5694,N_3949,N_3864);
nor U5695 (N_5695,N_4796,N_2834);
nor U5696 (N_5696,N_4466,N_4205);
or U5697 (N_5697,N_2516,N_4341);
nand U5698 (N_5698,N_3338,N_2909);
nor U5699 (N_5699,N_3731,N_4154);
nor U5700 (N_5700,N_3735,N_2917);
nand U5701 (N_5701,N_2999,N_3249);
or U5702 (N_5702,N_2534,N_4521);
or U5703 (N_5703,N_3658,N_4841);
and U5704 (N_5704,N_2807,N_3976);
nand U5705 (N_5705,N_2732,N_3406);
nand U5706 (N_5706,N_2612,N_4618);
nand U5707 (N_5707,N_3769,N_4373);
and U5708 (N_5708,N_2842,N_3173);
nand U5709 (N_5709,N_3392,N_4474);
nand U5710 (N_5710,N_3631,N_4045);
or U5711 (N_5711,N_4444,N_3301);
nand U5712 (N_5712,N_3289,N_3014);
and U5713 (N_5713,N_4106,N_3451);
xnor U5714 (N_5714,N_3403,N_4677);
nand U5715 (N_5715,N_3232,N_4717);
and U5716 (N_5716,N_3191,N_4203);
nand U5717 (N_5717,N_4260,N_2881);
nand U5718 (N_5718,N_2972,N_3067);
nand U5719 (N_5719,N_3865,N_4879);
nand U5720 (N_5720,N_3168,N_4276);
nor U5721 (N_5721,N_3405,N_4064);
nand U5722 (N_5722,N_4247,N_3553);
or U5723 (N_5723,N_3584,N_2849);
and U5724 (N_5724,N_4297,N_4795);
and U5725 (N_5725,N_4416,N_3171);
nand U5726 (N_5726,N_4955,N_3131);
nor U5727 (N_5727,N_3798,N_4700);
xor U5728 (N_5728,N_3259,N_3427);
nand U5729 (N_5729,N_4270,N_2788);
or U5730 (N_5730,N_4692,N_2850);
or U5731 (N_5731,N_4775,N_3357);
or U5732 (N_5732,N_3227,N_3397);
nand U5733 (N_5733,N_4685,N_4590);
or U5734 (N_5734,N_3711,N_2737);
and U5735 (N_5735,N_4958,N_4765);
nand U5736 (N_5736,N_3998,N_2581);
nand U5737 (N_5737,N_3610,N_4546);
nand U5738 (N_5738,N_4791,N_4873);
or U5739 (N_5739,N_4941,N_4492);
or U5740 (N_5740,N_3906,N_3991);
nor U5741 (N_5741,N_3329,N_3589);
nand U5742 (N_5742,N_4414,N_3728);
or U5743 (N_5743,N_3860,N_3608);
and U5744 (N_5744,N_4090,N_4544);
xor U5745 (N_5745,N_4407,N_3235);
or U5746 (N_5746,N_3579,N_3293);
or U5747 (N_5747,N_2889,N_2861);
nor U5748 (N_5748,N_3581,N_4888);
nand U5749 (N_5749,N_3381,N_4294);
or U5750 (N_5750,N_4489,N_4625);
or U5751 (N_5751,N_2976,N_4735);
and U5752 (N_5752,N_3144,N_3082);
or U5753 (N_5753,N_3862,N_3587);
and U5754 (N_5754,N_3832,N_4125);
nand U5755 (N_5755,N_3186,N_3039);
nor U5756 (N_5756,N_4452,N_2987);
or U5757 (N_5757,N_3028,N_4385);
or U5758 (N_5758,N_2703,N_3279);
nand U5759 (N_5759,N_4267,N_3917);
nor U5760 (N_5760,N_2912,N_3369);
nor U5761 (N_5761,N_4507,N_4042);
nor U5762 (N_5762,N_3347,N_4112);
or U5763 (N_5763,N_3684,N_4976);
or U5764 (N_5764,N_4595,N_3747);
and U5765 (N_5765,N_3120,N_4614);
nor U5766 (N_5766,N_4111,N_4296);
or U5767 (N_5767,N_3508,N_4108);
xor U5768 (N_5768,N_2611,N_3879);
or U5769 (N_5769,N_3472,N_2679);
and U5770 (N_5770,N_2528,N_4273);
or U5771 (N_5771,N_3888,N_3696);
or U5772 (N_5772,N_3899,N_3107);
nand U5773 (N_5773,N_3910,N_3874);
or U5774 (N_5774,N_4339,N_3312);
and U5775 (N_5775,N_3378,N_4615);
and U5776 (N_5776,N_3180,N_2743);
nor U5777 (N_5777,N_4293,N_4100);
or U5778 (N_5778,N_3341,N_3604);
and U5779 (N_5779,N_2954,N_3996);
and U5780 (N_5780,N_2773,N_4475);
or U5781 (N_5781,N_4331,N_4105);
nand U5782 (N_5782,N_2651,N_3580);
nand U5783 (N_5783,N_4383,N_2721);
nand U5784 (N_5784,N_4650,N_3195);
nor U5785 (N_5785,N_3593,N_4161);
and U5786 (N_5786,N_4274,N_3866);
or U5787 (N_5787,N_4215,N_3007);
or U5788 (N_5788,N_2890,N_3460);
or U5789 (N_5789,N_2798,N_4074);
and U5790 (N_5790,N_2896,N_4970);
and U5791 (N_5791,N_4062,N_4880);
and U5792 (N_5792,N_4242,N_3479);
nor U5793 (N_5793,N_3162,N_4171);
xnor U5794 (N_5794,N_4287,N_4213);
or U5795 (N_5795,N_4178,N_3469);
nor U5796 (N_5796,N_2872,N_3623);
xnor U5797 (N_5797,N_4232,N_4075);
nand U5798 (N_5798,N_2555,N_2907);
nor U5799 (N_5799,N_4004,N_4436);
nand U5800 (N_5800,N_3105,N_4032);
and U5801 (N_5801,N_3520,N_2845);
or U5802 (N_5802,N_3015,N_4944);
nor U5803 (N_5803,N_4481,N_4978);
nor U5804 (N_5804,N_3343,N_2781);
or U5805 (N_5805,N_4078,N_4912);
nand U5806 (N_5806,N_3614,N_3123);
or U5807 (N_5807,N_2720,N_4258);
or U5808 (N_5808,N_3835,N_4185);
nand U5809 (N_5809,N_3687,N_2982);
nand U5810 (N_5810,N_4520,N_4086);
nand U5811 (N_5811,N_3535,N_4989);
xnor U5812 (N_5812,N_3844,N_4468);
nand U5813 (N_5813,N_4491,N_4623);
or U5814 (N_5814,N_3055,N_3755);
nand U5815 (N_5815,N_4644,N_3934);
xnor U5816 (N_5816,N_3911,N_2563);
nor U5817 (N_5817,N_2895,N_3740);
nor U5818 (N_5818,N_2813,N_4714);
and U5819 (N_5819,N_3300,N_4547);
or U5820 (N_5820,N_4016,N_4307);
xor U5821 (N_5821,N_3206,N_2957);
or U5822 (N_5822,N_4406,N_4593);
and U5823 (N_5823,N_4504,N_3924);
or U5824 (N_5824,N_4768,N_3281);
nor U5825 (N_5825,N_3376,N_4512);
and U5826 (N_5826,N_2500,N_4557);
nand U5827 (N_5827,N_3240,N_4522);
nor U5828 (N_5828,N_4403,N_3775);
xor U5829 (N_5829,N_4855,N_3514);
or U5830 (N_5830,N_4844,N_3734);
nor U5831 (N_5831,N_4233,N_3829);
and U5832 (N_5832,N_4981,N_4697);
nand U5833 (N_5833,N_3944,N_4542);
or U5834 (N_5834,N_3638,N_3506);
and U5835 (N_5835,N_3940,N_3177);
or U5836 (N_5836,N_2980,N_4636);
xor U5837 (N_5837,N_4886,N_3718);
nor U5838 (N_5838,N_2649,N_4138);
nand U5839 (N_5839,N_3895,N_2756);
or U5840 (N_5840,N_3166,N_3314);
nor U5841 (N_5841,N_4804,N_2707);
nand U5842 (N_5842,N_3184,N_4336);
nand U5843 (N_5843,N_3634,N_3733);
and U5844 (N_5844,N_4420,N_2547);
or U5845 (N_5845,N_3088,N_2966);
nand U5846 (N_5846,N_4174,N_3964);
and U5847 (N_5847,N_2921,N_3439);
or U5848 (N_5848,N_2905,N_2691);
xor U5849 (N_5849,N_4103,N_3296);
nand U5850 (N_5850,N_2935,N_3661);
and U5851 (N_5851,N_3501,N_2820);
and U5852 (N_5852,N_4359,N_3867);
nand U5853 (N_5853,N_4057,N_4305);
nand U5854 (N_5854,N_3465,N_4220);
and U5855 (N_5855,N_4606,N_3307);
nand U5856 (N_5856,N_3974,N_2836);
xnor U5857 (N_5857,N_3642,N_4158);
or U5858 (N_5858,N_4585,N_4917);
nand U5859 (N_5859,N_3676,N_4789);
or U5860 (N_5860,N_3404,N_3315);
nor U5861 (N_5861,N_3550,N_4227);
nor U5862 (N_5862,N_2531,N_3834);
or U5863 (N_5863,N_4968,N_4848);
and U5864 (N_5864,N_4919,N_4807);
nand U5865 (N_5865,N_4221,N_3124);
nand U5866 (N_5866,N_4246,N_3672);
nor U5867 (N_5867,N_3246,N_2853);
nand U5868 (N_5868,N_4021,N_2590);
xor U5869 (N_5869,N_2965,N_2780);
nand U5870 (N_5870,N_4104,N_4803);
nand U5871 (N_5871,N_3639,N_3770);
or U5872 (N_5872,N_2754,N_2610);
nor U5873 (N_5873,N_3004,N_3480);
nor U5874 (N_5874,N_2705,N_3673);
nand U5875 (N_5875,N_3629,N_4943);
nand U5876 (N_5876,N_4607,N_4069);
xor U5877 (N_5877,N_2559,N_4300);
nor U5878 (N_5878,N_3231,N_3548);
or U5879 (N_5879,N_3499,N_3855);
nor U5880 (N_5880,N_2874,N_4890);
nor U5881 (N_5881,N_4219,N_4012);
nand U5882 (N_5882,N_4610,N_2804);
nor U5883 (N_5883,N_3256,N_4224);
and U5884 (N_5884,N_3000,N_2597);
xnor U5885 (N_5885,N_3379,N_4669);
nand U5886 (N_5886,N_2653,N_3121);
nor U5887 (N_5887,N_4136,N_4054);
nor U5888 (N_5888,N_2518,N_3062);
and U5889 (N_5889,N_4695,N_3628);
nor U5890 (N_5890,N_3251,N_2768);
and U5891 (N_5891,N_3442,N_3768);
nor U5892 (N_5892,N_4338,N_3417);
and U5893 (N_5893,N_3784,N_4725);
and U5894 (N_5894,N_4281,N_3370);
or U5895 (N_5895,N_3532,N_4825);
or U5896 (N_5896,N_3918,N_4434);
nor U5897 (N_5897,N_4655,N_3852);
nor U5898 (N_5898,N_4712,N_3425);
nand U5899 (N_5899,N_3117,N_4200);
nand U5900 (N_5900,N_3806,N_4132);
nand U5901 (N_5901,N_4101,N_2900);
nor U5902 (N_5902,N_4773,N_4376);
nor U5903 (N_5903,N_2685,N_2829);
nor U5904 (N_5904,N_4552,N_3221);
and U5905 (N_5905,N_3539,N_3678);
nor U5906 (N_5906,N_2943,N_2978);
and U5907 (N_5907,N_3133,N_3922);
and U5908 (N_5908,N_2884,N_3527);
and U5909 (N_5909,N_3685,N_3223);
nand U5910 (N_5910,N_4044,N_4812);
xnor U5911 (N_5911,N_3577,N_3873);
nor U5912 (N_5912,N_2990,N_3882);
nor U5913 (N_5913,N_4997,N_2837);
and U5914 (N_5914,N_3342,N_2561);
and U5915 (N_5915,N_2799,N_2698);
nor U5916 (N_5916,N_3081,N_4641);
nand U5917 (N_5917,N_3099,N_2809);
nand U5918 (N_5918,N_3083,N_3601);
nand U5919 (N_5919,N_2753,N_3932);
xnor U5920 (N_5920,N_3154,N_3010);
and U5921 (N_5921,N_3756,N_4904);
nand U5922 (N_5922,N_4218,N_2695);
xnor U5923 (N_5923,N_2678,N_4811);
xor U5924 (N_5924,N_2938,N_4646);
nor U5925 (N_5925,N_4668,N_3774);
or U5926 (N_5926,N_3363,N_4191);
nand U5927 (N_5927,N_3633,N_3652);
nor U5928 (N_5928,N_4328,N_3178);
xor U5929 (N_5929,N_3045,N_2763);
nand U5930 (N_5930,N_2794,N_3471);
and U5931 (N_5931,N_4534,N_2543);
or U5932 (N_5932,N_3390,N_2833);
or U5933 (N_5933,N_4654,N_4903);
and U5934 (N_5934,N_3876,N_4195);
xor U5935 (N_5935,N_4217,N_4907);
nand U5936 (N_5936,N_3989,N_4988);
nor U5937 (N_5937,N_3999,N_4001);
and U5938 (N_5938,N_2627,N_3029);
and U5939 (N_5939,N_3358,N_4645);
or U5940 (N_5940,N_2501,N_3431);
xnor U5941 (N_5941,N_2504,N_2761);
xor U5942 (N_5942,N_2508,N_3109);
nand U5943 (N_5943,N_4036,N_3575);
nor U5944 (N_5944,N_4680,N_2887);
nand U5945 (N_5945,N_3356,N_4705);
xnor U5946 (N_5946,N_3710,N_4211);
nor U5947 (N_5947,N_4509,N_3496);
nor U5948 (N_5948,N_4372,N_3826);
and U5949 (N_5949,N_2733,N_4899);
and U5950 (N_5950,N_4288,N_3020);
nand U5951 (N_5951,N_2551,N_4400);
xnor U5952 (N_5952,N_3662,N_4806);
nand U5953 (N_5953,N_3732,N_4759);
nand U5954 (N_5954,N_2701,N_3904);
nand U5955 (N_5955,N_3688,N_3207);
nor U5956 (N_5956,N_4578,N_3702);
or U5957 (N_5957,N_4702,N_4747);
or U5958 (N_5958,N_4993,N_4537);
or U5959 (N_5959,N_3011,N_3692);
nand U5960 (N_5960,N_3851,N_2723);
nand U5961 (N_5961,N_2812,N_3886);
and U5962 (N_5962,N_3098,N_2644);
or U5963 (N_5963,N_4399,N_4239);
nand U5964 (N_5964,N_4514,N_4330);
and U5965 (N_5965,N_3306,N_3925);
nor U5966 (N_5966,N_3757,N_4493);
nor U5967 (N_5967,N_3666,N_4678);
nor U5968 (N_5968,N_4635,N_3640);
nor U5969 (N_5969,N_3132,N_2961);
xor U5970 (N_5970,N_2724,N_3615);
or U5971 (N_5971,N_4034,N_4188);
xor U5972 (N_5972,N_2941,N_4429);
nand U5973 (N_5973,N_2931,N_4126);
xnor U5974 (N_5974,N_3602,N_4099);
nor U5975 (N_5975,N_3179,N_2708);
nand U5976 (N_5976,N_3945,N_4388);
nor U5977 (N_5977,N_2835,N_4501);
or U5978 (N_5978,N_4885,N_4146);
and U5979 (N_5979,N_3689,N_4987);
nor U5980 (N_5980,N_4961,N_4515);
xnor U5981 (N_5981,N_3101,N_2643);
or U5982 (N_5982,N_3304,N_4865);
or U5983 (N_5983,N_4168,N_2586);
and U5984 (N_5984,N_4150,N_4562);
and U5985 (N_5985,N_4152,N_4401);
nor U5986 (N_5986,N_2621,N_4072);
or U5987 (N_5987,N_4788,N_4361);
xor U5988 (N_5988,N_4555,N_4783);
or U5989 (N_5989,N_3003,N_4882);
and U5990 (N_5990,N_2729,N_4632);
xnor U5991 (N_5991,N_4234,N_2766);
nor U5992 (N_5992,N_4508,N_3956);
nor U5993 (N_5993,N_4122,N_4752);
and U5994 (N_5994,N_4225,N_4782);
nand U5995 (N_5995,N_2502,N_4592);
or U5996 (N_5996,N_2856,N_4574);
nand U5997 (N_5997,N_2992,N_3308);
nand U5998 (N_5998,N_2667,N_4433);
nor U5999 (N_5999,N_4411,N_2869);
nor U6000 (N_6000,N_2545,N_3926);
nand U6001 (N_6001,N_2519,N_4409);
nand U6002 (N_6002,N_2877,N_4991);
and U6003 (N_6003,N_3975,N_3933);
or U6004 (N_6004,N_3151,N_4369);
nor U6005 (N_6005,N_3916,N_4393);
and U6006 (N_6006,N_4289,N_4911);
nor U6007 (N_6007,N_3825,N_2893);
or U6008 (N_6008,N_4500,N_3921);
and U6009 (N_6009,N_4482,N_4298);
and U6010 (N_6010,N_2847,N_3052);
or U6011 (N_6011,N_3455,N_3349);
nor U6012 (N_6012,N_4673,N_4314);
or U6013 (N_6013,N_4846,N_3509);
or U6014 (N_6014,N_2854,N_4640);
and U6015 (N_6015,N_4335,N_3969);
and U6016 (N_6016,N_3566,N_3458);
nand U6017 (N_6017,N_3084,N_3570);
nor U6018 (N_6018,N_4430,N_4271);
nor U6019 (N_6019,N_2552,N_4887);
nand U6020 (N_6020,N_2742,N_3412);
and U6021 (N_6021,N_2841,N_4358);
nand U6022 (N_6022,N_4165,N_3053);
nor U6023 (N_6023,N_3958,N_4742);
or U6024 (N_6024,N_3928,N_3068);
or U6025 (N_6025,N_4387,N_4706);
and U6026 (N_6026,N_3582,N_3954);
xnor U6027 (N_6027,N_3278,N_4003);
nor U6028 (N_6028,N_3856,N_4724);
or U6029 (N_6029,N_2882,N_4755);
nor U6030 (N_6030,N_3528,N_4055);
and U6031 (N_6031,N_3977,N_2618);
nor U6032 (N_6032,N_4465,N_3429);
nand U6033 (N_6033,N_4145,N_2933);
nor U6034 (N_6034,N_3318,N_2596);
xor U6035 (N_6035,N_2760,N_4905);
nand U6036 (N_6036,N_4320,N_3182);
or U6037 (N_6037,N_3699,N_2719);
or U6038 (N_6038,N_4164,N_3226);
nor U6039 (N_6039,N_3244,N_4053);
and U6040 (N_6040,N_3205,N_4167);
or U6041 (N_6041,N_3837,N_4480);
or U6042 (N_6042,N_4402,N_2952);
nand U6043 (N_6043,N_3878,N_2870);
nor U6044 (N_6044,N_3019,N_4893);
and U6045 (N_6045,N_4292,N_4252);
or U6046 (N_6046,N_3794,N_4204);
nand U6047 (N_6047,N_4442,N_3270);
nand U6048 (N_6048,N_2512,N_3230);
nand U6049 (N_6049,N_4612,N_4836);
and U6050 (N_6050,N_3241,N_3313);
nand U6051 (N_6051,N_2713,N_3097);
or U6052 (N_6052,N_2950,N_4485);
xnor U6053 (N_6053,N_4151,N_4318);
nor U6054 (N_6054,N_4653,N_4845);
nand U6055 (N_6055,N_3729,N_2779);
or U6056 (N_6056,N_4039,N_2795);
nand U6057 (N_6057,N_4777,N_2647);
nand U6058 (N_6058,N_4866,N_4484);
and U6059 (N_6059,N_3636,N_4709);
or U6060 (N_6060,N_4394,N_2574);
nand U6061 (N_6061,N_3018,N_4349);
nand U6062 (N_6062,N_4477,N_3713);
or U6063 (N_6063,N_4498,N_3497);
or U6064 (N_6064,N_3618,N_4346);
or U6065 (N_6065,N_2738,N_2631);
nand U6066 (N_6066,N_3250,N_2554);
or U6067 (N_6067,N_3766,N_3477);
and U6068 (N_6068,N_3181,N_2585);
nand U6069 (N_6069,N_4908,N_2704);
nand U6070 (N_6070,N_2658,N_2751);
or U6071 (N_6071,N_2879,N_3238);
and U6072 (N_6072,N_3402,N_3510);
or U6073 (N_6073,N_2897,N_3242);
nand U6074 (N_6074,N_4304,N_4020);
or U6075 (N_6075,N_2700,N_4869);
or U6076 (N_6076,N_3074,N_3410);
nor U6077 (N_6077,N_2711,N_4497);
and U6078 (N_6078,N_4116,N_3046);
or U6079 (N_6079,N_3060,N_4437);
or U6080 (N_6080,N_4275,N_3902);
nand U6081 (N_6081,N_3980,N_3529);
or U6082 (N_6082,N_3994,N_3839);
or U6083 (N_6083,N_3237,N_3262);
xnor U6084 (N_6084,N_4462,N_2645);
nand U6085 (N_6085,N_4956,N_4990);
or U6086 (N_6086,N_4463,N_3421);
nor U6087 (N_6087,N_3536,N_4671);
nand U6088 (N_6088,N_4867,N_3654);
and U6089 (N_6089,N_4056,N_2770);
nor U6090 (N_6090,N_3193,N_2934);
nand U6091 (N_6091,N_2883,N_4637);
nand U6092 (N_6092,N_4716,N_4354);
and U6093 (N_6093,N_3448,N_3648);
nand U6094 (N_6094,N_4432,N_2514);
xor U6095 (N_6095,N_4098,N_2624);
nand U6096 (N_6096,N_2564,N_2663);
and U6097 (N_6097,N_4505,N_4030);
and U6098 (N_6098,N_4621,N_4503);
and U6099 (N_6099,N_3386,N_3807);
nor U6100 (N_6100,N_4856,N_3302);
nor U6101 (N_6101,N_4740,N_2793);
or U6102 (N_6102,N_4365,N_4472);
or U6103 (N_6103,N_2775,N_4753);
or U6104 (N_6104,N_2569,N_3219);
and U6105 (N_6105,N_3901,N_3037);
or U6106 (N_6106,N_2958,N_4541);
and U6107 (N_6107,N_3597,N_3059);
or U6108 (N_6108,N_2752,N_3987);
or U6109 (N_6109,N_4652,N_3819);
nor U6110 (N_6110,N_2568,N_3391);
nand U6111 (N_6111,N_2755,N_4235);
or U6112 (N_6112,N_2786,N_4025);
or U6113 (N_6113,N_2671,N_2745);
or U6114 (N_6114,N_3533,N_3982);
nor U6115 (N_6115,N_2906,N_3311);
nor U6116 (N_6116,N_3885,N_3809);
nand U6117 (N_6117,N_3430,N_4043);
nor U6118 (N_6118,N_2757,N_4568);
nand U6119 (N_6119,N_4516,N_4110);
nor U6120 (N_6120,N_4581,N_2864);
nand U6121 (N_6121,N_3353,N_3569);
nand U6122 (N_6122,N_3411,N_4017);
nand U6123 (N_6123,N_4302,N_3563);
and U6124 (N_6124,N_3094,N_4877);
or U6125 (N_6125,N_4450,N_4322);
or U6126 (N_6126,N_4906,N_3280);
nor U6127 (N_6127,N_4236,N_4441);
nand U6128 (N_6128,N_2662,N_3953);
nor U6129 (N_6129,N_4749,N_4603);
nand U6130 (N_6130,N_3194,N_4876);
nand U6131 (N_6131,N_3075,N_3064);
or U6132 (N_6132,N_3317,N_4774);
xnor U6133 (N_6133,N_3106,N_2852);
nand U6134 (N_6134,N_2595,N_2878);
nand U6135 (N_6135,N_2953,N_3463);
or U6136 (N_6136,N_4147,N_3437);
and U6137 (N_6137,N_2851,N_3695);
or U6138 (N_6138,N_2535,N_4563);
and U6139 (N_6139,N_4309,N_4779);
or U6140 (N_6140,N_2689,N_4038);
nand U6141 (N_6141,N_2926,N_3622);
nor U6142 (N_6142,N_2797,N_3089);
or U6143 (N_6143,N_3036,N_2718);
and U6144 (N_6144,N_2913,N_3027);
or U6145 (N_6145,N_3167,N_4980);
nor U6146 (N_6146,N_3394,N_2550);
nor U6147 (N_6147,N_2873,N_3190);
nor U6148 (N_6148,N_3268,N_4035);
nand U6149 (N_6149,N_3759,N_2560);
nand U6150 (N_6150,N_2521,N_2526);
nor U6151 (N_6151,N_3407,N_3040);
or U6152 (N_6152,N_4175,N_3466);
nand U6153 (N_6153,N_3066,N_4531);
or U6154 (N_6154,N_3305,N_4726);
nand U6155 (N_6155,N_4878,N_3668);
or U6156 (N_6156,N_4459,N_4415);
and U6157 (N_6157,N_3985,N_2875);
xnor U6158 (N_6158,N_2638,N_4909);
or U6159 (N_6159,N_2843,N_3763);
and U6160 (N_6160,N_3285,N_2511);
nand U6161 (N_6161,N_3006,N_2553);
and U6162 (N_6162,N_4245,N_4007);
nor U6163 (N_6163,N_4999,N_4602);
and U6164 (N_6164,N_3324,N_4769);
and U6165 (N_6165,N_2814,N_4208);
nor U6166 (N_6166,N_4662,N_3730);
or U6167 (N_6167,N_4550,N_4617);
nor U6168 (N_6168,N_4113,N_4207);
and U6169 (N_6169,N_2650,N_2709);
nand U6170 (N_6170,N_4006,N_2924);
nand U6171 (N_6171,N_3287,N_2641);
and U6172 (N_6172,N_3716,N_3630);
nor U6173 (N_6173,N_3643,N_3800);
and U6174 (N_6174,N_2672,N_3524);
or U6175 (N_6175,N_2868,N_3100);
and U6176 (N_6176,N_4094,N_2584);
nand U6177 (N_6177,N_2988,N_2994);
nand U6178 (N_6178,N_3127,N_3898);
nor U6179 (N_6179,N_3323,N_4756);
nand U6180 (N_6180,N_4770,N_3503);
nor U6181 (N_6181,N_3229,N_4767);
or U6182 (N_6182,N_4972,N_3005);
or U6183 (N_6183,N_3276,N_3978);
nor U6184 (N_6184,N_4262,N_4189);
and U6185 (N_6185,N_3041,N_2506);
or U6186 (N_6186,N_3600,N_3599);
and U6187 (N_6187,N_4676,N_3624);
or U6188 (N_6188,N_4681,N_2515);
nor U6189 (N_6189,N_3868,N_2817);
and U6190 (N_6190,N_3493,N_3023);
or U6191 (N_6191,N_3952,N_3559);
nor U6192 (N_6192,N_2894,N_4794);
and U6193 (N_6193,N_3322,N_3586);
xor U6194 (N_6194,N_4591,N_4052);
and U6195 (N_6195,N_3930,N_3804);
nor U6196 (N_6196,N_3896,N_4089);
nand U6197 (N_6197,N_3607,N_3335);
nand U6198 (N_6198,N_2925,N_3517);
xnor U6199 (N_6199,N_4554,N_3257);
nor U6200 (N_6200,N_4310,N_3545);
nor U6201 (N_6201,N_4378,N_2787);
nand U6202 (N_6202,N_4874,N_2684);
xor U6203 (N_6203,N_4533,N_3008);
and U6204 (N_6204,N_4850,N_3395);
nor U6205 (N_6205,N_3247,N_4971);
nor U6206 (N_6206,N_2830,N_2682);
nand U6207 (N_6207,N_4778,N_4710);
nor U6208 (N_6208,N_4457,N_4763);
or U6209 (N_6209,N_4588,N_2969);
nand U6210 (N_6210,N_4496,N_4088);
nand U6211 (N_6211,N_3616,N_4413);
or U6212 (N_6212,N_4049,N_4923);
nand U6213 (N_6213,N_3339,N_4835);
nor U6214 (N_6214,N_3290,N_4093);
and U6215 (N_6215,N_2613,N_4397);
or U6216 (N_6216,N_2942,N_2944);
nor U6217 (N_6217,N_4326,N_4137);
and U6218 (N_6218,N_3072,N_3360);
nand U6219 (N_6219,N_4842,N_4525);
nor U6220 (N_6220,N_3500,N_3523);
nand U6221 (N_6221,N_3175,N_4823);
nor U6222 (N_6222,N_3515,N_4133);
and U6223 (N_6223,N_3090,N_3201);
nor U6224 (N_6224,N_3291,N_3679);
xnor U6225 (N_6225,N_4959,N_3309);
and U6226 (N_6226,N_3328,N_3919);
or U6227 (N_6227,N_4408,N_4119);
nor U6228 (N_6228,N_3641,N_4675);
nor U6229 (N_6229,N_4295,N_4076);
nand U6230 (N_6230,N_3146,N_4139);
nand U6231 (N_6231,N_2608,N_3344);
or U6232 (N_6232,N_4925,N_4490);
and U6233 (N_6233,N_3811,N_3222);
or U6234 (N_6234,N_3413,N_4587);
or U6235 (N_6235,N_3822,N_4721);
nand U6236 (N_6236,N_2801,N_4852);
nand U6237 (N_6237,N_3374,N_3516);
xnor U6238 (N_6238,N_3069,N_4370);
or U6239 (N_6239,N_3384,N_3032);
and U6240 (N_6240,N_2714,N_3842);
xnor U6241 (N_6241,N_2736,N_3091);
nand U6242 (N_6242,N_4350,N_4157);
nor U6243 (N_6243,N_4744,N_4095);
and U6244 (N_6244,N_3220,N_4128);
nor U6245 (N_6245,N_3115,N_3979);
and U6246 (N_6246,N_3035,N_3016);
and U6247 (N_6247,N_4889,N_3836);
nor U6248 (N_6248,N_4634,N_4622);
or U6249 (N_6249,N_3436,N_3362);
and U6250 (N_6250,N_3497,N_2893);
and U6251 (N_6251,N_4140,N_3500);
or U6252 (N_6252,N_4670,N_4099);
nand U6253 (N_6253,N_2780,N_4812);
nand U6254 (N_6254,N_4209,N_2559);
nand U6255 (N_6255,N_4011,N_3844);
or U6256 (N_6256,N_4019,N_2840);
or U6257 (N_6257,N_4263,N_3068);
and U6258 (N_6258,N_4141,N_3648);
nor U6259 (N_6259,N_4139,N_2882);
nor U6260 (N_6260,N_4447,N_3860);
nand U6261 (N_6261,N_3907,N_2986);
and U6262 (N_6262,N_4370,N_4499);
and U6263 (N_6263,N_3269,N_3937);
nand U6264 (N_6264,N_3085,N_3035);
and U6265 (N_6265,N_2962,N_2628);
xnor U6266 (N_6266,N_4898,N_3285);
and U6267 (N_6267,N_3051,N_3712);
or U6268 (N_6268,N_3758,N_3320);
nor U6269 (N_6269,N_4901,N_3194);
nor U6270 (N_6270,N_4013,N_3146);
nor U6271 (N_6271,N_3911,N_4478);
or U6272 (N_6272,N_2696,N_2776);
nand U6273 (N_6273,N_4037,N_4620);
and U6274 (N_6274,N_3775,N_3386);
and U6275 (N_6275,N_3067,N_2911);
and U6276 (N_6276,N_4744,N_2861);
nand U6277 (N_6277,N_4896,N_3091);
nor U6278 (N_6278,N_2862,N_3133);
nor U6279 (N_6279,N_4443,N_3880);
nand U6280 (N_6280,N_2977,N_3106);
nor U6281 (N_6281,N_3776,N_2504);
nand U6282 (N_6282,N_3152,N_3191);
or U6283 (N_6283,N_2648,N_4502);
and U6284 (N_6284,N_2737,N_4575);
nand U6285 (N_6285,N_3941,N_4944);
and U6286 (N_6286,N_2574,N_3541);
or U6287 (N_6287,N_2857,N_3692);
or U6288 (N_6288,N_3101,N_2522);
xor U6289 (N_6289,N_4421,N_4215);
nor U6290 (N_6290,N_3423,N_2541);
nor U6291 (N_6291,N_3206,N_4346);
and U6292 (N_6292,N_3750,N_4821);
and U6293 (N_6293,N_3999,N_4252);
or U6294 (N_6294,N_3134,N_3162);
nand U6295 (N_6295,N_3580,N_2702);
nand U6296 (N_6296,N_3721,N_2568);
nor U6297 (N_6297,N_2788,N_4324);
nand U6298 (N_6298,N_3138,N_3196);
or U6299 (N_6299,N_2799,N_3681);
nor U6300 (N_6300,N_3278,N_4712);
or U6301 (N_6301,N_2654,N_4969);
nand U6302 (N_6302,N_4817,N_2973);
nor U6303 (N_6303,N_4733,N_3709);
and U6304 (N_6304,N_3030,N_3855);
xor U6305 (N_6305,N_4877,N_4806);
and U6306 (N_6306,N_4782,N_4005);
or U6307 (N_6307,N_3854,N_4265);
or U6308 (N_6308,N_3378,N_2577);
or U6309 (N_6309,N_4438,N_3952);
or U6310 (N_6310,N_3745,N_3287);
and U6311 (N_6311,N_4263,N_3032);
or U6312 (N_6312,N_2547,N_4823);
nor U6313 (N_6313,N_3542,N_3820);
nand U6314 (N_6314,N_2963,N_2933);
or U6315 (N_6315,N_3543,N_4255);
and U6316 (N_6316,N_3485,N_3903);
or U6317 (N_6317,N_4363,N_4096);
nand U6318 (N_6318,N_4922,N_4212);
or U6319 (N_6319,N_3198,N_3157);
or U6320 (N_6320,N_4375,N_2562);
nand U6321 (N_6321,N_2908,N_4346);
or U6322 (N_6322,N_3295,N_4282);
and U6323 (N_6323,N_3903,N_2831);
and U6324 (N_6324,N_3177,N_4010);
and U6325 (N_6325,N_4142,N_2697);
nand U6326 (N_6326,N_2885,N_2661);
and U6327 (N_6327,N_2979,N_4451);
nor U6328 (N_6328,N_2790,N_3272);
and U6329 (N_6329,N_4701,N_3430);
xnor U6330 (N_6330,N_4708,N_4792);
nor U6331 (N_6331,N_4908,N_4058);
nand U6332 (N_6332,N_3854,N_4397);
and U6333 (N_6333,N_2580,N_4819);
or U6334 (N_6334,N_3134,N_2656);
nand U6335 (N_6335,N_4151,N_2638);
nor U6336 (N_6336,N_3525,N_4479);
nand U6337 (N_6337,N_2532,N_4868);
nor U6338 (N_6338,N_2787,N_3397);
and U6339 (N_6339,N_4150,N_3599);
or U6340 (N_6340,N_3937,N_2984);
and U6341 (N_6341,N_2954,N_4794);
nor U6342 (N_6342,N_4619,N_4285);
and U6343 (N_6343,N_3110,N_4113);
nand U6344 (N_6344,N_4605,N_4788);
and U6345 (N_6345,N_2843,N_4439);
nand U6346 (N_6346,N_3209,N_3840);
and U6347 (N_6347,N_3631,N_3747);
or U6348 (N_6348,N_4975,N_4326);
nor U6349 (N_6349,N_4255,N_2790);
nand U6350 (N_6350,N_3280,N_2553);
nor U6351 (N_6351,N_3854,N_3674);
or U6352 (N_6352,N_2897,N_4512);
nand U6353 (N_6353,N_3887,N_4875);
and U6354 (N_6354,N_3605,N_4564);
nor U6355 (N_6355,N_4902,N_3658);
nand U6356 (N_6356,N_4697,N_2875);
nor U6357 (N_6357,N_2612,N_4574);
nand U6358 (N_6358,N_4916,N_4555);
nand U6359 (N_6359,N_2713,N_4175);
nor U6360 (N_6360,N_4054,N_4064);
nand U6361 (N_6361,N_2512,N_4184);
nand U6362 (N_6362,N_4940,N_4233);
nand U6363 (N_6363,N_2903,N_3989);
nand U6364 (N_6364,N_4909,N_3588);
and U6365 (N_6365,N_3132,N_4079);
nand U6366 (N_6366,N_3664,N_2702);
and U6367 (N_6367,N_3343,N_4619);
and U6368 (N_6368,N_4571,N_3048);
nand U6369 (N_6369,N_4364,N_2858);
and U6370 (N_6370,N_4072,N_3521);
nand U6371 (N_6371,N_3268,N_2821);
and U6372 (N_6372,N_3916,N_3792);
nand U6373 (N_6373,N_4456,N_3762);
and U6374 (N_6374,N_4310,N_4592);
nand U6375 (N_6375,N_3797,N_4891);
nand U6376 (N_6376,N_4514,N_4270);
and U6377 (N_6377,N_3219,N_3205);
and U6378 (N_6378,N_4350,N_4023);
nand U6379 (N_6379,N_4539,N_4147);
xnor U6380 (N_6380,N_4721,N_2700);
or U6381 (N_6381,N_2875,N_3272);
xor U6382 (N_6382,N_4794,N_4696);
nor U6383 (N_6383,N_3505,N_4639);
nor U6384 (N_6384,N_3163,N_4614);
nor U6385 (N_6385,N_3029,N_2728);
or U6386 (N_6386,N_2557,N_3546);
nand U6387 (N_6387,N_3110,N_4773);
nor U6388 (N_6388,N_3409,N_3223);
nand U6389 (N_6389,N_2530,N_4830);
nand U6390 (N_6390,N_4901,N_4301);
nor U6391 (N_6391,N_4925,N_4246);
and U6392 (N_6392,N_3356,N_2566);
or U6393 (N_6393,N_3541,N_3694);
and U6394 (N_6394,N_4015,N_4899);
or U6395 (N_6395,N_4140,N_4538);
and U6396 (N_6396,N_3359,N_3702);
and U6397 (N_6397,N_4367,N_2890);
nor U6398 (N_6398,N_2704,N_3454);
or U6399 (N_6399,N_4651,N_3789);
nand U6400 (N_6400,N_2525,N_2717);
or U6401 (N_6401,N_4421,N_2823);
nand U6402 (N_6402,N_4118,N_2889);
nand U6403 (N_6403,N_4113,N_4780);
and U6404 (N_6404,N_3852,N_2815);
nand U6405 (N_6405,N_4876,N_2827);
nand U6406 (N_6406,N_3231,N_4486);
nand U6407 (N_6407,N_4723,N_4258);
or U6408 (N_6408,N_4397,N_3176);
and U6409 (N_6409,N_4439,N_4405);
nor U6410 (N_6410,N_4289,N_3513);
xnor U6411 (N_6411,N_4669,N_3123);
or U6412 (N_6412,N_4425,N_4823);
or U6413 (N_6413,N_4415,N_4793);
nor U6414 (N_6414,N_3044,N_2688);
and U6415 (N_6415,N_4889,N_4417);
nand U6416 (N_6416,N_4597,N_3046);
or U6417 (N_6417,N_3033,N_3133);
nand U6418 (N_6418,N_4149,N_3886);
and U6419 (N_6419,N_3978,N_3179);
nand U6420 (N_6420,N_3206,N_4911);
and U6421 (N_6421,N_2627,N_2613);
nand U6422 (N_6422,N_3781,N_3705);
nand U6423 (N_6423,N_3968,N_4911);
nor U6424 (N_6424,N_2826,N_4177);
or U6425 (N_6425,N_4275,N_3860);
and U6426 (N_6426,N_4342,N_2737);
nand U6427 (N_6427,N_4030,N_3427);
or U6428 (N_6428,N_2576,N_4594);
nand U6429 (N_6429,N_2511,N_4303);
or U6430 (N_6430,N_4043,N_3003);
or U6431 (N_6431,N_2817,N_3701);
nand U6432 (N_6432,N_2642,N_2836);
and U6433 (N_6433,N_4817,N_3789);
and U6434 (N_6434,N_3099,N_2692);
and U6435 (N_6435,N_3809,N_4325);
nand U6436 (N_6436,N_3927,N_2529);
or U6437 (N_6437,N_4853,N_3323);
nand U6438 (N_6438,N_4370,N_2894);
nand U6439 (N_6439,N_2770,N_3214);
and U6440 (N_6440,N_4873,N_3750);
or U6441 (N_6441,N_3285,N_4283);
nor U6442 (N_6442,N_2978,N_4319);
nor U6443 (N_6443,N_4840,N_3601);
xnor U6444 (N_6444,N_4734,N_3976);
nor U6445 (N_6445,N_3349,N_4006);
nand U6446 (N_6446,N_4957,N_4375);
and U6447 (N_6447,N_2656,N_3142);
or U6448 (N_6448,N_4320,N_4975);
nor U6449 (N_6449,N_4921,N_4949);
nor U6450 (N_6450,N_2813,N_3883);
nand U6451 (N_6451,N_2798,N_2819);
nand U6452 (N_6452,N_4725,N_4694);
nand U6453 (N_6453,N_4245,N_3959);
nor U6454 (N_6454,N_4297,N_3837);
or U6455 (N_6455,N_3342,N_4234);
nor U6456 (N_6456,N_3162,N_3840);
nor U6457 (N_6457,N_4159,N_3238);
and U6458 (N_6458,N_3212,N_4014);
nand U6459 (N_6459,N_4620,N_2524);
nand U6460 (N_6460,N_4519,N_3378);
and U6461 (N_6461,N_3841,N_2983);
nand U6462 (N_6462,N_4888,N_2704);
nor U6463 (N_6463,N_4651,N_3915);
nor U6464 (N_6464,N_3232,N_3744);
and U6465 (N_6465,N_3544,N_3470);
nand U6466 (N_6466,N_3508,N_4163);
nor U6467 (N_6467,N_2547,N_4163);
nor U6468 (N_6468,N_4284,N_3972);
and U6469 (N_6469,N_2943,N_3211);
or U6470 (N_6470,N_4747,N_3680);
nor U6471 (N_6471,N_2624,N_2837);
and U6472 (N_6472,N_3299,N_4051);
nor U6473 (N_6473,N_4301,N_4232);
and U6474 (N_6474,N_3983,N_4158);
nor U6475 (N_6475,N_2531,N_4097);
nand U6476 (N_6476,N_3324,N_3427);
xnor U6477 (N_6477,N_4822,N_3634);
nor U6478 (N_6478,N_3207,N_3521);
nor U6479 (N_6479,N_4849,N_4390);
or U6480 (N_6480,N_3833,N_4692);
nor U6481 (N_6481,N_2569,N_2810);
nor U6482 (N_6482,N_4384,N_4827);
or U6483 (N_6483,N_3377,N_3717);
nand U6484 (N_6484,N_4172,N_3563);
or U6485 (N_6485,N_4804,N_4183);
xor U6486 (N_6486,N_4552,N_4238);
and U6487 (N_6487,N_2856,N_3643);
and U6488 (N_6488,N_3066,N_3632);
nand U6489 (N_6489,N_3413,N_4874);
and U6490 (N_6490,N_2615,N_4272);
and U6491 (N_6491,N_2543,N_3483);
nand U6492 (N_6492,N_4861,N_2923);
or U6493 (N_6493,N_2521,N_3638);
nor U6494 (N_6494,N_4165,N_3552);
nand U6495 (N_6495,N_4124,N_4955);
and U6496 (N_6496,N_2934,N_4512);
nand U6497 (N_6497,N_2988,N_3098);
xor U6498 (N_6498,N_3144,N_4911);
and U6499 (N_6499,N_4227,N_4698);
xnor U6500 (N_6500,N_3935,N_4025);
or U6501 (N_6501,N_2571,N_4505);
and U6502 (N_6502,N_2769,N_3249);
nand U6503 (N_6503,N_4354,N_3776);
and U6504 (N_6504,N_4045,N_2855);
and U6505 (N_6505,N_2609,N_3038);
nand U6506 (N_6506,N_3812,N_2605);
nand U6507 (N_6507,N_4274,N_4447);
nor U6508 (N_6508,N_2763,N_2778);
xor U6509 (N_6509,N_2776,N_3067);
and U6510 (N_6510,N_4911,N_4366);
and U6511 (N_6511,N_2835,N_4865);
and U6512 (N_6512,N_3041,N_3419);
or U6513 (N_6513,N_2564,N_3196);
or U6514 (N_6514,N_2684,N_4768);
or U6515 (N_6515,N_4013,N_3024);
and U6516 (N_6516,N_4273,N_3212);
nand U6517 (N_6517,N_4149,N_3984);
xnor U6518 (N_6518,N_3277,N_3392);
and U6519 (N_6519,N_2972,N_3126);
or U6520 (N_6520,N_4242,N_4721);
nor U6521 (N_6521,N_4278,N_2584);
or U6522 (N_6522,N_4436,N_3605);
nor U6523 (N_6523,N_3751,N_4634);
nand U6524 (N_6524,N_4328,N_2558);
and U6525 (N_6525,N_3448,N_4355);
or U6526 (N_6526,N_3636,N_4767);
or U6527 (N_6527,N_2761,N_2856);
nor U6528 (N_6528,N_4954,N_4220);
nor U6529 (N_6529,N_3279,N_4191);
nand U6530 (N_6530,N_3219,N_3074);
nor U6531 (N_6531,N_3555,N_3176);
nor U6532 (N_6532,N_3301,N_2834);
or U6533 (N_6533,N_3074,N_4018);
and U6534 (N_6534,N_3556,N_3752);
or U6535 (N_6535,N_3005,N_3198);
nor U6536 (N_6536,N_4471,N_4748);
nand U6537 (N_6537,N_3134,N_3519);
and U6538 (N_6538,N_4633,N_4287);
and U6539 (N_6539,N_3058,N_3739);
nand U6540 (N_6540,N_3316,N_2564);
nand U6541 (N_6541,N_3012,N_3951);
nand U6542 (N_6542,N_4017,N_2765);
and U6543 (N_6543,N_4347,N_3067);
nor U6544 (N_6544,N_3030,N_3013);
xor U6545 (N_6545,N_2690,N_4343);
or U6546 (N_6546,N_4713,N_3905);
nand U6547 (N_6547,N_2652,N_2544);
nor U6548 (N_6548,N_4670,N_4742);
or U6549 (N_6549,N_2599,N_2781);
xnor U6550 (N_6550,N_4519,N_4317);
or U6551 (N_6551,N_4034,N_3543);
nor U6552 (N_6552,N_4805,N_3563);
nand U6553 (N_6553,N_3455,N_3239);
or U6554 (N_6554,N_4885,N_4721);
and U6555 (N_6555,N_3731,N_3958);
or U6556 (N_6556,N_4291,N_4854);
nor U6557 (N_6557,N_4139,N_4500);
xnor U6558 (N_6558,N_4941,N_2829);
or U6559 (N_6559,N_2979,N_2890);
or U6560 (N_6560,N_2673,N_4539);
nor U6561 (N_6561,N_3121,N_4502);
nand U6562 (N_6562,N_3314,N_4632);
nand U6563 (N_6563,N_4347,N_2897);
nor U6564 (N_6564,N_3032,N_3395);
nor U6565 (N_6565,N_3835,N_3507);
and U6566 (N_6566,N_3665,N_2844);
or U6567 (N_6567,N_4844,N_4554);
xnor U6568 (N_6568,N_2808,N_3514);
nor U6569 (N_6569,N_4223,N_3695);
nand U6570 (N_6570,N_2587,N_4095);
or U6571 (N_6571,N_3465,N_4069);
or U6572 (N_6572,N_3348,N_4677);
and U6573 (N_6573,N_2979,N_3938);
and U6574 (N_6574,N_3172,N_3503);
or U6575 (N_6575,N_4536,N_4318);
nor U6576 (N_6576,N_3609,N_4286);
nand U6577 (N_6577,N_4409,N_4687);
nand U6578 (N_6578,N_3382,N_3740);
nand U6579 (N_6579,N_4945,N_4633);
nor U6580 (N_6580,N_4051,N_4433);
and U6581 (N_6581,N_4179,N_4072);
and U6582 (N_6582,N_2539,N_4483);
nand U6583 (N_6583,N_2744,N_3302);
nand U6584 (N_6584,N_2605,N_4849);
xnor U6585 (N_6585,N_2807,N_2968);
or U6586 (N_6586,N_3714,N_4103);
and U6587 (N_6587,N_2702,N_4696);
nand U6588 (N_6588,N_4493,N_3224);
nor U6589 (N_6589,N_4858,N_4690);
or U6590 (N_6590,N_2653,N_4014);
and U6591 (N_6591,N_3801,N_2530);
and U6592 (N_6592,N_2693,N_3096);
nand U6593 (N_6593,N_4729,N_3023);
and U6594 (N_6594,N_3203,N_3021);
and U6595 (N_6595,N_3239,N_3589);
or U6596 (N_6596,N_3375,N_3280);
nor U6597 (N_6597,N_3949,N_2990);
nor U6598 (N_6598,N_4688,N_4287);
nor U6599 (N_6599,N_4815,N_3229);
xnor U6600 (N_6600,N_3909,N_3704);
and U6601 (N_6601,N_4401,N_3608);
or U6602 (N_6602,N_3039,N_3357);
xor U6603 (N_6603,N_4675,N_2789);
nor U6604 (N_6604,N_3413,N_4830);
nor U6605 (N_6605,N_4445,N_3411);
nand U6606 (N_6606,N_3334,N_4510);
nor U6607 (N_6607,N_3487,N_4341);
nor U6608 (N_6608,N_3212,N_3770);
and U6609 (N_6609,N_4901,N_4593);
nand U6610 (N_6610,N_3446,N_4806);
and U6611 (N_6611,N_2880,N_3375);
nand U6612 (N_6612,N_4921,N_2958);
nand U6613 (N_6613,N_3754,N_2678);
and U6614 (N_6614,N_3532,N_4095);
xnor U6615 (N_6615,N_4030,N_4322);
xor U6616 (N_6616,N_3365,N_3183);
xnor U6617 (N_6617,N_3121,N_4710);
and U6618 (N_6618,N_3912,N_2749);
nand U6619 (N_6619,N_4773,N_2995);
or U6620 (N_6620,N_2699,N_2552);
and U6621 (N_6621,N_4552,N_3034);
xnor U6622 (N_6622,N_3793,N_4129);
or U6623 (N_6623,N_2880,N_3441);
nand U6624 (N_6624,N_4559,N_3291);
nand U6625 (N_6625,N_4352,N_3777);
and U6626 (N_6626,N_4208,N_4219);
and U6627 (N_6627,N_4184,N_2992);
and U6628 (N_6628,N_4093,N_4943);
and U6629 (N_6629,N_3712,N_2567);
or U6630 (N_6630,N_3903,N_2854);
or U6631 (N_6631,N_3901,N_3205);
xnor U6632 (N_6632,N_4052,N_2621);
nor U6633 (N_6633,N_4709,N_2674);
nor U6634 (N_6634,N_4101,N_3745);
nand U6635 (N_6635,N_2603,N_4345);
xnor U6636 (N_6636,N_4146,N_3346);
nand U6637 (N_6637,N_4496,N_2505);
xor U6638 (N_6638,N_4406,N_4918);
or U6639 (N_6639,N_3164,N_4896);
or U6640 (N_6640,N_3049,N_4977);
xnor U6641 (N_6641,N_3266,N_3225);
nand U6642 (N_6642,N_2538,N_4590);
nor U6643 (N_6643,N_2684,N_3822);
nor U6644 (N_6644,N_4863,N_3489);
nand U6645 (N_6645,N_4659,N_3173);
xor U6646 (N_6646,N_4424,N_3020);
or U6647 (N_6647,N_4067,N_2844);
nand U6648 (N_6648,N_4353,N_4528);
and U6649 (N_6649,N_2500,N_3936);
nand U6650 (N_6650,N_4108,N_3217);
nor U6651 (N_6651,N_3337,N_2852);
nand U6652 (N_6652,N_3762,N_2741);
xor U6653 (N_6653,N_4355,N_4158);
and U6654 (N_6654,N_4807,N_4086);
and U6655 (N_6655,N_3578,N_4412);
or U6656 (N_6656,N_4697,N_3467);
and U6657 (N_6657,N_3930,N_3905);
nand U6658 (N_6658,N_3029,N_4287);
nand U6659 (N_6659,N_2807,N_4628);
nor U6660 (N_6660,N_3655,N_4465);
nand U6661 (N_6661,N_2909,N_4451);
nand U6662 (N_6662,N_3990,N_4296);
or U6663 (N_6663,N_3366,N_3244);
xnor U6664 (N_6664,N_2839,N_3016);
nand U6665 (N_6665,N_4556,N_2584);
nor U6666 (N_6666,N_2818,N_4006);
and U6667 (N_6667,N_4613,N_2726);
nand U6668 (N_6668,N_3526,N_2788);
nor U6669 (N_6669,N_2561,N_3434);
xnor U6670 (N_6670,N_3473,N_4204);
nand U6671 (N_6671,N_3578,N_2811);
or U6672 (N_6672,N_2541,N_3908);
and U6673 (N_6673,N_4724,N_4460);
or U6674 (N_6674,N_4588,N_4839);
nand U6675 (N_6675,N_3238,N_3875);
nand U6676 (N_6676,N_4825,N_2523);
xor U6677 (N_6677,N_3266,N_4346);
nor U6678 (N_6678,N_4447,N_3522);
nand U6679 (N_6679,N_4815,N_2853);
nor U6680 (N_6680,N_3623,N_4667);
nor U6681 (N_6681,N_4769,N_4756);
or U6682 (N_6682,N_3301,N_3160);
nand U6683 (N_6683,N_3119,N_4298);
nor U6684 (N_6684,N_4913,N_2623);
nor U6685 (N_6685,N_4700,N_3110);
or U6686 (N_6686,N_4245,N_4374);
nand U6687 (N_6687,N_4752,N_4766);
xor U6688 (N_6688,N_3704,N_4129);
nand U6689 (N_6689,N_3441,N_4453);
or U6690 (N_6690,N_4490,N_4717);
or U6691 (N_6691,N_3127,N_2764);
and U6692 (N_6692,N_3803,N_3565);
or U6693 (N_6693,N_3097,N_2774);
and U6694 (N_6694,N_2745,N_4782);
or U6695 (N_6695,N_4605,N_3686);
and U6696 (N_6696,N_4685,N_3017);
nor U6697 (N_6697,N_4341,N_2871);
nand U6698 (N_6698,N_3122,N_4797);
nand U6699 (N_6699,N_2952,N_3218);
nand U6700 (N_6700,N_3758,N_3512);
or U6701 (N_6701,N_2823,N_2869);
nor U6702 (N_6702,N_4463,N_2514);
or U6703 (N_6703,N_2531,N_4590);
xnor U6704 (N_6704,N_3138,N_4742);
nor U6705 (N_6705,N_2924,N_3136);
or U6706 (N_6706,N_3056,N_3149);
and U6707 (N_6707,N_2980,N_4063);
nor U6708 (N_6708,N_4527,N_4205);
nand U6709 (N_6709,N_4423,N_3389);
and U6710 (N_6710,N_4303,N_4429);
nor U6711 (N_6711,N_3615,N_4293);
nand U6712 (N_6712,N_4031,N_4175);
nor U6713 (N_6713,N_4507,N_3367);
or U6714 (N_6714,N_2776,N_3952);
nand U6715 (N_6715,N_2802,N_4077);
xor U6716 (N_6716,N_4808,N_4304);
nand U6717 (N_6717,N_3632,N_4539);
nor U6718 (N_6718,N_4726,N_3369);
nor U6719 (N_6719,N_3559,N_4847);
and U6720 (N_6720,N_2773,N_3386);
or U6721 (N_6721,N_3318,N_4318);
nand U6722 (N_6722,N_4250,N_4553);
or U6723 (N_6723,N_2997,N_4335);
and U6724 (N_6724,N_3910,N_3603);
nand U6725 (N_6725,N_4983,N_2574);
or U6726 (N_6726,N_3182,N_4996);
nor U6727 (N_6727,N_4530,N_4582);
nand U6728 (N_6728,N_3986,N_3713);
xnor U6729 (N_6729,N_3733,N_3097);
and U6730 (N_6730,N_2525,N_2907);
nand U6731 (N_6731,N_3824,N_3760);
or U6732 (N_6732,N_4734,N_4418);
and U6733 (N_6733,N_4467,N_2812);
or U6734 (N_6734,N_3036,N_2560);
nor U6735 (N_6735,N_4976,N_3307);
nand U6736 (N_6736,N_3111,N_4565);
and U6737 (N_6737,N_4864,N_3649);
or U6738 (N_6738,N_4181,N_4205);
or U6739 (N_6739,N_4924,N_3541);
xnor U6740 (N_6740,N_4798,N_4489);
nor U6741 (N_6741,N_4168,N_4202);
nand U6742 (N_6742,N_2813,N_3005);
nor U6743 (N_6743,N_3177,N_3525);
and U6744 (N_6744,N_4509,N_3497);
nand U6745 (N_6745,N_4092,N_4511);
nor U6746 (N_6746,N_4316,N_4096);
or U6747 (N_6747,N_4343,N_4212);
or U6748 (N_6748,N_3361,N_3170);
or U6749 (N_6749,N_3650,N_4421);
and U6750 (N_6750,N_3954,N_2906);
nor U6751 (N_6751,N_3267,N_3374);
or U6752 (N_6752,N_4189,N_3563);
nor U6753 (N_6753,N_2809,N_4418);
nand U6754 (N_6754,N_3642,N_4693);
or U6755 (N_6755,N_4936,N_4814);
and U6756 (N_6756,N_3789,N_4180);
nand U6757 (N_6757,N_4749,N_2763);
nor U6758 (N_6758,N_3500,N_3166);
and U6759 (N_6759,N_2618,N_4595);
and U6760 (N_6760,N_3175,N_2945);
or U6761 (N_6761,N_2561,N_2658);
nand U6762 (N_6762,N_3035,N_3461);
xor U6763 (N_6763,N_3434,N_2693);
and U6764 (N_6764,N_2890,N_3835);
or U6765 (N_6765,N_3297,N_4967);
xor U6766 (N_6766,N_2876,N_4153);
nand U6767 (N_6767,N_4119,N_3981);
nor U6768 (N_6768,N_3874,N_3496);
nand U6769 (N_6769,N_3980,N_4902);
nand U6770 (N_6770,N_4323,N_4621);
nand U6771 (N_6771,N_3654,N_4567);
nand U6772 (N_6772,N_3096,N_2500);
xor U6773 (N_6773,N_3377,N_3462);
nor U6774 (N_6774,N_2818,N_4991);
and U6775 (N_6775,N_2525,N_4805);
or U6776 (N_6776,N_4817,N_4793);
nor U6777 (N_6777,N_3350,N_3503);
nand U6778 (N_6778,N_3876,N_3633);
nor U6779 (N_6779,N_3860,N_2844);
nand U6780 (N_6780,N_3751,N_3465);
nand U6781 (N_6781,N_4431,N_3627);
nand U6782 (N_6782,N_4596,N_3605);
nor U6783 (N_6783,N_4097,N_4625);
nor U6784 (N_6784,N_3318,N_4087);
or U6785 (N_6785,N_2860,N_2959);
nor U6786 (N_6786,N_4981,N_3450);
nor U6787 (N_6787,N_4534,N_3055);
or U6788 (N_6788,N_3747,N_2959);
nor U6789 (N_6789,N_2896,N_3828);
and U6790 (N_6790,N_3921,N_3979);
and U6791 (N_6791,N_4142,N_4614);
nand U6792 (N_6792,N_3810,N_3113);
or U6793 (N_6793,N_3241,N_3149);
nand U6794 (N_6794,N_3806,N_3411);
nor U6795 (N_6795,N_4375,N_3870);
nand U6796 (N_6796,N_3587,N_2636);
nand U6797 (N_6797,N_2994,N_3802);
and U6798 (N_6798,N_3679,N_4163);
nor U6799 (N_6799,N_4374,N_3390);
nor U6800 (N_6800,N_4814,N_3963);
nand U6801 (N_6801,N_2638,N_2851);
or U6802 (N_6802,N_4612,N_4791);
and U6803 (N_6803,N_2661,N_2915);
xnor U6804 (N_6804,N_4538,N_4452);
xor U6805 (N_6805,N_2918,N_3504);
nor U6806 (N_6806,N_3070,N_4637);
and U6807 (N_6807,N_4808,N_3312);
or U6808 (N_6808,N_3823,N_3891);
or U6809 (N_6809,N_4257,N_3702);
nand U6810 (N_6810,N_2650,N_4074);
and U6811 (N_6811,N_3164,N_2793);
and U6812 (N_6812,N_4263,N_2838);
nand U6813 (N_6813,N_3997,N_4669);
and U6814 (N_6814,N_3272,N_3237);
nand U6815 (N_6815,N_3224,N_3621);
xnor U6816 (N_6816,N_4842,N_3277);
nor U6817 (N_6817,N_2637,N_2698);
or U6818 (N_6818,N_3696,N_2845);
and U6819 (N_6819,N_4108,N_2779);
and U6820 (N_6820,N_2938,N_4647);
nand U6821 (N_6821,N_2715,N_3359);
or U6822 (N_6822,N_3538,N_2887);
or U6823 (N_6823,N_3434,N_3375);
or U6824 (N_6824,N_4160,N_3969);
and U6825 (N_6825,N_4622,N_2728);
or U6826 (N_6826,N_3089,N_3855);
and U6827 (N_6827,N_4382,N_3082);
nor U6828 (N_6828,N_2810,N_3267);
nand U6829 (N_6829,N_3603,N_4038);
or U6830 (N_6830,N_4741,N_3653);
or U6831 (N_6831,N_3031,N_2706);
xnor U6832 (N_6832,N_2520,N_3825);
nor U6833 (N_6833,N_3502,N_4468);
xor U6834 (N_6834,N_4404,N_4531);
nand U6835 (N_6835,N_3265,N_3373);
and U6836 (N_6836,N_3999,N_4879);
nand U6837 (N_6837,N_3626,N_2616);
or U6838 (N_6838,N_2704,N_4264);
or U6839 (N_6839,N_3931,N_4072);
or U6840 (N_6840,N_2570,N_2970);
or U6841 (N_6841,N_4811,N_3411);
nand U6842 (N_6842,N_2977,N_2879);
xor U6843 (N_6843,N_4646,N_3758);
and U6844 (N_6844,N_4356,N_2872);
nor U6845 (N_6845,N_3797,N_3445);
and U6846 (N_6846,N_4963,N_2688);
nand U6847 (N_6847,N_3096,N_2855);
and U6848 (N_6848,N_3202,N_2613);
and U6849 (N_6849,N_4500,N_3377);
nor U6850 (N_6850,N_3787,N_2573);
nor U6851 (N_6851,N_4897,N_3503);
nor U6852 (N_6852,N_4802,N_4167);
or U6853 (N_6853,N_3872,N_3032);
and U6854 (N_6854,N_3421,N_4701);
nand U6855 (N_6855,N_3594,N_3531);
nor U6856 (N_6856,N_4651,N_3838);
and U6857 (N_6857,N_4766,N_3970);
or U6858 (N_6858,N_4308,N_3646);
and U6859 (N_6859,N_4065,N_3497);
or U6860 (N_6860,N_3288,N_2798);
or U6861 (N_6861,N_3511,N_4803);
and U6862 (N_6862,N_4786,N_3183);
nand U6863 (N_6863,N_4973,N_3781);
nand U6864 (N_6864,N_2731,N_4587);
or U6865 (N_6865,N_3018,N_4810);
and U6866 (N_6866,N_3590,N_4999);
or U6867 (N_6867,N_4819,N_4815);
nand U6868 (N_6868,N_3171,N_3994);
nor U6869 (N_6869,N_3558,N_4203);
nor U6870 (N_6870,N_4775,N_3147);
xnor U6871 (N_6871,N_4291,N_2980);
or U6872 (N_6872,N_4590,N_4775);
and U6873 (N_6873,N_4490,N_4590);
nand U6874 (N_6874,N_3051,N_4578);
nand U6875 (N_6875,N_3138,N_2798);
or U6876 (N_6876,N_3354,N_3686);
or U6877 (N_6877,N_3949,N_4138);
nand U6878 (N_6878,N_3272,N_4011);
nand U6879 (N_6879,N_3103,N_3320);
or U6880 (N_6880,N_3922,N_4514);
nand U6881 (N_6881,N_4100,N_3092);
and U6882 (N_6882,N_3457,N_3907);
or U6883 (N_6883,N_3343,N_3733);
xor U6884 (N_6884,N_4391,N_2894);
and U6885 (N_6885,N_3126,N_4056);
xor U6886 (N_6886,N_4133,N_3147);
nor U6887 (N_6887,N_4001,N_4714);
nand U6888 (N_6888,N_4451,N_4593);
or U6889 (N_6889,N_2532,N_3915);
nor U6890 (N_6890,N_3794,N_3078);
nor U6891 (N_6891,N_4431,N_2604);
nand U6892 (N_6892,N_4678,N_4569);
and U6893 (N_6893,N_3274,N_2529);
nand U6894 (N_6894,N_4999,N_4696);
nor U6895 (N_6895,N_2586,N_4175);
xnor U6896 (N_6896,N_4637,N_3880);
or U6897 (N_6897,N_3142,N_4486);
nand U6898 (N_6898,N_3048,N_4759);
or U6899 (N_6899,N_4172,N_4671);
nand U6900 (N_6900,N_4488,N_3873);
nor U6901 (N_6901,N_2711,N_4500);
and U6902 (N_6902,N_2524,N_3881);
and U6903 (N_6903,N_2928,N_3289);
nor U6904 (N_6904,N_2963,N_3186);
nand U6905 (N_6905,N_3363,N_2752);
nor U6906 (N_6906,N_2755,N_2716);
nor U6907 (N_6907,N_4366,N_3022);
xnor U6908 (N_6908,N_4972,N_4880);
xnor U6909 (N_6909,N_3036,N_4603);
nor U6910 (N_6910,N_3937,N_2585);
nand U6911 (N_6911,N_4720,N_3104);
nor U6912 (N_6912,N_4337,N_4426);
and U6913 (N_6913,N_4753,N_3222);
and U6914 (N_6914,N_4126,N_3312);
and U6915 (N_6915,N_3302,N_4148);
nor U6916 (N_6916,N_2818,N_4359);
nand U6917 (N_6917,N_3528,N_4421);
nand U6918 (N_6918,N_3541,N_4297);
nor U6919 (N_6919,N_4886,N_2626);
xor U6920 (N_6920,N_2610,N_4251);
and U6921 (N_6921,N_3702,N_2616);
nor U6922 (N_6922,N_2672,N_3057);
nor U6923 (N_6923,N_4759,N_2792);
nand U6924 (N_6924,N_4481,N_3372);
or U6925 (N_6925,N_4209,N_4880);
or U6926 (N_6926,N_4388,N_2713);
or U6927 (N_6927,N_4546,N_4510);
nor U6928 (N_6928,N_3121,N_4702);
and U6929 (N_6929,N_3947,N_3992);
nand U6930 (N_6930,N_4822,N_3761);
nand U6931 (N_6931,N_3514,N_2536);
or U6932 (N_6932,N_4867,N_2762);
and U6933 (N_6933,N_3447,N_3381);
nand U6934 (N_6934,N_4019,N_4081);
nor U6935 (N_6935,N_2971,N_2865);
nand U6936 (N_6936,N_3821,N_3018);
or U6937 (N_6937,N_2694,N_4051);
or U6938 (N_6938,N_3578,N_4456);
nor U6939 (N_6939,N_2705,N_3290);
and U6940 (N_6940,N_4133,N_4674);
or U6941 (N_6941,N_4208,N_2992);
or U6942 (N_6942,N_4705,N_3629);
and U6943 (N_6943,N_2639,N_4283);
nand U6944 (N_6944,N_4964,N_3784);
and U6945 (N_6945,N_3306,N_3800);
and U6946 (N_6946,N_4437,N_4203);
nand U6947 (N_6947,N_3129,N_3069);
nand U6948 (N_6948,N_4250,N_4547);
or U6949 (N_6949,N_4861,N_3243);
nand U6950 (N_6950,N_4643,N_3749);
nand U6951 (N_6951,N_3396,N_2884);
nor U6952 (N_6952,N_3593,N_4498);
nand U6953 (N_6953,N_4310,N_2623);
nor U6954 (N_6954,N_4501,N_4581);
and U6955 (N_6955,N_4920,N_3663);
or U6956 (N_6956,N_4998,N_4337);
nand U6957 (N_6957,N_4435,N_3079);
nor U6958 (N_6958,N_4845,N_3029);
nor U6959 (N_6959,N_4359,N_2741);
or U6960 (N_6960,N_3737,N_4408);
nor U6961 (N_6961,N_2845,N_4084);
and U6962 (N_6962,N_3764,N_3546);
xnor U6963 (N_6963,N_4167,N_3795);
or U6964 (N_6964,N_4215,N_4563);
nor U6965 (N_6965,N_3506,N_3970);
and U6966 (N_6966,N_4608,N_3690);
and U6967 (N_6967,N_3820,N_2732);
or U6968 (N_6968,N_3437,N_4308);
nor U6969 (N_6969,N_3826,N_4467);
or U6970 (N_6970,N_3251,N_3468);
nor U6971 (N_6971,N_2724,N_3864);
or U6972 (N_6972,N_4979,N_2795);
nor U6973 (N_6973,N_2794,N_2759);
and U6974 (N_6974,N_2578,N_2542);
or U6975 (N_6975,N_4103,N_4736);
nor U6976 (N_6976,N_4391,N_4010);
and U6977 (N_6977,N_4967,N_4341);
or U6978 (N_6978,N_2806,N_3648);
nor U6979 (N_6979,N_3176,N_4186);
and U6980 (N_6980,N_2733,N_4021);
nor U6981 (N_6981,N_3035,N_4634);
or U6982 (N_6982,N_4608,N_3645);
nand U6983 (N_6983,N_3336,N_4338);
or U6984 (N_6984,N_3390,N_4055);
and U6985 (N_6985,N_3644,N_2567);
nand U6986 (N_6986,N_2984,N_3563);
or U6987 (N_6987,N_4525,N_3728);
and U6988 (N_6988,N_2594,N_2578);
or U6989 (N_6989,N_4629,N_4677);
xor U6990 (N_6990,N_4087,N_2710);
nor U6991 (N_6991,N_4950,N_4244);
or U6992 (N_6992,N_3664,N_4318);
or U6993 (N_6993,N_3400,N_3408);
nand U6994 (N_6994,N_3561,N_4435);
and U6995 (N_6995,N_3485,N_3017);
nor U6996 (N_6996,N_3101,N_2774);
nor U6997 (N_6997,N_2841,N_4172);
and U6998 (N_6998,N_4055,N_2655);
and U6999 (N_6999,N_3424,N_3087);
and U7000 (N_7000,N_4863,N_4708);
or U7001 (N_7001,N_3366,N_4129);
nor U7002 (N_7002,N_2981,N_4037);
and U7003 (N_7003,N_3454,N_2983);
or U7004 (N_7004,N_2519,N_3590);
nand U7005 (N_7005,N_3988,N_4509);
nand U7006 (N_7006,N_4849,N_3864);
nor U7007 (N_7007,N_3947,N_3278);
nor U7008 (N_7008,N_3222,N_4676);
nor U7009 (N_7009,N_3571,N_4055);
or U7010 (N_7010,N_4977,N_4229);
and U7011 (N_7011,N_3585,N_3165);
nand U7012 (N_7012,N_4728,N_3661);
or U7013 (N_7013,N_3809,N_3633);
and U7014 (N_7014,N_4695,N_3371);
xor U7015 (N_7015,N_4391,N_2821);
nor U7016 (N_7016,N_3333,N_4548);
nand U7017 (N_7017,N_3629,N_2884);
or U7018 (N_7018,N_3183,N_4245);
or U7019 (N_7019,N_2836,N_2666);
and U7020 (N_7020,N_3607,N_3250);
nor U7021 (N_7021,N_3784,N_3558);
xnor U7022 (N_7022,N_4287,N_2933);
and U7023 (N_7023,N_3419,N_2986);
xnor U7024 (N_7024,N_4504,N_3161);
or U7025 (N_7025,N_4647,N_4575);
or U7026 (N_7026,N_4833,N_3147);
nand U7027 (N_7027,N_4388,N_4632);
nand U7028 (N_7028,N_4760,N_2633);
xnor U7029 (N_7029,N_4164,N_3557);
and U7030 (N_7030,N_4170,N_4622);
xor U7031 (N_7031,N_4283,N_4749);
nand U7032 (N_7032,N_3585,N_3879);
or U7033 (N_7033,N_4086,N_4369);
nor U7034 (N_7034,N_3262,N_4331);
nand U7035 (N_7035,N_3087,N_3669);
nor U7036 (N_7036,N_3969,N_4483);
or U7037 (N_7037,N_3624,N_2760);
nand U7038 (N_7038,N_3097,N_4528);
or U7039 (N_7039,N_4681,N_2518);
or U7040 (N_7040,N_2545,N_4406);
and U7041 (N_7041,N_2658,N_3441);
or U7042 (N_7042,N_2540,N_3461);
xnor U7043 (N_7043,N_4367,N_3026);
or U7044 (N_7044,N_2662,N_2996);
and U7045 (N_7045,N_2760,N_3266);
and U7046 (N_7046,N_3820,N_4289);
nor U7047 (N_7047,N_3869,N_4747);
and U7048 (N_7048,N_2932,N_4918);
and U7049 (N_7049,N_2859,N_2855);
nor U7050 (N_7050,N_4529,N_2843);
or U7051 (N_7051,N_4664,N_4496);
or U7052 (N_7052,N_2925,N_2900);
xnor U7053 (N_7053,N_3072,N_4682);
or U7054 (N_7054,N_2998,N_4858);
xor U7055 (N_7055,N_2998,N_3788);
nand U7056 (N_7056,N_4886,N_3462);
or U7057 (N_7057,N_3017,N_4704);
nand U7058 (N_7058,N_4202,N_3981);
and U7059 (N_7059,N_4084,N_2517);
or U7060 (N_7060,N_3709,N_3119);
nor U7061 (N_7061,N_3449,N_2562);
nand U7062 (N_7062,N_3680,N_4145);
and U7063 (N_7063,N_4505,N_3291);
and U7064 (N_7064,N_3712,N_4385);
nand U7065 (N_7065,N_4404,N_3153);
nand U7066 (N_7066,N_3708,N_4390);
or U7067 (N_7067,N_3269,N_3617);
and U7068 (N_7068,N_3316,N_4614);
or U7069 (N_7069,N_4009,N_4319);
or U7070 (N_7070,N_3704,N_4029);
or U7071 (N_7071,N_4937,N_3950);
or U7072 (N_7072,N_4849,N_4322);
and U7073 (N_7073,N_3474,N_4490);
nand U7074 (N_7074,N_3259,N_3585);
xnor U7075 (N_7075,N_4680,N_3269);
nor U7076 (N_7076,N_2808,N_4626);
nor U7077 (N_7077,N_4197,N_4960);
and U7078 (N_7078,N_3842,N_4966);
or U7079 (N_7079,N_4614,N_4701);
or U7080 (N_7080,N_4400,N_2787);
or U7081 (N_7081,N_3669,N_4533);
nand U7082 (N_7082,N_3199,N_4753);
and U7083 (N_7083,N_3105,N_3396);
xnor U7084 (N_7084,N_3643,N_4241);
or U7085 (N_7085,N_2624,N_4725);
and U7086 (N_7086,N_4459,N_3794);
nor U7087 (N_7087,N_4653,N_3659);
nor U7088 (N_7088,N_4548,N_4733);
nor U7089 (N_7089,N_3625,N_3952);
and U7090 (N_7090,N_4443,N_4177);
nor U7091 (N_7091,N_3336,N_4529);
and U7092 (N_7092,N_3741,N_4166);
nor U7093 (N_7093,N_3531,N_2859);
and U7094 (N_7094,N_2532,N_2950);
nor U7095 (N_7095,N_2980,N_2680);
or U7096 (N_7096,N_4514,N_3538);
and U7097 (N_7097,N_3218,N_4611);
nand U7098 (N_7098,N_2579,N_4638);
nand U7099 (N_7099,N_3963,N_3265);
or U7100 (N_7100,N_3164,N_2648);
xor U7101 (N_7101,N_3969,N_2696);
nand U7102 (N_7102,N_4717,N_3392);
or U7103 (N_7103,N_4326,N_4274);
nor U7104 (N_7104,N_4630,N_3510);
and U7105 (N_7105,N_4264,N_3549);
xor U7106 (N_7106,N_4796,N_4108);
xor U7107 (N_7107,N_3410,N_4293);
or U7108 (N_7108,N_4491,N_3599);
nand U7109 (N_7109,N_3310,N_3853);
xor U7110 (N_7110,N_4042,N_4162);
nor U7111 (N_7111,N_2823,N_3240);
and U7112 (N_7112,N_3308,N_3566);
or U7113 (N_7113,N_3139,N_3875);
or U7114 (N_7114,N_3590,N_2905);
or U7115 (N_7115,N_3692,N_3113);
and U7116 (N_7116,N_4530,N_3900);
and U7117 (N_7117,N_3779,N_2972);
or U7118 (N_7118,N_3480,N_4322);
or U7119 (N_7119,N_4252,N_2759);
nor U7120 (N_7120,N_3912,N_4865);
and U7121 (N_7121,N_3574,N_3120);
and U7122 (N_7122,N_2565,N_3170);
nor U7123 (N_7123,N_4561,N_4205);
nor U7124 (N_7124,N_4525,N_3501);
nor U7125 (N_7125,N_3704,N_3059);
or U7126 (N_7126,N_4375,N_3852);
nand U7127 (N_7127,N_3795,N_3017);
and U7128 (N_7128,N_3798,N_3618);
nor U7129 (N_7129,N_4240,N_4834);
nor U7130 (N_7130,N_2707,N_4350);
nand U7131 (N_7131,N_4360,N_3053);
and U7132 (N_7132,N_4431,N_4675);
xor U7133 (N_7133,N_4565,N_4877);
nor U7134 (N_7134,N_4597,N_2811);
and U7135 (N_7135,N_3857,N_3047);
or U7136 (N_7136,N_2800,N_2625);
xnor U7137 (N_7137,N_4525,N_4500);
and U7138 (N_7138,N_3190,N_3201);
or U7139 (N_7139,N_2840,N_3602);
and U7140 (N_7140,N_2512,N_4672);
or U7141 (N_7141,N_4514,N_4122);
nor U7142 (N_7142,N_4783,N_4946);
or U7143 (N_7143,N_2662,N_3972);
or U7144 (N_7144,N_3345,N_3085);
nand U7145 (N_7145,N_4474,N_4254);
nand U7146 (N_7146,N_4408,N_3219);
xor U7147 (N_7147,N_3396,N_4220);
or U7148 (N_7148,N_2847,N_2845);
or U7149 (N_7149,N_3892,N_4670);
or U7150 (N_7150,N_3225,N_2617);
nand U7151 (N_7151,N_2525,N_4023);
or U7152 (N_7152,N_4882,N_4947);
or U7153 (N_7153,N_4604,N_4723);
or U7154 (N_7154,N_4325,N_4068);
or U7155 (N_7155,N_4305,N_4001);
nand U7156 (N_7156,N_3349,N_3944);
and U7157 (N_7157,N_4676,N_3076);
and U7158 (N_7158,N_4296,N_2967);
and U7159 (N_7159,N_3118,N_3496);
nor U7160 (N_7160,N_3607,N_4953);
and U7161 (N_7161,N_3249,N_4809);
xor U7162 (N_7162,N_4077,N_3996);
nand U7163 (N_7163,N_4852,N_3300);
nand U7164 (N_7164,N_4833,N_3226);
and U7165 (N_7165,N_3354,N_4687);
and U7166 (N_7166,N_4717,N_3154);
or U7167 (N_7167,N_4662,N_4675);
and U7168 (N_7168,N_3968,N_4204);
and U7169 (N_7169,N_2807,N_3944);
and U7170 (N_7170,N_3838,N_3259);
and U7171 (N_7171,N_3188,N_3512);
nand U7172 (N_7172,N_2708,N_3416);
nor U7173 (N_7173,N_4559,N_4775);
and U7174 (N_7174,N_4735,N_3582);
and U7175 (N_7175,N_4923,N_2993);
nor U7176 (N_7176,N_3939,N_4500);
or U7177 (N_7177,N_4611,N_4160);
or U7178 (N_7178,N_3796,N_3141);
nand U7179 (N_7179,N_3278,N_2973);
nand U7180 (N_7180,N_2944,N_4283);
nor U7181 (N_7181,N_4405,N_3658);
and U7182 (N_7182,N_2917,N_3497);
nor U7183 (N_7183,N_4893,N_3020);
and U7184 (N_7184,N_4872,N_3921);
or U7185 (N_7185,N_3823,N_3200);
or U7186 (N_7186,N_2939,N_4795);
or U7187 (N_7187,N_3343,N_3359);
xnor U7188 (N_7188,N_3059,N_4602);
nand U7189 (N_7189,N_4843,N_3744);
nor U7190 (N_7190,N_4977,N_4488);
or U7191 (N_7191,N_3945,N_4791);
nor U7192 (N_7192,N_4198,N_2999);
nand U7193 (N_7193,N_4747,N_3539);
or U7194 (N_7194,N_4788,N_4693);
nor U7195 (N_7195,N_2615,N_3132);
and U7196 (N_7196,N_3169,N_3026);
and U7197 (N_7197,N_3910,N_4746);
and U7198 (N_7198,N_2964,N_3351);
nor U7199 (N_7199,N_4211,N_2765);
or U7200 (N_7200,N_4950,N_3006);
nand U7201 (N_7201,N_3474,N_2617);
and U7202 (N_7202,N_2690,N_4548);
or U7203 (N_7203,N_4335,N_4825);
nand U7204 (N_7204,N_4769,N_2984);
and U7205 (N_7205,N_3665,N_4463);
and U7206 (N_7206,N_3797,N_3742);
and U7207 (N_7207,N_4105,N_4947);
and U7208 (N_7208,N_4463,N_3266);
and U7209 (N_7209,N_3306,N_3571);
xor U7210 (N_7210,N_3047,N_3490);
or U7211 (N_7211,N_4387,N_4846);
nand U7212 (N_7212,N_2715,N_3833);
nand U7213 (N_7213,N_3019,N_2601);
or U7214 (N_7214,N_3787,N_4772);
or U7215 (N_7215,N_2589,N_3203);
or U7216 (N_7216,N_4023,N_4104);
nor U7217 (N_7217,N_4109,N_2595);
or U7218 (N_7218,N_4761,N_2552);
nor U7219 (N_7219,N_3566,N_4274);
or U7220 (N_7220,N_3381,N_3912);
nor U7221 (N_7221,N_4872,N_2850);
xor U7222 (N_7222,N_4476,N_4853);
or U7223 (N_7223,N_3196,N_3277);
or U7224 (N_7224,N_4153,N_2713);
nand U7225 (N_7225,N_3699,N_3094);
nand U7226 (N_7226,N_3279,N_2941);
nor U7227 (N_7227,N_3013,N_2726);
nand U7228 (N_7228,N_4279,N_4373);
or U7229 (N_7229,N_4721,N_3028);
nand U7230 (N_7230,N_4376,N_3585);
or U7231 (N_7231,N_2714,N_3843);
xor U7232 (N_7232,N_2691,N_4554);
nand U7233 (N_7233,N_2918,N_4816);
nand U7234 (N_7234,N_4713,N_2857);
and U7235 (N_7235,N_4049,N_3164);
or U7236 (N_7236,N_3183,N_3196);
nand U7237 (N_7237,N_3848,N_4728);
nand U7238 (N_7238,N_4962,N_2957);
and U7239 (N_7239,N_3771,N_2657);
and U7240 (N_7240,N_3602,N_4764);
nor U7241 (N_7241,N_4804,N_2708);
nand U7242 (N_7242,N_2931,N_4149);
or U7243 (N_7243,N_4905,N_4027);
nand U7244 (N_7244,N_4733,N_3157);
or U7245 (N_7245,N_2901,N_2905);
and U7246 (N_7246,N_2569,N_4186);
nor U7247 (N_7247,N_4697,N_3664);
nor U7248 (N_7248,N_4666,N_3478);
or U7249 (N_7249,N_4709,N_3676);
nand U7250 (N_7250,N_3669,N_4526);
xnor U7251 (N_7251,N_2626,N_3925);
and U7252 (N_7252,N_4588,N_2778);
nand U7253 (N_7253,N_2984,N_3305);
nor U7254 (N_7254,N_4161,N_4967);
and U7255 (N_7255,N_2699,N_3706);
xor U7256 (N_7256,N_3663,N_4071);
or U7257 (N_7257,N_4772,N_2818);
and U7258 (N_7258,N_3485,N_4331);
nor U7259 (N_7259,N_3670,N_4663);
nand U7260 (N_7260,N_4421,N_4943);
nor U7261 (N_7261,N_3555,N_4855);
xor U7262 (N_7262,N_3644,N_2515);
nand U7263 (N_7263,N_4452,N_4443);
nand U7264 (N_7264,N_4141,N_3377);
and U7265 (N_7265,N_3282,N_4969);
and U7266 (N_7266,N_3245,N_3910);
nor U7267 (N_7267,N_4926,N_2813);
and U7268 (N_7268,N_4211,N_4731);
xor U7269 (N_7269,N_4412,N_2622);
nor U7270 (N_7270,N_4706,N_4258);
and U7271 (N_7271,N_3220,N_4171);
nand U7272 (N_7272,N_4437,N_4093);
and U7273 (N_7273,N_4816,N_3940);
and U7274 (N_7274,N_4801,N_4345);
nand U7275 (N_7275,N_4737,N_3340);
or U7276 (N_7276,N_3264,N_2898);
nand U7277 (N_7277,N_3091,N_3156);
nand U7278 (N_7278,N_4178,N_4621);
nand U7279 (N_7279,N_4564,N_3794);
nand U7280 (N_7280,N_3916,N_4448);
or U7281 (N_7281,N_4321,N_2842);
and U7282 (N_7282,N_3106,N_3338);
or U7283 (N_7283,N_4787,N_4032);
nor U7284 (N_7284,N_3671,N_4857);
xnor U7285 (N_7285,N_2681,N_4709);
xor U7286 (N_7286,N_3125,N_3588);
nand U7287 (N_7287,N_3124,N_4402);
nand U7288 (N_7288,N_4758,N_3006);
nor U7289 (N_7289,N_3905,N_2681);
nor U7290 (N_7290,N_3853,N_2873);
nor U7291 (N_7291,N_4086,N_2647);
or U7292 (N_7292,N_2571,N_3741);
nor U7293 (N_7293,N_4972,N_3701);
or U7294 (N_7294,N_2623,N_4014);
nor U7295 (N_7295,N_4356,N_4722);
and U7296 (N_7296,N_4543,N_3840);
or U7297 (N_7297,N_3999,N_3566);
and U7298 (N_7298,N_3079,N_4982);
or U7299 (N_7299,N_2665,N_4127);
and U7300 (N_7300,N_3760,N_3507);
nor U7301 (N_7301,N_3119,N_3075);
nor U7302 (N_7302,N_4438,N_4005);
and U7303 (N_7303,N_4208,N_3256);
xor U7304 (N_7304,N_4670,N_3697);
or U7305 (N_7305,N_4176,N_3483);
xor U7306 (N_7306,N_4667,N_2966);
nand U7307 (N_7307,N_4718,N_4305);
nor U7308 (N_7308,N_3007,N_4177);
xor U7309 (N_7309,N_3304,N_4552);
or U7310 (N_7310,N_2918,N_4799);
nand U7311 (N_7311,N_3541,N_4855);
nor U7312 (N_7312,N_2585,N_4639);
xor U7313 (N_7313,N_4651,N_4745);
nor U7314 (N_7314,N_4333,N_3229);
nand U7315 (N_7315,N_4983,N_3523);
or U7316 (N_7316,N_4306,N_3044);
xor U7317 (N_7317,N_3953,N_2599);
and U7318 (N_7318,N_3210,N_2657);
nand U7319 (N_7319,N_4297,N_3781);
nor U7320 (N_7320,N_2889,N_3006);
nand U7321 (N_7321,N_3691,N_4964);
nand U7322 (N_7322,N_4395,N_2811);
nand U7323 (N_7323,N_3766,N_4006);
or U7324 (N_7324,N_3947,N_4081);
nand U7325 (N_7325,N_2586,N_3230);
nand U7326 (N_7326,N_4340,N_3380);
or U7327 (N_7327,N_4871,N_3460);
and U7328 (N_7328,N_4911,N_2624);
and U7329 (N_7329,N_4388,N_4345);
nor U7330 (N_7330,N_4798,N_3089);
nand U7331 (N_7331,N_2885,N_4937);
nand U7332 (N_7332,N_3824,N_2716);
nand U7333 (N_7333,N_4848,N_3297);
or U7334 (N_7334,N_3265,N_3458);
and U7335 (N_7335,N_4203,N_3861);
xor U7336 (N_7336,N_4311,N_3109);
and U7337 (N_7337,N_4122,N_4645);
or U7338 (N_7338,N_3656,N_4244);
or U7339 (N_7339,N_3786,N_4001);
and U7340 (N_7340,N_2956,N_4882);
and U7341 (N_7341,N_3969,N_3482);
nor U7342 (N_7342,N_3641,N_2637);
nor U7343 (N_7343,N_2815,N_3728);
nor U7344 (N_7344,N_2558,N_3671);
or U7345 (N_7345,N_3924,N_3502);
nand U7346 (N_7346,N_3100,N_4099);
or U7347 (N_7347,N_2701,N_2972);
nor U7348 (N_7348,N_3306,N_4060);
nand U7349 (N_7349,N_4728,N_3854);
nor U7350 (N_7350,N_3624,N_4096);
and U7351 (N_7351,N_3856,N_2712);
nor U7352 (N_7352,N_4148,N_2688);
xnor U7353 (N_7353,N_2578,N_4502);
or U7354 (N_7354,N_3541,N_3962);
nor U7355 (N_7355,N_3678,N_4652);
xnor U7356 (N_7356,N_2639,N_3801);
nor U7357 (N_7357,N_4536,N_3491);
nor U7358 (N_7358,N_3334,N_4980);
nand U7359 (N_7359,N_4374,N_2546);
nor U7360 (N_7360,N_4358,N_3683);
nor U7361 (N_7361,N_2697,N_3471);
and U7362 (N_7362,N_3858,N_4081);
or U7363 (N_7363,N_3926,N_3663);
nor U7364 (N_7364,N_4817,N_2523);
or U7365 (N_7365,N_3781,N_2547);
and U7366 (N_7366,N_4987,N_4761);
nor U7367 (N_7367,N_2735,N_3290);
or U7368 (N_7368,N_4018,N_4413);
or U7369 (N_7369,N_4125,N_3996);
or U7370 (N_7370,N_3724,N_4843);
nor U7371 (N_7371,N_2500,N_3952);
or U7372 (N_7372,N_4786,N_3756);
and U7373 (N_7373,N_3616,N_3539);
xor U7374 (N_7374,N_4032,N_4472);
nor U7375 (N_7375,N_3820,N_4142);
nand U7376 (N_7376,N_3078,N_3777);
and U7377 (N_7377,N_3203,N_4030);
nor U7378 (N_7378,N_4652,N_4666);
or U7379 (N_7379,N_4743,N_4344);
nor U7380 (N_7380,N_3070,N_3759);
xor U7381 (N_7381,N_3301,N_3549);
nand U7382 (N_7382,N_3755,N_3023);
nor U7383 (N_7383,N_4652,N_2685);
xor U7384 (N_7384,N_3910,N_2564);
and U7385 (N_7385,N_3316,N_2962);
or U7386 (N_7386,N_4619,N_3416);
and U7387 (N_7387,N_4756,N_4409);
or U7388 (N_7388,N_2797,N_2612);
nand U7389 (N_7389,N_4602,N_4834);
and U7390 (N_7390,N_2529,N_3179);
nand U7391 (N_7391,N_3728,N_4502);
nor U7392 (N_7392,N_4865,N_2537);
or U7393 (N_7393,N_2845,N_3388);
or U7394 (N_7394,N_2991,N_4939);
xnor U7395 (N_7395,N_3521,N_3969);
nand U7396 (N_7396,N_4013,N_3877);
nand U7397 (N_7397,N_3694,N_4638);
and U7398 (N_7398,N_3378,N_4178);
nand U7399 (N_7399,N_4948,N_4942);
nand U7400 (N_7400,N_3737,N_4772);
xor U7401 (N_7401,N_3789,N_3172);
nor U7402 (N_7402,N_3935,N_3333);
xor U7403 (N_7403,N_4838,N_3200);
nor U7404 (N_7404,N_3575,N_3960);
nand U7405 (N_7405,N_4669,N_4030);
and U7406 (N_7406,N_3165,N_3915);
nor U7407 (N_7407,N_4093,N_3034);
nand U7408 (N_7408,N_3585,N_3094);
nor U7409 (N_7409,N_3261,N_4235);
nand U7410 (N_7410,N_3175,N_3982);
or U7411 (N_7411,N_4096,N_3074);
or U7412 (N_7412,N_3116,N_4330);
nor U7413 (N_7413,N_4509,N_4004);
and U7414 (N_7414,N_3676,N_3500);
nor U7415 (N_7415,N_4799,N_4388);
nor U7416 (N_7416,N_4340,N_4298);
and U7417 (N_7417,N_4314,N_4109);
nor U7418 (N_7418,N_4246,N_4563);
nand U7419 (N_7419,N_4038,N_4758);
nand U7420 (N_7420,N_3615,N_3706);
nor U7421 (N_7421,N_3050,N_4170);
nor U7422 (N_7422,N_3310,N_4527);
and U7423 (N_7423,N_3406,N_4552);
nand U7424 (N_7424,N_4687,N_2620);
nand U7425 (N_7425,N_3431,N_2833);
and U7426 (N_7426,N_2709,N_2728);
nor U7427 (N_7427,N_4193,N_4020);
or U7428 (N_7428,N_4015,N_2852);
nor U7429 (N_7429,N_3117,N_4611);
nor U7430 (N_7430,N_3676,N_3790);
or U7431 (N_7431,N_2909,N_4263);
nor U7432 (N_7432,N_3441,N_3650);
nand U7433 (N_7433,N_4501,N_3671);
and U7434 (N_7434,N_2566,N_2753);
xnor U7435 (N_7435,N_3193,N_3679);
nand U7436 (N_7436,N_4754,N_4650);
nand U7437 (N_7437,N_4366,N_4572);
nor U7438 (N_7438,N_2835,N_3256);
xor U7439 (N_7439,N_4972,N_3031);
and U7440 (N_7440,N_3115,N_4021);
nor U7441 (N_7441,N_3513,N_2831);
or U7442 (N_7442,N_3141,N_3436);
nand U7443 (N_7443,N_3568,N_2961);
and U7444 (N_7444,N_2836,N_4371);
nor U7445 (N_7445,N_2556,N_4574);
or U7446 (N_7446,N_2947,N_3702);
or U7447 (N_7447,N_3787,N_3618);
nor U7448 (N_7448,N_4182,N_4346);
and U7449 (N_7449,N_3323,N_2949);
nand U7450 (N_7450,N_3251,N_4271);
xor U7451 (N_7451,N_4488,N_3275);
nand U7452 (N_7452,N_3662,N_3797);
and U7453 (N_7453,N_4176,N_4241);
nand U7454 (N_7454,N_4990,N_3514);
and U7455 (N_7455,N_3925,N_3641);
xnor U7456 (N_7456,N_2987,N_3206);
and U7457 (N_7457,N_3197,N_2735);
xnor U7458 (N_7458,N_3841,N_2547);
and U7459 (N_7459,N_3109,N_3093);
nor U7460 (N_7460,N_4793,N_3421);
and U7461 (N_7461,N_4376,N_4228);
nor U7462 (N_7462,N_4989,N_3289);
nor U7463 (N_7463,N_4257,N_3171);
nand U7464 (N_7464,N_4756,N_2912);
nand U7465 (N_7465,N_3074,N_4645);
or U7466 (N_7466,N_2773,N_4524);
or U7467 (N_7467,N_2811,N_4651);
nand U7468 (N_7468,N_2893,N_3817);
and U7469 (N_7469,N_4440,N_4101);
and U7470 (N_7470,N_4588,N_3622);
nand U7471 (N_7471,N_2704,N_3315);
xor U7472 (N_7472,N_2671,N_3898);
xor U7473 (N_7473,N_3593,N_3113);
nand U7474 (N_7474,N_2955,N_4095);
and U7475 (N_7475,N_2736,N_4800);
nor U7476 (N_7476,N_3171,N_4218);
xor U7477 (N_7477,N_3280,N_3938);
xor U7478 (N_7478,N_3544,N_4457);
or U7479 (N_7479,N_4549,N_3028);
nand U7480 (N_7480,N_2849,N_3549);
nand U7481 (N_7481,N_3338,N_3281);
and U7482 (N_7482,N_2630,N_3438);
and U7483 (N_7483,N_4680,N_4124);
or U7484 (N_7484,N_4894,N_3032);
nand U7485 (N_7485,N_2801,N_4364);
nand U7486 (N_7486,N_2683,N_4935);
xnor U7487 (N_7487,N_4470,N_3560);
nor U7488 (N_7488,N_3936,N_4058);
nand U7489 (N_7489,N_4979,N_2753);
nor U7490 (N_7490,N_3065,N_2555);
nand U7491 (N_7491,N_4840,N_4455);
xnor U7492 (N_7492,N_3480,N_3777);
nor U7493 (N_7493,N_4307,N_3756);
and U7494 (N_7494,N_4941,N_3431);
or U7495 (N_7495,N_3616,N_3620);
nor U7496 (N_7496,N_3723,N_3062);
and U7497 (N_7497,N_4524,N_3044);
and U7498 (N_7498,N_2824,N_4381);
nor U7499 (N_7499,N_4917,N_4425);
nor U7500 (N_7500,N_7357,N_5578);
or U7501 (N_7501,N_6173,N_5735);
or U7502 (N_7502,N_6825,N_6777);
nand U7503 (N_7503,N_5413,N_7122);
nand U7504 (N_7504,N_6548,N_5652);
nor U7505 (N_7505,N_7178,N_6263);
or U7506 (N_7506,N_6215,N_7024);
and U7507 (N_7507,N_6086,N_7318);
nor U7508 (N_7508,N_6708,N_7190);
or U7509 (N_7509,N_6151,N_6061);
and U7510 (N_7510,N_5936,N_6671);
nand U7511 (N_7511,N_6901,N_7220);
nand U7512 (N_7512,N_7197,N_6774);
or U7513 (N_7513,N_7141,N_5016);
nand U7514 (N_7514,N_6821,N_6762);
xnor U7515 (N_7515,N_5873,N_7235);
or U7516 (N_7516,N_6957,N_5497);
nor U7517 (N_7517,N_5834,N_7078);
and U7518 (N_7518,N_5668,N_6141);
or U7519 (N_7519,N_5988,N_5934);
or U7520 (N_7520,N_6233,N_6104);
and U7521 (N_7521,N_5386,N_5704);
nand U7522 (N_7522,N_6315,N_5822);
and U7523 (N_7523,N_6601,N_6186);
or U7524 (N_7524,N_6721,N_6359);
xor U7525 (N_7525,N_6341,N_5629);
xnor U7526 (N_7526,N_7345,N_6972);
or U7527 (N_7527,N_5533,N_6660);
xnor U7528 (N_7528,N_7031,N_5498);
nor U7529 (N_7529,N_6096,N_7027);
nor U7530 (N_7530,N_5898,N_7300);
nor U7531 (N_7531,N_5775,N_5681);
nor U7532 (N_7532,N_7095,N_5983);
and U7533 (N_7533,N_6227,N_6007);
or U7534 (N_7534,N_6192,N_5452);
or U7535 (N_7535,N_5846,N_5731);
nor U7536 (N_7536,N_6140,N_6406);
xor U7537 (N_7537,N_6254,N_6318);
nand U7538 (N_7538,N_5955,N_5601);
xor U7539 (N_7539,N_6996,N_6164);
nand U7540 (N_7540,N_5277,N_6154);
nor U7541 (N_7541,N_7407,N_5012);
xor U7542 (N_7542,N_6223,N_5338);
and U7543 (N_7543,N_7090,N_5826);
nor U7544 (N_7544,N_5930,N_7081);
nand U7545 (N_7545,N_7030,N_7114);
or U7546 (N_7546,N_5303,N_7194);
nor U7547 (N_7547,N_7209,N_6260);
or U7548 (N_7548,N_6745,N_6685);
nand U7549 (N_7549,N_5737,N_6894);
or U7550 (N_7550,N_6617,N_7364);
and U7551 (N_7551,N_6329,N_7173);
nor U7552 (N_7552,N_6010,N_5758);
xnor U7553 (N_7553,N_6541,N_6313);
or U7554 (N_7554,N_5700,N_5763);
and U7555 (N_7555,N_7453,N_6103);
and U7556 (N_7556,N_6664,N_7098);
and U7557 (N_7557,N_6609,N_7032);
nand U7558 (N_7558,N_6792,N_5496);
nand U7559 (N_7559,N_7283,N_6966);
or U7560 (N_7560,N_7377,N_6564);
nand U7561 (N_7561,N_6712,N_7099);
nor U7562 (N_7562,N_5744,N_5856);
xnor U7563 (N_7563,N_7189,N_5573);
or U7564 (N_7564,N_6064,N_5053);
nand U7565 (N_7565,N_5669,N_5109);
or U7566 (N_7566,N_7390,N_6780);
and U7567 (N_7567,N_6177,N_6603);
nor U7568 (N_7568,N_5257,N_5130);
nor U7569 (N_7569,N_7076,N_5490);
nor U7570 (N_7570,N_7080,N_5858);
xnor U7571 (N_7571,N_6445,N_5305);
xnor U7572 (N_7572,N_5371,N_6420);
or U7573 (N_7573,N_5990,N_6840);
or U7574 (N_7574,N_6955,N_6931);
nor U7575 (N_7575,N_6039,N_6448);
nor U7576 (N_7576,N_5029,N_5952);
xnor U7577 (N_7577,N_5269,N_6421);
nor U7578 (N_7578,N_6596,N_6057);
nand U7579 (N_7579,N_6600,N_5807);
and U7580 (N_7580,N_7026,N_5838);
nand U7581 (N_7581,N_5918,N_5508);
and U7582 (N_7582,N_6265,N_7128);
or U7583 (N_7583,N_7199,N_7291);
or U7584 (N_7584,N_5633,N_6816);
and U7585 (N_7585,N_6650,N_7137);
nand U7586 (N_7586,N_7091,N_7191);
and U7587 (N_7587,N_6506,N_6466);
or U7588 (N_7588,N_6314,N_7158);
nand U7589 (N_7589,N_7392,N_7202);
nor U7590 (N_7590,N_7472,N_5294);
and U7591 (N_7591,N_5131,N_6148);
or U7592 (N_7592,N_7142,N_5865);
or U7593 (N_7593,N_5612,N_5541);
nand U7594 (N_7594,N_7496,N_6951);
nor U7595 (N_7595,N_7260,N_5992);
nand U7596 (N_7596,N_6638,N_6826);
nor U7597 (N_7597,N_7337,N_6903);
or U7598 (N_7598,N_5581,N_5556);
nand U7599 (N_7599,N_7008,N_5068);
or U7600 (N_7600,N_7249,N_5026);
xnor U7601 (N_7601,N_5264,N_5719);
and U7602 (N_7602,N_5870,N_5975);
or U7603 (N_7603,N_5032,N_5423);
nor U7604 (N_7604,N_7000,N_6939);
nor U7605 (N_7605,N_7428,N_5558);
nand U7606 (N_7606,N_5977,N_6447);
and U7607 (N_7607,N_5392,N_7421);
or U7608 (N_7608,N_5646,N_7229);
and U7609 (N_7609,N_7304,N_6252);
and U7610 (N_7610,N_6725,N_7490);
xnor U7611 (N_7611,N_5214,N_6839);
nor U7612 (N_7612,N_5575,N_6045);
nor U7613 (N_7613,N_7104,N_6312);
and U7614 (N_7614,N_6942,N_6900);
and U7615 (N_7615,N_5090,N_6538);
xnor U7616 (N_7616,N_5745,N_5583);
or U7617 (N_7617,N_7072,N_5117);
and U7618 (N_7618,N_7383,N_6180);
nor U7619 (N_7619,N_6817,N_6455);
and U7620 (N_7620,N_6077,N_6449);
nand U7621 (N_7621,N_5966,N_6129);
and U7622 (N_7622,N_5343,N_6283);
or U7623 (N_7623,N_5086,N_7074);
and U7624 (N_7624,N_7239,N_5649);
nand U7625 (N_7625,N_5788,N_6153);
or U7626 (N_7626,N_5276,N_7156);
nand U7627 (N_7627,N_6991,N_6733);
and U7628 (N_7628,N_6552,N_5723);
nor U7629 (N_7629,N_7038,N_6851);
or U7630 (N_7630,N_6946,N_6789);
or U7631 (N_7631,N_5429,N_7481);
nand U7632 (N_7632,N_5391,N_5367);
nand U7633 (N_7633,N_5144,N_5805);
or U7634 (N_7634,N_5548,N_6612);
nor U7635 (N_7635,N_6912,N_7361);
xor U7636 (N_7636,N_5076,N_6968);
and U7637 (N_7637,N_5140,N_6847);
xnor U7638 (N_7638,N_6083,N_7398);
and U7639 (N_7639,N_6349,N_5417);
xor U7640 (N_7640,N_7075,N_7084);
or U7641 (N_7641,N_7052,N_5440);
or U7642 (N_7642,N_5804,N_6806);
nor U7643 (N_7643,N_5085,N_5657);
nand U7644 (N_7644,N_6945,N_6531);
and U7645 (N_7645,N_6068,N_7131);
and U7646 (N_7646,N_7323,N_5770);
nand U7647 (N_7647,N_7063,N_5660);
nand U7648 (N_7648,N_5783,N_5639);
or U7649 (N_7649,N_5126,N_5688);
nand U7650 (N_7650,N_6679,N_6749);
or U7651 (N_7651,N_6990,N_5241);
or U7652 (N_7652,N_5613,N_7284);
nor U7653 (N_7653,N_7417,N_5926);
nand U7654 (N_7654,N_6978,N_5041);
nand U7655 (N_7655,N_6843,N_5353);
and U7656 (N_7656,N_5978,N_5526);
nand U7657 (N_7657,N_7376,N_6740);
nand U7658 (N_7658,N_7321,N_5015);
nand U7659 (N_7659,N_7427,N_6624);
and U7660 (N_7660,N_5162,N_6948);
or U7661 (N_7661,N_6094,N_5844);
nor U7662 (N_7662,N_5954,N_6284);
xnor U7663 (N_7663,N_5505,N_5451);
and U7664 (N_7664,N_6386,N_5267);
nand U7665 (N_7665,N_6256,N_6289);
or U7666 (N_7666,N_6493,N_7480);
and U7667 (N_7667,N_7223,N_5079);
nand U7668 (N_7668,N_7044,N_6917);
or U7669 (N_7669,N_5196,N_7314);
xnor U7670 (N_7670,N_5246,N_6275);
and U7671 (N_7671,N_5872,N_7192);
nand U7672 (N_7672,N_5237,N_7255);
and U7673 (N_7673,N_7266,N_6684);
nand U7674 (N_7674,N_6998,N_5519);
or U7675 (N_7675,N_6756,N_5236);
or U7676 (N_7676,N_6979,N_5564);
and U7677 (N_7677,N_5445,N_6428);
and U7678 (N_7678,N_6926,N_6967);
xnor U7679 (N_7679,N_6793,N_5782);
nand U7680 (N_7680,N_6288,N_6222);
nand U7681 (N_7681,N_5538,N_6323);
or U7682 (N_7682,N_5348,N_7441);
and U7683 (N_7683,N_6442,N_6522);
and U7684 (N_7684,N_7251,N_7051);
and U7685 (N_7685,N_7350,N_5081);
xor U7686 (N_7686,N_6909,N_7097);
xor U7687 (N_7687,N_5570,N_5462);
or U7688 (N_7688,N_7048,N_5106);
or U7689 (N_7689,N_6344,N_7134);
nand U7690 (N_7690,N_5841,N_6138);
xor U7691 (N_7691,N_5271,N_5132);
nor U7692 (N_7692,N_5852,N_7014);
and U7693 (N_7693,N_7464,N_5874);
nand U7694 (N_7694,N_7174,N_5024);
nor U7695 (N_7695,N_5774,N_6881);
and U7696 (N_7696,N_7144,N_5861);
and U7697 (N_7697,N_5361,N_6109);
nand U7698 (N_7698,N_6179,N_5395);
nor U7699 (N_7699,N_6079,N_5096);
or U7700 (N_7700,N_5453,N_5714);
and U7701 (N_7701,N_6044,N_6472);
nand U7702 (N_7702,N_5333,N_7019);
nand U7703 (N_7703,N_6408,N_5599);
nor U7704 (N_7704,N_6231,N_6135);
and U7705 (N_7705,N_5280,N_6673);
nor U7706 (N_7706,N_6781,N_6370);
nand U7707 (N_7707,N_7461,N_6120);
nand U7708 (N_7708,N_6719,N_6997);
xnor U7709 (N_7709,N_5000,N_7277);
or U7710 (N_7710,N_5715,N_6869);
and U7711 (N_7711,N_5039,N_5891);
nor U7712 (N_7712,N_5710,N_5998);
or U7713 (N_7713,N_7294,N_6099);
and U7714 (N_7714,N_5040,N_5640);
nor U7715 (N_7715,N_7150,N_5400);
and U7716 (N_7716,N_6499,N_7047);
and U7717 (N_7717,N_6131,N_5849);
and U7718 (N_7718,N_5278,N_6628);
or U7719 (N_7719,N_6433,N_6262);
and U7720 (N_7720,N_5127,N_6102);
nand U7721 (N_7721,N_5717,N_6053);
nand U7722 (N_7722,N_6732,N_6711);
nor U7723 (N_7723,N_5957,N_5212);
nand U7724 (N_7724,N_5254,N_5396);
nand U7725 (N_7725,N_7405,N_6845);
or U7726 (N_7726,N_5410,N_6403);
nand U7727 (N_7727,N_6389,N_6150);
or U7728 (N_7728,N_6454,N_5382);
nor U7729 (N_7729,N_5209,N_6773);
nor U7730 (N_7730,N_6842,N_5919);
or U7731 (N_7731,N_7397,N_5943);
or U7732 (N_7732,N_7272,N_5215);
nor U7733 (N_7733,N_6272,N_5881);
or U7734 (N_7734,N_5565,N_6768);
nand U7735 (N_7735,N_6739,N_7491);
or U7736 (N_7736,N_5671,N_6354);
or U7737 (N_7737,N_5142,N_5240);
nand U7738 (N_7738,N_5065,N_7325);
nor U7739 (N_7739,N_5173,N_5456);
nor U7740 (N_7740,N_6571,N_7415);
and U7741 (N_7741,N_6819,N_6597);
nand U7742 (N_7742,N_6870,N_6006);
nand U7743 (N_7743,N_6385,N_6608);
or U7744 (N_7744,N_6994,N_5562);
xor U7745 (N_7745,N_6735,N_6828);
nor U7746 (N_7746,N_5938,N_5454);
nor U7747 (N_7747,N_6280,N_6623);
nand U7748 (N_7748,N_6297,N_7403);
or U7749 (N_7749,N_5523,N_5547);
and U7750 (N_7750,N_5426,N_7469);
nand U7751 (N_7751,N_7413,N_5634);
xnor U7752 (N_7752,N_5860,N_6703);
or U7753 (N_7753,N_5949,N_7252);
or U7754 (N_7754,N_5535,N_7324);
or U7755 (N_7755,N_5001,N_5568);
and U7756 (N_7756,N_6391,N_6824);
nor U7757 (N_7757,N_5885,N_6090);
and U7758 (N_7758,N_5747,N_5506);
and U7759 (N_7759,N_7382,N_5840);
xnor U7760 (N_7760,N_5370,N_7457);
nor U7761 (N_7761,N_5932,N_7017);
or U7762 (N_7762,N_7149,N_6761);
nand U7763 (N_7763,N_6510,N_5190);
xor U7764 (N_7764,N_6534,N_6074);
nor U7765 (N_7765,N_5686,N_7298);
or U7766 (N_7766,N_5554,N_5513);
and U7767 (N_7767,N_5042,N_5650);
or U7768 (N_7768,N_5195,N_7434);
and U7769 (N_7769,N_7366,N_6490);
nand U7770 (N_7770,N_5302,N_6054);
or U7771 (N_7771,N_6070,N_6904);
and U7772 (N_7772,N_7247,N_6118);
nor U7773 (N_7773,N_6962,N_6518);
xor U7774 (N_7774,N_5584,N_6937);
and U7775 (N_7775,N_6040,N_7475);
nand U7776 (N_7776,N_6143,N_6627);
nand U7777 (N_7777,N_6863,N_6799);
or U7778 (N_7778,N_6091,N_7351);
nor U7779 (N_7779,N_6366,N_5373);
xnor U7780 (N_7780,N_6414,N_5808);
xnor U7781 (N_7781,N_7211,N_6126);
nand U7782 (N_7782,N_5743,N_6521);
and U7783 (N_7783,N_6683,N_7162);
and U7784 (N_7784,N_5438,N_6720);
xor U7785 (N_7785,N_5482,N_6658);
nor U7786 (N_7786,N_6369,N_5569);
nor U7787 (N_7787,N_6633,N_7280);
and U7788 (N_7788,N_5159,N_5110);
nand U7789 (N_7789,N_6033,N_5799);
or U7790 (N_7790,N_6337,N_6834);
and U7791 (N_7791,N_5151,N_5813);
or U7792 (N_7792,N_5848,N_6914);
nor U7793 (N_7793,N_5610,N_6823);
xor U7794 (N_7794,N_5307,N_7391);
or U7795 (N_7795,N_7039,N_6278);
nand U7796 (N_7796,N_7065,N_5384);
or U7797 (N_7797,N_6832,N_5060);
nor U7798 (N_7798,N_7393,N_5468);
and U7799 (N_7799,N_5093,N_5336);
or U7800 (N_7800,N_5285,N_5530);
nand U7801 (N_7801,N_5324,N_5408);
and U7802 (N_7802,N_6100,N_6194);
nor U7803 (N_7803,N_5532,N_6885);
nand U7804 (N_7804,N_5164,N_6417);
or U7805 (N_7805,N_7271,N_6804);
nor U7806 (N_7806,N_6622,N_5958);
and U7807 (N_7807,N_6095,N_6388);
or U7808 (N_7808,N_5457,N_5114);
nor U7809 (N_7809,N_7020,N_6975);
nand U7810 (N_7810,N_7409,N_5796);
nand U7811 (N_7811,N_7400,N_7317);
nor U7812 (N_7812,N_5208,N_5608);
nor U7813 (N_7813,N_7045,N_5136);
nand U7814 (N_7814,N_5851,N_6307);
or U7815 (N_7815,N_6229,N_6050);
or U7816 (N_7816,N_5956,N_6540);
xnor U7817 (N_7817,N_5691,N_7226);
or U7818 (N_7818,N_6444,N_5871);
and U7819 (N_7819,N_6224,N_5542);
nor U7820 (N_7820,N_6663,N_5066);
nor U7821 (N_7821,N_5292,N_7408);
and U7822 (N_7822,N_7328,N_6829);
xnor U7823 (N_7823,N_7136,N_5626);
nand U7824 (N_7824,N_5019,N_5561);
nand U7825 (N_7825,N_6021,N_5328);
and U7826 (N_7826,N_7333,N_5027);
nor U7827 (N_7827,N_6764,N_6782);
or U7828 (N_7828,N_6430,N_6776);
nor U7829 (N_7829,N_6133,N_5446);
nand U7830 (N_7830,N_5033,N_5036);
and U7831 (N_7831,N_5797,N_7116);
nor U7832 (N_7832,N_6020,N_6573);
and U7833 (N_7833,N_5732,N_5928);
nand U7834 (N_7834,N_7015,N_6497);
or U7835 (N_7835,N_5900,N_6360);
or U7836 (N_7836,N_6911,N_6365);
and U7837 (N_7837,N_6182,N_6424);
or U7838 (N_7838,N_5402,N_6013);
or U7839 (N_7839,N_6738,N_5986);
nand U7840 (N_7840,N_7103,N_5916);
nand U7841 (N_7841,N_6983,N_5077);
nand U7842 (N_7842,N_7006,N_6795);
nand U7843 (N_7843,N_6482,N_6471);
or U7844 (N_7844,N_5405,N_5133);
xnor U7845 (N_7845,N_6836,N_5366);
nand U7846 (N_7846,N_6970,N_6729);
and U7847 (N_7847,N_6000,N_6085);
or U7848 (N_7848,N_6432,N_7218);
nand U7849 (N_7849,N_7442,N_5050);
or U7850 (N_7850,N_6766,N_5707);
nand U7851 (N_7851,N_6958,N_6561);
or U7852 (N_7852,N_6483,N_6858);
and U7853 (N_7853,N_5394,N_6121);
xnor U7854 (N_7854,N_5028,N_7499);
and U7855 (N_7855,N_5961,N_6145);
nand U7856 (N_7856,N_5301,N_6038);
xor U7857 (N_7857,N_5101,N_7494);
or U7858 (N_7858,N_6240,N_6770);
xnor U7859 (N_7859,N_6960,N_5166);
nor U7860 (N_7860,N_5622,N_5647);
nand U7861 (N_7861,N_6470,N_6401);
and U7862 (N_7862,N_5518,N_5833);
and U7863 (N_7863,N_7269,N_5697);
nand U7864 (N_7864,N_5663,N_6175);
or U7865 (N_7865,N_7127,N_5178);
and U7866 (N_7866,N_5102,N_6264);
and U7867 (N_7867,N_6328,N_7359);
and U7868 (N_7868,N_7085,N_6755);
nand U7869 (N_7869,N_6977,N_6503);
or U7870 (N_7870,N_5945,N_5537);
nand U7871 (N_7871,N_5135,N_6635);
nand U7872 (N_7872,N_6055,N_6512);
or U7873 (N_7873,N_5730,N_7079);
nor U7874 (N_7874,N_6568,N_6507);
nand U7875 (N_7875,N_5795,N_6481);
nand U7876 (N_7876,N_6460,N_5924);
nand U7877 (N_7877,N_5123,N_6775);
nor U7878 (N_7878,N_5866,N_6362);
or U7879 (N_7879,N_5901,N_6204);
nand U7880 (N_7880,N_6257,N_6744);
nand U7881 (N_7881,N_6043,N_5592);
or U7882 (N_7882,N_5359,N_5013);
and U7883 (N_7883,N_7089,N_6317);
or U7884 (N_7884,N_6202,N_5399);
or U7885 (N_7885,N_6004,N_5062);
xnor U7886 (N_7886,N_6221,N_5205);
and U7887 (N_7887,N_5931,N_6641);
nand U7888 (N_7888,N_5054,N_6759);
and U7889 (N_7889,N_7240,N_7165);
and U7890 (N_7890,N_6950,N_6715);
xnor U7891 (N_7891,N_7320,N_6751);
and U7892 (N_7892,N_6974,N_6463);
xnor U7893 (N_7893,N_5174,N_5722);
or U7894 (N_7894,N_6809,N_6029);
and U7895 (N_7895,N_5820,N_6498);
nand U7896 (N_7896,N_5913,N_6253);
nand U7897 (N_7897,N_5644,N_5487);
nor U7898 (N_7898,N_7021,N_7281);
nand U7899 (N_7899,N_7436,N_5406);
nand U7900 (N_7900,N_5605,N_7492);
xnor U7901 (N_7901,N_5158,N_6107);
and U7902 (N_7902,N_5489,N_5880);
or U7903 (N_7903,N_5607,N_5709);
and U7904 (N_7904,N_6737,N_5520);
and U7905 (N_7905,N_6213,N_6160);
and U7906 (N_7906,N_7055,N_6363);
xnor U7907 (N_7907,N_6785,N_5772);
xor U7908 (N_7908,N_5525,N_5416);
xor U7909 (N_7909,N_6158,N_6191);
or U7910 (N_7910,N_5818,N_5682);
and U7911 (N_7911,N_6290,N_5769);
nor U7912 (N_7912,N_6984,N_6677);
nand U7913 (N_7913,N_6404,N_7381);
nand U7914 (N_7914,N_6963,N_7111);
and U7915 (N_7915,N_6680,N_6211);
nor U7916 (N_7916,N_6206,N_6611);
nor U7917 (N_7917,N_7438,N_5339);
or U7918 (N_7918,N_6450,N_6117);
or U7919 (N_7919,N_6101,N_6333);
nor U7920 (N_7920,N_7347,N_5767);
or U7921 (N_7921,N_6338,N_7456);
nor U7922 (N_7922,N_6525,N_7476);
and U7923 (N_7923,N_5794,N_7447);
and U7924 (N_7924,N_5694,N_5120);
and U7925 (N_7925,N_5198,N_6783);
nand U7926 (N_7926,N_6713,N_5685);
nand U7927 (N_7927,N_5238,N_5281);
xor U7928 (N_7928,N_6168,N_7286);
nand U7929 (N_7929,N_5300,N_7443);
or U7930 (N_7930,N_6921,N_6956);
or U7931 (N_7931,N_6357,N_6487);
or U7932 (N_7932,N_7454,N_6644);
nor U7933 (N_7933,N_6862,N_5229);
nand U7934 (N_7934,N_7430,N_6837);
and U7935 (N_7935,N_6798,N_7278);
nor U7936 (N_7936,N_5058,N_5727);
or U7937 (N_7937,N_5256,N_5604);
nand U7938 (N_7938,N_5527,N_5202);
or U7939 (N_7939,N_5893,N_6698);
or U7940 (N_7940,N_6545,N_5980);
nand U7941 (N_7941,N_6636,N_5511);
and U7942 (N_7942,N_5611,N_6352);
or U7943 (N_7943,N_5441,N_6412);
nand U7944 (N_7944,N_5628,N_6028);
nand U7945 (N_7945,N_6877,N_6249);
nand U7946 (N_7946,N_7452,N_7358);
nor U7947 (N_7947,N_7297,N_6989);
nand U7948 (N_7948,N_5586,N_5232);
or U7949 (N_7949,N_7117,N_5403);
nand U7950 (N_7950,N_5119,N_6875);
nor U7951 (N_7951,N_5552,N_6932);
xnor U7952 (N_7952,N_5470,N_5574);
and U7953 (N_7953,N_6704,N_6281);
nand U7954 (N_7954,N_5398,N_7422);
and U7955 (N_7955,N_7336,N_6155);
or U7956 (N_7956,N_6818,N_5100);
and U7957 (N_7957,N_5486,N_5897);
nor U7958 (N_7958,N_7465,N_5811);
nor U7959 (N_7959,N_5588,N_5326);
nor U7960 (N_7960,N_6582,N_6516);
nand U7961 (N_7961,N_7395,N_5969);
or U7962 (N_7962,N_7151,N_7082);
nor U7963 (N_7963,N_6898,N_5284);
and U7964 (N_7964,N_6724,N_5206);
and U7965 (N_7965,N_6577,N_7205);
xnor U7966 (N_7966,N_6566,N_6508);
or U7967 (N_7967,N_6927,N_6852);
or U7968 (N_7968,N_5156,N_7295);
nand U7969 (N_7969,N_6195,N_5203);
nand U7970 (N_7970,N_6550,N_7228);
or U7971 (N_7971,N_7132,N_5200);
or U7972 (N_7972,N_7375,N_5543);
nand U7973 (N_7973,N_6277,N_5684);
or U7974 (N_7974,N_6859,N_5141);
or U7975 (N_7975,N_7354,N_6648);
or U7976 (N_7976,N_6916,N_6459);
nand U7977 (N_7977,N_6159,N_5516);
xor U7978 (N_7978,N_7148,N_5806);
and U7979 (N_7979,N_6579,N_5389);
and U7980 (N_7980,N_6473,N_5037);
nor U7981 (N_7981,N_5340,N_6981);
nand U7982 (N_7982,N_7301,N_6261);
or U7983 (N_7983,N_6505,N_7402);
and U7984 (N_7984,N_5055,N_5145);
and U7985 (N_7985,N_6119,N_6146);
nand U7986 (N_7986,N_5597,N_5803);
xor U7987 (N_7987,N_7034,N_7374);
nor U7988 (N_7988,N_7265,N_6811);
nand U7989 (N_7989,N_5662,N_6382);
nand U7990 (N_7990,N_6938,N_5869);
and U7991 (N_7991,N_7313,N_6754);
nand U7992 (N_7992,N_7088,N_5344);
nand U7993 (N_7993,N_5828,N_7470);
or U7994 (N_7994,N_7264,N_7025);
or U7995 (N_7995,N_7215,N_6351);
nor U7996 (N_7996,N_6098,N_5658);
and U7997 (N_7997,N_5274,N_5448);
xor U7998 (N_7998,N_5981,N_6504);
or U7999 (N_7999,N_7221,N_6169);
nor U8000 (N_8000,N_6554,N_5404);
xnor U8001 (N_8001,N_6062,N_5252);
nand U8002 (N_8002,N_6092,N_6236);
or U8003 (N_8003,N_7167,N_5545);
xnor U8004 (N_8004,N_7348,N_5331);
and U8005 (N_8005,N_6399,N_5310);
xor U8006 (N_8006,N_7455,N_5721);
nor U8007 (N_8007,N_6426,N_7478);
and U8008 (N_8008,N_5920,N_5968);
nor U8009 (N_8009,N_5350,N_5754);
or U8010 (N_8010,N_7468,N_5982);
and U8011 (N_8011,N_7367,N_7384);
nand U8012 (N_8012,N_6198,N_6319);
or U8013 (N_8013,N_6659,N_5887);
nand U8014 (N_8014,N_7035,N_5847);
nor U8015 (N_8015,N_5593,N_6619);
xnor U8016 (N_8016,N_7179,N_7061);
nor U8017 (N_8017,N_6743,N_6947);
or U8018 (N_8018,N_5149,N_6849);
or U8019 (N_8019,N_5606,N_5810);
nand U8020 (N_8020,N_5247,N_7483);
nor U8021 (N_8021,N_7003,N_6187);
nand U8022 (N_8022,N_6702,N_5876);
nor U8023 (N_8023,N_6855,N_5666);
and U8024 (N_8024,N_5903,N_6496);
nand U8025 (N_8025,N_5046,N_6392);
and U8026 (N_8026,N_5509,N_5177);
and U8027 (N_8027,N_6985,N_6431);
nand U8028 (N_8028,N_5948,N_6614);
and U8029 (N_8029,N_6864,N_5699);
nor U8030 (N_8030,N_6590,N_5749);
and U8031 (N_8031,N_7203,N_6896);
or U8032 (N_8032,N_6411,N_5321);
nand U8033 (N_8033,N_6791,N_6714);
or U8034 (N_8034,N_5021,N_5253);
nand U8035 (N_8035,N_5069,N_7037);
nor U8036 (N_8036,N_5143,N_5314);
nand U8037 (N_8037,N_5034,N_5430);
and U8038 (N_8038,N_6396,N_5003);
nor U8039 (N_8039,N_6669,N_5375);
and U8040 (N_8040,N_6815,N_7273);
xnor U8041 (N_8041,N_6779,N_5939);
nor U8042 (N_8042,N_5007,N_5244);
nor U8043 (N_8043,N_5676,N_6796);
and U8044 (N_8044,N_6457,N_6181);
or U8045 (N_8045,N_5995,N_5989);
or U8046 (N_8046,N_6670,N_7412);
nand U8047 (N_8047,N_6913,N_5892);
nor U8048 (N_8048,N_6405,N_5741);
or U8049 (N_8049,N_5155,N_6434);
or U8050 (N_8050,N_7204,N_5207);
and U8051 (N_8051,N_7498,N_6316);
or U8052 (N_8052,N_5465,N_5474);
nand U8053 (N_8053,N_7231,N_7423);
or U8054 (N_8054,N_5631,N_6572);
and U8055 (N_8055,N_7440,N_5337);
xor U8056 (N_8056,N_5376,N_6695);
or U8057 (N_8057,N_5967,N_5125);
nand U8058 (N_8058,N_5167,N_5687);
nor U8059 (N_8059,N_5473,N_6273);
or U8060 (N_8060,N_5619,N_6170);
xor U8061 (N_8061,N_6928,N_6258);
nand U8062 (N_8062,N_5814,N_5842);
xnor U8063 (N_8063,N_6458,N_5170);
or U8064 (N_8064,N_5351,N_7410);
and U8065 (N_8065,N_5553,N_6621);
nor U8066 (N_8066,N_5354,N_6848);
or U8067 (N_8067,N_6286,N_6515);
and U8068 (N_8068,N_6034,N_6872);
and U8069 (N_8069,N_7296,N_6152);
xor U8070 (N_8070,N_6124,N_6585);
or U8071 (N_8071,N_6694,N_5827);
and U8072 (N_8072,N_5579,N_7257);
or U8073 (N_8073,N_6524,N_6246);
nor U8074 (N_8074,N_6557,N_6747);
and U8075 (N_8075,N_6347,N_6539);
nor U8076 (N_8076,N_6395,N_5134);
and U8077 (N_8077,N_6478,N_7334);
nand U8078 (N_8078,N_7282,N_6439);
nand U8079 (N_8079,N_7289,N_5225);
nand U8080 (N_8080,N_6452,N_5725);
nor U8081 (N_8081,N_6583,N_7309);
nor U8082 (N_8082,N_6285,N_6185);
nand U8083 (N_8083,N_6924,N_6248);
nand U8084 (N_8084,N_5759,N_6477);
nand U8085 (N_8085,N_7344,N_5449);
and U8086 (N_8086,N_7096,N_5194);
and U8087 (N_8087,N_5638,N_7355);
nor U8088 (N_8088,N_6551,N_7049);
nand U8089 (N_8089,N_7279,N_5680);
nand U8090 (N_8090,N_5309,N_6212);
or U8091 (N_8091,N_6108,N_5695);
and U8092 (N_8092,N_6024,N_5025);
and U8093 (N_8093,N_5008,N_7473);
and U8094 (N_8094,N_7346,N_7054);
or U8095 (N_8095,N_7100,N_7426);
nor U8096 (N_8096,N_6610,N_6188);
xor U8097 (N_8097,N_7138,N_6736);
and U8098 (N_8098,N_6309,N_6345);
nand U8099 (N_8099,N_7371,N_6905);
nor U8100 (N_8100,N_6906,N_5341);
nand U8101 (N_8101,N_5854,N_7356);
or U8102 (N_8102,N_5491,N_6165);
nor U8103 (N_8103,N_6861,N_5780);
nor U8104 (N_8104,N_5661,N_6607);
or U8105 (N_8105,N_5139,N_6933);
nand U8106 (N_8106,N_5625,N_7449);
nor U8107 (N_8107,N_7331,N_5996);
and U8108 (N_8108,N_5286,N_5724);
or U8109 (N_8109,N_7130,N_7372);
nor U8110 (N_8110,N_5539,N_6892);
nand U8111 (N_8111,N_6226,N_6718);
nor U8112 (N_8112,N_6331,N_6130);
nor U8113 (N_8113,N_6731,N_7467);
and U8114 (N_8114,N_7224,N_6003);
nor U8115 (N_8115,N_6210,N_6325);
or U8116 (N_8116,N_5922,N_6786);
nand U8117 (N_8117,N_5227,N_6063);
nor U8118 (N_8118,N_5674,N_7246);
xor U8119 (N_8119,N_7460,N_7254);
nand U8120 (N_8120,N_6778,N_5129);
or U8121 (N_8121,N_5412,N_6001);
nor U8122 (N_8122,N_5507,N_6270);
and U8123 (N_8123,N_5180,N_5418);
and U8124 (N_8124,N_6476,N_5004);
and U8125 (N_8125,N_6041,N_6655);
xor U8126 (N_8126,N_5192,N_6709);
and U8127 (N_8127,N_6139,N_6758);
nand U8128 (N_8128,N_7486,N_6513);
nor U8129 (N_8129,N_6699,N_7484);
xnor U8130 (N_8130,N_5884,N_6820);
and U8131 (N_8131,N_7145,N_5911);
and U8132 (N_8132,N_6479,N_5843);
nor U8133 (N_8133,N_6009,N_6769);
nand U8134 (N_8134,N_6536,N_6046);
xor U8135 (N_8135,N_5250,N_5991);
or U8136 (N_8136,N_5984,N_7338);
and U8137 (N_8137,N_5559,N_5381);
and U8138 (N_8138,N_7115,N_5461);
nor U8139 (N_8139,N_6511,N_5999);
nor U8140 (N_8140,N_5739,N_6813);
nand U8141 (N_8141,N_5970,N_6653);
nand U8142 (N_8142,N_6115,N_5550);
nor U8143 (N_8143,N_5283,N_5540);
or U8144 (N_8144,N_5414,N_5216);
or U8145 (N_8145,N_5057,N_5478);
nor U8146 (N_8146,N_5346,N_6569);
and U8147 (N_8147,N_6008,N_6184);
nor U8148 (N_8148,N_5809,N_7083);
nor U8149 (N_8149,N_5693,N_5484);
or U8150 (N_8150,N_5378,N_5768);
and U8151 (N_8151,N_5435,N_6348);
or U8152 (N_8152,N_6995,N_5994);
and U8153 (N_8153,N_5659,N_5641);
nand U8154 (N_8154,N_5362,N_6056);
and U8155 (N_8155,N_6075,N_5312);
xor U8156 (N_8156,N_6532,N_5083);
or U8157 (N_8157,N_6017,N_6048);
nand U8158 (N_8158,N_5667,N_7005);
nor U8159 (N_8159,N_7029,N_5544);
nand U8160 (N_8160,N_6805,N_6543);
nor U8161 (N_8161,N_7379,N_7140);
nand U8162 (N_8162,N_7157,N_6378);
nor U8163 (N_8163,N_7168,N_6682);
nand U8164 (N_8164,N_5510,N_7175);
nand U8165 (N_8165,N_5757,N_6298);
nor U8166 (N_8166,N_6646,N_5315);
and U8167 (N_8167,N_5228,N_5904);
and U8168 (N_8168,N_7155,N_6080);
and U8169 (N_8169,N_7216,N_6292);
and U8170 (N_8170,N_7013,N_6005);
nand U8171 (N_8171,N_5740,N_5380);
and U8172 (N_8172,N_7068,N_5425);
nor U8173 (N_8173,N_5587,N_6446);
xor U8174 (N_8174,N_7010,N_6690);
or U8175 (N_8175,N_6822,N_5655);
nor U8176 (N_8176,N_6376,N_7164);
and U8177 (N_8177,N_5293,N_5492);
or U8178 (N_8178,N_5450,N_6961);
and U8179 (N_8179,N_6178,N_6250);
and U8180 (N_8180,N_7066,N_5014);
or U8181 (N_8181,N_6716,N_6196);
nor U8182 (N_8182,N_5690,N_6423);
or U8183 (N_8183,N_6752,N_7077);
or U8184 (N_8184,N_6943,N_6067);
or U8185 (N_8185,N_6311,N_6850);
and U8186 (N_8186,N_6689,N_7471);
and U8187 (N_8187,N_6697,N_5829);
or U8188 (N_8188,N_5352,N_7352);
nor U8189 (N_8189,N_5706,N_6189);
and U8190 (N_8190,N_5355,N_6419);
or U8191 (N_8191,N_5878,N_5793);
xor U8192 (N_8192,N_6110,N_5387);
nand U8193 (N_8193,N_6241,N_5460);
nand U8194 (N_8194,N_5635,N_6372);
xnor U8195 (N_8195,N_6576,N_5147);
nand U8196 (N_8196,N_7234,N_5557);
or U8197 (N_8197,N_6052,N_6626);
or U8198 (N_8198,N_5643,N_6171);
nor U8199 (N_8199,N_6701,N_6047);
nor U8200 (N_8200,N_6830,N_7479);
and U8201 (N_8201,N_5422,N_7394);
and U8202 (N_8202,N_6897,N_6023);
or U8203 (N_8203,N_5317,N_6320);
and U8204 (N_8204,N_5153,N_5464);
and U8205 (N_8205,N_7250,N_6375);
nor U8206 (N_8206,N_5193,N_5729);
or U8207 (N_8207,N_5488,N_6666);
nor U8208 (N_8208,N_6353,N_7237);
nor U8209 (N_8209,N_5500,N_6305);
nand U8210 (N_8210,N_6436,N_5219);
nor U8211 (N_8211,N_5411,N_5673);
or U8212 (N_8212,N_5617,N_6865);
xor U8213 (N_8213,N_5620,N_7056);
xnor U8214 (N_8214,N_7267,N_7120);
nand U8215 (N_8215,N_5211,N_6243);
nor U8216 (N_8216,N_6529,N_7060);
nor U8217 (N_8217,N_6765,N_6734);
nand U8218 (N_8218,N_5572,N_7485);
and U8219 (N_8219,N_7482,N_7343);
nand U8220 (N_8220,N_5297,N_5678);
nand U8221 (N_8221,N_7439,N_5974);
nand U8222 (N_8222,N_6604,N_6889);
and U8223 (N_8223,N_6553,N_6071);
nor U8224 (N_8224,N_5296,N_6944);
xnor U8225 (N_8225,N_6592,N_5927);
or U8226 (N_8226,N_7433,N_5789);
nand U8227 (N_8227,N_5882,N_5917);
nand U8228 (N_8228,N_5480,N_5845);
or U8229 (N_8229,N_5602,N_5349);
nand U8230 (N_8230,N_5325,N_7125);
nand U8231 (N_8231,N_6334,N_6220);
xnor U8232 (N_8232,N_7488,N_6549);
nor U8233 (N_8233,N_5197,N_5061);
or U8234 (N_8234,N_5976,N_5689);
and U8235 (N_8235,N_5273,N_6802);
nor U8236 (N_8236,N_7123,N_7106);
and U8237 (N_8237,N_6302,N_5191);
or U8238 (N_8238,N_5536,N_5105);
and U8239 (N_8239,N_7193,N_6501);
xor U8240 (N_8240,N_5591,N_6574);
nand U8241 (N_8241,N_6330,N_6570);
nor U8242 (N_8242,N_7270,N_5172);
nand U8243 (N_8243,N_5726,N_5698);
nor U8244 (N_8244,N_7414,N_6595);
or U8245 (N_8245,N_5683,N_5204);
nand U8246 (N_8246,N_5035,N_5585);
or U8247 (N_8247,N_5363,N_6072);
or U8248 (N_8248,N_5692,N_6546);
or U8249 (N_8249,N_5475,N_5360);
nand U8250 (N_8250,N_6502,N_5942);
nand U8251 (N_8251,N_6287,N_5765);
and U8252 (N_8252,N_7368,N_5836);
and U8253 (N_8253,N_6727,N_5175);
nand U8254 (N_8254,N_6163,N_5696);
nand U8255 (N_8255,N_6544,N_6559);
and U8256 (N_8256,N_5899,N_7258);
nand U8257 (N_8257,N_6293,N_6147);
nor U8258 (N_8258,N_5221,N_6973);
or U8259 (N_8259,N_6267,N_5122);
nor U8260 (N_8260,N_6907,N_5862);
nor U8261 (N_8261,N_5103,N_6687);
or U8262 (N_8262,N_5596,N_6925);
and U8263 (N_8263,N_5792,N_7036);
or U8264 (N_8264,N_5358,N_5239);
nand U8265 (N_8265,N_6157,N_7069);
and U8266 (N_8266,N_5746,N_6763);
and U8267 (N_8267,N_7135,N_5108);
or U8268 (N_8268,N_5790,N_5442);
or U8269 (N_8269,N_5374,N_6910);
or U8270 (N_8270,N_6336,N_5260);
or U8271 (N_8271,N_5272,N_6705);
and U8272 (N_8272,N_5761,N_5415);
nor U8273 (N_8273,N_7419,N_6217);
or U8274 (N_8274,N_6190,N_5877);
nor U8275 (N_8275,N_6238,N_5883);
nor U8276 (N_8276,N_6692,N_6486);
nand U8277 (N_8277,N_6980,N_5902);
nand U8278 (N_8278,N_5632,N_6976);
nand U8279 (N_8279,N_6707,N_5379);
nand U8280 (N_8280,N_5437,N_7259);
or U8281 (N_8281,N_6002,N_5388);
and U8282 (N_8282,N_7101,N_5316);
and U8283 (N_8283,N_6717,N_5773);
xnor U8284 (N_8284,N_5030,N_7420);
and U8285 (N_8285,N_5589,N_5063);
nor U8286 (N_8286,N_5905,N_5642);
or U8287 (N_8287,N_5816,N_7139);
or U8288 (N_8288,N_6868,N_7110);
or U8289 (N_8289,N_5169,N_6339);
nor U8290 (N_8290,N_7236,N_6651);
xor U8291 (N_8291,N_5888,N_6200);
nor U8292 (N_8292,N_5049,N_7330);
xor U8293 (N_8293,N_5483,N_5915);
nand U8294 (N_8294,N_5185,N_6025);
nor U8295 (N_8295,N_5347,N_5791);
xor U8296 (N_8296,N_6199,N_5436);
xnor U8297 (N_8297,N_6810,N_5677);
and U8298 (N_8298,N_6833,N_5072);
nor U8299 (N_8299,N_6547,N_5369);
nor U8300 (N_8300,N_6073,N_5289);
nand U8301 (N_8301,N_7362,N_5751);
xor U8302 (N_8302,N_6183,N_6492);
or U8303 (N_8303,N_5466,N_7329);
nor U8304 (N_8304,N_6259,N_6465);
or U8305 (N_8305,N_6234,N_5784);
nor U8306 (N_8306,N_6027,N_7196);
or U8307 (N_8307,N_5424,N_6588);
xor U8308 (N_8308,N_7293,N_5863);
or U8309 (N_8309,N_5393,N_5112);
xor U8310 (N_8310,N_5823,N_5923);
nor U8311 (N_8311,N_5290,N_6686);
nand U8312 (N_8312,N_6381,N_6867);
or U8313 (N_8313,N_5265,N_5567);
nor U8314 (N_8314,N_6533,N_5815);
nor U8315 (N_8315,N_5261,N_5334);
xor U8316 (N_8316,N_6741,N_6880);
xnor U8317 (N_8317,N_6632,N_6631);
nor U8318 (N_8318,N_5637,N_5327);
nor U8319 (N_8319,N_5563,N_5598);
or U8320 (N_8320,N_5009,N_7303);
or U8321 (N_8321,N_6555,N_6014);
and U8322 (N_8322,N_6602,N_5987);
nand U8323 (N_8323,N_6422,N_6676);
nor U8324 (N_8324,N_5670,N_5471);
nand U8325 (N_8325,N_5421,N_6228);
or U8326 (N_8326,N_6332,N_6383);
or U8327 (N_8327,N_6239,N_5258);
nand U8328 (N_8328,N_6485,N_5245);
nor U8329 (N_8329,N_6672,N_6988);
nor U8330 (N_8330,N_7124,N_5043);
and U8331 (N_8331,N_5501,N_5979);
and U8332 (N_8332,N_6484,N_6575);
and U8333 (N_8333,N_5798,N_6594);
or U8334 (N_8334,N_7340,N_6355);
or U8335 (N_8335,N_7243,N_6599);
or U8336 (N_8336,N_6857,N_6437);
and U8337 (N_8337,N_6031,N_6468);
xor U8338 (N_8338,N_6296,N_6992);
nand U8339 (N_8339,N_5266,N_6556);
or U8340 (N_8340,N_5018,N_5047);
and U8341 (N_8341,N_6218,N_6402);
or U8342 (N_8342,N_6652,N_7233);
and U8343 (N_8343,N_6757,N_5182);
or U8344 (N_8344,N_6474,N_6871);
nor U8345 (N_8345,N_5288,N_5184);
or U8346 (N_8346,N_5766,N_6242);
or U8347 (N_8347,N_7353,N_5124);
xnor U8348 (N_8348,N_6598,N_5675);
nand U8349 (N_8349,N_6986,N_5906);
nand U8350 (N_8350,N_6301,N_7105);
nand U8351 (N_8351,N_5113,N_7349);
nand U8352 (N_8352,N_7166,N_5091);
nand U8353 (N_8353,N_7308,N_5529);
or U8354 (N_8354,N_6874,N_5595);
and U8355 (N_8355,N_5534,N_5837);
nor U8356 (N_8356,N_6884,N_7172);
or U8357 (N_8357,N_5472,N_5577);
nand U8358 (N_8358,N_5555,N_7238);
or U8359 (N_8359,N_6321,N_7058);
nand U8360 (N_8360,N_7437,N_7087);
nand U8361 (N_8361,N_5154,N_7497);
nor U8362 (N_8362,N_7424,N_7425);
xnor U8363 (N_8363,N_5210,N_7444);
or U8364 (N_8364,N_7086,N_7133);
nand U8365 (N_8365,N_5299,N_6088);
or U8366 (N_8366,N_5251,N_6380);
or U8367 (N_8367,N_7171,N_5867);
and U8368 (N_8368,N_7022,N_6886);
nand U8369 (N_8369,N_6954,N_5656);
xnor U8370 (N_8370,N_7380,N_5255);
and U8371 (N_8371,N_7305,N_7225);
nand U8372 (N_8372,N_5270,N_5963);
nand U8373 (N_8373,N_5427,N_7256);
and U8374 (N_8374,N_5051,N_7435);
nor U8375 (N_8375,N_5163,N_7363);
or U8376 (N_8376,N_7302,N_5365);
xor U8377 (N_8377,N_7200,N_5094);
nor U8378 (N_8378,N_6866,N_6642);
nor U8379 (N_8379,N_6019,N_5521);
xnor U8380 (N_8380,N_7458,N_5099);
xnor U8381 (N_8381,N_5875,N_6730);
and U8382 (N_8382,N_6310,N_5010);
nand U8383 (N_8383,N_5679,N_5711);
and U8384 (N_8384,N_6846,N_5821);
and U8385 (N_8385,N_7183,N_6379);
nor U8386 (N_8386,N_7232,N_6675);
or U8387 (N_8387,N_5703,N_5493);
and U8388 (N_8388,N_5912,N_6681);
nor U8389 (N_8389,N_5220,N_5017);
nor U8390 (N_8390,N_7459,N_6398);
xnor U8391 (N_8391,N_6882,N_5636);
xnor U8392 (N_8392,N_5973,N_5104);
or U8393 (N_8393,N_6142,N_5756);
nor U8394 (N_8394,N_7245,N_6410);
nand U8395 (N_8395,N_7418,N_5830);
nor U8396 (N_8396,N_6123,N_7290);
or U8397 (N_8397,N_6443,N_6245);
or U8398 (N_8398,N_7401,N_6902);
nor U8399 (N_8399,N_7004,N_7062);
nor U8400 (N_8400,N_7432,N_5282);
or U8401 (N_8401,N_5006,N_6461);
and U8402 (N_8402,N_5223,N_7041);
nor U8403 (N_8403,N_5779,N_6230);
or U8404 (N_8404,N_7495,N_5896);
and U8405 (N_8405,N_7059,N_6367);
and U8406 (N_8406,N_5005,N_7208);
xnor U8407 (N_8407,N_7207,N_5023);
or U8408 (N_8408,N_5098,N_6049);
or U8409 (N_8409,N_6526,N_5268);
or U8410 (N_8410,N_5073,N_5070);
nand U8411 (N_8411,N_6581,N_6373);
nand U8412 (N_8412,N_6668,N_6409);
or U8413 (N_8413,N_5095,N_5752);
nor U8414 (N_8414,N_6606,N_6371);
nand U8415 (N_8415,N_5409,N_7185);
or U8416 (N_8416,N_5665,N_5432);
and U8417 (N_8417,N_6418,N_5263);
nor U8418 (N_8418,N_5582,N_6327);
xor U8419 (N_8419,N_6887,N_5097);
nand U8420 (N_8420,N_7493,N_5224);
nor U8421 (N_8421,N_5121,N_6772);
and U8422 (N_8422,N_5420,N_5189);
and U8423 (N_8423,N_6657,N_5528);
nor U8424 (N_8424,N_7248,N_7431);
or U8425 (N_8425,N_7386,N_7143);
and U8426 (N_8426,N_6578,N_7180);
xnor U8427 (N_8427,N_5653,N_5469);
and U8428 (N_8428,N_5020,N_6368);
xnor U8429 (N_8429,N_6279,N_6374);
and U8430 (N_8430,N_6613,N_5549);
nand U8431 (N_8431,N_5243,N_6959);
and U8432 (N_8432,N_6794,N_6134);
or U8433 (N_8433,N_5786,N_5455);
or U8434 (N_8434,N_6808,N_7108);
or U8435 (N_8435,N_6161,N_5614);
nand U8436 (N_8436,N_5868,N_6841);
and U8437 (N_8437,N_6207,N_6356);
and U8438 (N_8438,N_5953,N_6214);
nor U8439 (N_8439,N_5812,N_5825);
or U8440 (N_8440,N_6879,N_6084);
nand U8441 (N_8441,N_7399,N_6208);
and U8442 (N_8442,N_6467,N_6271);
nand U8443 (N_8443,N_5304,N_5357);
nand U8444 (N_8444,N_5802,N_7001);
and U8445 (N_8445,N_6105,N_5502);
and U8446 (N_8446,N_6746,N_6728);
nor U8447 (N_8447,N_7152,N_7307);
or U8448 (N_8448,N_6920,N_5323);
nor U8449 (N_8449,N_5431,N_5929);
nor U8450 (N_8450,N_5933,N_5801);
or U8451 (N_8451,N_6197,N_5839);
nor U8452 (N_8452,N_5546,N_6137);
xnor U8453 (N_8453,N_5907,N_5148);
or U8454 (N_8454,N_7227,N_6475);
or U8455 (N_8455,N_6587,N_5311);
and U8456 (N_8456,N_7446,N_5171);
nor U8457 (N_8457,N_6688,N_5495);
nand U8458 (N_8458,N_5044,N_7378);
and U8459 (N_8459,N_6643,N_6742);
and U8460 (N_8460,N_6953,N_7230);
nor U8461 (N_8461,N_7326,N_6814);
and U8462 (N_8462,N_5627,N_5712);
and U8463 (N_8463,N_6647,N_6247);
nor U8464 (N_8464,N_5504,N_5390);
and U8465 (N_8465,N_5962,N_5950);
nor U8466 (N_8466,N_5160,N_7016);
nand U8467 (N_8467,N_5831,N_5576);
and U8468 (N_8468,N_5603,N_7070);
nand U8469 (N_8469,N_7146,N_5045);
nand U8470 (N_8470,N_7261,N_7102);
nor U8471 (N_8471,N_5718,N_6384);
or U8472 (N_8472,N_5082,N_6888);
nand U8473 (N_8473,N_6645,N_5295);
nand U8474 (N_8474,N_5951,N_5781);
nand U8475 (N_8475,N_7170,N_5092);
and U8476 (N_8476,N_5762,N_5499);
nor U8477 (N_8477,N_5459,N_5512);
nor U8478 (N_8478,N_5738,N_6753);
nor U8479 (N_8479,N_7274,N_6637);
xnor U8480 (N_8480,N_6949,N_7445);
or U8481 (N_8481,N_5946,N_6413);
nand U8482 (N_8482,N_6035,N_5235);
xor U8483 (N_8483,N_6930,N_5463);
or U8484 (N_8484,N_6537,N_7241);
or U8485 (N_8485,N_7163,N_5997);
or U8486 (N_8486,N_6873,N_6274);
or U8487 (N_8487,N_6710,N_7332);
or U8488 (N_8488,N_7064,N_5150);
or U8489 (N_8489,N_7214,N_6125);
and U8490 (N_8490,N_6965,N_5397);
nor U8491 (N_8491,N_5494,N_7222);
or U8492 (N_8492,N_7311,N_5372);
and U8493 (N_8493,N_5985,N_7176);
xor U8494 (N_8494,N_6162,N_6069);
xnor U8495 (N_8495,N_6018,N_6844);
and U8496 (N_8496,N_5479,N_7073);
nor U8497 (N_8497,N_6415,N_7287);
or U8498 (N_8498,N_7129,N_5895);
nor U8499 (N_8499,N_5087,N_5183);
nand U8500 (N_8500,N_6042,N_5476);
nor U8501 (N_8501,N_7285,N_5964);
and U8502 (N_8502,N_6377,N_7195);
or U8503 (N_8503,N_5819,N_5778);
xnor U8504 (N_8504,N_7042,N_5080);
xor U8505 (N_8505,N_5879,N_7119);
nand U8506 (N_8506,N_6167,N_5067);
or U8507 (N_8507,N_7023,N_5385);
nor U8508 (N_8508,N_5443,N_6922);
nand U8509 (N_8509,N_5921,N_7043);
nor U8510 (N_8510,N_6335,N_6562);
nor U8511 (N_8511,N_6589,N_5910);
or U8512 (N_8512,N_5089,N_5356);
or U8513 (N_8513,N_6801,N_6722);
and U8514 (N_8514,N_7448,N_6174);
nand U8515 (N_8515,N_5059,N_6156);
and U8516 (N_8516,N_7341,N_5111);
and U8517 (N_8517,N_7147,N_6453);
and U8518 (N_8518,N_5434,N_5908);
or U8519 (N_8519,N_6251,N_5777);
and U8520 (N_8520,N_7206,N_6923);
nand U8521 (N_8521,N_7389,N_7092);
nor U8522 (N_8522,N_6565,N_7160);
or U8523 (N_8523,N_6856,N_5074);
or U8524 (N_8524,N_6971,N_6558);
nand U8525 (N_8525,N_6225,N_5648);
nor U8526 (N_8526,N_5320,N_5600);
xor U8527 (N_8527,N_5377,N_6166);
and U8528 (N_8528,N_5181,N_5318);
nor U8529 (N_8529,N_7385,N_7342);
nand U8530 (N_8530,N_6788,N_5971);
nor U8531 (N_8531,N_5330,N_5708);
nand U8532 (N_8532,N_6488,N_5755);
and U8533 (N_8533,N_7474,N_6235);
nand U8534 (N_8534,N_5419,N_7388);
or U8535 (N_8535,N_5517,N_6416);
and U8536 (N_8536,N_5855,N_5179);
nand U8537 (N_8537,N_6563,N_6082);
nand U8538 (N_8538,N_6520,N_6387);
and U8539 (N_8539,N_5439,N_5234);
nand U8540 (N_8540,N_7373,N_5407);
or U8541 (N_8541,N_6929,N_5313);
xor U8542 (N_8542,N_6269,N_6678);
nand U8543 (N_8543,N_6853,N_5817);
nor U8544 (N_8544,N_5701,N_5894);
and U8545 (N_8545,N_5242,N_6244);
xor U8546 (N_8546,N_5233,N_6803);
nand U8547 (N_8547,N_6831,N_5217);
nor U8548 (N_8548,N_6216,N_6936);
nor U8549 (N_8549,N_7169,N_6219);
or U8550 (N_8550,N_6058,N_5128);
nand U8551 (N_8551,N_5623,N_6517);
or U8552 (N_8552,N_5188,N_5654);
nor U8553 (N_8553,N_6860,N_7370);
or U8554 (N_8554,N_7012,N_6696);
nor U8555 (N_8555,N_7046,N_6066);
or U8556 (N_8556,N_5705,N_7093);
and U8557 (N_8557,N_6771,N_5306);
or U8558 (N_8558,N_7387,N_5993);
nand U8559 (N_8559,N_5853,N_6495);
nor U8560 (N_8560,N_6022,N_5048);
and U8561 (N_8561,N_5477,N_5753);
nand U8562 (N_8562,N_6128,N_6306);
and U8563 (N_8563,N_6918,N_6893);
or U8564 (N_8564,N_6935,N_6790);
and U8565 (N_8565,N_7339,N_6203);
xnor U8566 (N_8566,N_5728,N_7107);
xor U8567 (N_8567,N_6835,N_5199);
xor U8568 (N_8568,N_6097,N_7201);
and U8569 (N_8569,N_6500,N_5342);
nor U8570 (N_8570,N_7319,N_5279);
nor U8571 (N_8571,N_6464,N_5168);
or U8572 (N_8572,N_6528,N_7288);
nor U8573 (N_8573,N_6237,N_7217);
or U8574 (N_8574,N_5291,N_6649);
and U8575 (N_8575,N_5088,N_6883);
xor U8576 (N_8576,N_5481,N_5152);
and U8577 (N_8577,N_7184,N_7112);
nand U8578 (N_8578,N_5800,N_6106);
or U8579 (N_8579,N_7360,N_5075);
nor U8580 (N_8580,N_5201,N_7212);
and U8581 (N_8581,N_5760,N_6114);
or U8582 (N_8582,N_7011,N_5231);
nand U8583 (N_8583,N_6654,N_6542);
or U8584 (N_8584,N_5514,N_6787);
nand U8585 (N_8585,N_5503,N_6032);
or U8586 (N_8586,N_5322,N_5116);
nor U8587 (N_8587,N_6667,N_6616);
nor U8588 (N_8588,N_6051,N_7121);
nor U8589 (N_8589,N_6266,N_6586);
xnor U8590 (N_8590,N_5914,N_5118);
nand U8591 (N_8591,N_5734,N_5002);
nand U8592 (N_8592,N_6691,N_5832);
or U8593 (N_8593,N_6827,N_6993);
nor U8594 (N_8594,N_7177,N_6393);
nor U8595 (N_8595,N_7253,N_6469);
nor U8596 (N_8596,N_5935,N_7018);
nand U8597 (N_8597,N_6390,N_7159);
or U8598 (N_8598,N_6076,N_7299);
or U8599 (N_8599,N_6193,N_7316);
nand U8600 (N_8600,N_6639,N_7188);
nor U8601 (N_8601,N_6509,N_7406);
or U8602 (N_8602,N_6397,N_5467);
nor U8603 (N_8603,N_7187,N_6451);
nor U8604 (N_8604,N_5551,N_7306);
and U8605 (N_8605,N_6615,N_6394);
nor U8606 (N_8606,N_6030,N_5941);
nor U8607 (N_8607,N_6605,N_6629);
and U8608 (N_8608,N_6304,N_6760);
nand U8609 (N_8609,N_5287,N_6530);
and U8610 (N_8610,N_5716,N_5859);
xor U8611 (N_8611,N_5485,N_6291);
and U8612 (N_8612,N_6149,N_5645);
and U8613 (N_8613,N_5890,N_5146);
and U8614 (N_8614,N_6519,N_7094);
and U8615 (N_8615,N_5590,N_7126);
nor U8616 (N_8616,N_6176,N_7154);
nand U8617 (N_8617,N_5345,N_5161);
and U8618 (N_8618,N_5319,N_6016);
nor U8619 (N_8619,N_7161,N_5447);
nor U8620 (N_8620,N_6060,N_5651);
and U8621 (N_8621,N_6037,N_5368);
and U8622 (N_8622,N_5560,N_7263);
and U8623 (N_8623,N_6295,N_6999);
nand U8624 (N_8624,N_7335,N_6089);
or U8625 (N_8625,N_5226,N_7365);
nand U8626 (N_8626,N_7219,N_6116);
or U8627 (N_8627,N_5886,N_6300);
nor U8628 (N_8628,N_5329,N_6440);
nor U8629 (N_8629,N_7462,N_5138);
or U8630 (N_8630,N_6127,N_5566);
xor U8631 (N_8631,N_5332,N_5947);
and U8632 (N_8632,N_5909,N_6593);
nor U8633 (N_8633,N_6435,N_6299);
and U8634 (N_8634,N_6940,N_5672);
and U8635 (N_8635,N_6112,N_5248);
and U8636 (N_8636,N_6342,N_5764);
nor U8637 (N_8637,N_6640,N_7451);
or U8638 (N_8638,N_5222,N_5249);
nor U8639 (N_8639,N_5937,N_6429);
or U8640 (N_8640,N_6322,N_5084);
or U8641 (N_8641,N_6987,N_5618);
and U8642 (N_8642,N_6111,N_6620);
xor U8643 (N_8643,N_7450,N_5750);
and U8644 (N_8644,N_5776,N_5736);
or U8645 (N_8645,N_5213,N_5458);
or U8646 (N_8646,N_7213,N_7477);
nor U8647 (N_8647,N_6693,N_7416);
or U8648 (N_8648,N_6876,N_5850);
nor U8649 (N_8649,N_5889,N_5515);
nor U8650 (N_8650,N_7404,N_5580);
or U8651 (N_8651,N_6491,N_5298);
nand U8652 (N_8652,N_5275,N_6630);
nor U8653 (N_8653,N_6427,N_5785);
and U8654 (N_8654,N_7242,N_6350);
xnor U8655 (N_8655,N_5038,N_7002);
xnor U8656 (N_8656,N_6232,N_5137);
or U8657 (N_8657,N_6364,N_5720);
nor U8658 (N_8658,N_6462,N_7113);
nor U8659 (N_8659,N_6303,N_6276);
or U8660 (N_8660,N_6011,N_6915);
nand U8661 (N_8661,N_5022,N_5335);
nand U8662 (N_8662,N_5308,N_6891);
nand U8663 (N_8663,N_6919,N_5064);
nor U8664 (N_8664,N_6294,N_6807);
nand U8665 (N_8665,N_7312,N_7262);
or U8666 (N_8666,N_5011,N_6400);
nand U8667 (N_8667,N_5364,N_6908);
nand U8668 (N_8668,N_6201,N_7463);
or U8669 (N_8669,N_6326,N_5071);
nor U8670 (N_8670,N_6324,N_6723);
and U8671 (N_8671,N_5383,N_6748);
and U8672 (N_8672,N_7244,N_7315);
nand U8673 (N_8673,N_7487,N_5972);
nor U8674 (N_8674,N_6618,N_5944);
and U8675 (N_8675,N_5052,N_7028);
nand U8676 (N_8676,N_7153,N_6982);
nand U8677 (N_8677,N_5433,N_6969);
and U8678 (N_8678,N_6343,N_6584);
nor U8679 (N_8679,N_6172,N_5630);
and U8680 (N_8680,N_6093,N_6750);
nand U8681 (N_8681,N_6784,N_6255);
or U8682 (N_8682,N_5428,N_7033);
nand U8683 (N_8683,N_6087,N_6560);
nand U8684 (N_8684,N_6580,N_7322);
nand U8685 (N_8685,N_6308,N_5609);
and U8686 (N_8686,N_5864,N_6952);
nor U8687 (N_8687,N_6700,N_6941);
nor U8688 (N_8688,N_6706,N_6425);
xor U8689 (N_8689,N_6567,N_5940);
nand U8690 (N_8690,N_6136,N_6340);
nand U8691 (N_8691,N_5230,N_5524);
nor U8692 (N_8692,N_6878,N_6078);
nor U8693 (N_8693,N_6661,N_6059);
nand U8694 (N_8694,N_5925,N_5733);
xnor U8695 (N_8695,N_6012,N_5615);
xnor U8696 (N_8696,N_6144,N_5165);
or U8697 (N_8697,N_6268,N_6209);
or U8698 (N_8698,N_5078,N_5835);
nor U8699 (N_8699,N_5664,N_6523);
nor U8700 (N_8700,N_7292,N_6767);
nor U8701 (N_8701,N_5218,N_5259);
and U8702 (N_8702,N_5857,N_5742);
xor U8703 (N_8703,N_5787,N_7067);
nand U8704 (N_8704,N_6934,N_6113);
xnor U8705 (N_8705,N_6514,N_6480);
or U8706 (N_8706,N_5107,N_6438);
nand U8707 (N_8707,N_6036,N_6838);
nand U8708 (N_8708,N_7275,N_6132);
or U8709 (N_8709,N_6591,N_6282);
and U8710 (N_8710,N_5702,N_5031);
and U8711 (N_8711,N_7310,N_6634);
nor U8712 (N_8712,N_6361,N_7071);
nand U8713 (N_8713,N_7429,N_6662);
or U8714 (N_8714,N_6665,N_5444);
xnor U8715 (N_8715,N_5056,N_7040);
or U8716 (N_8716,N_5594,N_5571);
xor U8717 (N_8717,N_6205,N_7369);
and U8718 (N_8718,N_5960,N_5965);
or U8719 (N_8719,N_5157,N_6407);
nand U8720 (N_8720,N_5771,N_5959);
or U8721 (N_8721,N_6527,N_7118);
and U8722 (N_8722,N_6674,N_6812);
or U8723 (N_8723,N_6890,N_7489);
xor U8724 (N_8724,N_7053,N_7057);
nand U8725 (N_8725,N_6489,N_7186);
or U8726 (N_8726,N_6081,N_7466);
nand U8727 (N_8727,N_6456,N_5176);
and U8728 (N_8728,N_6358,N_7268);
and U8729 (N_8729,N_7396,N_5624);
and U8730 (N_8730,N_6015,N_7210);
nand U8731 (N_8731,N_7109,N_7009);
nor U8732 (N_8732,N_7327,N_7007);
nor U8733 (N_8733,N_7050,N_6854);
nor U8734 (N_8734,N_7411,N_6065);
nand U8735 (N_8735,N_5115,N_5748);
nor U8736 (N_8736,N_6441,N_6726);
nor U8737 (N_8737,N_7181,N_6800);
nor U8738 (N_8738,N_6535,N_5262);
and U8739 (N_8739,N_7182,N_6656);
nor U8740 (N_8740,N_6899,N_7198);
or U8741 (N_8741,N_5713,N_5616);
nor U8742 (N_8742,N_6895,N_5531);
nand U8743 (N_8743,N_5824,N_5522);
xor U8744 (N_8744,N_5187,N_6346);
nand U8745 (N_8745,N_6122,N_7276);
nand U8746 (N_8746,N_6797,N_6494);
xor U8747 (N_8747,N_6964,N_5621);
or U8748 (N_8748,N_5186,N_6625);
and U8749 (N_8749,N_5401,N_6026);
nor U8750 (N_8750,N_5819,N_7349);
nand U8751 (N_8751,N_5931,N_5381);
nor U8752 (N_8752,N_6435,N_5076);
xor U8753 (N_8753,N_6048,N_5152);
and U8754 (N_8754,N_6712,N_5752);
nand U8755 (N_8755,N_6053,N_7082);
and U8756 (N_8756,N_6236,N_6721);
nand U8757 (N_8757,N_6015,N_5056);
and U8758 (N_8758,N_6503,N_7188);
or U8759 (N_8759,N_7315,N_7455);
nor U8760 (N_8760,N_5397,N_6380);
xnor U8761 (N_8761,N_6409,N_5677);
or U8762 (N_8762,N_5857,N_6027);
or U8763 (N_8763,N_6729,N_5395);
and U8764 (N_8764,N_6888,N_7079);
or U8765 (N_8765,N_7087,N_5922);
xnor U8766 (N_8766,N_6097,N_7319);
and U8767 (N_8767,N_5127,N_5335);
xnor U8768 (N_8768,N_6108,N_6030);
nand U8769 (N_8769,N_6685,N_5135);
nand U8770 (N_8770,N_5048,N_5571);
nor U8771 (N_8771,N_6098,N_6913);
nor U8772 (N_8772,N_7189,N_6601);
nor U8773 (N_8773,N_5878,N_6626);
or U8774 (N_8774,N_5851,N_7015);
nand U8775 (N_8775,N_7152,N_5246);
nor U8776 (N_8776,N_6145,N_6029);
nand U8777 (N_8777,N_6031,N_5242);
or U8778 (N_8778,N_6678,N_5508);
nand U8779 (N_8779,N_6517,N_5514);
and U8780 (N_8780,N_6004,N_5029);
nand U8781 (N_8781,N_7400,N_5404);
or U8782 (N_8782,N_6844,N_5840);
and U8783 (N_8783,N_6934,N_7090);
nor U8784 (N_8784,N_7057,N_5262);
nand U8785 (N_8785,N_6077,N_5334);
and U8786 (N_8786,N_6195,N_5770);
nor U8787 (N_8787,N_5391,N_5761);
nor U8788 (N_8788,N_5261,N_5801);
nor U8789 (N_8789,N_6004,N_7137);
or U8790 (N_8790,N_7395,N_6150);
xor U8791 (N_8791,N_6458,N_6537);
nand U8792 (N_8792,N_5509,N_6633);
or U8793 (N_8793,N_5010,N_7343);
or U8794 (N_8794,N_6766,N_6850);
nand U8795 (N_8795,N_5636,N_5340);
nand U8796 (N_8796,N_6728,N_6670);
nor U8797 (N_8797,N_6148,N_6505);
or U8798 (N_8798,N_6186,N_5245);
nand U8799 (N_8799,N_6351,N_6347);
or U8800 (N_8800,N_5953,N_7111);
and U8801 (N_8801,N_5059,N_5688);
or U8802 (N_8802,N_7132,N_6415);
and U8803 (N_8803,N_6513,N_5814);
xor U8804 (N_8804,N_7196,N_5637);
and U8805 (N_8805,N_6723,N_5925);
and U8806 (N_8806,N_7045,N_6358);
or U8807 (N_8807,N_6390,N_5720);
nor U8808 (N_8808,N_5751,N_6018);
nor U8809 (N_8809,N_7045,N_6899);
and U8810 (N_8810,N_6393,N_7219);
or U8811 (N_8811,N_5278,N_7353);
nand U8812 (N_8812,N_6192,N_6297);
nor U8813 (N_8813,N_6773,N_6441);
and U8814 (N_8814,N_6099,N_7100);
nor U8815 (N_8815,N_6485,N_5234);
or U8816 (N_8816,N_6618,N_5464);
or U8817 (N_8817,N_5932,N_7121);
or U8818 (N_8818,N_6373,N_5234);
or U8819 (N_8819,N_6856,N_5657);
and U8820 (N_8820,N_6290,N_6025);
nand U8821 (N_8821,N_7404,N_6890);
and U8822 (N_8822,N_7455,N_5889);
nor U8823 (N_8823,N_6147,N_5408);
nor U8824 (N_8824,N_6574,N_5528);
nor U8825 (N_8825,N_5385,N_5507);
and U8826 (N_8826,N_5200,N_7182);
nand U8827 (N_8827,N_5674,N_6044);
or U8828 (N_8828,N_5032,N_6934);
xnor U8829 (N_8829,N_5252,N_6499);
or U8830 (N_8830,N_5975,N_6835);
nor U8831 (N_8831,N_6937,N_6070);
or U8832 (N_8832,N_5429,N_6482);
nand U8833 (N_8833,N_5646,N_6594);
or U8834 (N_8834,N_6900,N_6665);
xnor U8835 (N_8835,N_6199,N_6049);
nor U8836 (N_8836,N_5063,N_5404);
or U8837 (N_8837,N_6268,N_5233);
xor U8838 (N_8838,N_5318,N_6987);
nand U8839 (N_8839,N_6028,N_5050);
or U8840 (N_8840,N_7310,N_5095);
or U8841 (N_8841,N_6174,N_6537);
and U8842 (N_8842,N_5084,N_5780);
or U8843 (N_8843,N_6937,N_6800);
nor U8844 (N_8844,N_6365,N_6319);
nand U8845 (N_8845,N_5435,N_5517);
nand U8846 (N_8846,N_7028,N_7146);
or U8847 (N_8847,N_5057,N_6344);
nand U8848 (N_8848,N_6526,N_7321);
nor U8849 (N_8849,N_5541,N_5033);
and U8850 (N_8850,N_7377,N_5406);
or U8851 (N_8851,N_6784,N_5627);
and U8852 (N_8852,N_5165,N_5803);
nor U8853 (N_8853,N_5758,N_7340);
or U8854 (N_8854,N_5917,N_6643);
nand U8855 (N_8855,N_5466,N_5799);
nor U8856 (N_8856,N_5824,N_7145);
xor U8857 (N_8857,N_5418,N_5268);
nand U8858 (N_8858,N_6236,N_5511);
nor U8859 (N_8859,N_5613,N_6725);
or U8860 (N_8860,N_5786,N_6741);
or U8861 (N_8861,N_7418,N_5538);
and U8862 (N_8862,N_6614,N_6307);
nor U8863 (N_8863,N_6059,N_5187);
or U8864 (N_8864,N_6480,N_5901);
and U8865 (N_8865,N_7074,N_7492);
nor U8866 (N_8866,N_5726,N_5236);
nor U8867 (N_8867,N_6970,N_5528);
nor U8868 (N_8868,N_6469,N_6182);
or U8869 (N_8869,N_6997,N_7049);
xnor U8870 (N_8870,N_7323,N_5798);
nand U8871 (N_8871,N_5175,N_6754);
nand U8872 (N_8872,N_5740,N_6998);
xor U8873 (N_8873,N_5002,N_6030);
nor U8874 (N_8874,N_5759,N_5428);
xnor U8875 (N_8875,N_5252,N_7030);
nor U8876 (N_8876,N_6078,N_5372);
nor U8877 (N_8877,N_7112,N_5306);
nand U8878 (N_8878,N_5240,N_6133);
or U8879 (N_8879,N_5610,N_6568);
nand U8880 (N_8880,N_5010,N_5099);
nor U8881 (N_8881,N_7245,N_5837);
nor U8882 (N_8882,N_6634,N_6868);
nand U8883 (N_8883,N_6507,N_5609);
nand U8884 (N_8884,N_5883,N_5963);
and U8885 (N_8885,N_5753,N_5808);
nor U8886 (N_8886,N_6810,N_6740);
and U8887 (N_8887,N_5559,N_6291);
nor U8888 (N_8888,N_5681,N_6213);
and U8889 (N_8889,N_7110,N_7331);
nor U8890 (N_8890,N_6066,N_6794);
nand U8891 (N_8891,N_5200,N_6790);
and U8892 (N_8892,N_7394,N_7037);
or U8893 (N_8893,N_6066,N_5146);
nand U8894 (N_8894,N_6108,N_6396);
nand U8895 (N_8895,N_7365,N_7161);
or U8896 (N_8896,N_6717,N_6202);
nor U8897 (N_8897,N_5939,N_7471);
and U8898 (N_8898,N_7493,N_5222);
nand U8899 (N_8899,N_6577,N_6836);
nor U8900 (N_8900,N_6698,N_5911);
or U8901 (N_8901,N_5213,N_6409);
or U8902 (N_8902,N_7129,N_5810);
and U8903 (N_8903,N_5052,N_6287);
nor U8904 (N_8904,N_6691,N_6251);
or U8905 (N_8905,N_5666,N_6698);
nor U8906 (N_8906,N_6638,N_7339);
and U8907 (N_8907,N_5622,N_7355);
nand U8908 (N_8908,N_5776,N_5280);
and U8909 (N_8909,N_6087,N_6420);
xnor U8910 (N_8910,N_7161,N_5244);
or U8911 (N_8911,N_5592,N_6045);
nor U8912 (N_8912,N_6465,N_5170);
nor U8913 (N_8913,N_6445,N_5433);
nor U8914 (N_8914,N_6937,N_6045);
nand U8915 (N_8915,N_5176,N_6625);
nand U8916 (N_8916,N_6093,N_6738);
or U8917 (N_8917,N_6759,N_7110);
nand U8918 (N_8918,N_6002,N_6229);
and U8919 (N_8919,N_5450,N_5233);
nor U8920 (N_8920,N_6033,N_5909);
nor U8921 (N_8921,N_5687,N_6981);
nand U8922 (N_8922,N_6653,N_6934);
or U8923 (N_8923,N_5740,N_7050);
nor U8924 (N_8924,N_6040,N_6218);
or U8925 (N_8925,N_7266,N_6822);
or U8926 (N_8926,N_6537,N_5986);
nor U8927 (N_8927,N_5537,N_5229);
nor U8928 (N_8928,N_6896,N_5535);
nand U8929 (N_8929,N_7097,N_6719);
nand U8930 (N_8930,N_7150,N_6995);
or U8931 (N_8931,N_6895,N_5090);
xnor U8932 (N_8932,N_6889,N_6308);
nor U8933 (N_8933,N_6956,N_5122);
nor U8934 (N_8934,N_6593,N_5046);
or U8935 (N_8935,N_6116,N_5376);
nand U8936 (N_8936,N_5362,N_6788);
xnor U8937 (N_8937,N_7365,N_6100);
and U8938 (N_8938,N_5186,N_7448);
nor U8939 (N_8939,N_5833,N_5486);
nand U8940 (N_8940,N_6769,N_7017);
nor U8941 (N_8941,N_7442,N_6231);
nand U8942 (N_8942,N_5396,N_6343);
and U8943 (N_8943,N_6992,N_6990);
and U8944 (N_8944,N_6288,N_5013);
and U8945 (N_8945,N_6504,N_5817);
or U8946 (N_8946,N_5994,N_6917);
and U8947 (N_8947,N_5620,N_5971);
nor U8948 (N_8948,N_6728,N_6646);
nor U8949 (N_8949,N_6875,N_5989);
or U8950 (N_8950,N_5059,N_6696);
xor U8951 (N_8951,N_6091,N_5376);
nand U8952 (N_8952,N_6084,N_5514);
or U8953 (N_8953,N_7295,N_6271);
or U8954 (N_8954,N_6163,N_6413);
or U8955 (N_8955,N_7195,N_6152);
or U8956 (N_8956,N_5006,N_6473);
and U8957 (N_8957,N_5752,N_6529);
nand U8958 (N_8958,N_5715,N_7048);
nand U8959 (N_8959,N_7163,N_6635);
nand U8960 (N_8960,N_5219,N_6711);
or U8961 (N_8961,N_6133,N_5596);
nor U8962 (N_8962,N_6986,N_5271);
nand U8963 (N_8963,N_7056,N_5101);
nand U8964 (N_8964,N_7044,N_5381);
or U8965 (N_8965,N_5867,N_5049);
nand U8966 (N_8966,N_5999,N_7473);
nand U8967 (N_8967,N_5247,N_6994);
or U8968 (N_8968,N_5543,N_7488);
nand U8969 (N_8969,N_6857,N_6679);
nand U8970 (N_8970,N_5773,N_7028);
nand U8971 (N_8971,N_5532,N_5650);
nor U8972 (N_8972,N_5684,N_5627);
nand U8973 (N_8973,N_7345,N_6739);
or U8974 (N_8974,N_5534,N_7062);
and U8975 (N_8975,N_7304,N_5817);
nand U8976 (N_8976,N_7090,N_6050);
or U8977 (N_8977,N_6579,N_7002);
and U8978 (N_8978,N_5953,N_6234);
nand U8979 (N_8979,N_7499,N_7413);
nor U8980 (N_8980,N_6330,N_7075);
nand U8981 (N_8981,N_5024,N_6259);
nor U8982 (N_8982,N_5195,N_6670);
and U8983 (N_8983,N_7312,N_7046);
nand U8984 (N_8984,N_6291,N_6512);
nand U8985 (N_8985,N_6256,N_5013);
nor U8986 (N_8986,N_5858,N_6608);
nor U8987 (N_8987,N_6554,N_7242);
or U8988 (N_8988,N_6188,N_6983);
xor U8989 (N_8989,N_5329,N_5036);
xnor U8990 (N_8990,N_6875,N_6716);
and U8991 (N_8991,N_5995,N_6933);
or U8992 (N_8992,N_7318,N_6874);
nor U8993 (N_8993,N_7062,N_5490);
nand U8994 (N_8994,N_5239,N_6981);
nand U8995 (N_8995,N_5809,N_5040);
xnor U8996 (N_8996,N_5429,N_6551);
nand U8997 (N_8997,N_6111,N_5341);
or U8998 (N_8998,N_6685,N_6216);
xor U8999 (N_8999,N_7033,N_6339);
nand U9000 (N_9000,N_5204,N_6250);
nor U9001 (N_9001,N_7057,N_5532);
or U9002 (N_9002,N_5572,N_7031);
nor U9003 (N_9003,N_6508,N_6853);
or U9004 (N_9004,N_5719,N_6375);
nor U9005 (N_9005,N_7176,N_6375);
nor U9006 (N_9006,N_6087,N_6784);
and U9007 (N_9007,N_7391,N_6004);
nand U9008 (N_9008,N_6732,N_6466);
nand U9009 (N_9009,N_5376,N_5401);
nor U9010 (N_9010,N_5455,N_5919);
and U9011 (N_9011,N_6479,N_6983);
nand U9012 (N_9012,N_7398,N_5184);
or U9013 (N_9013,N_5151,N_5369);
nand U9014 (N_9014,N_6613,N_5816);
or U9015 (N_9015,N_5131,N_6701);
and U9016 (N_9016,N_5310,N_5762);
nor U9017 (N_9017,N_7437,N_6890);
nor U9018 (N_9018,N_5648,N_6580);
nor U9019 (N_9019,N_5654,N_5134);
nor U9020 (N_9020,N_5650,N_6641);
xor U9021 (N_9021,N_5665,N_6488);
nand U9022 (N_9022,N_5293,N_5617);
or U9023 (N_9023,N_6866,N_6497);
and U9024 (N_9024,N_6381,N_5194);
nor U9025 (N_9025,N_5624,N_6795);
or U9026 (N_9026,N_7342,N_6416);
and U9027 (N_9027,N_6700,N_6501);
and U9028 (N_9028,N_5712,N_5805);
and U9029 (N_9029,N_5131,N_7317);
nor U9030 (N_9030,N_5903,N_5181);
or U9031 (N_9031,N_6743,N_5222);
xor U9032 (N_9032,N_7054,N_5479);
nand U9033 (N_9033,N_6520,N_7261);
and U9034 (N_9034,N_7485,N_6281);
nor U9035 (N_9035,N_7375,N_6233);
nand U9036 (N_9036,N_6029,N_6336);
or U9037 (N_9037,N_6575,N_6050);
nand U9038 (N_9038,N_5132,N_6020);
xnor U9039 (N_9039,N_7076,N_7312);
nor U9040 (N_9040,N_6877,N_6770);
and U9041 (N_9041,N_6228,N_5425);
xor U9042 (N_9042,N_6157,N_6758);
and U9043 (N_9043,N_5425,N_5153);
and U9044 (N_9044,N_6167,N_5542);
and U9045 (N_9045,N_6087,N_6348);
or U9046 (N_9046,N_7130,N_5734);
nor U9047 (N_9047,N_6693,N_5697);
or U9048 (N_9048,N_6013,N_6398);
nor U9049 (N_9049,N_5674,N_7049);
nor U9050 (N_9050,N_7222,N_5285);
xor U9051 (N_9051,N_6030,N_6991);
nor U9052 (N_9052,N_6454,N_6367);
or U9053 (N_9053,N_7169,N_6446);
nor U9054 (N_9054,N_6009,N_5830);
nand U9055 (N_9055,N_6766,N_5015);
nor U9056 (N_9056,N_6379,N_5290);
nand U9057 (N_9057,N_6204,N_5944);
nand U9058 (N_9058,N_6712,N_6317);
nand U9059 (N_9059,N_6814,N_6534);
and U9060 (N_9060,N_6274,N_6938);
or U9061 (N_9061,N_6904,N_6590);
or U9062 (N_9062,N_5117,N_6808);
and U9063 (N_9063,N_6571,N_7312);
xnor U9064 (N_9064,N_5628,N_5083);
and U9065 (N_9065,N_5293,N_5812);
and U9066 (N_9066,N_7093,N_6018);
nand U9067 (N_9067,N_5812,N_6532);
nand U9068 (N_9068,N_5047,N_6946);
and U9069 (N_9069,N_7467,N_6908);
nand U9070 (N_9070,N_6808,N_5405);
xnor U9071 (N_9071,N_6862,N_7206);
and U9072 (N_9072,N_5108,N_5006);
or U9073 (N_9073,N_5263,N_5055);
nor U9074 (N_9074,N_7397,N_6497);
nor U9075 (N_9075,N_6463,N_6314);
nor U9076 (N_9076,N_5236,N_5014);
xnor U9077 (N_9077,N_5131,N_5353);
and U9078 (N_9078,N_6340,N_6437);
xnor U9079 (N_9079,N_5023,N_7410);
nor U9080 (N_9080,N_7370,N_7390);
or U9081 (N_9081,N_5186,N_7428);
nor U9082 (N_9082,N_7479,N_6925);
or U9083 (N_9083,N_6047,N_7043);
nor U9084 (N_9084,N_5697,N_6314);
or U9085 (N_9085,N_5142,N_6887);
or U9086 (N_9086,N_5764,N_6663);
nand U9087 (N_9087,N_5517,N_6831);
nor U9088 (N_9088,N_6617,N_6374);
nand U9089 (N_9089,N_7180,N_5890);
and U9090 (N_9090,N_5140,N_6693);
or U9091 (N_9091,N_5844,N_5531);
and U9092 (N_9092,N_6597,N_5524);
nor U9093 (N_9093,N_6644,N_5618);
nor U9094 (N_9094,N_5825,N_5864);
or U9095 (N_9095,N_5998,N_5940);
xnor U9096 (N_9096,N_7484,N_6653);
or U9097 (N_9097,N_5179,N_5299);
xnor U9098 (N_9098,N_6039,N_7159);
and U9099 (N_9099,N_5898,N_5388);
xor U9100 (N_9100,N_5426,N_5587);
nor U9101 (N_9101,N_7238,N_6641);
and U9102 (N_9102,N_6753,N_6837);
nand U9103 (N_9103,N_5541,N_7463);
or U9104 (N_9104,N_5084,N_5630);
xnor U9105 (N_9105,N_5493,N_7305);
nor U9106 (N_9106,N_5196,N_6094);
and U9107 (N_9107,N_6668,N_6041);
and U9108 (N_9108,N_5861,N_6360);
or U9109 (N_9109,N_5959,N_5839);
and U9110 (N_9110,N_6268,N_6897);
nand U9111 (N_9111,N_7086,N_5810);
nor U9112 (N_9112,N_7048,N_6352);
nand U9113 (N_9113,N_5507,N_5415);
or U9114 (N_9114,N_6967,N_5556);
nor U9115 (N_9115,N_6205,N_6437);
nand U9116 (N_9116,N_6088,N_6526);
and U9117 (N_9117,N_6615,N_7118);
nand U9118 (N_9118,N_6347,N_6374);
nor U9119 (N_9119,N_6725,N_5043);
or U9120 (N_9120,N_7242,N_5760);
and U9121 (N_9121,N_7311,N_6458);
or U9122 (N_9122,N_6403,N_7386);
or U9123 (N_9123,N_5719,N_6214);
or U9124 (N_9124,N_5346,N_6957);
nor U9125 (N_9125,N_6870,N_5595);
nand U9126 (N_9126,N_5223,N_6038);
nand U9127 (N_9127,N_6340,N_5348);
nor U9128 (N_9128,N_6986,N_5450);
nand U9129 (N_9129,N_5598,N_6051);
nor U9130 (N_9130,N_6869,N_6160);
or U9131 (N_9131,N_7437,N_5785);
and U9132 (N_9132,N_5451,N_6742);
nor U9133 (N_9133,N_6748,N_5642);
xor U9134 (N_9134,N_5307,N_7120);
xor U9135 (N_9135,N_5669,N_5739);
nand U9136 (N_9136,N_5968,N_5287);
or U9137 (N_9137,N_5559,N_5068);
xnor U9138 (N_9138,N_6915,N_5305);
and U9139 (N_9139,N_6983,N_7307);
or U9140 (N_9140,N_6932,N_5537);
nand U9141 (N_9141,N_6447,N_7465);
nor U9142 (N_9142,N_7346,N_5212);
nand U9143 (N_9143,N_6302,N_6842);
nand U9144 (N_9144,N_5788,N_7101);
or U9145 (N_9145,N_5072,N_6608);
nor U9146 (N_9146,N_7147,N_5374);
xnor U9147 (N_9147,N_6106,N_5742);
nor U9148 (N_9148,N_5175,N_5733);
nand U9149 (N_9149,N_6306,N_5580);
xor U9150 (N_9150,N_6431,N_6378);
nor U9151 (N_9151,N_5738,N_5407);
nor U9152 (N_9152,N_6645,N_5169);
and U9153 (N_9153,N_5697,N_7250);
nand U9154 (N_9154,N_6169,N_6188);
or U9155 (N_9155,N_6493,N_6762);
nor U9156 (N_9156,N_6589,N_6145);
or U9157 (N_9157,N_5833,N_7334);
xnor U9158 (N_9158,N_5964,N_5509);
and U9159 (N_9159,N_5108,N_5853);
or U9160 (N_9160,N_5978,N_5525);
or U9161 (N_9161,N_5263,N_7001);
or U9162 (N_9162,N_6780,N_7100);
or U9163 (N_9163,N_6441,N_6690);
or U9164 (N_9164,N_6590,N_7275);
xnor U9165 (N_9165,N_6963,N_7336);
nand U9166 (N_9166,N_5632,N_6439);
or U9167 (N_9167,N_6188,N_7287);
nor U9168 (N_9168,N_7159,N_6775);
nand U9169 (N_9169,N_7309,N_6432);
or U9170 (N_9170,N_6815,N_6894);
nand U9171 (N_9171,N_6941,N_6389);
nand U9172 (N_9172,N_6961,N_5773);
nor U9173 (N_9173,N_6709,N_6476);
and U9174 (N_9174,N_5344,N_5129);
nor U9175 (N_9175,N_7386,N_7430);
and U9176 (N_9176,N_6802,N_5822);
or U9177 (N_9177,N_7005,N_5953);
nor U9178 (N_9178,N_6171,N_5198);
nor U9179 (N_9179,N_6129,N_5213);
nor U9180 (N_9180,N_5995,N_5627);
xor U9181 (N_9181,N_5767,N_6160);
and U9182 (N_9182,N_6343,N_5543);
and U9183 (N_9183,N_6062,N_7124);
and U9184 (N_9184,N_5387,N_6652);
nor U9185 (N_9185,N_5799,N_6172);
and U9186 (N_9186,N_6004,N_5879);
nor U9187 (N_9187,N_5239,N_5401);
or U9188 (N_9188,N_6202,N_5951);
nand U9189 (N_9189,N_7170,N_5361);
and U9190 (N_9190,N_5364,N_5470);
xnor U9191 (N_9191,N_5422,N_5974);
nand U9192 (N_9192,N_6554,N_7356);
or U9193 (N_9193,N_6768,N_6204);
and U9194 (N_9194,N_5149,N_7172);
nor U9195 (N_9195,N_6840,N_5392);
nor U9196 (N_9196,N_5545,N_6949);
nor U9197 (N_9197,N_6243,N_5439);
or U9198 (N_9198,N_6239,N_5904);
nor U9199 (N_9199,N_6358,N_6293);
nor U9200 (N_9200,N_5824,N_6475);
and U9201 (N_9201,N_6541,N_5801);
nand U9202 (N_9202,N_5857,N_5513);
and U9203 (N_9203,N_6501,N_5056);
and U9204 (N_9204,N_5296,N_5044);
nor U9205 (N_9205,N_5545,N_5070);
and U9206 (N_9206,N_6147,N_6475);
and U9207 (N_9207,N_5603,N_5901);
and U9208 (N_9208,N_6231,N_7154);
xor U9209 (N_9209,N_5346,N_5233);
and U9210 (N_9210,N_5469,N_6181);
or U9211 (N_9211,N_5294,N_6353);
nand U9212 (N_9212,N_5984,N_6602);
and U9213 (N_9213,N_6471,N_6464);
or U9214 (N_9214,N_5025,N_5988);
nand U9215 (N_9215,N_5632,N_5537);
or U9216 (N_9216,N_7274,N_6620);
and U9217 (N_9217,N_5807,N_5330);
xor U9218 (N_9218,N_7160,N_6469);
or U9219 (N_9219,N_6770,N_5189);
nand U9220 (N_9220,N_6004,N_5999);
or U9221 (N_9221,N_5501,N_5335);
xor U9222 (N_9222,N_6450,N_6940);
or U9223 (N_9223,N_5872,N_6995);
nor U9224 (N_9224,N_6621,N_7035);
or U9225 (N_9225,N_5760,N_7023);
and U9226 (N_9226,N_5746,N_6677);
nor U9227 (N_9227,N_5793,N_5721);
or U9228 (N_9228,N_5154,N_7164);
and U9229 (N_9229,N_7337,N_5161);
nor U9230 (N_9230,N_5008,N_5230);
or U9231 (N_9231,N_6650,N_7393);
and U9232 (N_9232,N_5760,N_5246);
nor U9233 (N_9233,N_6145,N_5106);
nand U9234 (N_9234,N_5795,N_6466);
nand U9235 (N_9235,N_7163,N_5134);
and U9236 (N_9236,N_6779,N_6504);
nand U9237 (N_9237,N_6920,N_6233);
nor U9238 (N_9238,N_7116,N_5794);
nand U9239 (N_9239,N_6806,N_7459);
and U9240 (N_9240,N_5823,N_7232);
nor U9241 (N_9241,N_6552,N_6897);
nor U9242 (N_9242,N_7412,N_5204);
and U9243 (N_9243,N_6386,N_5791);
and U9244 (N_9244,N_6404,N_5890);
nand U9245 (N_9245,N_6825,N_7190);
and U9246 (N_9246,N_7397,N_5424);
nand U9247 (N_9247,N_5905,N_6933);
nand U9248 (N_9248,N_6460,N_6155);
nand U9249 (N_9249,N_6362,N_6816);
and U9250 (N_9250,N_5215,N_7134);
nor U9251 (N_9251,N_6044,N_5426);
or U9252 (N_9252,N_6545,N_5402);
or U9253 (N_9253,N_5903,N_5106);
and U9254 (N_9254,N_6474,N_5450);
xor U9255 (N_9255,N_6083,N_6404);
nor U9256 (N_9256,N_6825,N_6965);
nand U9257 (N_9257,N_6816,N_6939);
xnor U9258 (N_9258,N_5529,N_6456);
and U9259 (N_9259,N_5478,N_5099);
nor U9260 (N_9260,N_7459,N_5930);
nor U9261 (N_9261,N_6604,N_5738);
nor U9262 (N_9262,N_6686,N_7237);
nand U9263 (N_9263,N_6616,N_6030);
xor U9264 (N_9264,N_6301,N_7356);
nand U9265 (N_9265,N_6250,N_6814);
or U9266 (N_9266,N_6319,N_6682);
nand U9267 (N_9267,N_6568,N_6682);
and U9268 (N_9268,N_6655,N_6134);
or U9269 (N_9269,N_5125,N_6618);
or U9270 (N_9270,N_6225,N_7125);
nand U9271 (N_9271,N_6838,N_7228);
nand U9272 (N_9272,N_6016,N_6285);
and U9273 (N_9273,N_6845,N_7406);
nor U9274 (N_9274,N_7278,N_6406);
or U9275 (N_9275,N_5857,N_6249);
and U9276 (N_9276,N_5735,N_6486);
or U9277 (N_9277,N_7426,N_5248);
nor U9278 (N_9278,N_7214,N_7197);
nor U9279 (N_9279,N_7445,N_6024);
nor U9280 (N_9280,N_7221,N_5553);
nor U9281 (N_9281,N_6633,N_5050);
nand U9282 (N_9282,N_7142,N_5933);
and U9283 (N_9283,N_7262,N_5643);
nor U9284 (N_9284,N_6223,N_6550);
nor U9285 (N_9285,N_6815,N_6898);
nand U9286 (N_9286,N_5498,N_6767);
and U9287 (N_9287,N_6647,N_7026);
xnor U9288 (N_9288,N_7097,N_5018);
nand U9289 (N_9289,N_7266,N_6708);
or U9290 (N_9290,N_5960,N_7087);
nand U9291 (N_9291,N_6859,N_7398);
or U9292 (N_9292,N_6200,N_6934);
or U9293 (N_9293,N_5778,N_6769);
xor U9294 (N_9294,N_6487,N_6038);
nand U9295 (N_9295,N_5246,N_6677);
or U9296 (N_9296,N_7346,N_7297);
and U9297 (N_9297,N_5794,N_6830);
or U9298 (N_9298,N_6189,N_6840);
nand U9299 (N_9299,N_6612,N_5468);
and U9300 (N_9300,N_6414,N_6712);
nand U9301 (N_9301,N_6098,N_7467);
or U9302 (N_9302,N_5596,N_5434);
or U9303 (N_9303,N_6643,N_6603);
or U9304 (N_9304,N_5298,N_6840);
xnor U9305 (N_9305,N_7014,N_5269);
or U9306 (N_9306,N_6818,N_7386);
xor U9307 (N_9307,N_6607,N_6386);
or U9308 (N_9308,N_7227,N_6597);
nor U9309 (N_9309,N_6962,N_5426);
or U9310 (N_9310,N_5400,N_5997);
and U9311 (N_9311,N_5398,N_6942);
and U9312 (N_9312,N_5126,N_5481);
nand U9313 (N_9313,N_5163,N_5390);
nand U9314 (N_9314,N_5686,N_6146);
or U9315 (N_9315,N_6075,N_5797);
nand U9316 (N_9316,N_5670,N_5378);
and U9317 (N_9317,N_5154,N_5699);
nor U9318 (N_9318,N_5241,N_6168);
nor U9319 (N_9319,N_6005,N_5356);
or U9320 (N_9320,N_5244,N_5557);
or U9321 (N_9321,N_7065,N_5083);
and U9322 (N_9322,N_6379,N_5542);
and U9323 (N_9323,N_6301,N_5818);
or U9324 (N_9324,N_7244,N_5939);
or U9325 (N_9325,N_5631,N_7376);
or U9326 (N_9326,N_5881,N_6529);
and U9327 (N_9327,N_5098,N_5661);
and U9328 (N_9328,N_6263,N_7297);
xor U9329 (N_9329,N_7374,N_5531);
nand U9330 (N_9330,N_5653,N_5940);
or U9331 (N_9331,N_5906,N_6862);
nand U9332 (N_9332,N_6423,N_5676);
nand U9333 (N_9333,N_5051,N_6630);
and U9334 (N_9334,N_5170,N_7134);
nand U9335 (N_9335,N_7109,N_6707);
nand U9336 (N_9336,N_7214,N_5080);
nand U9337 (N_9337,N_6251,N_6153);
nand U9338 (N_9338,N_6333,N_6887);
nand U9339 (N_9339,N_6347,N_7176);
and U9340 (N_9340,N_7255,N_7278);
and U9341 (N_9341,N_5626,N_6653);
nor U9342 (N_9342,N_6389,N_7063);
nand U9343 (N_9343,N_6051,N_6790);
nand U9344 (N_9344,N_5347,N_6539);
or U9345 (N_9345,N_7412,N_7403);
nand U9346 (N_9346,N_5828,N_5834);
nor U9347 (N_9347,N_5812,N_5294);
or U9348 (N_9348,N_5913,N_5499);
nand U9349 (N_9349,N_6683,N_5225);
and U9350 (N_9350,N_7365,N_6654);
xor U9351 (N_9351,N_5152,N_6953);
and U9352 (N_9352,N_6591,N_5542);
or U9353 (N_9353,N_6246,N_6142);
xnor U9354 (N_9354,N_6642,N_5383);
nor U9355 (N_9355,N_6793,N_6116);
nor U9356 (N_9356,N_7278,N_6725);
and U9357 (N_9357,N_6138,N_6201);
nor U9358 (N_9358,N_6709,N_5610);
nand U9359 (N_9359,N_6596,N_7336);
and U9360 (N_9360,N_5612,N_5749);
xnor U9361 (N_9361,N_6533,N_6448);
nor U9362 (N_9362,N_7494,N_5366);
xor U9363 (N_9363,N_6481,N_5951);
nor U9364 (N_9364,N_7317,N_7451);
or U9365 (N_9365,N_6880,N_5384);
nand U9366 (N_9366,N_5889,N_5102);
or U9367 (N_9367,N_6537,N_5881);
or U9368 (N_9368,N_7123,N_6991);
or U9369 (N_9369,N_5603,N_6698);
nor U9370 (N_9370,N_6317,N_7381);
nand U9371 (N_9371,N_5069,N_6478);
nand U9372 (N_9372,N_6346,N_5111);
nor U9373 (N_9373,N_6633,N_7475);
nand U9374 (N_9374,N_5854,N_6747);
nor U9375 (N_9375,N_5227,N_7439);
and U9376 (N_9376,N_5601,N_6436);
or U9377 (N_9377,N_6003,N_6553);
xnor U9378 (N_9378,N_5782,N_6292);
and U9379 (N_9379,N_6847,N_6559);
xnor U9380 (N_9380,N_5257,N_5681);
nand U9381 (N_9381,N_5599,N_6528);
nand U9382 (N_9382,N_7006,N_7264);
or U9383 (N_9383,N_5389,N_5542);
nand U9384 (N_9384,N_5584,N_6691);
nand U9385 (N_9385,N_5925,N_6085);
xnor U9386 (N_9386,N_5633,N_6482);
nand U9387 (N_9387,N_6863,N_6970);
xnor U9388 (N_9388,N_7436,N_6356);
nand U9389 (N_9389,N_6586,N_7457);
and U9390 (N_9390,N_7454,N_6265);
nand U9391 (N_9391,N_6210,N_5633);
nand U9392 (N_9392,N_6085,N_5221);
xor U9393 (N_9393,N_5861,N_5568);
nand U9394 (N_9394,N_5358,N_6520);
xor U9395 (N_9395,N_7274,N_7361);
or U9396 (N_9396,N_7108,N_6693);
or U9397 (N_9397,N_5486,N_5856);
or U9398 (N_9398,N_5694,N_6378);
xor U9399 (N_9399,N_5217,N_6830);
nor U9400 (N_9400,N_6825,N_5629);
or U9401 (N_9401,N_7097,N_7129);
or U9402 (N_9402,N_6080,N_5201);
nand U9403 (N_9403,N_6273,N_6778);
or U9404 (N_9404,N_5389,N_6981);
nand U9405 (N_9405,N_6135,N_6882);
nor U9406 (N_9406,N_5701,N_7274);
or U9407 (N_9407,N_5654,N_7399);
and U9408 (N_9408,N_5381,N_6681);
nand U9409 (N_9409,N_6971,N_6723);
xor U9410 (N_9410,N_5479,N_5359);
or U9411 (N_9411,N_6762,N_7181);
nor U9412 (N_9412,N_7177,N_6284);
nor U9413 (N_9413,N_5898,N_5728);
or U9414 (N_9414,N_6998,N_7438);
or U9415 (N_9415,N_7200,N_7078);
or U9416 (N_9416,N_6238,N_5178);
or U9417 (N_9417,N_5622,N_5317);
nand U9418 (N_9418,N_5460,N_5316);
or U9419 (N_9419,N_7133,N_6214);
nor U9420 (N_9420,N_6696,N_5932);
nand U9421 (N_9421,N_6721,N_5563);
nand U9422 (N_9422,N_6266,N_6842);
nor U9423 (N_9423,N_7183,N_5188);
nand U9424 (N_9424,N_6708,N_5477);
or U9425 (N_9425,N_6917,N_5538);
nand U9426 (N_9426,N_6400,N_5549);
xnor U9427 (N_9427,N_6044,N_5583);
or U9428 (N_9428,N_6153,N_7327);
nor U9429 (N_9429,N_6497,N_5956);
and U9430 (N_9430,N_6738,N_5012);
xnor U9431 (N_9431,N_6906,N_6447);
and U9432 (N_9432,N_5149,N_6829);
or U9433 (N_9433,N_6633,N_5852);
nor U9434 (N_9434,N_6760,N_5517);
nor U9435 (N_9435,N_6444,N_6245);
or U9436 (N_9436,N_5859,N_6173);
or U9437 (N_9437,N_5116,N_6313);
nand U9438 (N_9438,N_6408,N_6114);
and U9439 (N_9439,N_5390,N_5126);
and U9440 (N_9440,N_5931,N_6309);
or U9441 (N_9441,N_6288,N_6816);
nor U9442 (N_9442,N_7377,N_7259);
and U9443 (N_9443,N_6078,N_5972);
nand U9444 (N_9444,N_5166,N_6852);
or U9445 (N_9445,N_6128,N_5494);
nor U9446 (N_9446,N_5745,N_5955);
or U9447 (N_9447,N_7318,N_6567);
and U9448 (N_9448,N_7330,N_6209);
or U9449 (N_9449,N_6162,N_5776);
xnor U9450 (N_9450,N_7250,N_5392);
nand U9451 (N_9451,N_6575,N_7406);
nor U9452 (N_9452,N_7247,N_5315);
nor U9453 (N_9453,N_7396,N_6469);
nand U9454 (N_9454,N_6276,N_6831);
nor U9455 (N_9455,N_7388,N_5664);
nand U9456 (N_9456,N_6543,N_6952);
or U9457 (N_9457,N_6320,N_6283);
or U9458 (N_9458,N_6331,N_5063);
and U9459 (N_9459,N_6383,N_5647);
and U9460 (N_9460,N_7057,N_7007);
nand U9461 (N_9461,N_5899,N_6322);
nor U9462 (N_9462,N_6362,N_5113);
xor U9463 (N_9463,N_5243,N_5612);
xnor U9464 (N_9464,N_7028,N_6209);
and U9465 (N_9465,N_6721,N_7272);
nor U9466 (N_9466,N_7030,N_6972);
nand U9467 (N_9467,N_5275,N_5067);
nand U9468 (N_9468,N_6969,N_7039);
nand U9469 (N_9469,N_6432,N_6558);
nor U9470 (N_9470,N_6939,N_5878);
and U9471 (N_9471,N_5859,N_7048);
and U9472 (N_9472,N_5888,N_5526);
nor U9473 (N_9473,N_6953,N_7049);
nor U9474 (N_9474,N_7304,N_6775);
and U9475 (N_9475,N_7103,N_6799);
nand U9476 (N_9476,N_6883,N_5471);
nand U9477 (N_9477,N_5603,N_5791);
nand U9478 (N_9478,N_7135,N_6747);
nor U9479 (N_9479,N_5470,N_5128);
and U9480 (N_9480,N_5512,N_5684);
or U9481 (N_9481,N_5493,N_6536);
and U9482 (N_9482,N_6222,N_7360);
nand U9483 (N_9483,N_6963,N_6474);
nand U9484 (N_9484,N_6627,N_5555);
xor U9485 (N_9485,N_6045,N_6496);
and U9486 (N_9486,N_6456,N_5839);
nand U9487 (N_9487,N_5670,N_6466);
nor U9488 (N_9488,N_5623,N_7320);
nor U9489 (N_9489,N_6553,N_5734);
xnor U9490 (N_9490,N_6027,N_5383);
nand U9491 (N_9491,N_6923,N_5314);
nand U9492 (N_9492,N_6215,N_5938);
xor U9493 (N_9493,N_5105,N_6225);
and U9494 (N_9494,N_5143,N_5064);
nor U9495 (N_9495,N_7340,N_6500);
and U9496 (N_9496,N_6714,N_5788);
or U9497 (N_9497,N_5104,N_6882);
xor U9498 (N_9498,N_6156,N_6094);
nor U9499 (N_9499,N_6564,N_5946);
and U9500 (N_9500,N_7058,N_6163);
and U9501 (N_9501,N_7053,N_6808);
and U9502 (N_9502,N_6156,N_5732);
nand U9503 (N_9503,N_6242,N_6126);
or U9504 (N_9504,N_5694,N_5439);
nand U9505 (N_9505,N_6492,N_6657);
or U9506 (N_9506,N_5978,N_6514);
nand U9507 (N_9507,N_7463,N_7229);
and U9508 (N_9508,N_5857,N_7080);
nand U9509 (N_9509,N_6900,N_5124);
or U9510 (N_9510,N_5998,N_5672);
and U9511 (N_9511,N_5691,N_6089);
nand U9512 (N_9512,N_6761,N_6942);
or U9513 (N_9513,N_6012,N_7047);
nand U9514 (N_9514,N_6652,N_5177);
and U9515 (N_9515,N_7337,N_6907);
and U9516 (N_9516,N_6182,N_5892);
and U9517 (N_9517,N_7256,N_6432);
or U9518 (N_9518,N_5714,N_5873);
nor U9519 (N_9519,N_6447,N_7306);
nand U9520 (N_9520,N_5272,N_6925);
xnor U9521 (N_9521,N_6142,N_7289);
and U9522 (N_9522,N_6920,N_5770);
nor U9523 (N_9523,N_5468,N_6594);
nand U9524 (N_9524,N_5039,N_6800);
or U9525 (N_9525,N_5975,N_7345);
xor U9526 (N_9526,N_5111,N_7312);
or U9527 (N_9527,N_7045,N_5841);
and U9528 (N_9528,N_6395,N_6884);
xor U9529 (N_9529,N_6435,N_5782);
or U9530 (N_9530,N_6420,N_6059);
and U9531 (N_9531,N_7124,N_7297);
nand U9532 (N_9532,N_7289,N_7295);
nor U9533 (N_9533,N_7457,N_5429);
xnor U9534 (N_9534,N_6413,N_7252);
xnor U9535 (N_9535,N_5108,N_5343);
nand U9536 (N_9536,N_7428,N_7180);
nor U9537 (N_9537,N_5990,N_6726);
nor U9538 (N_9538,N_5461,N_7286);
nand U9539 (N_9539,N_7455,N_5881);
or U9540 (N_9540,N_6104,N_5135);
nor U9541 (N_9541,N_5694,N_6251);
nand U9542 (N_9542,N_5517,N_7088);
or U9543 (N_9543,N_5240,N_6399);
nor U9544 (N_9544,N_6296,N_5655);
or U9545 (N_9545,N_6519,N_6845);
nand U9546 (N_9546,N_5891,N_6436);
xor U9547 (N_9547,N_7047,N_6389);
nand U9548 (N_9548,N_7074,N_6615);
and U9549 (N_9549,N_5871,N_5648);
or U9550 (N_9550,N_5327,N_5033);
nand U9551 (N_9551,N_6006,N_6726);
or U9552 (N_9552,N_5224,N_6330);
xnor U9553 (N_9553,N_5076,N_5126);
nor U9554 (N_9554,N_6578,N_7492);
nand U9555 (N_9555,N_7180,N_6918);
xor U9556 (N_9556,N_5414,N_6787);
and U9557 (N_9557,N_6581,N_5799);
nor U9558 (N_9558,N_5827,N_7316);
or U9559 (N_9559,N_7242,N_6801);
and U9560 (N_9560,N_6509,N_5709);
and U9561 (N_9561,N_6503,N_6432);
nand U9562 (N_9562,N_6158,N_6941);
and U9563 (N_9563,N_5582,N_7039);
nor U9564 (N_9564,N_5902,N_6497);
nand U9565 (N_9565,N_5631,N_6092);
or U9566 (N_9566,N_6312,N_6994);
nand U9567 (N_9567,N_6748,N_6680);
and U9568 (N_9568,N_7118,N_6159);
nor U9569 (N_9569,N_6468,N_7194);
and U9570 (N_9570,N_6507,N_6810);
or U9571 (N_9571,N_7183,N_7496);
xor U9572 (N_9572,N_5738,N_5657);
and U9573 (N_9573,N_5607,N_7317);
nand U9574 (N_9574,N_6617,N_7102);
nand U9575 (N_9575,N_7235,N_6607);
nand U9576 (N_9576,N_5320,N_5242);
or U9577 (N_9577,N_6489,N_5524);
nand U9578 (N_9578,N_6953,N_5764);
nor U9579 (N_9579,N_6652,N_6463);
nor U9580 (N_9580,N_5333,N_6444);
nor U9581 (N_9581,N_5953,N_6251);
or U9582 (N_9582,N_7331,N_6789);
nand U9583 (N_9583,N_7067,N_5207);
nor U9584 (N_9584,N_6468,N_5351);
nor U9585 (N_9585,N_7217,N_6790);
nand U9586 (N_9586,N_6328,N_5485);
or U9587 (N_9587,N_6731,N_5198);
xor U9588 (N_9588,N_5538,N_5158);
and U9589 (N_9589,N_5411,N_5622);
or U9590 (N_9590,N_5388,N_5073);
and U9591 (N_9591,N_6378,N_6210);
nand U9592 (N_9592,N_6921,N_7267);
nand U9593 (N_9593,N_5409,N_6632);
or U9594 (N_9594,N_5366,N_7228);
nand U9595 (N_9595,N_5342,N_6017);
nand U9596 (N_9596,N_7202,N_6076);
nand U9597 (N_9597,N_7169,N_6692);
xor U9598 (N_9598,N_5271,N_6776);
nand U9599 (N_9599,N_5696,N_6704);
and U9600 (N_9600,N_6019,N_5939);
xor U9601 (N_9601,N_6159,N_5577);
nand U9602 (N_9602,N_6685,N_5492);
or U9603 (N_9603,N_6358,N_5874);
and U9604 (N_9604,N_7084,N_6553);
nand U9605 (N_9605,N_7419,N_6306);
and U9606 (N_9606,N_5223,N_6699);
or U9607 (N_9607,N_6770,N_7081);
xor U9608 (N_9608,N_5926,N_6821);
nor U9609 (N_9609,N_6887,N_6472);
and U9610 (N_9610,N_6361,N_6683);
nor U9611 (N_9611,N_7401,N_5789);
nor U9612 (N_9612,N_6542,N_6807);
xnor U9613 (N_9613,N_5406,N_5933);
nand U9614 (N_9614,N_5758,N_6132);
or U9615 (N_9615,N_7245,N_6463);
nand U9616 (N_9616,N_6814,N_7222);
nand U9617 (N_9617,N_6277,N_5451);
and U9618 (N_9618,N_7471,N_6838);
nor U9619 (N_9619,N_7444,N_6622);
and U9620 (N_9620,N_6189,N_5473);
nand U9621 (N_9621,N_6594,N_5109);
nor U9622 (N_9622,N_6104,N_5524);
or U9623 (N_9623,N_5666,N_5104);
xor U9624 (N_9624,N_7021,N_6405);
nor U9625 (N_9625,N_5310,N_7193);
nor U9626 (N_9626,N_5318,N_5975);
nor U9627 (N_9627,N_5736,N_5392);
nor U9628 (N_9628,N_6815,N_5351);
or U9629 (N_9629,N_5633,N_6910);
nand U9630 (N_9630,N_6393,N_6930);
nor U9631 (N_9631,N_5425,N_7421);
nor U9632 (N_9632,N_7130,N_6298);
or U9633 (N_9633,N_5136,N_6242);
and U9634 (N_9634,N_7490,N_6581);
and U9635 (N_9635,N_5671,N_6482);
nor U9636 (N_9636,N_6074,N_5467);
nor U9637 (N_9637,N_6454,N_7275);
or U9638 (N_9638,N_6358,N_7029);
nand U9639 (N_9639,N_5143,N_7436);
nor U9640 (N_9640,N_7053,N_5029);
xor U9641 (N_9641,N_6922,N_6281);
xor U9642 (N_9642,N_6708,N_6769);
nand U9643 (N_9643,N_6790,N_7367);
nand U9644 (N_9644,N_6139,N_7053);
nand U9645 (N_9645,N_5728,N_5102);
nand U9646 (N_9646,N_5744,N_5040);
and U9647 (N_9647,N_7094,N_6476);
nand U9648 (N_9648,N_6702,N_5579);
nand U9649 (N_9649,N_5029,N_5237);
nor U9650 (N_9650,N_6888,N_7182);
or U9651 (N_9651,N_6769,N_6013);
nand U9652 (N_9652,N_5912,N_7009);
nand U9653 (N_9653,N_7259,N_5099);
xnor U9654 (N_9654,N_6868,N_6581);
nand U9655 (N_9655,N_5323,N_6264);
or U9656 (N_9656,N_5716,N_5120);
nand U9657 (N_9657,N_5047,N_6771);
and U9658 (N_9658,N_6625,N_7326);
nor U9659 (N_9659,N_5340,N_6994);
and U9660 (N_9660,N_6821,N_6409);
or U9661 (N_9661,N_6355,N_6302);
nand U9662 (N_9662,N_5395,N_6852);
nor U9663 (N_9663,N_6714,N_5092);
nand U9664 (N_9664,N_6687,N_6015);
or U9665 (N_9665,N_5908,N_6121);
nand U9666 (N_9666,N_5322,N_6273);
and U9667 (N_9667,N_5851,N_5614);
nand U9668 (N_9668,N_7042,N_6303);
or U9669 (N_9669,N_6230,N_5053);
and U9670 (N_9670,N_7199,N_7348);
nor U9671 (N_9671,N_5164,N_5339);
or U9672 (N_9672,N_5029,N_6016);
nor U9673 (N_9673,N_7331,N_5023);
or U9674 (N_9674,N_6217,N_6041);
nor U9675 (N_9675,N_7277,N_5550);
nor U9676 (N_9676,N_6593,N_6150);
or U9677 (N_9677,N_6408,N_5797);
and U9678 (N_9678,N_5298,N_6611);
and U9679 (N_9679,N_5758,N_6931);
or U9680 (N_9680,N_7155,N_6455);
nor U9681 (N_9681,N_5237,N_6003);
nand U9682 (N_9682,N_5224,N_7307);
or U9683 (N_9683,N_5651,N_6300);
or U9684 (N_9684,N_6370,N_6398);
nand U9685 (N_9685,N_6294,N_6448);
and U9686 (N_9686,N_5578,N_6268);
nor U9687 (N_9687,N_6332,N_6848);
or U9688 (N_9688,N_5550,N_6232);
nand U9689 (N_9689,N_5286,N_5039);
nor U9690 (N_9690,N_6179,N_5648);
nor U9691 (N_9691,N_7301,N_5175);
nand U9692 (N_9692,N_5291,N_6387);
or U9693 (N_9693,N_5541,N_6701);
xnor U9694 (N_9694,N_7429,N_5593);
nor U9695 (N_9695,N_5364,N_5657);
or U9696 (N_9696,N_5838,N_5659);
nor U9697 (N_9697,N_5119,N_6738);
nand U9698 (N_9698,N_5524,N_7437);
or U9699 (N_9699,N_5438,N_7240);
xnor U9700 (N_9700,N_5576,N_6665);
nand U9701 (N_9701,N_5108,N_5808);
nand U9702 (N_9702,N_6171,N_5917);
nor U9703 (N_9703,N_5512,N_6365);
and U9704 (N_9704,N_6842,N_5778);
xnor U9705 (N_9705,N_5621,N_6522);
and U9706 (N_9706,N_6707,N_5665);
xor U9707 (N_9707,N_6291,N_6950);
and U9708 (N_9708,N_6239,N_7264);
nand U9709 (N_9709,N_6657,N_5525);
xnor U9710 (N_9710,N_6949,N_5044);
and U9711 (N_9711,N_6546,N_5514);
and U9712 (N_9712,N_5932,N_6822);
nand U9713 (N_9713,N_6995,N_5198);
or U9714 (N_9714,N_5187,N_7022);
and U9715 (N_9715,N_5702,N_6719);
nor U9716 (N_9716,N_7392,N_6993);
and U9717 (N_9717,N_6030,N_6935);
nor U9718 (N_9718,N_6482,N_5262);
nor U9719 (N_9719,N_7280,N_5762);
nor U9720 (N_9720,N_5711,N_7248);
nand U9721 (N_9721,N_7472,N_6377);
or U9722 (N_9722,N_5958,N_5891);
or U9723 (N_9723,N_6938,N_6854);
nor U9724 (N_9724,N_7036,N_7396);
or U9725 (N_9725,N_5109,N_5808);
or U9726 (N_9726,N_5694,N_5378);
and U9727 (N_9727,N_5412,N_6655);
nor U9728 (N_9728,N_6174,N_5637);
xnor U9729 (N_9729,N_5437,N_5999);
nand U9730 (N_9730,N_7119,N_6354);
nand U9731 (N_9731,N_5602,N_6378);
nor U9732 (N_9732,N_6522,N_6303);
nand U9733 (N_9733,N_6292,N_5336);
nand U9734 (N_9734,N_6563,N_6660);
nor U9735 (N_9735,N_6777,N_7450);
or U9736 (N_9736,N_6422,N_5357);
xor U9737 (N_9737,N_6584,N_7282);
and U9738 (N_9738,N_6936,N_5278);
or U9739 (N_9739,N_7387,N_6895);
or U9740 (N_9740,N_5757,N_6324);
and U9741 (N_9741,N_6216,N_6112);
nand U9742 (N_9742,N_7323,N_6789);
nand U9743 (N_9743,N_6721,N_7267);
xor U9744 (N_9744,N_5398,N_6396);
xor U9745 (N_9745,N_7446,N_7266);
and U9746 (N_9746,N_6893,N_7277);
or U9747 (N_9747,N_5358,N_5166);
nand U9748 (N_9748,N_5599,N_5333);
xnor U9749 (N_9749,N_6721,N_7266);
nand U9750 (N_9750,N_5002,N_6952);
xor U9751 (N_9751,N_6038,N_5327);
or U9752 (N_9752,N_7303,N_7227);
or U9753 (N_9753,N_5011,N_5582);
nand U9754 (N_9754,N_5218,N_5299);
or U9755 (N_9755,N_6679,N_5823);
or U9756 (N_9756,N_6072,N_5253);
or U9757 (N_9757,N_5013,N_5364);
nand U9758 (N_9758,N_7453,N_6418);
and U9759 (N_9759,N_5025,N_7463);
nor U9760 (N_9760,N_6518,N_7408);
nor U9761 (N_9761,N_5434,N_6524);
or U9762 (N_9762,N_6914,N_5524);
or U9763 (N_9763,N_5565,N_5522);
and U9764 (N_9764,N_5283,N_7496);
or U9765 (N_9765,N_6048,N_5134);
nand U9766 (N_9766,N_5207,N_6078);
nor U9767 (N_9767,N_6900,N_6100);
nor U9768 (N_9768,N_7435,N_6422);
or U9769 (N_9769,N_5605,N_5239);
and U9770 (N_9770,N_5494,N_6964);
nand U9771 (N_9771,N_6032,N_5693);
nand U9772 (N_9772,N_6692,N_6570);
nand U9773 (N_9773,N_5358,N_7245);
nor U9774 (N_9774,N_6596,N_6677);
xnor U9775 (N_9775,N_5690,N_5478);
xor U9776 (N_9776,N_6946,N_5452);
nor U9777 (N_9777,N_5277,N_5102);
or U9778 (N_9778,N_5472,N_6700);
nand U9779 (N_9779,N_5698,N_6926);
nand U9780 (N_9780,N_6399,N_5535);
nand U9781 (N_9781,N_6448,N_6338);
or U9782 (N_9782,N_5662,N_5851);
nand U9783 (N_9783,N_6220,N_7250);
nand U9784 (N_9784,N_6324,N_6550);
nor U9785 (N_9785,N_5280,N_7355);
nor U9786 (N_9786,N_6057,N_7438);
xnor U9787 (N_9787,N_7116,N_7228);
nand U9788 (N_9788,N_6334,N_5541);
and U9789 (N_9789,N_6480,N_6269);
and U9790 (N_9790,N_5559,N_6796);
and U9791 (N_9791,N_6174,N_5357);
xor U9792 (N_9792,N_5779,N_5682);
and U9793 (N_9793,N_7389,N_6279);
or U9794 (N_9794,N_7406,N_6451);
nand U9795 (N_9795,N_7218,N_6895);
nand U9796 (N_9796,N_6172,N_6737);
or U9797 (N_9797,N_6078,N_6550);
or U9798 (N_9798,N_6081,N_6990);
or U9799 (N_9799,N_6832,N_6189);
nor U9800 (N_9800,N_5985,N_7214);
and U9801 (N_9801,N_6072,N_6838);
and U9802 (N_9802,N_7324,N_5389);
or U9803 (N_9803,N_7244,N_7388);
nor U9804 (N_9804,N_6227,N_6569);
nor U9805 (N_9805,N_6203,N_6526);
or U9806 (N_9806,N_6777,N_5758);
or U9807 (N_9807,N_6709,N_7368);
and U9808 (N_9808,N_5029,N_6473);
nor U9809 (N_9809,N_7109,N_6801);
xor U9810 (N_9810,N_5458,N_5944);
nand U9811 (N_9811,N_6683,N_5242);
nor U9812 (N_9812,N_7481,N_6414);
nor U9813 (N_9813,N_6480,N_7320);
or U9814 (N_9814,N_5683,N_7100);
nor U9815 (N_9815,N_5473,N_6186);
or U9816 (N_9816,N_5041,N_7055);
xor U9817 (N_9817,N_6499,N_5979);
and U9818 (N_9818,N_5606,N_7453);
nand U9819 (N_9819,N_7388,N_5660);
nor U9820 (N_9820,N_5355,N_6838);
nand U9821 (N_9821,N_6726,N_5255);
nand U9822 (N_9822,N_6241,N_5210);
or U9823 (N_9823,N_5099,N_6521);
nor U9824 (N_9824,N_5172,N_7072);
nor U9825 (N_9825,N_6100,N_6795);
or U9826 (N_9826,N_5731,N_5836);
xnor U9827 (N_9827,N_5081,N_5680);
or U9828 (N_9828,N_5910,N_6043);
nor U9829 (N_9829,N_7428,N_7077);
nor U9830 (N_9830,N_7300,N_7405);
or U9831 (N_9831,N_5700,N_6183);
nand U9832 (N_9832,N_7460,N_6959);
or U9833 (N_9833,N_6221,N_6536);
or U9834 (N_9834,N_6909,N_5179);
or U9835 (N_9835,N_5201,N_5946);
and U9836 (N_9836,N_5762,N_6274);
nor U9837 (N_9837,N_5941,N_5614);
or U9838 (N_9838,N_5467,N_6174);
nor U9839 (N_9839,N_5437,N_7145);
and U9840 (N_9840,N_5293,N_5513);
nor U9841 (N_9841,N_6301,N_6002);
xnor U9842 (N_9842,N_5691,N_5593);
xor U9843 (N_9843,N_7215,N_6755);
nand U9844 (N_9844,N_5546,N_6226);
and U9845 (N_9845,N_6726,N_5864);
nand U9846 (N_9846,N_6760,N_5345);
or U9847 (N_9847,N_5020,N_5647);
nand U9848 (N_9848,N_5294,N_5246);
nor U9849 (N_9849,N_5778,N_6805);
or U9850 (N_9850,N_7466,N_6587);
nand U9851 (N_9851,N_6625,N_6087);
or U9852 (N_9852,N_5047,N_6532);
nor U9853 (N_9853,N_6900,N_6742);
nand U9854 (N_9854,N_5874,N_5262);
and U9855 (N_9855,N_7224,N_7216);
nand U9856 (N_9856,N_5976,N_6286);
xnor U9857 (N_9857,N_5508,N_5291);
nor U9858 (N_9858,N_6960,N_5915);
nor U9859 (N_9859,N_7232,N_5272);
or U9860 (N_9860,N_5143,N_7415);
xnor U9861 (N_9861,N_7066,N_7450);
or U9862 (N_9862,N_5475,N_7305);
nand U9863 (N_9863,N_6421,N_6093);
nor U9864 (N_9864,N_6373,N_7058);
or U9865 (N_9865,N_7333,N_6414);
nor U9866 (N_9866,N_7060,N_5173);
and U9867 (N_9867,N_6720,N_6273);
or U9868 (N_9868,N_6030,N_5279);
or U9869 (N_9869,N_5348,N_5808);
or U9870 (N_9870,N_6393,N_5870);
xnor U9871 (N_9871,N_6298,N_5647);
or U9872 (N_9872,N_5120,N_5101);
or U9873 (N_9873,N_6884,N_6418);
and U9874 (N_9874,N_6920,N_5526);
nand U9875 (N_9875,N_5774,N_5945);
or U9876 (N_9876,N_6753,N_7448);
or U9877 (N_9877,N_7083,N_6721);
or U9878 (N_9878,N_6083,N_7450);
nor U9879 (N_9879,N_6139,N_6250);
nand U9880 (N_9880,N_5821,N_7234);
nor U9881 (N_9881,N_6140,N_5701);
nand U9882 (N_9882,N_5207,N_5706);
nor U9883 (N_9883,N_6432,N_6241);
nand U9884 (N_9884,N_6438,N_5305);
and U9885 (N_9885,N_7064,N_5404);
and U9886 (N_9886,N_7171,N_5280);
nand U9887 (N_9887,N_6558,N_6344);
and U9888 (N_9888,N_5789,N_6330);
and U9889 (N_9889,N_6453,N_6040);
nor U9890 (N_9890,N_6016,N_7270);
nor U9891 (N_9891,N_5914,N_7340);
and U9892 (N_9892,N_7388,N_6724);
and U9893 (N_9893,N_7064,N_6669);
and U9894 (N_9894,N_5945,N_6859);
nand U9895 (N_9895,N_6669,N_6899);
or U9896 (N_9896,N_6254,N_6807);
xor U9897 (N_9897,N_6083,N_6487);
or U9898 (N_9898,N_7110,N_7095);
nor U9899 (N_9899,N_5866,N_5326);
nand U9900 (N_9900,N_5417,N_5442);
and U9901 (N_9901,N_5256,N_7389);
or U9902 (N_9902,N_6410,N_6862);
and U9903 (N_9903,N_5513,N_7289);
nor U9904 (N_9904,N_5330,N_5107);
nand U9905 (N_9905,N_6220,N_6313);
and U9906 (N_9906,N_5618,N_5133);
xor U9907 (N_9907,N_5844,N_5842);
nand U9908 (N_9908,N_6121,N_5417);
and U9909 (N_9909,N_6205,N_6249);
nand U9910 (N_9910,N_6536,N_6942);
nand U9911 (N_9911,N_6635,N_6986);
nand U9912 (N_9912,N_7117,N_6749);
nor U9913 (N_9913,N_5599,N_6988);
or U9914 (N_9914,N_5376,N_7101);
nand U9915 (N_9915,N_6486,N_5234);
xnor U9916 (N_9916,N_5759,N_5304);
nor U9917 (N_9917,N_7261,N_6965);
or U9918 (N_9918,N_6416,N_5809);
nor U9919 (N_9919,N_6160,N_5760);
and U9920 (N_9920,N_6002,N_5777);
nor U9921 (N_9921,N_6296,N_6974);
and U9922 (N_9922,N_6022,N_5921);
nor U9923 (N_9923,N_7043,N_5453);
nor U9924 (N_9924,N_6759,N_7305);
or U9925 (N_9925,N_6061,N_5300);
nand U9926 (N_9926,N_5819,N_5132);
and U9927 (N_9927,N_5056,N_6327);
or U9928 (N_9928,N_5976,N_5542);
nor U9929 (N_9929,N_5345,N_5426);
nand U9930 (N_9930,N_6584,N_5336);
and U9931 (N_9931,N_7033,N_6473);
nand U9932 (N_9932,N_7159,N_6569);
nor U9933 (N_9933,N_7396,N_5192);
nand U9934 (N_9934,N_5315,N_5637);
nor U9935 (N_9935,N_6488,N_7285);
nand U9936 (N_9936,N_6705,N_5147);
or U9937 (N_9937,N_7053,N_6116);
or U9938 (N_9938,N_7297,N_7452);
nor U9939 (N_9939,N_6824,N_6677);
nand U9940 (N_9940,N_7250,N_5639);
nand U9941 (N_9941,N_5582,N_6147);
nor U9942 (N_9942,N_5314,N_6393);
and U9943 (N_9943,N_6018,N_6181);
nand U9944 (N_9944,N_6617,N_5460);
nand U9945 (N_9945,N_6177,N_6766);
nand U9946 (N_9946,N_7212,N_6740);
nor U9947 (N_9947,N_6546,N_6643);
nor U9948 (N_9948,N_7425,N_6024);
and U9949 (N_9949,N_6212,N_5902);
nand U9950 (N_9950,N_7186,N_5731);
nor U9951 (N_9951,N_5981,N_6453);
xnor U9952 (N_9952,N_5335,N_6762);
and U9953 (N_9953,N_6825,N_5859);
or U9954 (N_9954,N_5711,N_5991);
nand U9955 (N_9955,N_5310,N_6816);
nand U9956 (N_9956,N_6155,N_7237);
and U9957 (N_9957,N_6458,N_5326);
nand U9958 (N_9958,N_6733,N_6862);
nor U9959 (N_9959,N_6097,N_6614);
nand U9960 (N_9960,N_5376,N_6901);
nor U9961 (N_9961,N_6765,N_6436);
and U9962 (N_9962,N_5763,N_5878);
nor U9963 (N_9963,N_6838,N_6646);
nand U9964 (N_9964,N_6517,N_5796);
xor U9965 (N_9965,N_6000,N_6759);
nor U9966 (N_9966,N_6821,N_5945);
nand U9967 (N_9967,N_7429,N_7076);
nor U9968 (N_9968,N_5996,N_7025);
xnor U9969 (N_9969,N_5345,N_7239);
xor U9970 (N_9970,N_6584,N_6296);
nor U9971 (N_9971,N_6918,N_5726);
and U9972 (N_9972,N_5457,N_6093);
nor U9973 (N_9973,N_5872,N_6967);
nand U9974 (N_9974,N_7013,N_5415);
or U9975 (N_9975,N_6458,N_5450);
xnor U9976 (N_9976,N_5875,N_6284);
or U9977 (N_9977,N_6614,N_6803);
or U9978 (N_9978,N_6288,N_5927);
nor U9979 (N_9979,N_6054,N_7119);
and U9980 (N_9980,N_5785,N_7354);
and U9981 (N_9981,N_7282,N_5125);
or U9982 (N_9982,N_6084,N_5894);
nand U9983 (N_9983,N_5504,N_6616);
or U9984 (N_9984,N_5031,N_6097);
nand U9985 (N_9985,N_5078,N_5958);
and U9986 (N_9986,N_7497,N_7484);
nand U9987 (N_9987,N_6786,N_6158);
and U9988 (N_9988,N_5069,N_6702);
or U9989 (N_9989,N_5047,N_5809);
nor U9990 (N_9990,N_5306,N_6989);
nor U9991 (N_9991,N_5400,N_6112);
and U9992 (N_9992,N_6999,N_6236);
nand U9993 (N_9993,N_6303,N_5083);
nand U9994 (N_9994,N_5363,N_5634);
or U9995 (N_9995,N_5670,N_5867);
nand U9996 (N_9996,N_5194,N_7030);
and U9997 (N_9997,N_5599,N_6943);
or U9998 (N_9998,N_6540,N_5081);
or U9999 (N_9999,N_6083,N_6180);
nand UO_0 (O_0,N_8880,N_9319);
nor UO_1 (O_1,N_9686,N_9480);
or UO_2 (O_2,N_9427,N_7634);
and UO_3 (O_3,N_7824,N_9019);
nor UO_4 (O_4,N_9915,N_9815);
nand UO_5 (O_5,N_9360,N_8048);
nand UO_6 (O_6,N_9251,N_8052);
and UO_7 (O_7,N_7886,N_7922);
or UO_8 (O_8,N_8376,N_9781);
nand UO_9 (O_9,N_8711,N_7842);
xnor UO_10 (O_10,N_7846,N_7772);
nand UO_11 (O_11,N_7602,N_9637);
and UO_12 (O_12,N_8012,N_9991);
nor UO_13 (O_13,N_9266,N_7505);
or UO_14 (O_14,N_8783,N_9942);
xnor UO_15 (O_15,N_9627,N_9581);
xor UO_16 (O_16,N_7956,N_8175);
or UO_17 (O_17,N_8302,N_8737);
nand UO_18 (O_18,N_8490,N_7508);
xor UO_19 (O_19,N_8709,N_8437);
and UO_20 (O_20,N_9588,N_7542);
and UO_21 (O_21,N_8277,N_8982);
or UO_22 (O_22,N_9902,N_9587);
nand UO_23 (O_23,N_7896,N_8465);
or UO_24 (O_24,N_9458,N_7591);
or UO_25 (O_25,N_9344,N_9021);
or UO_26 (O_26,N_8295,N_8256);
or UO_27 (O_27,N_9534,N_7659);
and UO_28 (O_28,N_7798,N_7636);
nand UO_29 (O_29,N_7762,N_8249);
xor UO_30 (O_30,N_9394,N_9212);
and UO_31 (O_31,N_8863,N_7539);
or UO_32 (O_32,N_9105,N_8621);
nand UO_33 (O_33,N_9912,N_9625);
and UO_34 (O_34,N_8187,N_9530);
or UO_35 (O_35,N_8126,N_7708);
nand UO_36 (O_36,N_9146,N_7855);
nor UO_37 (O_37,N_8851,N_9052);
and UO_38 (O_38,N_7947,N_8733);
and UO_39 (O_39,N_7990,N_9846);
or UO_40 (O_40,N_7671,N_8518);
or UO_41 (O_41,N_7849,N_9432);
nor UO_42 (O_42,N_9058,N_9608);
nor UO_43 (O_43,N_9123,N_8955);
nand UO_44 (O_44,N_9579,N_9644);
or UO_45 (O_45,N_9658,N_7832);
and UO_46 (O_46,N_9434,N_9704);
or UO_47 (O_47,N_8207,N_9606);
xnor UO_48 (O_48,N_7519,N_8476);
nand UO_49 (O_49,N_8805,N_7581);
nor UO_50 (O_50,N_9059,N_8320);
and UO_51 (O_51,N_8576,N_8210);
and UO_52 (O_52,N_7700,N_8956);
nor UO_53 (O_53,N_9260,N_7517);
and UO_54 (O_54,N_9777,N_8875);
nand UO_55 (O_55,N_8753,N_8700);
and UO_56 (O_56,N_9814,N_7507);
nor UO_57 (O_57,N_8199,N_7993);
or UO_58 (O_58,N_7532,N_8230);
and UO_59 (O_59,N_8854,N_7652);
and UO_60 (O_60,N_8087,N_9366);
nand UO_61 (O_61,N_9927,N_7616);
and UO_62 (O_62,N_8767,N_8029);
or UO_63 (O_63,N_9520,N_9690);
and UO_64 (O_64,N_9693,N_8130);
nand UO_65 (O_65,N_8754,N_9538);
nor UO_66 (O_66,N_9092,N_9735);
nor UO_67 (O_67,N_9210,N_9167);
nor UO_68 (O_68,N_9916,N_7869);
or UO_69 (O_69,N_8962,N_9724);
or UO_70 (O_70,N_9555,N_9976);
xor UO_71 (O_71,N_8197,N_9208);
and UO_72 (O_72,N_8337,N_7523);
or UO_73 (O_73,N_7514,N_9727);
nor UO_74 (O_74,N_9160,N_7872);
nor UO_75 (O_75,N_8200,N_9609);
nand UO_76 (O_76,N_8185,N_9907);
or UO_77 (O_77,N_9221,N_7530);
or UO_78 (O_78,N_7687,N_9657);
or UO_79 (O_79,N_9411,N_7743);
and UO_80 (O_80,N_8608,N_8002);
or UO_81 (O_81,N_8685,N_8969);
xnor UO_82 (O_82,N_8074,N_7609);
nand UO_83 (O_83,N_7917,N_9115);
or UO_84 (O_84,N_8272,N_8995);
or UO_85 (O_85,N_9818,N_8707);
nand UO_86 (O_86,N_8375,N_8392);
nor UO_87 (O_87,N_8644,N_8368);
nand UO_88 (O_88,N_8591,N_9041);
or UO_89 (O_89,N_8109,N_8399);
and UO_90 (O_90,N_9946,N_8472);
and UO_91 (O_91,N_9447,N_9603);
nor UO_92 (O_92,N_9370,N_8104);
xor UO_93 (O_93,N_8744,N_7836);
xor UO_94 (O_94,N_8308,N_8022);
or UO_95 (O_95,N_9859,N_7590);
and UO_96 (O_96,N_8228,N_8484);
nor UO_97 (O_97,N_8931,N_9514);
nor UO_98 (O_98,N_8887,N_8263);
nor UO_99 (O_99,N_7538,N_9340);
nor UO_100 (O_100,N_8730,N_7510);
nor UO_101 (O_101,N_7870,N_7715);
xnor UO_102 (O_102,N_9300,N_8575);
or UO_103 (O_103,N_8936,N_8192);
and UO_104 (O_104,N_8920,N_9599);
nor UO_105 (O_105,N_8373,N_9073);
and UO_106 (O_106,N_9051,N_8541);
and UO_107 (O_107,N_8403,N_8319);
nor UO_108 (O_108,N_7978,N_8351);
xor UO_109 (O_109,N_8362,N_8856);
xnor UO_110 (O_110,N_8423,N_9793);
xnor UO_111 (O_111,N_8543,N_8118);
nand UO_112 (O_112,N_7705,N_7728);
nand UO_113 (O_113,N_9275,N_8299);
nor UO_114 (O_114,N_9496,N_8301);
or UO_115 (O_115,N_8911,N_9978);
nor UO_116 (O_116,N_8757,N_8326);
xnor UO_117 (O_117,N_9114,N_7768);
or UO_118 (O_118,N_8840,N_9591);
xnor UO_119 (O_119,N_9033,N_8238);
or UO_120 (O_120,N_7500,N_8222);
nand UO_121 (O_121,N_9756,N_9362);
nand UO_122 (O_122,N_8512,N_8958);
or UO_123 (O_123,N_9085,N_7977);
and UO_124 (O_124,N_9631,N_9699);
and UO_125 (O_125,N_8824,N_8629);
nor UO_126 (O_126,N_9175,N_8158);
or UO_127 (O_127,N_9833,N_7518);
nand UO_128 (O_128,N_8689,N_9656);
or UO_129 (O_129,N_7904,N_7674);
or UO_130 (O_130,N_7533,N_8105);
and UO_131 (O_131,N_7620,N_9101);
or UO_132 (O_132,N_9144,N_8164);
or UO_133 (O_133,N_8154,N_7724);
and UO_134 (O_134,N_9437,N_7516);
nor UO_135 (O_135,N_8357,N_9526);
nand UO_136 (O_136,N_9542,N_9905);
and UO_137 (O_137,N_8204,N_8620);
and UO_138 (O_138,N_9967,N_8823);
xor UO_139 (O_139,N_9225,N_9650);
nand UO_140 (O_140,N_9087,N_8945);
nor UO_141 (O_141,N_9107,N_8546);
nor UO_142 (O_142,N_7559,N_9182);
and UO_143 (O_143,N_8129,N_9855);
and UO_144 (O_144,N_8452,N_8719);
nand UO_145 (O_145,N_9013,N_7828);
and UO_146 (O_146,N_9474,N_9363);
and UO_147 (O_147,N_8374,N_8852);
nor UO_148 (O_148,N_8567,N_9931);
and UO_149 (O_149,N_9361,N_8128);
or UO_150 (O_150,N_7695,N_8183);
and UO_151 (O_151,N_8015,N_9575);
nand UO_152 (O_152,N_9749,N_8745);
or UO_153 (O_153,N_9076,N_9632);
nand UO_154 (O_154,N_9888,N_8321);
nor UO_155 (O_155,N_9497,N_7521);
or UO_156 (O_156,N_8798,N_9492);
or UO_157 (O_157,N_8897,N_9849);
or UO_158 (O_158,N_9418,N_9977);
nor UO_159 (O_159,N_7574,N_9238);
and UO_160 (O_160,N_9601,N_7604);
and UO_161 (O_161,N_8669,N_9446);
or UO_162 (O_162,N_9265,N_8985);
xor UO_163 (O_163,N_9816,N_9126);
nand UO_164 (O_164,N_8696,N_8214);
and UO_165 (O_165,N_9232,N_8957);
nor UO_166 (O_166,N_9923,N_9359);
nand UO_167 (O_167,N_7610,N_9342);
or UO_168 (O_168,N_8511,N_8708);
nand UO_169 (O_169,N_8485,N_7997);
nor UO_170 (O_170,N_9537,N_9436);
and UO_171 (O_171,N_9292,N_8035);
or UO_172 (O_172,N_7873,N_9765);
or UO_173 (O_173,N_9148,N_7885);
nor UO_174 (O_174,N_7642,N_8280);
nor UO_175 (O_175,N_8626,N_8628);
and UO_176 (O_176,N_8281,N_7918);
and UO_177 (O_177,N_8503,N_7792);
xor UO_178 (O_178,N_8358,N_7627);
or UO_179 (O_179,N_9773,N_7723);
nand UO_180 (O_180,N_9722,N_8789);
nor UO_181 (O_181,N_8092,N_7913);
nor UO_182 (O_182,N_9909,N_9270);
and UO_183 (O_183,N_8180,N_8554);
or UO_184 (O_184,N_8324,N_9760);
nand UO_185 (O_185,N_7683,N_8435);
nand UO_186 (O_186,N_9435,N_9847);
and UO_187 (O_187,N_8089,N_8998);
nand UO_188 (O_188,N_8542,N_7862);
nand UO_189 (O_189,N_9832,N_9757);
nor UO_190 (O_190,N_7761,N_9889);
nand UO_191 (O_191,N_9498,N_8217);
and UO_192 (O_192,N_9250,N_8966);
nand UO_193 (O_193,N_8746,N_8501);
and UO_194 (O_194,N_9896,N_7564);
nor UO_195 (O_195,N_8194,N_8066);
xnor UO_196 (O_196,N_8410,N_7621);
nand UO_197 (O_197,N_9307,N_9830);
nor UO_198 (O_198,N_7709,N_9471);
or UO_199 (O_199,N_8534,N_8876);
xor UO_200 (O_200,N_8869,N_9594);
nor UO_201 (O_201,N_8136,N_8046);
or UO_202 (O_202,N_8836,N_8287);
xor UO_203 (O_203,N_7554,N_9679);
and UO_204 (O_204,N_9367,N_8391);
or UO_205 (O_205,N_8994,N_8344);
or UO_206 (O_206,N_9928,N_8318);
nand UO_207 (O_207,N_8095,N_9120);
and UO_208 (O_208,N_7866,N_9844);
or UO_209 (O_209,N_9091,N_7607);
and UO_210 (O_210,N_7580,N_8273);
or UO_211 (O_211,N_9968,N_9950);
xor UO_212 (O_212,N_8528,N_9157);
and UO_213 (O_213,N_9553,N_9416);
nor UO_214 (O_214,N_8811,N_8504);
nand UO_215 (O_215,N_8563,N_9046);
nor UO_216 (O_216,N_9023,N_7865);
and UO_217 (O_217,N_8532,N_9166);
nand UO_218 (O_218,N_9487,N_7942);
and UO_219 (O_219,N_7596,N_9719);
or UO_220 (O_220,N_7688,N_8160);
nand UO_221 (O_221,N_9378,N_9505);
or UO_222 (O_222,N_8986,N_9034);
nand UO_223 (O_223,N_9053,N_8860);
nor UO_224 (O_224,N_7511,N_8247);
and UO_225 (O_225,N_7553,N_9673);
and UO_226 (O_226,N_8349,N_9209);
and UO_227 (O_227,N_9569,N_8414);
and UO_228 (O_228,N_7890,N_9503);
nor UO_229 (O_229,N_9116,N_7676);
and UO_230 (O_230,N_9834,N_7984);
and UO_231 (O_231,N_9429,N_7880);
and UO_232 (O_232,N_7910,N_7868);
and UO_233 (O_233,N_9707,N_9702);
or UO_234 (O_234,N_9242,N_8602);
or UO_235 (O_235,N_9277,N_9348);
nor UO_236 (O_236,N_9334,N_9419);
nand UO_237 (O_237,N_8115,N_9532);
nor UO_238 (O_238,N_7879,N_9188);
nor UO_239 (O_239,N_9140,N_9294);
and UO_240 (O_240,N_9223,N_9353);
nor UO_241 (O_241,N_9003,N_8143);
nand UO_242 (O_242,N_8397,N_7812);
or UO_243 (O_243,N_7887,N_8579);
nor UO_244 (O_244,N_7839,N_8728);
xor UO_245 (O_245,N_8792,N_8710);
or UO_246 (O_246,N_7637,N_8146);
and UO_247 (O_247,N_8270,N_8455);
xor UO_248 (O_248,N_8582,N_7949);
nand UO_249 (O_249,N_9835,N_8383);
and UO_250 (O_250,N_9689,N_8517);
or UO_251 (O_251,N_7502,N_9808);
nand UO_252 (O_252,N_8334,N_9320);
and UO_253 (O_253,N_9372,N_8965);
or UO_254 (O_254,N_8475,N_8699);
and UO_255 (O_255,N_7934,N_8165);
or UO_256 (O_256,N_9778,N_7749);
or UO_257 (O_257,N_9668,N_8742);
or UO_258 (O_258,N_8269,N_8429);
nor UO_259 (O_259,N_8097,N_9162);
and UO_260 (O_260,N_8463,N_7791);
and UO_261 (O_261,N_8583,N_7701);
xor UO_262 (O_262,N_9231,N_7623);
nor UO_263 (O_263,N_9128,N_9990);
or UO_264 (O_264,N_7883,N_7830);
nand UO_265 (O_265,N_9473,N_9462);
and UO_266 (O_266,N_9568,N_8186);
nor UO_267 (O_267,N_8330,N_8433);
or UO_268 (O_268,N_7874,N_9676);
nor UO_269 (O_269,N_7789,N_9386);
or UO_270 (O_270,N_8794,N_9851);
nand UO_271 (O_271,N_9999,N_9876);
nand UO_272 (O_272,N_8682,N_9864);
nand UO_273 (O_273,N_7650,N_9753);
or UO_274 (O_274,N_9891,N_9020);
nand UO_275 (O_275,N_8874,N_9789);
nand UO_276 (O_276,N_7905,N_8890);
nor UO_277 (O_277,N_8573,N_7794);
or UO_278 (O_278,N_8428,N_7631);
nand UO_279 (O_279,N_8963,N_9333);
and UO_280 (O_280,N_8834,N_9549);
and UO_281 (O_281,N_7527,N_9110);
nand UO_282 (O_282,N_8866,N_7649);
or UO_283 (O_283,N_7857,N_9806);
nand UO_284 (O_284,N_9438,N_9797);
or UO_285 (O_285,N_8359,N_7878);
and UO_286 (O_286,N_8350,N_9626);
or UO_287 (O_287,N_9878,N_7919);
or UO_288 (O_288,N_8690,N_9868);
nor UO_289 (O_289,N_9649,N_9567);
or UO_290 (O_290,N_8979,N_9564);
nand UO_291 (O_291,N_9352,N_8515);
and UO_292 (O_292,N_8076,N_9562);
or UO_293 (O_293,N_9820,N_9718);
nand UO_294 (O_294,N_8693,N_9397);
nor UO_295 (O_295,N_8044,N_7888);
nand UO_296 (O_296,N_9468,N_9129);
or UO_297 (O_297,N_8915,N_8014);
and UO_298 (O_298,N_8293,N_7766);
nand UO_299 (O_299,N_7987,N_8721);
and UO_300 (O_300,N_8818,N_9421);
nand UO_301 (O_301,N_8549,N_7658);
or UO_302 (O_302,N_9994,N_7531);
nor UO_303 (O_303,N_9399,N_8325);
and UO_304 (O_304,N_8364,N_8960);
nand UO_305 (O_305,N_8905,N_8658);
or UO_306 (O_306,N_8174,N_7966);
or UO_307 (O_307,N_8676,N_7786);
and UO_308 (O_308,N_7657,N_8071);
nor UO_309 (O_309,N_8973,N_9170);
and UO_310 (O_310,N_8625,N_9713);
and UO_311 (O_311,N_8533,N_9593);
nor UO_312 (O_312,N_8347,N_7776);
nand UO_313 (O_313,N_9596,N_9404);
nor UO_314 (O_314,N_8918,N_9893);
nand UO_315 (O_315,N_8303,N_9449);
nand UO_316 (O_316,N_8883,N_7867);
xor UO_317 (O_317,N_8891,N_8152);
or UO_318 (O_318,N_9181,N_9374);
xnor UO_319 (O_319,N_9130,N_7781);
or UO_320 (O_320,N_7967,N_8884);
xnor UO_321 (O_321,N_8677,N_7736);
or UO_322 (O_322,N_9848,N_9379);
nor UO_323 (O_323,N_8903,N_8121);
nor UO_324 (O_324,N_9748,N_7814);
nand UO_325 (O_325,N_8906,N_9234);
and UO_326 (O_326,N_9580,N_9222);
nand UO_327 (O_327,N_7600,N_8372);
and UO_328 (O_328,N_9484,N_9630);
nand UO_329 (O_329,N_7572,N_8929);
or UO_330 (O_330,N_7503,N_9299);
or UO_331 (O_331,N_8073,N_9618);
nor UO_332 (O_332,N_8479,N_9764);
xor UO_333 (O_333,N_8234,N_8723);
and UO_334 (O_334,N_9867,N_9281);
nand UO_335 (O_335,N_9393,N_7703);
and UO_336 (O_336,N_8913,N_7906);
and UO_337 (O_337,N_9733,N_8348);
or UO_338 (O_338,N_9743,N_8494);
and UO_339 (O_339,N_9671,N_9346);
xor UO_340 (O_340,N_8999,N_8288);
nor UO_341 (O_341,N_8952,N_7854);
nand UO_342 (O_342,N_9108,N_9813);
or UO_343 (O_343,N_8134,N_9457);
nor UO_344 (O_344,N_8027,N_8790);
nor UO_345 (O_345,N_8108,N_8064);
nand UO_346 (O_346,N_9736,N_8806);
nand UO_347 (O_347,N_7656,N_8246);
and UO_348 (O_348,N_8933,N_9422);
xnor UO_349 (O_349,N_8773,N_7968);
nand UO_350 (O_350,N_8233,N_9089);
and UO_351 (O_351,N_8361,N_8729);
nor UO_352 (O_352,N_9973,N_8694);
nor UO_353 (O_353,N_9924,N_8497);
nor UO_354 (O_354,N_8294,N_9259);
nand UO_355 (O_355,N_9758,N_7617);
xor UO_356 (O_356,N_8785,N_9708);
and UO_357 (O_357,N_8003,N_9226);
or UO_358 (O_358,N_9290,N_7624);
xnor UO_359 (O_359,N_8117,N_9911);
nand UO_360 (O_360,N_7647,N_7838);
nor UO_361 (O_361,N_9358,N_8764);
or UO_362 (O_362,N_8864,N_8007);
nor UO_363 (O_363,N_8650,N_9621);
nor UO_364 (O_364,N_8535,N_8271);
or UO_365 (O_365,N_9774,N_8502);
or UO_366 (O_366,N_7686,N_8923);
or UO_367 (O_367,N_8236,N_8144);
nor UO_368 (O_368,N_9804,N_9515);
and UO_369 (O_369,N_7663,N_8587);
or UO_370 (O_370,N_8695,N_9612);
or UO_371 (O_371,N_7944,N_9104);
or UO_372 (O_372,N_9857,N_8093);
xor UO_373 (O_373,N_8774,N_7809);
nand UO_374 (O_374,N_9957,N_9272);
and UO_375 (O_375,N_8436,N_8081);
and UO_376 (O_376,N_8120,N_8045);
and UO_377 (O_377,N_7744,N_9527);
or UO_378 (O_378,N_9391,N_8861);
nand UO_379 (O_379,N_9850,N_9694);
nor UO_380 (O_380,N_9246,N_8356);
nor UO_381 (O_381,N_9682,N_9099);
xnor UO_382 (O_382,N_9750,N_8981);
or UO_383 (O_383,N_7936,N_7588);
and UO_384 (O_384,N_8306,N_8259);
or UO_385 (O_385,N_8407,N_8379);
nor UO_386 (O_386,N_8190,N_7907);
or UO_387 (O_387,N_8566,N_9218);
and UO_388 (O_388,N_8371,N_9783);
nand UO_389 (O_389,N_8808,N_9405);
or UO_390 (O_390,N_7512,N_7690);
nor UO_391 (O_391,N_9584,N_8849);
xnor UO_392 (O_392,N_8396,N_8795);
or UO_393 (O_393,N_8980,N_9825);
nand UO_394 (O_394,N_9414,N_9018);
and UO_395 (O_395,N_9295,N_8645);
and UO_396 (O_396,N_9009,N_8099);
nand UO_397 (O_397,N_9563,N_9680);
nor UO_398 (O_398,N_9965,N_8031);
and UO_399 (O_399,N_9877,N_8545);
xor UO_400 (O_400,N_8151,N_7802);
and UO_401 (O_401,N_7679,N_8340);
and UO_402 (O_402,N_9293,N_7745);
nor UO_403 (O_403,N_9354,N_9728);
or UO_404 (O_404,N_7951,N_9088);
nor UO_405 (O_405,N_9066,N_7681);
and UO_406 (O_406,N_9745,N_9881);
and UO_407 (O_407,N_8637,N_7793);
nand UO_408 (O_408,N_9486,N_9604);
nand UO_409 (O_409,N_9516,N_8613);
nor UO_410 (O_410,N_9661,N_8859);
or UO_411 (O_411,N_7628,N_8385);
nand UO_412 (O_412,N_8937,N_9169);
nor UO_413 (O_413,N_7784,N_8972);
nor UO_414 (O_414,N_7654,N_8668);
nand UO_415 (O_415,N_7726,N_8848);
nand UO_416 (O_416,N_9706,N_9838);
and UO_417 (O_417,N_7833,N_7739);
nor UO_418 (O_418,N_7754,N_8345);
and UO_419 (O_419,N_9112,N_9064);
nand UO_420 (O_420,N_8569,N_8691);
or UO_421 (O_421,N_9959,N_8219);
nor UO_422 (O_422,N_7861,N_7982);
nand UO_423 (O_423,N_9636,N_7999);
or UO_424 (O_424,N_9356,N_9080);
or UO_425 (O_425,N_8529,N_7928);
or UO_426 (O_426,N_7950,N_8323);
nor UO_427 (O_427,N_7589,N_7645);
nand UO_428 (O_428,N_9096,N_9910);
and UO_429 (O_429,N_7528,N_8060);
xnor UO_430 (O_430,N_8950,N_8725);
nand UO_431 (O_431,N_7957,N_8850);
and UO_432 (O_432,N_9629,N_8291);
and UO_433 (O_433,N_9552,N_9106);
nor UO_434 (O_434,N_7567,N_8057);
nand UO_435 (O_435,N_9303,N_7955);
nor UO_436 (O_436,N_7815,N_9995);
nor UO_437 (O_437,N_9856,N_9925);
nor UO_438 (O_438,N_8008,N_7711);
nor UO_439 (O_439,N_9504,N_8283);
nor UO_440 (O_440,N_9577,N_7763);
nand UO_441 (O_441,N_8801,N_9841);
and UO_442 (O_442,N_8810,N_8862);
xnor UO_443 (O_443,N_8611,N_8701);
nand UO_444 (O_444,N_8341,N_7780);
or UO_445 (O_445,N_9006,N_8211);
or UO_446 (O_446,N_8469,N_7731);
nor UO_447 (O_447,N_9180,N_7980);
nand UO_448 (O_448,N_9351,N_8716);
nor UO_449 (O_449,N_7719,N_9817);
nand UO_450 (O_450,N_7613,N_8033);
xnor UO_451 (O_451,N_9842,N_7795);
nor UO_452 (O_452,N_9684,N_8432);
xnor UO_453 (O_453,N_9141,N_8736);
nor UO_454 (O_454,N_9944,N_8202);
and UO_455 (O_455,N_7626,N_9535);
and UO_456 (O_456,N_9075,N_8482);
xor UO_457 (O_457,N_9616,N_9477);
and UO_458 (O_458,N_9309,N_8732);
and UO_459 (O_459,N_8935,N_9664);
nand UO_460 (O_460,N_9558,N_8766);
nand UO_461 (O_461,N_9173,N_9079);
or UO_462 (O_462,N_9517,N_9895);
or UO_463 (O_463,N_7691,N_8527);
nor UO_464 (O_464,N_7525,N_8360);
and UO_465 (O_465,N_9213,N_8991);
nand UO_466 (O_466,N_9752,N_8643);
nor UO_467 (O_467,N_8760,N_9547);
and UO_468 (O_468,N_8687,N_7660);
nor UO_469 (O_469,N_7562,N_7779);
nand UO_470 (O_470,N_8775,N_9559);
and UO_471 (O_471,N_7742,N_9461);
or UO_472 (O_472,N_7756,N_8313);
nand UO_473 (O_473,N_9521,N_9714);
nand UO_474 (O_474,N_9768,N_9775);
and UO_475 (O_475,N_8235,N_8844);
nor UO_476 (O_476,N_9464,N_7875);
nor UO_477 (O_477,N_8201,N_8342);
or UO_478 (O_478,N_8227,N_8561);
xnor UO_479 (O_479,N_9103,N_8315);
nand UO_480 (O_480,N_8009,N_7773);
or UO_481 (O_481,N_8830,N_7770);
and UO_482 (O_482,N_9971,N_7557);
nor UO_483 (O_483,N_8899,N_7790);
nor UO_484 (O_484,N_8286,N_8928);
nor UO_485 (O_485,N_7550,N_7926);
nor UO_486 (O_486,N_8605,N_7785);
xor UO_487 (O_487,N_9192,N_8132);
and UO_488 (O_488,N_7829,N_9385);
and UO_489 (O_489,N_7900,N_7569);
nand UO_490 (O_490,N_9952,N_8352);
and UO_491 (O_491,N_7666,N_8697);
or UO_492 (O_492,N_8892,N_8404);
nor UO_493 (O_493,N_7587,N_9620);
nand UO_494 (O_494,N_9426,N_8713);
or UO_495 (O_495,N_9565,N_8505);
or UO_496 (O_496,N_8193,N_9171);
or UO_497 (O_497,N_7994,N_8635);
nor UO_498 (O_498,N_9002,N_7661);
and UO_499 (O_499,N_9413,N_8267);
nand UO_500 (O_500,N_8943,N_9219);
nor UO_501 (O_501,N_8080,N_9135);
nor UO_502 (O_502,N_8577,N_7689);
and UO_503 (O_503,N_9077,N_7767);
nor UO_504 (O_504,N_8274,N_9744);
or UO_505 (O_505,N_9328,N_8843);
xnor UO_506 (O_506,N_9685,N_8419);
nor UO_507 (O_507,N_7816,N_8179);
nand UO_508 (O_508,N_8593,N_8477);
or UO_509 (O_509,N_7976,N_7561);
or UO_510 (O_510,N_8380,N_8409);
nand UO_511 (O_511,N_7845,N_9335);
nand UO_512 (O_512,N_8817,N_8223);
nor UO_513 (O_513,N_8251,N_9015);
nor UO_514 (O_514,N_9642,N_8447);
and UO_515 (O_515,N_8879,N_9518);
nor UO_516 (O_516,N_9945,N_9139);
nor UO_517 (O_517,N_8393,N_9502);
nand UO_518 (O_518,N_7668,N_8872);
or UO_519 (O_519,N_7892,N_9189);
nand UO_520 (O_520,N_9044,N_8067);
or UO_521 (O_521,N_9132,N_9150);
nor UO_522 (O_522,N_8453,N_8420);
and UO_523 (O_523,N_8055,N_9669);
and UO_524 (O_524,N_8406,N_7605);
nor UO_525 (O_525,N_8026,N_9406);
or UO_526 (O_526,N_9381,N_9786);
or UO_527 (O_527,N_7548,N_8655);
nor UO_528 (O_528,N_8565,N_8917);
nand UO_529 (O_529,N_9528,N_8522);
nor UO_530 (O_530,N_9330,N_8103);
nand UO_531 (O_531,N_8594,N_9698);
nor UO_532 (O_532,N_9133,N_9283);
and UO_533 (O_533,N_8042,N_7710);
nor UO_534 (O_534,N_8405,N_7813);
nor UO_535 (O_535,N_8809,N_8498);
nor UO_536 (O_536,N_9955,N_9355);
nand UO_537 (O_537,N_9985,N_8984);
nor UO_538 (O_538,N_9322,N_7684);
and UO_539 (O_539,N_9751,N_8756);
and UO_540 (O_540,N_9903,N_9382);
or UO_541 (O_541,N_7541,N_8139);
nor UO_542 (O_542,N_9828,N_7592);
and UO_543 (O_543,N_7823,N_9176);
and UO_544 (O_544,N_9183,N_9741);
or UO_545 (O_545,N_8262,N_7852);
and UO_546 (O_546,N_8833,N_7902);
nand UO_547 (O_547,N_8604,N_8954);
nand UO_548 (O_548,N_9495,N_9341);
nand UO_549 (O_549,N_8221,N_7536);
or UO_550 (O_550,N_9441,N_9048);
nand UO_551 (O_551,N_9628,N_9324);
or UO_552 (O_552,N_8156,N_9081);
or UO_553 (O_553,N_8040,N_7757);
and UO_554 (O_554,N_7765,N_7669);
or UO_555 (O_555,N_7706,N_7840);
and UO_556 (O_556,N_8241,N_8752);
xor UO_557 (O_557,N_9121,N_8226);
nand UO_558 (O_558,N_8858,N_8133);
and UO_559 (O_559,N_7974,N_7943);
nand UO_560 (O_560,N_8603,N_7535);
and UO_561 (O_561,N_9501,N_9701);
nor UO_562 (O_562,N_7787,N_8032);
nand UO_563 (O_563,N_8855,N_9055);
xnor UO_564 (O_564,N_9245,N_7625);
or UO_565 (O_565,N_8148,N_7629);
and UO_566 (O_566,N_9769,N_8740);
nand UO_567 (O_567,N_9423,N_8720);
or UO_568 (O_568,N_8556,N_9983);
nand UO_569 (O_569,N_9926,N_9711);
or UO_570 (O_570,N_8135,N_7643);
nand UO_571 (O_571,N_8781,N_9090);
or UO_572 (O_572,N_9453,N_9936);
nor UO_573 (O_573,N_7544,N_8336);
and UO_574 (O_574,N_9998,N_7717);
xnor UO_575 (O_575,N_7964,N_8666);
nor UO_576 (O_576,N_7863,N_9879);
and UO_577 (O_577,N_8425,N_8084);
nand UO_578 (O_578,N_8590,N_7915);
or UO_579 (O_579,N_7635,N_8237);
nand UO_580 (O_580,N_7925,N_8034);
xor UO_581 (O_581,N_7734,N_9763);
nor UO_582 (O_582,N_8431,N_9024);
xor UO_583 (O_583,N_9964,N_8001);
nand UO_584 (O_584,N_7841,N_9710);
and UO_585 (O_585,N_8938,N_7667);
nand UO_586 (O_586,N_8846,N_7556);
nor UO_587 (O_587,N_9001,N_8167);
and UO_588 (O_588,N_9239,N_8119);
nor UO_589 (O_589,N_8623,N_8714);
or UO_590 (O_590,N_9310,N_8705);
nor UO_591 (O_591,N_7799,N_8717);
and UO_592 (O_592,N_7665,N_9403);
or UO_593 (O_593,N_9920,N_8459);
or UO_594 (O_594,N_8153,N_7558);
and UO_595 (O_595,N_8908,N_9331);
nand UO_596 (O_596,N_8053,N_7639);
nand UO_597 (O_597,N_8726,N_7638);
nor UO_598 (O_598,N_8328,N_7932);
or UO_599 (O_599,N_9483,N_9119);
or UO_600 (O_600,N_7764,N_9651);
and UO_601 (O_601,N_9493,N_8028);
xnor UO_602 (O_602,N_7702,N_8460);
nor UO_603 (O_603,N_8377,N_9969);
and UO_604 (O_604,N_9155,N_8877);
nand UO_605 (O_605,N_9415,N_7912);
nand UO_606 (O_606,N_9791,N_8282);
or UO_607 (O_607,N_8050,N_9984);
and UO_608 (O_608,N_9400,N_7575);
or UO_609 (O_609,N_8678,N_8090);
nor UO_610 (O_610,N_8589,N_7526);
nor UO_611 (O_611,N_8131,N_9919);
nand UO_612 (O_612,N_9819,N_9068);
nand UO_613 (O_613,N_8471,N_9980);
or UO_614 (O_614,N_9312,N_7971);
nand UO_615 (O_615,N_9276,N_9665);
xnor UO_616 (O_616,N_8088,N_9262);
nor UO_617 (O_617,N_8665,N_9729);
xnor UO_618 (O_618,N_8524,N_8261);
or UO_619 (O_619,N_8997,N_8434);
or UO_620 (O_620,N_8647,N_7537);
nor UO_621 (O_621,N_7633,N_9932);
nand UO_622 (O_622,N_8769,N_8025);
nor UO_623 (O_623,N_7992,N_8536);
and UO_624 (O_624,N_8513,N_9198);
nand UO_625 (O_625,N_7834,N_8389);
nand UO_626 (O_626,N_9043,N_8967);
and UO_627 (O_627,N_9993,N_8365);
nor UO_628 (O_628,N_8307,N_8332);
nor UO_629 (O_629,N_9301,N_7608);
nor UO_630 (O_630,N_8530,N_9913);
and UO_631 (O_631,N_8889,N_9541);
and UO_632 (O_632,N_9904,N_9659);
and UO_633 (O_633,N_9953,N_9574);
and UO_634 (O_634,N_8290,N_9573);
and UO_635 (O_635,N_7871,N_8615);
nor UO_636 (O_636,N_7672,N_9014);
nand UO_637 (O_637,N_8662,N_9038);
and UO_638 (O_638,N_8675,N_9070);
nor UO_639 (O_639,N_8616,N_7920);
or UO_640 (O_640,N_7775,N_8111);
xnor UO_641 (O_641,N_8487,N_9611);
nor UO_642 (O_642,N_7945,N_7595);
xnor UO_643 (O_643,N_7758,N_9605);
and UO_644 (O_644,N_8597,N_9554);
or UO_645 (O_645,N_8581,N_9963);
or UO_646 (O_646,N_8570,N_7963);
nand UO_647 (O_647,N_8101,N_8762);
nor UO_648 (O_648,N_9084,N_9417);
nor UO_649 (O_649,N_9705,N_7826);
nor UO_650 (O_650,N_9576,N_9313);
nand UO_651 (O_651,N_9204,N_8870);
or UO_652 (O_652,N_7782,N_8091);
nor UO_653 (O_653,N_7655,N_9884);
or UO_654 (O_654,N_8229,N_8150);
nor UO_655 (O_655,N_7718,N_9633);
xnor UO_656 (O_656,N_7953,N_8614);
nand UO_657 (O_657,N_9163,N_8782);
and UO_658 (O_658,N_9784,N_8553);
nand UO_659 (O_659,N_9958,N_8592);
nor UO_660 (O_660,N_9199,N_9185);
and UO_661 (O_661,N_9866,N_7583);
xnor UO_662 (O_662,N_8141,N_9653);
and UO_663 (O_663,N_7699,N_9589);
and UO_664 (O_664,N_8704,N_9648);
nor UO_665 (O_665,N_9345,N_9249);
nor UO_666 (O_666,N_8755,N_9887);
xnor UO_667 (O_667,N_7969,N_7820);
or UO_668 (O_668,N_7819,N_9460);
and UO_669 (O_669,N_9578,N_8831);
and UO_670 (O_670,N_9289,N_8547);
and UO_671 (O_671,N_9966,N_8322);
and UO_672 (O_672,N_9057,N_7565);
and UO_673 (O_673,N_9007,N_8243);
or UO_674 (O_674,N_8454,N_7696);
or UO_675 (O_675,N_7801,N_8402);
or UO_676 (O_676,N_7952,N_7612);
or UO_677 (O_677,N_9016,N_8049);
or UO_678 (O_678,N_8902,N_9635);
and UO_679 (O_679,N_9687,N_9854);
or UO_680 (O_680,N_7716,N_9428);
or UO_681 (O_681,N_7851,N_8017);
and UO_682 (O_682,N_8005,N_9224);
or UO_683 (O_683,N_9570,N_8191);
and UO_684 (O_684,N_7891,N_9060);
xnor UO_685 (O_685,N_9450,N_9329);
or UO_686 (O_686,N_9220,N_9615);
nor UO_687 (O_687,N_9083,N_9264);
xor UO_688 (O_688,N_8548,N_7520);
and UO_689 (O_689,N_9196,N_7504);
nand UO_690 (O_690,N_8398,N_9738);
nor UO_691 (O_691,N_8595,N_7680);
or UO_692 (O_692,N_9901,N_9398);
or UO_693 (O_693,N_8692,N_9882);
and UO_694 (O_694,N_8633,N_8260);
or UO_695 (O_695,N_9662,N_8242);
nor UO_696 (O_696,N_9045,N_8255);
nand UO_697 (O_697,N_9174,N_8638);
nand UO_698 (O_698,N_8763,N_7555);
and UO_699 (O_699,N_8619,N_9767);
and UO_700 (O_700,N_8948,N_9158);
nor UO_701 (O_701,N_9142,N_7741);
xor UO_702 (O_702,N_9646,N_9491);
nor UO_703 (O_703,N_9439,N_9470);
or UO_704 (O_704,N_8268,N_9805);
xor UO_705 (O_705,N_9478,N_8651);
or UO_706 (O_706,N_8250,N_8684);
and UO_707 (O_707,N_8715,N_9194);
xor UO_708 (O_708,N_8122,N_9005);
and UO_709 (O_709,N_8642,N_9287);
or UO_710 (O_710,N_9149,N_8559);
or UO_711 (O_711,N_9472,N_9102);
nand UO_712 (O_712,N_7931,N_9683);
nand UO_713 (O_713,N_8378,N_7962);
or UO_714 (O_714,N_7941,N_8041);
or UO_715 (O_715,N_8944,N_8069);
and UO_716 (O_716,N_8445,N_8671);
and UO_717 (O_717,N_9256,N_9590);
xnor UO_718 (O_718,N_7921,N_8514);
or UO_719 (O_719,N_8456,N_8748);
and UO_720 (O_720,N_8114,N_9771);
nor UO_721 (O_721,N_8750,N_9444);
or UO_722 (O_722,N_9566,N_8942);
and UO_723 (O_723,N_9430,N_7935);
or UO_724 (O_724,N_8568,N_7948);
nor UO_725 (O_725,N_8653,N_8670);
xor UO_726 (O_726,N_8660,N_9479);
and UO_727 (O_727,N_7707,N_9766);
nand UO_728 (O_728,N_7939,N_8927);
and UO_729 (O_729,N_8300,N_7881);
or UO_730 (O_730,N_8770,N_8343);
or UO_731 (O_731,N_8727,N_9723);
and UO_732 (O_732,N_8181,N_7972);
and UO_733 (O_733,N_8314,N_9047);
nor UO_734 (O_734,N_9782,N_7698);
nand UO_735 (O_735,N_9852,N_8971);
nor UO_736 (O_736,N_9996,N_8279);
nand UO_737 (O_737,N_7946,N_8438);
and UO_738 (O_738,N_9643,N_8632);
xnor UO_739 (O_739,N_8674,N_7970);
and UO_740 (O_740,N_9717,N_8304);
or UO_741 (O_741,N_8196,N_8468);
nor UO_742 (O_742,N_7882,N_8857);
nor UO_743 (O_743,N_7697,N_8363);
or UO_744 (O_744,N_9696,N_8483);
nor UO_745 (O_745,N_8523,N_9371);
xor UO_746 (O_746,N_8988,N_7755);
nand UO_747 (O_747,N_8083,N_9795);
nor UO_748 (O_748,N_8641,N_9655);
nor UO_749 (O_749,N_8925,N_8895);
and UO_750 (O_750,N_9207,N_9858);
or UO_751 (O_751,N_7778,N_7929);
xor UO_752 (O_752,N_9211,N_9153);
nor UO_753 (O_753,N_8312,N_9244);
nand UO_754 (O_754,N_8072,N_9551);
or UO_755 (O_755,N_7805,N_9305);
xnor UO_756 (O_756,N_7747,N_9408);
xnor UO_757 (O_757,N_8799,N_9347);
xor UO_758 (O_758,N_9762,N_9396);
and UO_759 (O_759,N_8683,N_8835);
or UO_760 (O_760,N_9754,N_8248);
and UO_761 (O_761,N_8292,N_9357);
nor UO_762 (O_762,N_9523,N_9557);
xor UO_763 (O_763,N_8170,N_8688);
and UO_764 (O_764,N_7817,N_8886);
nor UO_765 (O_765,N_9215,N_9237);
and UO_766 (O_766,N_8430,N_9004);
and UO_767 (O_767,N_8257,N_9248);
or UO_768 (O_768,N_8622,N_8169);
nor UO_769 (O_769,N_8310,N_9869);
and UO_770 (O_770,N_9890,N_9829);
and UO_771 (O_771,N_9598,N_9652);
nor UO_772 (O_772,N_8574,N_8731);
and UO_773 (O_773,N_8006,N_7899);
nand UO_774 (O_774,N_9065,N_9177);
nand UO_775 (O_775,N_8140,N_8244);
nand UO_776 (O_776,N_9445,N_9826);
and UO_777 (O_777,N_9800,N_9040);
and UO_778 (O_778,N_9732,N_8910);
nand UO_779 (O_779,N_9970,N_7540);
nand UO_780 (O_780,N_8610,N_7771);
or UO_781 (O_781,N_7584,N_8996);
xor UO_782 (O_782,N_9561,N_7858);
nor UO_783 (O_783,N_9921,N_7803);
xnor UO_784 (O_784,N_9660,N_8195);
xor UO_785 (O_785,N_9098,N_8634);
nand UO_786 (O_786,N_8868,N_9172);
xor UO_787 (O_787,N_8078,N_9350);
xor UO_788 (O_788,N_9304,N_9012);
or UO_789 (O_789,N_7909,N_9638);
nor UO_790 (O_790,N_9131,N_8220);
nor UO_791 (O_791,N_9233,N_8079);
and UO_792 (O_792,N_8070,N_9934);
nand UO_793 (O_793,N_9202,N_9136);
nand UO_794 (O_794,N_8388,N_9420);
or UO_795 (O_795,N_9241,N_8552);
nand UO_796 (O_796,N_9010,N_9759);
nand UO_797 (O_797,N_9228,N_7524);
nor UO_798 (O_798,N_8975,N_8627);
nand UO_799 (O_799,N_9582,N_9069);
nor UO_800 (O_800,N_8584,N_9647);
nand UO_801 (O_801,N_8338,N_9074);
nor UO_802 (O_802,N_9801,N_9823);
and UO_803 (O_803,N_9511,N_7594);
nor UO_804 (O_804,N_7837,N_8772);
nor UO_805 (O_805,N_9236,N_8949);
or UO_806 (O_806,N_9388,N_9022);
and UO_807 (O_807,N_9095,N_8412);
nand UO_808 (O_808,N_8698,N_9440);
nand UO_809 (O_809,N_9243,N_8618);
and UO_810 (O_810,N_7704,N_8839);
nand UO_811 (O_811,N_9639,N_8739);
nand UO_812 (O_812,N_8252,N_7850);
or UO_813 (O_813,N_8110,N_9390);
nor UO_814 (O_814,N_7856,N_8558);
nand UO_815 (O_815,N_9695,N_9124);
and UO_816 (O_816,N_7662,N_8075);
and UO_817 (O_817,N_9914,N_8464);
nand UO_818 (O_818,N_9071,N_9720);
nor UO_819 (O_819,N_9097,N_9201);
nor UO_820 (O_820,N_8355,N_9235);
nor UO_821 (O_821,N_9772,N_7777);
nand UO_822 (O_822,N_7685,N_8474);
xor UO_823 (O_823,N_9297,N_7563);
or UO_824 (O_824,N_8100,N_9296);
or UO_825 (O_825,N_9203,N_9798);
nor UO_826 (O_826,N_8063,N_8871);
xor UO_827 (O_827,N_9837,N_9494);
and UO_828 (O_828,N_8636,N_7601);
and UO_829 (O_829,N_8841,N_8520);
xor UO_830 (O_830,N_8457,N_8401);
nor UO_831 (O_831,N_9056,N_9513);
or UO_832 (O_832,N_9790,N_9122);
and UO_833 (O_833,N_8639,N_9454);
and UO_834 (O_834,N_8231,N_7853);
nand UO_835 (O_835,N_9227,N_8970);
nor UO_836 (O_836,N_7806,N_9061);
nand UO_837 (O_837,N_8448,N_8987);
or UO_838 (O_838,N_9929,N_9030);
nor UO_839 (O_839,N_9206,N_7522);
xnor UO_840 (O_840,N_7670,N_7664);
nand UO_841 (O_841,N_7981,N_7843);
and UO_842 (O_842,N_8061,N_9082);
nand UO_843 (O_843,N_9692,N_8961);
nand UO_844 (O_844,N_9886,N_9384);
nand UO_845 (O_845,N_8661,N_9402);
nor UO_846 (O_846,N_8791,N_9691);
xnor UO_847 (O_847,N_8571,N_7760);
nand UO_848 (O_848,N_8519,N_9118);
nor UO_849 (O_849,N_8013,N_9670);
nor UO_850 (O_850,N_8656,N_9885);
or UO_851 (O_851,N_8976,N_8894);
or UO_852 (O_852,N_8537,N_8059);
and UO_853 (O_853,N_8198,N_7733);
nor UO_854 (O_854,N_8296,N_9401);
and UO_855 (O_855,N_7752,N_7644);
nor UO_856 (O_856,N_8509,N_9831);
nor UO_857 (O_857,N_8580,N_8203);
or UO_858 (O_858,N_8047,N_9600);
or UO_859 (O_859,N_9697,N_7986);
nor UO_860 (O_860,N_9519,N_8123);
nor UO_861 (O_861,N_9897,N_8116);
nor UO_862 (O_862,N_8275,N_8912);
nor UO_863 (O_863,N_8804,N_8004);
and UO_864 (O_864,N_8415,N_8832);
nor UO_865 (O_865,N_9452,N_8417);
nand UO_866 (O_866,N_9546,N_8441);
and UO_867 (O_867,N_9737,N_9111);
and UO_868 (O_868,N_8681,N_9147);
nand UO_869 (O_869,N_8885,N_8085);
nor UO_870 (O_870,N_7720,N_9899);
nor UO_871 (O_871,N_9960,N_8743);
nand UO_872 (O_872,N_7818,N_8599);
xor UO_873 (O_873,N_8178,N_8540);
xor UO_874 (O_874,N_9407,N_9703);
nor UO_875 (O_875,N_8449,N_8735);
nor UO_876 (O_876,N_9337,N_9282);
nand UO_877 (O_877,N_7573,N_8664);
nor UO_878 (O_878,N_9861,N_8339);
nand UO_879 (O_879,N_8786,N_9377);
nand UO_880 (O_880,N_7678,N_8607);
xnor UO_881 (O_881,N_8168,N_9316);
and UO_882 (O_882,N_8919,N_9469);
nor UO_883 (O_883,N_9100,N_7973);
nand UO_884 (O_884,N_7860,N_9306);
nor UO_885 (O_885,N_8212,N_8422);
and UO_886 (O_886,N_9874,N_9037);
and UO_887 (O_887,N_8765,N_8157);
nor UO_888 (O_888,N_9883,N_8387);
xnor UO_889 (O_889,N_7646,N_8335);
and UO_890 (O_890,N_9311,N_8094);
nand UO_891 (O_891,N_8747,N_9529);
nor UO_892 (O_892,N_7566,N_8496);
nor UO_893 (O_893,N_9827,N_7552);
nor UO_894 (O_894,N_8137,N_9992);
nor UO_895 (O_895,N_9151,N_9217);
xor UO_896 (O_896,N_8646,N_7847);
or UO_897 (O_897,N_8450,N_9387);
xnor UO_898 (O_898,N_7729,N_8316);
xor UO_899 (O_899,N_9165,N_8758);
and UO_900 (O_900,N_8480,N_9338);
and UO_901 (O_901,N_8909,N_8443);
or UO_902 (O_902,N_9974,N_9134);
nor UO_903 (O_903,N_7675,N_8218);
and UO_904 (O_904,N_9349,N_8924);
nand UO_905 (O_905,N_8900,N_8163);
nor UO_906 (O_906,N_7727,N_8865);
and UO_907 (O_907,N_9865,N_8421);
nand UO_908 (O_908,N_7721,N_9533);
nor UO_909 (O_909,N_9730,N_9050);
and UO_910 (O_910,N_9476,N_8820);
nor UO_911 (O_911,N_9845,N_8718);
xnor UO_912 (O_912,N_9164,N_7730);
xnor UO_913 (O_913,N_8208,N_9940);
or UO_914 (O_914,N_7545,N_9137);
or UO_915 (O_915,N_8686,N_8213);
xnor UO_916 (O_916,N_7641,N_9000);
and UO_917 (O_917,N_9254,N_9216);
nand UO_918 (O_918,N_9332,N_9810);
nand UO_919 (O_919,N_7725,N_7998);
or UO_920 (O_920,N_9860,N_7597);
nand UO_921 (O_921,N_8802,N_9364);
nand UO_922 (O_922,N_8506,N_9257);
nand UO_923 (O_923,N_9339,N_8539);
and UO_924 (O_924,N_9510,N_8845);
nor UO_925 (O_925,N_8395,N_9981);
and UO_926 (O_926,N_8768,N_8572);
or UO_927 (O_927,N_9770,N_9032);
nand UO_928 (O_928,N_8024,N_9138);
nand UO_929 (O_929,N_8525,N_9962);
and UO_930 (O_930,N_7571,N_7753);
and UO_931 (O_931,N_9267,N_9943);
nand UO_932 (O_932,N_8065,N_9799);
or UO_933 (O_933,N_8125,N_8526);
nand UO_934 (O_934,N_8020,N_9677);
or UO_935 (O_935,N_7618,N_8914);
nand UO_936 (O_936,N_8416,N_8367);
and UO_937 (O_937,N_7844,N_8853);
nor UO_938 (O_938,N_8284,N_8354);
and UO_939 (O_939,N_8408,N_7831);
and UO_940 (O_940,N_8974,N_7937);
xnor UO_941 (O_941,N_8787,N_8184);
nand UO_942 (O_942,N_9822,N_7848);
and UO_943 (O_943,N_8964,N_8978);
nor UO_944 (O_944,N_8510,N_8826);
and UO_945 (O_945,N_8827,N_9193);
and UO_946 (O_946,N_8788,N_9159);
nand UO_947 (O_947,N_8825,N_9451);
nand UO_948 (O_948,N_8486,N_9531);
nor UO_949 (O_949,N_8166,N_9343);
nand UO_950 (O_950,N_8596,N_8102);
and UO_951 (O_951,N_8507,N_8882);
xor UO_952 (O_952,N_7578,N_8837);
or UO_953 (O_953,N_8276,N_8333);
nor UO_954 (O_954,N_9975,N_7606);
nor UO_955 (O_955,N_8010,N_9125);
nor UO_956 (O_956,N_9780,N_8807);
and UO_957 (O_957,N_8939,N_9456);
xor UO_958 (O_958,N_9836,N_9787);
nor UO_959 (O_959,N_9721,N_9093);
xnor UO_960 (O_960,N_9190,N_9917);
or UO_961 (O_961,N_9602,N_8586);
or UO_962 (O_962,N_8702,N_7560);
xor UO_963 (O_963,N_7693,N_8440);
xnor UO_964 (O_964,N_9663,N_9214);
nand UO_965 (O_965,N_9029,N_8331);
or UO_966 (O_966,N_8159,N_8082);
and UO_967 (O_967,N_8253,N_9986);
and UO_968 (O_968,N_7750,N_9409);
nor UO_969 (O_969,N_8800,N_8400);
or UO_970 (O_970,N_8491,N_9035);
nand UO_971 (O_971,N_8317,N_8381);
or UO_972 (O_972,N_9933,N_7821);
nand UO_973 (O_973,N_9152,N_9522);
xnor UO_974 (O_974,N_9918,N_7807);
and UO_975 (O_975,N_7893,N_7894);
nand UO_976 (O_976,N_7751,N_8424);
and UO_977 (O_977,N_8544,N_7908);
nand UO_978 (O_978,N_8500,N_7995);
nand UO_979 (O_979,N_8470,N_9870);
and UO_980 (O_980,N_9191,N_9543);
or UO_981 (O_981,N_7940,N_8953);
nor UO_982 (O_982,N_8000,N_8112);
xor UO_983 (O_983,N_9853,N_7546);
nor UO_984 (O_984,N_7835,N_9154);
or UO_985 (O_985,N_9811,N_7586);
or UO_986 (O_986,N_9792,N_8056);
nor UO_987 (O_987,N_7619,N_9674);
or UO_988 (O_988,N_9455,N_8309);
nor UO_989 (O_989,N_8369,N_9229);
or UO_990 (O_990,N_9506,N_8606);
and UO_991 (O_991,N_9205,N_8784);
and UO_992 (O_992,N_8461,N_7954);
and UO_993 (O_993,N_9373,N_8904);
or UO_994 (O_994,N_9078,N_9807);
and UO_995 (O_995,N_7615,N_9623);
and UO_996 (O_996,N_8451,N_8413);
nor UO_997 (O_997,N_9725,N_8266);
or UO_998 (O_998,N_8657,N_9273);
nor UO_999 (O_999,N_7501,N_9951);
or UO_1000 (O_1000,N_9424,N_9368);
nand UO_1001 (O_1001,N_9540,N_9873);
nand UO_1002 (O_1002,N_9586,N_9027);
xor UO_1003 (O_1003,N_7959,N_8265);
or UO_1004 (O_1004,N_8382,N_7632);
and UO_1005 (O_1005,N_9443,N_9490);
nor UO_1006 (O_1006,N_8096,N_9610);
or UO_1007 (O_1007,N_8989,N_9908);
or UO_1008 (O_1008,N_7877,N_9550);
and UO_1009 (O_1009,N_8127,N_7738);
or UO_1010 (O_1010,N_9302,N_8842);
and UO_1011 (O_1011,N_9184,N_8761);
nand UO_1012 (O_1012,N_8847,N_8993);
or UO_1013 (O_1013,N_9507,N_7903);
or UO_1014 (O_1014,N_8585,N_9336);
and UO_1015 (O_1015,N_8550,N_7827);
nor UO_1016 (O_1016,N_7985,N_7614);
nand UO_1017 (O_1017,N_8959,N_8672);
or UO_1018 (O_1018,N_7603,N_7808);
nand UO_1019 (O_1019,N_9619,N_8734);
nand UO_1020 (O_1020,N_8776,N_8161);
or UO_1021 (O_1021,N_9740,N_9431);
nor UO_1022 (O_1022,N_8038,N_9672);
nor UO_1023 (O_1023,N_8538,N_8466);
and UO_1024 (O_1024,N_7677,N_9072);
or UO_1025 (O_1025,N_9054,N_9839);
and UO_1026 (O_1026,N_9509,N_8601);
and UO_1027 (O_1027,N_9230,N_9025);
and UO_1028 (O_1028,N_9499,N_9326);
nand UO_1029 (O_1029,N_9067,N_9824);
xnor UO_1030 (O_1030,N_9794,N_8932);
xnor UO_1031 (O_1031,N_7585,N_9375);
xor UO_1032 (O_1032,N_8023,N_9127);
and UO_1033 (O_1033,N_9086,N_7547);
xor UO_1034 (O_1034,N_9261,N_8926);
nand UO_1035 (O_1035,N_9812,N_9314);
and UO_1036 (O_1036,N_9840,N_9572);
xor UO_1037 (O_1037,N_9937,N_7975);
and UO_1038 (O_1038,N_9017,N_9700);
and UO_1039 (O_1039,N_9585,N_9459);
nor UO_1040 (O_1040,N_9843,N_8822);
nand UO_1041 (O_1041,N_8921,N_8881);
xor UO_1042 (O_1042,N_8738,N_8209);
nand UO_1043 (O_1043,N_8149,N_9109);
or UO_1044 (O_1044,N_8815,N_8439);
nand UO_1045 (O_1045,N_7551,N_8813);
nand UO_1046 (O_1046,N_8649,N_9318);
nor UO_1047 (O_1047,N_8427,N_8442);
nor UO_1048 (O_1048,N_7916,N_8930);
or UO_1049 (O_1049,N_9525,N_8777);
nand UO_1050 (O_1050,N_8215,N_7737);
nor UO_1051 (O_1051,N_9571,N_7884);
nor UO_1052 (O_1052,N_9654,N_9709);
and UO_1053 (O_1053,N_9278,N_8147);
nor UO_1054 (O_1054,N_8977,N_7914);
nor UO_1055 (O_1055,N_8205,N_9678);
or UO_1056 (O_1056,N_9465,N_8481);
or UO_1057 (O_1057,N_8947,N_8759);
nor UO_1058 (O_1058,N_7804,N_7989);
nand UO_1059 (O_1059,N_8173,N_9168);
or UO_1060 (O_1060,N_8492,N_8142);
and UO_1061 (O_1061,N_9161,N_8171);
and UO_1062 (O_1062,N_9922,N_9641);
nor UO_1063 (O_1063,N_8145,N_8631);
nand UO_1064 (O_1064,N_9645,N_8021);
and UO_1065 (O_1065,N_8652,N_8353);
nor UO_1066 (O_1066,N_7735,N_7722);
or UO_1067 (O_1067,N_8043,N_8384);
nand UO_1068 (O_1068,N_8054,N_7930);
nand UO_1069 (O_1069,N_8298,N_8821);
or UO_1070 (O_1070,N_8327,N_9247);
xor UO_1071 (O_1071,N_8779,N_7673);
nor UO_1072 (O_1072,N_9433,N_9143);
nand UO_1073 (O_1073,N_8177,N_9548);
nor UO_1074 (O_1074,N_9979,N_7577);
nor UO_1075 (O_1075,N_9156,N_9466);
nand UO_1076 (O_1076,N_8941,N_8630);
xor UO_1077 (O_1077,N_9989,N_7740);
nor UO_1078 (O_1078,N_8819,N_7961);
or UO_1079 (O_1079,N_8893,N_9395);
and UO_1080 (O_1080,N_9026,N_9011);
or UO_1081 (O_1081,N_9524,N_7622);
and UO_1082 (O_1082,N_7825,N_9667);
and UO_1083 (O_1083,N_8030,N_7640);
and UO_1084 (O_1084,N_9442,N_9263);
or UO_1085 (O_1085,N_9008,N_8617);
or UO_1086 (O_1086,N_7864,N_8992);
and UO_1087 (O_1087,N_8816,N_8803);
nor UO_1088 (O_1088,N_7515,N_9258);
nand UO_1089 (O_1089,N_8311,N_9369);
nand UO_1090 (O_1090,N_8240,N_9279);
and UO_1091 (O_1091,N_9485,N_8551);
nand UO_1092 (O_1092,N_8703,N_8489);
nand UO_1093 (O_1093,N_8654,N_9796);
or UO_1094 (O_1094,N_9315,N_8712);
and UO_1095 (O_1095,N_9634,N_9560);
nand UO_1096 (O_1096,N_9240,N_8888);
nor UO_1097 (O_1097,N_8838,N_7648);
or UO_1098 (O_1098,N_7579,N_9481);
or UO_1099 (O_1099,N_8305,N_8667);
nand UO_1100 (O_1100,N_9747,N_9954);
nor UO_1101 (O_1101,N_8600,N_7543);
or UO_1102 (O_1102,N_8951,N_8036);
or UO_1103 (O_1103,N_8086,N_9252);
and UO_1104 (O_1104,N_7599,N_9746);
and UO_1105 (O_1105,N_9389,N_8106);
nor UO_1106 (O_1106,N_9031,N_8793);
nand UO_1107 (O_1107,N_8285,N_8562);
nand UO_1108 (O_1108,N_9063,N_9972);
nand UO_1109 (O_1109,N_9308,N_7983);
or UO_1110 (O_1110,N_9380,N_9286);
and UO_1111 (O_1111,N_7748,N_8462);
nand UO_1112 (O_1112,N_7598,N_9900);
or UO_1113 (O_1113,N_8990,N_9640);
or UO_1114 (O_1114,N_9412,N_8058);
nand UO_1115 (O_1115,N_8624,N_8751);
nor UO_1116 (O_1116,N_8019,N_8564);
or UO_1117 (O_1117,N_8473,N_8426);
or UO_1118 (O_1118,N_8796,N_7611);
and UO_1119 (O_1119,N_7593,N_8386);
and UO_1120 (O_1120,N_9197,N_8901);
or UO_1121 (O_1121,N_9317,N_7759);
and UO_1122 (O_1122,N_9592,N_9117);
nor UO_1123 (O_1123,N_7694,N_8797);
and UO_1124 (O_1124,N_7783,N_8588);
and UO_1125 (O_1125,N_9761,N_8264);
nor UO_1126 (O_1126,N_9675,N_9145);
nand UO_1127 (O_1127,N_9614,N_9742);
and UO_1128 (O_1128,N_7582,N_7911);
or UO_1129 (O_1129,N_8182,N_9712);
nand UO_1130 (O_1130,N_7788,N_8749);
and UO_1131 (O_1131,N_7651,N_9448);
or UO_1132 (O_1132,N_7692,N_7859);
xor UO_1133 (O_1133,N_9475,N_9482);
and UO_1134 (O_1134,N_7800,N_7889);
nor UO_1135 (O_1135,N_9376,N_7576);
or UO_1136 (O_1136,N_9949,N_9726);
nor UO_1137 (O_1137,N_8162,N_8458);
and UO_1138 (O_1138,N_9383,N_7506);
and UO_1139 (O_1139,N_7876,N_9755);
and UO_1140 (O_1140,N_8039,N_9734);
and UO_1141 (O_1141,N_8018,N_9988);
nand UO_1142 (O_1142,N_8390,N_7549);
nand UO_1143 (O_1143,N_9863,N_9788);
nand UO_1144 (O_1144,N_9288,N_8224);
and UO_1145 (O_1145,N_8278,N_8648);
nand UO_1146 (O_1146,N_8206,N_9871);
nor UO_1147 (O_1147,N_9255,N_8896);
or UO_1148 (O_1148,N_9028,N_9872);
and UO_1149 (O_1149,N_9280,N_9617);
and UO_1150 (O_1150,N_7682,N_9463);
nor UO_1151 (O_1151,N_8907,N_8828);
or UO_1152 (O_1152,N_9688,N_9323);
nand UO_1153 (O_1153,N_7653,N_9892);
nor UO_1154 (O_1154,N_9930,N_7901);
nor UO_1155 (O_1155,N_9583,N_7923);
or UO_1156 (O_1156,N_8155,N_7811);
or UO_1157 (O_1157,N_9624,N_9200);
nand UO_1158 (O_1158,N_8499,N_8495);
or UO_1159 (O_1159,N_8258,N_9875);
nand UO_1160 (O_1160,N_9898,N_9939);
or UO_1161 (O_1161,N_9113,N_9906);
or UO_1162 (O_1162,N_8531,N_9291);
and UO_1163 (O_1163,N_8983,N_9681);
xor UO_1164 (O_1164,N_9392,N_9779);
nand UO_1165 (O_1165,N_7797,N_9187);
or UO_1166 (O_1166,N_7714,N_9536);
nor UO_1167 (O_1167,N_7938,N_8516);
and UO_1168 (O_1168,N_9731,N_9508);
xor UO_1169 (O_1169,N_7924,N_9607);
nand UO_1170 (O_1170,N_7991,N_9425);
or UO_1171 (O_1171,N_8812,N_9880);
nor UO_1172 (O_1172,N_9544,N_9894);
nand UO_1173 (O_1173,N_7933,N_9982);
or UO_1174 (O_1174,N_8016,N_9049);
or UO_1175 (O_1175,N_8478,N_9595);
nor UO_1176 (O_1176,N_8673,N_9268);
nor UO_1177 (O_1177,N_8411,N_8778);
nand UO_1178 (O_1178,N_8297,N_9298);
xor UO_1179 (O_1179,N_8444,N_8098);
or UO_1180 (O_1180,N_9987,N_9186);
nand UO_1181 (O_1181,N_9271,N_7570);
nor UO_1182 (O_1182,N_7746,N_9489);
or UO_1183 (O_1183,N_7732,N_8521);
or UO_1184 (O_1184,N_9862,N_8189);
and UO_1185 (O_1185,N_9365,N_9274);
xor UO_1186 (O_1186,N_8780,N_8124);
nand UO_1187 (O_1187,N_8508,N_7810);
or UO_1188 (O_1188,N_7568,N_8329);
nand UO_1189 (O_1189,N_8051,N_8680);
nor UO_1190 (O_1190,N_8488,N_8493);
nor UO_1191 (O_1191,N_7769,N_9941);
xor UO_1192 (O_1192,N_7630,N_9956);
nor UO_1193 (O_1193,N_8722,N_7927);
or UO_1194 (O_1194,N_9948,N_8107);
nor UO_1195 (O_1195,N_8225,N_8814);
and UO_1196 (O_1196,N_8467,N_9597);
and UO_1197 (O_1197,N_8113,N_9042);
xor UO_1198 (O_1198,N_8062,N_9094);
nand UO_1199 (O_1199,N_7796,N_8724);
and UO_1200 (O_1200,N_7898,N_8370);
nor UO_1201 (O_1201,N_8446,N_9195);
xnor UO_1202 (O_1202,N_8232,N_7996);
and UO_1203 (O_1203,N_8077,N_7979);
or UO_1204 (O_1204,N_9739,N_7960);
or UO_1205 (O_1205,N_8289,N_9325);
nand UO_1206 (O_1206,N_8940,N_9821);
nand UO_1207 (O_1207,N_8609,N_8663);
nor UO_1208 (O_1208,N_9179,N_9284);
nor UO_1209 (O_1209,N_8916,N_9716);
or UO_1210 (O_1210,N_8188,N_7958);
nor UO_1211 (O_1211,N_9321,N_8771);
or UO_1212 (O_1212,N_7712,N_8640);
xor UO_1213 (O_1213,N_8934,N_8922);
nor UO_1214 (O_1214,N_9178,N_8346);
nand UO_1215 (O_1215,N_8216,N_9539);
nand UO_1216 (O_1216,N_8578,N_9666);
nand UO_1217 (O_1217,N_8138,N_7713);
nor UO_1218 (O_1218,N_9285,N_9500);
nor UO_1219 (O_1219,N_9776,N_9269);
or UO_1220 (O_1220,N_9961,N_9622);
nor UO_1221 (O_1221,N_8829,N_8254);
and UO_1222 (O_1222,N_8706,N_8037);
or UO_1223 (O_1223,N_8873,N_9715);
and UO_1224 (O_1224,N_8741,N_7529);
nand UO_1225 (O_1225,N_9512,N_9785);
and UO_1226 (O_1226,N_9613,N_8867);
nand UO_1227 (O_1227,N_8555,N_8366);
and UO_1228 (O_1228,N_8394,N_8679);
and UO_1229 (O_1229,N_7965,N_7513);
nand UO_1230 (O_1230,N_9809,N_8968);
and UO_1231 (O_1231,N_8898,N_7774);
nand UO_1232 (O_1232,N_7822,N_9938);
nand UO_1233 (O_1233,N_8172,N_8418);
nand UO_1234 (O_1234,N_9327,N_9803);
nor UO_1235 (O_1235,N_8557,N_9935);
nand UO_1236 (O_1236,N_8176,N_7988);
or UO_1237 (O_1237,N_8068,N_9410);
and UO_1238 (O_1238,N_9802,N_8659);
xor UO_1239 (O_1239,N_9545,N_9467);
nor UO_1240 (O_1240,N_8560,N_8612);
nand UO_1241 (O_1241,N_9556,N_9039);
nand UO_1242 (O_1242,N_9947,N_8946);
or UO_1243 (O_1243,N_9253,N_8878);
nor UO_1244 (O_1244,N_7534,N_7897);
or UO_1245 (O_1245,N_9997,N_7895);
nor UO_1246 (O_1246,N_8245,N_8011);
xor UO_1247 (O_1247,N_9488,N_7509);
xor UO_1248 (O_1248,N_9036,N_9062);
xor UO_1249 (O_1249,N_8598,N_8239);
or UO_1250 (O_1250,N_7912,N_7536);
or UO_1251 (O_1251,N_8682,N_9515);
or UO_1252 (O_1252,N_9805,N_7687);
and UO_1253 (O_1253,N_8587,N_8347);
nor UO_1254 (O_1254,N_9235,N_9752);
or UO_1255 (O_1255,N_9888,N_7684);
nor UO_1256 (O_1256,N_8072,N_8407);
xor UO_1257 (O_1257,N_9521,N_9672);
nor UO_1258 (O_1258,N_7697,N_8251);
nand UO_1259 (O_1259,N_9936,N_8515);
nor UO_1260 (O_1260,N_9148,N_8937);
or UO_1261 (O_1261,N_7513,N_9529);
nand UO_1262 (O_1262,N_7581,N_9578);
and UO_1263 (O_1263,N_7565,N_8372);
nand UO_1264 (O_1264,N_7899,N_8236);
nor UO_1265 (O_1265,N_9155,N_8014);
nand UO_1266 (O_1266,N_9969,N_8752);
or UO_1267 (O_1267,N_8078,N_7999);
xor UO_1268 (O_1268,N_8369,N_7589);
nor UO_1269 (O_1269,N_9247,N_8445);
nor UO_1270 (O_1270,N_9152,N_9642);
xnor UO_1271 (O_1271,N_9344,N_8982);
and UO_1272 (O_1272,N_9600,N_9221);
or UO_1273 (O_1273,N_9081,N_9875);
nor UO_1274 (O_1274,N_9633,N_8756);
and UO_1275 (O_1275,N_8859,N_8081);
and UO_1276 (O_1276,N_7658,N_9732);
nor UO_1277 (O_1277,N_9255,N_9524);
nor UO_1278 (O_1278,N_9766,N_8909);
nand UO_1279 (O_1279,N_8077,N_8571);
and UO_1280 (O_1280,N_7593,N_7805);
nand UO_1281 (O_1281,N_7988,N_9652);
and UO_1282 (O_1282,N_9764,N_9156);
nor UO_1283 (O_1283,N_8574,N_8052);
nor UO_1284 (O_1284,N_9958,N_9872);
or UO_1285 (O_1285,N_7803,N_9647);
xor UO_1286 (O_1286,N_8311,N_8675);
or UO_1287 (O_1287,N_9782,N_9020);
nor UO_1288 (O_1288,N_7513,N_8899);
nor UO_1289 (O_1289,N_7550,N_9432);
nand UO_1290 (O_1290,N_9517,N_9207);
nor UO_1291 (O_1291,N_9885,N_8311);
nand UO_1292 (O_1292,N_9488,N_8635);
and UO_1293 (O_1293,N_8447,N_7912);
and UO_1294 (O_1294,N_8692,N_9564);
nor UO_1295 (O_1295,N_7862,N_7742);
nand UO_1296 (O_1296,N_9305,N_9525);
and UO_1297 (O_1297,N_8349,N_9104);
nand UO_1298 (O_1298,N_9070,N_9616);
nand UO_1299 (O_1299,N_7917,N_7644);
nor UO_1300 (O_1300,N_8638,N_9512);
or UO_1301 (O_1301,N_9787,N_7999);
nand UO_1302 (O_1302,N_7950,N_7990);
and UO_1303 (O_1303,N_7833,N_9251);
or UO_1304 (O_1304,N_9304,N_7864);
nor UO_1305 (O_1305,N_8334,N_9383);
and UO_1306 (O_1306,N_8447,N_7741);
or UO_1307 (O_1307,N_9635,N_9744);
nand UO_1308 (O_1308,N_9324,N_9638);
and UO_1309 (O_1309,N_9281,N_9309);
and UO_1310 (O_1310,N_8507,N_9611);
nor UO_1311 (O_1311,N_7511,N_8655);
nand UO_1312 (O_1312,N_8378,N_9577);
or UO_1313 (O_1313,N_8485,N_9609);
and UO_1314 (O_1314,N_9808,N_8896);
nand UO_1315 (O_1315,N_8674,N_9840);
or UO_1316 (O_1316,N_9743,N_7913);
and UO_1317 (O_1317,N_9675,N_8941);
xnor UO_1318 (O_1318,N_8704,N_7642);
or UO_1319 (O_1319,N_9158,N_9319);
or UO_1320 (O_1320,N_9184,N_7991);
nand UO_1321 (O_1321,N_9965,N_8033);
nand UO_1322 (O_1322,N_9078,N_7507);
xnor UO_1323 (O_1323,N_7550,N_9781);
nor UO_1324 (O_1324,N_9820,N_8296);
or UO_1325 (O_1325,N_8032,N_8582);
or UO_1326 (O_1326,N_8385,N_8270);
or UO_1327 (O_1327,N_8609,N_8785);
nor UO_1328 (O_1328,N_9969,N_8790);
or UO_1329 (O_1329,N_7635,N_8235);
nand UO_1330 (O_1330,N_7793,N_9936);
nor UO_1331 (O_1331,N_8684,N_8237);
and UO_1332 (O_1332,N_9546,N_9630);
nand UO_1333 (O_1333,N_9255,N_9519);
and UO_1334 (O_1334,N_7760,N_8198);
nand UO_1335 (O_1335,N_7633,N_9525);
and UO_1336 (O_1336,N_8352,N_7630);
or UO_1337 (O_1337,N_8505,N_9159);
nand UO_1338 (O_1338,N_9051,N_9890);
nor UO_1339 (O_1339,N_9986,N_9338);
nor UO_1340 (O_1340,N_7877,N_7839);
nand UO_1341 (O_1341,N_8106,N_9089);
and UO_1342 (O_1342,N_9854,N_9175);
nor UO_1343 (O_1343,N_9761,N_9080);
nor UO_1344 (O_1344,N_8878,N_9575);
nand UO_1345 (O_1345,N_9240,N_7714);
or UO_1346 (O_1346,N_9495,N_8864);
and UO_1347 (O_1347,N_8452,N_7912);
and UO_1348 (O_1348,N_8205,N_8284);
nor UO_1349 (O_1349,N_9559,N_8970);
and UO_1350 (O_1350,N_8356,N_9073);
and UO_1351 (O_1351,N_8059,N_8419);
and UO_1352 (O_1352,N_7886,N_8685);
and UO_1353 (O_1353,N_8019,N_9743);
nor UO_1354 (O_1354,N_9831,N_8476);
nor UO_1355 (O_1355,N_9144,N_7716);
nor UO_1356 (O_1356,N_9410,N_9828);
or UO_1357 (O_1357,N_7808,N_8737);
nand UO_1358 (O_1358,N_9996,N_9227);
nand UO_1359 (O_1359,N_7849,N_8963);
and UO_1360 (O_1360,N_8744,N_9904);
and UO_1361 (O_1361,N_8772,N_8097);
nand UO_1362 (O_1362,N_8128,N_8854);
nor UO_1363 (O_1363,N_9392,N_8424);
nor UO_1364 (O_1364,N_9827,N_7576);
nor UO_1365 (O_1365,N_8035,N_7763);
nand UO_1366 (O_1366,N_9684,N_9566);
and UO_1367 (O_1367,N_9078,N_8312);
nor UO_1368 (O_1368,N_8582,N_9218);
and UO_1369 (O_1369,N_7831,N_8032);
and UO_1370 (O_1370,N_7547,N_8795);
nor UO_1371 (O_1371,N_8256,N_9857);
and UO_1372 (O_1372,N_8400,N_8522);
nor UO_1373 (O_1373,N_8630,N_7559);
nor UO_1374 (O_1374,N_9813,N_7679);
and UO_1375 (O_1375,N_9020,N_7745);
or UO_1376 (O_1376,N_8328,N_9287);
nand UO_1377 (O_1377,N_8538,N_7533);
or UO_1378 (O_1378,N_8562,N_8935);
or UO_1379 (O_1379,N_9011,N_8384);
nor UO_1380 (O_1380,N_9618,N_9924);
nand UO_1381 (O_1381,N_9476,N_7920);
xnor UO_1382 (O_1382,N_9046,N_9815);
nor UO_1383 (O_1383,N_8540,N_8139);
or UO_1384 (O_1384,N_7902,N_8407);
nor UO_1385 (O_1385,N_7789,N_8801);
or UO_1386 (O_1386,N_9992,N_8923);
xnor UO_1387 (O_1387,N_8336,N_8671);
nand UO_1388 (O_1388,N_8844,N_7584);
xnor UO_1389 (O_1389,N_9785,N_8285);
and UO_1390 (O_1390,N_9924,N_7726);
xnor UO_1391 (O_1391,N_8582,N_9312);
nand UO_1392 (O_1392,N_7574,N_8172);
nor UO_1393 (O_1393,N_8367,N_7745);
xor UO_1394 (O_1394,N_8224,N_8452);
nand UO_1395 (O_1395,N_7607,N_9075);
or UO_1396 (O_1396,N_8402,N_8193);
and UO_1397 (O_1397,N_7994,N_8536);
nor UO_1398 (O_1398,N_7590,N_9350);
xnor UO_1399 (O_1399,N_8714,N_8351);
or UO_1400 (O_1400,N_9008,N_9765);
and UO_1401 (O_1401,N_9452,N_8035);
nand UO_1402 (O_1402,N_7590,N_7874);
nor UO_1403 (O_1403,N_9948,N_9478);
xor UO_1404 (O_1404,N_7596,N_7844);
nor UO_1405 (O_1405,N_9430,N_9068);
nand UO_1406 (O_1406,N_8814,N_8705);
nor UO_1407 (O_1407,N_8464,N_8737);
nand UO_1408 (O_1408,N_8738,N_8436);
nand UO_1409 (O_1409,N_8879,N_8028);
xor UO_1410 (O_1410,N_7946,N_8138);
nand UO_1411 (O_1411,N_9000,N_7780);
and UO_1412 (O_1412,N_7634,N_9621);
and UO_1413 (O_1413,N_7780,N_9882);
and UO_1414 (O_1414,N_9035,N_8218);
and UO_1415 (O_1415,N_9091,N_9871);
nand UO_1416 (O_1416,N_9094,N_7914);
xor UO_1417 (O_1417,N_9694,N_9518);
or UO_1418 (O_1418,N_8334,N_8887);
and UO_1419 (O_1419,N_8153,N_7720);
nor UO_1420 (O_1420,N_7682,N_8367);
and UO_1421 (O_1421,N_8198,N_8821);
and UO_1422 (O_1422,N_7770,N_9385);
and UO_1423 (O_1423,N_7769,N_9872);
xnor UO_1424 (O_1424,N_9054,N_9150);
nand UO_1425 (O_1425,N_8787,N_9794);
nand UO_1426 (O_1426,N_9028,N_8985);
xor UO_1427 (O_1427,N_8773,N_9932);
or UO_1428 (O_1428,N_7914,N_9165);
nor UO_1429 (O_1429,N_9930,N_9331);
or UO_1430 (O_1430,N_7988,N_9170);
nor UO_1431 (O_1431,N_8090,N_7898);
xor UO_1432 (O_1432,N_7716,N_8556);
and UO_1433 (O_1433,N_9892,N_8479);
nand UO_1434 (O_1434,N_8067,N_8101);
or UO_1435 (O_1435,N_9238,N_8136);
or UO_1436 (O_1436,N_9163,N_9213);
and UO_1437 (O_1437,N_8970,N_7578);
nand UO_1438 (O_1438,N_9821,N_8750);
nand UO_1439 (O_1439,N_8333,N_8785);
nor UO_1440 (O_1440,N_8641,N_8927);
nand UO_1441 (O_1441,N_8493,N_8093);
nor UO_1442 (O_1442,N_8256,N_8692);
or UO_1443 (O_1443,N_9552,N_9990);
and UO_1444 (O_1444,N_9803,N_8234);
nand UO_1445 (O_1445,N_9680,N_8538);
nor UO_1446 (O_1446,N_9113,N_9977);
nor UO_1447 (O_1447,N_7987,N_7736);
or UO_1448 (O_1448,N_9385,N_7717);
nor UO_1449 (O_1449,N_8665,N_8151);
and UO_1450 (O_1450,N_7581,N_8573);
nor UO_1451 (O_1451,N_9459,N_9154);
nand UO_1452 (O_1452,N_7860,N_8260);
nor UO_1453 (O_1453,N_7808,N_7944);
or UO_1454 (O_1454,N_8153,N_8947);
nand UO_1455 (O_1455,N_8325,N_8668);
nand UO_1456 (O_1456,N_8270,N_9606);
or UO_1457 (O_1457,N_9528,N_9952);
nand UO_1458 (O_1458,N_7615,N_9556);
and UO_1459 (O_1459,N_9924,N_8390);
and UO_1460 (O_1460,N_9970,N_9743);
nand UO_1461 (O_1461,N_9669,N_9284);
and UO_1462 (O_1462,N_8466,N_7866);
and UO_1463 (O_1463,N_9698,N_9146);
nor UO_1464 (O_1464,N_8837,N_9849);
nor UO_1465 (O_1465,N_7689,N_9162);
nand UO_1466 (O_1466,N_7679,N_8127);
or UO_1467 (O_1467,N_9661,N_8714);
nand UO_1468 (O_1468,N_8052,N_7641);
xnor UO_1469 (O_1469,N_8847,N_8844);
or UO_1470 (O_1470,N_9818,N_7878);
and UO_1471 (O_1471,N_8458,N_8624);
nand UO_1472 (O_1472,N_8824,N_9388);
xnor UO_1473 (O_1473,N_9084,N_9499);
or UO_1474 (O_1474,N_7987,N_9421);
or UO_1475 (O_1475,N_8627,N_9524);
nand UO_1476 (O_1476,N_7911,N_9499);
nand UO_1477 (O_1477,N_9871,N_8923);
nand UO_1478 (O_1478,N_7847,N_8560);
nor UO_1479 (O_1479,N_9451,N_7744);
nor UO_1480 (O_1480,N_9576,N_8942);
nand UO_1481 (O_1481,N_7859,N_7812);
and UO_1482 (O_1482,N_9975,N_9709);
nand UO_1483 (O_1483,N_7697,N_8392);
and UO_1484 (O_1484,N_9109,N_9061);
xnor UO_1485 (O_1485,N_7829,N_8620);
nor UO_1486 (O_1486,N_9482,N_9127);
and UO_1487 (O_1487,N_9901,N_7673);
and UO_1488 (O_1488,N_8866,N_9522);
or UO_1489 (O_1489,N_8795,N_9398);
and UO_1490 (O_1490,N_8545,N_8519);
nand UO_1491 (O_1491,N_8441,N_7874);
or UO_1492 (O_1492,N_9015,N_9713);
or UO_1493 (O_1493,N_7685,N_9365);
and UO_1494 (O_1494,N_8086,N_9102);
nand UO_1495 (O_1495,N_8451,N_8099);
nand UO_1496 (O_1496,N_9102,N_8340);
nand UO_1497 (O_1497,N_9278,N_9891);
nand UO_1498 (O_1498,N_8678,N_9053);
and UO_1499 (O_1499,N_7653,N_8099);
endmodule