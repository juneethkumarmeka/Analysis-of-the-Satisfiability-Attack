module basic_2500_25000_3000_25_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
xor U0 (N_0,In_435,In_468);
and U1 (N_1,In_2460,In_2009);
and U2 (N_2,In_226,In_2369);
nor U3 (N_3,In_277,In_672);
and U4 (N_4,In_1716,In_1575);
or U5 (N_5,In_1913,In_2044);
and U6 (N_6,In_1070,In_2057);
and U7 (N_7,In_1188,In_1622);
xnor U8 (N_8,In_397,In_382);
nor U9 (N_9,In_232,In_1559);
nor U10 (N_10,In_420,In_1309);
xor U11 (N_11,In_1998,In_1325);
and U12 (N_12,In_1220,In_602);
nand U13 (N_13,In_791,In_2290);
nand U14 (N_14,In_850,In_1897);
nor U15 (N_15,In_266,In_831);
xnor U16 (N_16,In_809,In_2233);
or U17 (N_17,In_33,In_1671);
nor U18 (N_18,In_565,In_386);
nand U19 (N_19,In_1595,In_476);
nor U20 (N_20,In_985,In_1533);
nor U21 (N_21,In_1936,In_1753);
or U22 (N_22,In_1850,In_768);
and U23 (N_23,In_2109,In_1721);
nor U24 (N_24,In_2175,In_1683);
nand U25 (N_25,In_2160,In_921);
nand U26 (N_26,In_1316,In_16);
nand U27 (N_27,In_1051,In_2248);
nor U28 (N_28,In_2181,In_26);
or U29 (N_29,In_2449,In_629);
nand U30 (N_30,In_2465,In_1699);
nand U31 (N_31,In_754,In_1706);
or U32 (N_32,In_2336,In_883);
nor U33 (N_33,In_825,In_1226);
xnor U34 (N_34,In_1734,In_2285);
and U35 (N_35,In_2488,In_2348);
and U36 (N_36,In_1892,In_1270);
nand U37 (N_37,In_1926,In_1437);
and U38 (N_38,In_1567,In_379);
nor U39 (N_39,In_2183,In_628);
and U40 (N_40,In_2299,In_220);
nor U41 (N_41,In_1079,In_490);
or U42 (N_42,In_783,In_696);
or U43 (N_43,In_906,In_669);
nand U44 (N_44,In_1896,In_2218);
xnor U45 (N_45,In_836,In_1239);
xnor U46 (N_46,In_464,In_1159);
and U47 (N_47,In_199,In_1771);
or U48 (N_48,In_418,In_2026);
and U49 (N_49,In_1137,In_2088);
or U50 (N_50,In_853,In_733);
nand U51 (N_51,In_1023,In_119);
nand U52 (N_52,In_917,In_49);
nor U53 (N_53,In_374,In_2256);
nand U54 (N_54,In_2343,In_113);
nor U55 (N_55,In_747,In_1320);
and U56 (N_56,In_1800,In_1868);
xor U57 (N_57,In_1222,In_689);
nor U58 (N_58,In_1234,In_363);
nor U59 (N_59,In_903,In_2398);
and U60 (N_60,In_147,In_2410);
or U61 (N_61,In_781,In_326);
nand U62 (N_62,In_1828,In_803);
nor U63 (N_63,In_613,In_2433);
and U64 (N_64,In_1748,In_1003);
nor U65 (N_65,In_1708,In_404);
and U66 (N_66,In_1713,In_1784);
and U67 (N_67,In_563,In_503);
nor U68 (N_68,In_2113,In_601);
nor U69 (N_69,In_90,In_1738);
and U70 (N_70,In_982,In_802);
xnor U71 (N_71,In_805,In_2115);
nand U72 (N_72,In_1539,In_2456);
xor U73 (N_73,In_1047,In_1409);
nor U74 (N_74,In_1015,In_2487);
xnor U75 (N_75,In_341,In_2304);
nand U76 (N_76,In_723,In_826);
and U77 (N_77,In_2015,In_1025);
and U78 (N_78,In_1656,In_30);
or U79 (N_79,In_562,In_2119);
nor U80 (N_80,In_1093,In_1669);
nor U81 (N_81,In_1277,In_3);
or U82 (N_82,In_1942,In_56);
xor U83 (N_83,In_1366,In_1425);
or U84 (N_84,In_1958,In_1024);
nand U85 (N_85,In_51,In_1152);
nand U86 (N_86,In_1395,In_1731);
nor U87 (N_87,In_463,In_2326);
and U88 (N_88,In_1084,In_1755);
nand U89 (N_89,In_1767,In_814);
xnor U90 (N_90,In_1916,In_875);
xor U91 (N_91,In_1410,In_2154);
and U92 (N_92,In_2152,In_2394);
nand U93 (N_93,In_857,In_1008);
and U94 (N_94,In_966,In_2210);
xor U95 (N_95,In_429,In_2238);
and U96 (N_96,In_846,In_817);
and U97 (N_97,In_1485,In_1974);
xor U98 (N_98,In_2126,In_53);
and U99 (N_99,In_50,In_582);
xnor U100 (N_100,In_2325,In_1636);
xor U101 (N_101,In_2314,In_1690);
xor U102 (N_102,In_1351,In_2240);
nand U103 (N_103,In_904,In_958);
nor U104 (N_104,In_118,In_255);
nor U105 (N_105,In_1297,In_612);
nand U106 (N_106,In_440,In_1112);
and U107 (N_107,In_1117,In_384);
or U108 (N_108,In_605,In_842);
and U109 (N_109,In_899,In_1468);
xnor U110 (N_110,In_224,In_614);
and U111 (N_111,In_996,In_1643);
nor U112 (N_112,In_2013,In_711);
or U113 (N_113,In_287,In_598);
or U114 (N_114,In_1430,In_898);
nor U115 (N_115,In_1728,In_1332);
or U116 (N_116,In_866,In_372);
nand U117 (N_117,In_1081,In_1457);
and U118 (N_118,In_2089,In_716);
xnor U119 (N_119,In_247,In_577);
or U120 (N_120,In_1875,In_158);
nor U121 (N_121,In_1927,In_1106);
nand U122 (N_122,In_952,In_496);
nor U123 (N_123,In_1786,In_1306);
nand U124 (N_124,In_478,In_2423);
or U125 (N_125,In_1872,In_2367);
nand U126 (N_126,In_2370,In_1413);
or U127 (N_127,In_2083,In_532);
nor U128 (N_128,In_408,In_991);
nand U129 (N_129,In_123,In_1290);
xor U130 (N_130,In_1119,In_546);
xor U131 (N_131,In_1493,In_334);
nor U132 (N_132,In_2359,In_784);
and U133 (N_133,In_2142,In_986);
nand U134 (N_134,In_1995,In_1953);
and U135 (N_135,In_1519,In_342);
xnor U136 (N_136,In_1302,In_1861);
xor U137 (N_137,In_799,In_1596);
and U138 (N_138,In_892,In_2234);
or U139 (N_139,In_2194,In_1406);
xor U140 (N_140,In_68,In_362);
nand U141 (N_141,In_1807,In_455);
xor U142 (N_142,In_2138,In_391);
nand U143 (N_143,In_238,In_1857);
nand U144 (N_144,In_1951,In_2150);
nor U145 (N_145,In_1651,In_551);
and U146 (N_146,In_1253,In_2352);
xnor U147 (N_147,In_1764,In_1588);
xor U148 (N_148,In_2022,In_967);
or U149 (N_149,In_1216,In_2200);
xor U150 (N_150,In_137,In_84);
and U151 (N_151,In_1328,In_617);
nand U152 (N_152,In_1097,In_969);
nand U153 (N_153,In_1945,In_1167);
nor U154 (N_154,In_1355,In_1029);
or U155 (N_155,In_311,In_37);
or U156 (N_156,In_1369,In_1219);
nand U157 (N_157,In_1173,In_416);
nor U158 (N_158,In_2146,In_99);
nor U159 (N_159,In_1685,In_2086);
or U160 (N_160,In_1211,In_960);
nand U161 (N_161,In_1512,In_253);
and U162 (N_162,In_2269,In_2253);
nand U163 (N_163,In_2415,In_1455);
or U164 (N_164,In_951,In_43);
or U165 (N_165,In_2084,In_797);
nor U166 (N_166,In_21,In_1019);
xnor U167 (N_167,In_499,In_2262);
nand U168 (N_168,In_2267,In_1391);
and U169 (N_169,In_1223,In_1985);
xnor U170 (N_170,In_2176,In_2346);
xor U171 (N_171,In_446,In_2491);
and U172 (N_172,In_2090,In_970);
xor U173 (N_173,In_1091,In_1360);
nand U174 (N_174,In_1809,In_1675);
or U175 (N_175,In_516,In_316);
or U176 (N_176,In_299,In_1061);
xnor U177 (N_177,In_8,In_1885);
and U178 (N_178,In_2289,In_176);
nand U179 (N_179,In_1315,In_434);
nor U180 (N_180,In_1703,In_949);
or U181 (N_181,In_2364,In_432);
nand U182 (N_182,In_631,In_2206);
nand U183 (N_183,In_200,In_2403);
and U184 (N_184,In_111,In_1200);
nor U185 (N_185,In_1978,In_2192);
and U186 (N_186,In_1072,In_191);
xor U187 (N_187,In_1255,In_1460);
nand U188 (N_188,In_2486,In_1611);
or U189 (N_189,In_1531,In_500);
nand U190 (N_190,In_448,In_1578);
xnor U191 (N_191,In_1935,In_2496);
nor U192 (N_192,In_216,In_957);
nor U193 (N_193,In_2024,In_1359);
nor U194 (N_194,In_1915,In_366);
and U195 (N_195,In_356,In_548);
or U196 (N_196,In_804,In_798);
nand U197 (N_197,In_758,In_1311);
xor U198 (N_198,In_2258,In_322);
or U199 (N_199,In_242,In_1480);
xor U200 (N_200,In_881,In_593);
nor U201 (N_201,In_488,In_1415);
or U202 (N_202,In_2012,In_869);
nand U203 (N_203,In_679,In_2237);
and U204 (N_204,In_507,In_273);
and U205 (N_205,In_697,In_1839);
nor U206 (N_206,In_2094,In_330);
or U207 (N_207,In_732,In_1462);
or U208 (N_208,In_533,In_567);
and U209 (N_209,In_1647,In_1229);
nand U210 (N_210,In_1478,In_1298);
or U211 (N_211,In_2081,In_201);
nand U212 (N_212,In_1063,In_2072);
and U213 (N_213,In_2429,In_2096);
and U214 (N_214,In_620,In_2439);
nand U215 (N_215,In_1107,In_594);
xor U216 (N_216,In_292,In_5);
and U217 (N_217,In_728,In_743);
nor U218 (N_218,In_1544,In_196);
nand U219 (N_219,In_135,In_1546);
or U220 (N_220,In_1590,In_2328);
and U221 (N_221,In_310,In_1497);
xor U222 (N_222,In_2023,In_257);
nor U223 (N_223,In_1579,In_2475);
nand U224 (N_224,In_2362,In_1141);
or U225 (N_225,In_1765,In_1659);
nand U226 (N_226,In_108,In_2034);
xnor U227 (N_227,In_673,In_1775);
nand U228 (N_228,In_1192,In_719);
or U229 (N_229,In_729,In_2103);
xor U230 (N_230,In_1238,In_61);
nand U231 (N_231,In_1598,In_403);
nand U232 (N_232,In_639,In_1472);
nand U233 (N_233,In_2417,In_474);
xnor U234 (N_234,In_1465,In_2165);
nor U235 (N_235,In_11,In_1928);
or U236 (N_236,In_553,In_2467);
nand U237 (N_237,In_1608,In_793);
nand U238 (N_238,In_1274,In_720);
or U239 (N_239,In_771,In_369);
or U240 (N_240,In_888,In_1396);
nor U241 (N_241,In_1631,In_2291);
and U242 (N_242,In_1957,In_1910);
nor U243 (N_243,In_169,In_1130);
nand U244 (N_244,In_1550,In_710);
nor U245 (N_245,In_1944,In_355);
or U246 (N_246,In_1754,In_406);
nor U247 (N_247,In_1232,In_444);
nor U248 (N_248,In_782,In_1496);
nand U249 (N_249,In_1416,In_1248);
nand U250 (N_250,In_486,In_17);
and U251 (N_251,In_214,In_1028);
xor U252 (N_252,In_1210,In_1966);
xor U253 (N_253,In_428,In_1812);
nand U254 (N_254,In_632,In_1291);
xnor U255 (N_255,In_934,In_636);
or U256 (N_256,In_1421,In_570);
nor U257 (N_257,In_2177,In_2260);
and U258 (N_258,In_1847,In_942);
xor U259 (N_259,In_1445,In_762);
and U260 (N_260,In_926,In_2422);
nor U261 (N_261,In_1503,In_2116);
nor U262 (N_262,In_289,In_343);
nor U263 (N_263,In_1118,In_1278);
or U264 (N_264,In_1494,In_761);
nand U265 (N_265,In_1894,In_911);
or U266 (N_266,In_62,In_1640);
or U267 (N_267,In_1993,In_608);
and U268 (N_268,In_703,In_1766);
nand U269 (N_269,In_1515,In_886);
nand U270 (N_270,In_910,In_1664);
nand U271 (N_271,In_735,In_410);
or U272 (N_272,In_1433,In_1862);
xnor U273 (N_273,In_1403,In_1004);
nor U274 (N_274,In_2425,In_1076);
xor U275 (N_275,In_143,In_749);
nor U276 (N_276,In_419,In_2205);
and U277 (N_277,In_1001,In_1197);
xor U278 (N_278,In_1155,In_1481);
nand U279 (N_279,In_1573,In_2051);
xnor U280 (N_280,In_2391,In_1895);
xnor U281 (N_281,In_1536,In_1134);
and U282 (N_282,In_360,In_331);
nor U283 (N_283,In_979,In_742);
nand U284 (N_284,In_1123,In_2479);
or U285 (N_285,In_23,In_436);
xor U286 (N_286,In_513,In_439);
nor U287 (N_287,In_1920,In_447);
xor U288 (N_288,In_1148,In_1422);
and U289 (N_289,In_1735,In_752);
xnor U290 (N_290,In_2492,In_597);
xor U291 (N_291,In_1370,In_351);
nand U292 (N_292,In_1498,In_1529);
xnor U293 (N_293,In_2058,In_1792);
and U294 (N_294,In_642,In_1940);
or U295 (N_295,In_1644,In_915);
nor U296 (N_296,In_1122,In_709);
nand U297 (N_297,In_279,In_1697);
and U298 (N_298,In_1036,In_2451);
nand U299 (N_299,In_859,In_501);
xnor U300 (N_300,In_863,In_1435);
nor U301 (N_301,In_1300,In_988);
nand U302 (N_302,In_1012,In_997);
xor U303 (N_303,In_1090,In_1888);
nand U304 (N_304,In_1301,In_1228);
xnor U305 (N_305,In_1702,In_581);
nor U306 (N_306,In_1750,In_2186);
and U307 (N_307,In_1860,In_1987);
and U308 (N_308,In_340,In_759);
and U309 (N_309,In_1074,In_2278);
xnor U310 (N_310,In_1676,In_1242);
nor U311 (N_311,In_550,In_2466);
nand U312 (N_312,In_2167,In_534);
nand U313 (N_313,In_1668,In_36);
and U314 (N_314,In_1545,In_1844);
xnor U315 (N_315,In_1491,In_1905);
nor U316 (N_316,In_2190,In_338);
nor U317 (N_317,In_600,In_2317);
or U318 (N_318,In_2159,In_1712);
nor U319 (N_319,In_205,In_1217);
xor U320 (N_320,In_2202,In_422);
nor U321 (N_321,In_1401,In_2216);
xnor U322 (N_322,In_1532,In_2098);
nand U323 (N_323,In_1534,In_1674);
and U324 (N_324,In_2033,In_2478);
nor U325 (N_325,In_874,In_2135);
xor U326 (N_326,In_452,In_1372);
and U327 (N_327,In_2482,In_1020);
or U328 (N_328,In_1086,In_1040);
nand U329 (N_329,In_2063,In_2061);
xnor U330 (N_330,In_2408,In_1317);
nand U331 (N_331,In_170,In_1749);
and U332 (N_332,In_1438,In_818);
nand U333 (N_333,In_2,In_1243);
nand U334 (N_334,In_2179,In_2372);
nand U335 (N_335,In_1353,In_1762);
nor U336 (N_336,In_131,In_207);
and U337 (N_337,In_1808,In_1357);
xor U338 (N_338,In_198,In_1981);
or U339 (N_339,In_2211,In_1695);
and U340 (N_340,In_157,In_2373);
and U341 (N_341,In_332,In_1742);
and U342 (N_342,In_2312,In_827);
or U343 (N_343,In_1964,In_1027);
xor U344 (N_344,In_1296,In_1684);
xnor U345 (N_345,In_955,In_811);
and U346 (N_346,In_700,In_1751);
and U347 (N_347,In_1961,In_517);
or U348 (N_348,In_2108,In_2353);
nor U349 (N_349,In_2169,In_2386);
nand U350 (N_350,In_1058,In_458);
and U351 (N_351,In_1428,In_900);
nor U352 (N_352,In_497,In_664);
nand U353 (N_353,In_1602,In_763);
nor U354 (N_354,In_133,In_510);
xnor U355 (N_355,In_626,In_67);
nand U356 (N_356,In_1477,In_789);
nor U357 (N_357,In_395,In_564);
or U358 (N_358,In_2077,In_2302);
and U359 (N_359,In_107,In_544);
and U360 (N_360,In_136,In_1778);
or U361 (N_361,In_248,In_847);
nand U362 (N_362,In_424,In_2461);
nor U363 (N_363,In_261,In_1042);
nand U364 (N_364,In_1662,In_2100);
nand U365 (N_365,In_106,In_2092);
xnor U366 (N_366,In_890,In_2105);
and U367 (N_367,In_1518,In_1212);
and U368 (N_368,In_2301,In_897);
and U369 (N_369,In_670,In_1789);
xnor U370 (N_370,In_1615,In_554);
nand U371 (N_371,In_409,In_1113);
nand U372 (N_372,In_2266,In_1803);
and U373 (N_373,In_109,In_184);
nor U374 (N_374,In_114,In_725);
nor U375 (N_375,In_695,In_821);
xor U376 (N_376,In_76,In_1752);
xor U377 (N_377,In_1402,In_2436);
or U378 (N_378,In_1272,In_2318);
xor U379 (N_379,In_520,In_865);
and U380 (N_380,In_1543,In_2095);
nor U381 (N_381,In_990,In_2198);
xor U382 (N_382,In_1826,In_354);
nor U383 (N_383,In_1776,In_2404);
and U384 (N_384,In_1831,In_460);
or U385 (N_385,In_1833,In_1876);
and U386 (N_386,In_2313,In_1709);
or U387 (N_387,In_477,In_535);
and U388 (N_388,In_1740,In_877);
nand U389 (N_389,In_329,In_647);
nand U390 (N_390,In_2157,In_574);
and U391 (N_391,In_19,In_2279);
and U392 (N_392,In_365,In_1938);
nor U393 (N_393,In_481,In_2080);
or U394 (N_394,In_1194,In_1718);
or U395 (N_395,In_138,In_381);
or U396 (N_396,In_203,In_1879);
xor U397 (N_397,In_2184,In_1021);
nand U398 (N_398,In_168,In_2463);
xnor U399 (N_399,In_2383,In_1982);
nor U400 (N_400,In_901,In_15);
or U401 (N_401,In_524,In_1069);
nor U402 (N_402,In_838,In_1941);
nand U403 (N_403,In_1492,In_1185);
nand U404 (N_404,In_1707,In_920);
nor U405 (N_405,In_150,In_197);
nor U406 (N_406,In_1663,In_690);
and U407 (N_407,In_1479,In_1840);
and U408 (N_408,In_1680,In_280);
and U409 (N_409,In_2032,In_1250);
xnor U410 (N_410,In_2172,In_2384);
nand U411 (N_411,In_2280,In_1568);
and U412 (N_412,In_1429,In_389);
xor U413 (N_413,In_2356,In_1323);
or U414 (N_414,In_1172,In_820);
xor U415 (N_415,In_1555,In_2007);
and U416 (N_416,In_1612,In_375);
xor U417 (N_417,In_1976,In_2204);
xor U418 (N_418,In_1973,In_1537);
and U419 (N_419,In_1098,In_1347);
or U420 (N_420,In_1078,In_2474);
and U421 (N_421,In_44,In_1379);
nand U422 (N_422,In_1411,In_2321);
and U423 (N_423,In_1569,In_41);
xor U424 (N_424,In_2286,In_1960);
xor U425 (N_425,In_1770,In_1617);
or U426 (N_426,In_1334,In_515);
or U427 (N_427,In_1863,In_1346);
and U428 (N_428,In_940,In_1774);
xor U429 (N_429,In_1161,In_2283);
nor U430 (N_430,In_560,In_259);
or U431 (N_431,In_1135,In_69);
nand U432 (N_432,In_2239,In_245);
or U433 (N_433,In_649,In_1925);
or U434 (N_434,In_2068,In_2164);
nand U435 (N_435,In_2350,In_298);
nor U436 (N_436,In_1557,In_2246);
nor U437 (N_437,In_523,In_2495);
or U438 (N_438,In_1085,In_202);
xor U439 (N_439,In_1837,In_645);
xor U440 (N_440,In_740,In_206);
and U441 (N_441,In_2327,In_656);
nand U442 (N_442,In_1947,In_2339);
or U443 (N_443,In_2221,In_640);
nand U444 (N_444,In_1610,In_421);
nor U445 (N_445,In_183,In_1144);
xor U446 (N_446,In_1454,In_870);
and U447 (N_447,In_1132,In_660);
and U448 (N_448,In_1870,In_12);
nand U449 (N_449,In_2497,In_1000);
nor U450 (N_450,In_1109,In_2059);
xor U451 (N_451,In_2195,In_1902);
xor U452 (N_452,In_1089,In_2220);
xnor U453 (N_453,In_336,In_94);
nand U454 (N_454,In_2295,In_215);
or U455 (N_455,In_707,In_1698);
xnor U456 (N_456,In_2104,In_575);
nor U457 (N_457,In_156,In_1723);
nand U458 (N_458,In_992,In_1388);
nor U459 (N_459,In_675,In_1225);
or U460 (N_460,In_1714,In_1521);
or U461 (N_461,In_58,In_1830);
and U462 (N_462,In_213,In_1715);
or U463 (N_463,In_2021,In_572);
nor U464 (N_464,In_1,In_335);
and U465 (N_465,In_1205,In_918);
and U466 (N_466,In_1073,In_1358);
and U467 (N_467,In_536,In_175);
nor U468 (N_468,In_2387,In_858);
xnor U469 (N_469,In_687,In_348);
xnor U470 (N_470,In_2122,In_177);
and U471 (N_471,In_1653,In_518);
nor U472 (N_472,In_2399,In_1777);
and U473 (N_473,In_223,In_1287);
and U474 (N_474,In_1198,In_81);
nor U475 (N_475,In_18,In_1886);
and U476 (N_476,In_453,In_1158);
and U477 (N_477,In_285,In_263);
nor U478 (N_478,In_978,In_1609);
xnor U479 (N_479,In_1510,In_980);
nor U480 (N_480,In_2070,In_1585);
or U481 (N_481,In_1045,In_661);
or U482 (N_482,In_2292,In_624);
nor U483 (N_483,In_1279,In_1574);
or U484 (N_484,In_1570,In_293);
nand U485 (N_485,In_417,In_823);
and U486 (N_486,In_2255,In_530);
xnor U487 (N_487,In_315,In_361);
nand U488 (N_488,In_2121,In_1240);
and U489 (N_489,In_1845,In_317);
nor U490 (N_490,In_2274,In_674);
and U491 (N_491,In_71,In_909);
nand U492 (N_492,In_1991,In_1825);
xnor U493 (N_493,In_2131,In_1790);
xor U494 (N_494,In_88,In_1005);
xnor U495 (N_495,In_2323,In_508);
or U496 (N_496,In_1199,In_1948);
or U497 (N_497,In_2257,In_1393);
nand U498 (N_498,In_93,In_1952);
or U499 (N_499,In_1881,In_1067);
xor U500 (N_500,In_922,In_1431);
xor U501 (N_501,In_1405,In_2344);
nor U502 (N_502,In_1031,In_1427);
and U503 (N_503,In_2450,In_2380);
xor U504 (N_504,In_2432,In_678);
and U505 (N_505,In_2201,In_1619);
nor U506 (N_506,In_1377,In_1453);
nand U507 (N_507,In_2476,In_392);
nand U508 (N_508,In_2249,In_2360);
or U509 (N_509,In_1852,In_924);
nor U510 (N_510,In_295,In_1052);
or U511 (N_511,In_1760,In_2203);
or U512 (N_512,In_699,In_1711);
nor U513 (N_513,In_1154,In_1147);
nand U514 (N_514,In_1408,In_1542);
and U515 (N_515,In_2049,In_2430);
xnor U516 (N_516,In_1526,In_2259);
xor U517 (N_517,In_2128,In_1009);
nand U518 (N_518,In_130,In_2300);
xor U519 (N_519,In_1175,In_164);
nand U520 (N_520,In_125,In_646);
nor U521 (N_521,In_1517,In_1127);
and U522 (N_522,In_1145,In_1461);
and U523 (N_523,In_1835,In_873);
nand U524 (N_524,In_835,In_396);
or U525 (N_525,In_368,In_1832);
nand U526 (N_526,In_914,In_1180);
nand U527 (N_527,In_2355,In_1096);
nor U528 (N_528,In_989,In_225);
nand U529 (N_529,In_1151,In_2148);
xnor U530 (N_530,In_1330,In_357);
and U531 (N_531,In_219,In_2139);
nand U532 (N_532,In_1782,In_2050);
or U533 (N_533,In_1083,In_1996);
nand U534 (N_534,In_265,In_1068);
and U535 (N_535,In_2055,In_939);
or U536 (N_536,In_296,In_2390);
nand U537 (N_537,In_473,In_1989);
nand U538 (N_538,In_1691,In_1587);
or U539 (N_539,In_1992,In_1898);
nand U540 (N_540,In_126,In_1022);
and U541 (N_541,In_1524,In_1576);
xor U542 (N_542,In_2006,In_2245);
or U543 (N_543,In_2307,In_1094);
xnor U544 (N_544,In_1082,In_449);
or U545 (N_545,In_2188,In_1525);
or U546 (N_546,In_1246,In_2064);
and U547 (N_547,In_1303,In_537);
and U548 (N_548,In_1704,In_1417);
or U549 (N_549,In_2079,In_227);
nand U550 (N_550,In_1681,In_1439);
nor U551 (N_551,In_2110,In_1033);
and U552 (N_552,In_2143,In_461);
or U553 (N_553,In_808,In_769);
or U554 (N_554,In_1099,In_182);
xor U555 (N_555,In_1160,In_995);
xnor U556 (N_556,In_794,In_2168);
nand U557 (N_557,In_1384,In_2485);
nor U558 (N_558,In_2401,In_1464);
nand U559 (N_559,In_144,In_1324);
nand U560 (N_560,In_1917,In_977);
nand U561 (N_561,In_994,In_971);
xor U562 (N_562,In_65,In_2406);
xnor U563 (N_563,In_2231,In_1580);
xor U564 (N_564,In_953,In_92);
nor U565 (N_565,In_1686,In_584);
nand U566 (N_566,In_1489,In_1514);
nor U567 (N_567,In_1939,In_876);
or U568 (N_568,In_1934,In_1361);
nand U569 (N_569,In_1245,In_1980);
nand U570 (N_570,In_1584,In_659);
nor U571 (N_571,In_1983,In_1797);
nor U572 (N_572,In_324,In_35);
nor U573 (N_573,In_1269,In_1289);
nand U574 (N_574,In_1744,In_465);
nand U575 (N_575,In_845,In_1564);
and U576 (N_576,In_1900,In_837);
and U577 (N_577,In_1710,In_843);
nor U578 (N_578,In_2494,In_34);
nor U579 (N_579,In_806,In_339);
nand U580 (N_580,In_864,In_987);
and U581 (N_581,In_1930,In_1247);
or U582 (N_582,In_2112,In_1010);
or U583 (N_583,In_194,In_1440);
xnor U584 (N_584,In_179,In_1162);
nand U585 (N_585,In_2016,In_1380);
nand U586 (N_586,In_1563,In_451);
xnor U587 (N_587,In_1642,In_834);
or U588 (N_588,In_1387,In_1858);
or U589 (N_589,In_964,In_1006);
or U590 (N_590,In_2392,In_1997);
nor U591 (N_591,In_2263,In_1788);
or U592 (N_592,In_1463,In_1367);
nor U593 (N_593,In_32,In_89);
or U594 (N_594,In_2054,In_962);
or U595 (N_595,In_1108,In_2462);
nand U596 (N_596,In_2099,In_1719);
and U597 (N_597,In_976,In_1195);
nor U598 (N_598,In_1442,In_1678);
nor U599 (N_599,In_1968,In_1635);
nand U600 (N_600,In_1577,In_1268);
and U601 (N_601,In_1513,In_1092);
and U602 (N_602,In_1854,In_1582);
and U603 (N_603,In_155,In_394);
nor U604 (N_604,In_2224,In_941);
xor U605 (N_605,In_2296,In_2270);
nor U606 (N_606,In_592,In_2219);
nor U607 (N_607,In_963,In_1541);
and U608 (N_608,In_724,In_1914);
and U609 (N_609,In_1319,In_1745);
or U610 (N_610,In_2374,In_933);
and U611 (N_611,In_120,In_777);
or U612 (N_612,In_2078,In_1793);
nor U613 (N_613,In_2273,In_1412);
nor U614 (N_614,In_427,In_55);
and U615 (N_615,In_1060,In_66);
nor U616 (N_616,In_59,In_445);
or U617 (N_617,In_1768,In_2427);
xnor U618 (N_618,In_1652,In_736);
nor U619 (N_619,In_1037,In_110);
nor U620 (N_620,In_1679,In_2019);
nor U621 (N_621,In_583,In_217);
xnor U622 (N_622,In_433,In_294);
and U623 (N_623,In_912,In_561);
and U624 (N_624,In_1352,In_1648);
and U625 (N_625,In_891,In_772);
nor U626 (N_626,In_1561,In_2120);
xor U627 (N_627,In_1314,In_349);
or U628 (N_628,In_27,In_87);
and U629 (N_629,In_1115,In_321);
nand U630 (N_630,In_320,In_2371);
and U631 (N_631,In_1120,In_2178);
nand U632 (N_632,In_2144,In_2389);
xnor U633 (N_633,In_252,In_1943);
or U634 (N_634,In_2187,In_2041);
xor U635 (N_635,In_1589,In_829);
xor U636 (N_636,In_181,In_704);
xnor U637 (N_637,In_738,In_333);
xnor U638 (N_638,In_482,In_1507);
nand U639 (N_639,In_1390,In_905);
or U640 (N_640,In_1111,In_1164);
nand U641 (N_641,In_531,In_24);
or U642 (N_642,In_383,In_558);
nand U643 (N_643,In_1450,In_1252);
xnor U644 (N_644,In_1689,In_812);
or U645 (N_645,In_1385,In_393);
nor U646 (N_646,In_1834,In_1528);
or U647 (N_647,In_1383,In_300);
and U648 (N_648,In_275,In_730);
nor U649 (N_649,In_254,In_1979);
or U650 (N_650,In_2297,In_502);
or U651 (N_651,In_1955,In_286);
or U652 (N_652,In_1283,In_1634);
nor U653 (N_653,In_230,In_2303);
xor U654 (N_654,In_7,In_188);
nand U655 (N_655,In_1110,In_2191);
or U656 (N_656,In_9,In_816);
xor U657 (N_657,In_2347,In_1271);
nand U658 (N_658,In_1077,In_662);
nand U659 (N_659,In_1867,In_425);
nor U660 (N_660,In_48,In_2293);
nand U661 (N_661,In_1853,In_786);
or U662 (N_662,In_2132,In_1038);
nor U663 (N_663,In_229,In_1329);
and U664 (N_664,In_2130,In_204);
nor U665 (N_665,In_618,In_222);
nand U666 (N_666,In_1907,In_1694);
and U667 (N_667,In_1586,In_950);
or U668 (N_668,In_815,In_961);
nand U669 (N_669,In_2305,In_824);
nor U670 (N_670,In_456,In_1806);
nand U671 (N_671,In_174,In_1236);
or U672 (N_672,In_1449,In_2284);
nor U673 (N_673,In_1182,In_2298);
nand U674 (N_674,In_521,In_1827);
nor U675 (N_675,In_2133,In_210);
and U676 (N_676,In_2413,In_652);
xnor U677 (N_677,In_556,In_1142);
or U678 (N_678,In_1321,In_97);
or U679 (N_679,In_2226,In_1138);
and U680 (N_680,In_2337,In_737);
nor U681 (N_681,In_2140,In_1984);
xnor U682 (N_682,In_1044,In_2189);
nor U683 (N_683,In_1013,In_438);
or U684 (N_684,In_1203,In_122);
and U685 (N_685,In_872,In_1871);
and U686 (N_686,In_2046,In_1670);
xor U687 (N_687,In_2087,In_512);
xnor U688 (N_688,In_1904,In_1350);
nor U689 (N_689,In_2421,In_1994);
nand U690 (N_690,In_667,In_1554);
xor U691 (N_691,In_83,In_2014);
or U692 (N_692,In_2332,In_999);
nand U693 (N_693,In_1448,In_2446);
nor U694 (N_694,In_350,In_1382);
nor U695 (N_695,In_218,In_2342);
and U696 (N_696,In_655,In_2196);
or U697 (N_697,In_359,In_2418);
nor U698 (N_698,In_407,In_511);
and U699 (N_699,In_589,In_309);
nand U700 (N_700,In_454,In_237);
xor U701 (N_701,In_239,In_1065);
nor U702 (N_702,In_2225,In_2003);
nand U703 (N_703,In_1104,In_882);
nand U704 (N_704,In_1365,In_1150);
nand U705 (N_705,In_685,In_801);
xor U706 (N_706,In_1855,In_258);
and U707 (N_707,In_1178,In_146);
or U708 (N_708,In_965,In_671);
and U709 (N_709,In_2042,In_2228);
xnor U710 (N_710,In_919,In_2163);
or U711 (N_711,In_1432,In_727);
xnor U712 (N_712,In_790,In_1312);
nand U713 (N_713,In_1486,In_1444);
and U714 (N_714,In_2357,In_1102);
nand U715 (N_715,In_2162,In_956);
and U716 (N_716,In_1201,In_153);
xor U717 (N_717,In_607,In_2288);
nor U718 (N_718,In_2074,In_2158);
or U719 (N_719,In_2331,In_60);
xor U720 (N_720,In_2282,In_1345);
xnor U721 (N_721,In_2027,In_2137);
nand U722 (N_722,In_1343,In_1482);
nand U723 (N_723,In_1932,In_2490);
xnor U724 (N_724,In_2431,In_1179);
nor U725 (N_725,In_492,In_494);
xnor U726 (N_726,In_104,In_1629);
or U727 (N_727,In_272,In_149);
or U728 (N_728,In_462,In_498);
and U729 (N_729,In_2407,In_1874);
and U730 (N_730,In_1376,In_2464);
nand U731 (N_731,In_4,In_2277);
nand U732 (N_732,In_1658,In_590);
nor U733 (N_733,In_1547,In_2125);
nor U734 (N_734,In_134,In_1869);
xnor U735 (N_735,In_102,In_929);
nand U736 (N_736,In_1473,In_457);
or U737 (N_737,In_152,In_25);
nor U738 (N_738,In_916,In_1878);
xnor U739 (N_739,In_2477,In_833);
and U740 (N_740,In_637,In_2316);
nand U741 (N_741,In_2170,In_1055);
nand U742 (N_742,In_1344,In_1215);
xor U743 (N_743,In_676,In_2445);
nor U744 (N_744,In_2197,In_471);
and U745 (N_745,In_1340,In_2306);
and U746 (N_746,In_1729,In_1451);
nor U747 (N_747,In_1266,In_2414);
nor U748 (N_748,In_1267,In_756);
nor U749 (N_749,In_947,In_1121);
and U750 (N_750,In_1034,In_549);
nand U751 (N_751,In_2271,In_1282);
or U752 (N_752,In_430,In_1667);
xnor U753 (N_753,In_764,In_2376);
nand U754 (N_754,In_1139,In_1049);
and U755 (N_755,In_785,In_1285);
or U756 (N_756,In_271,In_2069);
or U757 (N_757,In_1308,In_1338);
and U758 (N_758,In_212,In_1923);
and U759 (N_759,In_1552,In_1397);
nand U760 (N_760,In_854,In_2010);
xnor U761 (N_761,In_208,In_1657);
and U762 (N_762,In_483,In_117);
nand U763 (N_763,In_1956,In_1739);
nor U764 (N_764,In_1891,In_1459);
nor U765 (N_765,In_1504,In_1820);
and U766 (N_766,In_1661,In_1780);
nand U767 (N_767,In_2471,In_879);
and U768 (N_768,In_1890,In_405);
nor U769 (N_769,In_1420,In_609);
or U770 (N_770,In_871,In_1424);
and U771 (N_771,In_2199,In_145);
or U772 (N_772,In_1458,In_1176);
xnor U773 (N_773,In_2043,In_1761);
or U774 (N_774,In_541,In_1349);
or U775 (N_775,In_1261,In_345);
or U776 (N_776,In_412,In_1284);
nor U777 (N_777,In_387,In_1551);
and U778 (N_778,In_2493,In_1466);
nor U779 (N_779,In_1373,In_1389);
xnor U780 (N_780,In_47,In_1169);
nor U781 (N_781,In_1275,In_1548);
and U782 (N_782,In_1398,In_1924);
nand U783 (N_783,In_2002,In_1404);
or U784 (N_784,In_1535,In_1183);
nand U785 (N_785,In_2000,In_1331);
and U786 (N_786,In_127,In_161);
or U787 (N_787,In_270,In_2333);
nor U788 (N_788,In_2229,In_450);
or U789 (N_789,In_2315,In_306);
nor U790 (N_790,In_1795,In_775);
or U791 (N_791,In_741,In_2469);
nor U792 (N_792,In_691,In_91);
and U793 (N_793,In_930,In_538);
nor U794 (N_794,In_896,In_1230);
nand U795 (N_795,In_2483,In_1693);
xnor U796 (N_796,In_1990,In_1889);
and U797 (N_797,In_1600,In_431);
nand U798 (N_798,In_2330,In_682);
and U799 (N_799,In_1965,In_1873);
or U800 (N_800,In_807,In_1333);
nand U801 (N_801,In_1500,In_1506);
or U802 (N_802,In_2053,In_193);
or U803 (N_803,In_973,In_1733);
xnor U804 (N_804,In_1214,In_1625);
nand U805 (N_805,In_1189,In_1313);
xor U806 (N_806,In_840,In_1262);
and U807 (N_807,In_353,In_1011);
and U808 (N_808,In_868,In_1660);
nand U809 (N_809,In_1838,In_160);
nand U810 (N_810,In_861,In_625);
and U811 (N_811,In_998,In_755);
nand U812 (N_812,In_1163,In_569);
xnor U813 (N_813,In_792,In_526);
and U814 (N_814,In_766,In_2093);
xor U815 (N_815,In_1950,In_1540);
or U816 (N_816,In_1864,In_650);
nand U817 (N_817,In_2025,In_1632);
xnor U818 (N_818,In_666,In_1153);
nor U819 (N_819,In_1769,In_1257);
nand U820 (N_820,In_1511,In_1866);
xnor U821 (N_821,In_1565,In_1562);
and U822 (N_822,In_1814,In_1204);
or U823 (N_823,In_717,In_2395);
or U824 (N_824,In_1342,In_1177);
xor U825 (N_825,In_2311,In_1665);
nor U826 (N_826,In_1621,In_493);
or U827 (N_827,In_2473,In_1599);
and U828 (N_828,In_1307,In_2275);
and U829 (N_829,In_303,In_555);
and U830 (N_830,In_1906,In_1251);
or U831 (N_831,In_64,In_1400);
or U832 (N_832,In_1883,In_1273);
nand U833 (N_833,In_819,In_1682);
nor U834 (N_834,In_1783,In_318);
and U835 (N_835,In_681,In_721);
or U836 (N_836,In_1791,In_2480);
or U837 (N_837,In_2111,In_2419);
xor U838 (N_838,In_1337,In_2379);
or U839 (N_839,In_770,In_1641);
nor U840 (N_840,In_1856,In_278);
nand U841 (N_841,In_1841,In_677);
nand U842 (N_842,In_1556,In_29);
xor U843 (N_843,In_1597,In_2366);
xnor U844 (N_844,In_1280,In_2222);
nand U845 (N_845,In_1071,In_162);
xnor U846 (N_846,In_1743,In_972);
or U847 (N_847,In_2149,In_2106);
or U848 (N_848,In_1156,In_851);
and U849 (N_849,In_2129,In_935);
or U850 (N_850,In_1732,In_1884);
nor U851 (N_851,In_1527,In_1977);
and U852 (N_852,In_2320,In_2045);
xor U853 (N_853,In_378,In_2242);
and U854 (N_854,In_2217,In_731);
nor U855 (N_855,In_1763,In_1399);
and U856 (N_856,In_1700,In_1779);
and U857 (N_857,In_312,In_665);
and U858 (N_858,In_974,In_1931);
or U859 (N_859,In_40,In_585);
or U860 (N_860,In_932,In_765);
nand U861 (N_861,In_778,In_1630);
and U862 (N_862,In_1362,In_2232);
and U863 (N_863,In_2272,In_908);
and U864 (N_864,In_1050,In_788);
nand U865 (N_865,In_2117,In_2151);
nand U866 (N_866,In_95,In_2381);
or U867 (N_867,In_1818,In_1184);
or U868 (N_868,In_688,In_1143);
nor U869 (N_869,In_1374,In_1483);
nor U870 (N_870,In_855,In_1474);
xnor U871 (N_871,In_1281,In_587);
xnor U872 (N_872,In_337,In_1218);
or U873 (N_873,In_2388,In_2349);
nand U874 (N_874,In_1919,In_2308);
xnor U875 (N_875,In_2247,In_443);
nand U876 (N_876,In_2124,In_1655);
and U877 (N_877,In_2067,In_63);
and U878 (N_878,In_2004,In_46);
or U879 (N_879,In_1717,In_780);
xnor U880 (N_880,In_442,In_1075);
nand U881 (N_881,In_525,In_413);
nor U882 (N_882,In_1186,In_1613);
and U883 (N_883,In_2438,In_2039);
xnor U884 (N_884,In_1949,In_249);
or U885 (N_885,In_1341,In_895);
nand U886 (N_886,In_884,In_1487);
xor U887 (N_887,In_1294,In_894);
nor U888 (N_888,In_1418,In_1456);
or U889 (N_889,In_1035,In_604);
nor U890 (N_890,In_2402,In_246);
nor U891 (N_891,In_98,In_633);
nor U892 (N_892,In_1520,In_1196);
or U893 (N_893,In_1348,In_297);
or U894 (N_894,In_491,In_1901);
nand U895 (N_895,In_1558,In_85);
nor U896 (N_896,In_2241,In_680);
and U897 (N_897,In_2470,In_2261);
xor U898 (N_898,In_1128,In_314);
or U899 (N_899,In_1819,In_1171);
or U900 (N_900,In_1508,In_328);
and U901 (N_901,In_195,In_578);
xor U902 (N_902,In_506,In_327);
nor U903 (N_903,In_1623,In_2319);
xor U904 (N_904,In_2118,In_893);
nor U905 (N_905,In_1231,In_82);
nor U906 (N_906,In_1627,In_757);
or U907 (N_907,In_1688,In_358);
nand U908 (N_908,In_1041,In_276);
and U909 (N_909,In_1759,In_240);
and U910 (N_910,In_1007,In_22);
nor U911 (N_911,In_654,In_634);
and U912 (N_912,In_2382,In_1241);
and U913 (N_913,In_936,In_1811);
nand U914 (N_914,In_1601,In_288);
nor U915 (N_915,In_96,In_1181);
nor U916 (N_916,In_573,In_72);
and U917 (N_917,In_45,In_2062);
nor U918 (N_918,In_399,In_1646);
xnor U919 (N_919,In_1672,In_1286);
nand U920 (N_920,In_469,In_367);
or U921 (N_921,In_1100,In_105);
nor U922 (N_922,In_2056,In_1057);
nor U923 (N_923,In_925,In_487);
and U924 (N_924,In_1207,In_2123);
nand U925 (N_925,In_485,In_2264);
nand U926 (N_926,In_722,In_1392);
and U927 (N_927,In_1467,In_2444);
xor U928 (N_928,In_623,In_559);
nand U929 (N_929,In_1887,In_70);
xnor U930 (N_930,In_1849,In_945);
and U931 (N_931,In_2341,In_100);
nor U932 (N_932,In_1654,In_1963);
or U933 (N_933,In_698,In_571);
nand U934 (N_934,In_2435,In_2489);
or U935 (N_935,In_1581,In_2442);
xnor U936 (N_936,In_1095,In_547);
nor U937 (N_937,In_2047,In_1799);
nand U938 (N_938,In_2037,In_1639);
nor U939 (N_939,In_302,In_653);
or U940 (N_940,In_2145,In_2397);
xnor U941 (N_941,In_103,In_595);
and U942 (N_942,In_576,In_2136);
nor U943 (N_943,In_1605,In_1447);
or U944 (N_944,In_993,In_1785);
nand U945 (N_945,In_2038,In_241);
or U946 (N_946,In_1295,In_1452);
nor U947 (N_947,In_20,In_1798);
or U948 (N_948,In_619,In_2018);
xor U949 (N_949,In_1469,In_2455);
and U950 (N_950,In_1843,In_1484);
xor U951 (N_951,In_1165,In_1962);
and U952 (N_952,In_52,In_1363);
or U953 (N_953,In_1583,In_968);
nor U954 (N_954,In_1490,In_566);
nor U955 (N_955,In_701,In_2396);
or U956 (N_956,In_2268,In_638);
xor U957 (N_957,In_2005,In_1727);
and U958 (N_958,In_591,In_1129);
nand U959 (N_959,In_1501,In_1815);
xor U960 (N_960,In_2065,In_776);
nor U961 (N_961,In_552,In_694);
nand U962 (N_962,In_1824,In_2060);
or U963 (N_963,In_1048,In_466);
nor U964 (N_964,In_2207,In_714);
nand U965 (N_965,In_1053,In_1495);
xor U966 (N_966,In_1292,In_423);
xor U967 (N_967,In_364,In_305);
nand U968 (N_968,In_1614,In_2368);
or U969 (N_969,In_1796,In_2251);
nand U970 (N_970,In_2011,In_1794);
nand U971 (N_971,In_1039,In_414);
xnor U972 (N_972,In_923,In_112);
or U973 (N_973,In_1757,In_2254);
and U974 (N_974,In_1470,In_504);
and U975 (N_975,In_1133,In_1899);
nor U976 (N_976,In_2020,In_1722);
or U977 (N_977,In_1059,In_1265);
nand U978 (N_978,In_1516,In_1032);
nor U979 (N_979,In_1946,In_2230);
nor U980 (N_980,In_2365,In_684);
nor U981 (N_981,In_529,In_522);
or U982 (N_982,In_2393,In_543);
or U983 (N_983,In_1209,In_1126);
or U984 (N_984,In_643,In_148);
xnor U985 (N_985,In_1823,In_1381);
nand U986 (N_986,In_28,In_2017);
xor U987 (N_987,In_2097,In_1730);
and U988 (N_988,In_1736,In_291);
or U989 (N_989,In_621,In_1310);
or U990 (N_990,In_189,In_1969);
nor U991 (N_991,In_519,In_1746);
nor U992 (N_992,In_1882,In_2335);
and U993 (N_993,In_1339,In_373);
nor U994 (N_994,In_1781,In_2001);
nand U995 (N_995,In_713,In_1628);
and U996 (N_996,In_1975,In_2400);
nand U997 (N_997,In_839,In_2340);
nor U998 (N_998,In_860,In_568);
nand U999 (N_999,In_1509,In_1187);
or U1000 (N_1000,In_178,In_141);
and U1001 (N_1001,In_1146,N_990);
nand U1002 (N_1002,In_753,N_189);
or U1003 (N_1003,In_325,N_372);
nor U1004 (N_1004,In_2085,N_610);
or U1005 (N_1005,N_248,In_1592);
nor U1006 (N_1006,N_780,In_1356);
xnor U1007 (N_1007,In_165,N_337);
xor U1008 (N_1008,In_1970,N_379);
xor U1009 (N_1009,In_800,N_487);
nand U1010 (N_1010,N_529,N_109);
nand U1011 (N_1011,N_30,N_844);
and U1012 (N_1012,N_50,In_878);
and U1013 (N_1013,In_1893,N_570);
xor U1014 (N_1014,N_434,N_206);
and U1015 (N_1015,N_985,N_754);
xnor U1016 (N_1016,N_21,In_13);
nand U1017 (N_1017,In_1014,N_286);
nor U1018 (N_1018,N_840,N_751);
and U1019 (N_1019,N_69,N_967);
xor U1020 (N_1020,N_942,N_141);
nand U1021 (N_1021,In_236,N_876);
nor U1022 (N_1022,N_635,N_897);
xor U1023 (N_1023,N_393,In_927);
and U1024 (N_1024,N_224,N_604);
nand U1025 (N_1025,In_2416,In_1737);
nand U1026 (N_1026,In_2294,N_811);
nand U1027 (N_1027,N_165,In_1414);
xnor U1028 (N_1028,In_268,N_386);
nand U1029 (N_1029,N_582,In_2161);
xor U1030 (N_1030,N_166,N_752);
nand U1031 (N_1031,N_258,N_546);
xor U1032 (N_1032,N_228,N_781);
nor U1033 (N_1033,In_79,In_151);
and U1034 (N_1034,In_1030,N_328);
nand U1035 (N_1035,N_830,N_678);
nand U1036 (N_1036,In_376,In_648);
nand U1037 (N_1037,N_605,N_325);
nor U1038 (N_1038,N_525,In_1624);
or U1039 (N_1039,In_1846,In_718);
xor U1040 (N_1040,N_991,N_730);
and U1041 (N_1041,N_647,N_531);
nand U1042 (N_1042,N_9,In_1805);
or U1043 (N_1043,N_798,N_800);
nand U1044 (N_1044,N_571,In_712);
nor U1045 (N_1045,N_187,N_3);
nor U1046 (N_1046,In_2185,In_371);
or U1047 (N_1047,N_958,N_22);
nand U1048 (N_1048,N_824,In_509);
nor U1049 (N_1049,N_979,N_607);
and U1050 (N_1050,N_231,In_1304);
nand U1051 (N_1051,In_1933,N_787);
and U1052 (N_1052,In_274,N_32);
nor U1053 (N_1053,In_74,N_542);
nor U1054 (N_1054,N_164,In_902);
xor U1055 (N_1055,In_1816,N_913);
and U1056 (N_1056,N_756,In_1880);
and U1057 (N_1057,N_191,In_231);
xnor U1058 (N_1058,In_708,N_223);
and U1059 (N_1059,N_322,N_335);
nor U1060 (N_1060,In_1701,In_774);
and U1061 (N_1061,N_160,In_128);
nand U1062 (N_1062,In_2453,N_691);
and U1063 (N_1063,N_731,N_359);
or U1064 (N_1064,N_839,N_995);
and U1065 (N_1065,In_1062,In_2156);
nor U1066 (N_1066,In_588,In_1593);
nor U1067 (N_1067,N_956,N_597);
and U1068 (N_1068,In_2375,N_430);
or U1069 (N_1069,In_726,In_2073);
or U1070 (N_1070,In_810,N_974);
nor U1071 (N_1071,N_299,N_457);
nand U1072 (N_1072,N_360,N_274);
nor U1073 (N_1073,In_2412,In_2101);
and U1074 (N_1074,N_867,In_1725);
and U1075 (N_1075,N_528,N_578);
nor U1076 (N_1076,N_220,N_85);
and U1077 (N_1077,N_671,N_616);
or U1078 (N_1078,N_414,In_1821);
nand U1079 (N_1079,N_126,N_447);
nand U1080 (N_1080,N_427,In_1326);
and U1081 (N_1081,N_733,In_495);
nor U1082 (N_1082,N_945,In_1375);
xnor U1083 (N_1083,N_878,N_633);
nand U1084 (N_1084,In_946,N_266);
and U1085 (N_1085,N_855,N_885);
nor U1086 (N_1086,N_433,In_1087);
or U1087 (N_1087,N_947,N_688);
nand U1088 (N_1088,N_930,N_680);
and U1089 (N_1089,In_2075,In_1233);
or U1090 (N_1090,N_177,N_820);
nand U1091 (N_1091,N_676,N_152);
nor U1092 (N_1092,N_895,N_881);
nor U1093 (N_1093,N_481,N_284);
or U1094 (N_1094,In_2076,In_1080);
nor U1095 (N_1095,N_832,In_748);
or U1096 (N_1096,N_298,N_494);
nor U1097 (N_1097,N_342,N_116);
nand U1098 (N_1098,N_724,In_1263);
nor U1099 (N_1099,In_981,N_746);
and U1100 (N_1100,In_610,N_596);
nand U1101 (N_1101,N_460,N_861);
nand U1102 (N_1102,N_240,In_1986);
and U1103 (N_1103,In_1136,In_750);
nor U1104 (N_1104,N_67,N_162);
and U1105 (N_1105,In_186,In_1476);
or U1106 (N_1106,N_426,In_2153);
and U1107 (N_1107,N_216,N_203);
nand U1108 (N_1108,N_768,In_1848);
nand U1109 (N_1109,N_188,N_180);
or U1110 (N_1110,In_2441,N_176);
nor U1111 (N_1111,N_934,N_370);
and U1112 (N_1112,N_743,In_1264);
nand U1113 (N_1113,N_236,N_167);
or U1114 (N_1114,N_685,N_273);
xnor U1115 (N_1115,N_470,N_27);
or U1116 (N_1116,N_163,In_211);
or U1117 (N_1117,N_835,In_686);
nand U1118 (N_1118,N_79,N_559);
xnor U1119 (N_1119,N_239,N_455);
nand U1120 (N_1120,N_399,N_606);
nand U1121 (N_1121,N_723,N_106);
nor U1122 (N_1122,N_617,In_1174);
nand U1123 (N_1123,N_789,N_57);
xnor U1124 (N_1124,N_233,N_437);
nand U1125 (N_1125,N_416,N_194);
nand U1126 (N_1126,N_410,In_644);
nand U1127 (N_1127,N_686,N_874);
nand U1128 (N_1128,N_613,In_796);
or U1129 (N_1129,In_352,N_618);
and U1130 (N_1130,In_1937,N_968);
or U1131 (N_1131,N_52,N_900);
nor U1132 (N_1132,In_1801,N_883);
and U1133 (N_1133,In_2447,N_654);
nor U1134 (N_1134,N_999,N_658);
nor U1135 (N_1135,N_420,In_209);
nand U1136 (N_1136,In_77,In_984);
nor U1137 (N_1137,In_2378,N_518);
nand U1138 (N_1138,In_290,In_2155);
or U1139 (N_1139,N_146,In_1364);
nor U1140 (N_1140,N_125,N_234);
xor U1141 (N_1141,N_716,N_406);
nor U1142 (N_1142,N_879,N_677);
nor U1143 (N_1143,N_476,N_961);
or U1144 (N_1144,N_408,N_212);
and U1145 (N_1145,N_112,In_140);
or U1146 (N_1146,N_612,N_20);
nand U1147 (N_1147,N_290,N_454);
xnor U1148 (N_1148,In_1929,N_963);
nand U1149 (N_1149,In_2363,N_232);
or U1150 (N_1150,N_827,N_615);
nor U1151 (N_1151,N_837,N_681);
nand U1152 (N_1152,N_651,N_438);
nand U1153 (N_1153,In_734,N_23);
nand U1154 (N_1154,N_75,N_173);
nand U1155 (N_1155,In_2454,N_828);
or U1156 (N_1156,N_285,N_415);
or U1157 (N_1157,In_907,In_80);
or U1158 (N_1158,N_375,N_851);
or U1159 (N_1159,N_114,In_2276);
and U1160 (N_1160,N_356,N_564);
or U1161 (N_1161,N_45,In_1443);
or U1162 (N_1162,N_402,In_234);
and U1163 (N_1163,In_2227,N_478);
or U1164 (N_1164,In_2008,N_729);
and U1165 (N_1165,In_630,N_117);
nand U1166 (N_1166,N_648,N_64);
nor U1167 (N_1167,N_380,In_739);
nand U1168 (N_1168,N_252,N_110);
nor U1169 (N_1169,N_770,N_169);
and U1170 (N_1170,N_255,N_100);
xnor U1171 (N_1171,In_1836,N_854);
nand U1172 (N_1172,In_658,In_313);
and U1173 (N_1173,N_297,N_697);
and U1174 (N_1174,N_763,In_1043);
or U1175 (N_1175,N_280,N_905);
nand U1176 (N_1176,N_906,N_857);
nor U1177 (N_1177,N_92,N_89);
nand U1178 (N_1178,N_355,N_504);
and U1179 (N_1179,N_765,N_972);
nor U1180 (N_1180,N_382,N_701);
or U1181 (N_1181,N_692,N_148);
and U1182 (N_1182,In_2420,N_254);
xnor U1183 (N_1183,N_46,N_407);
or U1184 (N_1184,N_432,N_965);
nand U1185 (N_1185,N_706,In_388);
and U1186 (N_1186,In_2361,In_1607);
and U1187 (N_1187,N_818,In_2448);
and U1188 (N_1188,N_367,In_528);
xor U1189 (N_1189,In_57,In_651);
nor U1190 (N_1190,N_514,N_130);
xor U1191 (N_1191,N_804,N_270);
and U1192 (N_1192,In_1522,N_465);
or U1193 (N_1193,N_603,In_400);
nand U1194 (N_1194,In_828,In_2173);
nand U1195 (N_1195,N_541,N_7);
nand U1196 (N_1196,In_867,In_42);
nor U1197 (N_1197,N_184,N_915);
and U1198 (N_1198,N_522,In_627);
nor U1199 (N_1199,In_2091,N_761);
nor U1200 (N_1200,In_415,N_251);
or U1201 (N_1201,N_244,N_91);
and U1202 (N_1202,N_96,N_652);
nand U1203 (N_1203,N_636,N_138);
or U1204 (N_1204,N_534,In_115);
xor U1205 (N_1205,N_667,N_424);
nand U1206 (N_1206,In_1327,N_943);
or U1207 (N_1207,N_575,In_2310);
and U1208 (N_1208,In_2458,N_679);
nor U1209 (N_1209,N_352,In_284);
nor U1210 (N_1210,In_1696,In_2252);
xnor U1211 (N_1211,N_737,N_343);
xnor U1212 (N_1212,N_949,In_1394);
nand U1213 (N_1213,N_93,In_1606);
nand U1214 (N_1214,N_97,N_35);
xnor U1215 (N_1215,In_2472,In_154);
or U1216 (N_1216,N_823,N_859);
nor U1217 (N_1217,N_916,N_826);
nand U1218 (N_1218,In_1190,In_1747);
nand U1219 (N_1219,In_1817,N_361);
nor U1220 (N_1220,N_533,In_1903);
and U1221 (N_1221,N_267,N_750);
xor U1222 (N_1222,N_102,N_941);
or U1223 (N_1223,N_29,N_953);
and U1224 (N_1224,N_278,In_2102);
nor U1225 (N_1225,N_735,N_238);
nand U1226 (N_1226,N_179,N_98);
nand U1227 (N_1227,N_769,N_512);
nand U1228 (N_1228,N_627,N_25);
xnor U1229 (N_1229,N_741,N_49);
nand U1230 (N_1230,In_539,N_799);
xnor U1231 (N_1231,In_1720,N_887);
xor U1232 (N_1232,In_192,In_844);
nor U1233 (N_1233,N_229,N_373);
nand U1234 (N_1234,N_168,N_301);
nand U1235 (N_1235,In_1168,In_1224);
xnor U1236 (N_1236,N_235,In_398);
nand U1237 (N_1237,N_966,N_535);
nor U1238 (N_1238,N_642,N_901);
nor U1239 (N_1239,N_14,N_923);
nor U1240 (N_1240,N_866,In_1972);
nand U1241 (N_1241,N_264,In_1378);
or U1242 (N_1242,N_256,In_1724);
and U1243 (N_1243,N_120,In_308);
or U1244 (N_1244,N_333,N_241);
xor U1245 (N_1245,N_547,In_683);
nand U1246 (N_1246,N_845,In_1446);
or U1247 (N_1247,N_157,N_70);
nand U1248 (N_1248,N_475,N_329);
xnor U1249 (N_1249,N_969,In_187);
or U1250 (N_1250,N_350,N_601);
and U1251 (N_1251,N_124,N_374);
xor U1252 (N_1252,In_1140,In_1213);
xnor U1253 (N_1253,N_272,In_380);
nand U1254 (N_1254,N_12,In_1829);
and U1255 (N_1255,N_53,In_2481);
or U1256 (N_1256,N_918,N_712);
nor U1257 (N_1257,N_803,In_166);
nor U1258 (N_1258,In_1131,N_135);
nor U1259 (N_1259,N_496,N_200);
nand U1260 (N_1260,In_1988,N_421);
and U1261 (N_1261,In_603,In_1208);
nor U1262 (N_1262,N_121,N_326);
and U1263 (N_1263,In_2141,N_912);
xnor U1264 (N_1264,In_78,N_417);
and U1265 (N_1265,In_441,N_592);
nor U1266 (N_1266,N_161,In_1859);
nor U1267 (N_1267,In_1523,In_307);
or U1268 (N_1268,N_60,In_1258);
nor U1269 (N_1269,N_577,N_672);
xnor U1270 (N_1270,N_381,N_33);
nor U1271 (N_1271,In_2338,N_892);
nor U1272 (N_1272,N_338,In_1288);
xor U1273 (N_1273,N_634,N_626);
nand U1274 (N_1274,N_872,N_351);
xor U1275 (N_1275,N_668,N_922);
and U1276 (N_1276,In_931,N_515);
or U1277 (N_1277,N_503,In_390);
nand U1278 (N_1278,N_62,N_491);
xnor U1279 (N_1279,In_2498,N_865);
nand U1280 (N_1280,N_611,N_819);
or U1281 (N_1281,N_246,In_2212);
xor U1282 (N_1282,N_445,In_2107);
or U1283 (N_1283,N_88,In_1191);
nor U1284 (N_1284,N_502,In_2223);
nor U1285 (N_1285,N_181,N_305);
nor U1286 (N_1286,N_580,N_755);
and U1287 (N_1287,N_588,In_751);
nor U1288 (N_1288,N_925,N_468);
nand U1289 (N_1289,N_449,N_140);
nor U1290 (N_1290,N_219,In_2040);
nand U1291 (N_1291,N_566,N_962);
or U1292 (N_1292,N_221,N_624);
nand U1293 (N_1293,In_2180,N_10);
nand U1294 (N_1294,N_2,N_924);
nand U1295 (N_1295,In_1237,In_579);
nand U1296 (N_1296,In_1235,N_183);
and U1297 (N_1297,N_815,N_283);
nand U1298 (N_1298,N_790,In_1538);
xor U1299 (N_1299,N_122,In_2147);
xor U1300 (N_1300,N_703,N_170);
nor U1301 (N_1301,N_719,N_482);
nor U1302 (N_1302,N_732,N_562);
nor U1303 (N_1303,In_1125,In_1016);
nand U1304 (N_1304,N_759,In_101);
nand U1305 (N_1305,N_26,In_635);
or U1306 (N_1306,In_1804,N_920);
or U1307 (N_1307,N_321,In_959);
nor U1308 (N_1308,N_208,N_489);
and U1309 (N_1309,N_107,In_937);
nand U1310 (N_1310,N_767,N_527);
nand U1311 (N_1311,N_599,N_726);
nor U1312 (N_1312,In_1426,N_926);
xnor U1313 (N_1313,N_650,In_983);
nor U1314 (N_1314,In_641,N_341);
nor U1315 (N_1315,N_83,In_1909);
nor U1316 (N_1316,N_975,N_108);
and U1317 (N_1317,N_670,N_536);
nand U1318 (N_1318,N_0,N_142);
nand U1319 (N_1319,In_599,In_1502);
nand U1320 (N_1320,In_480,N_401);
and U1321 (N_1321,N_453,N_707);
xnor U1322 (N_1322,N_809,N_282);
or U1323 (N_1323,In_1101,N_419);
xnor U1324 (N_1324,N_838,N_47);
and U1325 (N_1325,N_911,In_2287);
or U1326 (N_1326,In_1026,N_981);
or U1327 (N_1327,In_2443,N_257);
or U1328 (N_1328,N_492,In_1572);
or U1329 (N_1329,N_847,N_795);
nand U1330 (N_1330,N_538,N_622);
or U1331 (N_1331,N_131,N_269);
and U1332 (N_1332,N_806,N_526);
or U1333 (N_1333,In_668,N_291);
xor U1334 (N_1334,N_620,In_256);
and U1335 (N_1335,N_391,In_1959);
xor U1336 (N_1336,In_841,In_437);
or U1337 (N_1337,In_1054,N_581);
nand U1338 (N_1338,In_1305,N_472);
nand U1339 (N_1339,N_144,N_65);
nand U1340 (N_1340,N_714,N_51);
nor U1341 (N_1341,N_779,N_349);
xor U1342 (N_1342,N_158,N_657);
and U1343 (N_1343,N_193,N_663);
nor U1344 (N_1344,N_971,N_345);
nor U1345 (N_1345,N_662,N_311);
or U1346 (N_1346,N_946,N_182);
and U1347 (N_1347,In_527,In_889);
and U1348 (N_1348,In_39,N_630);
and U1349 (N_1349,N_507,N_268);
nor U1350 (N_1350,In_1017,In_1371);
nor U1351 (N_1351,In_385,N_682);
or U1352 (N_1352,In_2035,In_124);
xnor U1353 (N_1353,N_858,N_940);
or U1354 (N_1354,In_1549,In_2440);
and U1355 (N_1355,In_262,N_5);
nand U1356 (N_1356,In_1249,N_499);
and U1357 (N_1357,In_1908,N_293);
nor U1358 (N_1358,N_978,N_99);
nor U1359 (N_1359,N_888,N_175);
or U1360 (N_1360,N_11,N_997);
or U1361 (N_1361,N_772,In_1633);
and U1362 (N_1362,In_1650,N_794);
or U1363 (N_1363,In_1773,N_970);
nor U1364 (N_1364,N_760,In_10);
xnor U1365 (N_1365,N_998,N_902);
or U1366 (N_1366,N_385,N_78);
nand U1367 (N_1367,N_816,In_913);
nor U1368 (N_1368,N_28,In_693);
nand U1369 (N_1369,N_656,N_791);
nand U1370 (N_1370,N_841,In_173);
nor U1371 (N_1371,In_479,In_2354);
xnor U1372 (N_1372,In_411,N_554);
or U1373 (N_1373,N_801,N_384);
xor U1374 (N_1374,N_950,N_745);
xnor U1375 (N_1375,N_890,In_1822);
nor U1376 (N_1376,N_927,N_485);
or U1377 (N_1377,N_704,In_159);
xnor U1378 (N_1378,N_42,N_348);
nor U1379 (N_1379,N_459,In_2171);
or U1380 (N_1380,N_748,N_728);
nand U1381 (N_1381,N_497,N_318);
nand U1382 (N_1382,N_443,N_551);
and U1383 (N_1383,N_145,N_689);
and U1384 (N_1384,N_749,N_831);
nor U1385 (N_1385,N_364,N_38);
xor U1386 (N_1386,In_1488,N_186);
and U1387 (N_1387,N_931,N_16);
xnor U1388 (N_1388,N_237,In_86);
and U1389 (N_1389,In_283,In_606);
and U1390 (N_1390,In_233,In_264);
xnor U1391 (N_1391,N_637,N_19);
nor U1392 (N_1392,In_1244,N_327);
or U1393 (N_1393,N_115,N_230);
nand U1394 (N_1394,N_951,N_172);
and U1395 (N_1395,In_1865,In_1299);
and U1396 (N_1396,N_330,N_908);
nor U1397 (N_1397,In_1002,In_540);
nand U1398 (N_1398,In_744,N_440);
nand U1399 (N_1399,N_877,In_185);
nor U1400 (N_1400,N_242,N_209);
nand U1401 (N_1401,N_548,N_134);
or U1402 (N_1402,In_2209,N_105);
or U1403 (N_1403,In_557,In_38);
and U1404 (N_1404,N_675,In_1620);
xor U1405 (N_1405,N_669,N_608);
and U1406 (N_1406,N_690,N_987);
nand U1407 (N_1407,In_1368,N_856);
and U1408 (N_1408,In_849,N_834);
or U1409 (N_1409,N_247,N_411);
nand U1410 (N_1410,In_1741,N_24);
nor U1411 (N_1411,In_1594,In_760);
and U1412 (N_1412,N_448,N_446);
nor U1413 (N_1413,N_295,In_1921);
and U1414 (N_1414,N_625,In_2082);
nand U1415 (N_1415,N_409,In_1571);
or U1416 (N_1416,N_339,N_340);
nand U1417 (N_1417,N_563,In_459);
nor U1418 (N_1418,N_213,N_959);
nor U1419 (N_1419,N_400,N_899);
or U1420 (N_1420,N_136,In_1954);
nor U1421 (N_1421,N_572,In_2235);
nand U1422 (N_1422,In_426,In_1645);
nor U1423 (N_1423,In_663,N_185);
and U1424 (N_1424,N_584,N_747);
and U1425 (N_1425,N_4,In_6);
xnor U1426 (N_1426,In_1149,N_674);
xor U1427 (N_1427,N_505,N_313);
and U1428 (N_1428,N_955,N_253);
nor U1429 (N_1429,N_467,N_174);
nand U1430 (N_1430,N_784,N_521);
and U1431 (N_1431,N_127,In_848);
or U1432 (N_1432,In_2071,In_938);
and U1433 (N_1433,N_593,N_619);
and U1434 (N_1434,N_708,N_429);
and U1435 (N_1435,N_928,N_740);
nor U1436 (N_1436,In_2134,N_628);
or U1437 (N_1437,N_614,N_388);
or U1438 (N_1438,N_553,N_404);
or U1439 (N_1439,In_2457,In_2213);
nor U1440 (N_1440,In_1677,In_1322);
nor U1441 (N_1441,In_1386,N_776);
xnor U1442 (N_1442,N_812,N_353);
nor U1443 (N_1443,N_989,N_797);
nor U1444 (N_1444,N_556,In_2052);
or U1445 (N_1445,N_308,N_591);
nor U1446 (N_1446,N_644,N_435);
nand U1447 (N_1447,N_451,N_276);
nor U1448 (N_1448,N_484,N_609);
or U1449 (N_1449,N_332,In_1637);
or U1450 (N_1450,N_933,N_48);
nand U1451 (N_1451,N_243,N_623);
nand U1452 (N_1452,In_616,N_486);
or U1453 (N_1453,In_235,N_314);
nand U1454 (N_1454,N_773,N_225);
and U1455 (N_1455,N_156,N_319);
xor U1456 (N_1456,N_464,In_346);
nor U1457 (N_1457,N_699,N_569);
nor U1458 (N_1458,In_943,In_1553);
and U1459 (N_1459,N_18,N_523);
xnor U1460 (N_1460,N_629,N_90);
xor U1461 (N_1461,In_1692,N_218);
or U1462 (N_1462,N_762,N_640);
and U1463 (N_1463,N_81,N_76);
or U1464 (N_1464,N_506,N_227);
xnor U1465 (N_1465,N_192,In_1475);
xor U1466 (N_1466,N_41,N_211);
and U1467 (N_1467,N_771,N_101);
and U1468 (N_1468,N_957,In_1591);
nand U1469 (N_1469,N_993,N_937);
or U1470 (N_1470,In_1787,N_825);
nor U1471 (N_1471,In_1638,N_250);
or U1472 (N_1472,N_394,In_706);
and U1473 (N_1473,N_873,N_696);
and U1474 (N_1474,N_139,N_396);
or U1475 (N_1475,N_821,In_1726);
nand U1476 (N_1476,N_598,N_552);
or U1477 (N_1477,N_785,In_54);
or U1478 (N_1478,N_589,In_954);
nor U1479 (N_1479,N_471,N_720);
nand U1480 (N_1480,N_147,In_116);
and U1481 (N_1481,N_641,N_539);
and U1482 (N_1482,In_1877,In_1202);
nand U1483 (N_1483,N_111,In_260);
and U1484 (N_1484,N_271,In_1407);
xnor U1485 (N_1485,In_251,In_2066);
nand U1486 (N_1486,N_198,In_484);
and U1487 (N_1487,N_532,N_882);
and U1488 (N_1488,N_513,N_713);
or U1489 (N_1489,N_738,N_568);
and U1490 (N_1490,N_423,N_555);
and U1491 (N_1491,In_1499,N_129);
or U1492 (N_1492,In_344,In_1560);
nor U1493 (N_1493,N_155,N_736);
nor U1494 (N_1494,N_316,In_880);
or U1495 (N_1495,N_132,N_422);
nor U1496 (N_1496,In_1116,N_621);
nor U1497 (N_1497,In_0,N_764);
xor U1498 (N_1498,In_1758,N_383);
and U1499 (N_1499,N_984,In_2358);
xnor U1500 (N_1500,In_1705,N_698);
or U1501 (N_1501,N_403,N_574);
and U1502 (N_1502,N_277,In_2028);
or U1503 (N_1503,N_894,N_263);
nand U1504 (N_1504,In_928,In_2174);
xor U1505 (N_1505,N_944,N_807);
nand U1506 (N_1506,N_980,In_163);
or U1507 (N_1507,N_378,N_705);
xnor U1508 (N_1508,N_34,N_306);
nand U1509 (N_1509,In_2411,N_387);
or U1510 (N_1510,N_583,In_282);
xnor U1511 (N_1511,N_660,N_565);
or U1512 (N_1512,N_317,N_994);
and U1513 (N_1513,N_304,N_500);
or U1514 (N_1514,N_61,N_479);
nand U1515 (N_1515,In_1227,N_442);
and U1516 (N_1516,N_366,N_54);
or U1517 (N_1517,In_2468,N_412);
nor U1518 (N_1518,In_514,N_793);
or U1519 (N_1519,N_17,N_848);
nor U1520 (N_1520,In_1851,In_746);
nor U1521 (N_1521,In_139,In_586);
nand U1522 (N_1522,In_1256,N_520);
and U1523 (N_1523,N_977,In_2434);
or U1524 (N_1524,N_36,In_862);
and U1525 (N_1525,N_323,N_477);
and U1526 (N_1526,N_871,N_104);
or U1527 (N_1527,In_370,N_149);
nand U1528 (N_1528,In_472,In_2484);
nand U1529 (N_1529,In_244,In_1810);
xnor U1530 (N_1530,N_498,In_2029);
and U1531 (N_1531,N_655,N_405);
nand U1532 (N_1532,N_77,N_792);
xnor U1533 (N_1533,In_2309,N_217);
and U1534 (N_1534,In_542,N_702);
nand U1535 (N_1535,N_365,In_1046);
and U1536 (N_1536,N_586,In_401);
xor U1537 (N_1537,N_813,N_932);
nand U1538 (N_1538,N_986,N_143);
nand U1539 (N_1539,N_501,N_118);
nor U1540 (N_1540,N_444,In_304);
nor U1541 (N_1541,In_243,N_725);
or U1542 (N_1542,In_2405,In_2166);
nand U1543 (N_1543,N_664,N_153);
and U1544 (N_1544,In_545,N_880);
and U1545 (N_1545,N_6,In_1354);
xnor U1546 (N_1546,In_795,N_860);
or U1547 (N_1547,N_917,In_692);
or U1548 (N_1548,In_813,N_205);
nand U1549 (N_1549,N_259,N_490);
nor U1550 (N_1550,In_1616,N_659);
nor U1551 (N_1551,In_1103,N_37);
or U1552 (N_1552,In_323,In_2329);
and U1553 (N_1553,In_2193,In_657);
and U1554 (N_1554,N_178,N_510);
and U1555 (N_1555,N_907,N_742);
nor U1556 (N_1556,N_390,N_646);
nand U1557 (N_1557,N_1,N_197);
xor U1558 (N_1558,N_261,In_1259);
and U1559 (N_1559,N_929,N_84);
nand U1560 (N_1560,N_288,N_315);
xnor U1561 (N_1561,N_123,N_836);
or U1562 (N_1562,N_694,N_331);
and U1563 (N_1563,N_898,N_590);
xor U1564 (N_1564,In_832,N_281);
nand U1565 (N_1565,N_73,N_886);
xnor U1566 (N_1566,N_921,N_296);
xnor U1567 (N_1567,N_869,N_909);
nand U1568 (N_1568,N_560,N_201);
and U1569 (N_1569,N_954,N_693);
and U1570 (N_1570,N_893,N_549);
xor U1571 (N_1571,In_1436,N_8);
nor U1572 (N_1572,N_517,N_700);
or U1573 (N_1573,N_910,N_853);
nor U1574 (N_1574,N_312,In_2031);
xnor U1575 (N_1575,N_389,N_474);
nand U1576 (N_1576,In_2030,In_1911);
or U1577 (N_1577,N_684,N_519);
or U1578 (N_1578,N_56,N_265);
and U1579 (N_1579,In_2250,N_347);
xor U1580 (N_1580,N_95,N_550);
xnor U1581 (N_1581,In_2127,N_948);
nor U1582 (N_1582,In_171,In_1967);
nand U1583 (N_1583,In_142,N_862);
xor U1584 (N_1584,N_524,N_673);
nand U1585 (N_1585,N_71,N_94);
and U1586 (N_1586,N_204,N_868);
nand U1587 (N_1587,N_849,N_567);
and U1588 (N_1588,N_561,N_846);
nor U1589 (N_1589,In_1114,N_425);
xnor U1590 (N_1590,In_14,N_44);
or U1591 (N_1591,N_309,N_150);
nand U1592 (N_1592,In_1813,In_1626);
xor U1593 (N_1593,N_665,N_558);
or U1594 (N_1594,N_461,N_805);
nand U1595 (N_1595,N_303,In_2048);
nand U1596 (N_1596,In_1434,In_402);
nor U1597 (N_1597,N_66,In_1471);
xnor U1598 (N_1598,In_1912,N_573);
nor U1599 (N_1599,N_939,In_1105);
nand U1600 (N_1600,N_307,In_2265);
nor U1601 (N_1601,In_2322,N_159);
nor U1602 (N_1602,N_919,In_2385);
and U1603 (N_1603,N_822,N_441);
or U1604 (N_1604,N_310,In_1221);
and U1605 (N_1605,N_788,N_456);
and U1606 (N_1606,N_74,N_709);
nand U1607 (N_1607,N_766,N_717);
nor U1608 (N_1608,N_40,N_336);
or U1609 (N_1609,In_1419,N_783);
nor U1610 (N_1610,In_887,N_936);
xnor U1611 (N_1611,N_775,N_711);
xor U1612 (N_1612,In_1293,N_392);
or U1613 (N_1613,N_439,N_202);
and U1614 (N_1614,N_357,N_86);
nand U1615 (N_1615,N_289,In_2345);
nand U1616 (N_1616,N_436,In_1157);
and U1617 (N_1617,N_544,N_870);
or U1618 (N_1618,N_545,N_557);
xor U1619 (N_1619,N_796,N_511);
or U1620 (N_1620,N_683,N_262);
nor U1621 (N_1621,In_467,In_2214);
and U1622 (N_1622,N_450,In_944);
nor U1623 (N_1623,In_1276,N_579);
or U1624 (N_1624,N_275,N_537);
nor U1625 (N_1625,N_695,In_1318);
or U1626 (N_1626,N_802,N_344);
nor U1627 (N_1627,N_988,In_830);
and U1628 (N_1628,In_2215,In_611);
or U1629 (N_1629,In_2351,In_705);
nand U1630 (N_1630,In_885,N_744);
nor U1631 (N_1631,N_358,N_829);
or U1632 (N_1632,N_631,In_2114);
nor U1633 (N_1633,N_128,N_63);
nand U1634 (N_1634,In_475,In_301);
nand U1635 (N_1635,In_2424,N_395);
nor U1636 (N_1636,N_643,N_516);
or U1637 (N_1637,In_2499,In_190);
or U1638 (N_1638,N_368,N_727);
or U1639 (N_1639,N_354,In_2452);
xor U1640 (N_1640,N_369,In_1018);
nor U1641 (N_1641,N_903,N_778);
nand U1642 (N_1642,N_377,In_1066);
or U1643 (N_1643,N_810,N_469);
nand U1644 (N_1644,N_463,N_576);
or U1645 (N_1645,N_782,In_975);
or U1646 (N_1646,N_137,N_215);
and U1647 (N_1647,In_2208,N_602);
xnor U1648 (N_1648,N_171,N_58);
and U1649 (N_1649,N_587,In_745);
nor U1650 (N_1650,In_2437,N_722);
xor U1651 (N_1651,N_488,In_615);
nor U1652 (N_1652,N_59,N_294);
xor U1653 (N_1653,N_245,In_180);
or U1654 (N_1654,N_462,N_774);
nand U1655 (N_1655,In_1687,In_281);
and U1656 (N_1656,In_2236,N_638);
or U1657 (N_1657,N_777,N_896);
or U1658 (N_1658,N_72,In_2182);
xor U1659 (N_1659,N_935,In_1842);
and U1660 (N_1660,In_773,In_250);
xor U1661 (N_1661,N_260,N_80);
nand U1662 (N_1662,In_1603,N_645);
nor U1663 (N_1663,In_1566,In_1922);
or U1664 (N_1664,In_1604,In_73);
nand U1665 (N_1665,N_39,In_1505);
and U1666 (N_1666,In_1124,N_666);
nand U1667 (N_1667,In_1260,N_884);
nor U1668 (N_1668,In_1056,N_418);
nor U1669 (N_1669,N_996,N_718);
nand U1670 (N_1670,N_151,N_739);
and U1671 (N_1671,In_2324,In_767);
nand U1672 (N_1672,In_1206,In_31);
xor U1673 (N_1673,N_753,N_734);
and U1674 (N_1674,N_904,In_1772);
or U1675 (N_1675,N_302,N_595);
or U1676 (N_1676,N_473,N_983);
xor U1677 (N_1677,N_431,In_856);
xnor U1678 (N_1678,In_2243,In_1802);
xor U1679 (N_1679,N_82,N_850);
xor U1680 (N_1680,In_787,In_1618);
and U1681 (N_1681,N_585,In_1254);
nand U1682 (N_1682,N_207,In_269);
and U1683 (N_1683,N_757,In_596);
and U1684 (N_1684,In_1335,N_334);
and U1685 (N_1685,In_1756,N_324);
xnor U1686 (N_1686,N_214,In_948);
nor U1687 (N_1687,In_1441,N_458);
nand U1688 (N_1688,N_68,In_129);
or U1689 (N_1689,In_228,N_889);
and U1690 (N_1690,N_833,In_1530);
or U1691 (N_1691,N_398,N_842);
and U1692 (N_1692,N_495,In_489);
and U1693 (N_1693,N_758,N_808);
xnor U1694 (N_1694,N_864,N_973);
nand U1695 (N_1695,N_362,In_470);
and U1696 (N_1696,N_964,In_622);
or U1697 (N_1697,N_891,N_87);
and U1698 (N_1698,In_2334,N_31);
nor U1699 (N_1699,In_1193,N_715);
nor U1700 (N_1700,N_413,N_279);
xor U1701 (N_1701,In_1666,In_852);
or U1702 (N_1702,N_196,N_952);
or U1703 (N_1703,N_452,N_287);
and U1704 (N_1704,In_172,In_2244);
or U1705 (N_1705,N_508,N_653);
nor U1706 (N_1706,N_190,In_1088);
nor U1707 (N_1707,N_154,In_779);
xnor U1708 (N_1708,N_543,N_863);
nand U1709 (N_1709,N_661,N_843);
or U1710 (N_1710,In_75,N_594);
nor U1711 (N_1711,In_377,N_15);
and U1712 (N_1712,N_721,In_1336);
nand U1713 (N_1713,N_397,N_300);
or U1714 (N_1714,N_992,N_786);
nor U1715 (N_1715,N_710,In_2036);
nand U1716 (N_1716,N_493,N_371);
nand U1717 (N_1717,N_483,In_1971);
or U1718 (N_1718,N_530,N_13);
and U1719 (N_1719,In_267,N_639);
xor U1720 (N_1720,N_938,N_466);
and U1721 (N_1721,N_960,N_428);
xnor U1722 (N_1722,In_2281,In_2428);
or U1723 (N_1723,N_852,In_2377);
xor U1724 (N_1724,N_222,In_1423);
nand U1725 (N_1725,N_540,N_226);
nand U1726 (N_1726,N_346,N_103);
nor U1727 (N_1727,N_875,N_292);
xor U1728 (N_1728,N_687,In_1170);
nor U1729 (N_1729,N_480,In_702);
nor U1730 (N_1730,N_119,In_132);
xnor U1731 (N_1731,In_1999,In_1166);
xor U1732 (N_1732,N_320,N_133);
nor U1733 (N_1733,In_347,N_600);
or U1734 (N_1734,N_509,N_376);
xor U1735 (N_1735,In_121,N_817);
and U1736 (N_1736,N_195,In_715);
and U1737 (N_1737,N_814,In_1064);
and U1738 (N_1738,In_2426,N_43);
nand U1739 (N_1739,In_2459,In_505);
nand U1740 (N_1740,In_1649,N_210);
nand U1741 (N_1741,N_249,In_1918);
nor U1742 (N_1742,In_167,N_55);
nand U1743 (N_1743,In_221,In_580);
or U1744 (N_1744,N_914,N_982);
xnor U1745 (N_1745,In_319,N_199);
and U1746 (N_1746,In_2409,N_976);
nand U1747 (N_1747,In_822,N_632);
and U1748 (N_1748,N_363,In_1673);
nand U1749 (N_1749,N_649,N_113);
and U1750 (N_1750,In_1522,In_1056);
nor U1751 (N_1751,In_2481,N_449);
xnor U1752 (N_1752,N_593,N_376);
or U1753 (N_1753,N_609,N_829);
nor U1754 (N_1754,N_95,In_1851);
or U1755 (N_1755,N_103,In_1441);
nor U1756 (N_1756,In_1087,N_102);
and U1757 (N_1757,N_870,N_837);
nand U1758 (N_1758,N_718,In_1326);
xnor U1759 (N_1759,In_401,N_583);
and U1760 (N_1760,In_370,In_1638);
and U1761 (N_1761,N_937,N_212);
nor U1762 (N_1762,N_189,In_2040);
and U1763 (N_1763,N_214,In_2448);
nor U1764 (N_1764,N_448,N_403);
nor U1765 (N_1765,In_946,N_184);
nor U1766 (N_1766,In_1259,N_756);
xor U1767 (N_1767,N_957,N_317);
or U1768 (N_1768,N_891,N_460);
or U1769 (N_1769,In_380,In_867);
or U1770 (N_1770,N_801,N_144);
nand U1771 (N_1771,N_95,N_15);
nor U1772 (N_1772,N_148,In_14);
or U1773 (N_1773,N_571,N_97);
or U1774 (N_1774,N_631,N_350);
nand U1775 (N_1775,N_492,N_255);
nor U1776 (N_1776,In_1103,In_192);
nand U1777 (N_1777,In_401,N_83);
or U1778 (N_1778,N_868,N_105);
nand U1779 (N_1779,N_440,N_473);
nor U1780 (N_1780,In_1101,In_2071);
nand U1781 (N_1781,N_319,N_420);
nor U1782 (N_1782,N_13,In_2085);
xor U1783 (N_1783,N_36,N_377);
and U1784 (N_1784,N_536,In_599);
or U1785 (N_1785,N_833,N_395);
nor U1786 (N_1786,In_267,N_23);
nand U1787 (N_1787,N_381,N_339);
xnor U1788 (N_1788,N_166,In_1221);
and U1789 (N_1789,N_205,N_373);
or U1790 (N_1790,N_74,In_2028);
xnor U1791 (N_1791,In_1549,N_404);
and U1792 (N_1792,N_36,N_811);
or U1793 (N_1793,N_992,N_411);
nor U1794 (N_1794,N_425,N_915);
nor U1795 (N_1795,N_356,N_39);
nor U1796 (N_1796,N_830,In_1522);
and U1797 (N_1797,N_482,In_116);
or U1798 (N_1798,N_804,N_48);
or U1799 (N_1799,In_1880,N_47);
nand U1800 (N_1800,N_684,N_936);
nand U1801 (N_1801,N_808,N_283);
or U1802 (N_1802,N_918,N_736);
nand U1803 (N_1803,N_856,In_557);
and U1804 (N_1804,In_2354,N_823);
xor U1805 (N_1805,N_774,N_144);
xor U1806 (N_1806,N_285,N_83);
xnor U1807 (N_1807,In_1530,N_106);
nor U1808 (N_1808,In_1865,N_445);
xor U1809 (N_1809,In_1124,In_1244);
xnor U1810 (N_1810,N_102,N_651);
nand U1811 (N_1811,N_291,N_77);
nor U1812 (N_1812,N_743,In_2193);
nor U1813 (N_1813,N_719,N_739);
nand U1814 (N_1814,N_355,In_739);
nor U1815 (N_1815,In_1988,N_598);
nand U1816 (N_1816,N_812,N_625);
nand U1817 (N_1817,N_447,In_1233);
nand U1818 (N_1818,N_844,N_412);
or U1819 (N_1819,In_264,N_725);
nand U1820 (N_1820,N_586,N_261);
or U1821 (N_1821,N_507,N_265);
nand U1822 (N_1822,In_2409,In_301);
xnor U1823 (N_1823,In_841,N_995);
xnor U1824 (N_1824,In_1859,N_146);
or U1825 (N_1825,N_501,N_83);
nor U1826 (N_1826,N_794,N_29);
and U1827 (N_1827,N_142,N_118);
or U1828 (N_1828,N_529,N_953);
and U1829 (N_1829,In_2082,In_2441);
or U1830 (N_1830,N_566,In_1821);
nand U1831 (N_1831,N_197,N_157);
or U1832 (N_1832,N_995,N_581);
nor U1833 (N_1833,In_1741,N_282);
or U1834 (N_1834,N_647,N_773);
xor U1835 (N_1835,N_561,N_507);
or U1836 (N_1836,N_850,In_1737);
nor U1837 (N_1837,N_502,N_28);
nor U1838 (N_1838,N_905,N_784);
xor U1839 (N_1839,N_703,N_943);
nor U1840 (N_1840,N_535,N_103);
xnor U1841 (N_1841,In_86,In_2351);
xor U1842 (N_1842,N_727,N_815);
or U1843 (N_1843,In_2127,In_385);
nor U1844 (N_1844,N_770,N_96);
xor U1845 (N_1845,N_836,In_1553);
or U1846 (N_1846,N_445,In_290);
nand U1847 (N_1847,N_141,N_851);
nor U1848 (N_1848,In_745,N_382);
xor U1849 (N_1849,N_354,N_818);
nor U1850 (N_1850,In_1149,N_307);
or U1851 (N_1851,N_936,N_961);
or U1852 (N_1852,In_1645,N_640);
and U1853 (N_1853,N_107,In_2437);
nor U1854 (N_1854,N_575,N_542);
nor U1855 (N_1855,N_863,N_426);
xor U1856 (N_1856,N_236,N_175);
or U1857 (N_1857,N_532,In_1530);
and U1858 (N_1858,N_107,N_591);
nand U1859 (N_1859,N_898,N_178);
or U1860 (N_1860,In_115,N_613);
or U1861 (N_1861,N_905,N_779);
and U1862 (N_1862,N_592,N_514);
and U1863 (N_1863,In_244,In_1264);
xor U1864 (N_1864,In_622,N_573);
nor U1865 (N_1865,N_709,N_177);
xnor U1866 (N_1866,N_670,N_785);
nor U1867 (N_1867,N_7,N_540);
and U1868 (N_1868,N_606,In_1434);
nand U1869 (N_1869,N_796,N_897);
xnor U1870 (N_1870,In_1725,N_524);
xnor U1871 (N_1871,N_413,N_190);
nand U1872 (N_1872,In_1213,N_832);
and U1873 (N_1873,In_2102,In_2134);
nor U1874 (N_1874,N_849,N_310);
nor U1875 (N_1875,In_2294,N_989);
or U1876 (N_1876,N_846,N_168);
nor U1877 (N_1877,In_983,In_2472);
nor U1878 (N_1878,N_393,N_290);
or U1879 (N_1879,In_228,In_2294);
nor U1880 (N_1880,In_1101,N_388);
nor U1881 (N_1881,N_534,In_1999);
xnor U1882 (N_1882,N_851,In_1692);
nand U1883 (N_1883,In_1604,In_2481);
nand U1884 (N_1884,N_446,N_684);
or U1885 (N_1885,N_349,N_707);
or U1886 (N_1886,In_1747,In_1136);
or U1887 (N_1887,In_415,N_192);
nand U1888 (N_1888,N_898,In_1116);
nor U1889 (N_1889,N_541,N_127);
or U1890 (N_1890,In_1224,N_925);
xnor U1891 (N_1891,In_1157,N_643);
nor U1892 (N_1892,N_357,N_432);
xor U1893 (N_1893,N_100,N_690);
xor U1894 (N_1894,N_155,N_904);
nand U1895 (N_1895,N_749,In_1419);
nor U1896 (N_1896,N_199,N_737);
and U1897 (N_1897,N_622,N_444);
xnor U1898 (N_1898,N_397,In_140);
nand U1899 (N_1899,N_137,N_853);
and U1900 (N_1900,N_340,N_537);
or U1901 (N_1901,In_2309,In_2052);
or U1902 (N_1902,N_533,In_2424);
or U1903 (N_1903,N_624,In_1103);
and U1904 (N_1904,N_218,N_314);
and U1905 (N_1905,N_644,In_1758);
nand U1906 (N_1906,N_55,N_820);
nand U1907 (N_1907,N_20,N_261);
nor U1908 (N_1908,N_881,N_7);
xnor U1909 (N_1909,N_406,N_273);
xnor U1910 (N_1910,N_866,N_217);
xor U1911 (N_1911,In_172,N_601);
and U1912 (N_1912,In_209,N_184);
and U1913 (N_1913,N_505,N_335);
nor U1914 (N_1914,N_852,In_1371);
or U1915 (N_1915,N_857,In_1475);
xnor U1916 (N_1916,N_286,In_693);
or U1917 (N_1917,N_885,In_1505);
nand U1918 (N_1918,In_753,In_828);
xnor U1919 (N_1919,N_695,N_981);
or U1920 (N_1920,In_1787,In_615);
xnor U1921 (N_1921,In_1305,N_774);
xor U1922 (N_1922,N_402,N_878);
nor U1923 (N_1923,N_243,In_580);
nand U1924 (N_1924,N_651,N_324);
or U1925 (N_1925,N_624,In_1371);
xnor U1926 (N_1926,N_8,N_453);
nor U1927 (N_1927,N_572,N_208);
xnor U1928 (N_1928,N_963,N_871);
nor U1929 (N_1929,N_75,In_2082);
or U1930 (N_1930,N_429,N_771);
and U1931 (N_1931,In_57,In_260);
nor U1932 (N_1932,N_576,N_902);
or U1933 (N_1933,N_688,N_861);
nand U1934 (N_1934,In_251,N_170);
or U1935 (N_1935,In_209,N_424);
xor U1936 (N_1936,N_100,N_505);
nor U1937 (N_1937,N_152,N_859);
or U1938 (N_1938,In_1322,N_394);
nand U1939 (N_1939,N_69,N_653);
nor U1940 (N_1940,In_190,N_577);
or U1941 (N_1941,N_186,N_586);
nor U1942 (N_1942,N_945,In_467);
nor U1943 (N_1943,N_890,N_134);
nor U1944 (N_1944,N_209,N_597);
xnor U1945 (N_1945,N_774,N_305);
and U1946 (N_1946,In_459,N_500);
xnor U1947 (N_1947,N_418,N_704);
nor U1948 (N_1948,N_291,In_1170);
xnor U1949 (N_1949,N_512,N_486);
nand U1950 (N_1950,N_554,N_459);
or U1951 (N_1951,N_118,N_641);
xor U1952 (N_1952,N_960,N_616);
or U1953 (N_1953,N_225,In_2075);
or U1954 (N_1954,In_101,N_398);
and U1955 (N_1955,In_712,N_429);
and U1956 (N_1956,N_467,N_264);
nand U1957 (N_1957,N_435,N_724);
nand U1958 (N_1958,N_487,N_690);
nand U1959 (N_1959,N_461,In_748);
or U1960 (N_1960,In_74,N_259);
and U1961 (N_1961,N_912,In_849);
or U1962 (N_1962,N_545,In_744);
or U1963 (N_1963,N_809,N_201);
nor U1964 (N_1964,In_1802,N_952);
and U1965 (N_1965,In_630,N_387);
or U1966 (N_1966,N_292,In_1064);
and U1967 (N_1967,N_931,N_142);
nor U1968 (N_1968,In_889,N_849);
nand U1969 (N_1969,In_377,N_443);
nor U1970 (N_1970,N_137,N_712);
nor U1971 (N_1971,N_414,N_426);
xor U1972 (N_1972,In_1773,N_536);
nor U1973 (N_1973,N_622,In_250);
and U1974 (N_1974,N_689,N_418);
xor U1975 (N_1975,N_323,N_720);
nor U1976 (N_1976,N_257,N_321);
or U1977 (N_1977,In_1502,N_519);
nand U1978 (N_1978,N_368,N_924);
and U1979 (N_1979,N_145,N_398);
xnor U1980 (N_1980,N_302,N_894);
or U1981 (N_1981,In_830,In_1737);
xnor U1982 (N_1982,In_1193,In_1375);
xnor U1983 (N_1983,N_513,In_773);
xnor U1984 (N_1984,N_558,N_446);
xor U1985 (N_1985,In_2447,N_67);
xor U1986 (N_1986,In_1821,N_754);
or U1987 (N_1987,In_1318,N_626);
nand U1988 (N_1988,N_75,N_156);
nand U1989 (N_1989,N_245,N_197);
nand U1990 (N_1990,N_527,N_482);
nor U1991 (N_1991,N_734,In_78);
xnor U1992 (N_1992,In_2147,N_417);
or U1993 (N_1993,N_2,N_796);
nor U1994 (N_1994,N_811,N_651);
nor U1995 (N_1995,N_402,In_1356);
xnor U1996 (N_1996,In_347,N_893);
xor U1997 (N_1997,N_133,N_22);
nand U1998 (N_1998,N_37,In_1030);
nand U1999 (N_1999,In_262,N_175);
nor U2000 (N_2000,N_1348,N_1697);
or U2001 (N_2001,N_1313,N_1492);
nor U2002 (N_2002,N_1165,N_1247);
nand U2003 (N_2003,N_1833,N_1890);
xor U2004 (N_2004,N_1608,N_1319);
nor U2005 (N_2005,N_1813,N_1748);
or U2006 (N_2006,N_1283,N_1181);
nor U2007 (N_2007,N_1870,N_1256);
nor U2008 (N_2008,N_1409,N_1618);
xor U2009 (N_2009,N_1801,N_1856);
and U2010 (N_2010,N_1630,N_1321);
or U2011 (N_2011,N_1255,N_1167);
xnor U2012 (N_2012,N_1043,N_1209);
nand U2013 (N_2013,N_1616,N_1170);
xor U2014 (N_2014,N_1772,N_1658);
xnor U2015 (N_2015,N_1547,N_1713);
nor U2016 (N_2016,N_1314,N_1597);
or U2017 (N_2017,N_1031,N_1602);
or U2018 (N_2018,N_1325,N_1470);
xor U2019 (N_2019,N_1228,N_1480);
nand U2020 (N_2020,N_1806,N_1795);
and U2021 (N_2021,N_1930,N_1961);
or U2022 (N_2022,N_1387,N_1947);
xnor U2023 (N_2023,N_1650,N_1768);
nor U2024 (N_2024,N_1148,N_1477);
nor U2025 (N_2025,N_1909,N_1566);
nand U2026 (N_2026,N_1593,N_1157);
or U2027 (N_2027,N_1021,N_1497);
nand U2028 (N_2028,N_1496,N_1192);
or U2029 (N_2029,N_1441,N_1107);
and U2030 (N_2030,N_1360,N_1932);
or U2031 (N_2031,N_1604,N_1421);
or U2032 (N_2032,N_1967,N_1464);
xor U2033 (N_2033,N_1797,N_1361);
or U2034 (N_2034,N_1123,N_1263);
and U2035 (N_2035,N_1504,N_1163);
and U2036 (N_2036,N_1219,N_1615);
nand U2037 (N_2037,N_1201,N_1337);
or U2038 (N_2038,N_1149,N_1814);
nand U2039 (N_2039,N_1137,N_1030);
and U2040 (N_2040,N_1840,N_1934);
or U2041 (N_2041,N_1037,N_1548);
or U2042 (N_2042,N_1972,N_1308);
nor U2043 (N_2043,N_1982,N_1029);
xor U2044 (N_2044,N_1689,N_1382);
and U2045 (N_2045,N_1385,N_1686);
or U2046 (N_2046,N_1681,N_1472);
nand U2047 (N_2047,N_1519,N_1394);
xnor U2048 (N_2048,N_1749,N_1558);
and U2049 (N_2049,N_1076,N_1637);
xnor U2050 (N_2050,N_1668,N_1834);
xnor U2051 (N_2051,N_1702,N_1927);
or U2052 (N_2052,N_1956,N_1483);
and U2053 (N_2053,N_1111,N_1493);
nor U2054 (N_2054,N_1996,N_1941);
and U2055 (N_2055,N_1708,N_1950);
xor U2056 (N_2056,N_1855,N_1775);
and U2057 (N_2057,N_1572,N_1272);
or U2058 (N_2058,N_1306,N_1859);
nor U2059 (N_2059,N_1286,N_1766);
nand U2060 (N_2060,N_1907,N_1282);
xor U2061 (N_2061,N_1380,N_1869);
nor U2062 (N_2062,N_1059,N_1067);
nor U2063 (N_2063,N_1931,N_1627);
and U2064 (N_2064,N_1260,N_1525);
nor U2065 (N_2065,N_1841,N_1114);
nor U2066 (N_2066,N_1543,N_1459);
and U2067 (N_2067,N_1638,N_1402);
nand U2068 (N_2068,N_1036,N_1747);
and U2069 (N_2069,N_1992,N_1551);
nand U2070 (N_2070,N_1077,N_1010);
nand U2071 (N_2071,N_1224,N_1046);
xnor U2072 (N_2072,N_1744,N_1629);
or U2073 (N_2073,N_1264,N_1753);
nand U2074 (N_2074,N_1861,N_1530);
nor U2075 (N_2075,N_1634,N_1968);
or U2076 (N_2076,N_1230,N_1805);
nor U2077 (N_2077,N_1478,N_1068);
xnor U2078 (N_2078,N_1151,N_1742);
nand U2079 (N_2079,N_1871,N_1590);
and U2080 (N_2080,N_1412,N_1916);
xor U2081 (N_2081,N_1475,N_1112);
nor U2082 (N_2082,N_1052,N_1993);
nand U2083 (N_2083,N_1202,N_1523);
or U2084 (N_2084,N_1568,N_1518);
xor U2085 (N_2085,N_1507,N_1463);
nor U2086 (N_2086,N_1177,N_1751);
xor U2087 (N_2087,N_1734,N_1442);
or U2088 (N_2088,N_1220,N_1549);
nand U2089 (N_2089,N_1688,N_1559);
or U2090 (N_2090,N_1635,N_1746);
nor U2091 (N_2091,N_1487,N_1132);
nand U2092 (N_2092,N_1414,N_1513);
nand U2093 (N_2093,N_1115,N_1088);
and U2094 (N_2094,N_1745,N_1245);
xnor U2095 (N_2095,N_1860,N_1583);
or U2096 (N_2096,N_1910,N_1207);
nor U2097 (N_2097,N_1914,N_1295);
nand U2098 (N_2098,N_1574,N_1644);
and U2099 (N_2099,N_1539,N_1456);
nor U2100 (N_2100,N_1677,N_1083);
nand U2101 (N_2101,N_1505,N_1328);
nand U2102 (N_2102,N_1905,N_1375);
or U2103 (N_2103,N_1595,N_1884);
and U2104 (N_2104,N_1320,N_1318);
xor U2105 (N_2105,N_1189,N_1705);
nor U2106 (N_2106,N_1527,N_1218);
xor U2107 (N_2107,N_1099,N_1130);
and U2108 (N_2108,N_1128,N_1235);
nand U2109 (N_2109,N_1449,N_1390);
and U2110 (N_2110,N_1039,N_1854);
nand U2111 (N_2111,N_1988,N_1820);
nor U2112 (N_2112,N_1617,N_1999);
xnor U2113 (N_2113,N_1471,N_1926);
nor U2114 (N_2114,N_1490,N_1079);
xnor U2115 (N_2115,N_1995,N_1004);
nand U2116 (N_2116,N_1345,N_1420);
xor U2117 (N_2117,N_1034,N_1138);
nand U2118 (N_2118,N_1266,N_1237);
nor U2119 (N_2119,N_1935,N_1919);
xnor U2120 (N_2120,N_1399,N_1655);
nand U2121 (N_2121,N_1675,N_1397);
or U2122 (N_2122,N_1529,N_1821);
nand U2123 (N_2123,N_1178,N_1000);
and U2124 (N_2124,N_1270,N_1729);
xor U2125 (N_2125,N_1550,N_1054);
xnor U2126 (N_2126,N_1569,N_1761);
nor U2127 (N_2127,N_1511,N_1233);
nand U2128 (N_2128,N_1389,N_1489);
nor U2129 (N_2129,N_1769,N_1579);
and U2130 (N_2130,N_1001,N_1810);
nand U2131 (N_2131,N_1060,N_1093);
nand U2132 (N_2132,N_1271,N_1829);
xor U2133 (N_2133,N_1923,N_1843);
xnor U2134 (N_2134,N_1468,N_1791);
nand U2135 (N_2135,N_1508,N_1285);
nand U2136 (N_2136,N_1398,N_1051);
nand U2137 (N_2137,N_1169,N_1101);
nand U2138 (N_2138,N_1661,N_1610);
nand U2139 (N_2139,N_1249,N_1153);
and U2140 (N_2140,N_1994,N_1622);
xnor U2141 (N_2141,N_1837,N_1291);
nor U2142 (N_2142,N_1868,N_1809);
nand U2143 (N_2143,N_1591,N_1048);
and U2144 (N_2144,N_1279,N_1150);
and U2145 (N_2145,N_1817,N_1939);
nand U2146 (N_2146,N_1055,N_1918);
or U2147 (N_2147,N_1561,N_1469);
or U2148 (N_2148,N_1700,N_1857);
nor U2149 (N_2149,N_1824,N_1594);
nor U2150 (N_2150,N_1780,N_1373);
or U2151 (N_2151,N_1739,N_1023);
and U2152 (N_2152,N_1240,N_1364);
nor U2153 (N_2153,N_1792,N_1684);
xnor U2154 (N_2154,N_1844,N_1517);
nand U2155 (N_2155,N_1141,N_1011);
xnor U2156 (N_2156,N_1913,N_1071);
nor U2157 (N_2157,N_1646,N_1427);
xor U2158 (N_2158,N_1783,N_1050);
or U2159 (N_2159,N_1155,N_1546);
nor U2160 (N_2160,N_1522,N_1670);
nor U2161 (N_2161,N_1198,N_1903);
or U2162 (N_2162,N_1885,N_1624);
and U2163 (N_2163,N_1381,N_1014);
or U2164 (N_2164,N_1296,N_1243);
nand U2165 (N_2165,N_1006,N_1691);
nor U2166 (N_2166,N_1576,N_1987);
or U2167 (N_2167,N_1038,N_1556);
or U2168 (N_2168,N_1210,N_1288);
nor U2169 (N_2169,N_1632,N_1392);
or U2170 (N_2170,N_1304,N_1045);
xnor U2171 (N_2171,N_1898,N_1537);
or U2172 (N_2172,N_1952,N_1452);
or U2173 (N_2173,N_1351,N_1370);
nor U2174 (N_2174,N_1336,N_1356);
or U2175 (N_2175,N_1185,N_1359);
or U2176 (N_2176,N_1186,N_1600);
nand U2177 (N_2177,N_1440,N_1433);
nor U2178 (N_2178,N_1631,N_1231);
or U2179 (N_2179,N_1582,N_1921);
nand U2180 (N_2180,N_1589,N_1598);
xnor U2181 (N_2181,N_1180,N_1252);
xor U2182 (N_2182,N_1659,N_1728);
nand U2183 (N_2183,N_1925,N_1109);
nand U2184 (N_2184,N_1732,N_1984);
or U2185 (N_2185,N_1097,N_1825);
nor U2186 (N_2186,N_1940,N_1888);
nand U2187 (N_2187,N_1278,N_1486);
nor U2188 (N_2188,N_1152,N_1722);
and U2189 (N_2189,N_1378,N_1835);
nand U2190 (N_2190,N_1353,N_1665);
nand U2191 (N_2191,N_1120,N_1754);
nor U2192 (N_2192,N_1807,N_1404);
nand U2193 (N_2193,N_1300,N_1289);
nor U2194 (N_2194,N_1455,N_1401);
xor U2195 (N_2195,N_1958,N_1764);
xor U2196 (N_2196,N_1563,N_1042);
nor U2197 (N_2197,N_1415,N_1715);
nand U2198 (N_2198,N_1232,N_1485);
xnor U2199 (N_2199,N_1985,N_1727);
and U2200 (N_2200,N_1127,N_1267);
and U2201 (N_2201,N_1040,N_1838);
nor U2202 (N_2202,N_1265,N_1586);
or U2203 (N_2203,N_1396,N_1366);
xor U2204 (N_2204,N_1437,N_1113);
nor U2205 (N_2205,N_1474,N_1199);
or U2206 (N_2206,N_1896,N_1811);
nor U2207 (N_2207,N_1080,N_1828);
xnor U2208 (N_2208,N_1866,N_1020);
nor U2209 (N_2209,N_1154,N_1242);
or U2210 (N_2210,N_1332,N_1078);
nor U2211 (N_2211,N_1058,N_1438);
nor U2212 (N_2212,N_1534,N_1317);
nand U2213 (N_2213,N_1693,N_1822);
nand U2214 (N_2214,N_1592,N_1706);
nand U2215 (N_2215,N_1892,N_1405);
or U2216 (N_2216,N_1403,N_1425);
or U2217 (N_2217,N_1103,N_1831);
xnor U2218 (N_2218,N_1897,N_1462);
or U2219 (N_2219,N_1570,N_1092);
nor U2220 (N_2220,N_1718,N_1363);
or U2221 (N_2221,N_1799,N_1599);
or U2222 (N_2222,N_1662,N_1851);
nand U2223 (N_2223,N_1384,N_1253);
nand U2224 (N_2224,N_1977,N_1965);
xor U2225 (N_2225,N_1022,N_1719);
or U2226 (N_2226,N_1287,N_1945);
and U2227 (N_2227,N_1676,N_1625);
nor U2228 (N_2228,N_1976,N_1057);
xor U2229 (N_2229,N_1391,N_1696);
xnor U2230 (N_2230,N_1793,N_1491);
xor U2231 (N_2231,N_1917,N_1195);
nand U2232 (N_2232,N_1429,N_1274);
or U2233 (N_2233,N_1139,N_1110);
and U2234 (N_2234,N_1221,N_1090);
or U2235 (N_2235,N_1346,N_1347);
or U2236 (N_2236,N_1262,N_1002);
xnor U2237 (N_2237,N_1636,N_1555);
xor U2238 (N_2238,N_1545,N_1663);
xnor U2239 (N_2239,N_1881,N_1575);
and U2240 (N_2240,N_1488,N_1937);
or U2241 (N_2241,N_1408,N_1701);
and U2242 (N_2242,N_1763,N_1294);
xor U2243 (N_2243,N_1257,N_1657);
or U2244 (N_2244,N_1407,N_1639);
xor U2245 (N_2245,N_1400,N_1528);
nand U2246 (N_2246,N_1187,N_1275);
nand U2247 (N_2247,N_1091,N_1738);
nor U2248 (N_2248,N_1643,N_1121);
xor U2249 (N_2249,N_1538,N_1654);
or U2250 (N_2250,N_1454,N_1277);
or U2251 (N_2251,N_1803,N_1193);
or U2252 (N_2252,N_1516,N_1331);
xnor U2253 (N_2253,N_1571,N_1899);
or U2254 (N_2254,N_1105,N_1307);
nand U2255 (N_2255,N_1682,N_1889);
nor U2256 (N_2256,N_1443,N_1710);
nor U2257 (N_2257,N_1482,N_1808);
and U2258 (N_2258,N_1203,N_1015);
or U2259 (N_2259,N_1891,N_1862);
and U2260 (N_2260,N_1075,N_1258);
xnor U2261 (N_2261,N_1466,N_1816);
nor U2262 (N_2262,N_1369,N_1502);
nor U2263 (N_2263,N_1339,N_1760);
or U2264 (N_2264,N_1322,N_1943);
and U2265 (N_2265,N_1479,N_1554);
xor U2266 (N_2266,N_1096,N_1229);
and U2267 (N_2267,N_1188,N_1125);
or U2268 (N_2268,N_1311,N_1619);
nand U2269 (N_2269,N_1225,N_1197);
or U2270 (N_2270,N_1131,N_1327);
nand U2271 (N_2271,N_1933,N_1303);
xor U2272 (N_2272,N_1721,N_1104);
nor U2273 (N_2273,N_1750,N_1779);
nor U2274 (N_2274,N_1172,N_1316);
xor U2275 (N_2275,N_1371,N_1461);
and U2276 (N_2276,N_1334,N_1895);
or U2277 (N_2277,N_1874,N_1781);
and U2278 (N_2278,N_1166,N_1865);
and U2279 (N_2279,N_1964,N_1305);
nand U2280 (N_2280,N_1969,N_1158);
xnor U2281 (N_2281,N_1035,N_1259);
or U2282 (N_2282,N_1007,N_1515);
xnor U2283 (N_2283,N_1978,N_1827);
and U2284 (N_2284,N_1794,N_1126);
or U2285 (N_2285,N_1755,N_1330);
nor U2286 (N_2286,N_1413,N_1236);
and U2287 (N_2287,N_1847,N_1607);
xor U2288 (N_2288,N_1714,N_1611);
and U2289 (N_2289,N_1374,N_1499);
xnor U2290 (N_2290,N_1877,N_1435);
xnor U2291 (N_2291,N_1122,N_1009);
or U2292 (N_2292,N_1144,N_1293);
nand U2293 (N_2293,N_1342,N_1326);
or U2294 (N_2294,N_1019,N_1609);
or U2295 (N_2295,N_1119,N_1560);
and U2296 (N_2296,N_1161,N_1074);
or U2297 (N_2297,N_1072,N_1695);
xor U2298 (N_2298,N_1648,N_1213);
xnor U2299 (N_2299,N_1395,N_1906);
nand U2300 (N_2300,N_1116,N_1842);
nand U2301 (N_2301,N_1542,N_1687);
nor U2302 (N_2302,N_1852,N_1182);
xnor U2303 (N_2303,N_1142,N_1882);
or U2304 (N_2304,N_1447,N_1674);
or U2305 (N_2305,N_1312,N_1983);
and U2306 (N_2306,N_1873,N_1786);
and U2307 (N_2307,N_1357,N_1770);
xor U2308 (N_2308,N_1268,N_1500);
xnor U2309 (N_2309,N_1887,N_1944);
xnor U2310 (N_2310,N_1717,N_1893);
nor U2311 (N_2311,N_1016,N_1422);
or U2312 (N_2312,N_1510,N_1184);
nand U2313 (N_2313,N_1535,N_1241);
and U2314 (N_2314,N_1222,N_1901);
and U2315 (N_2315,N_1883,N_1234);
and U2316 (N_2316,N_1778,N_1973);
nor U2317 (N_2317,N_1372,N_1915);
or U2318 (N_2318,N_1056,N_1553);
or U2319 (N_2319,N_1849,N_1061);
nand U2320 (N_2320,N_1953,N_1424);
and U2321 (N_2321,N_1005,N_1206);
nand U2322 (N_2322,N_1026,N_1073);
nor U2323 (N_2323,N_1215,N_1876);
and U2324 (N_2324,N_1106,N_1419);
nand U2325 (N_2325,N_1666,N_1208);
nor U2326 (N_2326,N_1341,N_1790);
xnor U2327 (N_2327,N_1416,N_1614);
or U2328 (N_2328,N_1875,N_1911);
and U2329 (N_2329,N_1752,N_1736);
and U2330 (N_2330,N_1960,N_1924);
nor U2331 (N_2331,N_1564,N_1724);
nand U2332 (N_2332,N_1044,N_1532);
nand U2333 (N_2333,N_1920,N_1164);
or U2334 (N_2334,N_1217,N_1143);
xnor U2335 (N_2335,N_1990,N_1227);
nor U2336 (N_2336,N_1212,N_1853);
nor U2337 (N_2337,N_1756,N_1818);
and U2338 (N_2338,N_1606,N_1678);
nand U2339 (N_2339,N_1509,N_1740);
nand U2340 (N_2340,N_1084,N_1848);
and U2341 (N_2341,N_1033,N_1928);
or U2342 (N_2342,N_1388,N_1640);
or U2343 (N_2343,N_1584,N_1226);
or U2344 (N_2344,N_1309,N_1191);
nor U2345 (N_2345,N_1991,N_1418);
nor U2346 (N_2346,N_1070,N_1018);
xnor U2347 (N_2347,N_1254,N_1129);
xnor U2348 (N_2348,N_1660,N_1467);
and U2349 (N_2349,N_1411,N_1823);
or U2350 (N_2350,N_1417,N_1613);
and U2351 (N_2351,N_1900,N_1368);
and U2352 (N_2352,N_1726,N_1102);
xnor U2353 (N_2353,N_1481,N_1878);
or U2354 (N_2354,N_1577,N_1520);
nand U2355 (N_2355,N_1290,N_1703);
and U2356 (N_2356,N_1066,N_1017);
or U2357 (N_2357,N_1273,N_1297);
or U2358 (N_2358,N_1365,N_1782);
nand U2359 (N_2359,N_1281,N_1867);
and U2360 (N_2360,N_1216,N_1773);
xor U2361 (N_2361,N_1176,N_1064);
nor U2362 (N_2362,N_1621,N_1501);
or U2363 (N_2363,N_1626,N_1671);
or U2364 (N_2364,N_1200,N_1839);
nand U2365 (N_2365,N_1248,N_1503);
and U2366 (N_2366,N_1211,N_1980);
nand U2367 (N_2367,N_1159,N_1439);
nand U2368 (N_2368,N_1386,N_1628);
and U2369 (N_2369,N_1767,N_1098);
nand U2370 (N_2370,N_1776,N_1473);
nand U2371 (N_2371,N_1434,N_1494);
and U2372 (N_2372,N_1680,N_1694);
or U2373 (N_2373,N_1759,N_1377);
or U2374 (N_2374,N_1450,N_1730);
nand U2375 (N_2375,N_1383,N_1725);
xor U2376 (N_2376,N_1698,N_1445);
or U2377 (N_2377,N_1565,N_1205);
nor U2378 (N_2378,N_1938,N_1707);
and U2379 (N_2379,N_1690,N_1785);
and U2380 (N_2380,N_1065,N_1041);
and U2381 (N_2381,N_1376,N_1812);
and U2382 (N_2382,N_1647,N_1024);
or U2383 (N_2383,N_1832,N_1942);
nor U2384 (N_2384,N_1118,N_1951);
and U2385 (N_2385,N_1175,N_1393);
or U2386 (N_2386,N_1298,N_1966);
and U2387 (N_2387,N_1085,N_1758);
nand U2388 (N_2388,N_1174,N_1652);
xnor U2389 (N_2389,N_1135,N_1013);
nand U2390 (N_2390,N_1850,N_1735);
xnor U2391 (N_2391,N_1214,N_1536);
nand U2392 (N_2392,N_1133,N_1787);
or U2393 (N_2393,N_1190,N_1557);
or U2394 (N_2394,N_1804,N_1436);
or U2395 (N_2395,N_1012,N_1183);
or U2396 (N_2396,N_1989,N_1959);
and U2397 (N_2397,N_1292,N_1086);
xor U2398 (N_2398,N_1246,N_1406);
xor U2399 (N_2399,N_1284,N_1970);
or U2400 (N_2400,N_1335,N_1664);
nand U2401 (N_2401,N_1446,N_1929);
and U2402 (N_2402,N_1460,N_1651);
or U2403 (N_2403,N_1062,N_1239);
xor U2404 (N_2404,N_1476,N_1338);
and U2405 (N_2405,N_1997,N_1845);
and U2406 (N_2406,N_1465,N_1100);
or U2407 (N_2407,N_1904,N_1025);
nor U2408 (N_2408,N_1008,N_1147);
or U2409 (N_2409,N_1349,N_1484);
or U2410 (N_2410,N_1301,N_1367);
nand U2411 (N_2411,N_1082,N_1692);
or U2412 (N_2412,N_1063,N_1633);
nor U2413 (N_2413,N_1521,N_1712);
and U2414 (N_2414,N_1581,N_1936);
xor U2415 (N_2415,N_1514,N_1423);
nor U2416 (N_2416,N_1975,N_1134);
nor U2417 (N_2417,N_1863,N_1354);
nor U2418 (N_2418,N_1498,N_1587);
and U2419 (N_2419,N_1605,N_1315);
nor U2420 (N_2420,N_1324,N_1789);
nand U2421 (N_2421,N_1981,N_1788);
xor U2422 (N_2422,N_1580,N_1667);
nor U2423 (N_2423,N_1765,N_1032);
nor U2424 (N_2424,N_1998,N_1524);
xnor U2425 (N_2425,N_1094,N_1800);
xor U2426 (N_2426,N_1986,N_1173);
or U2427 (N_2427,N_1495,N_1124);
nand U2428 (N_2428,N_1087,N_1344);
and U2429 (N_2429,N_1620,N_1578);
or U2430 (N_2430,N_1623,N_1458);
xnor U2431 (N_2431,N_1003,N_1596);
nand U2432 (N_2432,N_1815,N_1673);
and U2433 (N_2433,N_1448,N_1880);
nor U2434 (N_2434,N_1974,N_1720);
and U2435 (N_2435,N_1089,N_1140);
nor U2436 (N_2436,N_1963,N_1879);
nand U2437 (N_2437,N_1922,N_1612);
and U2438 (N_2438,N_1711,N_1771);
xor U2439 (N_2439,N_1340,N_1379);
and U2440 (N_2440,N_1774,N_1836);
or U2441 (N_2441,N_1709,N_1955);
or U2442 (N_2442,N_1117,N_1741);
and U2443 (N_2443,N_1430,N_1585);
nand U2444 (N_2444,N_1156,N_1194);
or U2445 (N_2445,N_1830,N_1047);
nor U2446 (N_2446,N_1957,N_1160);
and U2447 (N_2447,N_1355,N_1223);
or U2448 (N_2448,N_1081,N_1762);
xor U2449 (N_2449,N_1656,N_1872);
nor U2450 (N_2450,N_1802,N_1451);
or U2451 (N_2451,N_1567,N_1683);
xor U2452 (N_2452,N_1672,N_1444);
and U2453 (N_2453,N_1146,N_1276);
and U2454 (N_2454,N_1962,N_1541);
xnor U2455 (N_2455,N_1261,N_1601);
xnor U2456 (N_2456,N_1269,N_1136);
nand U2457 (N_2457,N_1588,N_1168);
nor U2458 (N_2458,N_1573,N_1552);
xor U2459 (N_2459,N_1027,N_1971);
and U2460 (N_2460,N_1053,N_1028);
nand U2461 (N_2461,N_1826,N_1310);
and U2462 (N_2462,N_1979,N_1908);
nor U2463 (N_2463,N_1352,N_1362);
or U2464 (N_2464,N_1244,N_1685);
and U2465 (N_2465,N_1894,N_1864);
nand U2466 (N_2466,N_1653,N_1743);
nor U2467 (N_2467,N_1251,N_1049);
nor U2468 (N_2468,N_1095,N_1846);
xnor U2469 (N_2469,N_1716,N_1358);
xnor U2470 (N_2470,N_1886,N_1679);
xor U2471 (N_2471,N_1302,N_1645);
and U2472 (N_2472,N_1333,N_1731);
nand U2473 (N_2473,N_1533,N_1453);
or U2474 (N_2474,N_1704,N_1145);
xnor U2475 (N_2475,N_1280,N_1343);
xnor U2476 (N_2476,N_1179,N_1162);
nand U2477 (N_2477,N_1642,N_1649);
nand U2478 (N_2478,N_1069,N_1948);
or U2479 (N_2479,N_1784,N_1540);
nand U2480 (N_2480,N_1108,N_1902);
or U2481 (N_2481,N_1949,N_1329);
nand U2482 (N_2482,N_1562,N_1723);
xor U2483 (N_2483,N_1798,N_1531);
nor U2484 (N_2484,N_1603,N_1431);
and U2485 (N_2485,N_1544,N_1250);
nand U2486 (N_2486,N_1699,N_1526);
and U2487 (N_2487,N_1669,N_1238);
nand U2488 (N_2488,N_1426,N_1777);
and U2489 (N_2489,N_1737,N_1428);
xnor U2490 (N_2490,N_1733,N_1506);
or U2491 (N_2491,N_1757,N_1299);
nand U2492 (N_2492,N_1432,N_1819);
nand U2493 (N_2493,N_1858,N_1946);
or U2494 (N_2494,N_1204,N_1171);
or U2495 (N_2495,N_1350,N_1641);
nor U2496 (N_2496,N_1954,N_1410);
or U2497 (N_2497,N_1796,N_1457);
nand U2498 (N_2498,N_1912,N_1196);
nor U2499 (N_2499,N_1323,N_1512);
nor U2500 (N_2500,N_1639,N_1373);
and U2501 (N_2501,N_1739,N_1294);
and U2502 (N_2502,N_1290,N_1569);
and U2503 (N_2503,N_1952,N_1548);
or U2504 (N_2504,N_1108,N_1596);
and U2505 (N_2505,N_1399,N_1188);
nand U2506 (N_2506,N_1130,N_1603);
and U2507 (N_2507,N_1107,N_1480);
xor U2508 (N_2508,N_1010,N_1799);
nand U2509 (N_2509,N_1342,N_1736);
and U2510 (N_2510,N_1775,N_1935);
nand U2511 (N_2511,N_1944,N_1160);
and U2512 (N_2512,N_1998,N_1681);
and U2513 (N_2513,N_1626,N_1001);
nand U2514 (N_2514,N_1247,N_1895);
and U2515 (N_2515,N_1892,N_1168);
xor U2516 (N_2516,N_1564,N_1006);
nand U2517 (N_2517,N_1329,N_1071);
xor U2518 (N_2518,N_1257,N_1158);
or U2519 (N_2519,N_1976,N_1326);
nand U2520 (N_2520,N_1597,N_1344);
xor U2521 (N_2521,N_1021,N_1616);
nor U2522 (N_2522,N_1246,N_1635);
nand U2523 (N_2523,N_1007,N_1739);
nor U2524 (N_2524,N_1161,N_1568);
and U2525 (N_2525,N_1784,N_1161);
xnor U2526 (N_2526,N_1149,N_1477);
nor U2527 (N_2527,N_1741,N_1660);
and U2528 (N_2528,N_1429,N_1854);
or U2529 (N_2529,N_1231,N_1611);
nand U2530 (N_2530,N_1017,N_1522);
xnor U2531 (N_2531,N_1255,N_1887);
xor U2532 (N_2532,N_1060,N_1774);
nand U2533 (N_2533,N_1430,N_1584);
or U2534 (N_2534,N_1864,N_1230);
nor U2535 (N_2535,N_1492,N_1403);
xor U2536 (N_2536,N_1260,N_1737);
nor U2537 (N_2537,N_1377,N_1038);
xnor U2538 (N_2538,N_1395,N_1348);
xor U2539 (N_2539,N_1966,N_1174);
nor U2540 (N_2540,N_1180,N_1542);
nor U2541 (N_2541,N_1355,N_1214);
nand U2542 (N_2542,N_1533,N_1103);
or U2543 (N_2543,N_1285,N_1627);
xor U2544 (N_2544,N_1495,N_1980);
and U2545 (N_2545,N_1420,N_1809);
nand U2546 (N_2546,N_1190,N_1267);
or U2547 (N_2547,N_1173,N_1336);
or U2548 (N_2548,N_1356,N_1343);
and U2549 (N_2549,N_1292,N_1335);
xnor U2550 (N_2550,N_1908,N_1447);
xnor U2551 (N_2551,N_1683,N_1800);
and U2552 (N_2552,N_1776,N_1366);
nand U2553 (N_2553,N_1859,N_1126);
or U2554 (N_2554,N_1459,N_1329);
or U2555 (N_2555,N_1261,N_1998);
xor U2556 (N_2556,N_1092,N_1844);
nand U2557 (N_2557,N_1317,N_1592);
xor U2558 (N_2558,N_1864,N_1527);
or U2559 (N_2559,N_1479,N_1728);
nand U2560 (N_2560,N_1125,N_1343);
or U2561 (N_2561,N_1770,N_1453);
or U2562 (N_2562,N_1170,N_1887);
or U2563 (N_2563,N_1157,N_1791);
nor U2564 (N_2564,N_1116,N_1266);
nand U2565 (N_2565,N_1651,N_1257);
nand U2566 (N_2566,N_1867,N_1815);
xor U2567 (N_2567,N_1782,N_1690);
xor U2568 (N_2568,N_1637,N_1306);
or U2569 (N_2569,N_1349,N_1523);
and U2570 (N_2570,N_1636,N_1853);
nand U2571 (N_2571,N_1758,N_1877);
and U2572 (N_2572,N_1731,N_1410);
nor U2573 (N_2573,N_1487,N_1423);
nor U2574 (N_2574,N_1203,N_1294);
nand U2575 (N_2575,N_1942,N_1330);
and U2576 (N_2576,N_1148,N_1949);
xor U2577 (N_2577,N_1953,N_1115);
and U2578 (N_2578,N_1992,N_1456);
and U2579 (N_2579,N_1376,N_1635);
nor U2580 (N_2580,N_1673,N_1170);
or U2581 (N_2581,N_1037,N_1705);
nand U2582 (N_2582,N_1350,N_1370);
xor U2583 (N_2583,N_1115,N_1888);
or U2584 (N_2584,N_1021,N_1774);
nor U2585 (N_2585,N_1368,N_1329);
or U2586 (N_2586,N_1841,N_1080);
nor U2587 (N_2587,N_1349,N_1827);
nor U2588 (N_2588,N_1396,N_1943);
or U2589 (N_2589,N_1135,N_1487);
nor U2590 (N_2590,N_1861,N_1318);
nand U2591 (N_2591,N_1471,N_1150);
nand U2592 (N_2592,N_1473,N_1325);
nor U2593 (N_2593,N_1016,N_1370);
and U2594 (N_2594,N_1992,N_1451);
and U2595 (N_2595,N_1373,N_1949);
nor U2596 (N_2596,N_1681,N_1671);
and U2597 (N_2597,N_1990,N_1257);
xnor U2598 (N_2598,N_1566,N_1605);
xor U2599 (N_2599,N_1457,N_1125);
xnor U2600 (N_2600,N_1005,N_1925);
nor U2601 (N_2601,N_1454,N_1333);
nand U2602 (N_2602,N_1558,N_1489);
nand U2603 (N_2603,N_1745,N_1012);
nand U2604 (N_2604,N_1446,N_1452);
or U2605 (N_2605,N_1649,N_1627);
nor U2606 (N_2606,N_1527,N_1548);
nand U2607 (N_2607,N_1031,N_1089);
and U2608 (N_2608,N_1019,N_1508);
nor U2609 (N_2609,N_1531,N_1380);
and U2610 (N_2610,N_1233,N_1540);
xnor U2611 (N_2611,N_1939,N_1371);
or U2612 (N_2612,N_1530,N_1951);
xor U2613 (N_2613,N_1679,N_1581);
nor U2614 (N_2614,N_1080,N_1168);
nor U2615 (N_2615,N_1431,N_1380);
nand U2616 (N_2616,N_1204,N_1822);
and U2617 (N_2617,N_1278,N_1347);
nor U2618 (N_2618,N_1461,N_1028);
or U2619 (N_2619,N_1556,N_1647);
xor U2620 (N_2620,N_1063,N_1112);
and U2621 (N_2621,N_1940,N_1659);
and U2622 (N_2622,N_1921,N_1104);
and U2623 (N_2623,N_1594,N_1642);
and U2624 (N_2624,N_1038,N_1638);
and U2625 (N_2625,N_1038,N_1628);
nand U2626 (N_2626,N_1446,N_1813);
xnor U2627 (N_2627,N_1859,N_1115);
nor U2628 (N_2628,N_1662,N_1078);
nor U2629 (N_2629,N_1047,N_1836);
nor U2630 (N_2630,N_1676,N_1269);
or U2631 (N_2631,N_1114,N_1296);
xor U2632 (N_2632,N_1957,N_1590);
nor U2633 (N_2633,N_1294,N_1066);
xor U2634 (N_2634,N_1432,N_1434);
nor U2635 (N_2635,N_1232,N_1631);
xor U2636 (N_2636,N_1740,N_1408);
nor U2637 (N_2637,N_1560,N_1081);
xor U2638 (N_2638,N_1475,N_1748);
nand U2639 (N_2639,N_1939,N_1411);
and U2640 (N_2640,N_1279,N_1494);
and U2641 (N_2641,N_1207,N_1952);
xor U2642 (N_2642,N_1561,N_1701);
nor U2643 (N_2643,N_1471,N_1710);
nor U2644 (N_2644,N_1102,N_1764);
nor U2645 (N_2645,N_1095,N_1477);
xnor U2646 (N_2646,N_1272,N_1191);
and U2647 (N_2647,N_1216,N_1676);
nand U2648 (N_2648,N_1401,N_1494);
nand U2649 (N_2649,N_1460,N_1859);
or U2650 (N_2650,N_1917,N_1208);
nand U2651 (N_2651,N_1024,N_1149);
nor U2652 (N_2652,N_1868,N_1507);
nand U2653 (N_2653,N_1208,N_1007);
nor U2654 (N_2654,N_1231,N_1911);
xnor U2655 (N_2655,N_1480,N_1148);
nor U2656 (N_2656,N_1442,N_1586);
nand U2657 (N_2657,N_1685,N_1696);
or U2658 (N_2658,N_1046,N_1854);
nor U2659 (N_2659,N_1864,N_1582);
or U2660 (N_2660,N_1424,N_1338);
nand U2661 (N_2661,N_1805,N_1331);
xnor U2662 (N_2662,N_1506,N_1503);
nand U2663 (N_2663,N_1042,N_1439);
nand U2664 (N_2664,N_1600,N_1281);
xor U2665 (N_2665,N_1494,N_1864);
nand U2666 (N_2666,N_1674,N_1854);
nor U2667 (N_2667,N_1697,N_1564);
xnor U2668 (N_2668,N_1709,N_1138);
or U2669 (N_2669,N_1673,N_1878);
nor U2670 (N_2670,N_1056,N_1557);
xnor U2671 (N_2671,N_1348,N_1350);
or U2672 (N_2672,N_1565,N_1443);
nand U2673 (N_2673,N_1845,N_1349);
and U2674 (N_2674,N_1857,N_1169);
xor U2675 (N_2675,N_1054,N_1807);
or U2676 (N_2676,N_1292,N_1043);
or U2677 (N_2677,N_1065,N_1739);
nand U2678 (N_2678,N_1146,N_1904);
xor U2679 (N_2679,N_1396,N_1928);
xnor U2680 (N_2680,N_1234,N_1868);
or U2681 (N_2681,N_1393,N_1292);
and U2682 (N_2682,N_1938,N_1953);
or U2683 (N_2683,N_1191,N_1231);
or U2684 (N_2684,N_1950,N_1136);
or U2685 (N_2685,N_1617,N_1216);
nor U2686 (N_2686,N_1259,N_1197);
or U2687 (N_2687,N_1981,N_1809);
nor U2688 (N_2688,N_1661,N_1472);
nand U2689 (N_2689,N_1221,N_1102);
and U2690 (N_2690,N_1507,N_1137);
xor U2691 (N_2691,N_1609,N_1772);
xor U2692 (N_2692,N_1553,N_1788);
or U2693 (N_2693,N_1492,N_1280);
nand U2694 (N_2694,N_1989,N_1028);
and U2695 (N_2695,N_1172,N_1117);
xor U2696 (N_2696,N_1439,N_1623);
or U2697 (N_2697,N_1544,N_1331);
xor U2698 (N_2698,N_1664,N_1398);
nand U2699 (N_2699,N_1245,N_1969);
or U2700 (N_2700,N_1225,N_1404);
or U2701 (N_2701,N_1635,N_1882);
nor U2702 (N_2702,N_1492,N_1206);
nand U2703 (N_2703,N_1695,N_1115);
nand U2704 (N_2704,N_1560,N_1287);
nor U2705 (N_2705,N_1487,N_1411);
and U2706 (N_2706,N_1560,N_1340);
nand U2707 (N_2707,N_1728,N_1513);
nor U2708 (N_2708,N_1582,N_1695);
xnor U2709 (N_2709,N_1712,N_1037);
and U2710 (N_2710,N_1401,N_1820);
and U2711 (N_2711,N_1819,N_1867);
or U2712 (N_2712,N_1733,N_1809);
or U2713 (N_2713,N_1790,N_1949);
nand U2714 (N_2714,N_1440,N_1046);
xnor U2715 (N_2715,N_1971,N_1172);
nand U2716 (N_2716,N_1898,N_1285);
xnor U2717 (N_2717,N_1677,N_1496);
and U2718 (N_2718,N_1816,N_1687);
or U2719 (N_2719,N_1586,N_1343);
nor U2720 (N_2720,N_1623,N_1397);
nand U2721 (N_2721,N_1541,N_1132);
xor U2722 (N_2722,N_1442,N_1609);
or U2723 (N_2723,N_1027,N_1994);
or U2724 (N_2724,N_1078,N_1126);
or U2725 (N_2725,N_1433,N_1038);
and U2726 (N_2726,N_1351,N_1055);
xor U2727 (N_2727,N_1861,N_1835);
or U2728 (N_2728,N_1247,N_1603);
nand U2729 (N_2729,N_1571,N_1742);
or U2730 (N_2730,N_1263,N_1689);
xnor U2731 (N_2731,N_1629,N_1873);
nand U2732 (N_2732,N_1015,N_1141);
and U2733 (N_2733,N_1924,N_1340);
nand U2734 (N_2734,N_1697,N_1969);
or U2735 (N_2735,N_1904,N_1648);
nor U2736 (N_2736,N_1998,N_1776);
or U2737 (N_2737,N_1639,N_1656);
nor U2738 (N_2738,N_1627,N_1956);
xnor U2739 (N_2739,N_1811,N_1694);
or U2740 (N_2740,N_1115,N_1276);
and U2741 (N_2741,N_1942,N_1601);
xor U2742 (N_2742,N_1137,N_1403);
xor U2743 (N_2743,N_1652,N_1625);
xnor U2744 (N_2744,N_1599,N_1607);
and U2745 (N_2745,N_1690,N_1320);
nand U2746 (N_2746,N_1443,N_1746);
nor U2747 (N_2747,N_1950,N_1968);
and U2748 (N_2748,N_1083,N_1218);
nor U2749 (N_2749,N_1741,N_1859);
and U2750 (N_2750,N_1830,N_1815);
nand U2751 (N_2751,N_1404,N_1060);
and U2752 (N_2752,N_1777,N_1546);
and U2753 (N_2753,N_1890,N_1668);
nor U2754 (N_2754,N_1582,N_1455);
nor U2755 (N_2755,N_1242,N_1367);
or U2756 (N_2756,N_1078,N_1675);
nand U2757 (N_2757,N_1970,N_1710);
xor U2758 (N_2758,N_1812,N_1379);
nor U2759 (N_2759,N_1172,N_1823);
xor U2760 (N_2760,N_1840,N_1963);
and U2761 (N_2761,N_1942,N_1275);
and U2762 (N_2762,N_1483,N_1677);
or U2763 (N_2763,N_1237,N_1415);
nor U2764 (N_2764,N_1713,N_1785);
nand U2765 (N_2765,N_1391,N_1519);
xor U2766 (N_2766,N_1056,N_1921);
nor U2767 (N_2767,N_1742,N_1548);
nor U2768 (N_2768,N_1881,N_1031);
or U2769 (N_2769,N_1567,N_1275);
xnor U2770 (N_2770,N_1130,N_1192);
xor U2771 (N_2771,N_1562,N_1927);
xnor U2772 (N_2772,N_1384,N_1868);
or U2773 (N_2773,N_1822,N_1956);
or U2774 (N_2774,N_1847,N_1196);
xor U2775 (N_2775,N_1025,N_1618);
xor U2776 (N_2776,N_1760,N_1171);
and U2777 (N_2777,N_1963,N_1050);
and U2778 (N_2778,N_1127,N_1573);
nor U2779 (N_2779,N_1722,N_1818);
xnor U2780 (N_2780,N_1893,N_1529);
or U2781 (N_2781,N_1214,N_1322);
nand U2782 (N_2782,N_1497,N_1034);
xor U2783 (N_2783,N_1912,N_1767);
or U2784 (N_2784,N_1791,N_1241);
nor U2785 (N_2785,N_1908,N_1311);
nand U2786 (N_2786,N_1729,N_1847);
xor U2787 (N_2787,N_1983,N_1991);
nand U2788 (N_2788,N_1529,N_1386);
nor U2789 (N_2789,N_1174,N_1447);
or U2790 (N_2790,N_1928,N_1390);
nor U2791 (N_2791,N_1918,N_1880);
xor U2792 (N_2792,N_1911,N_1262);
nand U2793 (N_2793,N_1194,N_1607);
nand U2794 (N_2794,N_1495,N_1402);
xor U2795 (N_2795,N_1505,N_1625);
or U2796 (N_2796,N_1717,N_1839);
xnor U2797 (N_2797,N_1528,N_1550);
nand U2798 (N_2798,N_1611,N_1148);
nor U2799 (N_2799,N_1092,N_1660);
xor U2800 (N_2800,N_1159,N_1281);
or U2801 (N_2801,N_1642,N_1396);
and U2802 (N_2802,N_1044,N_1027);
and U2803 (N_2803,N_1775,N_1361);
xor U2804 (N_2804,N_1295,N_1325);
and U2805 (N_2805,N_1843,N_1534);
nand U2806 (N_2806,N_1248,N_1587);
nor U2807 (N_2807,N_1017,N_1151);
nand U2808 (N_2808,N_1537,N_1486);
xnor U2809 (N_2809,N_1921,N_1434);
xnor U2810 (N_2810,N_1404,N_1820);
xnor U2811 (N_2811,N_1908,N_1261);
or U2812 (N_2812,N_1946,N_1909);
nand U2813 (N_2813,N_1897,N_1683);
or U2814 (N_2814,N_1629,N_1867);
nor U2815 (N_2815,N_1699,N_1774);
xor U2816 (N_2816,N_1415,N_1911);
xnor U2817 (N_2817,N_1044,N_1042);
and U2818 (N_2818,N_1623,N_1910);
xnor U2819 (N_2819,N_1756,N_1462);
nor U2820 (N_2820,N_1493,N_1199);
nand U2821 (N_2821,N_1222,N_1783);
nor U2822 (N_2822,N_1283,N_1031);
nand U2823 (N_2823,N_1401,N_1604);
xor U2824 (N_2824,N_1810,N_1795);
xnor U2825 (N_2825,N_1048,N_1340);
nand U2826 (N_2826,N_1382,N_1753);
nand U2827 (N_2827,N_1076,N_1999);
nor U2828 (N_2828,N_1172,N_1597);
or U2829 (N_2829,N_1262,N_1702);
and U2830 (N_2830,N_1005,N_1350);
nor U2831 (N_2831,N_1603,N_1465);
nor U2832 (N_2832,N_1439,N_1182);
nor U2833 (N_2833,N_1148,N_1711);
xor U2834 (N_2834,N_1534,N_1725);
and U2835 (N_2835,N_1092,N_1908);
xnor U2836 (N_2836,N_1680,N_1835);
nand U2837 (N_2837,N_1277,N_1226);
nor U2838 (N_2838,N_1756,N_1121);
nor U2839 (N_2839,N_1554,N_1978);
xor U2840 (N_2840,N_1334,N_1522);
and U2841 (N_2841,N_1490,N_1259);
and U2842 (N_2842,N_1496,N_1486);
nor U2843 (N_2843,N_1372,N_1837);
or U2844 (N_2844,N_1194,N_1464);
nor U2845 (N_2845,N_1562,N_1575);
nor U2846 (N_2846,N_1120,N_1262);
xor U2847 (N_2847,N_1187,N_1712);
nand U2848 (N_2848,N_1524,N_1188);
xnor U2849 (N_2849,N_1069,N_1144);
and U2850 (N_2850,N_1842,N_1196);
nor U2851 (N_2851,N_1249,N_1452);
and U2852 (N_2852,N_1935,N_1466);
nand U2853 (N_2853,N_1637,N_1332);
or U2854 (N_2854,N_1867,N_1261);
or U2855 (N_2855,N_1189,N_1186);
nor U2856 (N_2856,N_1652,N_1258);
xor U2857 (N_2857,N_1594,N_1763);
or U2858 (N_2858,N_1608,N_1671);
nor U2859 (N_2859,N_1559,N_1893);
and U2860 (N_2860,N_1431,N_1072);
or U2861 (N_2861,N_1343,N_1776);
nand U2862 (N_2862,N_1602,N_1434);
or U2863 (N_2863,N_1067,N_1239);
nand U2864 (N_2864,N_1085,N_1587);
or U2865 (N_2865,N_1522,N_1333);
and U2866 (N_2866,N_1779,N_1936);
nand U2867 (N_2867,N_1468,N_1750);
or U2868 (N_2868,N_1540,N_1228);
nand U2869 (N_2869,N_1965,N_1306);
and U2870 (N_2870,N_1096,N_1909);
and U2871 (N_2871,N_1335,N_1347);
nor U2872 (N_2872,N_1192,N_1928);
nor U2873 (N_2873,N_1189,N_1619);
xnor U2874 (N_2874,N_1369,N_1616);
and U2875 (N_2875,N_1761,N_1641);
and U2876 (N_2876,N_1027,N_1848);
xor U2877 (N_2877,N_1927,N_1972);
and U2878 (N_2878,N_1990,N_1149);
xnor U2879 (N_2879,N_1896,N_1771);
xnor U2880 (N_2880,N_1438,N_1971);
nand U2881 (N_2881,N_1769,N_1649);
or U2882 (N_2882,N_1750,N_1605);
xor U2883 (N_2883,N_1907,N_1123);
and U2884 (N_2884,N_1534,N_1520);
nor U2885 (N_2885,N_1047,N_1283);
and U2886 (N_2886,N_1213,N_1221);
nand U2887 (N_2887,N_1199,N_1953);
and U2888 (N_2888,N_1148,N_1142);
nor U2889 (N_2889,N_1326,N_1150);
nor U2890 (N_2890,N_1373,N_1820);
and U2891 (N_2891,N_1693,N_1050);
nor U2892 (N_2892,N_1188,N_1444);
or U2893 (N_2893,N_1038,N_1957);
nand U2894 (N_2894,N_1416,N_1780);
nand U2895 (N_2895,N_1236,N_1378);
xnor U2896 (N_2896,N_1203,N_1594);
xnor U2897 (N_2897,N_1753,N_1174);
nor U2898 (N_2898,N_1599,N_1738);
and U2899 (N_2899,N_1723,N_1876);
nor U2900 (N_2900,N_1577,N_1323);
nor U2901 (N_2901,N_1715,N_1486);
or U2902 (N_2902,N_1278,N_1473);
or U2903 (N_2903,N_1650,N_1213);
nand U2904 (N_2904,N_1330,N_1116);
and U2905 (N_2905,N_1431,N_1230);
or U2906 (N_2906,N_1381,N_1623);
nand U2907 (N_2907,N_1473,N_1370);
nand U2908 (N_2908,N_1207,N_1532);
nor U2909 (N_2909,N_1207,N_1815);
and U2910 (N_2910,N_1516,N_1224);
nand U2911 (N_2911,N_1287,N_1367);
nand U2912 (N_2912,N_1549,N_1906);
or U2913 (N_2913,N_1925,N_1811);
nor U2914 (N_2914,N_1807,N_1796);
or U2915 (N_2915,N_1314,N_1426);
xnor U2916 (N_2916,N_1106,N_1200);
xor U2917 (N_2917,N_1265,N_1574);
or U2918 (N_2918,N_1270,N_1945);
nor U2919 (N_2919,N_1063,N_1126);
or U2920 (N_2920,N_1938,N_1091);
nand U2921 (N_2921,N_1264,N_1696);
nor U2922 (N_2922,N_1532,N_1275);
xnor U2923 (N_2923,N_1640,N_1574);
or U2924 (N_2924,N_1353,N_1190);
xor U2925 (N_2925,N_1849,N_1216);
xor U2926 (N_2926,N_1203,N_1787);
and U2927 (N_2927,N_1786,N_1266);
or U2928 (N_2928,N_1895,N_1164);
nand U2929 (N_2929,N_1076,N_1789);
nand U2930 (N_2930,N_1667,N_1934);
and U2931 (N_2931,N_1344,N_1686);
and U2932 (N_2932,N_1119,N_1251);
and U2933 (N_2933,N_1906,N_1997);
or U2934 (N_2934,N_1117,N_1616);
or U2935 (N_2935,N_1730,N_1092);
nand U2936 (N_2936,N_1251,N_1834);
xor U2937 (N_2937,N_1843,N_1398);
xor U2938 (N_2938,N_1673,N_1096);
and U2939 (N_2939,N_1496,N_1029);
or U2940 (N_2940,N_1539,N_1437);
and U2941 (N_2941,N_1130,N_1051);
and U2942 (N_2942,N_1059,N_1253);
nor U2943 (N_2943,N_1361,N_1140);
nor U2944 (N_2944,N_1092,N_1404);
or U2945 (N_2945,N_1632,N_1993);
and U2946 (N_2946,N_1280,N_1038);
and U2947 (N_2947,N_1929,N_1651);
and U2948 (N_2948,N_1170,N_1480);
or U2949 (N_2949,N_1126,N_1438);
nand U2950 (N_2950,N_1985,N_1173);
nand U2951 (N_2951,N_1501,N_1750);
nor U2952 (N_2952,N_1965,N_1788);
and U2953 (N_2953,N_1326,N_1766);
xor U2954 (N_2954,N_1419,N_1224);
nor U2955 (N_2955,N_1358,N_1344);
nand U2956 (N_2956,N_1683,N_1677);
xor U2957 (N_2957,N_1485,N_1850);
nand U2958 (N_2958,N_1106,N_1631);
nand U2959 (N_2959,N_1488,N_1003);
xnor U2960 (N_2960,N_1739,N_1495);
xnor U2961 (N_2961,N_1299,N_1407);
and U2962 (N_2962,N_1654,N_1447);
or U2963 (N_2963,N_1283,N_1115);
nor U2964 (N_2964,N_1685,N_1150);
nand U2965 (N_2965,N_1877,N_1202);
nand U2966 (N_2966,N_1801,N_1037);
and U2967 (N_2967,N_1999,N_1305);
or U2968 (N_2968,N_1805,N_1512);
or U2969 (N_2969,N_1901,N_1519);
nor U2970 (N_2970,N_1988,N_1594);
xnor U2971 (N_2971,N_1678,N_1624);
or U2972 (N_2972,N_1715,N_1876);
nand U2973 (N_2973,N_1075,N_1009);
or U2974 (N_2974,N_1741,N_1784);
nand U2975 (N_2975,N_1719,N_1362);
and U2976 (N_2976,N_1074,N_1085);
nor U2977 (N_2977,N_1259,N_1401);
or U2978 (N_2978,N_1183,N_1984);
or U2979 (N_2979,N_1495,N_1210);
and U2980 (N_2980,N_1299,N_1625);
nand U2981 (N_2981,N_1325,N_1677);
nand U2982 (N_2982,N_1952,N_1139);
nor U2983 (N_2983,N_1195,N_1823);
xnor U2984 (N_2984,N_1021,N_1083);
and U2985 (N_2985,N_1584,N_1489);
xor U2986 (N_2986,N_1280,N_1091);
nor U2987 (N_2987,N_1758,N_1407);
and U2988 (N_2988,N_1731,N_1328);
and U2989 (N_2989,N_1579,N_1529);
or U2990 (N_2990,N_1636,N_1134);
nand U2991 (N_2991,N_1257,N_1211);
or U2992 (N_2992,N_1648,N_1519);
xnor U2993 (N_2993,N_1154,N_1989);
and U2994 (N_2994,N_1129,N_1654);
nand U2995 (N_2995,N_1369,N_1387);
xnor U2996 (N_2996,N_1992,N_1164);
or U2997 (N_2997,N_1185,N_1422);
and U2998 (N_2998,N_1538,N_1960);
xor U2999 (N_2999,N_1956,N_1599);
nor U3000 (N_3000,N_2602,N_2546);
and U3001 (N_3001,N_2469,N_2919);
and U3002 (N_3002,N_2764,N_2097);
nor U3003 (N_3003,N_2346,N_2292);
nor U3004 (N_3004,N_2307,N_2338);
xnor U3005 (N_3005,N_2399,N_2704);
and U3006 (N_3006,N_2630,N_2114);
and U3007 (N_3007,N_2597,N_2531);
or U3008 (N_3008,N_2418,N_2043);
and U3009 (N_3009,N_2818,N_2411);
and U3010 (N_3010,N_2805,N_2789);
nand U3011 (N_3011,N_2389,N_2500);
xnor U3012 (N_3012,N_2001,N_2695);
xor U3013 (N_3013,N_2787,N_2589);
or U3014 (N_3014,N_2314,N_2950);
and U3015 (N_3015,N_2693,N_2134);
nand U3016 (N_3016,N_2288,N_2372);
or U3017 (N_3017,N_2094,N_2203);
or U3018 (N_3018,N_2154,N_2379);
nand U3019 (N_3019,N_2049,N_2781);
nor U3020 (N_3020,N_2893,N_2096);
nand U3021 (N_3021,N_2223,N_2383);
nor U3022 (N_3022,N_2827,N_2552);
xor U3023 (N_3023,N_2286,N_2968);
or U3024 (N_3024,N_2743,N_2617);
nand U3025 (N_3025,N_2477,N_2975);
or U3026 (N_3026,N_2926,N_2988);
and U3027 (N_3027,N_2929,N_2304);
or U3028 (N_3028,N_2783,N_2875);
nor U3029 (N_3029,N_2637,N_2221);
xor U3030 (N_3030,N_2146,N_2867);
nor U3031 (N_3031,N_2756,N_2032);
or U3032 (N_3032,N_2191,N_2080);
xnor U3033 (N_3033,N_2023,N_2568);
and U3034 (N_3034,N_2206,N_2464);
and U3035 (N_3035,N_2976,N_2941);
xnor U3036 (N_3036,N_2315,N_2566);
or U3037 (N_3037,N_2054,N_2512);
nor U3038 (N_3038,N_2732,N_2339);
or U3039 (N_3039,N_2966,N_2684);
or U3040 (N_3040,N_2616,N_2951);
or U3041 (N_3041,N_2239,N_2425);
nor U3042 (N_3042,N_2141,N_2227);
and U3043 (N_3043,N_2669,N_2010);
xnor U3044 (N_3044,N_2034,N_2224);
or U3045 (N_3045,N_2924,N_2618);
nand U3046 (N_3046,N_2368,N_2397);
and U3047 (N_3047,N_2916,N_2879);
xor U3048 (N_3048,N_2085,N_2216);
xor U3049 (N_3049,N_2747,N_2712);
and U3050 (N_3050,N_2538,N_2742);
or U3051 (N_3051,N_2579,N_2631);
or U3052 (N_3052,N_2614,N_2654);
xor U3053 (N_3053,N_2907,N_2682);
xor U3054 (N_3054,N_2553,N_2884);
nand U3055 (N_3055,N_2825,N_2246);
or U3056 (N_3056,N_2606,N_2865);
xnor U3057 (N_3057,N_2840,N_2746);
and U3058 (N_3058,N_2470,N_2355);
xnor U3059 (N_3059,N_2584,N_2777);
nand U3060 (N_3060,N_2605,N_2357);
or U3061 (N_3061,N_2430,N_2878);
or U3062 (N_3062,N_2164,N_2360);
or U3063 (N_3063,N_2779,N_2627);
and U3064 (N_3064,N_2252,N_2822);
or U3065 (N_3065,N_2115,N_2422);
xnor U3066 (N_3066,N_2690,N_2086);
xnor U3067 (N_3067,N_2133,N_2258);
or U3068 (N_3068,N_2237,N_2255);
or U3069 (N_3069,N_2969,N_2895);
and U3070 (N_3070,N_2248,N_2956);
and U3071 (N_3071,N_2636,N_2699);
and U3072 (N_3072,N_2264,N_2433);
nor U3073 (N_3073,N_2717,N_2738);
nand U3074 (N_3074,N_2317,N_2110);
or U3075 (N_3075,N_2646,N_2476);
nor U3076 (N_3076,N_2665,N_2651);
or U3077 (N_3077,N_2539,N_2808);
nand U3078 (N_3078,N_2388,N_2853);
nor U3079 (N_3079,N_2656,N_2963);
nand U3080 (N_3080,N_2562,N_2015);
nor U3081 (N_3081,N_2974,N_2382);
xnor U3082 (N_3082,N_2318,N_2572);
nor U3083 (N_3083,N_2081,N_2344);
xnor U3084 (N_3084,N_2971,N_2236);
xnor U3085 (N_3085,N_2208,N_2960);
xor U3086 (N_3086,N_2782,N_2837);
xnor U3087 (N_3087,N_2495,N_2519);
nor U3088 (N_3088,N_2913,N_2809);
or U3089 (N_3089,N_2736,N_2072);
or U3090 (N_3090,N_2019,N_2432);
and U3091 (N_3091,N_2478,N_2920);
or U3092 (N_3092,N_2268,N_2269);
and U3093 (N_3093,N_2235,N_2930);
nor U3094 (N_3094,N_2554,N_2401);
xor U3095 (N_3095,N_2957,N_2600);
or U3096 (N_3096,N_2607,N_2829);
xnor U3097 (N_3097,N_2989,N_2316);
and U3098 (N_3098,N_2748,N_2226);
nor U3099 (N_3099,N_2964,N_2509);
or U3100 (N_3100,N_2551,N_2813);
xnor U3101 (N_3101,N_2250,N_2659);
nand U3102 (N_3102,N_2555,N_2864);
and U3103 (N_3103,N_2352,N_2140);
nand U3104 (N_3104,N_2341,N_2322);
or U3105 (N_3105,N_2333,N_2063);
xnor U3106 (N_3106,N_2965,N_2413);
or U3107 (N_3107,N_2168,N_2062);
and U3108 (N_3108,N_2159,N_2869);
and U3109 (N_3109,N_2726,N_2485);
and U3110 (N_3110,N_2610,N_2792);
and U3111 (N_3111,N_2423,N_2858);
nand U3112 (N_3112,N_2241,N_2267);
and U3113 (N_3113,N_2385,N_2806);
and U3114 (N_3114,N_2161,N_2922);
xnor U3115 (N_3115,N_2280,N_2508);
nand U3116 (N_3116,N_2376,N_2112);
nor U3117 (N_3117,N_2370,N_2549);
nand U3118 (N_3118,N_2045,N_2819);
nor U3119 (N_3119,N_2276,N_2939);
nor U3120 (N_3120,N_2983,N_2407);
nand U3121 (N_3121,N_2676,N_2724);
and U3122 (N_3122,N_2943,N_2300);
nor U3123 (N_3123,N_2776,N_2437);
nor U3124 (N_3124,N_2135,N_2426);
xor U3125 (N_3125,N_2127,N_2524);
or U3126 (N_3126,N_2130,N_2698);
nand U3127 (N_3127,N_2625,N_2473);
or U3128 (N_3128,N_2155,N_2612);
and U3129 (N_3129,N_2859,N_2655);
nor U3130 (N_3130,N_2163,N_2909);
xor U3131 (N_3131,N_2739,N_2041);
and U3132 (N_3132,N_2689,N_2772);
nor U3133 (N_3133,N_2728,N_2621);
nand U3134 (N_3134,N_2132,N_2557);
xnor U3135 (N_3135,N_2523,N_2028);
and U3136 (N_3136,N_2733,N_2981);
or U3137 (N_3137,N_2463,N_2752);
nor U3138 (N_3138,N_2791,N_2649);
nor U3139 (N_3139,N_2537,N_2639);
nand U3140 (N_3140,N_2103,N_2412);
nor U3141 (N_3141,N_2873,N_2369);
nor U3142 (N_3142,N_2944,N_2986);
nor U3143 (N_3143,N_2016,N_2815);
and U3144 (N_3144,N_2295,N_2581);
nor U3145 (N_3145,N_2442,N_2287);
or U3146 (N_3146,N_2243,N_2384);
or U3147 (N_3147,N_2244,N_2395);
or U3148 (N_3148,N_2079,N_2734);
nor U3149 (N_3149,N_2946,N_2457);
or U3150 (N_3150,N_2710,N_2923);
and U3151 (N_3151,N_2468,N_2414);
nor U3152 (N_3152,N_2165,N_2660);
nand U3153 (N_3153,N_2973,N_2004);
xor U3154 (N_3154,N_2011,N_2898);
nor U3155 (N_3155,N_2088,N_2419);
or U3156 (N_3156,N_2106,N_2375);
and U3157 (N_3157,N_2586,N_2018);
and U3158 (N_3158,N_2831,N_2984);
nand U3159 (N_3159,N_2679,N_2954);
or U3160 (N_3160,N_2427,N_2720);
nand U3161 (N_3161,N_2120,N_2773);
xor U3162 (N_3162,N_2598,N_2177);
xnor U3163 (N_3163,N_2501,N_2970);
nor U3164 (N_3164,N_2077,N_2632);
and U3165 (N_3165,N_2730,N_2780);
nor U3166 (N_3166,N_2441,N_2263);
or U3167 (N_3167,N_2794,N_2585);
nor U3168 (N_3168,N_2713,N_2574);
nor U3169 (N_3169,N_2703,N_2948);
xnor U3170 (N_3170,N_2741,N_2021);
or U3171 (N_3171,N_2249,N_2642);
or U3172 (N_3172,N_2569,N_2852);
and U3173 (N_3173,N_2897,N_2933);
or U3174 (N_3174,N_2047,N_2152);
xor U3175 (N_3175,N_2993,N_2391);
xor U3176 (N_3176,N_2778,N_2420);
or U3177 (N_3177,N_2821,N_2697);
nand U3178 (N_3178,N_2284,N_2325);
nand U3179 (N_3179,N_2529,N_2937);
xnor U3180 (N_3180,N_2390,N_2949);
and U3181 (N_3181,N_2836,N_2520);
or U3182 (N_3182,N_2200,N_2359);
xnor U3183 (N_3183,N_2735,N_2424);
xor U3184 (N_3184,N_2565,N_2331);
or U3185 (N_3185,N_2716,N_2417);
nor U3186 (N_3186,N_2619,N_2308);
and U3187 (N_3187,N_2351,N_2886);
and U3188 (N_3188,N_2214,N_2057);
nor U3189 (N_3189,N_2672,N_2319);
nor U3190 (N_3190,N_2447,N_2124);
xor U3191 (N_3191,N_2647,N_2013);
xnor U3192 (N_3192,N_2481,N_2256);
and U3193 (N_3193,N_2488,N_2580);
and U3194 (N_3194,N_2109,N_2222);
xor U3195 (N_3195,N_2262,N_2035);
and U3196 (N_3196,N_2193,N_2406);
and U3197 (N_3197,N_2215,N_2784);
nor U3198 (N_3198,N_2828,N_2843);
xnor U3199 (N_3199,N_2230,N_2938);
nor U3200 (N_3200,N_2686,N_2460);
xor U3201 (N_3201,N_2259,N_2876);
nand U3202 (N_3202,N_2449,N_2036);
nand U3203 (N_3203,N_2452,N_2991);
xnor U3204 (N_3204,N_2052,N_2309);
and U3205 (N_3205,N_2762,N_2816);
xnor U3206 (N_3206,N_2234,N_2472);
and U3207 (N_3207,N_2078,N_2064);
or U3208 (N_3208,N_2482,N_2877);
xor U3209 (N_3209,N_2334,N_2179);
and U3210 (N_3210,N_2925,N_2274);
and U3211 (N_3211,N_2279,N_2291);
or U3212 (N_3212,N_2595,N_2350);
xor U3213 (N_3213,N_2297,N_2148);
xor U3214 (N_3214,N_2144,N_2799);
nor U3215 (N_3215,N_2030,N_2727);
or U3216 (N_3216,N_2719,N_2910);
xor U3217 (N_3217,N_2870,N_2136);
xnor U3218 (N_3218,N_2217,N_2723);
xor U3219 (N_3219,N_2116,N_2918);
xor U3220 (N_3220,N_2113,N_2475);
nor U3221 (N_3221,N_2615,N_2498);
xor U3222 (N_3222,N_2590,N_2996);
and U3223 (N_3223,N_2891,N_2089);
and U3224 (N_3224,N_2139,N_2440);
or U3225 (N_3225,N_2471,N_2196);
nor U3226 (N_3226,N_2205,N_2172);
and U3227 (N_3227,N_2378,N_2567);
and U3228 (N_3228,N_2801,N_2131);
or U3229 (N_3229,N_2111,N_2587);
xor U3230 (N_3230,N_2219,N_2483);
or U3231 (N_3231,N_2272,N_2192);
xnor U3232 (N_3232,N_2367,N_2745);
or U3233 (N_3233,N_2305,N_2157);
or U3234 (N_3234,N_2453,N_2366);
nor U3235 (N_3235,N_2025,N_2841);
and U3236 (N_3236,N_2917,N_2622);
or U3237 (N_3237,N_2683,N_2666);
or U3238 (N_3238,N_2953,N_2521);
xor U3239 (N_3239,N_2544,N_2125);
nand U3240 (N_3240,N_2436,N_2560);
or U3241 (N_3241,N_2883,N_2990);
or U3242 (N_3242,N_2007,N_2848);
nor U3243 (N_3243,N_2181,N_2911);
nand U3244 (N_3244,N_2294,N_2972);
and U3245 (N_3245,N_2289,N_2373);
nand U3246 (N_3246,N_2790,N_2480);
and U3247 (N_3247,N_2066,N_2392);
nor U3248 (N_3248,N_2073,N_2623);
or U3249 (N_3249,N_2348,N_2663);
nand U3250 (N_3250,N_2548,N_2454);
nand U3251 (N_3251,N_2921,N_2101);
nor U3252 (N_3252,N_2074,N_2982);
xnor U3253 (N_3253,N_2564,N_2265);
nor U3254 (N_3254,N_2231,N_2402);
xor U3255 (N_3255,N_2186,N_2039);
nor U3256 (N_3256,N_2643,N_2467);
xnor U3257 (N_3257,N_2082,N_2563);
nor U3258 (N_3258,N_2980,N_2575);
or U3259 (N_3259,N_2486,N_2050);
nand U3260 (N_3260,N_2067,N_2667);
xor U3261 (N_3261,N_2635,N_2121);
xnor U3262 (N_3262,N_2516,N_2721);
xnor U3263 (N_3263,N_2296,N_2908);
and U3264 (N_3264,N_2489,N_2761);
or U3265 (N_3265,N_2823,N_2652);
and U3266 (N_3266,N_2169,N_2582);
and U3267 (N_3267,N_2803,N_2439);
nor U3268 (N_3268,N_2708,N_2505);
and U3269 (N_3269,N_2160,N_2800);
and U3270 (N_3270,N_2356,N_2814);
xnor U3271 (N_3271,N_2797,N_2995);
xnor U3272 (N_3272,N_2832,N_2588);
nor U3273 (N_3273,N_2349,N_2151);
xnor U3274 (N_3274,N_2518,N_2492);
xor U3275 (N_3275,N_2403,N_2849);
and U3276 (N_3276,N_2490,N_2942);
and U3277 (N_3277,N_2075,N_2706);
nand U3278 (N_3278,N_2012,N_2793);
nor U3279 (N_3279,N_2674,N_2170);
and U3280 (N_3280,N_2329,N_2240);
xnor U3281 (N_3281,N_2700,N_2446);
or U3282 (N_3282,N_2670,N_2664);
and U3283 (N_3283,N_2577,N_2303);
nor U3284 (N_3284,N_2657,N_2725);
and U3285 (N_3285,N_2311,N_2484);
and U3286 (N_3286,N_2648,N_2421);
and U3287 (N_3287,N_2902,N_2817);
or U3288 (N_3288,N_2961,N_2129);
or U3289 (N_3289,N_2149,N_2673);
nand U3290 (N_3290,N_2839,N_2641);
xor U3291 (N_3291,N_2099,N_2507);
nor U3292 (N_3292,N_2861,N_2466);
or U3293 (N_3293,N_2358,N_2451);
nor U3294 (N_3294,N_2091,N_2844);
xnor U3295 (N_3295,N_2601,N_2556);
xnor U3296 (N_3296,N_2962,N_2293);
and U3297 (N_3297,N_2158,N_2985);
and U3298 (N_3298,N_2765,N_2024);
and U3299 (N_3299,N_2715,N_2461);
nand U3300 (N_3300,N_2270,N_2826);
xnor U3301 (N_3301,N_2978,N_2824);
xnor U3302 (N_3302,N_2633,N_2688);
nor U3303 (N_3303,N_2225,N_2150);
or U3304 (N_3304,N_2530,N_2095);
nor U3305 (N_3305,N_2434,N_2046);
nor U3306 (N_3306,N_2999,N_2448);
nor U3307 (N_3307,N_2198,N_2330);
and U3308 (N_3308,N_2137,N_2934);
nor U3309 (N_3309,N_2044,N_2758);
xnor U3310 (N_3310,N_2261,N_2583);
and U3311 (N_3311,N_2108,N_2324);
or U3312 (N_3312,N_2428,N_2210);
or U3313 (N_3313,N_2802,N_2202);
nand U3314 (N_3314,N_2894,N_2438);
nor U3315 (N_3315,N_2662,N_2611);
nor U3316 (N_3316,N_2009,N_2854);
or U3317 (N_3317,N_2228,N_2107);
nand U3318 (N_3318,N_2887,N_2740);
xnor U3319 (N_3319,N_2055,N_2415);
xnor U3320 (N_3320,N_2022,N_2026);
nand U3321 (N_3321,N_2098,N_2709);
nor U3322 (N_3322,N_2685,N_2872);
or U3323 (N_3323,N_2851,N_2638);
or U3324 (N_3324,N_2644,N_2737);
xor U3325 (N_3325,N_2257,N_2603);
nor U3326 (N_3326,N_2014,N_2543);
nand U3327 (N_3327,N_2533,N_2232);
and U3328 (N_3328,N_2207,N_2932);
nor U3329 (N_3329,N_2213,N_2871);
nand U3330 (N_3330,N_2393,N_2608);
nor U3331 (N_3331,N_2573,N_2834);
and U3332 (N_3332,N_2184,N_2763);
and U3333 (N_3333,N_2542,N_2194);
nand U3334 (N_3334,N_2211,N_2889);
and U3335 (N_3335,N_2326,N_2890);
nand U3336 (N_3336,N_2313,N_2197);
xor U3337 (N_3337,N_2040,N_2405);
xor U3338 (N_3338,N_2795,N_2218);
nor U3339 (N_3339,N_2510,N_2102);
nand U3340 (N_3340,N_2253,N_2431);
and U3341 (N_3341,N_2061,N_2714);
nand U3342 (N_3342,N_2002,N_2335);
nand U3343 (N_3343,N_2347,N_2327);
xor U3344 (N_3344,N_2178,N_2033);
nand U3345 (N_3345,N_2354,N_2857);
nand U3346 (N_3346,N_2628,N_2275);
nor U3347 (N_3347,N_2759,N_2084);
nor U3348 (N_3348,N_2842,N_2398);
nor U3349 (N_3349,N_2076,N_2337);
and U3350 (N_3350,N_2320,N_2374);
or U3351 (N_3351,N_2912,N_2535);
nand U3352 (N_3352,N_2229,N_2811);
xor U3353 (N_3353,N_2020,N_2201);
and U3354 (N_3354,N_2513,N_2173);
and U3355 (N_3355,N_2182,N_2506);
and U3356 (N_3356,N_2245,N_2497);
nand U3357 (N_3357,N_2195,N_2070);
and U3358 (N_3358,N_2687,N_2408);
or U3359 (N_3359,N_2266,N_2845);
or U3360 (N_3360,N_2053,N_2282);
nand U3361 (N_3361,N_2429,N_2927);
nor U3362 (N_3362,N_2435,N_2754);
or U3363 (N_3363,N_2576,N_2692);
xor U3364 (N_3364,N_2896,N_2145);
xnor U3365 (N_3365,N_2947,N_2517);
xnor U3366 (N_3366,N_2380,N_2534);
and U3367 (N_3367,N_2166,N_2042);
xnor U3368 (N_3368,N_2238,N_2138);
xnor U3369 (N_3369,N_2998,N_2955);
nor U3370 (N_3370,N_2992,N_2882);
nand U3371 (N_3371,N_2979,N_2561);
nand U3372 (N_3372,N_2705,N_2658);
xnor U3373 (N_3373,N_2536,N_2550);
and U3374 (N_3374,N_2892,N_2959);
or U3375 (N_3375,N_2456,N_2702);
or U3376 (N_3376,N_2522,N_2846);
nand U3377 (N_3377,N_2620,N_2167);
nor U3378 (N_3378,N_2087,N_2915);
nand U3379 (N_3379,N_2885,N_2190);
or U3380 (N_3380,N_2571,N_2031);
or U3381 (N_3381,N_2812,N_2596);
nor U3382 (N_3382,N_2353,N_2547);
xor U3383 (N_3383,N_2301,N_2668);
and U3384 (N_3384,N_2377,N_2162);
and U3385 (N_3385,N_2526,N_2122);
xor U3386 (N_3386,N_2835,N_2796);
and U3387 (N_3387,N_2410,N_2008);
and U3388 (N_3388,N_2958,N_2068);
nand U3389 (N_3389,N_2459,N_2903);
nor U3390 (N_3390,N_2465,N_2528);
xnor U3391 (N_3391,N_2675,N_2254);
nand U3392 (N_3392,N_2770,N_2174);
nor U3393 (N_3393,N_2092,N_2499);
and U3394 (N_3394,N_2940,N_2118);
xnor U3395 (N_3395,N_2694,N_2204);
xor U3396 (N_3396,N_2545,N_2126);
nand U3397 (N_3397,N_2455,N_2677);
nor U3398 (N_3398,N_2409,N_2065);
nand U3399 (N_3399,N_2786,N_2570);
or U3400 (N_3400,N_2931,N_2678);
or U3401 (N_3401,N_2212,N_2005);
and U3402 (N_3402,N_2462,N_2775);
or U3403 (N_3403,N_2807,N_2365);
nor U3404 (N_3404,N_2302,N_2967);
xnor U3405 (N_3405,N_2119,N_2310);
nor U3406 (N_3406,N_2833,N_2592);
and U3407 (N_3407,N_2640,N_2935);
xnor U3408 (N_3408,N_2634,N_2624);
xnor U3409 (N_3409,N_2671,N_2604);
nand U3410 (N_3410,N_2880,N_2502);
xnor U3411 (N_3411,N_2128,N_2900);
and U3412 (N_3412,N_2850,N_2711);
nand U3413 (N_3413,N_2593,N_2363);
xnor U3414 (N_3414,N_2771,N_2707);
xor U3415 (N_3415,N_2729,N_2613);
nand U3416 (N_3416,N_2491,N_2209);
or U3417 (N_3417,N_2540,N_2340);
or U3418 (N_3418,N_2856,N_2220);
and U3419 (N_3419,N_2760,N_2650);
xnor U3420 (N_3420,N_2281,N_2361);
and U3421 (N_3421,N_2977,N_2751);
and U3422 (N_3422,N_2629,N_2945);
and U3423 (N_3423,N_2874,N_2810);
nor U3424 (N_3424,N_2493,N_2285);
nand U3425 (N_3425,N_2060,N_2450);
and U3426 (N_3426,N_2290,N_2804);
nand U3427 (N_3427,N_2645,N_2404);
nor U3428 (N_3428,N_2994,N_2444);
nand U3429 (N_3429,N_2371,N_2511);
xnor U3430 (N_3430,N_2003,N_2183);
nand U3431 (N_3431,N_2006,N_2525);
nand U3432 (N_3432,N_2798,N_2474);
nand U3433 (N_3433,N_2416,N_2038);
or U3434 (N_3434,N_2680,N_2071);
and U3435 (N_3435,N_2323,N_2386);
and U3436 (N_3436,N_2866,N_2503);
xor U3437 (N_3437,N_2000,N_2626);
nor U3438 (N_3438,N_2901,N_2189);
nand U3439 (N_3439,N_2153,N_2271);
and U3440 (N_3440,N_2863,N_2744);
nand U3441 (N_3441,N_2753,N_2928);
nor U3442 (N_3442,N_2769,N_2750);
or U3443 (N_3443,N_2188,N_2396);
or U3444 (N_3444,N_2987,N_2105);
nor U3445 (N_3445,N_2532,N_2862);
xor U3446 (N_3446,N_2696,N_2722);
xor U3447 (N_3447,N_2661,N_2701);
and U3448 (N_3448,N_2278,N_2653);
or U3449 (N_3449,N_2343,N_2541);
nor U3450 (N_3450,N_2336,N_2906);
xor U3451 (N_3451,N_2069,N_2381);
xnor U3452 (N_3452,N_2306,N_2599);
nor U3453 (N_3453,N_2233,N_2051);
and U3454 (N_3454,N_2594,N_2558);
or U3455 (N_3455,N_2820,N_2914);
nor U3456 (N_3456,N_2283,N_2838);
or U3457 (N_3457,N_2056,N_2156);
nor U3458 (N_3458,N_2242,N_2952);
or U3459 (N_3459,N_2731,N_2090);
nor U3460 (N_3460,N_2847,N_2123);
and U3461 (N_3461,N_2681,N_2117);
and U3462 (N_3462,N_2504,N_2027);
and U3463 (N_3463,N_2479,N_2768);
or U3464 (N_3464,N_2048,N_2345);
xnor U3465 (N_3465,N_2171,N_2199);
nor U3466 (N_3466,N_2691,N_2757);
and U3467 (N_3467,N_2364,N_2273);
and U3468 (N_3468,N_2868,N_2609);
or U3469 (N_3469,N_2394,N_2527);
nand U3470 (N_3470,N_2029,N_2904);
nand U3471 (N_3471,N_2083,N_2591);
nor U3472 (N_3472,N_2888,N_2362);
xnor U3473 (N_3473,N_2514,N_2830);
nand U3474 (N_3474,N_2755,N_2312);
xnor U3475 (N_3475,N_2142,N_2881);
nor U3476 (N_3476,N_2342,N_2104);
and U3477 (N_3477,N_2443,N_2147);
or U3478 (N_3478,N_2905,N_2515);
or U3479 (N_3479,N_2037,N_2718);
and U3480 (N_3480,N_2767,N_2785);
and U3481 (N_3481,N_2017,N_2321);
and U3482 (N_3482,N_2185,N_2277);
xor U3483 (N_3483,N_2774,N_2059);
nand U3484 (N_3484,N_2400,N_2855);
or U3485 (N_3485,N_2387,N_2445);
or U3486 (N_3486,N_2180,N_2175);
and U3487 (N_3487,N_2860,N_2559);
nor U3488 (N_3488,N_2458,N_2766);
nand U3489 (N_3489,N_2260,N_2058);
and U3490 (N_3490,N_2899,N_2247);
nand U3491 (N_3491,N_2494,N_2251);
and U3492 (N_3492,N_2749,N_2176);
and U3493 (N_3493,N_2487,N_2332);
xor U3494 (N_3494,N_2936,N_2298);
nor U3495 (N_3495,N_2997,N_2578);
and U3496 (N_3496,N_2093,N_2328);
and U3497 (N_3497,N_2143,N_2788);
and U3498 (N_3498,N_2100,N_2496);
xnor U3499 (N_3499,N_2299,N_2187);
or U3500 (N_3500,N_2198,N_2151);
and U3501 (N_3501,N_2064,N_2283);
and U3502 (N_3502,N_2020,N_2960);
or U3503 (N_3503,N_2172,N_2244);
xnor U3504 (N_3504,N_2213,N_2459);
and U3505 (N_3505,N_2090,N_2785);
nor U3506 (N_3506,N_2506,N_2241);
and U3507 (N_3507,N_2192,N_2649);
xor U3508 (N_3508,N_2862,N_2915);
nand U3509 (N_3509,N_2351,N_2111);
or U3510 (N_3510,N_2310,N_2885);
and U3511 (N_3511,N_2917,N_2143);
nor U3512 (N_3512,N_2837,N_2430);
nand U3513 (N_3513,N_2936,N_2520);
xnor U3514 (N_3514,N_2633,N_2591);
and U3515 (N_3515,N_2170,N_2604);
nor U3516 (N_3516,N_2145,N_2937);
nand U3517 (N_3517,N_2892,N_2523);
nor U3518 (N_3518,N_2674,N_2196);
nand U3519 (N_3519,N_2437,N_2212);
and U3520 (N_3520,N_2550,N_2527);
xnor U3521 (N_3521,N_2891,N_2099);
nand U3522 (N_3522,N_2002,N_2870);
and U3523 (N_3523,N_2607,N_2429);
nand U3524 (N_3524,N_2687,N_2837);
or U3525 (N_3525,N_2865,N_2908);
nand U3526 (N_3526,N_2676,N_2742);
and U3527 (N_3527,N_2760,N_2077);
xnor U3528 (N_3528,N_2078,N_2050);
or U3529 (N_3529,N_2062,N_2865);
nor U3530 (N_3530,N_2847,N_2900);
or U3531 (N_3531,N_2753,N_2888);
xnor U3532 (N_3532,N_2616,N_2701);
xnor U3533 (N_3533,N_2090,N_2320);
nor U3534 (N_3534,N_2434,N_2548);
or U3535 (N_3535,N_2542,N_2471);
and U3536 (N_3536,N_2346,N_2591);
nor U3537 (N_3537,N_2988,N_2024);
nor U3538 (N_3538,N_2920,N_2493);
nor U3539 (N_3539,N_2199,N_2368);
and U3540 (N_3540,N_2145,N_2128);
nor U3541 (N_3541,N_2353,N_2133);
nand U3542 (N_3542,N_2762,N_2130);
xor U3543 (N_3543,N_2592,N_2714);
nand U3544 (N_3544,N_2739,N_2934);
and U3545 (N_3545,N_2825,N_2151);
nor U3546 (N_3546,N_2905,N_2612);
nand U3547 (N_3547,N_2760,N_2216);
xnor U3548 (N_3548,N_2896,N_2887);
or U3549 (N_3549,N_2920,N_2357);
and U3550 (N_3550,N_2050,N_2984);
nand U3551 (N_3551,N_2386,N_2142);
and U3552 (N_3552,N_2387,N_2222);
nor U3553 (N_3553,N_2765,N_2445);
or U3554 (N_3554,N_2318,N_2965);
nor U3555 (N_3555,N_2634,N_2064);
xnor U3556 (N_3556,N_2803,N_2849);
nand U3557 (N_3557,N_2618,N_2204);
nor U3558 (N_3558,N_2052,N_2331);
nor U3559 (N_3559,N_2248,N_2478);
or U3560 (N_3560,N_2137,N_2886);
nand U3561 (N_3561,N_2856,N_2136);
and U3562 (N_3562,N_2604,N_2759);
xnor U3563 (N_3563,N_2726,N_2408);
nor U3564 (N_3564,N_2809,N_2976);
and U3565 (N_3565,N_2639,N_2168);
xor U3566 (N_3566,N_2762,N_2427);
xnor U3567 (N_3567,N_2190,N_2396);
nand U3568 (N_3568,N_2610,N_2764);
xnor U3569 (N_3569,N_2902,N_2005);
nand U3570 (N_3570,N_2056,N_2594);
xnor U3571 (N_3571,N_2994,N_2760);
and U3572 (N_3572,N_2404,N_2316);
nor U3573 (N_3573,N_2151,N_2704);
nand U3574 (N_3574,N_2376,N_2718);
nand U3575 (N_3575,N_2189,N_2026);
and U3576 (N_3576,N_2592,N_2467);
xnor U3577 (N_3577,N_2798,N_2887);
nor U3578 (N_3578,N_2273,N_2901);
nand U3579 (N_3579,N_2050,N_2815);
xor U3580 (N_3580,N_2129,N_2142);
nor U3581 (N_3581,N_2056,N_2475);
nand U3582 (N_3582,N_2766,N_2660);
nand U3583 (N_3583,N_2137,N_2286);
nor U3584 (N_3584,N_2453,N_2887);
and U3585 (N_3585,N_2641,N_2018);
nor U3586 (N_3586,N_2131,N_2471);
nand U3587 (N_3587,N_2482,N_2864);
nand U3588 (N_3588,N_2638,N_2989);
or U3589 (N_3589,N_2548,N_2839);
or U3590 (N_3590,N_2173,N_2768);
and U3591 (N_3591,N_2653,N_2395);
and U3592 (N_3592,N_2238,N_2773);
or U3593 (N_3593,N_2307,N_2495);
nor U3594 (N_3594,N_2053,N_2414);
xnor U3595 (N_3595,N_2034,N_2392);
or U3596 (N_3596,N_2681,N_2708);
and U3597 (N_3597,N_2019,N_2497);
nand U3598 (N_3598,N_2650,N_2947);
or U3599 (N_3599,N_2326,N_2826);
and U3600 (N_3600,N_2585,N_2789);
or U3601 (N_3601,N_2984,N_2014);
or U3602 (N_3602,N_2574,N_2807);
nor U3603 (N_3603,N_2594,N_2535);
nor U3604 (N_3604,N_2655,N_2925);
and U3605 (N_3605,N_2077,N_2130);
nor U3606 (N_3606,N_2841,N_2440);
xnor U3607 (N_3607,N_2583,N_2189);
nand U3608 (N_3608,N_2145,N_2534);
or U3609 (N_3609,N_2704,N_2365);
nand U3610 (N_3610,N_2251,N_2896);
nand U3611 (N_3611,N_2629,N_2704);
xnor U3612 (N_3612,N_2707,N_2017);
xor U3613 (N_3613,N_2391,N_2972);
and U3614 (N_3614,N_2977,N_2832);
nand U3615 (N_3615,N_2051,N_2218);
nor U3616 (N_3616,N_2838,N_2557);
or U3617 (N_3617,N_2424,N_2535);
or U3618 (N_3618,N_2640,N_2539);
nor U3619 (N_3619,N_2137,N_2843);
and U3620 (N_3620,N_2700,N_2280);
nor U3621 (N_3621,N_2577,N_2835);
or U3622 (N_3622,N_2312,N_2619);
or U3623 (N_3623,N_2560,N_2448);
and U3624 (N_3624,N_2853,N_2510);
and U3625 (N_3625,N_2196,N_2693);
or U3626 (N_3626,N_2176,N_2209);
nand U3627 (N_3627,N_2248,N_2624);
or U3628 (N_3628,N_2666,N_2633);
nand U3629 (N_3629,N_2830,N_2074);
nand U3630 (N_3630,N_2733,N_2311);
nand U3631 (N_3631,N_2726,N_2569);
nor U3632 (N_3632,N_2301,N_2971);
and U3633 (N_3633,N_2639,N_2503);
nand U3634 (N_3634,N_2960,N_2635);
or U3635 (N_3635,N_2305,N_2201);
nor U3636 (N_3636,N_2754,N_2495);
or U3637 (N_3637,N_2576,N_2467);
or U3638 (N_3638,N_2780,N_2134);
nor U3639 (N_3639,N_2324,N_2032);
or U3640 (N_3640,N_2814,N_2730);
xnor U3641 (N_3641,N_2473,N_2813);
nor U3642 (N_3642,N_2257,N_2552);
nand U3643 (N_3643,N_2630,N_2853);
xnor U3644 (N_3644,N_2402,N_2305);
nand U3645 (N_3645,N_2401,N_2742);
or U3646 (N_3646,N_2769,N_2487);
and U3647 (N_3647,N_2931,N_2871);
and U3648 (N_3648,N_2409,N_2053);
xnor U3649 (N_3649,N_2088,N_2878);
nor U3650 (N_3650,N_2554,N_2786);
or U3651 (N_3651,N_2611,N_2179);
xor U3652 (N_3652,N_2358,N_2910);
nand U3653 (N_3653,N_2306,N_2804);
nor U3654 (N_3654,N_2733,N_2970);
nand U3655 (N_3655,N_2383,N_2081);
nor U3656 (N_3656,N_2400,N_2762);
or U3657 (N_3657,N_2508,N_2755);
or U3658 (N_3658,N_2280,N_2241);
and U3659 (N_3659,N_2750,N_2251);
nor U3660 (N_3660,N_2476,N_2301);
nor U3661 (N_3661,N_2614,N_2767);
nor U3662 (N_3662,N_2850,N_2848);
or U3663 (N_3663,N_2144,N_2822);
or U3664 (N_3664,N_2661,N_2386);
and U3665 (N_3665,N_2183,N_2958);
nand U3666 (N_3666,N_2743,N_2064);
nor U3667 (N_3667,N_2101,N_2395);
and U3668 (N_3668,N_2015,N_2732);
or U3669 (N_3669,N_2754,N_2809);
nor U3670 (N_3670,N_2979,N_2246);
xor U3671 (N_3671,N_2845,N_2531);
nor U3672 (N_3672,N_2291,N_2342);
nor U3673 (N_3673,N_2028,N_2856);
nor U3674 (N_3674,N_2103,N_2476);
xnor U3675 (N_3675,N_2587,N_2030);
or U3676 (N_3676,N_2495,N_2524);
xnor U3677 (N_3677,N_2645,N_2300);
xnor U3678 (N_3678,N_2048,N_2136);
nand U3679 (N_3679,N_2283,N_2746);
nor U3680 (N_3680,N_2538,N_2062);
or U3681 (N_3681,N_2494,N_2421);
or U3682 (N_3682,N_2566,N_2304);
nand U3683 (N_3683,N_2310,N_2438);
and U3684 (N_3684,N_2322,N_2135);
nand U3685 (N_3685,N_2422,N_2186);
and U3686 (N_3686,N_2590,N_2534);
nand U3687 (N_3687,N_2460,N_2557);
nor U3688 (N_3688,N_2639,N_2287);
xor U3689 (N_3689,N_2425,N_2746);
nor U3690 (N_3690,N_2059,N_2989);
xor U3691 (N_3691,N_2462,N_2900);
nor U3692 (N_3692,N_2106,N_2535);
xor U3693 (N_3693,N_2655,N_2443);
xor U3694 (N_3694,N_2237,N_2163);
or U3695 (N_3695,N_2447,N_2482);
or U3696 (N_3696,N_2544,N_2035);
xor U3697 (N_3697,N_2797,N_2348);
nor U3698 (N_3698,N_2171,N_2524);
nand U3699 (N_3699,N_2185,N_2152);
or U3700 (N_3700,N_2506,N_2835);
xnor U3701 (N_3701,N_2273,N_2380);
xor U3702 (N_3702,N_2243,N_2798);
nand U3703 (N_3703,N_2296,N_2318);
nor U3704 (N_3704,N_2972,N_2053);
xor U3705 (N_3705,N_2792,N_2277);
and U3706 (N_3706,N_2339,N_2158);
xnor U3707 (N_3707,N_2633,N_2614);
nor U3708 (N_3708,N_2380,N_2790);
xor U3709 (N_3709,N_2858,N_2120);
nor U3710 (N_3710,N_2694,N_2332);
xnor U3711 (N_3711,N_2046,N_2655);
nor U3712 (N_3712,N_2013,N_2572);
nor U3713 (N_3713,N_2286,N_2203);
or U3714 (N_3714,N_2480,N_2091);
nor U3715 (N_3715,N_2369,N_2612);
nand U3716 (N_3716,N_2215,N_2369);
nor U3717 (N_3717,N_2533,N_2393);
nand U3718 (N_3718,N_2409,N_2640);
xor U3719 (N_3719,N_2832,N_2055);
xor U3720 (N_3720,N_2201,N_2527);
and U3721 (N_3721,N_2721,N_2563);
xor U3722 (N_3722,N_2148,N_2545);
or U3723 (N_3723,N_2863,N_2564);
nor U3724 (N_3724,N_2994,N_2338);
and U3725 (N_3725,N_2316,N_2162);
and U3726 (N_3726,N_2726,N_2459);
xor U3727 (N_3727,N_2895,N_2100);
or U3728 (N_3728,N_2322,N_2497);
and U3729 (N_3729,N_2796,N_2939);
nor U3730 (N_3730,N_2299,N_2471);
nand U3731 (N_3731,N_2318,N_2292);
nand U3732 (N_3732,N_2405,N_2918);
and U3733 (N_3733,N_2415,N_2366);
nand U3734 (N_3734,N_2265,N_2493);
and U3735 (N_3735,N_2443,N_2908);
nor U3736 (N_3736,N_2918,N_2825);
nor U3737 (N_3737,N_2341,N_2067);
or U3738 (N_3738,N_2631,N_2742);
xnor U3739 (N_3739,N_2374,N_2005);
and U3740 (N_3740,N_2332,N_2728);
nor U3741 (N_3741,N_2055,N_2241);
and U3742 (N_3742,N_2584,N_2478);
nand U3743 (N_3743,N_2281,N_2962);
nor U3744 (N_3744,N_2556,N_2830);
xnor U3745 (N_3745,N_2300,N_2668);
nand U3746 (N_3746,N_2337,N_2149);
or U3747 (N_3747,N_2336,N_2150);
and U3748 (N_3748,N_2708,N_2001);
nand U3749 (N_3749,N_2113,N_2359);
nand U3750 (N_3750,N_2188,N_2624);
nand U3751 (N_3751,N_2165,N_2787);
nand U3752 (N_3752,N_2206,N_2304);
nor U3753 (N_3753,N_2688,N_2839);
and U3754 (N_3754,N_2011,N_2579);
nand U3755 (N_3755,N_2736,N_2194);
xnor U3756 (N_3756,N_2685,N_2328);
nand U3757 (N_3757,N_2856,N_2083);
and U3758 (N_3758,N_2365,N_2453);
and U3759 (N_3759,N_2689,N_2532);
xnor U3760 (N_3760,N_2969,N_2677);
nand U3761 (N_3761,N_2895,N_2431);
and U3762 (N_3762,N_2931,N_2877);
nor U3763 (N_3763,N_2516,N_2947);
nand U3764 (N_3764,N_2512,N_2850);
and U3765 (N_3765,N_2930,N_2908);
or U3766 (N_3766,N_2797,N_2067);
nor U3767 (N_3767,N_2054,N_2034);
nand U3768 (N_3768,N_2424,N_2654);
nor U3769 (N_3769,N_2849,N_2282);
and U3770 (N_3770,N_2494,N_2391);
xnor U3771 (N_3771,N_2994,N_2116);
nor U3772 (N_3772,N_2668,N_2752);
xor U3773 (N_3773,N_2888,N_2078);
nor U3774 (N_3774,N_2027,N_2859);
or U3775 (N_3775,N_2888,N_2704);
nor U3776 (N_3776,N_2418,N_2830);
and U3777 (N_3777,N_2250,N_2162);
and U3778 (N_3778,N_2212,N_2014);
nor U3779 (N_3779,N_2355,N_2917);
nor U3780 (N_3780,N_2773,N_2905);
or U3781 (N_3781,N_2265,N_2803);
nor U3782 (N_3782,N_2483,N_2833);
nand U3783 (N_3783,N_2070,N_2939);
and U3784 (N_3784,N_2896,N_2639);
or U3785 (N_3785,N_2970,N_2212);
nand U3786 (N_3786,N_2935,N_2663);
xnor U3787 (N_3787,N_2894,N_2469);
nor U3788 (N_3788,N_2962,N_2412);
or U3789 (N_3789,N_2439,N_2419);
nand U3790 (N_3790,N_2064,N_2620);
nand U3791 (N_3791,N_2741,N_2313);
nand U3792 (N_3792,N_2488,N_2148);
or U3793 (N_3793,N_2108,N_2684);
nand U3794 (N_3794,N_2759,N_2501);
and U3795 (N_3795,N_2076,N_2802);
nor U3796 (N_3796,N_2719,N_2169);
xor U3797 (N_3797,N_2825,N_2863);
nand U3798 (N_3798,N_2303,N_2706);
nand U3799 (N_3799,N_2904,N_2512);
or U3800 (N_3800,N_2809,N_2753);
xnor U3801 (N_3801,N_2505,N_2861);
nand U3802 (N_3802,N_2873,N_2344);
nor U3803 (N_3803,N_2478,N_2301);
nand U3804 (N_3804,N_2217,N_2132);
nand U3805 (N_3805,N_2592,N_2063);
and U3806 (N_3806,N_2534,N_2780);
or U3807 (N_3807,N_2612,N_2213);
and U3808 (N_3808,N_2697,N_2429);
xor U3809 (N_3809,N_2769,N_2022);
xnor U3810 (N_3810,N_2605,N_2983);
xnor U3811 (N_3811,N_2302,N_2303);
xnor U3812 (N_3812,N_2089,N_2615);
and U3813 (N_3813,N_2173,N_2778);
or U3814 (N_3814,N_2645,N_2349);
nor U3815 (N_3815,N_2242,N_2415);
xnor U3816 (N_3816,N_2664,N_2360);
nor U3817 (N_3817,N_2833,N_2107);
or U3818 (N_3818,N_2790,N_2218);
or U3819 (N_3819,N_2333,N_2540);
nand U3820 (N_3820,N_2322,N_2665);
nor U3821 (N_3821,N_2998,N_2402);
nor U3822 (N_3822,N_2809,N_2080);
or U3823 (N_3823,N_2218,N_2652);
and U3824 (N_3824,N_2024,N_2968);
and U3825 (N_3825,N_2818,N_2559);
xor U3826 (N_3826,N_2920,N_2312);
and U3827 (N_3827,N_2778,N_2247);
nor U3828 (N_3828,N_2080,N_2670);
and U3829 (N_3829,N_2988,N_2820);
nand U3830 (N_3830,N_2569,N_2727);
nor U3831 (N_3831,N_2293,N_2156);
and U3832 (N_3832,N_2089,N_2579);
nand U3833 (N_3833,N_2290,N_2725);
nor U3834 (N_3834,N_2902,N_2768);
xor U3835 (N_3835,N_2478,N_2854);
and U3836 (N_3836,N_2124,N_2081);
nor U3837 (N_3837,N_2764,N_2070);
nor U3838 (N_3838,N_2075,N_2499);
and U3839 (N_3839,N_2313,N_2419);
xnor U3840 (N_3840,N_2379,N_2988);
nor U3841 (N_3841,N_2895,N_2838);
or U3842 (N_3842,N_2817,N_2115);
or U3843 (N_3843,N_2270,N_2137);
or U3844 (N_3844,N_2786,N_2442);
or U3845 (N_3845,N_2608,N_2132);
nor U3846 (N_3846,N_2849,N_2864);
and U3847 (N_3847,N_2195,N_2412);
and U3848 (N_3848,N_2976,N_2754);
nor U3849 (N_3849,N_2375,N_2809);
and U3850 (N_3850,N_2649,N_2772);
nand U3851 (N_3851,N_2520,N_2618);
nand U3852 (N_3852,N_2750,N_2372);
nand U3853 (N_3853,N_2962,N_2789);
or U3854 (N_3854,N_2198,N_2608);
and U3855 (N_3855,N_2702,N_2818);
and U3856 (N_3856,N_2331,N_2303);
xnor U3857 (N_3857,N_2075,N_2128);
xnor U3858 (N_3858,N_2814,N_2385);
or U3859 (N_3859,N_2168,N_2773);
nor U3860 (N_3860,N_2911,N_2327);
or U3861 (N_3861,N_2521,N_2477);
or U3862 (N_3862,N_2470,N_2636);
nand U3863 (N_3863,N_2424,N_2119);
nor U3864 (N_3864,N_2383,N_2681);
xor U3865 (N_3865,N_2607,N_2659);
nand U3866 (N_3866,N_2643,N_2723);
nor U3867 (N_3867,N_2866,N_2380);
nand U3868 (N_3868,N_2311,N_2408);
nor U3869 (N_3869,N_2340,N_2498);
and U3870 (N_3870,N_2241,N_2209);
xor U3871 (N_3871,N_2337,N_2558);
or U3872 (N_3872,N_2680,N_2306);
or U3873 (N_3873,N_2196,N_2003);
nor U3874 (N_3874,N_2836,N_2011);
nor U3875 (N_3875,N_2065,N_2672);
xor U3876 (N_3876,N_2143,N_2815);
xor U3877 (N_3877,N_2131,N_2052);
xnor U3878 (N_3878,N_2776,N_2804);
xor U3879 (N_3879,N_2672,N_2662);
xnor U3880 (N_3880,N_2991,N_2444);
or U3881 (N_3881,N_2998,N_2267);
xor U3882 (N_3882,N_2404,N_2012);
and U3883 (N_3883,N_2506,N_2485);
and U3884 (N_3884,N_2627,N_2700);
xnor U3885 (N_3885,N_2216,N_2391);
nor U3886 (N_3886,N_2912,N_2074);
xnor U3887 (N_3887,N_2208,N_2713);
or U3888 (N_3888,N_2133,N_2950);
nand U3889 (N_3889,N_2337,N_2207);
nand U3890 (N_3890,N_2924,N_2369);
or U3891 (N_3891,N_2779,N_2935);
xor U3892 (N_3892,N_2024,N_2653);
or U3893 (N_3893,N_2258,N_2002);
nor U3894 (N_3894,N_2063,N_2389);
or U3895 (N_3895,N_2942,N_2525);
or U3896 (N_3896,N_2339,N_2618);
xor U3897 (N_3897,N_2767,N_2086);
or U3898 (N_3898,N_2736,N_2535);
nand U3899 (N_3899,N_2596,N_2253);
nor U3900 (N_3900,N_2549,N_2134);
nand U3901 (N_3901,N_2178,N_2967);
nand U3902 (N_3902,N_2260,N_2561);
or U3903 (N_3903,N_2494,N_2294);
nand U3904 (N_3904,N_2935,N_2061);
nor U3905 (N_3905,N_2220,N_2799);
nand U3906 (N_3906,N_2341,N_2664);
nand U3907 (N_3907,N_2994,N_2344);
xor U3908 (N_3908,N_2118,N_2953);
and U3909 (N_3909,N_2262,N_2259);
nor U3910 (N_3910,N_2839,N_2030);
xnor U3911 (N_3911,N_2565,N_2359);
and U3912 (N_3912,N_2487,N_2912);
nand U3913 (N_3913,N_2012,N_2050);
and U3914 (N_3914,N_2954,N_2470);
or U3915 (N_3915,N_2969,N_2194);
xnor U3916 (N_3916,N_2683,N_2445);
nor U3917 (N_3917,N_2051,N_2710);
or U3918 (N_3918,N_2099,N_2607);
and U3919 (N_3919,N_2533,N_2794);
nand U3920 (N_3920,N_2126,N_2726);
and U3921 (N_3921,N_2966,N_2372);
nand U3922 (N_3922,N_2396,N_2098);
or U3923 (N_3923,N_2709,N_2555);
nor U3924 (N_3924,N_2936,N_2246);
or U3925 (N_3925,N_2542,N_2107);
nor U3926 (N_3926,N_2026,N_2519);
nand U3927 (N_3927,N_2844,N_2348);
xor U3928 (N_3928,N_2479,N_2375);
and U3929 (N_3929,N_2945,N_2691);
nand U3930 (N_3930,N_2123,N_2308);
and U3931 (N_3931,N_2107,N_2140);
nor U3932 (N_3932,N_2834,N_2271);
and U3933 (N_3933,N_2133,N_2592);
nand U3934 (N_3934,N_2386,N_2845);
or U3935 (N_3935,N_2332,N_2106);
or U3936 (N_3936,N_2448,N_2675);
nor U3937 (N_3937,N_2402,N_2166);
nand U3938 (N_3938,N_2914,N_2562);
nand U3939 (N_3939,N_2601,N_2912);
nand U3940 (N_3940,N_2984,N_2421);
or U3941 (N_3941,N_2149,N_2729);
or U3942 (N_3942,N_2976,N_2494);
xor U3943 (N_3943,N_2111,N_2353);
xnor U3944 (N_3944,N_2102,N_2638);
xor U3945 (N_3945,N_2872,N_2806);
or U3946 (N_3946,N_2705,N_2695);
and U3947 (N_3947,N_2681,N_2303);
nor U3948 (N_3948,N_2999,N_2733);
xnor U3949 (N_3949,N_2981,N_2569);
and U3950 (N_3950,N_2820,N_2467);
and U3951 (N_3951,N_2058,N_2722);
and U3952 (N_3952,N_2693,N_2618);
nor U3953 (N_3953,N_2133,N_2955);
xor U3954 (N_3954,N_2863,N_2094);
nor U3955 (N_3955,N_2063,N_2584);
or U3956 (N_3956,N_2308,N_2175);
or U3957 (N_3957,N_2229,N_2017);
and U3958 (N_3958,N_2772,N_2036);
or U3959 (N_3959,N_2197,N_2368);
nand U3960 (N_3960,N_2684,N_2762);
and U3961 (N_3961,N_2149,N_2889);
and U3962 (N_3962,N_2060,N_2541);
nor U3963 (N_3963,N_2745,N_2162);
and U3964 (N_3964,N_2008,N_2123);
and U3965 (N_3965,N_2712,N_2951);
nand U3966 (N_3966,N_2712,N_2918);
or U3967 (N_3967,N_2986,N_2521);
nor U3968 (N_3968,N_2464,N_2944);
and U3969 (N_3969,N_2143,N_2027);
or U3970 (N_3970,N_2314,N_2011);
nand U3971 (N_3971,N_2410,N_2342);
xnor U3972 (N_3972,N_2904,N_2500);
nor U3973 (N_3973,N_2919,N_2766);
and U3974 (N_3974,N_2572,N_2041);
xor U3975 (N_3975,N_2425,N_2798);
xnor U3976 (N_3976,N_2988,N_2417);
and U3977 (N_3977,N_2509,N_2337);
xor U3978 (N_3978,N_2766,N_2212);
and U3979 (N_3979,N_2043,N_2310);
nand U3980 (N_3980,N_2896,N_2088);
nand U3981 (N_3981,N_2595,N_2938);
and U3982 (N_3982,N_2089,N_2989);
xor U3983 (N_3983,N_2598,N_2911);
xnor U3984 (N_3984,N_2947,N_2332);
and U3985 (N_3985,N_2412,N_2932);
or U3986 (N_3986,N_2020,N_2245);
and U3987 (N_3987,N_2316,N_2433);
xor U3988 (N_3988,N_2724,N_2982);
and U3989 (N_3989,N_2442,N_2078);
nand U3990 (N_3990,N_2174,N_2533);
nor U3991 (N_3991,N_2072,N_2633);
xor U3992 (N_3992,N_2769,N_2464);
nand U3993 (N_3993,N_2577,N_2579);
nand U3994 (N_3994,N_2946,N_2714);
or U3995 (N_3995,N_2329,N_2764);
xnor U3996 (N_3996,N_2907,N_2892);
nor U3997 (N_3997,N_2004,N_2991);
and U3998 (N_3998,N_2150,N_2118);
xnor U3999 (N_3999,N_2042,N_2843);
nor U4000 (N_4000,N_3734,N_3726);
and U4001 (N_4001,N_3652,N_3105);
nor U4002 (N_4002,N_3352,N_3379);
xnor U4003 (N_4003,N_3749,N_3826);
nand U4004 (N_4004,N_3074,N_3954);
xnor U4005 (N_4005,N_3023,N_3697);
xor U4006 (N_4006,N_3350,N_3910);
or U4007 (N_4007,N_3143,N_3678);
xnor U4008 (N_4008,N_3134,N_3591);
nand U4009 (N_4009,N_3761,N_3084);
nor U4010 (N_4010,N_3784,N_3263);
xnor U4011 (N_4011,N_3363,N_3545);
nor U4012 (N_4012,N_3748,N_3767);
nand U4013 (N_4013,N_3716,N_3231);
and U4014 (N_4014,N_3326,N_3790);
or U4015 (N_4015,N_3179,N_3488);
nand U4016 (N_4016,N_3099,N_3013);
nor U4017 (N_4017,N_3290,N_3430);
nor U4018 (N_4018,N_3653,N_3088);
xor U4019 (N_4019,N_3832,N_3542);
xor U4020 (N_4020,N_3825,N_3329);
and U4021 (N_4021,N_3167,N_3119);
nor U4022 (N_4022,N_3950,N_3815);
nor U4023 (N_4023,N_3448,N_3838);
or U4024 (N_4024,N_3598,N_3333);
nor U4025 (N_4025,N_3746,N_3554);
and U4026 (N_4026,N_3229,N_3233);
nand U4027 (N_4027,N_3250,N_3853);
nand U4028 (N_4028,N_3934,N_3920);
xor U4029 (N_4029,N_3570,N_3972);
nor U4030 (N_4030,N_3559,N_3523);
xor U4031 (N_4031,N_3687,N_3961);
nor U4032 (N_4032,N_3087,N_3345);
nor U4033 (N_4033,N_3650,N_3235);
nor U4034 (N_4034,N_3303,N_3993);
or U4035 (N_4035,N_3863,N_3899);
xor U4036 (N_4036,N_3492,N_3422);
nor U4037 (N_4037,N_3358,N_3258);
nand U4038 (N_4038,N_3247,N_3259);
and U4039 (N_4039,N_3799,N_3061);
nor U4040 (N_4040,N_3412,N_3260);
nor U4041 (N_4041,N_3288,N_3765);
nand U4042 (N_4042,N_3080,N_3228);
xor U4043 (N_4043,N_3314,N_3571);
nor U4044 (N_4044,N_3042,N_3720);
and U4045 (N_4045,N_3403,N_3774);
and U4046 (N_4046,N_3880,N_3752);
xor U4047 (N_4047,N_3710,N_3184);
nor U4048 (N_4048,N_3103,N_3789);
and U4049 (N_4049,N_3963,N_3548);
nand U4050 (N_4050,N_3613,N_3661);
or U4051 (N_4051,N_3091,N_3140);
nand U4052 (N_4052,N_3969,N_3063);
or U4053 (N_4053,N_3249,N_3419);
or U4054 (N_4054,N_3193,N_3246);
xor U4055 (N_4055,N_3616,N_3460);
xor U4056 (N_4056,N_3271,N_3700);
nor U4057 (N_4057,N_3067,N_3036);
or U4058 (N_4058,N_3465,N_3861);
or U4059 (N_4059,N_3267,N_3704);
nor U4060 (N_4060,N_3619,N_3321);
or U4061 (N_4061,N_3956,N_3865);
xnor U4062 (N_4062,N_3445,N_3311);
nor U4063 (N_4063,N_3668,N_3810);
and U4064 (N_4064,N_3402,N_3762);
or U4065 (N_4065,N_3791,N_3092);
or U4066 (N_4066,N_3718,N_3577);
or U4067 (N_4067,N_3395,N_3755);
nand U4068 (N_4068,N_3451,N_3129);
or U4069 (N_4069,N_3398,N_3138);
and U4070 (N_4070,N_3908,N_3918);
or U4071 (N_4071,N_3497,N_3112);
nor U4072 (N_4072,N_3164,N_3751);
or U4073 (N_4073,N_3924,N_3513);
xnor U4074 (N_4074,N_3776,N_3521);
nor U4075 (N_4075,N_3557,N_3933);
nand U4076 (N_4076,N_3592,N_3868);
and U4077 (N_4077,N_3636,N_3928);
and U4078 (N_4078,N_3121,N_3086);
nor U4079 (N_4079,N_3538,N_3778);
and U4080 (N_4080,N_3420,N_3888);
nor U4081 (N_4081,N_3461,N_3628);
or U4082 (N_4082,N_3578,N_3053);
and U4083 (N_4083,N_3703,N_3962);
nand U4084 (N_4084,N_3917,N_3104);
and U4085 (N_4085,N_3931,N_3362);
nor U4086 (N_4086,N_3317,N_3527);
and U4087 (N_4087,N_3546,N_3889);
or U4088 (N_4088,N_3926,N_3381);
and U4089 (N_4089,N_3742,N_3261);
nand U4090 (N_4090,N_3560,N_3262);
or U4091 (N_4091,N_3045,N_3837);
nor U4092 (N_4092,N_3584,N_3443);
nor U4093 (N_4093,N_3551,N_3077);
or U4094 (N_4094,N_3268,N_3930);
nand U4095 (N_4095,N_3974,N_3425);
nor U4096 (N_4096,N_3029,N_3300);
and U4097 (N_4097,N_3606,N_3429);
or U4098 (N_4098,N_3894,N_3992);
and U4099 (N_4099,N_3265,N_3168);
or U4100 (N_4100,N_3620,N_3985);
nand U4101 (N_4101,N_3284,N_3328);
and U4102 (N_4102,N_3965,N_3226);
or U4103 (N_4103,N_3558,N_3048);
or U4104 (N_4104,N_3499,N_3209);
nor U4105 (N_4105,N_3565,N_3396);
nor U4106 (N_4106,N_3625,N_3895);
or U4107 (N_4107,N_3535,N_3866);
or U4108 (N_4108,N_3253,N_3622);
and U4109 (N_4109,N_3444,N_3191);
and U4110 (N_4110,N_3923,N_3713);
nor U4111 (N_4111,N_3058,N_3709);
xnor U4112 (N_4112,N_3970,N_3517);
or U4113 (N_4113,N_3941,N_3436);
nor U4114 (N_4114,N_3563,N_3222);
xor U4115 (N_4115,N_3296,N_3891);
or U4116 (N_4116,N_3310,N_3605);
nor U4117 (N_4117,N_3217,N_3686);
nor U4118 (N_4118,N_3039,N_3905);
nor U4119 (N_4119,N_3122,N_3407);
and U4120 (N_4120,N_3561,N_3618);
and U4121 (N_4121,N_3166,N_3475);
and U4122 (N_4122,N_3236,N_3427);
nor U4123 (N_4123,N_3732,N_3814);
and U4124 (N_4124,N_3032,N_3758);
nor U4125 (N_4125,N_3051,N_3449);
and U4126 (N_4126,N_3839,N_3325);
xnor U4127 (N_4127,N_3025,N_3681);
and U4128 (N_4128,N_3146,N_3293);
and U4129 (N_4129,N_3254,N_3501);
xnor U4130 (N_4130,N_3163,N_3977);
nor U4131 (N_4131,N_3135,N_3907);
or U4132 (N_4132,N_3028,N_3816);
nand U4133 (N_4133,N_3632,N_3079);
nor U4134 (N_4134,N_3877,N_3198);
nand U4135 (N_4135,N_3936,N_3364);
or U4136 (N_4136,N_3733,N_3286);
xor U4137 (N_4137,N_3024,N_3034);
nor U4138 (N_4138,N_3056,N_3990);
nand U4139 (N_4139,N_3937,N_3353);
nor U4140 (N_4140,N_3149,N_3520);
nor U4141 (N_4141,N_3308,N_3817);
and U4142 (N_4142,N_3484,N_3116);
nor U4143 (N_4143,N_3351,N_3553);
nand U4144 (N_4144,N_3848,N_3400);
xnor U4145 (N_4145,N_3737,N_3008);
and U4146 (N_4146,N_3912,N_3083);
xnor U4147 (N_4147,N_3289,N_3438);
nand U4148 (N_4148,N_3070,N_3071);
xor U4149 (N_4149,N_3169,N_3922);
or U4150 (N_4150,N_3902,N_3648);
nor U4151 (N_4151,N_3213,N_3638);
or U4152 (N_4152,N_3374,N_3630);
and U4153 (N_4153,N_3833,N_3531);
xor U4154 (N_4154,N_3844,N_3187);
or U4155 (N_4155,N_3512,N_3676);
and U4156 (N_4156,N_3579,N_3684);
xor U4157 (N_4157,N_3879,N_3552);
or U4158 (N_4158,N_3415,N_3344);
xor U4159 (N_4159,N_3323,N_3875);
xnor U4160 (N_4160,N_3723,N_3524);
xnor U4161 (N_4161,N_3275,N_3525);
nor U4162 (N_4162,N_3324,N_3884);
or U4163 (N_4163,N_3354,N_3137);
xnor U4164 (N_4164,N_3157,N_3892);
nor U4165 (N_4165,N_3347,N_3141);
xor U4166 (N_4166,N_3971,N_3585);
or U4167 (N_4167,N_3629,N_3901);
and U4168 (N_4168,N_3496,N_3366);
or U4169 (N_4169,N_3470,N_3530);
nor U4170 (N_4170,N_3820,N_3821);
nand U4171 (N_4171,N_3020,N_3463);
and U4172 (N_4172,N_3780,N_3312);
nand U4173 (N_4173,N_3022,N_3887);
nand U4174 (N_4174,N_3779,N_3212);
and U4175 (N_4175,N_3583,N_3124);
and U4176 (N_4176,N_3408,N_3054);
xor U4177 (N_4177,N_3979,N_3624);
or U4178 (N_4178,N_3355,N_3234);
or U4179 (N_4179,N_3110,N_3389);
nand U4180 (N_4180,N_3251,N_3480);
nor U4181 (N_4181,N_3478,N_3867);
or U4182 (N_4182,N_3454,N_3197);
nand U4183 (N_4183,N_3243,N_3428);
and U4184 (N_4184,N_3299,N_3763);
and U4185 (N_4185,N_3691,N_3801);
or U4186 (N_4186,N_3988,N_3126);
nor U4187 (N_4187,N_3117,N_3671);
and U4188 (N_4188,N_3831,N_3515);
nor U4189 (N_4189,N_3727,N_3128);
xnor U4190 (N_4190,N_3757,N_3044);
or U4191 (N_4191,N_3824,N_3062);
nor U4192 (N_4192,N_3014,N_3432);
or U4193 (N_4193,N_3370,N_3404);
and U4194 (N_4194,N_3830,N_3781);
nand U4195 (N_4195,N_3634,N_3647);
xnor U4196 (N_4196,N_3015,N_3665);
nor U4197 (N_4197,N_3159,N_3696);
nor U4198 (N_4198,N_3456,N_3847);
nor U4199 (N_4199,N_3683,N_3494);
nor U4200 (N_4200,N_3599,N_3967);
or U4201 (N_4201,N_3330,N_3335);
xnor U4202 (N_4202,N_3037,N_3139);
and U4203 (N_4203,N_3132,N_3596);
nor U4204 (N_4204,N_3946,N_3411);
or U4205 (N_4205,N_3431,N_3190);
and U4206 (N_4206,N_3828,N_3911);
nor U4207 (N_4207,N_3998,N_3747);
nor U4208 (N_4208,N_3667,N_3274);
nand U4209 (N_4209,N_3012,N_3199);
nand U4210 (N_4210,N_3241,N_3383);
xor U4211 (N_4211,N_3909,N_3893);
nand U4212 (N_4212,N_3855,N_3802);
nor U4213 (N_4213,N_3369,N_3773);
nor U4214 (N_4214,N_3211,N_3473);
or U4215 (N_4215,N_3097,N_3534);
nor U4216 (N_4216,N_3320,N_3481);
nor U4217 (N_4217,N_3148,N_3813);
nor U4218 (N_4218,N_3509,N_3007);
or U4219 (N_4219,N_3597,N_3073);
nor U4220 (N_4220,N_3675,N_3479);
nand U4221 (N_4221,N_3978,N_3796);
and U4222 (N_4222,N_3822,N_3204);
xor U4223 (N_4223,N_3698,N_3966);
xnor U4224 (N_4224,N_3147,N_3230);
and U4225 (N_4225,N_3659,N_3567);
nand U4226 (N_4226,N_3232,N_3556);
nor U4227 (N_4227,N_3872,N_3170);
nand U4228 (N_4228,N_3123,N_3336);
xor U4229 (N_4229,N_3614,N_3215);
and U4230 (N_4230,N_3502,N_3279);
nand U4231 (N_4231,N_3359,N_3850);
and U4232 (N_4232,N_3223,N_3171);
nand U4233 (N_4233,N_3717,N_3544);
or U4234 (N_4234,N_3298,N_3414);
nor U4235 (N_4235,N_3797,N_3541);
and U4236 (N_4236,N_3322,N_3437);
xor U4237 (N_4237,N_3981,N_3176);
nor U4238 (N_4238,N_3655,N_3455);
or U4239 (N_4239,N_3754,N_3468);
xor U4240 (N_4240,N_3756,N_3196);
nor U4241 (N_4241,N_3679,N_3098);
nor U4242 (N_4242,N_3670,N_3471);
and U4243 (N_4243,N_3151,N_3150);
nand U4244 (N_4244,N_3631,N_3959);
or U4245 (N_4245,N_3107,N_3741);
or U4246 (N_4246,N_3804,N_3027);
xor U4247 (N_4247,N_3674,N_3185);
and U4248 (N_4248,N_3935,N_3873);
and U4249 (N_4249,N_3342,N_3851);
xor U4250 (N_4250,N_3547,N_3607);
or U4251 (N_4251,N_3294,N_3252);
xnor U4252 (N_4252,N_3118,N_3133);
or U4253 (N_4253,N_3069,N_3845);
and U4254 (N_4254,N_3886,N_3794);
nand U4255 (N_4255,N_3782,N_3127);
and U4256 (N_4256,N_3929,N_3722);
nor U4257 (N_4257,N_3050,N_3368);
and U4258 (N_4258,N_3216,N_3949);
nor U4259 (N_4259,N_3611,N_3372);
nand U4260 (N_4260,N_3808,N_3082);
nor U4261 (N_4261,N_3540,N_3770);
nor U4262 (N_4262,N_3297,N_3573);
xor U4263 (N_4263,N_3812,N_3108);
nor U4264 (N_4264,N_3562,N_3273);
xnor U4265 (N_4265,N_3142,N_3278);
xor U4266 (N_4266,N_3218,N_3040);
or U4267 (N_4267,N_3656,N_3391);
xnor U4268 (N_4268,N_3490,N_3604);
nand U4269 (N_4269,N_3052,N_3952);
or U4270 (N_4270,N_3388,N_3493);
nand U4271 (N_4271,N_3242,N_3764);
nor U4272 (N_4272,N_3750,N_3595);
and U4273 (N_4273,N_3633,N_3919);
nand U4274 (N_4274,N_3162,N_3951);
and U4275 (N_4275,N_3771,N_3192);
xor U4276 (N_4276,N_3503,N_3532);
nand U4277 (N_4277,N_3405,N_3367);
nor U4278 (N_4278,N_3663,N_3030);
xor U4279 (N_4279,N_3154,N_3386);
nand U4280 (N_4280,N_3536,N_3476);
nand U4281 (N_4281,N_3702,N_3440);
nand U4282 (N_4282,N_3417,N_3009);
xor U4283 (N_4283,N_3640,N_3315);
xor U4284 (N_4284,N_3462,N_3421);
nor U4285 (N_4285,N_3180,N_3113);
nor U4286 (N_4286,N_3095,N_3982);
nor U4287 (N_4287,N_3453,N_3001);
and U4288 (N_4288,N_3487,N_3593);
and U4289 (N_4289,N_3011,N_3753);
and U4290 (N_4290,N_3257,N_3819);
xor U4291 (N_4291,N_3221,N_3806);
or U4292 (N_4292,N_3302,N_3201);
and U4293 (N_4293,N_3459,N_3021);
nor U4294 (N_4294,N_3626,N_3057);
or U4295 (N_4295,N_3621,N_3610);
nand U4296 (N_4296,N_3188,N_3735);
xnor U4297 (N_4297,N_3055,N_3307);
xnor U4298 (N_4298,N_3885,N_3569);
nor U4299 (N_4299,N_3182,N_3955);
or U4300 (N_4300,N_3474,N_3183);
nand U4301 (N_4301,N_3944,N_3669);
and U4302 (N_4302,N_3859,N_3466);
nor U4303 (N_4303,N_3401,N_3266);
or U4304 (N_4304,N_3006,N_3270);
and U4305 (N_4305,N_3313,N_3106);
and U4306 (N_4306,N_3537,N_3356);
xnor U4307 (N_4307,N_3576,N_3846);
or U4308 (N_4308,N_3608,N_3694);
nand U4309 (N_4309,N_3768,N_3526);
nor U4310 (N_4310,N_3393,N_3081);
and U4311 (N_4311,N_3996,N_3504);
or U4312 (N_4312,N_3047,N_3662);
and U4313 (N_4313,N_3072,N_3334);
nor U4314 (N_4314,N_3373,N_3729);
nand U4315 (N_4315,N_3019,N_3130);
nor U4316 (N_4316,N_3983,N_3076);
nand U4317 (N_4317,N_3786,N_3840);
nor U4318 (N_4318,N_3158,N_3377);
nor U4319 (N_4319,N_3360,N_3093);
xor U4320 (N_4320,N_3177,N_3682);
and U4321 (N_4321,N_3738,N_3469);
or U4322 (N_4322,N_3477,N_3600);
or U4323 (N_4323,N_3413,N_3602);
nor U4324 (N_4324,N_3685,N_3482);
and U4325 (N_4325,N_3100,N_3409);
nand U4326 (N_4326,N_3382,N_3125);
nand U4327 (N_4327,N_3916,N_3214);
or U4328 (N_4328,N_3575,N_3987);
nor U4329 (N_4329,N_3059,N_3915);
and U4330 (N_4330,N_3361,N_3574);
or U4331 (N_4331,N_3940,N_3999);
nand U4332 (N_4332,N_3304,N_3740);
or U4333 (N_4333,N_3380,N_3617);
nand U4334 (N_4334,N_3433,N_3500);
nand U4335 (N_4335,N_3639,N_3277);
nand U4336 (N_4336,N_3658,N_3707);
xnor U4337 (N_4337,N_3305,N_3017);
xnor U4338 (N_4338,N_3498,N_3219);
xnor U4339 (N_4339,N_3787,N_3564);
xnor U4340 (N_4340,N_3085,N_3173);
nor U4341 (N_4341,N_3060,N_3793);
xor U4342 (N_4342,N_3339,N_3309);
xnor U4343 (N_4343,N_3724,N_3491);
nand U4344 (N_4344,N_3064,N_3018);
xor U4345 (N_4345,N_3695,N_3739);
and U4346 (N_4346,N_3385,N_3896);
xor U4347 (N_4347,N_3483,N_3882);
xnor U4348 (N_4348,N_3510,N_3280);
nand U4349 (N_4349,N_3870,N_3446);
nand U4350 (N_4350,N_3094,N_3096);
nand U4351 (N_4351,N_3349,N_3829);
or U4352 (N_4352,N_3220,N_3701);
or U4353 (N_4353,N_3964,N_3410);
xnor U4354 (N_4354,N_3664,N_3172);
nor U4355 (N_4355,N_3458,N_3705);
nand U4356 (N_4356,N_3033,N_3225);
nor U4357 (N_4357,N_3533,N_3900);
nand U4358 (N_4358,N_3890,N_3208);
or U4359 (N_4359,N_3672,N_3818);
nor U4360 (N_4360,N_3111,N_3871);
xnor U4361 (N_4361,N_3874,N_3807);
nand U4362 (N_4362,N_3588,N_3316);
nand U4363 (N_4363,N_3506,N_3272);
nand U4364 (N_4364,N_3205,N_3078);
nand U4365 (N_4365,N_3953,N_3472);
nand U4366 (N_4366,N_3282,N_3376);
xor U4367 (N_4367,N_3643,N_3623);
and U4368 (N_4368,N_3237,N_3785);
nor U4369 (N_4369,N_3939,N_3276);
or U4370 (N_4370,N_3348,N_3744);
xnor U4371 (N_4371,N_3635,N_3397);
and U4372 (N_4372,N_3340,N_3745);
and U4373 (N_4373,N_3712,N_3856);
and U4374 (N_4374,N_3809,N_3109);
nand U4375 (N_4375,N_3156,N_3114);
nor U4376 (N_4376,N_3423,N_3522);
or U4377 (N_4377,N_3589,N_3450);
or U4378 (N_4378,N_3186,N_3357);
and U4379 (N_4379,N_3772,N_3153);
or U4380 (N_4380,N_3485,N_3646);
nor U4381 (N_4381,N_3898,N_3792);
nor U4382 (N_4382,N_3580,N_3841);
nand U4383 (N_4383,N_3467,N_3673);
nand U4384 (N_4384,N_3046,N_3906);
nor U4385 (N_4385,N_3677,N_3914);
xnor U4386 (N_4386,N_3160,N_3392);
xnor U4387 (N_4387,N_3043,N_3207);
nand U4388 (N_4388,N_3654,N_3508);
and U4389 (N_4389,N_3144,N_3255);
or U4390 (N_4390,N_3507,N_3035);
nand U4391 (N_4391,N_3943,N_3759);
and U4392 (N_4392,N_3292,N_3692);
xor U4393 (N_4393,N_3715,N_3306);
or U4394 (N_4394,N_3439,N_3447);
nand U4395 (N_4395,N_3003,N_3876);
or U4396 (N_4396,N_3452,N_3615);
nand U4397 (N_4397,N_3031,N_3783);
nand U4398 (N_4398,N_3418,N_3945);
or U4399 (N_4399,N_3337,N_3948);
nand U4400 (N_4400,N_3331,N_3178);
nand U4401 (N_4401,N_3991,N_3457);
nor U4402 (N_4402,N_3644,N_3957);
xnor U4403 (N_4403,N_3155,N_3248);
xor U4404 (N_4404,N_3161,N_3174);
nand U4405 (N_4405,N_3719,N_3775);
or U4406 (N_4406,N_3849,N_3000);
or U4407 (N_4407,N_3224,N_3601);
or U4408 (N_4408,N_3878,N_3341);
and U4409 (N_4409,N_3346,N_3986);
nand U4410 (N_4410,N_3200,N_3582);
nor U4411 (N_4411,N_3424,N_3239);
nand U4412 (N_4412,N_3864,N_3827);
nor U4413 (N_4413,N_3511,N_3406);
nor U4414 (N_4414,N_3399,N_3989);
xnor U4415 (N_4415,N_3203,N_3441);
nor U4416 (N_4416,N_3175,N_3516);
xor U4417 (N_4417,N_3938,N_3811);
nor U4418 (N_4418,N_3769,N_3690);
and U4419 (N_4419,N_3927,N_3041);
nor U4420 (N_4420,N_3721,N_3195);
xnor U4421 (N_4421,N_3968,N_3416);
nand U4422 (N_4422,N_3711,N_3743);
nor U4423 (N_4423,N_3730,N_3038);
xor U4424 (N_4424,N_3529,N_3843);
nor U4425 (N_4425,N_3505,N_3903);
nand U4426 (N_4426,N_3295,N_3731);
and U4427 (N_4427,N_3852,N_3995);
nor U4428 (N_4428,N_3005,N_3823);
or U4429 (N_4429,N_3378,N_3435);
or U4430 (N_4430,N_3269,N_3555);
and U4431 (N_4431,N_3587,N_3390);
or U4432 (N_4432,N_3657,N_3464);
and U4433 (N_4433,N_3495,N_3365);
nor U4434 (N_4434,N_3777,N_3131);
xnor U4435 (N_4435,N_3202,N_3343);
nand U4436 (N_4436,N_3913,N_3115);
nor U4437 (N_4437,N_3835,N_3594);
or U4438 (N_4438,N_3002,N_3921);
and U4439 (N_4439,N_3736,N_3102);
nand U4440 (N_4440,N_3714,N_3026);
and U4441 (N_4441,N_3689,N_3068);
and U4442 (N_4442,N_3539,N_3514);
nor U4443 (N_4443,N_3860,N_3904);
and U4444 (N_4444,N_3836,N_3004);
xnor U4445 (N_4445,N_3728,N_3394);
or U4446 (N_4446,N_3291,N_3245);
nand U4447 (N_4447,N_3206,N_3760);
xnor U4448 (N_4448,N_3660,N_3612);
or U4449 (N_4449,N_3375,N_3609);
xnor U4450 (N_4450,N_3881,N_3858);
or U4451 (N_4451,N_3994,N_3680);
or U4452 (N_4452,N_3800,N_3332);
xor U4453 (N_4453,N_3238,N_3136);
xor U4454 (N_4454,N_3645,N_3975);
xnor U4455 (N_4455,N_3066,N_3442);
xor U4456 (N_4456,N_3932,N_3590);
and U4457 (N_4457,N_3572,N_3264);
and U4458 (N_4458,N_3287,N_3240);
xnor U4459 (N_4459,N_3942,N_3549);
xnor U4460 (N_4460,N_3181,N_3642);
nor U4461 (N_4461,N_3795,N_3869);
or U4462 (N_4462,N_3854,N_3285);
xor U4463 (N_4463,N_3947,N_3958);
and U4464 (N_4464,N_3489,N_3244);
xnor U4465 (N_4465,N_3997,N_3519);
and U4466 (N_4466,N_3834,N_3883);
xor U4467 (N_4467,N_3566,N_3194);
nor U4468 (N_4468,N_3486,N_3803);
nand U4469 (N_4469,N_3842,N_3227);
xor U4470 (N_4470,N_3010,N_3805);
and U4471 (N_4471,N_3976,N_3387);
nor U4472 (N_4472,N_3649,N_3075);
nor U4473 (N_4473,N_3798,N_3973);
or U4474 (N_4474,N_3766,N_3603);
nor U4475 (N_4475,N_3708,N_3550);
or U4476 (N_4476,N_3788,N_3384);
nand U4477 (N_4477,N_3543,N_3101);
and U4478 (N_4478,N_3699,N_3528);
nor U4479 (N_4479,N_3145,N_3090);
or U4480 (N_4480,N_3301,N_3518);
nand U4481 (N_4481,N_3706,N_3862);
nor U4482 (N_4482,N_3256,N_3434);
nand U4483 (N_4483,N_3581,N_3980);
or U4484 (N_4484,N_3641,N_3651);
nand U4485 (N_4485,N_3857,N_3586);
nor U4486 (N_4486,N_3318,N_3897);
and U4487 (N_4487,N_3189,N_3984);
and U4488 (N_4488,N_3688,N_3960);
nand U4489 (N_4489,N_3049,N_3693);
xnor U4490 (N_4490,N_3281,N_3120);
and U4491 (N_4491,N_3283,N_3725);
or U4492 (N_4492,N_3089,N_3568);
nor U4493 (N_4493,N_3338,N_3165);
nand U4494 (N_4494,N_3016,N_3327);
and U4495 (N_4495,N_3152,N_3371);
nand U4496 (N_4496,N_3637,N_3065);
xnor U4497 (N_4497,N_3319,N_3925);
xnor U4498 (N_4498,N_3627,N_3210);
xnor U4499 (N_4499,N_3666,N_3426);
or U4500 (N_4500,N_3090,N_3209);
or U4501 (N_4501,N_3459,N_3173);
and U4502 (N_4502,N_3359,N_3283);
and U4503 (N_4503,N_3767,N_3849);
or U4504 (N_4504,N_3051,N_3079);
nor U4505 (N_4505,N_3357,N_3168);
and U4506 (N_4506,N_3118,N_3780);
xnor U4507 (N_4507,N_3822,N_3400);
nand U4508 (N_4508,N_3525,N_3208);
nor U4509 (N_4509,N_3532,N_3263);
nor U4510 (N_4510,N_3417,N_3040);
nand U4511 (N_4511,N_3905,N_3066);
nor U4512 (N_4512,N_3025,N_3552);
and U4513 (N_4513,N_3625,N_3060);
nand U4514 (N_4514,N_3679,N_3803);
nand U4515 (N_4515,N_3567,N_3205);
and U4516 (N_4516,N_3968,N_3084);
xor U4517 (N_4517,N_3192,N_3298);
nor U4518 (N_4518,N_3698,N_3334);
and U4519 (N_4519,N_3351,N_3115);
nand U4520 (N_4520,N_3392,N_3293);
xnor U4521 (N_4521,N_3536,N_3884);
xor U4522 (N_4522,N_3846,N_3175);
nand U4523 (N_4523,N_3849,N_3721);
and U4524 (N_4524,N_3670,N_3637);
nand U4525 (N_4525,N_3609,N_3768);
nand U4526 (N_4526,N_3035,N_3957);
and U4527 (N_4527,N_3500,N_3654);
xnor U4528 (N_4528,N_3612,N_3977);
xnor U4529 (N_4529,N_3126,N_3880);
nor U4530 (N_4530,N_3854,N_3257);
and U4531 (N_4531,N_3723,N_3266);
xor U4532 (N_4532,N_3229,N_3953);
or U4533 (N_4533,N_3029,N_3547);
nor U4534 (N_4534,N_3603,N_3849);
and U4535 (N_4535,N_3639,N_3275);
nor U4536 (N_4536,N_3517,N_3885);
nand U4537 (N_4537,N_3767,N_3910);
nand U4538 (N_4538,N_3869,N_3883);
or U4539 (N_4539,N_3465,N_3818);
xor U4540 (N_4540,N_3268,N_3551);
xnor U4541 (N_4541,N_3649,N_3982);
and U4542 (N_4542,N_3384,N_3990);
or U4543 (N_4543,N_3405,N_3951);
nand U4544 (N_4544,N_3671,N_3156);
or U4545 (N_4545,N_3233,N_3413);
and U4546 (N_4546,N_3995,N_3344);
or U4547 (N_4547,N_3484,N_3247);
and U4548 (N_4548,N_3507,N_3232);
or U4549 (N_4549,N_3219,N_3105);
and U4550 (N_4550,N_3050,N_3643);
nand U4551 (N_4551,N_3021,N_3210);
nand U4552 (N_4552,N_3351,N_3354);
and U4553 (N_4553,N_3537,N_3778);
nor U4554 (N_4554,N_3376,N_3116);
nor U4555 (N_4555,N_3195,N_3819);
or U4556 (N_4556,N_3170,N_3859);
nand U4557 (N_4557,N_3074,N_3111);
nand U4558 (N_4558,N_3481,N_3982);
xor U4559 (N_4559,N_3592,N_3655);
xnor U4560 (N_4560,N_3587,N_3105);
nor U4561 (N_4561,N_3657,N_3214);
nand U4562 (N_4562,N_3134,N_3513);
nand U4563 (N_4563,N_3256,N_3898);
nor U4564 (N_4564,N_3280,N_3735);
xnor U4565 (N_4565,N_3663,N_3100);
xor U4566 (N_4566,N_3589,N_3733);
nor U4567 (N_4567,N_3093,N_3464);
or U4568 (N_4568,N_3927,N_3937);
nand U4569 (N_4569,N_3927,N_3200);
nand U4570 (N_4570,N_3592,N_3792);
nor U4571 (N_4571,N_3732,N_3900);
and U4572 (N_4572,N_3686,N_3925);
xnor U4573 (N_4573,N_3139,N_3195);
nand U4574 (N_4574,N_3478,N_3497);
nand U4575 (N_4575,N_3746,N_3505);
nand U4576 (N_4576,N_3787,N_3637);
xnor U4577 (N_4577,N_3125,N_3594);
and U4578 (N_4578,N_3881,N_3735);
nor U4579 (N_4579,N_3609,N_3870);
and U4580 (N_4580,N_3742,N_3917);
nand U4581 (N_4581,N_3373,N_3519);
and U4582 (N_4582,N_3096,N_3255);
or U4583 (N_4583,N_3147,N_3525);
nor U4584 (N_4584,N_3442,N_3256);
xnor U4585 (N_4585,N_3663,N_3486);
or U4586 (N_4586,N_3346,N_3041);
or U4587 (N_4587,N_3169,N_3438);
or U4588 (N_4588,N_3666,N_3773);
and U4589 (N_4589,N_3102,N_3061);
and U4590 (N_4590,N_3035,N_3217);
nand U4591 (N_4591,N_3272,N_3698);
or U4592 (N_4592,N_3788,N_3754);
and U4593 (N_4593,N_3992,N_3630);
or U4594 (N_4594,N_3585,N_3505);
nor U4595 (N_4595,N_3923,N_3944);
nor U4596 (N_4596,N_3784,N_3544);
nor U4597 (N_4597,N_3673,N_3962);
nand U4598 (N_4598,N_3140,N_3249);
nor U4599 (N_4599,N_3623,N_3286);
and U4600 (N_4600,N_3013,N_3194);
nand U4601 (N_4601,N_3846,N_3116);
nand U4602 (N_4602,N_3959,N_3949);
nand U4603 (N_4603,N_3127,N_3537);
nand U4604 (N_4604,N_3032,N_3932);
xnor U4605 (N_4605,N_3254,N_3550);
and U4606 (N_4606,N_3284,N_3746);
xor U4607 (N_4607,N_3130,N_3037);
nand U4608 (N_4608,N_3070,N_3254);
xor U4609 (N_4609,N_3049,N_3721);
xor U4610 (N_4610,N_3898,N_3042);
or U4611 (N_4611,N_3557,N_3210);
nand U4612 (N_4612,N_3108,N_3366);
nand U4613 (N_4613,N_3195,N_3987);
xnor U4614 (N_4614,N_3470,N_3757);
nand U4615 (N_4615,N_3436,N_3240);
and U4616 (N_4616,N_3153,N_3690);
nor U4617 (N_4617,N_3932,N_3750);
xnor U4618 (N_4618,N_3954,N_3764);
nand U4619 (N_4619,N_3602,N_3379);
xnor U4620 (N_4620,N_3917,N_3850);
nor U4621 (N_4621,N_3166,N_3285);
or U4622 (N_4622,N_3964,N_3012);
or U4623 (N_4623,N_3230,N_3222);
and U4624 (N_4624,N_3848,N_3617);
xnor U4625 (N_4625,N_3159,N_3782);
nand U4626 (N_4626,N_3332,N_3183);
nor U4627 (N_4627,N_3283,N_3353);
and U4628 (N_4628,N_3153,N_3733);
or U4629 (N_4629,N_3769,N_3681);
or U4630 (N_4630,N_3312,N_3431);
xnor U4631 (N_4631,N_3232,N_3317);
nand U4632 (N_4632,N_3010,N_3521);
nor U4633 (N_4633,N_3527,N_3520);
xnor U4634 (N_4634,N_3918,N_3033);
nor U4635 (N_4635,N_3899,N_3469);
and U4636 (N_4636,N_3556,N_3842);
or U4637 (N_4637,N_3022,N_3029);
nor U4638 (N_4638,N_3254,N_3829);
xor U4639 (N_4639,N_3153,N_3835);
nor U4640 (N_4640,N_3018,N_3444);
or U4641 (N_4641,N_3506,N_3061);
nor U4642 (N_4642,N_3569,N_3203);
or U4643 (N_4643,N_3613,N_3337);
or U4644 (N_4644,N_3016,N_3213);
xnor U4645 (N_4645,N_3645,N_3222);
xnor U4646 (N_4646,N_3218,N_3368);
and U4647 (N_4647,N_3326,N_3926);
xnor U4648 (N_4648,N_3808,N_3016);
nor U4649 (N_4649,N_3929,N_3496);
nand U4650 (N_4650,N_3242,N_3228);
or U4651 (N_4651,N_3335,N_3538);
nor U4652 (N_4652,N_3570,N_3199);
nor U4653 (N_4653,N_3948,N_3914);
nand U4654 (N_4654,N_3053,N_3791);
and U4655 (N_4655,N_3422,N_3174);
nand U4656 (N_4656,N_3581,N_3634);
or U4657 (N_4657,N_3577,N_3752);
or U4658 (N_4658,N_3823,N_3729);
xor U4659 (N_4659,N_3938,N_3097);
nor U4660 (N_4660,N_3437,N_3716);
nand U4661 (N_4661,N_3103,N_3524);
or U4662 (N_4662,N_3245,N_3049);
and U4663 (N_4663,N_3308,N_3278);
xor U4664 (N_4664,N_3644,N_3280);
nand U4665 (N_4665,N_3072,N_3157);
nor U4666 (N_4666,N_3741,N_3878);
or U4667 (N_4667,N_3657,N_3277);
and U4668 (N_4668,N_3963,N_3270);
nor U4669 (N_4669,N_3620,N_3763);
or U4670 (N_4670,N_3690,N_3986);
or U4671 (N_4671,N_3891,N_3574);
or U4672 (N_4672,N_3261,N_3854);
and U4673 (N_4673,N_3585,N_3447);
and U4674 (N_4674,N_3155,N_3870);
or U4675 (N_4675,N_3743,N_3953);
nor U4676 (N_4676,N_3340,N_3820);
xnor U4677 (N_4677,N_3366,N_3109);
nor U4678 (N_4678,N_3027,N_3674);
and U4679 (N_4679,N_3357,N_3521);
and U4680 (N_4680,N_3671,N_3840);
or U4681 (N_4681,N_3286,N_3284);
and U4682 (N_4682,N_3383,N_3457);
xor U4683 (N_4683,N_3501,N_3512);
nor U4684 (N_4684,N_3492,N_3412);
nand U4685 (N_4685,N_3320,N_3027);
nand U4686 (N_4686,N_3466,N_3702);
and U4687 (N_4687,N_3447,N_3697);
or U4688 (N_4688,N_3138,N_3308);
or U4689 (N_4689,N_3401,N_3319);
and U4690 (N_4690,N_3857,N_3686);
and U4691 (N_4691,N_3454,N_3192);
and U4692 (N_4692,N_3936,N_3658);
and U4693 (N_4693,N_3059,N_3375);
or U4694 (N_4694,N_3126,N_3949);
and U4695 (N_4695,N_3377,N_3154);
xnor U4696 (N_4696,N_3979,N_3557);
or U4697 (N_4697,N_3422,N_3340);
nand U4698 (N_4698,N_3857,N_3571);
nor U4699 (N_4699,N_3600,N_3559);
nand U4700 (N_4700,N_3475,N_3836);
and U4701 (N_4701,N_3887,N_3103);
and U4702 (N_4702,N_3007,N_3759);
nor U4703 (N_4703,N_3257,N_3182);
or U4704 (N_4704,N_3895,N_3428);
xnor U4705 (N_4705,N_3796,N_3673);
or U4706 (N_4706,N_3335,N_3080);
nor U4707 (N_4707,N_3042,N_3529);
xor U4708 (N_4708,N_3329,N_3323);
xnor U4709 (N_4709,N_3394,N_3710);
nor U4710 (N_4710,N_3305,N_3393);
or U4711 (N_4711,N_3477,N_3552);
and U4712 (N_4712,N_3575,N_3416);
nand U4713 (N_4713,N_3526,N_3689);
nand U4714 (N_4714,N_3496,N_3091);
and U4715 (N_4715,N_3251,N_3448);
and U4716 (N_4716,N_3261,N_3989);
nand U4717 (N_4717,N_3887,N_3402);
or U4718 (N_4718,N_3020,N_3625);
nor U4719 (N_4719,N_3004,N_3919);
and U4720 (N_4720,N_3062,N_3503);
nand U4721 (N_4721,N_3527,N_3319);
nand U4722 (N_4722,N_3900,N_3498);
nor U4723 (N_4723,N_3237,N_3540);
or U4724 (N_4724,N_3799,N_3749);
nor U4725 (N_4725,N_3201,N_3185);
nand U4726 (N_4726,N_3842,N_3629);
xnor U4727 (N_4727,N_3531,N_3635);
and U4728 (N_4728,N_3095,N_3733);
and U4729 (N_4729,N_3783,N_3352);
nor U4730 (N_4730,N_3056,N_3312);
or U4731 (N_4731,N_3175,N_3293);
or U4732 (N_4732,N_3172,N_3629);
and U4733 (N_4733,N_3595,N_3749);
nand U4734 (N_4734,N_3805,N_3743);
nor U4735 (N_4735,N_3654,N_3188);
nor U4736 (N_4736,N_3863,N_3408);
nand U4737 (N_4737,N_3914,N_3229);
nand U4738 (N_4738,N_3000,N_3731);
xnor U4739 (N_4739,N_3371,N_3657);
or U4740 (N_4740,N_3567,N_3675);
and U4741 (N_4741,N_3178,N_3674);
nor U4742 (N_4742,N_3057,N_3418);
xnor U4743 (N_4743,N_3998,N_3961);
or U4744 (N_4744,N_3091,N_3181);
nor U4745 (N_4745,N_3583,N_3827);
nand U4746 (N_4746,N_3806,N_3283);
nand U4747 (N_4747,N_3952,N_3656);
nor U4748 (N_4748,N_3584,N_3679);
nor U4749 (N_4749,N_3795,N_3623);
nor U4750 (N_4750,N_3182,N_3019);
nor U4751 (N_4751,N_3231,N_3489);
and U4752 (N_4752,N_3701,N_3491);
or U4753 (N_4753,N_3988,N_3331);
nand U4754 (N_4754,N_3872,N_3137);
and U4755 (N_4755,N_3243,N_3876);
nor U4756 (N_4756,N_3486,N_3044);
nor U4757 (N_4757,N_3819,N_3503);
and U4758 (N_4758,N_3436,N_3180);
or U4759 (N_4759,N_3079,N_3771);
or U4760 (N_4760,N_3272,N_3363);
and U4761 (N_4761,N_3622,N_3931);
nor U4762 (N_4762,N_3961,N_3299);
xnor U4763 (N_4763,N_3170,N_3951);
and U4764 (N_4764,N_3647,N_3472);
or U4765 (N_4765,N_3813,N_3940);
or U4766 (N_4766,N_3639,N_3839);
xor U4767 (N_4767,N_3142,N_3530);
or U4768 (N_4768,N_3978,N_3440);
nand U4769 (N_4769,N_3678,N_3234);
nand U4770 (N_4770,N_3626,N_3330);
nor U4771 (N_4771,N_3387,N_3342);
nor U4772 (N_4772,N_3029,N_3875);
nand U4773 (N_4773,N_3896,N_3841);
nand U4774 (N_4774,N_3575,N_3997);
xor U4775 (N_4775,N_3499,N_3032);
nand U4776 (N_4776,N_3283,N_3056);
or U4777 (N_4777,N_3570,N_3345);
nor U4778 (N_4778,N_3140,N_3104);
nor U4779 (N_4779,N_3988,N_3377);
nand U4780 (N_4780,N_3057,N_3264);
nor U4781 (N_4781,N_3716,N_3232);
or U4782 (N_4782,N_3183,N_3560);
nand U4783 (N_4783,N_3325,N_3708);
and U4784 (N_4784,N_3948,N_3561);
or U4785 (N_4785,N_3584,N_3010);
or U4786 (N_4786,N_3340,N_3092);
nor U4787 (N_4787,N_3120,N_3111);
and U4788 (N_4788,N_3773,N_3892);
or U4789 (N_4789,N_3978,N_3118);
xnor U4790 (N_4790,N_3568,N_3985);
and U4791 (N_4791,N_3628,N_3222);
and U4792 (N_4792,N_3711,N_3502);
nor U4793 (N_4793,N_3728,N_3130);
nand U4794 (N_4794,N_3019,N_3889);
xor U4795 (N_4795,N_3072,N_3634);
and U4796 (N_4796,N_3695,N_3628);
or U4797 (N_4797,N_3786,N_3417);
xnor U4798 (N_4798,N_3733,N_3001);
nand U4799 (N_4799,N_3370,N_3895);
or U4800 (N_4800,N_3935,N_3024);
nand U4801 (N_4801,N_3406,N_3216);
nor U4802 (N_4802,N_3590,N_3318);
xnor U4803 (N_4803,N_3323,N_3463);
xnor U4804 (N_4804,N_3032,N_3074);
nor U4805 (N_4805,N_3744,N_3767);
nor U4806 (N_4806,N_3050,N_3031);
xnor U4807 (N_4807,N_3283,N_3832);
xnor U4808 (N_4808,N_3714,N_3737);
nand U4809 (N_4809,N_3235,N_3004);
and U4810 (N_4810,N_3160,N_3124);
xnor U4811 (N_4811,N_3712,N_3396);
or U4812 (N_4812,N_3029,N_3033);
nor U4813 (N_4813,N_3513,N_3256);
and U4814 (N_4814,N_3818,N_3222);
or U4815 (N_4815,N_3275,N_3522);
xnor U4816 (N_4816,N_3394,N_3037);
nand U4817 (N_4817,N_3064,N_3124);
xnor U4818 (N_4818,N_3663,N_3321);
or U4819 (N_4819,N_3278,N_3693);
or U4820 (N_4820,N_3077,N_3360);
nor U4821 (N_4821,N_3366,N_3648);
and U4822 (N_4822,N_3061,N_3597);
and U4823 (N_4823,N_3643,N_3206);
or U4824 (N_4824,N_3765,N_3849);
or U4825 (N_4825,N_3960,N_3656);
nor U4826 (N_4826,N_3115,N_3506);
xnor U4827 (N_4827,N_3498,N_3704);
and U4828 (N_4828,N_3204,N_3949);
xor U4829 (N_4829,N_3672,N_3340);
nand U4830 (N_4830,N_3710,N_3266);
xor U4831 (N_4831,N_3009,N_3819);
xnor U4832 (N_4832,N_3322,N_3308);
nor U4833 (N_4833,N_3654,N_3280);
or U4834 (N_4834,N_3434,N_3953);
or U4835 (N_4835,N_3336,N_3293);
or U4836 (N_4836,N_3469,N_3003);
xnor U4837 (N_4837,N_3751,N_3515);
nand U4838 (N_4838,N_3926,N_3814);
xnor U4839 (N_4839,N_3044,N_3599);
and U4840 (N_4840,N_3274,N_3717);
and U4841 (N_4841,N_3526,N_3248);
xor U4842 (N_4842,N_3605,N_3066);
xnor U4843 (N_4843,N_3046,N_3620);
nand U4844 (N_4844,N_3547,N_3667);
and U4845 (N_4845,N_3238,N_3019);
and U4846 (N_4846,N_3126,N_3438);
or U4847 (N_4847,N_3521,N_3972);
or U4848 (N_4848,N_3532,N_3195);
xnor U4849 (N_4849,N_3347,N_3123);
and U4850 (N_4850,N_3158,N_3468);
or U4851 (N_4851,N_3751,N_3396);
nor U4852 (N_4852,N_3325,N_3735);
or U4853 (N_4853,N_3917,N_3901);
nand U4854 (N_4854,N_3586,N_3131);
nor U4855 (N_4855,N_3284,N_3589);
nand U4856 (N_4856,N_3200,N_3208);
nor U4857 (N_4857,N_3160,N_3236);
xnor U4858 (N_4858,N_3031,N_3554);
nor U4859 (N_4859,N_3176,N_3549);
nand U4860 (N_4860,N_3518,N_3384);
and U4861 (N_4861,N_3029,N_3740);
xor U4862 (N_4862,N_3068,N_3952);
and U4863 (N_4863,N_3087,N_3655);
or U4864 (N_4864,N_3896,N_3628);
xnor U4865 (N_4865,N_3801,N_3203);
or U4866 (N_4866,N_3794,N_3091);
or U4867 (N_4867,N_3542,N_3662);
nor U4868 (N_4868,N_3627,N_3877);
nor U4869 (N_4869,N_3134,N_3092);
or U4870 (N_4870,N_3063,N_3179);
xnor U4871 (N_4871,N_3584,N_3864);
nor U4872 (N_4872,N_3028,N_3347);
and U4873 (N_4873,N_3608,N_3985);
or U4874 (N_4874,N_3118,N_3535);
and U4875 (N_4875,N_3113,N_3283);
or U4876 (N_4876,N_3768,N_3691);
or U4877 (N_4877,N_3727,N_3943);
nor U4878 (N_4878,N_3991,N_3004);
nand U4879 (N_4879,N_3189,N_3732);
and U4880 (N_4880,N_3340,N_3476);
nand U4881 (N_4881,N_3799,N_3442);
nor U4882 (N_4882,N_3913,N_3524);
and U4883 (N_4883,N_3031,N_3477);
or U4884 (N_4884,N_3158,N_3084);
or U4885 (N_4885,N_3804,N_3353);
or U4886 (N_4886,N_3771,N_3193);
xor U4887 (N_4887,N_3070,N_3800);
nor U4888 (N_4888,N_3112,N_3870);
and U4889 (N_4889,N_3513,N_3674);
nand U4890 (N_4890,N_3237,N_3843);
or U4891 (N_4891,N_3775,N_3526);
or U4892 (N_4892,N_3661,N_3336);
nand U4893 (N_4893,N_3295,N_3190);
xnor U4894 (N_4894,N_3333,N_3891);
or U4895 (N_4895,N_3753,N_3136);
and U4896 (N_4896,N_3803,N_3034);
nand U4897 (N_4897,N_3095,N_3470);
nor U4898 (N_4898,N_3501,N_3106);
nor U4899 (N_4899,N_3485,N_3374);
xor U4900 (N_4900,N_3217,N_3518);
and U4901 (N_4901,N_3615,N_3143);
nand U4902 (N_4902,N_3694,N_3159);
and U4903 (N_4903,N_3752,N_3993);
xor U4904 (N_4904,N_3629,N_3447);
nor U4905 (N_4905,N_3698,N_3417);
nor U4906 (N_4906,N_3109,N_3443);
nor U4907 (N_4907,N_3406,N_3004);
nor U4908 (N_4908,N_3151,N_3275);
xnor U4909 (N_4909,N_3450,N_3033);
or U4910 (N_4910,N_3664,N_3193);
or U4911 (N_4911,N_3303,N_3188);
or U4912 (N_4912,N_3402,N_3356);
nor U4913 (N_4913,N_3474,N_3318);
nand U4914 (N_4914,N_3613,N_3531);
or U4915 (N_4915,N_3695,N_3697);
and U4916 (N_4916,N_3002,N_3742);
or U4917 (N_4917,N_3414,N_3897);
nand U4918 (N_4918,N_3972,N_3670);
nand U4919 (N_4919,N_3265,N_3978);
xor U4920 (N_4920,N_3294,N_3457);
and U4921 (N_4921,N_3070,N_3857);
xor U4922 (N_4922,N_3392,N_3651);
or U4923 (N_4923,N_3333,N_3658);
and U4924 (N_4924,N_3521,N_3941);
and U4925 (N_4925,N_3059,N_3336);
xor U4926 (N_4926,N_3010,N_3854);
and U4927 (N_4927,N_3673,N_3142);
xnor U4928 (N_4928,N_3895,N_3877);
nand U4929 (N_4929,N_3723,N_3652);
and U4930 (N_4930,N_3122,N_3984);
nor U4931 (N_4931,N_3449,N_3472);
and U4932 (N_4932,N_3727,N_3151);
and U4933 (N_4933,N_3572,N_3341);
xnor U4934 (N_4934,N_3307,N_3634);
or U4935 (N_4935,N_3187,N_3900);
and U4936 (N_4936,N_3446,N_3375);
nand U4937 (N_4937,N_3328,N_3866);
nor U4938 (N_4938,N_3839,N_3890);
nand U4939 (N_4939,N_3969,N_3442);
nand U4940 (N_4940,N_3100,N_3565);
or U4941 (N_4941,N_3039,N_3127);
xor U4942 (N_4942,N_3277,N_3857);
nand U4943 (N_4943,N_3172,N_3353);
nor U4944 (N_4944,N_3697,N_3728);
and U4945 (N_4945,N_3212,N_3772);
xor U4946 (N_4946,N_3834,N_3142);
xnor U4947 (N_4947,N_3738,N_3319);
or U4948 (N_4948,N_3936,N_3419);
nor U4949 (N_4949,N_3447,N_3986);
nor U4950 (N_4950,N_3059,N_3936);
or U4951 (N_4951,N_3099,N_3247);
nor U4952 (N_4952,N_3234,N_3830);
nand U4953 (N_4953,N_3412,N_3875);
and U4954 (N_4954,N_3706,N_3251);
and U4955 (N_4955,N_3849,N_3267);
xor U4956 (N_4956,N_3459,N_3748);
or U4957 (N_4957,N_3464,N_3853);
and U4958 (N_4958,N_3249,N_3761);
nand U4959 (N_4959,N_3445,N_3018);
nor U4960 (N_4960,N_3471,N_3143);
xnor U4961 (N_4961,N_3483,N_3182);
and U4962 (N_4962,N_3224,N_3090);
xnor U4963 (N_4963,N_3402,N_3022);
or U4964 (N_4964,N_3365,N_3335);
xor U4965 (N_4965,N_3658,N_3830);
or U4966 (N_4966,N_3001,N_3833);
xnor U4967 (N_4967,N_3814,N_3856);
xnor U4968 (N_4968,N_3521,N_3328);
or U4969 (N_4969,N_3908,N_3513);
nor U4970 (N_4970,N_3219,N_3996);
nand U4971 (N_4971,N_3307,N_3138);
nor U4972 (N_4972,N_3388,N_3844);
nor U4973 (N_4973,N_3629,N_3678);
and U4974 (N_4974,N_3583,N_3649);
or U4975 (N_4975,N_3896,N_3745);
nand U4976 (N_4976,N_3794,N_3940);
or U4977 (N_4977,N_3715,N_3792);
and U4978 (N_4978,N_3618,N_3456);
xnor U4979 (N_4979,N_3856,N_3883);
xor U4980 (N_4980,N_3621,N_3128);
and U4981 (N_4981,N_3136,N_3894);
nor U4982 (N_4982,N_3540,N_3535);
and U4983 (N_4983,N_3496,N_3182);
nand U4984 (N_4984,N_3191,N_3199);
or U4985 (N_4985,N_3965,N_3060);
nor U4986 (N_4986,N_3847,N_3824);
nand U4987 (N_4987,N_3378,N_3236);
nand U4988 (N_4988,N_3229,N_3090);
xor U4989 (N_4989,N_3436,N_3002);
nor U4990 (N_4990,N_3638,N_3796);
nor U4991 (N_4991,N_3552,N_3662);
and U4992 (N_4992,N_3695,N_3405);
nand U4993 (N_4993,N_3923,N_3773);
nand U4994 (N_4994,N_3168,N_3069);
nand U4995 (N_4995,N_3056,N_3420);
xor U4996 (N_4996,N_3305,N_3284);
or U4997 (N_4997,N_3191,N_3293);
nor U4998 (N_4998,N_3987,N_3792);
nand U4999 (N_4999,N_3975,N_3763);
and U5000 (N_5000,N_4421,N_4508);
nor U5001 (N_5001,N_4476,N_4569);
nor U5002 (N_5002,N_4218,N_4768);
nor U5003 (N_5003,N_4622,N_4153);
and U5004 (N_5004,N_4752,N_4095);
nor U5005 (N_5005,N_4662,N_4681);
nor U5006 (N_5006,N_4015,N_4939);
nor U5007 (N_5007,N_4193,N_4774);
nand U5008 (N_5008,N_4607,N_4370);
and U5009 (N_5009,N_4783,N_4860);
or U5010 (N_5010,N_4328,N_4778);
or U5011 (N_5011,N_4532,N_4758);
and U5012 (N_5012,N_4110,N_4912);
or U5013 (N_5013,N_4143,N_4924);
nand U5014 (N_5014,N_4235,N_4058);
xnor U5015 (N_5015,N_4736,N_4066);
xor U5016 (N_5016,N_4424,N_4333);
xor U5017 (N_5017,N_4555,N_4059);
or U5018 (N_5018,N_4200,N_4352);
or U5019 (N_5019,N_4971,N_4790);
and U5020 (N_5020,N_4477,N_4678);
or U5021 (N_5021,N_4544,N_4405);
and U5022 (N_5022,N_4220,N_4417);
or U5023 (N_5023,N_4668,N_4787);
nor U5024 (N_5024,N_4760,N_4517);
and U5025 (N_5025,N_4265,N_4561);
xnor U5026 (N_5026,N_4208,N_4547);
nand U5027 (N_5027,N_4531,N_4753);
xor U5028 (N_5028,N_4746,N_4088);
or U5029 (N_5029,N_4779,N_4267);
xor U5030 (N_5030,N_4604,N_4827);
and U5031 (N_5031,N_4441,N_4907);
or U5032 (N_5032,N_4070,N_4588);
or U5033 (N_5033,N_4254,N_4534);
nor U5034 (N_5034,N_4603,N_4763);
nand U5035 (N_5035,N_4712,N_4455);
and U5036 (N_5036,N_4640,N_4967);
nor U5037 (N_5037,N_4324,N_4238);
xnor U5038 (N_5038,N_4909,N_4710);
xor U5039 (N_5039,N_4705,N_4770);
and U5040 (N_5040,N_4145,N_4935);
nor U5041 (N_5041,N_4700,N_4557);
nand U5042 (N_5042,N_4180,N_4849);
nor U5043 (N_5043,N_4359,N_4574);
xnor U5044 (N_5044,N_4259,N_4762);
and U5045 (N_5045,N_4624,N_4519);
nor U5046 (N_5046,N_4635,N_4985);
nor U5047 (N_5047,N_4659,N_4643);
nor U5048 (N_5048,N_4910,N_4196);
and U5049 (N_5049,N_4229,N_4191);
xor U5050 (N_5050,N_4123,N_4055);
and U5051 (N_5051,N_4564,N_4577);
and U5052 (N_5052,N_4018,N_4396);
or U5053 (N_5053,N_4704,N_4387);
nand U5054 (N_5054,N_4261,N_4187);
xnor U5055 (N_5055,N_4579,N_4136);
or U5056 (N_5056,N_4116,N_4642);
nor U5057 (N_5057,N_4067,N_4959);
nand U5058 (N_5058,N_4669,N_4583);
or U5059 (N_5059,N_4269,N_4843);
nand U5060 (N_5060,N_4848,N_4799);
and U5061 (N_5061,N_4231,N_4587);
nand U5062 (N_5062,N_4245,N_4166);
nor U5063 (N_5063,N_4483,N_4862);
xor U5064 (N_5064,N_4791,N_4820);
or U5065 (N_5065,N_4498,N_4479);
nor U5066 (N_5066,N_4402,N_4741);
nor U5067 (N_5067,N_4284,N_4727);
and U5068 (N_5068,N_4380,N_4696);
and U5069 (N_5069,N_4751,N_4335);
nor U5070 (N_5070,N_4020,N_4953);
or U5071 (N_5071,N_4992,N_4296);
or U5072 (N_5072,N_4307,N_4771);
xor U5073 (N_5073,N_4309,N_4589);
nand U5074 (N_5074,N_4379,N_4950);
nor U5075 (N_5075,N_4899,N_4318);
xnor U5076 (N_5076,N_4454,N_4581);
xor U5077 (N_5077,N_4052,N_4027);
nand U5078 (N_5078,N_4797,N_4809);
nor U5079 (N_5079,N_4528,N_4829);
nor U5080 (N_5080,N_4845,N_4775);
and U5081 (N_5081,N_4492,N_4051);
nor U5082 (N_5082,N_4369,N_4701);
nand U5083 (N_5083,N_4693,N_4942);
or U5084 (N_5084,N_4853,N_4375);
nand U5085 (N_5085,N_4515,N_4157);
or U5086 (N_5086,N_4553,N_4175);
xor U5087 (N_5087,N_4916,N_4716);
nand U5088 (N_5088,N_4888,N_4425);
nor U5089 (N_5089,N_4340,N_4349);
xor U5090 (N_5090,N_4486,N_4748);
and U5091 (N_5091,N_4445,N_4937);
and U5092 (N_5092,N_4972,N_4135);
or U5093 (N_5093,N_4004,N_4329);
nor U5094 (N_5094,N_4825,N_4986);
or U5095 (N_5095,N_4543,N_4851);
nor U5096 (N_5096,N_4154,N_4976);
nand U5097 (N_5097,N_4708,N_4767);
xor U5098 (N_5098,N_4031,N_4895);
nand U5099 (N_5099,N_4086,N_4317);
or U5100 (N_5100,N_4687,N_4538);
or U5101 (N_5101,N_4459,N_4563);
or U5102 (N_5102,N_4398,N_4788);
nand U5103 (N_5103,N_4395,N_4620);
and U5104 (N_5104,N_4392,N_4679);
xor U5105 (N_5105,N_4203,N_4279);
and U5106 (N_5106,N_4142,N_4499);
and U5107 (N_5107,N_4955,N_4242);
xor U5108 (N_5108,N_4949,N_4868);
nand U5109 (N_5109,N_4163,N_4990);
or U5110 (N_5110,N_4209,N_4301);
nand U5111 (N_5111,N_4570,N_4817);
xor U5112 (N_5112,N_4761,N_4830);
or U5113 (N_5113,N_4994,N_4075);
nor U5114 (N_5114,N_4198,N_4054);
nand U5115 (N_5115,N_4101,N_4729);
and U5116 (N_5116,N_4453,N_4996);
xor U5117 (N_5117,N_4093,N_4199);
and U5118 (N_5118,N_4133,N_4128);
or U5119 (N_5119,N_4011,N_4444);
or U5120 (N_5120,N_4155,N_4420);
xor U5121 (N_5121,N_4661,N_4697);
and U5122 (N_5122,N_4702,N_4523);
xor U5123 (N_5123,N_4594,N_4390);
nor U5124 (N_5124,N_4602,N_4836);
nor U5125 (N_5125,N_4368,N_4458);
or U5126 (N_5126,N_4546,N_4513);
xor U5127 (N_5127,N_4393,N_4367);
nor U5128 (N_5128,N_4177,N_4344);
nor U5129 (N_5129,N_4091,N_4025);
nand U5130 (N_5130,N_4934,N_4426);
or U5131 (N_5131,N_4832,N_4718);
and U5132 (N_5132,N_4884,N_4595);
or U5133 (N_5133,N_4898,N_4422);
nand U5134 (N_5134,N_4789,N_4504);
or U5135 (N_5135,N_4695,N_4673);
nor U5136 (N_5136,N_4464,N_4008);
or U5137 (N_5137,N_4326,N_4711);
or U5138 (N_5138,N_4999,N_4130);
nor U5139 (N_5139,N_4389,N_4707);
xor U5140 (N_5140,N_4260,N_4432);
and U5141 (N_5141,N_4501,N_4472);
nand U5142 (N_5142,N_4096,N_4026);
nand U5143 (N_5143,N_4403,N_4858);
nor U5144 (N_5144,N_4150,N_4740);
nor U5145 (N_5145,N_4911,N_4883);
and U5146 (N_5146,N_4225,N_4354);
nor U5147 (N_5147,N_4295,N_4300);
or U5148 (N_5148,N_4981,N_4212);
nand U5149 (N_5149,N_4724,N_4733);
and U5150 (N_5150,N_4435,N_4144);
or U5151 (N_5151,N_4772,N_4965);
nand U5152 (N_5152,N_4902,N_4289);
or U5153 (N_5153,N_4062,N_4222);
nand U5154 (N_5154,N_4415,N_4140);
or U5155 (N_5155,N_4606,N_4512);
xor U5156 (N_5156,N_4958,N_4106);
nand U5157 (N_5157,N_4255,N_4944);
and U5158 (N_5158,N_4005,N_4892);
or U5159 (N_5159,N_4671,N_4630);
nor U5160 (N_5160,N_4615,N_4009);
or U5161 (N_5161,N_4164,N_4539);
nor U5162 (N_5162,N_4725,N_4514);
nand U5163 (N_5163,N_4690,N_4619);
nand U5164 (N_5164,N_4556,N_4548);
nand U5165 (N_5165,N_4361,N_4156);
or U5166 (N_5166,N_4112,N_4754);
and U5167 (N_5167,N_4223,N_4074);
nand U5168 (N_5168,N_4795,N_4475);
or U5169 (N_5169,N_4131,N_4675);
or U5170 (N_5170,N_4565,N_4184);
nand U5171 (N_5171,N_4102,N_4765);
xor U5172 (N_5172,N_4505,N_4645);
xor U5173 (N_5173,N_4174,N_4171);
or U5174 (N_5174,N_4713,N_4646);
xnor U5175 (N_5175,N_4806,N_4400);
and U5176 (N_5176,N_4998,N_4658);
or U5177 (N_5177,N_4306,N_4134);
nand U5178 (N_5178,N_4566,N_4535);
nand U5179 (N_5179,N_4285,N_4777);
or U5180 (N_5180,N_4489,N_4537);
xnor U5181 (N_5181,N_4315,N_4742);
xnor U5182 (N_5182,N_4350,N_4703);
nor U5183 (N_5183,N_4889,N_4536);
or U5184 (N_5184,N_4650,N_4068);
or U5185 (N_5185,N_4132,N_4064);
xnor U5186 (N_5186,N_4356,N_4372);
xnor U5187 (N_5187,N_4663,N_4172);
or U5188 (N_5188,N_4303,N_4197);
nor U5189 (N_5189,N_4709,N_4666);
and U5190 (N_5190,N_4342,N_4946);
or U5191 (N_5191,N_4804,N_4207);
nand U5192 (N_5192,N_4629,N_4921);
nand U5193 (N_5193,N_4069,N_4217);
nor U5194 (N_5194,N_4966,N_4931);
xnor U5195 (N_5195,N_4462,N_4964);
nand U5196 (N_5196,N_4919,N_4449);
nor U5197 (N_5197,N_4468,N_4183);
or U5198 (N_5198,N_4840,N_4573);
nor U5199 (N_5199,N_4006,N_4117);
nor U5200 (N_5200,N_4757,N_4168);
nand U5201 (N_5201,N_4842,N_4147);
nand U5202 (N_5202,N_4305,N_4865);
nand U5203 (N_5203,N_4118,N_4854);
and U5204 (N_5204,N_4381,N_4287);
nand U5205 (N_5205,N_4078,N_4228);
or U5206 (N_5206,N_4451,N_4507);
nand U5207 (N_5207,N_4818,N_4816);
or U5208 (N_5208,N_4029,N_4126);
or U5209 (N_5209,N_4003,N_4580);
or U5210 (N_5210,N_4060,N_4181);
and U5211 (N_5211,N_4363,N_4439);
or U5212 (N_5212,N_4520,N_4796);
xnor U5213 (N_5213,N_4518,N_4234);
nand U5214 (N_5214,N_4657,N_4600);
xnor U5215 (N_5215,N_4291,N_4221);
or U5216 (N_5216,N_4276,N_4979);
and U5217 (N_5217,N_4429,N_4723);
xnor U5218 (N_5218,N_4022,N_4855);
nor U5219 (N_5219,N_4469,N_4956);
nand U5220 (N_5220,N_4694,N_4169);
and U5221 (N_5221,N_4656,N_4272);
xnor U5222 (N_5222,N_4598,N_4104);
and U5223 (N_5223,N_4253,N_4744);
nand U5224 (N_5224,N_4378,N_4347);
and U5225 (N_5225,N_4404,N_4418);
nand U5226 (N_5226,N_4552,N_4735);
and U5227 (N_5227,N_4745,N_4802);
and U5228 (N_5228,N_4590,N_4807);
and U5229 (N_5229,N_4491,N_4618);
nor U5230 (N_5230,N_4685,N_4576);
nand U5231 (N_5231,N_4360,N_4391);
nor U5232 (N_5232,N_4083,N_4894);
xor U5233 (N_5233,N_4857,N_4991);
nand U5234 (N_5234,N_4812,N_4293);
nor U5235 (N_5235,N_4384,N_4339);
nand U5236 (N_5236,N_4323,N_4412);
nand U5237 (N_5237,N_4097,N_4664);
nand U5238 (N_5238,N_4028,N_4322);
xor U5239 (N_5239,N_4376,N_4691);
nor U5240 (N_5240,N_4672,N_4948);
and U5241 (N_5241,N_4636,N_4159);
nor U5242 (N_5242,N_4905,N_4252);
nand U5243 (N_5243,N_4877,N_4073);
and U5244 (N_5244,N_4080,N_4227);
nor U5245 (N_5245,N_4192,N_4962);
and U5246 (N_5246,N_4871,N_4194);
xnor U5247 (N_5247,N_4283,N_4906);
nand U5248 (N_5248,N_4431,N_4401);
xnor U5249 (N_5249,N_4461,N_4639);
nand U5250 (N_5250,N_4353,N_4012);
nor U5251 (N_5251,N_4286,N_4688);
nor U5252 (N_5252,N_4633,N_4509);
nand U5253 (N_5253,N_4822,N_4978);
and U5254 (N_5254,N_4731,N_4852);
or U5255 (N_5255,N_4511,N_4021);
or U5256 (N_5256,N_4719,N_4918);
nor U5257 (N_5257,N_4016,N_4933);
or U5258 (N_5258,N_4647,N_4188);
nand U5259 (N_5259,N_4108,N_4148);
nor U5260 (N_5260,N_4500,N_4968);
nand U5261 (N_5261,N_4626,N_4308);
or U5262 (N_5262,N_4875,N_4035);
xor U5263 (N_5263,N_4699,N_4533);
and U5264 (N_5264,N_4450,N_4794);
nand U5265 (N_5265,N_4575,N_4559);
nor U5266 (N_5266,N_4219,N_4264);
nor U5267 (N_5267,N_4119,N_4407);
nand U5268 (N_5268,N_4487,N_4081);
nand U5269 (N_5269,N_4571,N_4438);
and U5270 (N_5270,N_4542,N_4204);
nand U5271 (N_5271,N_4605,N_4951);
or U5272 (N_5272,N_4747,N_4715);
nand U5273 (N_5273,N_4427,N_4230);
xnor U5274 (N_5274,N_4808,N_4529);
nand U5275 (N_5275,N_4525,N_4879);
nor U5276 (N_5276,N_4961,N_4516);
or U5277 (N_5277,N_4541,N_4125);
nand U5278 (N_5278,N_4792,N_4304);
and U5279 (N_5279,N_4692,N_4819);
or U5280 (N_5280,N_4103,N_4292);
xnor U5281 (N_5281,N_4258,N_4210);
or U5282 (N_5282,N_4846,N_4170);
nor U5283 (N_5283,N_4482,N_4969);
or U5284 (N_5284,N_4162,N_4313);
or U5285 (N_5285,N_4769,N_4087);
or U5286 (N_5286,N_4365,N_4109);
or U5287 (N_5287,N_4443,N_4540);
and U5288 (N_5288,N_4382,N_4874);
nand U5289 (N_5289,N_4176,N_4625);
xor U5290 (N_5290,N_4474,N_4173);
and U5291 (N_5291,N_4152,N_4090);
xnor U5292 (N_5292,N_4338,N_4728);
xor U5293 (N_5293,N_4608,N_4811);
nor U5294 (N_5294,N_4341,N_4885);
nor U5295 (N_5295,N_4017,N_4383);
nor U5296 (N_5296,N_4179,N_4205);
nor U5297 (N_5297,N_4881,N_4586);
and U5298 (N_5298,N_4739,N_4050);
xnor U5299 (N_5299,N_4801,N_4810);
or U5300 (N_5300,N_4866,N_4038);
xnor U5301 (N_5301,N_4226,N_4936);
or U5302 (N_5302,N_4914,N_4121);
and U5303 (N_5303,N_4730,N_4684);
nor U5304 (N_5304,N_4861,N_4214);
or U5305 (N_5305,N_4495,N_4077);
nor U5306 (N_5306,N_4872,N_4092);
or U5307 (N_5307,N_4036,N_4995);
or U5308 (N_5308,N_4397,N_4567);
nand U5309 (N_5309,N_4655,N_4616);
nand U5310 (N_5310,N_4446,N_4030);
or U5311 (N_5311,N_4257,N_4913);
nor U5312 (N_5312,N_4290,N_4545);
and U5313 (N_5313,N_4677,N_4270);
nand U5314 (N_5314,N_4037,N_4977);
or U5315 (N_5315,N_4847,N_4798);
nand U5316 (N_5316,N_4274,N_4190);
nor U5317 (N_5317,N_4597,N_4465);
and U5318 (N_5318,N_4249,N_4720);
nand U5319 (N_5319,N_4185,N_4355);
and U5320 (N_5320,N_4149,N_4882);
or U5321 (N_5321,N_4759,N_4273);
nand U5322 (N_5322,N_4281,N_4165);
xor U5323 (N_5323,N_4325,N_4084);
nand U5324 (N_5324,N_4665,N_4637);
xor U5325 (N_5325,N_4129,N_4813);
nand U5326 (N_5326,N_4114,N_4923);
or U5327 (N_5327,N_4714,N_4621);
nand U5328 (N_5328,N_4124,N_4063);
nor U5329 (N_5329,N_4034,N_4294);
nand U5330 (N_5330,N_4593,N_4984);
or U5331 (N_5331,N_4271,N_4330);
and U5332 (N_5332,N_4473,N_4319);
nand U5333 (N_5333,N_4072,N_4526);
and U5334 (N_5334,N_4146,N_4357);
and U5335 (N_5335,N_4332,N_4952);
xnor U5336 (N_5336,N_4151,N_4000);
nand U5337 (N_5337,N_4244,N_4929);
nor U5338 (N_5338,N_4189,N_4614);
nand U5339 (N_5339,N_4127,N_4256);
and U5340 (N_5340,N_4388,N_4945);
nor U5341 (N_5341,N_4764,N_4056);
or U5342 (N_5342,N_4698,N_4887);
nand U5343 (N_5343,N_4886,N_4240);
and U5344 (N_5344,N_4496,N_4239);
nor U5345 (N_5345,N_4631,N_4299);
xnor U5346 (N_5346,N_4442,N_4298);
nor U5347 (N_5347,N_4467,N_4480);
xor U5348 (N_5348,N_4917,N_4850);
nor U5349 (N_5349,N_4987,N_4649);
xnor U5350 (N_5350,N_4766,N_4551);
and U5351 (N_5351,N_4206,N_4686);
and U5352 (N_5352,N_4925,N_4471);
nand U5353 (N_5353,N_4841,N_4139);
xnor U5354 (N_5354,N_4186,N_4568);
nand U5355 (N_5355,N_4793,N_4111);
xnor U5356 (N_5356,N_4824,N_4839);
nor U5357 (N_5357,N_4947,N_4364);
nand U5358 (N_5358,N_4867,N_4706);
xnor U5359 (N_5359,N_4048,N_4043);
xnor U5360 (N_5360,N_4901,N_4503);
nor U5361 (N_5361,N_4282,N_4033);
xnor U5362 (N_5362,N_4302,N_4896);
nor U5363 (N_5363,N_4076,N_4628);
or U5364 (N_5364,N_4413,N_4634);
nor U5365 (N_5365,N_4447,N_4178);
and U5366 (N_5366,N_4236,N_4821);
nand U5367 (N_5367,N_4457,N_4488);
nand U5368 (N_5368,N_4859,N_4115);
and U5369 (N_5369,N_4416,N_4044);
nand U5370 (N_5370,N_4558,N_4927);
xor U5371 (N_5371,N_4202,N_4419);
nor U5372 (N_5372,N_4611,N_4960);
nor U5373 (N_5373,N_4920,N_4617);
or U5374 (N_5374,N_4311,N_4410);
and U5375 (N_5375,N_4478,N_4932);
nand U5376 (N_5376,N_4988,N_4079);
and U5377 (N_5377,N_4481,N_4609);
or U5378 (N_5378,N_4348,N_4366);
nand U5379 (N_5379,N_4786,N_4232);
or U5380 (N_5380,N_4247,N_4652);
xnor U5381 (N_5381,N_4592,N_4835);
xor U5382 (N_5382,N_4737,N_4963);
and U5383 (N_5383,N_4434,N_4343);
nand U5384 (N_5384,N_4160,N_4041);
nor U5385 (N_5385,N_4312,N_4674);
xnor U5386 (N_5386,N_4893,N_4408);
nor U5387 (N_5387,N_4336,N_4900);
nand U5388 (N_5388,N_4904,N_4237);
or U5389 (N_5389,N_4823,N_4627);
nand U5390 (N_5390,N_4107,N_4406);
and U5391 (N_5391,N_4409,N_4833);
xnor U5392 (N_5392,N_4922,N_4394);
xnor U5393 (N_5393,N_4834,N_4930);
and U5394 (N_5394,N_4463,N_4989);
and U5395 (N_5395,N_4680,N_4785);
xnor U5396 (N_5396,N_4550,N_4195);
and U5397 (N_5397,N_4549,N_4099);
nor U5398 (N_5398,N_4601,N_4815);
nand U5399 (N_5399,N_4460,N_4980);
xor U5400 (N_5400,N_4094,N_4456);
xor U5401 (N_5401,N_4466,N_4399);
and U5402 (N_5402,N_4982,N_4873);
or U5403 (N_5403,N_4734,N_4373);
nand U5404 (N_5404,N_4554,N_4584);
nand U5405 (N_5405,N_4277,N_4032);
nand U5406 (N_5406,N_4440,N_4938);
nand U5407 (N_5407,N_4120,N_4870);
and U5408 (N_5408,N_4057,N_4660);
and U5409 (N_5409,N_4493,N_4891);
nand U5410 (N_5410,N_4497,N_4137);
xnor U5411 (N_5411,N_4053,N_4755);
nor U5412 (N_5412,N_4837,N_4585);
nor U5413 (N_5413,N_4975,N_4738);
and U5414 (N_5414,N_4844,N_4013);
nand U5415 (N_5415,N_4897,N_4262);
nor U5416 (N_5416,N_4831,N_4250);
nor U5417 (N_5417,N_4863,N_4122);
nand U5418 (N_5418,N_4334,N_4377);
xor U5419 (N_5419,N_4828,N_4803);
or U5420 (N_5420,N_4374,N_4638);
and U5421 (N_5421,N_4411,N_4327);
or U5422 (N_5422,N_4019,N_4141);
or U5423 (N_5423,N_4161,N_4527);
nand U5424 (N_5424,N_4623,N_4158);
nor U5425 (N_5425,N_4266,N_4732);
xor U5426 (N_5426,N_4014,N_4437);
nand U5427 (N_5427,N_4805,N_4610);
nor U5428 (N_5428,N_4098,N_4908);
and U5429 (N_5429,N_4082,N_4915);
xnor U5430 (N_5430,N_4814,N_4780);
xnor U5431 (N_5431,N_4876,N_4903);
xor U5432 (N_5432,N_4138,N_4484);
or U5433 (N_5433,N_4040,N_4670);
xnor U5434 (N_5434,N_4530,N_4448);
and U5435 (N_5435,N_4973,N_4248);
nand U5436 (N_5436,N_4049,N_4275);
nor U5437 (N_5437,N_4717,N_4251);
nor U5438 (N_5438,N_4337,N_4560);
or U5439 (N_5439,N_4452,N_4345);
and U5440 (N_5440,N_4878,N_4351);
xnor U5441 (N_5441,N_4926,N_4582);
or U5442 (N_5442,N_4683,N_4838);
xnor U5443 (N_5443,N_4423,N_4726);
and U5444 (N_5444,N_4320,N_4105);
and U5445 (N_5445,N_4268,N_4494);
nor U5446 (N_5446,N_4782,N_4100);
and U5447 (N_5447,N_4502,N_4689);
and U5448 (N_5448,N_4721,N_4648);
xnor U5449 (N_5449,N_4596,N_4023);
or U5450 (N_5450,N_4215,N_4784);
xnor U5451 (N_5451,N_4224,N_4773);
nor U5452 (N_5452,N_4045,N_4297);
nor U5453 (N_5453,N_4362,N_4243);
nand U5454 (N_5454,N_4007,N_4386);
xnor U5455 (N_5455,N_4433,N_4957);
nand U5456 (N_5456,N_4941,N_4321);
and U5457 (N_5457,N_4167,N_4997);
or U5458 (N_5458,N_4983,N_4358);
or U5459 (N_5459,N_4233,N_4263);
and U5460 (N_5460,N_4346,N_4993);
and U5461 (N_5461,N_4940,N_4385);
xnor U5462 (N_5462,N_4470,N_4521);
nand U5463 (N_5463,N_4241,N_4316);
nand U5464 (N_5464,N_4641,N_4781);
and U5465 (N_5465,N_4667,N_4880);
nor U5466 (N_5466,N_4201,N_4756);
or U5467 (N_5467,N_4061,N_4800);
xnor U5468 (N_5468,N_4750,N_4613);
nor U5469 (N_5469,N_4001,N_4213);
and U5470 (N_5470,N_4591,N_4651);
nor U5471 (N_5471,N_4869,N_4371);
xnor U5472 (N_5472,N_4042,N_4414);
or U5473 (N_5473,N_4522,N_4211);
xnor U5474 (N_5474,N_4722,N_4485);
nand U5475 (N_5475,N_4599,N_4182);
nor U5476 (N_5476,N_4676,N_4749);
xnor U5477 (N_5477,N_4644,N_4943);
or U5478 (N_5478,N_4970,N_4024);
xnor U5479 (N_5479,N_4436,N_4524);
xnor U5480 (N_5480,N_4632,N_4928);
nand U5481 (N_5481,N_4089,N_4331);
nand U5482 (N_5482,N_4510,N_4246);
and U5483 (N_5483,N_4654,N_4002);
xor U5484 (N_5484,N_4954,N_4278);
or U5485 (N_5485,N_4776,N_4826);
xnor U5486 (N_5486,N_4743,N_4314);
nor U5487 (N_5487,N_4280,N_4039);
or U5488 (N_5488,N_4310,N_4065);
nor U5489 (N_5489,N_4490,N_4612);
xor U5490 (N_5490,N_4430,N_4071);
nor U5491 (N_5491,N_4288,N_4572);
or U5492 (N_5492,N_4856,N_4562);
nand U5493 (N_5493,N_4864,N_4653);
xor U5494 (N_5494,N_4506,N_4578);
and U5495 (N_5495,N_4113,N_4216);
nand U5496 (N_5496,N_4010,N_4890);
nor U5497 (N_5497,N_4085,N_4047);
or U5498 (N_5498,N_4046,N_4428);
xor U5499 (N_5499,N_4974,N_4682);
xor U5500 (N_5500,N_4611,N_4747);
nand U5501 (N_5501,N_4419,N_4944);
and U5502 (N_5502,N_4562,N_4021);
xor U5503 (N_5503,N_4146,N_4304);
and U5504 (N_5504,N_4792,N_4288);
or U5505 (N_5505,N_4145,N_4891);
nor U5506 (N_5506,N_4838,N_4116);
nand U5507 (N_5507,N_4916,N_4509);
xnor U5508 (N_5508,N_4703,N_4453);
or U5509 (N_5509,N_4790,N_4322);
nand U5510 (N_5510,N_4233,N_4482);
xor U5511 (N_5511,N_4481,N_4094);
nand U5512 (N_5512,N_4131,N_4998);
nand U5513 (N_5513,N_4909,N_4779);
or U5514 (N_5514,N_4910,N_4521);
xnor U5515 (N_5515,N_4495,N_4913);
or U5516 (N_5516,N_4790,N_4687);
and U5517 (N_5517,N_4032,N_4314);
nor U5518 (N_5518,N_4850,N_4939);
nor U5519 (N_5519,N_4077,N_4371);
xnor U5520 (N_5520,N_4020,N_4623);
nand U5521 (N_5521,N_4549,N_4504);
nand U5522 (N_5522,N_4603,N_4485);
nor U5523 (N_5523,N_4911,N_4371);
xnor U5524 (N_5524,N_4636,N_4187);
and U5525 (N_5525,N_4509,N_4959);
nand U5526 (N_5526,N_4792,N_4922);
xor U5527 (N_5527,N_4502,N_4267);
nand U5528 (N_5528,N_4135,N_4534);
and U5529 (N_5529,N_4784,N_4424);
nand U5530 (N_5530,N_4239,N_4823);
and U5531 (N_5531,N_4701,N_4404);
or U5532 (N_5532,N_4761,N_4125);
nor U5533 (N_5533,N_4759,N_4416);
nor U5534 (N_5534,N_4090,N_4773);
xor U5535 (N_5535,N_4276,N_4545);
nand U5536 (N_5536,N_4793,N_4328);
nand U5537 (N_5537,N_4863,N_4826);
and U5538 (N_5538,N_4300,N_4722);
nor U5539 (N_5539,N_4701,N_4706);
or U5540 (N_5540,N_4122,N_4991);
nor U5541 (N_5541,N_4022,N_4407);
xnor U5542 (N_5542,N_4848,N_4319);
nor U5543 (N_5543,N_4826,N_4468);
or U5544 (N_5544,N_4597,N_4412);
nand U5545 (N_5545,N_4898,N_4665);
and U5546 (N_5546,N_4692,N_4563);
and U5547 (N_5547,N_4399,N_4732);
nor U5548 (N_5548,N_4843,N_4461);
xnor U5549 (N_5549,N_4808,N_4652);
and U5550 (N_5550,N_4688,N_4658);
or U5551 (N_5551,N_4540,N_4992);
xor U5552 (N_5552,N_4532,N_4374);
nand U5553 (N_5553,N_4449,N_4845);
nand U5554 (N_5554,N_4857,N_4483);
xnor U5555 (N_5555,N_4802,N_4070);
nand U5556 (N_5556,N_4506,N_4831);
xor U5557 (N_5557,N_4135,N_4224);
or U5558 (N_5558,N_4972,N_4585);
xor U5559 (N_5559,N_4662,N_4886);
and U5560 (N_5560,N_4242,N_4041);
or U5561 (N_5561,N_4435,N_4306);
and U5562 (N_5562,N_4143,N_4290);
nand U5563 (N_5563,N_4108,N_4994);
nand U5564 (N_5564,N_4326,N_4508);
and U5565 (N_5565,N_4444,N_4190);
and U5566 (N_5566,N_4573,N_4518);
xor U5567 (N_5567,N_4747,N_4826);
xnor U5568 (N_5568,N_4741,N_4159);
nand U5569 (N_5569,N_4218,N_4395);
nor U5570 (N_5570,N_4694,N_4064);
xor U5571 (N_5571,N_4992,N_4210);
xor U5572 (N_5572,N_4287,N_4394);
nor U5573 (N_5573,N_4367,N_4573);
nand U5574 (N_5574,N_4479,N_4771);
or U5575 (N_5575,N_4591,N_4666);
nor U5576 (N_5576,N_4287,N_4555);
and U5577 (N_5577,N_4018,N_4213);
nand U5578 (N_5578,N_4361,N_4837);
nand U5579 (N_5579,N_4415,N_4688);
nand U5580 (N_5580,N_4542,N_4447);
nand U5581 (N_5581,N_4758,N_4338);
or U5582 (N_5582,N_4064,N_4418);
nor U5583 (N_5583,N_4084,N_4892);
or U5584 (N_5584,N_4926,N_4558);
xnor U5585 (N_5585,N_4430,N_4117);
or U5586 (N_5586,N_4919,N_4751);
nor U5587 (N_5587,N_4553,N_4023);
or U5588 (N_5588,N_4370,N_4041);
nor U5589 (N_5589,N_4790,N_4510);
xnor U5590 (N_5590,N_4183,N_4137);
xnor U5591 (N_5591,N_4709,N_4190);
and U5592 (N_5592,N_4850,N_4711);
nand U5593 (N_5593,N_4000,N_4563);
or U5594 (N_5594,N_4164,N_4743);
or U5595 (N_5595,N_4259,N_4458);
or U5596 (N_5596,N_4839,N_4886);
or U5597 (N_5597,N_4834,N_4868);
xnor U5598 (N_5598,N_4895,N_4253);
and U5599 (N_5599,N_4149,N_4577);
xor U5600 (N_5600,N_4155,N_4343);
or U5601 (N_5601,N_4320,N_4373);
or U5602 (N_5602,N_4966,N_4882);
xnor U5603 (N_5603,N_4392,N_4043);
nor U5604 (N_5604,N_4290,N_4107);
xor U5605 (N_5605,N_4329,N_4592);
nand U5606 (N_5606,N_4303,N_4872);
xor U5607 (N_5607,N_4250,N_4983);
or U5608 (N_5608,N_4205,N_4323);
and U5609 (N_5609,N_4526,N_4641);
xor U5610 (N_5610,N_4741,N_4102);
nand U5611 (N_5611,N_4945,N_4856);
and U5612 (N_5612,N_4114,N_4186);
xor U5613 (N_5613,N_4909,N_4682);
and U5614 (N_5614,N_4330,N_4388);
nor U5615 (N_5615,N_4276,N_4533);
nand U5616 (N_5616,N_4750,N_4618);
and U5617 (N_5617,N_4881,N_4134);
and U5618 (N_5618,N_4689,N_4018);
nand U5619 (N_5619,N_4183,N_4094);
nor U5620 (N_5620,N_4240,N_4479);
or U5621 (N_5621,N_4592,N_4126);
and U5622 (N_5622,N_4345,N_4915);
xnor U5623 (N_5623,N_4511,N_4146);
nor U5624 (N_5624,N_4023,N_4043);
xor U5625 (N_5625,N_4304,N_4474);
nor U5626 (N_5626,N_4129,N_4075);
nor U5627 (N_5627,N_4534,N_4787);
nand U5628 (N_5628,N_4000,N_4908);
xnor U5629 (N_5629,N_4678,N_4025);
xnor U5630 (N_5630,N_4683,N_4681);
xnor U5631 (N_5631,N_4886,N_4979);
xnor U5632 (N_5632,N_4725,N_4026);
xnor U5633 (N_5633,N_4787,N_4285);
or U5634 (N_5634,N_4727,N_4384);
or U5635 (N_5635,N_4658,N_4636);
or U5636 (N_5636,N_4159,N_4983);
or U5637 (N_5637,N_4625,N_4736);
or U5638 (N_5638,N_4862,N_4215);
and U5639 (N_5639,N_4691,N_4604);
and U5640 (N_5640,N_4428,N_4985);
nand U5641 (N_5641,N_4249,N_4231);
xor U5642 (N_5642,N_4106,N_4999);
xnor U5643 (N_5643,N_4292,N_4306);
and U5644 (N_5644,N_4654,N_4425);
xnor U5645 (N_5645,N_4768,N_4611);
or U5646 (N_5646,N_4854,N_4766);
xnor U5647 (N_5647,N_4810,N_4272);
or U5648 (N_5648,N_4208,N_4136);
or U5649 (N_5649,N_4362,N_4521);
and U5650 (N_5650,N_4472,N_4243);
or U5651 (N_5651,N_4171,N_4415);
and U5652 (N_5652,N_4015,N_4252);
nor U5653 (N_5653,N_4916,N_4139);
nor U5654 (N_5654,N_4297,N_4321);
and U5655 (N_5655,N_4749,N_4962);
nor U5656 (N_5656,N_4678,N_4879);
nor U5657 (N_5657,N_4131,N_4251);
xnor U5658 (N_5658,N_4438,N_4699);
and U5659 (N_5659,N_4608,N_4806);
nor U5660 (N_5660,N_4479,N_4077);
nor U5661 (N_5661,N_4457,N_4857);
and U5662 (N_5662,N_4144,N_4380);
and U5663 (N_5663,N_4099,N_4594);
nand U5664 (N_5664,N_4544,N_4438);
nor U5665 (N_5665,N_4575,N_4739);
nand U5666 (N_5666,N_4492,N_4472);
xor U5667 (N_5667,N_4354,N_4531);
nor U5668 (N_5668,N_4197,N_4044);
nand U5669 (N_5669,N_4669,N_4761);
xnor U5670 (N_5670,N_4963,N_4137);
nand U5671 (N_5671,N_4448,N_4647);
and U5672 (N_5672,N_4794,N_4900);
nand U5673 (N_5673,N_4003,N_4615);
nand U5674 (N_5674,N_4247,N_4601);
and U5675 (N_5675,N_4324,N_4027);
nand U5676 (N_5676,N_4385,N_4171);
xor U5677 (N_5677,N_4197,N_4533);
nor U5678 (N_5678,N_4014,N_4314);
xor U5679 (N_5679,N_4820,N_4774);
or U5680 (N_5680,N_4953,N_4622);
nor U5681 (N_5681,N_4173,N_4388);
or U5682 (N_5682,N_4671,N_4922);
xor U5683 (N_5683,N_4020,N_4831);
nor U5684 (N_5684,N_4788,N_4231);
xnor U5685 (N_5685,N_4335,N_4269);
nor U5686 (N_5686,N_4495,N_4213);
or U5687 (N_5687,N_4083,N_4693);
nor U5688 (N_5688,N_4481,N_4923);
nand U5689 (N_5689,N_4621,N_4351);
xnor U5690 (N_5690,N_4906,N_4440);
nand U5691 (N_5691,N_4621,N_4249);
xnor U5692 (N_5692,N_4092,N_4647);
or U5693 (N_5693,N_4277,N_4267);
xnor U5694 (N_5694,N_4512,N_4705);
nand U5695 (N_5695,N_4401,N_4921);
nand U5696 (N_5696,N_4348,N_4060);
xor U5697 (N_5697,N_4793,N_4563);
nor U5698 (N_5698,N_4520,N_4399);
nor U5699 (N_5699,N_4371,N_4155);
or U5700 (N_5700,N_4363,N_4116);
nand U5701 (N_5701,N_4561,N_4858);
or U5702 (N_5702,N_4430,N_4491);
and U5703 (N_5703,N_4607,N_4034);
nor U5704 (N_5704,N_4292,N_4386);
nand U5705 (N_5705,N_4539,N_4802);
nand U5706 (N_5706,N_4244,N_4246);
xor U5707 (N_5707,N_4153,N_4484);
nand U5708 (N_5708,N_4211,N_4665);
xnor U5709 (N_5709,N_4121,N_4525);
nor U5710 (N_5710,N_4056,N_4571);
and U5711 (N_5711,N_4696,N_4535);
nor U5712 (N_5712,N_4141,N_4543);
nand U5713 (N_5713,N_4243,N_4036);
nor U5714 (N_5714,N_4409,N_4639);
and U5715 (N_5715,N_4490,N_4282);
or U5716 (N_5716,N_4876,N_4166);
or U5717 (N_5717,N_4844,N_4734);
xor U5718 (N_5718,N_4874,N_4344);
nand U5719 (N_5719,N_4472,N_4801);
nand U5720 (N_5720,N_4590,N_4871);
and U5721 (N_5721,N_4639,N_4764);
xnor U5722 (N_5722,N_4870,N_4503);
xnor U5723 (N_5723,N_4524,N_4837);
nor U5724 (N_5724,N_4060,N_4628);
or U5725 (N_5725,N_4113,N_4287);
nor U5726 (N_5726,N_4523,N_4940);
nor U5727 (N_5727,N_4086,N_4791);
nor U5728 (N_5728,N_4101,N_4395);
and U5729 (N_5729,N_4599,N_4342);
or U5730 (N_5730,N_4577,N_4061);
or U5731 (N_5731,N_4945,N_4501);
xor U5732 (N_5732,N_4125,N_4089);
and U5733 (N_5733,N_4497,N_4548);
nand U5734 (N_5734,N_4563,N_4565);
xnor U5735 (N_5735,N_4532,N_4573);
nand U5736 (N_5736,N_4075,N_4119);
and U5737 (N_5737,N_4329,N_4783);
or U5738 (N_5738,N_4878,N_4971);
xor U5739 (N_5739,N_4107,N_4839);
nand U5740 (N_5740,N_4138,N_4576);
or U5741 (N_5741,N_4050,N_4543);
nor U5742 (N_5742,N_4827,N_4073);
or U5743 (N_5743,N_4647,N_4187);
and U5744 (N_5744,N_4127,N_4416);
or U5745 (N_5745,N_4440,N_4799);
and U5746 (N_5746,N_4990,N_4245);
xnor U5747 (N_5747,N_4152,N_4506);
and U5748 (N_5748,N_4416,N_4155);
nand U5749 (N_5749,N_4351,N_4014);
nor U5750 (N_5750,N_4371,N_4305);
and U5751 (N_5751,N_4513,N_4573);
or U5752 (N_5752,N_4439,N_4880);
nor U5753 (N_5753,N_4577,N_4095);
and U5754 (N_5754,N_4498,N_4559);
xor U5755 (N_5755,N_4353,N_4977);
or U5756 (N_5756,N_4872,N_4413);
nor U5757 (N_5757,N_4889,N_4967);
nand U5758 (N_5758,N_4333,N_4663);
xor U5759 (N_5759,N_4221,N_4005);
nor U5760 (N_5760,N_4403,N_4847);
xor U5761 (N_5761,N_4096,N_4892);
nor U5762 (N_5762,N_4006,N_4082);
nor U5763 (N_5763,N_4208,N_4903);
and U5764 (N_5764,N_4315,N_4578);
and U5765 (N_5765,N_4770,N_4188);
nor U5766 (N_5766,N_4257,N_4817);
xnor U5767 (N_5767,N_4809,N_4660);
and U5768 (N_5768,N_4351,N_4237);
xnor U5769 (N_5769,N_4681,N_4610);
and U5770 (N_5770,N_4865,N_4620);
nand U5771 (N_5771,N_4702,N_4618);
xor U5772 (N_5772,N_4300,N_4101);
xnor U5773 (N_5773,N_4860,N_4712);
and U5774 (N_5774,N_4353,N_4849);
and U5775 (N_5775,N_4742,N_4680);
xnor U5776 (N_5776,N_4987,N_4728);
and U5777 (N_5777,N_4198,N_4183);
or U5778 (N_5778,N_4926,N_4832);
xnor U5779 (N_5779,N_4360,N_4579);
and U5780 (N_5780,N_4994,N_4248);
nand U5781 (N_5781,N_4969,N_4816);
and U5782 (N_5782,N_4406,N_4131);
nand U5783 (N_5783,N_4101,N_4124);
and U5784 (N_5784,N_4842,N_4388);
nor U5785 (N_5785,N_4690,N_4073);
and U5786 (N_5786,N_4309,N_4523);
and U5787 (N_5787,N_4796,N_4590);
nor U5788 (N_5788,N_4172,N_4728);
or U5789 (N_5789,N_4926,N_4080);
nor U5790 (N_5790,N_4736,N_4763);
and U5791 (N_5791,N_4606,N_4541);
and U5792 (N_5792,N_4512,N_4360);
or U5793 (N_5793,N_4386,N_4619);
or U5794 (N_5794,N_4258,N_4025);
nor U5795 (N_5795,N_4875,N_4000);
xor U5796 (N_5796,N_4440,N_4247);
or U5797 (N_5797,N_4061,N_4943);
and U5798 (N_5798,N_4963,N_4295);
nand U5799 (N_5799,N_4604,N_4247);
and U5800 (N_5800,N_4040,N_4820);
nand U5801 (N_5801,N_4751,N_4912);
nor U5802 (N_5802,N_4416,N_4987);
xor U5803 (N_5803,N_4711,N_4855);
xnor U5804 (N_5804,N_4593,N_4020);
and U5805 (N_5805,N_4671,N_4788);
or U5806 (N_5806,N_4602,N_4333);
or U5807 (N_5807,N_4229,N_4875);
and U5808 (N_5808,N_4802,N_4333);
nand U5809 (N_5809,N_4547,N_4706);
nor U5810 (N_5810,N_4435,N_4527);
nor U5811 (N_5811,N_4677,N_4866);
nor U5812 (N_5812,N_4781,N_4913);
nand U5813 (N_5813,N_4030,N_4313);
nor U5814 (N_5814,N_4237,N_4723);
and U5815 (N_5815,N_4640,N_4701);
nor U5816 (N_5816,N_4198,N_4888);
nor U5817 (N_5817,N_4918,N_4035);
nor U5818 (N_5818,N_4796,N_4442);
nand U5819 (N_5819,N_4416,N_4452);
or U5820 (N_5820,N_4039,N_4387);
and U5821 (N_5821,N_4339,N_4129);
nor U5822 (N_5822,N_4975,N_4780);
nand U5823 (N_5823,N_4142,N_4282);
or U5824 (N_5824,N_4190,N_4720);
or U5825 (N_5825,N_4285,N_4679);
xor U5826 (N_5826,N_4522,N_4800);
or U5827 (N_5827,N_4636,N_4178);
xnor U5828 (N_5828,N_4783,N_4976);
nor U5829 (N_5829,N_4114,N_4017);
or U5830 (N_5830,N_4950,N_4622);
xnor U5831 (N_5831,N_4356,N_4462);
nand U5832 (N_5832,N_4571,N_4369);
and U5833 (N_5833,N_4264,N_4571);
nor U5834 (N_5834,N_4329,N_4228);
nor U5835 (N_5835,N_4617,N_4139);
nand U5836 (N_5836,N_4559,N_4231);
xor U5837 (N_5837,N_4606,N_4991);
nor U5838 (N_5838,N_4533,N_4322);
nor U5839 (N_5839,N_4125,N_4146);
or U5840 (N_5840,N_4698,N_4435);
nor U5841 (N_5841,N_4661,N_4626);
and U5842 (N_5842,N_4203,N_4756);
nand U5843 (N_5843,N_4796,N_4477);
xor U5844 (N_5844,N_4960,N_4070);
and U5845 (N_5845,N_4016,N_4707);
xnor U5846 (N_5846,N_4874,N_4490);
xnor U5847 (N_5847,N_4444,N_4037);
xnor U5848 (N_5848,N_4489,N_4947);
or U5849 (N_5849,N_4458,N_4909);
nor U5850 (N_5850,N_4510,N_4156);
and U5851 (N_5851,N_4762,N_4546);
nand U5852 (N_5852,N_4987,N_4025);
xnor U5853 (N_5853,N_4412,N_4962);
xor U5854 (N_5854,N_4148,N_4761);
or U5855 (N_5855,N_4394,N_4977);
or U5856 (N_5856,N_4908,N_4726);
and U5857 (N_5857,N_4249,N_4516);
nor U5858 (N_5858,N_4204,N_4230);
nor U5859 (N_5859,N_4795,N_4309);
xnor U5860 (N_5860,N_4147,N_4256);
nor U5861 (N_5861,N_4821,N_4515);
xnor U5862 (N_5862,N_4967,N_4703);
or U5863 (N_5863,N_4705,N_4098);
or U5864 (N_5864,N_4490,N_4323);
and U5865 (N_5865,N_4001,N_4239);
nor U5866 (N_5866,N_4764,N_4020);
and U5867 (N_5867,N_4448,N_4816);
xnor U5868 (N_5868,N_4719,N_4811);
and U5869 (N_5869,N_4310,N_4379);
and U5870 (N_5870,N_4851,N_4347);
and U5871 (N_5871,N_4330,N_4883);
nand U5872 (N_5872,N_4256,N_4067);
nor U5873 (N_5873,N_4824,N_4538);
and U5874 (N_5874,N_4044,N_4921);
or U5875 (N_5875,N_4093,N_4487);
or U5876 (N_5876,N_4561,N_4086);
nor U5877 (N_5877,N_4338,N_4852);
and U5878 (N_5878,N_4712,N_4460);
and U5879 (N_5879,N_4169,N_4157);
nor U5880 (N_5880,N_4113,N_4373);
nand U5881 (N_5881,N_4115,N_4574);
or U5882 (N_5882,N_4629,N_4102);
xnor U5883 (N_5883,N_4730,N_4593);
and U5884 (N_5884,N_4536,N_4979);
xnor U5885 (N_5885,N_4799,N_4701);
nor U5886 (N_5886,N_4737,N_4566);
or U5887 (N_5887,N_4212,N_4214);
nor U5888 (N_5888,N_4562,N_4748);
nor U5889 (N_5889,N_4375,N_4345);
nor U5890 (N_5890,N_4868,N_4540);
xnor U5891 (N_5891,N_4474,N_4492);
or U5892 (N_5892,N_4529,N_4114);
nand U5893 (N_5893,N_4676,N_4416);
nand U5894 (N_5894,N_4959,N_4619);
xnor U5895 (N_5895,N_4072,N_4340);
nor U5896 (N_5896,N_4771,N_4840);
nand U5897 (N_5897,N_4313,N_4900);
xnor U5898 (N_5898,N_4604,N_4832);
or U5899 (N_5899,N_4944,N_4731);
or U5900 (N_5900,N_4004,N_4821);
nor U5901 (N_5901,N_4687,N_4889);
nand U5902 (N_5902,N_4140,N_4346);
or U5903 (N_5903,N_4002,N_4323);
or U5904 (N_5904,N_4015,N_4144);
xor U5905 (N_5905,N_4114,N_4845);
and U5906 (N_5906,N_4460,N_4621);
xnor U5907 (N_5907,N_4592,N_4271);
and U5908 (N_5908,N_4876,N_4265);
or U5909 (N_5909,N_4857,N_4649);
xnor U5910 (N_5910,N_4478,N_4852);
or U5911 (N_5911,N_4455,N_4872);
nor U5912 (N_5912,N_4147,N_4429);
xor U5913 (N_5913,N_4044,N_4096);
and U5914 (N_5914,N_4879,N_4869);
nand U5915 (N_5915,N_4982,N_4652);
or U5916 (N_5916,N_4573,N_4471);
xor U5917 (N_5917,N_4318,N_4840);
xor U5918 (N_5918,N_4214,N_4763);
or U5919 (N_5919,N_4365,N_4316);
nor U5920 (N_5920,N_4476,N_4215);
and U5921 (N_5921,N_4181,N_4828);
xor U5922 (N_5922,N_4771,N_4675);
and U5923 (N_5923,N_4776,N_4326);
nand U5924 (N_5924,N_4828,N_4831);
or U5925 (N_5925,N_4009,N_4798);
nand U5926 (N_5926,N_4216,N_4132);
nor U5927 (N_5927,N_4074,N_4852);
and U5928 (N_5928,N_4459,N_4337);
and U5929 (N_5929,N_4109,N_4165);
and U5930 (N_5930,N_4704,N_4959);
xor U5931 (N_5931,N_4703,N_4563);
or U5932 (N_5932,N_4882,N_4828);
and U5933 (N_5933,N_4198,N_4708);
nor U5934 (N_5934,N_4877,N_4380);
xnor U5935 (N_5935,N_4516,N_4346);
and U5936 (N_5936,N_4647,N_4186);
nand U5937 (N_5937,N_4957,N_4201);
nor U5938 (N_5938,N_4727,N_4501);
and U5939 (N_5939,N_4570,N_4122);
nand U5940 (N_5940,N_4161,N_4132);
nor U5941 (N_5941,N_4867,N_4255);
xnor U5942 (N_5942,N_4917,N_4086);
and U5943 (N_5943,N_4231,N_4450);
or U5944 (N_5944,N_4331,N_4925);
or U5945 (N_5945,N_4405,N_4524);
or U5946 (N_5946,N_4168,N_4512);
or U5947 (N_5947,N_4533,N_4025);
and U5948 (N_5948,N_4146,N_4840);
or U5949 (N_5949,N_4394,N_4742);
nand U5950 (N_5950,N_4568,N_4609);
nand U5951 (N_5951,N_4653,N_4932);
xor U5952 (N_5952,N_4628,N_4135);
or U5953 (N_5953,N_4912,N_4080);
or U5954 (N_5954,N_4162,N_4754);
and U5955 (N_5955,N_4572,N_4233);
or U5956 (N_5956,N_4810,N_4044);
or U5957 (N_5957,N_4568,N_4382);
or U5958 (N_5958,N_4616,N_4061);
xnor U5959 (N_5959,N_4023,N_4617);
or U5960 (N_5960,N_4780,N_4338);
and U5961 (N_5961,N_4310,N_4264);
and U5962 (N_5962,N_4270,N_4958);
and U5963 (N_5963,N_4225,N_4652);
or U5964 (N_5964,N_4205,N_4050);
nor U5965 (N_5965,N_4651,N_4947);
or U5966 (N_5966,N_4921,N_4344);
or U5967 (N_5967,N_4462,N_4691);
or U5968 (N_5968,N_4920,N_4951);
xor U5969 (N_5969,N_4912,N_4055);
and U5970 (N_5970,N_4263,N_4281);
and U5971 (N_5971,N_4255,N_4131);
or U5972 (N_5972,N_4093,N_4252);
nand U5973 (N_5973,N_4412,N_4528);
and U5974 (N_5974,N_4941,N_4010);
xnor U5975 (N_5975,N_4875,N_4882);
and U5976 (N_5976,N_4494,N_4647);
or U5977 (N_5977,N_4704,N_4579);
and U5978 (N_5978,N_4278,N_4223);
nor U5979 (N_5979,N_4362,N_4913);
nor U5980 (N_5980,N_4519,N_4673);
and U5981 (N_5981,N_4649,N_4724);
nand U5982 (N_5982,N_4761,N_4702);
nor U5983 (N_5983,N_4399,N_4066);
nor U5984 (N_5984,N_4925,N_4536);
and U5985 (N_5985,N_4713,N_4613);
nor U5986 (N_5986,N_4355,N_4792);
nand U5987 (N_5987,N_4130,N_4969);
or U5988 (N_5988,N_4525,N_4554);
nand U5989 (N_5989,N_4060,N_4767);
xor U5990 (N_5990,N_4836,N_4091);
nor U5991 (N_5991,N_4359,N_4384);
or U5992 (N_5992,N_4861,N_4021);
nand U5993 (N_5993,N_4853,N_4331);
or U5994 (N_5994,N_4584,N_4487);
xor U5995 (N_5995,N_4869,N_4527);
nor U5996 (N_5996,N_4778,N_4653);
nor U5997 (N_5997,N_4689,N_4064);
and U5998 (N_5998,N_4857,N_4130);
nand U5999 (N_5999,N_4519,N_4980);
nand U6000 (N_6000,N_5266,N_5260);
or U6001 (N_6001,N_5982,N_5727);
xor U6002 (N_6002,N_5544,N_5675);
and U6003 (N_6003,N_5463,N_5219);
xor U6004 (N_6004,N_5587,N_5687);
nand U6005 (N_6005,N_5865,N_5488);
xor U6006 (N_6006,N_5254,N_5674);
or U6007 (N_6007,N_5434,N_5561);
nor U6008 (N_6008,N_5791,N_5469);
xor U6009 (N_6009,N_5609,N_5740);
nand U6010 (N_6010,N_5338,N_5844);
nand U6011 (N_6011,N_5214,N_5778);
and U6012 (N_6012,N_5783,N_5101);
xor U6013 (N_6013,N_5155,N_5639);
nand U6014 (N_6014,N_5619,N_5987);
or U6015 (N_6015,N_5459,N_5978);
or U6016 (N_6016,N_5393,N_5025);
or U6017 (N_6017,N_5658,N_5610);
and U6018 (N_6018,N_5756,N_5073);
or U6019 (N_6019,N_5611,N_5672);
nand U6020 (N_6020,N_5774,N_5819);
nand U6021 (N_6021,N_5122,N_5713);
and U6022 (N_6022,N_5929,N_5663);
xnor U6023 (N_6023,N_5613,N_5557);
nand U6024 (N_6024,N_5055,N_5239);
nand U6025 (N_6025,N_5919,N_5681);
or U6026 (N_6026,N_5457,N_5837);
xor U6027 (N_6027,N_5784,N_5960);
xnor U6028 (N_6028,N_5213,N_5891);
nor U6029 (N_6029,N_5848,N_5703);
or U6030 (N_6030,N_5077,N_5066);
and U6031 (N_6031,N_5424,N_5014);
nor U6032 (N_6032,N_5976,N_5612);
and U6033 (N_6033,N_5462,N_5192);
nand U6034 (N_6034,N_5545,N_5624);
xnor U6035 (N_6035,N_5735,N_5886);
nand U6036 (N_6036,N_5645,N_5023);
or U6037 (N_6037,N_5331,N_5945);
xor U6038 (N_6038,N_5660,N_5364);
and U6039 (N_6039,N_5438,N_5707);
nor U6040 (N_6040,N_5076,N_5964);
xor U6041 (N_6041,N_5592,N_5946);
nand U6042 (N_6042,N_5177,N_5107);
nand U6043 (N_6043,N_5706,N_5975);
xnor U6044 (N_6044,N_5692,N_5882);
nand U6045 (N_6045,N_5165,N_5518);
xor U6046 (N_6046,N_5563,N_5902);
and U6047 (N_6047,N_5862,N_5597);
or U6048 (N_6048,N_5500,N_5095);
nor U6049 (N_6049,N_5845,N_5932);
nand U6050 (N_6050,N_5253,N_5303);
nor U6051 (N_6051,N_5157,N_5836);
or U6052 (N_6052,N_5661,N_5471);
or U6053 (N_6053,N_5470,N_5382);
nor U6054 (N_6054,N_5234,N_5396);
nor U6055 (N_6055,N_5069,N_5637);
xor U6056 (N_6056,N_5512,N_5598);
nand U6057 (N_6057,N_5720,N_5898);
nand U6058 (N_6058,N_5472,N_5595);
xnor U6059 (N_6059,N_5568,N_5761);
xnor U6060 (N_6060,N_5885,N_5843);
xnor U6061 (N_6061,N_5558,N_5605);
or U6062 (N_6062,N_5136,N_5638);
nor U6063 (N_6063,N_5241,N_5632);
nand U6064 (N_6064,N_5662,N_5894);
and U6065 (N_6065,N_5667,N_5256);
and U6066 (N_6066,N_5087,N_5428);
or U6067 (N_6067,N_5630,N_5496);
xnor U6068 (N_6068,N_5517,N_5020);
nor U6069 (N_6069,N_5230,N_5082);
nor U6070 (N_6070,N_5152,N_5041);
or U6071 (N_6071,N_5161,N_5896);
xnor U6072 (N_6072,N_5231,N_5944);
and U6073 (N_6073,N_5917,N_5583);
xor U6074 (N_6074,N_5410,N_5120);
nor U6075 (N_6075,N_5813,N_5402);
nand U6076 (N_6076,N_5349,N_5990);
nor U6077 (N_6077,N_5255,N_5246);
nor U6078 (N_6078,N_5388,N_5543);
and U6079 (N_6079,N_5800,N_5053);
and U6080 (N_6080,N_5655,N_5357);
or U6081 (N_6081,N_5831,N_5934);
xor U6082 (N_6082,N_5233,N_5359);
or U6083 (N_6083,N_5252,N_5133);
xor U6084 (N_6084,N_5064,N_5810);
or U6085 (N_6085,N_5763,N_5323);
or U6086 (N_6086,N_5280,N_5555);
and U6087 (N_6087,N_5940,N_5311);
and U6088 (N_6088,N_5342,N_5738);
and U6089 (N_6089,N_5447,N_5059);
nand U6090 (N_6090,N_5140,N_5038);
xnor U6091 (N_6091,N_5390,N_5981);
or U6092 (N_6092,N_5935,N_5355);
and U6093 (N_6093,N_5847,N_5730);
nor U6094 (N_6094,N_5603,N_5635);
xnor U6095 (N_6095,N_5614,N_5823);
or U6096 (N_6096,N_5374,N_5985);
and U6097 (N_6097,N_5185,N_5271);
or U6098 (N_6098,N_5356,N_5998);
xnor U6099 (N_6099,N_5754,N_5001);
nor U6100 (N_6100,N_5045,N_5283);
and U6101 (N_6101,N_5895,N_5371);
nand U6102 (N_6102,N_5086,N_5709);
nand U6103 (N_6103,N_5771,N_5273);
or U6104 (N_6104,N_5372,N_5980);
and U6105 (N_6105,N_5839,N_5593);
nand U6106 (N_6106,N_5866,N_5433);
nand U6107 (N_6107,N_5695,N_5315);
nor U6108 (N_6108,N_5552,N_5223);
nor U6109 (N_6109,N_5868,N_5261);
xnor U6110 (N_6110,N_5394,N_5979);
nor U6111 (N_6111,N_5668,N_5298);
or U6112 (N_6112,N_5006,N_5058);
xor U6113 (N_6113,N_5016,N_5292);
nor U6114 (N_6114,N_5710,N_5715);
nor U6115 (N_6115,N_5456,N_5164);
xor U6116 (N_6116,N_5248,N_5959);
xor U6117 (N_6117,N_5577,N_5135);
and U6118 (N_6118,N_5716,N_5096);
xor U6119 (N_6119,N_5251,N_5257);
nor U6120 (N_6120,N_5576,N_5536);
or U6121 (N_6121,N_5793,N_5322);
or U6122 (N_6122,N_5093,N_5907);
xor U6123 (N_6123,N_5546,N_5098);
or U6124 (N_6124,N_5967,N_5453);
xor U6125 (N_6125,N_5367,N_5790);
and U6126 (N_6126,N_5582,N_5510);
and U6127 (N_6127,N_5176,N_5770);
xor U6128 (N_6128,N_5003,N_5081);
and U6129 (N_6129,N_5739,N_5033);
or U6130 (N_6130,N_5365,N_5392);
nand U6131 (N_6131,N_5621,N_5160);
nor U6132 (N_6132,N_5785,N_5391);
nand U6133 (N_6133,N_5075,N_5103);
nor U6134 (N_6134,N_5175,N_5736);
nand U6135 (N_6135,N_5872,N_5318);
nand U6136 (N_6136,N_5262,N_5495);
nand U6137 (N_6137,N_5719,N_5201);
or U6138 (N_6138,N_5189,N_5139);
nand U6139 (N_6139,N_5397,N_5291);
nor U6140 (N_6140,N_5024,N_5431);
or U6141 (N_6141,N_5051,N_5585);
xor U6142 (N_6142,N_5869,N_5377);
and U6143 (N_6143,N_5994,N_5806);
nand U6144 (N_6144,N_5969,N_5748);
or U6145 (N_6145,N_5010,N_5207);
nor U6146 (N_6146,N_5503,N_5217);
xor U6147 (N_6147,N_5203,N_5615);
nor U6148 (N_6148,N_5767,N_5962);
xnor U6149 (N_6149,N_5194,N_5276);
or U6150 (N_6150,N_5853,N_5634);
nand U6151 (N_6151,N_5743,N_5788);
xor U6152 (N_6152,N_5851,N_5956);
nand U6153 (N_6153,N_5515,N_5700);
or U6154 (N_6154,N_5553,N_5274);
nand U6155 (N_6155,N_5955,N_5330);
or U6156 (N_6156,N_5511,N_5734);
nand U6157 (N_6157,N_5070,N_5487);
nand U6158 (N_6158,N_5329,N_5524);
nor U6159 (N_6159,N_5090,N_5924);
nand U6160 (N_6160,N_5429,N_5650);
nor U6161 (N_6161,N_5733,N_5047);
nor U6162 (N_6162,N_5494,N_5030);
xnor U6163 (N_6163,N_5308,N_5746);
nand U6164 (N_6164,N_5474,N_5646);
and U6165 (N_6165,N_5272,N_5811);
or U6166 (N_6166,N_5741,N_5640);
or U6167 (N_6167,N_5212,N_5467);
nor U6168 (N_6168,N_5893,N_5466);
or U6169 (N_6169,N_5861,N_5608);
or U6170 (N_6170,N_5590,N_5389);
nand U6171 (N_6171,N_5912,N_5123);
and U6172 (N_6172,N_5400,N_5768);
and U6173 (N_6173,N_5671,N_5921);
or U6174 (N_6174,N_5225,N_5530);
and U6175 (N_6175,N_5554,N_5285);
xnor U6176 (N_6176,N_5153,N_5972);
and U6177 (N_6177,N_5387,N_5363);
and U6178 (N_6178,N_5647,N_5776);
nand U6179 (N_6179,N_5617,N_5422);
nor U6180 (N_6180,N_5996,N_5685);
or U6181 (N_6181,N_5817,N_5012);
nand U6182 (N_6182,N_5731,N_5306);
nand U6183 (N_6183,N_5581,N_5265);
nand U6184 (N_6184,N_5501,N_5221);
or U6185 (N_6185,N_5887,N_5689);
and U6186 (N_6186,N_5297,N_5504);
or U6187 (N_6187,N_5174,N_5589);
nor U6188 (N_6188,N_5642,N_5618);
and U6189 (N_6189,N_5683,N_5973);
nor U6190 (N_6190,N_5875,N_5673);
nor U6191 (N_6191,N_5523,N_5796);
or U6192 (N_6192,N_5759,N_5247);
nor U6193 (N_6193,N_5680,N_5726);
nor U6194 (N_6194,N_5521,N_5477);
and U6195 (N_6195,N_5777,N_5398);
and U6196 (N_6196,N_5013,N_5879);
nand U6197 (N_6197,N_5369,N_5008);
nand U6198 (N_6198,N_5780,N_5729);
xnor U6199 (N_6199,N_5441,N_5295);
xnor U6200 (N_6200,N_5760,N_5749);
nor U6201 (N_6201,N_5415,N_5911);
or U6202 (N_6202,N_5953,N_5037);
nand U6203 (N_6203,N_5420,N_5999);
nand U6204 (N_6204,N_5114,N_5573);
or U6205 (N_6205,N_5325,N_5282);
xnor U6206 (N_6206,N_5017,N_5931);
xor U6207 (N_6207,N_5751,N_5278);
and U6208 (N_6208,N_5379,N_5002);
nor U6209 (N_6209,N_5682,N_5287);
nor U6210 (N_6210,N_5578,N_5159);
and U6211 (N_6211,N_5856,N_5168);
and U6212 (N_6212,N_5947,N_5240);
nor U6213 (N_6213,N_5992,N_5178);
nor U6214 (N_6214,N_5526,N_5350);
nor U6215 (N_6215,N_5316,N_5963);
or U6216 (N_6216,N_5481,N_5222);
and U6217 (N_6217,N_5307,N_5781);
nor U6218 (N_6218,N_5513,N_5057);
or U6219 (N_6219,N_5537,N_5354);
nand U6220 (N_6220,N_5850,N_5814);
nor U6221 (N_6221,N_5065,N_5732);
nor U6222 (N_6222,N_5533,N_5224);
and U6223 (N_6223,N_5901,N_5113);
nor U6224 (N_6224,N_5991,N_5294);
or U6225 (N_6225,N_5208,N_5301);
nand U6226 (N_6226,N_5275,N_5816);
nor U6227 (N_6227,N_5631,N_5300);
nand U6228 (N_6228,N_5314,N_5195);
nand U6229 (N_6229,N_5717,N_5508);
nor U6230 (N_6230,N_5607,N_5529);
xor U6231 (N_6231,N_5304,N_5188);
or U6232 (N_6232,N_5535,N_5591);
and U6233 (N_6233,N_5551,N_5421);
nor U6234 (N_6234,N_5473,N_5957);
nor U6235 (N_6235,N_5186,N_5881);
nor U6236 (N_6236,N_5840,N_5809);
nand U6237 (N_6237,N_5958,N_5403);
and U6238 (N_6238,N_5833,N_5676);
nand U6239 (N_6239,N_5797,N_5149);
nor U6240 (N_6240,N_5199,N_5211);
or U6241 (N_6241,N_5050,N_5489);
or U6242 (N_6242,N_5627,N_5099);
nor U6243 (N_6243,N_5567,N_5035);
xor U6244 (N_6244,N_5191,N_5039);
nor U6245 (N_6245,N_5779,N_5859);
and U6246 (N_6246,N_5426,N_5021);
xnor U6247 (N_6247,N_5205,N_5516);
nand U6248 (N_6248,N_5908,N_5408);
nor U6249 (N_6249,N_5599,N_5916);
xor U6250 (N_6250,N_5828,N_5444);
and U6251 (N_6251,N_5485,N_5876);
and U6252 (N_6252,N_5131,N_5337);
xor U6253 (N_6253,N_5803,N_5965);
and U6254 (N_6254,N_5029,N_5413);
or U6255 (N_6255,N_5542,N_5903);
nand U6256 (N_6256,N_5293,N_5319);
nor U6257 (N_6257,N_5401,N_5368);
xor U6258 (N_6258,N_5943,N_5118);
nand U6259 (N_6259,N_5268,N_5827);
xor U6260 (N_6260,N_5228,N_5805);
nor U6261 (N_6261,N_5666,N_5514);
xor U6262 (N_6262,N_5659,N_5183);
and U6263 (N_6263,N_5015,N_5936);
nor U6264 (N_6264,N_5063,N_5562);
nand U6265 (N_6265,N_5450,N_5725);
xnor U6266 (N_6266,N_5941,N_5137);
nor U6267 (N_6267,N_5116,N_5332);
and U6268 (N_6268,N_5430,N_5678);
or U6269 (N_6269,N_5309,N_5150);
nand U6270 (N_6270,N_5480,N_5242);
or U6271 (N_6271,N_5375,N_5712);
and U6272 (N_6272,N_5130,N_5714);
nand U6273 (N_6273,N_5154,N_5102);
or U6274 (N_6274,N_5445,N_5170);
nand U6275 (N_6275,N_5146,N_5449);
nor U6276 (N_6276,N_5011,N_5288);
nand U6277 (N_6277,N_5046,N_5616);
or U6278 (N_6278,N_5566,N_5948);
and U6279 (N_6279,N_5117,N_5920);
xnor U6280 (N_6280,N_5966,N_5302);
or U6281 (N_6281,N_5062,N_5484);
and U6282 (N_6282,N_5905,N_5547);
or U6283 (N_6283,N_5755,N_5807);
nor U6284 (N_6284,N_5718,N_5156);
or U6285 (N_6285,N_5841,N_5918);
nor U6286 (N_6286,N_5180,N_5742);
xnor U6287 (N_6287,N_5949,N_5290);
and U6288 (N_6288,N_5766,N_5060);
nand U6289 (N_6289,N_5079,N_5448);
xor U6290 (N_6290,N_5792,N_5405);
nand U6291 (N_6291,N_5344,N_5336);
and U6292 (N_6292,N_5664,N_5834);
and U6293 (N_6293,N_5572,N_5772);
xnor U6294 (N_6294,N_5009,N_5376);
and U6295 (N_6295,N_5933,N_5475);
and U6296 (N_6296,N_5412,N_5418);
or U6297 (N_6297,N_5028,N_5238);
and U6298 (N_6298,N_5343,N_5310);
nor U6299 (N_6299,N_5758,N_5830);
or U6300 (N_6300,N_5004,N_5440);
nor U6301 (N_6301,N_5381,N_5520);
xnor U6302 (N_6302,N_5145,N_5723);
nor U6303 (N_6303,N_5838,N_5928);
and U6304 (N_6304,N_5798,N_5250);
nor U6305 (N_6305,N_5702,N_5753);
xnor U6306 (N_6306,N_5550,N_5031);
or U6307 (N_6307,N_5378,N_5922);
and U6308 (N_6308,N_5083,N_5068);
xor U6309 (N_6309,N_5125,N_5427);
and U6310 (N_6310,N_5335,N_5042);
and U6311 (N_6311,N_5857,N_5395);
nand U6312 (N_6312,N_5106,N_5899);
and U6313 (N_6313,N_5799,N_5437);
or U6314 (N_6314,N_5049,N_5399);
nand U6315 (N_6315,N_5370,N_5926);
or U6316 (N_6316,N_5651,N_5822);
or U6317 (N_6317,N_5479,N_5750);
nand U6318 (N_6318,N_5386,N_5997);
and U6319 (N_6319,N_5124,N_5559);
nand U6320 (N_6320,N_5824,N_5040);
xor U6321 (N_6321,N_5166,N_5328);
and U6322 (N_6322,N_5765,N_5334);
and U6323 (N_6323,N_5032,N_5232);
or U6324 (N_6324,N_5870,N_5084);
and U6325 (N_6325,N_5313,N_5406);
or U6326 (N_6326,N_5198,N_5220);
nand U6327 (N_6327,N_5108,N_5600);
xor U6328 (N_6328,N_5100,N_5158);
and U6329 (N_6329,N_5622,N_5277);
nor U6330 (N_6330,N_5961,N_5571);
or U6331 (N_6331,N_5867,N_5643);
xor U6332 (N_6332,N_5984,N_5110);
xnor U6333 (N_6333,N_5109,N_5633);
nand U6334 (N_6334,N_5018,N_5832);
or U6335 (N_6335,N_5324,N_5476);
nand U6336 (N_6336,N_5236,N_5596);
nor U6337 (N_6337,N_5121,N_5942);
and U6338 (N_6338,N_5539,N_5854);
or U6339 (N_6339,N_5464,N_5423);
and U6340 (N_6340,N_5988,N_5132);
xnor U6341 (N_6341,N_5696,N_5148);
or U6342 (N_6342,N_5229,N_5034);
nor U6343 (N_6343,N_5801,N_5531);
nand U6344 (N_6344,N_5812,N_5482);
or U6345 (N_6345,N_5606,N_5339);
nor U6346 (N_6346,N_5134,N_5665);
nor U6347 (N_6347,N_5022,N_5089);
or U6348 (N_6348,N_5173,N_5909);
nor U6349 (N_6349,N_5721,N_5588);
xor U6350 (N_6350,N_5442,N_5877);
xor U6351 (N_6351,N_5525,N_5620);
nor U6352 (N_6352,N_5143,N_5258);
or U6353 (N_6353,N_5358,N_5200);
nor U6354 (N_6354,N_5690,N_5182);
nor U6355 (N_6355,N_5968,N_5602);
nand U6356 (N_6356,N_5362,N_5091);
and U6357 (N_6357,N_5360,N_5305);
xor U6358 (N_6358,N_5519,N_5507);
nand U6359 (N_6359,N_5452,N_5565);
nand U6360 (N_6360,N_5353,N_5569);
xor U6361 (N_6361,N_5509,N_5993);
xnor U6362 (N_6362,N_5794,N_5461);
nor U6363 (N_6363,N_5737,N_5187);
nor U6364 (N_6364,N_5915,N_5227);
and U6365 (N_6365,N_5088,N_5669);
xor U6366 (N_6366,N_5052,N_5263);
nor U6367 (N_6367,N_5204,N_5141);
and U6368 (N_6368,N_5522,N_5641);
xnor U6369 (N_6369,N_5206,N_5701);
and U6370 (N_6370,N_5216,N_5056);
or U6371 (N_6371,N_5179,N_5910);
xnor U6372 (N_6372,N_5490,N_5094);
xor U6373 (N_6373,N_5326,N_5728);
nand U6374 (N_6374,N_5871,N_5184);
xnor U6375 (N_6375,N_5863,N_5048);
or U6376 (N_6376,N_5264,N_5722);
and U6377 (N_6377,N_5939,N_5815);
or U6378 (N_6378,N_5505,N_5270);
xor U6379 (N_6379,N_5654,N_5541);
xnor U6380 (N_6380,N_5986,N_5974);
nor U6381 (N_6381,N_5534,N_5345);
or U6382 (N_6382,N_5105,N_5636);
nand U6383 (N_6383,N_5026,N_5119);
xnor U6384 (N_6384,N_5190,N_5925);
xnor U6385 (N_6385,N_5243,N_5226);
xor U6386 (N_6386,N_5686,N_5465);
or U6387 (N_6387,N_5209,N_5197);
nand U6388 (N_6388,N_5327,N_5267);
nor U6389 (N_6389,N_5970,N_5527);
or U6390 (N_6390,N_5483,N_5044);
xnor U6391 (N_6391,N_5460,N_5601);
or U6392 (N_6392,N_5938,N_5849);
and U6393 (N_6393,N_5604,N_5071);
nand U6394 (N_6394,N_5693,N_5652);
or U6395 (N_6395,N_5983,N_5147);
nand U6396 (N_6396,N_5072,N_5657);
or U6397 (N_6397,N_5584,N_5499);
xnor U6398 (N_6398,N_5027,N_5744);
or U6399 (N_6399,N_5825,N_5468);
or U6400 (N_6400,N_5906,N_5549);
xor U6401 (N_6401,N_5312,N_5128);
and U6402 (N_6402,N_5952,N_5691);
or U6403 (N_6403,N_5913,N_5679);
nor U6404 (N_6404,N_5502,N_5914);
or U6405 (N_6405,N_5829,N_5745);
nand U6406 (N_6406,N_5000,N_5846);
and U6407 (N_6407,N_5923,N_5670);
or U6408 (N_6408,N_5787,N_5889);
nand U6409 (N_6409,N_5884,N_5820);
nor U6410 (N_6410,N_5804,N_5162);
nand U6411 (N_6411,N_5129,N_5883);
or U6412 (N_6412,N_5404,N_5644);
or U6413 (N_6413,N_5900,N_5532);
and U6414 (N_6414,N_5244,N_5432);
or U6415 (N_6415,N_5172,N_5361);
xnor U6416 (N_6416,N_5142,N_5786);
and U6417 (N_6417,N_5419,N_5078);
nand U6418 (N_6418,N_5085,N_5492);
xnor U6419 (N_6419,N_5169,N_5625);
nand U6420 (N_6420,N_5711,N_5705);
and U6421 (N_6421,N_5193,N_5340);
or U6422 (N_6422,N_5491,N_5138);
and U6423 (N_6423,N_5005,N_5351);
nor U6424 (N_6424,N_5826,N_5564);
nor U6425 (N_6425,N_5210,N_5281);
or U6426 (N_6426,N_5855,N_5950);
and U6427 (N_6427,N_5486,N_5259);
nor U6428 (N_6428,N_5299,N_5384);
nand U6429 (N_6429,N_5092,N_5904);
xor U6430 (N_6430,N_5019,N_5348);
and U6431 (N_6431,N_5757,N_5628);
and U6432 (N_6432,N_5629,N_5104);
and U6433 (N_6433,N_5498,N_5575);
and U6434 (N_6434,N_5446,N_5775);
xnor U6435 (N_6435,N_5080,N_5144);
xor U6436 (N_6436,N_5373,N_5385);
nand U6437 (N_6437,N_5540,N_5127);
xor U6438 (N_6438,N_5163,N_5007);
and U6439 (N_6439,N_5808,N_5954);
or U6440 (N_6440,N_5789,N_5842);
xor U6441 (N_6441,N_5995,N_5594);
nand U6442 (N_6442,N_5296,N_5989);
nand U6443 (N_6443,N_5383,N_5880);
nor U6444 (N_6444,N_5764,N_5237);
and U6445 (N_6445,N_5317,N_5245);
nand U6446 (N_6446,N_5411,N_5126);
nor U6447 (N_6447,N_5623,N_5352);
nor U6448 (N_6448,N_5802,N_5821);
nor U6449 (N_6449,N_5435,N_5586);
nor U6450 (N_6450,N_5218,N_5858);
and U6451 (N_6451,N_5626,N_5454);
nand U6452 (N_6452,N_5697,N_5333);
and U6453 (N_6453,N_5366,N_5436);
and U6454 (N_6454,N_5115,N_5579);
or U6455 (N_6455,N_5708,N_5704);
nor U6456 (N_6456,N_5548,N_5458);
nand U6457 (N_6457,N_5407,N_5752);
or U6458 (N_6458,N_5202,N_5181);
xor U6459 (N_6459,N_5574,N_5414);
xor U6460 (N_6460,N_5528,N_5249);
and U6461 (N_6461,N_5648,N_5971);
and U6462 (N_6462,N_5688,N_5560);
nand U6463 (N_6463,N_5698,N_5782);
and U6464 (N_6464,N_5196,N_5930);
or U6465 (N_6465,N_5656,N_5416);
nand U6466 (N_6466,N_5346,N_5897);
xnor U6467 (N_6467,N_5067,N_5874);
nand U6468 (N_6468,N_5653,N_5769);
nor U6469 (N_6469,N_5892,N_5890);
or U6470 (N_6470,N_5506,N_5497);
or U6471 (N_6471,N_5269,N_5289);
and U6472 (N_6472,N_5747,N_5762);
or U6473 (N_6473,N_5538,N_5951);
nand U6474 (N_6474,N_5580,N_5493);
xnor U6475 (N_6475,N_5279,N_5036);
nand U6476 (N_6476,N_5451,N_5852);
nand U6477 (N_6477,N_5795,N_5171);
xnor U6478 (N_6478,N_5167,N_5677);
or U6479 (N_6479,N_5860,N_5347);
and U6480 (N_6480,N_5818,N_5409);
or U6481 (N_6481,N_5888,N_5556);
xor U6482 (N_6482,N_5724,N_5061);
and U6483 (N_6483,N_5864,N_5977);
or U6484 (N_6484,N_5443,N_5417);
nand U6485 (N_6485,N_5151,N_5111);
and U6486 (N_6486,N_5215,N_5043);
nor U6487 (N_6487,N_5684,N_5074);
nand U6488 (N_6488,N_5699,N_5054);
or U6489 (N_6489,N_5873,N_5694);
nor U6490 (N_6490,N_5478,N_5320);
xor U6491 (N_6491,N_5937,N_5380);
nor U6492 (N_6492,N_5649,N_5425);
xor U6493 (N_6493,N_5455,N_5570);
xor U6494 (N_6494,N_5286,N_5439);
nor U6495 (N_6495,N_5341,N_5112);
and U6496 (N_6496,N_5835,N_5284);
and U6497 (N_6497,N_5321,N_5927);
nor U6498 (N_6498,N_5773,N_5878);
and U6499 (N_6499,N_5235,N_5097);
or U6500 (N_6500,N_5536,N_5037);
and U6501 (N_6501,N_5926,N_5750);
or U6502 (N_6502,N_5120,N_5034);
or U6503 (N_6503,N_5262,N_5950);
or U6504 (N_6504,N_5987,N_5252);
nand U6505 (N_6505,N_5583,N_5629);
and U6506 (N_6506,N_5063,N_5331);
xor U6507 (N_6507,N_5454,N_5376);
or U6508 (N_6508,N_5207,N_5657);
nor U6509 (N_6509,N_5676,N_5191);
nand U6510 (N_6510,N_5657,N_5402);
and U6511 (N_6511,N_5651,N_5943);
nor U6512 (N_6512,N_5983,N_5946);
nand U6513 (N_6513,N_5363,N_5552);
xnor U6514 (N_6514,N_5382,N_5695);
and U6515 (N_6515,N_5403,N_5906);
or U6516 (N_6516,N_5475,N_5970);
nand U6517 (N_6517,N_5216,N_5764);
xnor U6518 (N_6518,N_5309,N_5655);
or U6519 (N_6519,N_5895,N_5907);
nor U6520 (N_6520,N_5286,N_5786);
xnor U6521 (N_6521,N_5375,N_5987);
xor U6522 (N_6522,N_5511,N_5227);
and U6523 (N_6523,N_5516,N_5092);
and U6524 (N_6524,N_5876,N_5657);
nor U6525 (N_6525,N_5431,N_5448);
xor U6526 (N_6526,N_5923,N_5027);
nand U6527 (N_6527,N_5590,N_5374);
and U6528 (N_6528,N_5921,N_5293);
xor U6529 (N_6529,N_5936,N_5210);
nand U6530 (N_6530,N_5057,N_5359);
nor U6531 (N_6531,N_5115,N_5226);
and U6532 (N_6532,N_5715,N_5664);
xnor U6533 (N_6533,N_5487,N_5300);
and U6534 (N_6534,N_5767,N_5761);
nor U6535 (N_6535,N_5795,N_5921);
or U6536 (N_6536,N_5043,N_5644);
nor U6537 (N_6537,N_5977,N_5530);
xor U6538 (N_6538,N_5013,N_5722);
and U6539 (N_6539,N_5955,N_5158);
and U6540 (N_6540,N_5152,N_5976);
nor U6541 (N_6541,N_5196,N_5301);
xnor U6542 (N_6542,N_5961,N_5403);
and U6543 (N_6543,N_5987,N_5918);
xnor U6544 (N_6544,N_5374,N_5129);
nand U6545 (N_6545,N_5503,N_5118);
and U6546 (N_6546,N_5469,N_5471);
nand U6547 (N_6547,N_5306,N_5534);
nor U6548 (N_6548,N_5592,N_5514);
xnor U6549 (N_6549,N_5214,N_5488);
nand U6550 (N_6550,N_5035,N_5512);
and U6551 (N_6551,N_5885,N_5348);
xor U6552 (N_6552,N_5624,N_5802);
nor U6553 (N_6553,N_5283,N_5665);
nor U6554 (N_6554,N_5212,N_5058);
and U6555 (N_6555,N_5456,N_5212);
nand U6556 (N_6556,N_5477,N_5444);
xor U6557 (N_6557,N_5373,N_5805);
xor U6558 (N_6558,N_5957,N_5665);
xor U6559 (N_6559,N_5079,N_5455);
nand U6560 (N_6560,N_5913,N_5037);
nand U6561 (N_6561,N_5986,N_5595);
or U6562 (N_6562,N_5371,N_5612);
or U6563 (N_6563,N_5797,N_5515);
nor U6564 (N_6564,N_5291,N_5317);
nand U6565 (N_6565,N_5317,N_5356);
xor U6566 (N_6566,N_5223,N_5565);
and U6567 (N_6567,N_5988,N_5247);
and U6568 (N_6568,N_5916,N_5469);
xnor U6569 (N_6569,N_5434,N_5235);
nand U6570 (N_6570,N_5291,N_5414);
xnor U6571 (N_6571,N_5149,N_5823);
and U6572 (N_6572,N_5195,N_5135);
or U6573 (N_6573,N_5164,N_5320);
nand U6574 (N_6574,N_5802,N_5106);
or U6575 (N_6575,N_5861,N_5042);
and U6576 (N_6576,N_5525,N_5075);
xnor U6577 (N_6577,N_5412,N_5625);
or U6578 (N_6578,N_5071,N_5442);
nand U6579 (N_6579,N_5555,N_5499);
and U6580 (N_6580,N_5387,N_5348);
nor U6581 (N_6581,N_5396,N_5014);
nand U6582 (N_6582,N_5711,N_5432);
xnor U6583 (N_6583,N_5514,N_5947);
nand U6584 (N_6584,N_5473,N_5173);
or U6585 (N_6585,N_5875,N_5883);
or U6586 (N_6586,N_5429,N_5569);
xor U6587 (N_6587,N_5682,N_5936);
nand U6588 (N_6588,N_5321,N_5379);
nand U6589 (N_6589,N_5083,N_5109);
and U6590 (N_6590,N_5710,N_5985);
nor U6591 (N_6591,N_5022,N_5306);
xor U6592 (N_6592,N_5272,N_5254);
or U6593 (N_6593,N_5372,N_5276);
nor U6594 (N_6594,N_5766,N_5736);
and U6595 (N_6595,N_5599,N_5105);
and U6596 (N_6596,N_5478,N_5952);
and U6597 (N_6597,N_5944,N_5862);
and U6598 (N_6598,N_5163,N_5182);
or U6599 (N_6599,N_5432,N_5933);
nor U6600 (N_6600,N_5798,N_5433);
and U6601 (N_6601,N_5425,N_5622);
nand U6602 (N_6602,N_5893,N_5282);
nor U6603 (N_6603,N_5520,N_5447);
xnor U6604 (N_6604,N_5964,N_5757);
nand U6605 (N_6605,N_5256,N_5455);
nor U6606 (N_6606,N_5255,N_5741);
xnor U6607 (N_6607,N_5552,N_5965);
nor U6608 (N_6608,N_5376,N_5825);
nor U6609 (N_6609,N_5944,N_5949);
and U6610 (N_6610,N_5182,N_5463);
xnor U6611 (N_6611,N_5617,N_5332);
and U6612 (N_6612,N_5952,N_5720);
xnor U6613 (N_6613,N_5819,N_5192);
and U6614 (N_6614,N_5014,N_5066);
or U6615 (N_6615,N_5743,N_5883);
nor U6616 (N_6616,N_5528,N_5870);
and U6617 (N_6617,N_5884,N_5934);
nand U6618 (N_6618,N_5194,N_5780);
nand U6619 (N_6619,N_5205,N_5808);
nor U6620 (N_6620,N_5514,N_5118);
nor U6621 (N_6621,N_5150,N_5509);
and U6622 (N_6622,N_5860,N_5119);
xnor U6623 (N_6623,N_5800,N_5310);
or U6624 (N_6624,N_5526,N_5848);
xor U6625 (N_6625,N_5306,N_5639);
or U6626 (N_6626,N_5390,N_5545);
nor U6627 (N_6627,N_5929,N_5306);
xor U6628 (N_6628,N_5982,N_5415);
and U6629 (N_6629,N_5373,N_5658);
xor U6630 (N_6630,N_5736,N_5087);
or U6631 (N_6631,N_5868,N_5981);
nand U6632 (N_6632,N_5574,N_5753);
nor U6633 (N_6633,N_5265,N_5110);
xnor U6634 (N_6634,N_5128,N_5619);
and U6635 (N_6635,N_5320,N_5255);
or U6636 (N_6636,N_5360,N_5329);
nor U6637 (N_6637,N_5724,N_5869);
and U6638 (N_6638,N_5188,N_5362);
xnor U6639 (N_6639,N_5512,N_5749);
or U6640 (N_6640,N_5498,N_5209);
nor U6641 (N_6641,N_5325,N_5882);
xor U6642 (N_6642,N_5611,N_5052);
or U6643 (N_6643,N_5394,N_5464);
xnor U6644 (N_6644,N_5988,N_5067);
or U6645 (N_6645,N_5916,N_5083);
nor U6646 (N_6646,N_5868,N_5742);
nor U6647 (N_6647,N_5888,N_5833);
xor U6648 (N_6648,N_5338,N_5262);
nand U6649 (N_6649,N_5654,N_5545);
nor U6650 (N_6650,N_5879,N_5378);
or U6651 (N_6651,N_5274,N_5004);
or U6652 (N_6652,N_5719,N_5757);
nand U6653 (N_6653,N_5946,N_5941);
and U6654 (N_6654,N_5974,N_5838);
or U6655 (N_6655,N_5135,N_5626);
or U6656 (N_6656,N_5200,N_5334);
or U6657 (N_6657,N_5137,N_5891);
and U6658 (N_6658,N_5673,N_5608);
nor U6659 (N_6659,N_5360,N_5363);
nor U6660 (N_6660,N_5874,N_5472);
nand U6661 (N_6661,N_5308,N_5991);
nand U6662 (N_6662,N_5975,N_5470);
nor U6663 (N_6663,N_5262,N_5028);
nor U6664 (N_6664,N_5445,N_5411);
or U6665 (N_6665,N_5706,N_5384);
xor U6666 (N_6666,N_5480,N_5980);
nand U6667 (N_6667,N_5869,N_5865);
nor U6668 (N_6668,N_5469,N_5770);
nand U6669 (N_6669,N_5297,N_5471);
xor U6670 (N_6670,N_5736,N_5950);
nor U6671 (N_6671,N_5270,N_5776);
nor U6672 (N_6672,N_5276,N_5592);
nor U6673 (N_6673,N_5896,N_5446);
nor U6674 (N_6674,N_5433,N_5956);
nand U6675 (N_6675,N_5551,N_5216);
and U6676 (N_6676,N_5770,N_5143);
xor U6677 (N_6677,N_5609,N_5508);
or U6678 (N_6678,N_5611,N_5871);
xor U6679 (N_6679,N_5108,N_5904);
xor U6680 (N_6680,N_5744,N_5885);
xor U6681 (N_6681,N_5120,N_5325);
xnor U6682 (N_6682,N_5832,N_5655);
and U6683 (N_6683,N_5390,N_5498);
or U6684 (N_6684,N_5929,N_5351);
nand U6685 (N_6685,N_5415,N_5405);
nor U6686 (N_6686,N_5225,N_5365);
and U6687 (N_6687,N_5294,N_5591);
nand U6688 (N_6688,N_5418,N_5245);
nand U6689 (N_6689,N_5270,N_5113);
xnor U6690 (N_6690,N_5559,N_5916);
nand U6691 (N_6691,N_5588,N_5069);
nor U6692 (N_6692,N_5711,N_5520);
nand U6693 (N_6693,N_5367,N_5931);
xor U6694 (N_6694,N_5633,N_5951);
nand U6695 (N_6695,N_5928,N_5398);
or U6696 (N_6696,N_5050,N_5863);
nor U6697 (N_6697,N_5511,N_5137);
or U6698 (N_6698,N_5785,N_5234);
and U6699 (N_6699,N_5167,N_5959);
and U6700 (N_6700,N_5180,N_5184);
xor U6701 (N_6701,N_5316,N_5616);
nor U6702 (N_6702,N_5876,N_5044);
xor U6703 (N_6703,N_5754,N_5646);
and U6704 (N_6704,N_5885,N_5020);
nor U6705 (N_6705,N_5340,N_5274);
nand U6706 (N_6706,N_5865,N_5833);
xnor U6707 (N_6707,N_5500,N_5289);
or U6708 (N_6708,N_5959,N_5049);
and U6709 (N_6709,N_5527,N_5741);
or U6710 (N_6710,N_5651,N_5868);
nor U6711 (N_6711,N_5403,N_5641);
nor U6712 (N_6712,N_5427,N_5107);
nand U6713 (N_6713,N_5123,N_5752);
or U6714 (N_6714,N_5102,N_5391);
or U6715 (N_6715,N_5637,N_5580);
nand U6716 (N_6716,N_5360,N_5025);
nand U6717 (N_6717,N_5011,N_5846);
xnor U6718 (N_6718,N_5831,N_5725);
nand U6719 (N_6719,N_5584,N_5790);
nor U6720 (N_6720,N_5309,N_5099);
nand U6721 (N_6721,N_5493,N_5960);
or U6722 (N_6722,N_5191,N_5255);
nor U6723 (N_6723,N_5313,N_5058);
xor U6724 (N_6724,N_5799,N_5613);
nand U6725 (N_6725,N_5925,N_5033);
nor U6726 (N_6726,N_5434,N_5522);
xor U6727 (N_6727,N_5475,N_5642);
xnor U6728 (N_6728,N_5475,N_5882);
or U6729 (N_6729,N_5422,N_5454);
or U6730 (N_6730,N_5254,N_5153);
or U6731 (N_6731,N_5013,N_5211);
and U6732 (N_6732,N_5127,N_5519);
or U6733 (N_6733,N_5277,N_5942);
nand U6734 (N_6734,N_5554,N_5204);
nor U6735 (N_6735,N_5409,N_5776);
and U6736 (N_6736,N_5901,N_5560);
xor U6737 (N_6737,N_5129,N_5994);
nand U6738 (N_6738,N_5805,N_5583);
nand U6739 (N_6739,N_5149,N_5195);
and U6740 (N_6740,N_5406,N_5453);
and U6741 (N_6741,N_5944,N_5567);
nand U6742 (N_6742,N_5967,N_5785);
nand U6743 (N_6743,N_5138,N_5348);
or U6744 (N_6744,N_5660,N_5462);
nand U6745 (N_6745,N_5515,N_5858);
and U6746 (N_6746,N_5152,N_5742);
nand U6747 (N_6747,N_5738,N_5639);
or U6748 (N_6748,N_5663,N_5095);
xnor U6749 (N_6749,N_5417,N_5735);
and U6750 (N_6750,N_5206,N_5580);
or U6751 (N_6751,N_5851,N_5630);
or U6752 (N_6752,N_5032,N_5451);
and U6753 (N_6753,N_5802,N_5773);
and U6754 (N_6754,N_5800,N_5006);
nand U6755 (N_6755,N_5263,N_5711);
nor U6756 (N_6756,N_5695,N_5953);
and U6757 (N_6757,N_5475,N_5256);
nor U6758 (N_6758,N_5480,N_5173);
nand U6759 (N_6759,N_5415,N_5384);
or U6760 (N_6760,N_5565,N_5905);
nand U6761 (N_6761,N_5945,N_5554);
xnor U6762 (N_6762,N_5186,N_5244);
nor U6763 (N_6763,N_5744,N_5381);
nand U6764 (N_6764,N_5959,N_5142);
or U6765 (N_6765,N_5760,N_5853);
nor U6766 (N_6766,N_5384,N_5410);
nand U6767 (N_6767,N_5488,N_5215);
and U6768 (N_6768,N_5301,N_5313);
nand U6769 (N_6769,N_5270,N_5836);
nand U6770 (N_6770,N_5338,N_5860);
nor U6771 (N_6771,N_5326,N_5508);
nor U6772 (N_6772,N_5983,N_5559);
nand U6773 (N_6773,N_5403,N_5768);
or U6774 (N_6774,N_5486,N_5630);
and U6775 (N_6775,N_5833,N_5018);
and U6776 (N_6776,N_5431,N_5524);
and U6777 (N_6777,N_5652,N_5181);
nor U6778 (N_6778,N_5502,N_5711);
and U6779 (N_6779,N_5868,N_5055);
nor U6780 (N_6780,N_5066,N_5991);
or U6781 (N_6781,N_5819,N_5615);
nor U6782 (N_6782,N_5849,N_5540);
and U6783 (N_6783,N_5357,N_5345);
nand U6784 (N_6784,N_5730,N_5452);
nor U6785 (N_6785,N_5385,N_5088);
or U6786 (N_6786,N_5109,N_5098);
and U6787 (N_6787,N_5929,N_5468);
or U6788 (N_6788,N_5784,N_5370);
xnor U6789 (N_6789,N_5039,N_5721);
nand U6790 (N_6790,N_5030,N_5923);
nor U6791 (N_6791,N_5441,N_5705);
nor U6792 (N_6792,N_5309,N_5698);
or U6793 (N_6793,N_5701,N_5370);
nand U6794 (N_6794,N_5151,N_5226);
and U6795 (N_6795,N_5467,N_5772);
and U6796 (N_6796,N_5750,N_5298);
xnor U6797 (N_6797,N_5083,N_5873);
and U6798 (N_6798,N_5841,N_5420);
xnor U6799 (N_6799,N_5412,N_5345);
and U6800 (N_6800,N_5601,N_5921);
xnor U6801 (N_6801,N_5325,N_5108);
and U6802 (N_6802,N_5767,N_5674);
nand U6803 (N_6803,N_5068,N_5013);
nor U6804 (N_6804,N_5634,N_5366);
nor U6805 (N_6805,N_5248,N_5826);
xnor U6806 (N_6806,N_5778,N_5879);
nand U6807 (N_6807,N_5364,N_5249);
nand U6808 (N_6808,N_5582,N_5736);
nand U6809 (N_6809,N_5248,N_5919);
and U6810 (N_6810,N_5738,N_5813);
or U6811 (N_6811,N_5889,N_5646);
nor U6812 (N_6812,N_5862,N_5708);
or U6813 (N_6813,N_5892,N_5534);
xnor U6814 (N_6814,N_5741,N_5256);
nor U6815 (N_6815,N_5912,N_5962);
nor U6816 (N_6816,N_5613,N_5860);
xor U6817 (N_6817,N_5217,N_5940);
nor U6818 (N_6818,N_5600,N_5792);
xnor U6819 (N_6819,N_5440,N_5124);
nand U6820 (N_6820,N_5933,N_5834);
and U6821 (N_6821,N_5609,N_5966);
and U6822 (N_6822,N_5697,N_5885);
or U6823 (N_6823,N_5379,N_5733);
xor U6824 (N_6824,N_5549,N_5442);
xnor U6825 (N_6825,N_5531,N_5971);
xor U6826 (N_6826,N_5052,N_5470);
nand U6827 (N_6827,N_5286,N_5167);
nor U6828 (N_6828,N_5350,N_5599);
nor U6829 (N_6829,N_5959,N_5905);
or U6830 (N_6830,N_5373,N_5834);
nor U6831 (N_6831,N_5325,N_5721);
nor U6832 (N_6832,N_5734,N_5092);
nor U6833 (N_6833,N_5258,N_5655);
xor U6834 (N_6834,N_5463,N_5663);
or U6835 (N_6835,N_5373,N_5914);
or U6836 (N_6836,N_5236,N_5923);
nor U6837 (N_6837,N_5058,N_5323);
or U6838 (N_6838,N_5226,N_5599);
nor U6839 (N_6839,N_5224,N_5677);
or U6840 (N_6840,N_5594,N_5239);
nand U6841 (N_6841,N_5568,N_5339);
and U6842 (N_6842,N_5447,N_5333);
or U6843 (N_6843,N_5049,N_5285);
nand U6844 (N_6844,N_5811,N_5010);
nand U6845 (N_6845,N_5470,N_5665);
xor U6846 (N_6846,N_5468,N_5320);
nor U6847 (N_6847,N_5209,N_5049);
and U6848 (N_6848,N_5863,N_5848);
and U6849 (N_6849,N_5600,N_5404);
xor U6850 (N_6850,N_5431,N_5883);
nor U6851 (N_6851,N_5910,N_5153);
nor U6852 (N_6852,N_5270,N_5219);
nand U6853 (N_6853,N_5276,N_5830);
or U6854 (N_6854,N_5364,N_5471);
or U6855 (N_6855,N_5442,N_5561);
nor U6856 (N_6856,N_5785,N_5188);
xor U6857 (N_6857,N_5272,N_5455);
xor U6858 (N_6858,N_5174,N_5745);
xor U6859 (N_6859,N_5354,N_5964);
nand U6860 (N_6860,N_5154,N_5469);
xnor U6861 (N_6861,N_5644,N_5793);
and U6862 (N_6862,N_5660,N_5472);
nor U6863 (N_6863,N_5495,N_5440);
nor U6864 (N_6864,N_5193,N_5259);
or U6865 (N_6865,N_5372,N_5212);
xor U6866 (N_6866,N_5078,N_5541);
or U6867 (N_6867,N_5620,N_5200);
xnor U6868 (N_6868,N_5397,N_5670);
and U6869 (N_6869,N_5876,N_5079);
xnor U6870 (N_6870,N_5365,N_5023);
or U6871 (N_6871,N_5665,N_5593);
and U6872 (N_6872,N_5212,N_5416);
or U6873 (N_6873,N_5146,N_5458);
or U6874 (N_6874,N_5522,N_5262);
nor U6875 (N_6875,N_5767,N_5233);
nand U6876 (N_6876,N_5008,N_5001);
or U6877 (N_6877,N_5301,N_5589);
and U6878 (N_6878,N_5668,N_5635);
or U6879 (N_6879,N_5854,N_5198);
and U6880 (N_6880,N_5251,N_5688);
or U6881 (N_6881,N_5772,N_5409);
or U6882 (N_6882,N_5551,N_5366);
xnor U6883 (N_6883,N_5817,N_5812);
nand U6884 (N_6884,N_5498,N_5100);
nor U6885 (N_6885,N_5333,N_5930);
nand U6886 (N_6886,N_5360,N_5814);
nand U6887 (N_6887,N_5584,N_5254);
nand U6888 (N_6888,N_5927,N_5465);
xor U6889 (N_6889,N_5954,N_5292);
nand U6890 (N_6890,N_5794,N_5373);
and U6891 (N_6891,N_5038,N_5935);
and U6892 (N_6892,N_5540,N_5992);
xnor U6893 (N_6893,N_5681,N_5777);
and U6894 (N_6894,N_5419,N_5947);
nand U6895 (N_6895,N_5717,N_5651);
nand U6896 (N_6896,N_5280,N_5196);
and U6897 (N_6897,N_5332,N_5417);
nand U6898 (N_6898,N_5632,N_5543);
and U6899 (N_6899,N_5047,N_5568);
or U6900 (N_6900,N_5284,N_5649);
nand U6901 (N_6901,N_5906,N_5907);
xor U6902 (N_6902,N_5274,N_5487);
nor U6903 (N_6903,N_5686,N_5325);
nor U6904 (N_6904,N_5020,N_5469);
nor U6905 (N_6905,N_5305,N_5441);
xnor U6906 (N_6906,N_5501,N_5675);
nand U6907 (N_6907,N_5465,N_5976);
or U6908 (N_6908,N_5088,N_5910);
xnor U6909 (N_6909,N_5291,N_5637);
or U6910 (N_6910,N_5733,N_5525);
or U6911 (N_6911,N_5787,N_5267);
or U6912 (N_6912,N_5890,N_5352);
or U6913 (N_6913,N_5103,N_5025);
nand U6914 (N_6914,N_5713,N_5947);
xnor U6915 (N_6915,N_5197,N_5383);
or U6916 (N_6916,N_5233,N_5698);
nor U6917 (N_6917,N_5411,N_5985);
and U6918 (N_6918,N_5988,N_5694);
xor U6919 (N_6919,N_5088,N_5410);
or U6920 (N_6920,N_5693,N_5115);
nand U6921 (N_6921,N_5104,N_5558);
nand U6922 (N_6922,N_5079,N_5498);
or U6923 (N_6923,N_5600,N_5077);
xor U6924 (N_6924,N_5012,N_5982);
nand U6925 (N_6925,N_5664,N_5765);
nand U6926 (N_6926,N_5068,N_5736);
or U6927 (N_6927,N_5393,N_5052);
and U6928 (N_6928,N_5451,N_5158);
or U6929 (N_6929,N_5001,N_5818);
and U6930 (N_6930,N_5212,N_5692);
or U6931 (N_6931,N_5969,N_5479);
xor U6932 (N_6932,N_5136,N_5503);
or U6933 (N_6933,N_5585,N_5251);
and U6934 (N_6934,N_5623,N_5020);
nand U6935 (N_6935,N_5749,N_5778);
xnor U6936 (N_6936,N_5985,N_5600);
xnor U6937 (N_6937,N_5274,N_5524);
xor U6938 (N_6938,N_5573,N_5935);
xnor U6939 (N_6939,N_5299,N_5823);
xnor U6940 (N_6940,N_5460,N_5059);
xnor U6941 (N_6941,N_5082,N_5136);
nor U6942 (N_6942,N_5560,N_5282);
and U6943 (N_6943,N_5678,N_5107);
or U6944 (N_6944,N_5186,N_5891);
and U6945 (N_6945,N_5998,N_5891);
or U6946 (N_6946,N_5123,N_5272);
and U6947 (N_6947,N_5960,N_5965);
or U6948 (N_6948,N_5091,N_5106);
and U6949 (N_6949,N_5923,N_5836);
nor U6950 (N_6950,N_5650,N_5292);
nand U6951 (N_6951,N_5734,N_5356);
xnor U6952 (N_6952,N_5248,N_5451);
xor U6953 (N_6953,N_5818,N_5732);
or U6954 (N_6954,N_5712,N_5728);
nand U6955 (N_6955,N_5158,N_5124);
nand U6956 (N_6956,N_5891,N_5595);
or U6957 (N_6957,N_5689,N_5608);
and U6958 (N_6958,N_5415,N_5471);
nand U6959 (N_6959,N_5263,N_5438);
and U6960 (N_6960,N_5232,N_5930);
or U6961 (N_6961,N_5910,N_5953);
and U6962 (N_6962,N_5775,N_5455);
xor U6963 (N_6963,N_5470,N_5320);
xnor U6964 (N_6964,N_5796,N_5732);
and U6965 (N_6965,N_5503,N_5125);
nand U6966 (N_6966,N_5052,N_5035);
and U6967 (N_6967,N_5698,N_5574);
nor U6968 (N_6968,N_5199,N_5288);
xor U6969 (N_6969,N_5508,N_5307);
or U6970 (N_6970,N_5819,N_5629);
xnor U6971 (N_6971,N_5742,N_5917);
xor U6972 (N_6972,N_5261,N_5707);
nor U6973 (N_6973,N_5467,N_5746);
or U6974 (N_6974,N_5172,N_5309);
nand U6975 (N_6975,N_5103,N_5669);
or U6976 (N_6976,N_5456,N_5774);
nand U6977 (N_6977,N_5673,N_5219);
xnor U6978 (N_6978,N_5943,N_5477);
or U6979 (N_6979,N_5126,N_5896);
and U6980 (N_6980,N_5858,N_5875);
and U6981 (N_6981,N_5416,N_5075);
nand U6982 (N_6982,N_5185,N_5652);
and U6983 (N_6983,N_5458,N_5121);
xor U6984 (N_6984,N_5089,N_5860);
nand U6985 (N_6985,N_5288,N_5900);
nand U6986 (N_6986,N_5021,N_5023);
nand U6987 (N_6987,N_5420,N_5944);
and U6988 (N_6988,N_5720,N_5076);
and U6989 (N_6989,N_5159,N_5413);
and U6990 (N_6990,N_5927,N_5233);
nor U6991 (N_6991,N_5028,N_5393);
xnor U6992 (N_6992,N_5724,N_5059);
nand U6993 (N_6993,N_5788,N_5414);
nor U6994 (N_6994,N_5181,N_5266);
xor U6995 (N_6995,N_5068,N_5304);
or U6996 (N_6996,N_5276,N_5142);
nand U6997 (N_6997,N_5257,N_5394);
and U6998 (N_6998,N_5337,N_5313);
nor U6999 (N_6999,N_5735,N_5754);
or U7000 (N_7000,N_6002,N_6830);
nor U7001 (N_7001,N_6884,N_6901);
nand U7002 (N_7002,N_6091,N_6766);
nor U7003 (N_7003,N_6859,N_6338);
nand U7004 (N_7004,N_6512,N_6806);
and U7005 (N_7005,N_6336,N_6845);
and U7006 (N_7006,N_6122,N_6580);
xor U7007 (N_7007,N_6063,N_6049);
nor U7008 (N_7008,N_6251,N_6904);
xor U7009 (N_7009,N_6218,N_6438);
nor U7010 (N_7010,N_6761,N_6378);
or U7011 (N_7011,N_6341,N_6790);
nor U7012 (N_7012,N_6804,N_6750);
xor U7013 (N_7013,N_6763,N_6756);
and U7014 (N_7014,N_6616,N_6801);
nor U7015 (N_7015,N_6227,N_6686);
and U7016 (N_7016,N_6235,N_6943);
and U7017 (N_7017,N_6453,N_6687);
or U7018 (N_7018,N_6044,N_6051);
xor U7019 (N_7019,N_6427,N_6493);
or U7020 (N_7020,N_6148,N_6070);
xor U7021 (N_7021,N_6082,N_6005);
or U7022 (N_7022,N_6641,N_6660);
nand U7023 (N_7023,N_6244,N_6624);
and U7024 (N_7024,N_6054,N_6732);
xnor U7025 (N_7025,N_6899,N_6452);
or U7026 (N_7026,N_6062,N_6665);
or U7027 (N_7027,N_6929,N_6572);
and U7028 (N_7028,N_6131,N_6179);
nor U7029 (N_7029,N_6422,N_6673);
or U7030 (N_7030,N_6089,N_6731);
xnor U7031 (N_7031,N_6596,N_6125);
and U7032 (N_7032,N_6510,N_6282);
or U7033 (N_7033,N_6000,N_6206);
nor U7034 (N_7034,N_6600,N_6780);
xor U7035 (N_7035,N_6772,N_6306);
or U7036 (N_7036,N_6412,N_6886);
or U7037 (N_7037,N_6808,N_6141);
and U7038 (N_7038,N_6429,N_6987);
or U7039 (N_7039,N_6822,N_6875);
xor U7040 (N_7040,N_6507,N_6531);
nand U7041 (N_7041,N_6551,N_6670);
nand U7042 (N_7042,N_6405,N_6802);
and U7043 (N_7043,N_6966,N_6021);
or U7044 (N_7044,N_6478,N_6649);
nand U7045 (N_7045,N_6116,N_6284);
or U7046 (N_7046,N_6721,N_6432);
or U7047 (N_7047,N_6667,N_6240);
xnor U7048 (N_7048,N_6560,N_6525);
and U7049 (N_7049,N_6029,N_6204);
nor U7050 (N_7050,N_6094,N_6826);
xor U7051 (N_7051,N_6949,N_6158);
or U7052 (N_7052,N_6781,N_6150);
xor U7053 (N_7053,N_6272,N_6487);
nand U7054 (N_7054,N_6498,N_6417);
nor U7055 (N_7055,N_6410,N_6855);
and U7056 (N_7056,N_6085,N_6898);
xor U7057 (N_7057,N_6164,N_6080);
nor U7058 (N_7058,N_6605,N_6523);
nand U7059 (N_7059,N_6132,N_6144);
xor U7060 (N_7060,N_6773,N_6267);
nand U7061 (N_7061,N_6952,N_6262);
or U7062 (N_7062,N_6046,N_6757);
nand U7063 (N_7063,N_6746,N_6215);
and U7064 (N_7064,N_6947,N_6858);
and U7065 (N_7065,N_6574,N_6443);
or U7066 (N_7066,N_6703,N_6888);
nand U7067 (N_7067,N_6540,N_6851);
or U7068 (N_7068,N_6355,N_6546);
and U7069 (N_7069,N_6389,N_6294);
or U7070 (N_7070,N_6327,N_6839);
nand U7071 (N_7071,N_6558,N_6367);
nor U7072 (N_7072,N_6798,N_6118);
nand U7073 (N_7073,N_6878,N_6123);
nor U7074 (N_7074,N_6575,N_6059);
or U7075 (N_7075,N_6375,N_6400);
and U7076 (N_7076,N_6717,N_6060);
or U7077 (N_7077,N_6393,N_6360);
nand U7078 (N_7078,N_6979,N_6351);
xor U7079 (N_7079,N_6248,N_6800);
and U7080 (N_7080,N_6807,N_6101);
nand U7081 (N_7081,N_6787,N_6543);
xor U7082 (N_7082,N_6014,N_6301);
nand U7083 (N_7083,N_6853,N_6057);
nor U7084 (N_7084,N_6997,N_6145);
nand U7085 (N_7085,N_6106,N_6147);
nand U7086 (N_7086,N_6892,N_6420);
or U7087 (N_7087,N_6461,N_6208);
nor U7088 (N_7088,N_6406,N_6399);
xnor U7089 (N_7089,N_6656,N_6936);
xor U7090 (N_7090,N_6491,N_6706);
xor U7091 (N_7091,N_6096,N_6725);
and U7092 (N_7092,N_6371,N_6231);
and U7093 (N_7093,N_6197,N_6447);
xor U7094 (N_7094,N_6727,N_6829);
and U7095 (N_7095,N_6205,N_6786);
or U7096 (N_7096,N_6212,N_6981);
and U7097 (N_7097,N_6922,N_6648);
and U7098 (N_7098,N_6545,N_6710);
nor U7099 (N_7099,N_6916,N_6597);
nor U7100 (N_7100,N_6494,N_6562);
nand U7101 (N_7101,N_6277,N_6303);
nand U7102 (N_7102,N_6458,N_6852);
and U7103 (N_7103,N_6401,N_6655);
or U7104 (N_7104,N_6891,N_6874);
and U7105 (N_7105,N_6496,N_6905);
nand U7106 (N_7106,N_6637,N_6521);
or U7107 (N_7107,N_6941,N_6921);
and U7108 (N_7108,N_6867,N_6250);
and U7109 (N_7109,N_6102,N_6549);
and U7110 (N_7110,N_6996,N_6349);
nor U7111 (N_7111,N_6174,N_6236);
or U7112 (N_7112,N_6634,N_6926);
or U7113 (N_7113,N_6832,N_6245);
or U7114 (N_7114,N_6455,N_6473);
or U7115 (N_7115,N_6503,N_6961);
xnor U7116 (N_7116,N_6838,N_6385);
and U7117 (N_7117,N_6362,N_6735);
nand U7118 (N_7118,N_6121,N_6486);
nand U7119 (N_7119,N_6099,N_6210);
nand U7120 (N_7120,N_6998,N_6739);
nand U7121 (N_7121,N_6189,N_6668);
or U7122 (N_7122,N_6103,N_6664);
or U7123 (N_7123,N_6975,N_6843);
and U7124 (N_7124,N_6568,N_6237);
xor U7125 (N_7125,N_6595,N_6639);
nand U7126 (N_7126,N_6752,N_6383);
nand U7127 (N_7127,N_6069,N_6659);
xor U7128 (N_7128,N_6456,N_6482);
xnor U7129 (N_7129,N_6199,N_6940);
or U7130 (N_7130,N_6434,N_6675);
and U7131 (N_7131,N_6329,N_6618);
xnor U7132 (N_7132,N_6439,N_6469);
nor U7133 (N_7133,N_6354,N_6733);
and U7134 (N_7134,N_6226,N_6918);
or U7135 (N_7135,N_6071,N_6421);
xor U7136 (N_7136,N_6317,N_6139);
nor U7137 (N_7137,N_6599,N_6713);
nor U7138 (N_7138,N_6372,N_6247);
and U7139 (N_7139,N_6304,N_6740);
nor U7140 (N_7140,N_6969,N_6514);
xor U7141 (N_7141,N_6586,N_6584);
xnor U7142 (N_7142,N_6366,N_6948);
and U7143 (N_7143,N_6479,N_6423);
nor U7144 (N_7144,N_6263,N_6516);
xor U7145 (N_7145,N_6187,N_6462);
or U7146 (N_7146,N_6965,N_6047);
nor U7147 (N_7147,N_6913,N_6024);
nor U7148 (N_7148,N_6956,N_6292);
xnor U7149 (N_7149,N_6844,N_6261);
nand U7150 (N_7150,N_6223,N_6022);
nor U7151 (N_7151,N_6065,N_6636);
or U7152 (N_7152,N_6632,N_6993);
nor U7153 (N_7153,N_6138,N_6692);
or U7154 (N_7154,N_6621,N_6955);
or U7155 (N_7155,N_6629,N_6353);
or U7156 (N_7156,N_6056,N_6459);
nor U7157 (N_7157,N_6774,N_6419);
xor U7158 (N_7158,N_6533,N_6862);
and U7159 (N_7159,N_6885,N_6849);
and U7160 (N_7160,N_6296,N_6184);
nand U7161 (N_7161,N_6255,N_6676);
nor U7162 (N_7162,N_6477,N_6426);
nand U7163 (N_7163,N_6048,N_6652);
or U7164 (N_7164,N_6445,N_6391);
and U7165 (N_7165,N_6127,N_6093);
nor U7166 (N_7166,N_6111,N_6760);
or U7167 (N_7167,N_6628,N_6492);
xor U7168 (N_7168,N_6934,N_6522);
nor U7169 (N_7169,N_6741,N_6887);
and U7170 (N_7170,N_6620,N_6009);
xor U7171 (N_7171,N_6217,N_6475);
and U7172 (N_7172,N_6869,N_6027);
nand U7173 (N_7173,N_6889,N_6151);
or U7174 (N_7174,N_6571,N_6992);
or U7175 (N_7175,N_6092,N_6754);
and U7176 (N_7176,N_6015,N_6192);
xor U7177 (N_7177,N_6428,N_6819);
nor U7178 (N_7178,N_6042,N_6974);
or U7179 (N_7179,N_6895,N_6182);
nand U7180 (N_7180,N_6700,N_6359);
and U7181 (N_7181,N_6079,N_6058);
nand U7182 (N_7182,N_6016,N_6407);
or U7183 (N_7183,N_6257,N_6409);
nand U7184 (N_7184,N_6333,N_6191);
or U7185 (N_7185,N_6097,N_6561);
nor U7186 (N_7186,N_6076,N_6645);
nand U7187 (N_7187,N_6809,N_6653);
nor U7188 (N_7188,N_6394,N_6075);
xnor U7189 (N_7189,N_6290,N_6534);
or U7190 (N_7190,N_6113,N_6414);
xor U7191 (N_7191,N_6064,N_6081);
nor U7192 (N_7192,N_6630,N_6542);
and U7193 (N_7193,N_6134,N_6601);
and U7194 (N_7194,N_6654,N_6509);
nor U7195 (N_7195,N_6666,N_6638);
and U7196 (N_7196,N_6977,N_6203);
or U7197 (N_7197,N_6074,N_6988);
nor U7198 (N_7198,N_6007,N_6814);
nor U7199 (N_7199,N_6990,N_6045);
xor U7200 (N_7200,N_6034,N_6332);
and U7201 (N_7201,N_6233,N_6072);
nor U7202 (N_7202,N_6825,N_6963);
and U7203 (N_7203,N_6538,N_6457);
or U7204 (N_7204,N_6175,N_6281);
or U7205 (N_7205,N_6382,N_6036);
and U7206 (N_7206,N_6249,N_6611);
nand U7207 (N_7207,N_6403,N_6488);
or U7208 (N_7208,N_6931,N_6622);
and U7209 (N_7209,N_6124,N_6791);
nor U7210 (N_7210,N_6026,N_6265);
xnor U7211 (N_7211,N_6915,N_6536);
or U7212 (N_7212,N_6017,N_6783);
nor U7213 (N_7213,N_6982,N_6377);
nor U7214 (N_7214,N_6361,N_6490);
nand U7215 (N_7215,N_6577,N_6315);
nor U7216 (N_7216,N_6052,N_6278);
and U7217 (N_7217,N_6755,N_6954);
xnor U7218 (N_7218,N_6326,N_6207);
nand U7219 (N_7219,N_6310,N_6860);
and U7220 (N_7220,N_6865,N_6195);
nor U7221 (N_7221,N_6003,N_6300);
xnor U7222 (N_7222,N_6381,N_6827);
nor U7223 (N_7223,N_6778,N_6923);
xnor U7224 (N_7224,N_6770,N_6006);
nand U7225 (N_7225,N_6927,N_6751);
nor U7226 (N_7226,N_6155,N_6817);
xnor U7227 (N_7227,N_6243,N_6345);
and U7228 (N_7228,N_6681,N_6815);
nand U7229 (N_7229,N_6643,N_6259);
xnor U7230 (N_7230,N_6866,N_6095);
and U7231 (N_7231,N_6004,N_6685);
and U7232 (N_7232,N_6769,N_6672);
nand U7233 (N_7233,N_6087,N_6900);
and U7234 (N_7234,N_6232,N_6133);
nand U7235 (N_7235,N_6818,N_6626);
nand U7236 (N_7236,N_6258,N_6989);
nand U7237 (N_7237,N_6820,N_6214);
nand U7238 (N_7238,N_6796,N_6610);
or U7239 (N_7239,N_6962,N_6433);
nor U7240 (N_7240,N_6152,N_6154);
and U7241 (N_7241,N_6502,N_6376);
and U7242 (N_7242,N_6854,N_6168);
nor U7243 (N_7243,N_6167,N_6472);
and U7244 (N_7244,N_6220,N_6734);
and U7245 (N_7245,N_6368,N_6030);
nor U7246 (N_7246,N_6607,N_6526);
or U7247 (N_7247,N_6759,N_6454);
xnor U7248 (N_7248,N_6909,N_6912);
nand U7249 (N_7249,N_6719,N_6928);
nor U7250 (N_7250,N_6485,N_6194);
nor U7251 (N_7251,N_6318,N_6025);
xor U7252 (N_7252,N_6951,N_6067);
xnor U7253 (N_7253,N_6178,N_6295);
xnor U7254 (N_7254,N_6567,N_6117);
or U7255 (N_7255,N_6569,N_6505);
nor U7256 (N_7256,N_6877,N_6983);
xnor U7257 (N_7257,N_6906,N_6841);
or U7258 (N_7258,N_6484,N_6444);
or U7259 (N_7259,N_6229,N_6120);
and U7260 (N_7260,N_6209,N_6861);
nand U7261 (N_7261,N_6553,N_6720);
nand U7262 (N_7262,N_6647,N_6019);
nand U7263 (N_7263,N_6991,N_6441);
nand U7264 (N_7264,N_6728,N_6716);
nor U7265 (N_7265,N_6663,N_6615);
nor U7266 (N_7266,N_6784,N_6999);
nor U7267 (N_7267,N_6779,N_6153);
nand U7268 (N_7268,N_6169,N_6548);
nor U7269 (N_7269,N_6038,N_6810);
and U7270 (N_7270,N_6631,N_6451);
nand U7271 (N_7271,N_6564,N_6312);
xor U7272 (N_7272,N_6448,N_6342);
or U7273 (N_7273,N_6186,N_6471);
nand U7274 (N_7274,N_6264,N_6890);
nor U7275 (N_7275,N_6390,N_6320);
or U7276 (N_7276,N_6321,N_6379);
nand U7277 (N_7277,N_6785,N_6344);
xnor U7278 (N_7278,N_6911,N_6749);
nor U7279 (N_7279,N_6463,N_6268);
nor U7280 (N_7280,N_6253,N_6691);
xnor U7281 (N_7281,N_6520,N_6748);
and U7282 (N_7282,N_6340,N_6633);
and U7283 (N_7283,N_6589,N_6689);
and U7284 (N_7284,N_6397,N_6744);
or U7285 (N_7285,N_6346,N_6246);
nand U7286 (N_7286,N_6925,N_6585);
and U7287 (N_7287,N_6657,N_6055);
or U7288 (N_7288,N_6130,N_6537);
or U7289 (N_7289,N_6709,N_6722);
and U7290 (N_7290,N_6945,N_6950);
nand U7291 (N_7291,N_6010,N_6322);
nand U7292 (N_7292,N_6797,N_6782);
xnor U7293 (N_7293,N_6316,N_6881);
and U7294 (N_7294,N_6856,N_6411);
nand U7295 (N_7295,N_6053,N_6946);
nor U7296 (N_7296,N_6930,N_6697);
nor U7297 (N_7297,N_6588,N_6933);
xnor U7298 (N_7298,N_6698,N_6163);
or U7299 (N_7299,N_6324,N_6061);
or U7300 (N_7300,N_6793,N_6413);
and U7301 (N_7301,N_6373,N_6957);
nor U7302 (N_7302,N_6662,N_6557);
and U7303 (N_7303,N_6959,N_6870);
nand U7304 (N_7304,N_6651,N_6280);
nor U7305 (N_7305,N_6374,N_6497);
nor U7306 (N_7306,N_6500,N_6938);
or U7307 (N_7307,N_6224,N_6114);
xor U7308 (N_7308,N_6529,N_6742);
xnor U7309 (N_7309,N_6984,N_6335);
or U7310 (N_7310,N_6581,N_6446);
nand U7311 (N_7311,N_6041,N_6582);
xor U7312 (N_7312,N_6550,N_6978);
nand U7313 (N_7313,N_6105,N_6724);
and U7314 (N_7314,N_6180,N_6971);
and U7315 (N_7315,N_6813,N_6225);
nor U7316 (N_7316,N_6970,N_6942);
and U7317 (N_7317,N_6291,N_6960);
nand U7318 (N_7318,N_6894,N_6532);
nor U7319 (N_7319,N_6398,N_6623);
and U7320 (N_7320,N_6298,N_6937);
and U7321 (N_7321,N_6254,N_6098);
or U7322 (N_7322,N_6824,N_6823);
or U7323 (N_7323,N_6834,N_6518);
and U7324 (N_7324,N_6598,N_6068);
xor U7325 (N_7325,N_6392,N_6614);
and U7326 (N_7326,N_6435,N_6402);
nor U7327 (N_7327,N_6684,N_6216);
and U7328 (N_7328,N_6539,N_6967);
nand U7329 (N_7329,N_6704,N_6573);
xnor U7330 (N_7330,N_6450,N_6776);
or U7331 (N_7331,N_6256,N_6837);
nor U7332 (N_7332,N_6994,N_6736);
xnor U7333 (N_7333,N_6812,N_6530);
nand U7334 (N_7334,N_6508,N_6811);
and U7335 (N_7335,N_6415,N_6271);
or U7336 (N_7336,N_6188,N_6213);
nand U7337 (N_7337,N_6679,N_6260);
xnor U7338 (N_7338,N_6805,N_6517);
or U7339 (N_7339,N_6711,N_6737);
or U7340 (N_7340,N_6302,N_6602);
and U7341 (N_7341,N_6020,N_6501);
and U7342 (N_7342,N_6307,N_6897);
nand U7343 (N_7343,N_6460,N_6680);
or U7344 (N_7344,N_6701,N_6768);
xor U7345 (N_7345,N_6356,N_6464);
xor U7346 (N_7346,N_6288,N_6129);
nand U7347 (N_7347,N_6476,N_6836);
nand U7348 (N_7348,N_6939,N_6831);
and U7349 (N_7349,N_6050,N_6077);
and U7350 (N_7350,N_6495,N_6857);
and U7351 (N_7351,N_6640,N_6241);
nor U7352 (N_7352,N_6544,N_6995);
and U7353 (N_7353,N_6185,N_6771);
or U7354 (N_7354,N_6747,N_6364);
nor U7355 (N_7355,N_6847,N_6730);
or U7356 (N_7356,N_6788,N_6088);
nor U7357 (N_7357,N_6115,N_6160);
xnor U7358 (N_7358,N_6384,N_6350);
or U7359 (N_7359,N_6699,N_6201);
nor U7360 (N_7360,N_6033,N_6363);
xnor U7361 (N_7361,N_6323,N_6430);
or U7362 (N_7362,N_6576,N_6142);
or U7363 (N_7363,N_6156,N_6850);
or U7364 (N_7364,N_6674,N_6882);
nand U7365 (N_7365,N_6313,N_6176);
nor U7366 (N_7366,N_6985,N_6425);
and U7367 (N_7367,N_6126,N_6149);
xor U7368 (N_7368,N_6396,N_6308);
and U7369 (N_7369,N_6011,N_6172);
xor U7370 (N_7370,N_6489,N_6579);
nor U7371 (N_7371,N_6031,N_6694);
nand U7372 (N_7372,N_6339,N_6416);
nand U7373 (N_7373,N_6273,N_6696);
xor U7374 (N_7374,N_6297,N_6506);
and U7375 (N_7375,N_6683,N_6563);
nor U7376 (N_7376,N_6789,N_6758);
xor U7377 (N_7377,N_6466,N_6863);
nor U7378 (N_7378,N_6157,N_6729);
xor U7379 (N_7379,N_6775,N_6541);
or U7380 (N_7380,N_6792,N_6876);
xnor U7381 (N_7381,N_6196,N_6166);
nand U7382 (N_7382,N_6726,N_6879);
nor U7383 (N_7383,N_6404,N_6222);
nand U7384 (N_7384,N_6309,N_6380);
nand U7385 (N_7385,N_6617,N_6910);
nand U7386 (N_7386,N_6535,N_6591);
nor U7387 (N_7387,N_6883,N_6872);
and U7388 (N_7388,N_6436,N_6840);
nor U7389 (N_7389,N_6953,N_6110);
or U7390 (N_7390,N_6480,N_6128);
nor U7391 (N_7391,N_6604,N_6183);
and U7392 (N_7392,N_6311,N_6715);
xnor U7393 (N_7393,N_6504,N_6593);
or U7394 (N_7394,N_6334,N_6973);
xnor U7395 (N_7395,N_6644,N_6012);
and U7396 (N_7396,N_6762,N_6159);
or U7397 (N_7397,N_6465,N_6609);
nor U7398 (N_7398,N_6743,N_6028);
nor U7399 (N_7399,N_6037,N_6283);
xor U7400 (N_7400,N_6107,N_6442);
nor U7401 (N_7401,N_6864,N_6669);
or U7402 (N_7402,N_6221,N_6279);
nand U7403 (N_7403,N_6986,N_6100);
nand U7404 (N_7404,N_6499,N_6470);
and U7405 (N_7405,N_6357,N_6627);
xor U7406 (N_7406,N_6200,N_6109);
nor U7407 (N_7407,N_6902,N_6606);
nor U7408 (N_7408,N_6924,N_6958);
nor U7409 (N_7409,N_6305,N_6695);
nor U7410 (N_7410,N_6370,N_6202);
xnor U7411 (N_7411,N_6893,N_6707);
and U7412 (N_7412,N_6424,N_6833);
and U7413 (N_7413,N_6515,N_6777);
or U7414 (N_7414,N_6682,N_6646);
xor U7415 (N_7415,N_6702,N_6013);
xnor U7416 (N_7416,N_6619,N_6583);
or U7417 (N_7417,N_6972,N_6570);
nor U7418 (N_7418,N_6964,N_6745);
xor U7419 (N_7419,N_6285,N_6086);
nand U7420 (N_7420,N_6040,N_6348);
or U7421 (N_7421,N_6635,N_6252);
nor U7422 (N_7422,N_6347,N_6868);
and U7423 (N_7423,N_6511,N_6119);
nand U7424 (N_7424,N_6299,N_6211);
and U7425 (N_7425,N_6968,N_6608);
xor U7426 (N_7426,N_6143,N_6903);
nand U7427 (N_7427,N_6330,N_6828);
or U7428 (N_7428,N_6043,N_6270);
nor U7429 (N_7429,N_6039,N_6590);
nand U7430 (N_7430,N_6980,N_6035);
or U7431 (N_7431,N_6481,N_6896);
and U7432 (N_7432,N_6880,N_6276);
xor U7433 (N_7433,N_6613,N_6873);
nor U7434 (N_7434,N_6181,N_6935);
or U7435 (N_7435,N_6919,N_6198);
nand U7436 (N_7436,N_6688,N_6519);
nor U7437 (N_7437,N_6678,N_6528);
and U7438 (N_7438,N_6555,N_6112);
nor U7439 (N_7439,N_6848,N_6642);
nand U7440 (N_7440,N_6140,N_6556);
xor U7441 (N_7441,N_6431,N_6136);
or U7442 (N_7442,N_6908,N_6578);
or U7443 (N_7443,N_6083,N_6708);
nor U7444 (N_7444,N_6846,N_6712);
and U7445 (N_7445,N_6944,N_6816);
nand U7446 (N_7446,N_6269,N_6765);
nor U7447 (N_7447,N_6387,N_6337);
or U7448 (N_7448,N_6932,N_6907);
nor U7449 (N_7449,N_6266,N_6177);
xnor U7450 (N_7450,N_6803,N_6976);
or U7451 (N_7451,N_6594,N_6723);
or U7452 (N_7452,N_6032,N_6565);
and U7453 (N_7453,N_6483,N_6871);
or U7454 (N_7454,N_6238,N_6078);
nor U7455 (N_7455,N_6650,N_6690);
and U7456 (N_7456,N_6314,N_6671);
xnor U7457 (N_7457,N_6161,N_6275);
nand U7458 (N_7458,N_6474,N_6554);
nor U7459 (N_7459,N_6239,N_6625);
and U7460 (N_7460,N_6714,N_6705);
and U7461 (N_7461,N_6418,N_6795);
xnor U7462 (N_7462,N_6524,N_6821);
and U7463 (N_7463,N_6001,N_6234);
nand U7464 (N_7464,N_6592,N_6547);
xnor U7465 (N_7465,N_6319,N_6343);
nor U7466 (N_7466,N_6603,N_6799);
and U7467 (N_7467,N_6440,N_6173);
xnor U7468 (N_7468,N_6328,N_6146);
xnor U7469 (N_7469,N_6612,N_6293);
xnor U7470 (N_7470,N_6108,N_6193);
nor U7471 (N_7471,N_6219,N_6171);
or U7472 (N_7472,N_6917,N_6661);
nor U7473 (N_7473,N_6437,N_6228);
nor U7474 (N_7474,N_6325,N_6835);
nand U7475 (N_7475,N_6467,N_6023);
xor U7476 (N_7476,N_6162,N_6914);
and U7477 (N_7477,N_6718,N_6365);
or U7478 (N_7478,N_6794,N_6090);
and U7479 (N_7479,N_6527,N_6920);
and U7480 (N_7480,N_6287,N_6066);
or U7481 (N_7481,N_6513,N_6289);
nand U7482 (N_7482,N_6388,N_6677);
or U7483 (N_7483,N_6693,N_6764);
xor U7484 (N_7484,N_6286,N_6468);
and U7485 (N_7485,N_6767,N_6104);
or U7486 (N_7486,N_6587,N_6552);
and U7487 (N_7487,N_6230,N_6170);
nor U7488 (N_7488,N_6008,N_6842);
nand U7489 (N_7489,N_6753,N_6449);
or U7490 (N_7490,N_6073,N_6352);
and U7491 (N_7491,N_6190,N_6242);
and U7492 (N_7492,N_6084,N_6738);
or U7493 (N_7493,N_6559,N_6395);
and U7494 (N_7494,N_6165,N_6274);
xnor U7495 (N_7495,N_6358,N_6566);
nand U7496 (N_7496,N_6369,N_6658);
nand U7497 (N_7497,N_6408,N_6018);
nor U7498 (N_7498,N_6137,N_6135);
nor U7499 (N_7499,N_6386,N_6331);
nand U7500 (N_7500,N_6552,N_6081);
nor U7501 (N_7501,N_6300,N_6576);
or U7502 (N_7502,N_6064,N_6489);
xor U7503 (N_7503,N_6589,N_6940);
xnor U7504 (N_7504,N_6590,N_6691);
nor U7505 (N_7505,N_6365,N_6230);
or U7506 (N_7506,N_6436,N_6500);
or U7507 (N_7507,N_6778,N_6235);
or U7508 (N_7508,N_6251,N_6898);
xor U7509 (N_7509,N_6595,N_6052);
nor U7510 (N_7510,N_6979,N_6452);
or U7511 (N_7511,N_6913,N_6154);
and U7512 (N_7512,N_6725,N_6582);
nor U7513 (N_7513,N_6299,N_6061);
and U7514 (N_7514,N_6818,N_6892);
nand U7515 (N_7515,N_6428,N_6436);
and U7516 (N_7516,N_6223,N_6919);
xor U7517 (N_7517,N_6990,N_6154);
nor U7518 (N_7518,N_6655,N_6387);
or U7519 (N_7519,N_6820,N_6523);
or U7520 (N_7520,N_6169,N_6208);
and U7521 (N_7521,N_6684,N_6471);
xnor U7522 (N_7522,N_6467,N_6360);
nor U7523 (N_7523,N_6371,N_6227);
nor U7524 (N_7524,N_6536,N_6586);
xnor U7525 (N_7525,N_6393,N_6192);
nor U7526 (N_7526,N_6209,N_6653);
or U7527 (N_7527,N_6414,N_6745);
or U7528 (N_7528,N_6353,N_6800);
or U7529 (N_7529,N_6830,N_6172);
or U7530 (N_7530,N_6951,N_6260);
nor U7531 (N_7531,N_6190,N_6079);
and U7532 (N_7532,N_6989,N_6953);
and U7533 (N_7533,N_6934,N_6537);
and U7534 (N_7534,N_6442,N_6540);
nand U7535 (N_7535,N_6034,N_6375);
xnor U7536 (N_7536,N_6348,N_6927);
nor U7537 (N_7537,N_6068,N_6690);
and U7538 (N_7538,N_6079,N_6371);
nand U7539 (N_7539,N_6276,N_6348);
nor U7540 (N_7540,N_6622,N_6829);
nand U7541 (N_7541,N_6733,N_6248);
nand U7542 (N_7542,N_6202,N_6122);
xor U7543 (N_7543,N_6815,N_6891);
nor U7544 (N_7544,N_6130,N_6954);
nand U7545 (N_7545,N_6085,N_6452);
nand U7546 (N_7546,N_6635,N_6407);
xor U7547 (N_7547,N_6757,N_6145);
nand U7548 (N_7548,N_6720,N_6039);
nor U7549 (N_7549,N_6489,N_6338);
and U7550 (N_7550,N_6618,N_6498);
xor U7551 (N_7551,N_6212,N_6226);
or U7552 (N_7552,N_6884,N_6154);
and U7553 (N_7553,N_6208,N_6601);
xnor U7554 (N_7554,N_6208,N_6584);
xor U7555 (N_7555,N_6188,N_6241);
and U7556 (N_7556,N_6801,N_6174);
or U7557 (N_7557,N_6460,N_6823);
nor U7558 (N_7558,N_6792,N_6559);
nor U7559 (N_7559,N_6049,N_6882);
xor U7560 (N_7560,N_6878,N_6881);
or U7561 (N_7561,N_6765,N_6746);
and U7562 (N_7562,N_6618,N_6278);
and U7563 (N_7563,N_6401,N_6812);
and U7564 (N_7564,N_6855,N_6649);
and U7565 (N_7565,N_6661,N_6188);
nor U7566 (N_7566,N_6536,N_6860);
or U7567 (N_7567,N_6251,N_6658);
xor U7568 (N_7568,N_6953,N_6322);
nand U7569 (N_7569,N_6001,N_6802);
or U7570 (N_7570,N_6519,N_6535);
nor U7571 (N_7571,N_6778,N_6493);
nor U7572 (N_7572,N_6984,N_6439);
xnor U7573 (N_7573,N_6158,N_6952);
or U7574 (N_7574,N_6752,N_6770);
and U7575 (N_7575,N_6759,N_6745);
or U7576 (N_7576,N_6623,N_6817);
nor U7577 (N_7577,N_6686,N_6830);
nand U7578 (N_7578,N_6386,N_6956);
and U7579 (N_7579,N_6668,N_6236);
xnor U7580 (N_7580,N_6864,N_6748);
or U7581 (N_7581,N_6570,N_6111);
nor U7582 (N_7582,N_6260,N_6163);
and U7583 (N_7583,N_6085,N_6758);
nand U7584 (N_7584,N_6069,N_6669);
nand U7585 (N_7585,N_6024,N_6303);
xnor U7586 (N_7586,N_6109,N_6724);
xor U7587 (N_7587,N_6706,N_6278);
or U7588 (N_7588,N_6195,N_6220);
and U7589 (N_7589,N_6706,N_6321);
nand U7590 (N_7590,N_6529,N_6389);
nand U7591 (N_7591,N_6612,N_6127);
nor U7592 (N_7592,N_6662,N_6930);
xor U7593 (N_7593,N_6312,N_6675);
xnor U7594 (N_7594,N_6913,N_6512);
nand U7595 (N_7595,N_6920,N_6927);
and U7596 (N_7596,N_6471,N_6290);
or U7597 (N_7597,N_6997,N_6382);
xor U7598 (N_7598,N_6686,N_6792);
xnor U7599 (N_7599,N_6387,N_6173);
nor U7600 (N_7600,N_6766,N_6404);
xor U7601 (N_7601,N_6100,N_6072);
and U7602 (N_7602,N_6700,N_6776);
nand U7603 (N_7603,N_6062,N_6349);
nor U7604 (N_7604,N_6951,N_6952);
xor U7605 (N_7605,N_6759,N_6894);
and U7606 (N_7606,N_6154,N_6814);
xnor U7607 (N_7607,N_6903,N_6473);
and U7608 (N_7608,N_6725,N_6562);
nor U7609 (N_7609,N_6471,N_6783);
nor U7610 (N_7610,N_6159,N_6596);
or U7611 (N_7611,N_6959,N_6639);
and U7612 (N_7612,N_6018,N_6790);
nor U7613 (N_7613,N_6812,N_6807);
xor U7614 (N_7614,N_6488,N_6943);
or U7615 (N_7615,N_6316,N_6011);
and U7616 (N_7616,N_6124,N_6660);
or U7617 (N_7617,N_6947,N_6606);
nor U7618 (N_7618,N_6914,N_6651);
and U7619 (N_7619,N_6982,N_6909);
and U7620 (N_7620,N_6289,N_6387);
nor U7621 (N_7621,N_6446,N_6116);
nor U7622 (N_7622,N_6565,N_6449);
nand U7623 (N_7623,N_6377,N_6659);
nor U7624 (N_7624,N_6189,N_6489);
and U7625 (N_7625,N_6896,N_6138);
xnor U7626 (N_7626,N_6896,N_6472);
nor U7627 (N_7627,N_6014,N_6738);
and U7628 (N_7628,N_6531,N_6485);
nand U7629 (N_7629,N_6733,N_6948);
nand U7630 (N_7630,N_6279,N_6879);
nor U7631 (N_7631,N_6858,N_6388);
or U7632 (N_7632,N_6987,N_6968);
nor U7633 (N_7633,N_6852,N_6586);
nor U7634 (N_7634,N_6634,N_6981);
xnor U7635 (N_7635,N_6631,N_6076);
or U7636 (N_7636,N_6259,N_6115);
nand U7637 (N_7637,N_6069,N_6263);
nor U7638 (N_7638,N_6445,N_6787);
or U7639 (N_7639,N_6781,N_6071);
nor U7640 (N_7640,N_6343,N_6829);
or U7641 (N_7641,N_6445,N_6479);
or U7642 (N_7642,N_6686,N_6581);
xnor U7643 (N_7643,N_6663,N_6126);
xnor U7644 (N_7644,N_6691,N_6812);
and U7645 (N_7645,N_6281,N_6028);
nand U7646 (N_7646,N_6604,N_6654);
nand U7647 (N_7647,N_6812,N_6740);
xnor U7648 (N_7648,N_6866,N_6048);
nor U7649 (N_7649,N_6130,N_6050);
nand U7650 (N_7650,N_6934,N_6945);
and U7651 (N_7651,N_6805,N_6883);
nor U7652 (N_7652,N_6419,N_6224);
nor U7653 (N_7653,N_6853,N_6874);
and U7654 (N_7654,N_6423,N_6525);
nand U7655 (N_7655,N_6964,N_6179);
nand U7656 (N_7656,N_6325,N_6650);
nor U7657 (N_7657,N_6931,N_6558);
nor U7658 (N_7658,N_6598,N_6779);
and U7659 (N_7659,N_6271,N_6709);
xnor U7660 (N_7660,N_6575,N_6394);
xnor U7661 (N_7661,N_6746,N_6817);
and U7662 (N_7662,N_6981,N_6421);
and U7663 (N_7663,N_6854,N_6546);
nand U7664 (N_7664,N_6030,N_6120);
xor U7665 (N_7665,N_6474,N_6813);
or U7666 (N_7666,N_6148,N_6350);
nor U7667 (N_7667,N_6787,N_6122);
or U7668 (N_7668,N_6867,N_6477);
or U7669 (N_7669,N_6841,N_6944);
nand U7670 (N_7670,N_6584,N_6506);
or U7671 (N_7671,N_6423,N_6371);
or U7672 (N_7672,N_6111,N_6027);
nand U7673 (N_7673,N_6387,N_6032);
xnor U7674 (N_7674,N_6722,N_6893);
xor U7675 (N_7675,N_6426,N_6835);
and U7676 (N_7676,N_6536,N_6888);
nor U7677 (N_7677,N_6515,N_6809);
nor U7678 (N_7678,N_6789,N_6112);
nor U7679 (N_7679,N_6184,N_6359);
xnor U7680 (N_7680,N_6235,N_6200);
and U7681 (N_7681,N_6691,N_6814);
nand U7682 (N_7682,N_6960,N_6719);
xnor U7683 (N_7683,N_6709,N_6626);
nand U7684 (N_7684,N_6780,N_6882);
or U7685 (N_7685,N_6911,N_6529);
xnor U7686 (N_7686,N_6877,N_6701);
nand U7687 (N_7687,N_6160,N_6910);
nor U7688 (N_7688,N_6906,N_6080);
nand U7689 (N_7689,N_6433,N_6304);
nand U7690 (N_7690,N_6898,N_6633);
nand U7691 (N_7691,N_6492,N_6320);
nand U7692 (N_7692,N_6360,N_6547);
or U7693 (N_7693,N_6459,N_6920);
and U7694 (N_7694,N_6840,N_6515);
xnor U7695 (N_7695,N_6599,N_6746);
nor U7696 (N_7696,N_6615,N_6950);
nor U7697 (N_7697,N_6595,N_6177);
xor U7698 (N_7698,N_6743,N_6557);
xor U7699 (N_7699,N_6191,N_6276);
nand U7700 (N_7700,N_6098,N_6837);
or U7701 (N_7701,N_6343,N_6514);
nand U7702 (N_7702,N_6288,N_6623);
nor U7703 (N_7703,N_6349,N_6482);
nor U7704 (N_7704,N_6382,N_6489);
or U7705 (N_7705,N_6252,N_6200);
xor U7706 (N_7706,N_6162,N_6011);
xnor U7707 (N_7707,N_6763,N_6249);
and U7708 (N_7708,N_6426,N_6841);
nor U7709 (N_7709,N_6883,N_6313);
or U7710 (N_7710,N_6044,N_6043);
and U7711 (N_7711,N_6973,N_6710);
and U7712 (N_7712,N_6680,N_6428);
and U7713 (N_7713,N_6770,N_6262);
nand U7714 (N_7714,N_6601,N_6032);
xor U7715 (N_7715,N_6208,N_6799);
nor U7716 (N_7716,N_6755,N_6218);
and U7717 (N_7717,N_6659,N_6269);
xnor U7718 (N_7718,N_6731,N_6138);
nor U7719 (N_7719,N_6481,N_6665);
nand U7720 (N_7720,N_6108,N_6107);
and U7721 (N_7721,N_6557,N_6780);
nand U7722 (N_7722,N_6438,N_6030);
or U7723 (N_7723,N_6817,N_6232);
and U7724 (N_7724,N_6624,N_6838);
nor U7725 (N_7725,N_6502,N_6144);
nand U7726 (N_7726,N_6768,N_6106);
xor U7727 (N_7727,N_6419,N_6734);
and U7728 (N_7728,N_6861,N_6149);
nor U7729 (N_7729,N_6862,N_6066);
nand U7730 (N_7730,N_6776,N_6939);
or U7731 (N_7731,N_6885,N_6135);
xor U7732 (N_7732,N_6616,N_6706);
and U7733 (N_7733,N_6890,N_6646);
nor U7734 (N_7734,N_6068,N_6390);
nor U7735 (N_7735,N_6998,N_6963);
xnor U7736 (N_7736,N_6769,N_6939);
or U7737 (N_7737,N_6336,N_6760);
nor U7738 (N_7738,N_6817,N_6854);
nand U7739 (N_7739,N_6636,N_6183);
nor U7740 (N_7740,N_6689,N_6078);
or U7741 (N_7741,N_6906,N_6527);
xor U7742 (N_7742,N_6798,N_6200);
nor U7743 (N_7743,N_6204,N_6749);
or U7744 (N_7744,N_6720,N_6733);
nand U7745 (N_7745,N_6301,N_6365);
xor U7746 (N_7746,N_6591,N_6460);
and U7747 (N_7747,N_6572,N_6890);
or U7748 (N_7748,N_6526,N_6041);
xor U7749 (N_7749,N_6510,N_6964);
or U7750 (N_7750,N_6041,N_6131);
or U7751 (N_7751,N_6784,N_6232);
nor U7752 (N_7752,N_6818,N_6874);
and U7753 (N_7753,N_6398,N_6039);
xor U7754 (N_7754,N_6324,N_6526);
nand U7755 (N_7755,N_6384,N_6969);
nor U7756 (N_7756,N_6186,N_6142);
nor U7757 (N_7757,N_6474,N_6853);
and U7758 (N_7758,N_6537,N_6344);
nand U7759 (N_7759,N_6645,N_6127);
nor U7760 (N_7760,N_6220,N_6477);
and U7761 (N_7761,N_6417,N_6961);
and U7762 (N_7762,N_6815,N_6489);
nor U7763 (N_7763,N_6873,N_6335);
or U7764 (N_7764,N_6568,N_6072);
nand U7765 (N_7765,N_6352,N_6480);
and U7766 (N_7766,N_6680,N_6820);
or U7767 (N_7767,N_6938,N_6161);
and U7768 (N_7768,N_6000,N_6866);
xor U7769 (N_7769,N_6404,N_6584);
or U7770 (N_7770,N_6416,N_6212);
and U7771 (N_7771,N_6975,N_6974);
or U7772 (N_7772,N_6280,N_6510);
nor U7773 (N_7773,N_6929,N_6661);
xor U7774 (N_7774,N_6614,N_6328);
xnor U7775 (N_7775,N_6756,N_6197);
xor U7776 (N_7776,N_6908,N_6071);
nor U7777 (N_7777,N_6133,N_6942);
and U7778 (N_7778,N_6064,N_6956);
and U7779 (N_7779,N_6619,N_6184);
and U7780 (N_7780,N_6363,N_6837);
xor U7781 (N_7781,N_6144,N_6336);
and U7782 (N_7782,N_6253,N_6102);
or U7783 (N_7783,N_6844,N_6764);
or U7784 (N_7784,N_6645,N_6865);
nand U7785 (N_7785,N_6735,N_6084);
xnor U7786 (N_7786,N_6598,N_6921);
and U7787 (N_7787,N_6001,N_6107);
or U7788 (N_7788,N_6188,N_6910);
nor U7789 (N_7789,N_6623,N_6242);
nor U7790 (N_7790,N_6895,N_6288);
nor U7791 (N_7791,N_6042,N_6059);
or U7792 (N_7792,N_6855,N_6549);
nor U7793 (N_7793,N_6706,N_6403);
nor U7794 (N_7794,N_6024,N_6765);
nor U7795 (N_7795,N_6286,N_6068);
nand U7796 (N_7796,N_6402,N_6359);
or U7797 (N_7797,N_6804,N_6792);
or U7798 (N_7798,N_6536,N_6680);
nand U7799 (N_7799,N_6382,N_6981);
and U7800 (N_7800,N_6323,N_6477);
and U7801 (N_7801,N_6460,N_6022);
nor U7802 (N_7802,N_6284,N_6892);
or U7803 (N_7803,N_6457,N_6549);
and U7804 (N_7804,N_6898,N_6656);
nand U7805 (N_7805,N_6878,N_6966);
xnor U7806 (N_7806,N_6346,N_6201);
xor U7807 (N_7807,N_6179,N_6177);
xor U7808 (N_7808,N_6058,N_6450);
nand U7809 (N_7809,N_6185,N_6980);
and U7810 (N_7810,N_6109,N_6624);
nor U7811 (N_7811,N_6257,N_6582);
nand U7812 (N_7812,N_6472,N_6432);
nor U7813 (N_7813,N_6219,N_6812);
or U7814 (N_7814,N_6067,N_6153);
nand U7815 (N_7815,N_6121,N_6664);
and U7816 (N_7816,N_6452,N_6530);
nor U7817 (N_7817,N_6079,N_6099);
nor U7818 (N_7818,N_6001,N_6858);
and U7819 (N_7819,N_6918,N_6429);
and U7820 (N_7820,N_6949,N_6175);
nor U7821 (N_7821,N_6971,N_6689);
or U7822 (N_7822,N_6545,N_6045);
xnor U7823 (N_7823,N_6518,N_6237);
and U7824 (N_7824,N_6229,N_6598);
and U7825 (N_7825,N_6867,N_6855);
nor U7826 (N_7826,N_6579,N_6714);
nor U7827 (N_7827,N_6158,N_6879);
nor U7828 (N_7828,N_6651,N_6065);
and U7829 (N_7829,N_6347,N_6129);
or U7830 (N_7830,N_6210,N_6450);
and U7831 (N_7831,N_6983,N_6112);
nor U7832 (N_7832,N_6554,N_6034);
xor U7833 (N_7833,N_6161,N_6607);
nor U7834 (N_7834,N_6220,N_6369);
nor U7835 (N_7835,N_6303,N_6290);
or U7836 (N_7836,N_6595,N_6735);
nor U7837 (N_7837,N_6339,N_6273);
and U7838 (N_7838,N_6747,N_6394);
and U7839 (N_7839,N_6611,N_6951);
or U7840 (N_7840,N_6992,N_6491);
nor U7841 (N_7841,N_6366,N_6173);
nor U7842 (N_7842,N_6358,N_6128);
nand U7843 (N_7843,N_6562,N_6902);
or U7844 (N_7844,N_6854,N_6190);
nand U7845 (N_7845,N_6602,N_6514);
nor U7846 (N_7846,N_6363,N_6260);
nor U7847 (N_7847,N_6114,N_6137);
nor U7848 (N_7848,N_6701,N_6989);
or U7849 (N_7849,N_6773,N_6246);
and U7850 (N_7850,N_6635,N_6023);
nor U7851 (N_7851,N_6159,N_6347);
or U7852 (N_7852,N_6831,N_6677);
nand U7853 (N_7853,N_6647,N_6055);
and U7854 (N_7854,N_6542,N_6930);
and U7855 (N_7855,N_6356,N_6507);
xnor U7856 (N_7856,N_6653,N_6913);
or U7857 (N_7857,N_6233,N_6112);
and U7858 (N_7858,N_6845,N_6394);
or U7859 (N_7859,N_6337,N_6513);
xor U7860 (N_7860,N_6937,N_6956);
and U7861 (N_7861,N_6930,N_6185);
nor U7862 (N_7862,N_6972,N_6862);
nand U7863 (N_7863,N_6699,N_6820);
nor U7864 (N_7864,N_6027,N_6952);
xor U7865 (N_7865,N_6730,N_6810);
nor U7866 (N_7866,N_6651,N_6584);
and U7867 (N_7867,N_6773,N_6671);
nand U7868 (N_7868,N_6670,N_6348);
nor U7869 (N_7869,N_6902,N_6578);
xnor U7870 (N_7870,N_6916,N_6140);
and U7871 (N_7871,N_6734,N_6956);
nand U7872 (N_7872,N_6245,N_6845);
nand U7873 (N_7873,N_6133,N_6049);
or U7874 (N_7874,N_6706,N_6928);
or U7875 (N_7875,N_6779,N_6190);
nand U7876 (N_7876,N_6335,N_6851);
and U7877 (N_7877,N_6007,N_6044);
nor U7878 (N_7878,N_6471,N_6970);
xor U7879 (N_7879,N_6738,N_6366);
nor U7880 (N_7880,N_6303,N_6351);
and U7881 (N_7881,N_6247,N_6977);
and U7882 (N_7882,N_6665,N_6689);
xnor U7883 (N_7883,N_6816,N_6859);
nand U7884 (N_7884,N_6038,N_6432);
nor U7885 (N_7885,N_6984,N_6949);
or U7886 (N_7886,N_6092,N_6382);
nand U7887 (N_7887,N_6887,N_6916);
xor U7888 (N_7888,N_6082,N_6088);
nor U7889 (N_7889,N_6692,N_6108);
xnor U7890 (N_7890,N_6485,N_6777);
and U7891 (N_7891,N_6506,N_6136);
nand U7892 (N_7892,N_6117,N_6153);
and U7893 (N_7893,N_6190,N_6350);
nand U7894 (N_7894,N_6467,N_6608);
xor U7895 (N_7895,N_6476,N_6574);
nand U7896 (N_7896,N_6378,N_6434);
nand U7897 (N_7897,N_6906,N_6792);
nand U7898 (N_7898,N_6165,N_6337);
nor U7899 (N_7899,N_6832,N_6080);
and U7900 (N_7900,N_6366,N_6813);
nand U7901 (N_7901,N_6499,N_6261);
and U7902 (N_7902,N_6355,N_6213);
xnor U7903 (N_7903,N_6745,N_6917);
nor U7904 (N_7904,N_6843,N_6997);
xnor U7905 (N_7905,N_6663,N_6326);
and U7906 (N_7906,N_6740,N_6469);
nor U7907 (N_7907,N_6504,N_6122);
and U7908 (N_7908,N_6337,N_6875);
xnor U7909 (N_7909,N_6726,N_6685);
and U7910 (N_7910,N_6120,N_6075);
nor U7911 (N_7911,N_6483,N_6171);
xor U7912 (N_7912,N_6545,N_6739);
xor U7913 (N_7913,N_6124,N_6802);
or U7914 (N_7914,N_6996,N_6302);
or U7915 (N_7915,N_6030,N_6435);
nor U7916 (N_7916,N_6123,N_6355);
xnor U7917 (N_7917,N_6904,N_6128);
nand U7918 (N_7918,N_6708,N_6252);
xor U7919 (N_7919,N_6905,N_6007);
and U7920 (N_7920,N_6460,N_6649);
and U7921 (N_7921,N_6761,N_6936);
or U7922 (N_7922,N_6896,N_6643);
nor U7923 (N_7923,N_6261,N_6318);
nand U7924 (N_7924,N_6532,N_6951);
and U7925 (N_7925,N_6003,N_6333);
nand U7926 (N_7926,N_6052,N_6761);
nor U7927 (N_7927,N_6658,N_6724);
nand U7928 (N_7928,N_6366,N_6624);
nor U7929 (N_7929,N_6707,N_6325);
or U7930 (N_7930,N_6762,N_6900);
nor U7931 (N_7931,N_6602,N_6766);
xor U7932 (N_7932,N_6981,N_6736);
and U7933 (N_7933,N_6744,N_6407);
nor U7934 (N_7934,N_6301,N_6626);
xor U7935 (N_7935,N_6309,N_6533);
nor U7936 (N_7936,N_6832,N_6854);
nand U7937 (N_7937,N_6682,N_6142);
nor U7938 (N_7938,N_6453,N_6109);
and U7939 (N_7939,N_6226,N_6949);
nand U7940 (N_7940,N_6189,N_6741);
nand U7941 (N_7941,N_6124,N_6246);
and U7942 (N_7942,N_6233,N_6052);
xor U7943 (N_7943,N_6079,N_6771);
or U7944 (N_7944,N_6662,N_6417);
or U7945 (N_7945,N_6898,N_6924);
or U7946 (N_7946,N_6337,N_6941);
and U7947 (N_7947,N_6840,N_6260);
xor U7948 (N_7948,N_6150,N_6070);
xnor U7949 (N_7949,N_6694,N_6061);
nor U7950 (N_7950,N_6238,N_6076);
xor U7951 (N_7951,N_6750,N_6826);
or U7952 (N_7952,N_6039,N_6818);
nor U7953 (N_7953,N_6191,N_6628);
nor U7954 (N_7954,N_6019,N_6117);
or U7955 (N_7955,N_6266,N_6957);
nand U7956 (N_7956,N_6370,N_6883);
nand U7957 (N_7957,N_6840,N_6951);
and U7958 (N_7958,N_6658,N_6678);
nor U7959 (N_7959,N_6531,N_6785);
or U7960 (N_7960,N_6538,N_6851);
xnor U7961 (N_7961,N_6811,N_6034);
xnor U7962 (N_7962,N_6862,N_6628);
nand U7963 (N_7963,N_6931,N_6444);
and U7964 (N_7964,N_6604,N_6984);
nand U7965 (N_7965,N_6583,N_6569);
nand U7966 (N_7966,N_6167,N_6846);
or U7967 (N_7967,N_6374,N_6256);
and U7968 (N_7968,N_6959,N_6491);
xor U7969 (N_7969,N_6616,N_6124);
and U7970 (N_7970,N_6705,N_6745);
xor U7971 (N_7971,N_6351,N_6534);
or U7972 (N_7972,N_6013,N_6467);
xnor U7973 (N_7973,N_6588,N_6257);
nand U7974 (N_7974,N_6415,N_6999);
nand U7975 (N_7975,N_6274,N_6126);
and U7976 (N_7976,N_6895,N_6647);
and U7977 (N_7977,N_6254,N_6299);
nor U7978 (N_7978,N_6632,N_6550);
or U7979 (N_7979,N_6488,N_6819);
and U7980 (N_7980,N_6468,N_6151);
and U7981 (N_7981,N_6750,N_6486);
nand U7982 (N_7982,N_6204,N_6541);
nor U7983 (N_7983,N_6800,N_6419);
nand U7984 (N_7984,N_6594,N_6629);
nand U7985 (N_7985,N_6552,N_6070);
nor U7986 (N_7986,N_6430,N_6548);
nor U7987 (N_7987,N_6640,N_6810);
or U7988 (N_7988,N_6659,N_6154);
or U7989 (N_7989,N_6502,N_6611);
xnor U7990 (N_7990,N_6515,N_6223);
nand U7991 (N_7991,N_6648,N_6379);
nor U7992 (N_7992,N_6092,N_6051);
or U7993 (N_7993,N_6215,N_6828);
nand U7994 (N_7994,N_6268,N_6261);
or U7995 (N_7995,N_6549,N_6049);
xor U7996 (N_7996,N_6346,N_6866);
and U7997 (N_7997,N_6196,N_6009);
or U7998 (N_7998,N_6654,N_6957);
and U7999 (N_7999,N_6793,N_6275);
and U8000 (N_8000,N_7418,N_7864);
and U8001 (N_8001,N_7785,N_7288);
nand U8002 (N_8002,N_7954,N_7332);
nand U8003 (N_8003,N_7117,N_7669);
nor U8004 (N_8004,N_7446,N_7909);
or U8005 (N_8005,N_7336,N_7454);
nand U8006 (N_8006,N_7592,N_7077);
xnor U8007 (N_8007,N_7791,N_7170);
nor U8008 (N_8008,N_7005,N_7456);
and U8009 (N_8009,N_7687,N_7022);
or U8010 (N_8010,N_7775,N_7946);
and U8011 (N_8011,N_7874,N_7165);
and U8012 (N_8012,N_7373,N_7325);
nand U8013 (N_8013,N_7660,N_7303);
or U8014 (N_8014,N_7232,N_7227);
nand U8015 (N_8015,N_7981,N_7725);
and U8016 (N_8016,N_7943,N_7881);
nand U8017 (N_8017,N_7247,N_7366);
or U8018 (N_8018,N_7330,N_7289);
and U8019 (N_8019,N_7177,N_7891);
nand U8020 (N_8020,N_7050,N_7072);
nand U8021 (N_8021,N_7533,N_7640);
nor U8022 (N_8022,N_7416,N_7799);
xor U8023 (N_8023,N_7271,N_7906);
or U8024 (N_8024,N_7008,N_7442);
and U8025 (N_8025,N_7938,N_7402);
nor U8026 (N_8026,N_7195,N_7369);
xnor U8027 (N_8027,N_7720,N_7421);
and U8028 (N_8028,N_7635,N_7036);
or U8029 (N_8029,N_7190,N_7882);
and U8030 (N_8030,N_7989,N_7145);
and U8031 (N_8031,N_7007,N_7240);
or U8032 (N_8032,N_7595,N_7994);
nor U8033 (N_8033,N_7110,N_7063);
or U8034 (N_8034,N_7392,N_7738);
xnor U8035 (N_8035,N_7991,N_7593);
xor U8036 (N_8036,N_7098,N_7898);
nor U8037 (N_8037,N_7767,N_7108);
nand U8038 (N_8038,N_7228,N_7379);
nand U8039 (N_8039,N_7915,N_7001);
or U8040 (N_8040,N_7897,N_7286);
and U8041 (N_8041,N_7605,N_7269);
nor U8042 (N_8042,N_7718,N_7835);
nand U8043 (N_8043,N_7957,N_7493);
and U8044 (N_8044,N_7355,N_7252);
xnor U8045 (N_8045,N_7947,N_7322);
nor U8046 (N_8046,N_7320,N_7639);
or U8047 (N_8047,N_7284,N_7408);
or U8048 (N_8048,N_7612,N_7559);
or U8049 (N_8049,N_7041,N_7234);
nand U8050 (N_8050,N_7166,N_7914);
and U8051 (N_8051,N_7088,N_7282);
nand U8052 (N_8052,N_7849,N_7268);
xor U8053 (N_8053,N_7733,N_7224);
xor U8054 (N_8054,N_7144,N_7641);
nor U8055 (N_8055,N_7387,N_7751);
nand U8056 (N_8056,N_7798,N_7863);
and U8057 (N_8057,N_7780,N_7731);
and U8058 (N_8058,N_7934,N_7836);
or U8059 (N_8059,N_7074,N_7067);
and U8060 (N_8060,N_7122,N_7510);
xor U8061 (N_8061,N_7306,N_7528);
and U8062 (N_8062,N_7614,N_7766);
nor U8063 (N_8063,N_7423,N_7464);
or U8064 (N_8064,N_7637,N_7786);
or U8065 (N_8065,N_7087,N_7577);
nand U8066 (N_8066,N_7893,N_7099);
xnor U8067 (N_8067,N_7576,N_7011);
nand U8068 (N_8068,N_7484,N_7372);
xor U8069 (N_8069,N_7583,N_7211);
or U8070 (N_8070,N_7513,N_7018);
nand U8071 (N_8071,N_7212,N_7719);
or U8072 (N_8072,N_7382,N_7033);
xnor U8073 (N_8073,N_7796,N_7932);
and U8074 (N_8074,N_7668,N_7239);
or U8075 (N_8075,N_7105,N_7103);
xnor U8076 (N_8076,N_7710,N_7143);
nor U8077 (N_8077,N_7619,N_7205);
or U8078 (N_8078,N_7899,N_7429);
or U8079 (N_8079,N_7557,N_7753);
nor U8080 (N_8080,N_7942,N_7665);
xor U8081 (N_8081,N_7281,N_7830);
nor U8082 (N_8082,N_7956,N_7169);
and U8083 (N_8083,N_7648,N_7119);
xor U8084 (N_8084,N_7770,N_7193);
nor U8085 (N_8085,N_7304,N_7851);
and U8086 (N_8086,N_7186,N_7542);
xor U8087 (N_8087,N_7264,N_7340);
nand U8088 (N_8088,N_7101,N_7655);
nor U8089 (N_8089,N_7895,N_7734);
and U8090 (N_8090,N_7162,N_7521);
and U8091 (N_8091,N_7401,N_7541);
nor U8092 (N_8092,N_7196,N_7515);
nor U8093 (N_8093,N_7594,N_7996);
or U8094 (N_8094,N_7700,N_7532);
nor U8095 (N_8095,N_7266,N_7329);
or U8096 (N_8096,N_7376,N_7805);
xor U8097 (N_8097,N_7978,N_7817);
xor U8098 (N_8098,N_7457,N_7472);
nand U8099 (N_8099,N_7054,N_7121);
nor U8100 (N_8100,N_7537,N_7902);
nand U8101 (N_8101,N_7495,N_7862);
and U8102 (N_8102,N_7474,N_7032);
nand U8103 (N_8103,N_7507,N_7690);
nand U8104 (N_8104,N_7276,N_7903);
xnor U8105 (N_8105,N_7491,N_7176);
nand U8106 (N_8106,N_7255,N_7326);
nand U8107 (N_8107,N_7311,N_7468);
nand U8108 (N_8108,N_7590,N_7958);
nor U8109 (N_8109,N_7717,N_7709);
or U8110 (N_8110,N_7386,N_7707);
nand U8111 (N_8111,N_7527,N_7092);
or U8112 (N_8112,N_7682,N_7407);
xor U8113 (N_8113,N_7616,N_7986);
xnor U8114 (N_8114,N_7666,N_7979);
nor U8115 (N_8115,N_7302,N_7701);
and U8116 (N_8116,N_7927,N_7451);
and U8117 (N_8117,N_7560,N_7470);
and U8118 (N_8118,N_7524,N_7441);
xnor U8119 (N_8119,N_7997,N_7606);
nand U8120 (N_8120,N_7554,N_7191);
and U8121 (N_8121,N_7028,N_7959);
nand U8122 (N_8122,N_7853,N_7760);
and U8123 (N_8123,N_7926,N_7035);
and U8124 (N_8124,N_7543,N_7124);
or U8125 (N_8125,N_7130,N_7890);
nand U8126 (N_8126,N_7974,N_7246);
or U8127 (N_8127,N_7892,N_7625);
and U8128 (N_8128,N_7012,N_7622);
nor U8129 (N_8129,N_7395,N_7174);
xor U8130 (N_8130,N_7214,N_7218);
nor U8131 (N_8131,N_7797,N_7172);
nor U8132 (N_8132,N_7878,N_7125);
xor U8133 (N_8133,N_7132,N_7919);
xnor U8134 (N_8134,N_7222,N_7419);
and U8135 (N_8135,N_7743,N_7262);
and U8136 (N_8136,N_7683,N_7535);
xnor U8137 (N_8137,N_7434,N_7466);
and U8138 (N_8138,N_7458,N_7779);
nand U8139 (N_8139,N_7192,N_7829);
and U8140 (N_8140,N_7589,N_7275);
nor U8141 (N_8141,N_7764,N_7929);
and U8142 (N_8142,N_7358,N_7868);
or U8143 (N_8143,N_7643,N_7173);
nand U8144 (N_8144,N_7860,N_7925);
nor U8145 (N_8145,N_7531,N_7833);
xor U8146 (N_8146,N_7857,N_7681);
nor U8147 (N_8147,N_7597,N_7551);
xnor U8148 (N_8148,N_7217,N_7064);
nand U8149 (N_8149,N_7354,N_7931);
nand U8150 (N_8150,N_7935,N_7016);
and U8151 (N_8151,N_7280,N_7691);
and U8152 (N_8152,N_7397,N_7178);
xor U8153 (N_8153,N_7657,N_7100);
nand U8154 (N_8154,N_7522,N_7970);
or U8155 (N_8155,N_7658,N_7741);
nor U8156 (N_8156,N_7673,N_7735);
nor U8157 (N_8157,N_7448,N_7185);
or U8158 (N_8158,N_7726,N_7417);
nand U8159 (N_8159,N_7309,N_7327);
and U8160 (N_8160,N_7481,N_7852);
or U8161 (N_8161,N_7604,N_7566);
or U8162 (N_8162,N_7346,N_7952);
and U8163 (N_8163,N_7187,N_7115);
nand U8164 (N_8164,N_7500,N_7360);
and U8165 (N_8165,N_7085,N_7827);
xor U8166 (N_8166,N_7238,N_7343);
nor U8167 (N_8167,N_7285,N_7485);
nor U8168 (N_8168,N_7126,N_7905);
nor U8169 (N_8169,N_7519,N_7053);
or U8170 (N_8170,N_7722,N_7887);
and U8171 (N_8171,N_7420,N_7769);
nor U8172 (N_8172,N_7824,N_7563);
nor U8173 (N_8173,N_7603,N_7414);
xnor U8174 (N_8174,N_7645,N_7503);
nor U8175 (N_8175,N_7825,N_7759);
nor U8176 (N_8176,N_7861,N_7477);
and U8177 (N_8177,N_7618,N_7400);
xor U8178 (N_8178,N_7807,N_7591);
nand U8179 (N_8179,N_7138,N_7661);
or U8180 (N_8180,N_7509,N_7904);
nor U8181 (N_8181,N_7628,N_7998);
xnor U8182 (N_8182,N_7296,N_7870);
and U8183 (N_8183,N_7633,N_7936);
or U8184 (N_8184,N_7708,N_7570);
nand U8185 (N_8185,N_7514,N_7057);
xnor U8186 (N_8186,N_7381,N_7061);
nor U8187 (N_8187,N_7730,N_7802);
or U8188 (N_8188,N_7871,N_7702);
nand U8189 (N_8189,N_7911,N_7984);
nand U8190 (N_8190,N_7889,N_7896);
nand U8191 (N_8191,N_7368,N_7461);
nand U8192 (N_8192,N_7962,N_7746);
nor U8193 (N_8193,N_7312,N_7384);
xnor U8194 (N_8194,N_7651,N_7243);
xnor U8195 (N_8195,N_7610,N_7111);
or U8196 (N_8196,N_7762,N_7287);
nand U8197 (N_8197,N_7685,N_7081);
nor U8198 (N_8198,N_7784,N_7608);
and U8199 (N_8199,N_7804,N_7877);
nor U8200 (N_8200,N_7985,N_7250);
nor U8201 (N_8201,N_7757,N_7344);
nand U8202 (N_8202,N_7809,N_7965);
or U8203 (N_8203,N_7015,N_7654);
nand U8204 (N_8204,N_7009,N_7147);
xor U8205 (N_8205,N_7930,N_7244);
or U8206 (N_8206,N_7950,N_7237);
and U8207 (N_8207,N_7948,N_7412);
nor U8208 (N_8208,N_7353,N_7790);
and U8209 (N_8209,N_7728,N_7422);
xnor U8210 (N_8210,N_7025,N_7494);
xnor U8211 (N_8211,N_7501,N_7116);
and U8212 (N_8212,N_7127,N_7547);
nand U8213 (N_8213,N_7209,N_7571);
or U8214 (N_8214,N_7140,N_7567);
and U8215 (N_8215,N_7561,N_7980);
nand U8216 (N_8216,N_7960,N_7439);
or U8217 (N_8217,N_7480,N_7342);
and U8218 (N_8218,N_7265,N_7424);
or U8219 (N_8219,N_7436,N_7624);
nor U8220 (N_8220,N_7800,N_7273);
xor U8221 (N_8221,N_7686,N_7107);
xnor U8222 (N_8222,N_7114,N_7601);
and U8223 (N_8223,N_7109,N_7854);
or U8224 (N_8224,N_7945,N_7939);
nand U8225 (N_8225,N_7955,N_7774);
xor U8226 (N_8226,N_7729,N_7940);
or U8227 (N_8227,N_7155,N_7534);
xnor U8228 (N_8228,N_7553,N_7236);
nand U8229 (N_8229,N_7787,N_7199);
nand U8230 (N_8230,N_7748,N_7713);
xnor U8231 (N_8231,N_7506,N_7341);
nor U8232 (N_8232,N_7781,N_7813);
and U8233 (N_8233,N_7671,N_7812);
nor U8234 (N_8234,N_7314,N_7843);
nand U8235 (N_8235,N_7003,N_7575);
nand U8236 (N_8236,N_7093,N_7082);
nand U8237 (N_8237,N_7294,N_7982);
and U8238 (N_8238,N_7215,N_7638);
nor U8239 (N_8239,N_7617,N_7164);
xor U8240 (N_8240,N_7321,N_7095);
and U8241 (N_8241,N_7693,N_7399);
nand U8242 (N_8242,N_7462,N_7811);
or U8243 (N_8243,N_7789,N_7388);
or U8244 (N_8244,N_7675,N_7453);
and U8245 (N_8245,N_7473,N_7497);
nand U8246 (N_8246,N_7987,N_7014);
nor U8247 (N_8247,N_7377,N_7310);
or U8248 (N_8248,N_7581,N_7488);
nand U8249 (N_8249,N_7317,N_7113);
or U8250 (N_8250,N_7968,N_7133);
and U8251 (N_8251,N_7803,N_7578);
nand U8252 (N_8252,N_7391,N_7689);
and U8253 (N_8253,N_7696,N_7075);
and U8254 (N_8254,N_7405,N_7256);
nand U8255 (N_8255,N_7692,N_7818);
nand U8256 (N_8256,N_7027,N_7374);
nor U8257 (N_8257,N_7511,N_7846);
and U8258 (N_8258,N_7712,N_7971);
or U8259 (N_8259,N_7293,N_7150);
xor U8260 (N_8260,N_7837,N_7716);
and U8261 (N_8261,N_7705,N_7822);
nor U8262 (N_8262,N_7019,N_7703);
and U8263 (N_8263,N_7060,N_7794);
nor U8264 (N_8264,N_7875,N_7134);
xor U8265 (N_8265,N_7034,N_7990);
or U8266 (N_8266,N_7208,N_7175);
or U8267 (N_8267,N_7736,N_7248);
xor U8268 (N_8268,N_7739,N_7002);
xor U8269 (N_8269,N_7086,N_7051);
and U8270 (N_8270,N_7924,N_7385);
xnor U8271 (N_8271,N_7676,N_7880);
nor U8272 (N_8272,N_7684,N_7944);
nand U8273 (N_8273,N_7426,N_7972);
nor U8274 (N_8274,N_7646,N_7492);
nand U8275 (N_8275,N_7042,N_7367);
nand U8276 (N_8276,N_7204,N_7069);
xor U8277 (N_8277,N_7873,N_7425);
xor U8278 (N_8278,N_7520,N_7318);
nand U8279 (N_8279,N_7845,N_7525);
nand U8280 (N_8280,N_7146,N_7564);
nor U8281 (N_8281,N_7151,N_7023);
nand U8282 (N_8282,N_7806,N_7573);
or U8283 (N_8283,N_7352,N_7153);
or U8284 (N_8284,N_7450,N_7530);
nand U8285 (N_8285,N_7844,N_7058);
nand U8286 (N_8286,N_7776,N_7912);
xnor U8287 (N_8287,N_7197,N_7249);
and U8288 (N_8288,N_7884,N_7749);
nor U8289 (N_8289,N_7517,N_7337);
xnor U8290 (N_8290,N_7277,N_7308);
nand U8291 (N_8291,N_7200,N_7755);
or U8292 (N_8292,N_7476,N_7097);
xor U8293 (N_8293,N_7783,N_7923);
and U8294 (N_8294,N_7688,N_7771);
or U8295 (N_8295,N_7141,N_7350);
xnor U8296 (N_8296,N_7406,N_7832);
nor U8297 (N_8297,N_7482,N_7123);
nand U8298 (N_8298,N_7463,N_7580);
and U8299 (N_8299,N_7139,N_7663);
and U8300 (N_8300,N_7788,N_7096);
or U8301 (N_8301,N_7937,N_7052);
nor U8302 (N_8302,N_7071,N_7410);
and U8303 (N_8303,N_7516,N_7131);
xnor U8304 (N_8304,N_7740,N_7920);
or U8305 (N_8305,N_7378,N_7679);
or U8306 (N_8306,N_7210,N_7198);
or U8307 (N_8307,N_7297,N_7842);
or U8308 (N_8308,N_7398,N_7886);
and U8309 (N_8309,N_7536,N_7647);
or U8310 (N_8310,N_7548,N_7765);
and U8311 (N_8311,N_7274,N_7834);
nand U8312 (N_8312,N_7292,N_7489);
xnor U8313 (N_8313,N_7435,N_7756);
xor U8314 (N_8314,N_7992,N_7031);
nand U8315 (N_8315,N_7043,N_7662);
xor U8316 (N_8316,N_7855,N_7574);
or U8317 (N_8317,N_7216,N_7184);
nand U8318 (N_8318,N_7483,N_7221);
or U8319 (N_8319,N_7004,N_7182);
nor U8320 (N_8320,N_7869,N_7094);
and U8321 (N_8321,N_7859,N_7773);
or U8322 (N_8322,N_7431,N_7933);
xnor U8323 (N_8323,N_7727,N_7433);
or U8324 (N_8324,N_7445,N_7163);
nand U8325 (N_8325,N_7872,N_7251);
or U8326 (N_8326,N_7307,N_7747);
xor U8327 (N_8327,N_7430,N_7371);
or U8328 (N_8328,N_7118,N_7291);
or U8329 (N_8329,N_7112,N_7969);
xor U8330 (N_8330,N_7049,N_7226);
or U8331 (N_8331,N_7758,N_7951);
and U8332 (N_8332,N_7900,N_7549);
nand U8333 (N_8333,N_7518,N_7055);
or U8334 (N_8334,N_7778,N_7737);
nand U8335 (N_8335,N_7831,N_7370);
xnor U8336 (N_8336,N_7465,N_7588);
nand U8337 (N_8337,N_7242,N_7039);
or U8338 (N_8338,N_7207,N_7203);
or U8339 (N_8339,N_7335,N_7620);
nand U8340 (N_8340,N_7672,N_7404);
xnor U8341 (N_8341,N_7623,N_7079);
and U8342 (N_8342,N_7602,N_7586);
xnor U8343 (N_8343,N_7680,N_7467);
nor U8344 (N_8344,N_7415,N_7409);
xnor U8345 (N_8345,N_7848,N_7556);
and U8346 (N_8346,N_7089,N_7154);
nor U8347 (N_8347,N_7455,N_7711);
or U8348 (N_8348,N_7922,N_7910);
xor U8349 (N_8349,N_7697,N_7393);
and U8350 (N_8350,N_7677,N_7026);
or U8351 (N_8351,N_7656,N_7894);
and U8352 (N_8352,N_7148,N_7777);
xor U8353 (N_8353,N_7364,N_7331);
nor U8354 (N_8354,N_7883,N_7440);
nand U8355 (N_8355,N_7315,N_7512);
xnor U8356 (N_8356,N_7631,N_7587);
nand U8357 (N_8357,N_7821,N_7562);
nor U8358 (N_8358,N_7136,N_7629);
xnor U8359 (N_8359,N_7065,N_7636);
nor U8360 (N_8360,N_7539,N_7428);
and U8361 (N_8361,N_7615,N_7363);
nor U8362 (N_8362,N_7913,N_7847);
or U8363 (N_8363,N_7348,N_7828);
or U8364 (N_8364,N_7091,N_7714);
xor U8365 (N_8365,N_7283,N_7156);
nor U8366 (N_8366,N_7263,N_7850);
nand U8367 (N_8367,N_7867,N_7159);
nor U8368 (N_8368,N_7901,N_7632);
xor U8369 (N_8369,N_7475,N_7598);
nand U8370 (N_8370,N_7490,N_7976);
xor U8371 (N_8371,N_7356,N_7820);
nand U8372 (N_8372,N_7916,N_7678);
nor U8373 (N_8373,N_7865,N_7024);
nor U8374 (N_8374,N_7167,N_7070);
nor U8375 (N_8375,N_7323,N_7438);
xor U8376 (N_8376,N_7021,N_7840);
and U8377 (N_8377,N_7772,N_7839);
and U8378 (N_8378,N_7823,N_7826);
and U8379 (N_8379,N_7538,N_7102);
xnor U8380 (N_8380,N_7995,N_7219);
or U8381 (N_8381,N_7763,N_7667);
nor U8382 (N_8382,N_7254,N_7761);
nor U8383 (N_8383,N_7241,N_7963);
nand U8384 (N_8384,N_7301,N_7390);
nor U8385 (N_8385,N_7918,N_7964);
or U8386 (N_8386,N_7568,N_7270);
and U8387 (N_8387,N_7334,N_7258);
nand U8388 (N_8388,N_7611,N_7449);
nor U8389 (N_8389,N_7201,N_7202);
nand U8390 (N_8390,N_7841,N_7161);
and U8391 (N_8391,N_7706,N_7644);
and U8392 (N_8392,N_7260,N_7626);
nand U8393 (N_8393,N_7659,N_7104);
nand U8394 (N_8394,N_7444,N_7649);
or U8395 (N_8395,N_7585,N_7526);
and U8396 (N_8396,N_7447,N_7375);
and U8397 (N_8397,N_7966,N_7298);
nor U8398 (N_8398,N_7316,N_7715);
xnor U8399 (N_8399,N_7907,N_7856);
nor U8400 (N_8400,N_7609,N_7724);
and U8401 (N_8401,N_7469,N_7106);
or U8402 (N_8402,N_7782,N_7674);
and U8403 (N_8403,N_7471,N_7080);
and U8404 (N_8404,N_7128,N_7698);
xnor U8405 (N_8405,N_7630,N_7188);
nor U8406 (N_8406,N_7967,N_7020);
and U8407 (N_8407,N_7068,N_7090);
and U8408 (N_8408,N_7993,N_7858);
or U8409 (N_8409,N_7040,N_7479);
nand U8410 (N_8410,N_7555,N_7988);
or U8411 (N_8411,N_7816,N_7300);
and U8412 (N_8412,N_7029,N_7579);
nand U8413 (N_8413,N_7814,N_7885);
nand U8414 (N_8414,N_7059,N_7272);
nand U8415 (N_8415,N_7544,N_7582);
nand U8416 (N_8416,N_7838,N_7752);
nor U8417 (N_8417,N_7505,N_7349);
xor U8418 (N_8418,N_7152,N_7030);
xnor U8419 (N_8419,N_7487,N_7613);
nor U8420 (N_8420,N_7142,N_7013);
or U8421 (N_8421,N_7324,N_7653);
xor U8422 (N_8422,N_7704,N_7380);
and U8423 (N_8423,N_7084,N_7206);
nand U8424 (N_8424,N_7596,N_7313);
and U8425 (N_8425,N_7795,N_7973);
nand U8426 (N_8426,N_7650,N_7499);
nor U8427 (N_8427,N_7158,N_7921);
nor U8428 (N_8428,N_7745,N_7999);
nand U8429 (N_8429,N_7403,N_7267);
nand U8430 (N_8430,N_7584,N_7550);
and U8431 (N_8431,N_7365,N_7183);
nand U8432 (N_8432,N_7345,N_7694);
nand U8433 (N_8433,N_7552,N_7502);
or U8434 (N_8434,N_7225,N_7290);
nor U8435 (N_8435,N_7744,N_7160);
or U8436 (N_8436,N_7815,N_7545);
nand U8437 (N_8437,N_7621,N_7793);
nor U8438 (N_8438,N_7137,N_7220);
and U8439 (N_8439,N_7351,N_7496);
or U8440 (N_8440,N_7498,N_7006);
nor U8441 (N_8441,N_7044,N_7171);
nand U8442 (N_8442,N_7460,N_7888);
and U8443 (N_8443,N_7572,N_7664);
nand U8444 (N_8444,N_7486,N_7565);
and U8445 (N_8445,N_7078,N_7347);
or U8446 (N_8446,N_7866,N_7235);
and U8447 (N_8447,N_7048,N_7478);
and U8448 (N_8448,N_7168,N_7181);
nand U8449 (N_8449,N_7213,N_7357);
nor U8450 (N_8450,N_7459,N_7383);
and U8451 (N_8451,N_7389,N_7257);
xor U8452 (N_8452,N_7437,N_7699);
nand U8453 (N_8453,N_7073,N_7083);
or U8454 (N_8454,N_7917,N_7810);
nor U8455 (N_8455,N_7359,N_7362);
nand U8456 (N_8456,N_7299,N_7189);
xnor U8457 (N_8457,N_7231,N_7339);
or U8458 (N_8458,N_7278,N_7627);
or U8459 (N_8459,N_7792,N_7754);
xor U8460 (N_8460,N_7047,N_7319);
and U8461 (N_8461,N_7750,N_7961);
nor U8462 (N_8462,N_7695,N_7508);
or U8463 (N_8463,N_7056,N_7642);
nand U8464 (N_8464,N_7983,N_7540);
or U8465 (N_8465,N_7037,N_7452);
nand U8466 (N_8466,N_7928,N_7261);
nand U8467 (N_8467,N_7443,N_7194);
and U8468 (N_8468,N_7179,N_7180);
xor U8469 (N_8469,N_7908,N_7305);
xor U8470 (N_8470,N_7279,N_7338);
xnor U8471 (N_8471,N_7396,N_7977);
xor U8472 (N_8472,N_7017,N_7076);
xor U8473 (N_8473,N_7066,N_7361);
nor U8474 (N_8474,N_7010,N_7245);
nor U8475 (N_8475,N_7230,N_7259);
and U8476 (N_8476,N_7149,N_7295);
and U8477 (N_8477,N_7652,N_7432);
and U8478 (N_8478,N_7558,N_7879);
or U8479 (N_8479,N_7607,N_7670);
xnor U8480 (N_8480,N_7504,N_7120);
and U8481 (N_8481,N_7046,N_7721);
nand U8482 (N_8482,N_7546,N_7569);
and U8483 (N_8483,N_7876,N_7038);
and U8484 (N_8484,N_7333,N_7135);
xor U8485 (N_8485,N_7223,N_7732);
or U8486 (N_8486,N_7600,N_7941);
nand U8487 (N_8487,N_7819,N_7634);
xnor U8488 (N_8488,N_7413,N_7975);
or U8489 (N_8489,N_7808,N_7427);
nand U8490 (N_8490,N_7157,N_7000);
xnor U8491 (N_8491,N_7394,N_7599);
and U8492 (N_8492,N_7411,N_7045);
nand U8493 (N_8493,N_7529,N_7949);
nand U8494 (N_8494,N_7129,N_7953);
and U8495 (N_8495,N_7768,N_7233);
xnor U8496 (N_8496,N_7253,N_7229);
and U8497 (N_8497,N_7523,N_7742);
and U8498 (N_8498,N_7062,N_7801);
nand U8499 (N_8499,N_7328,N_7723);
and U8500 (N_8500,N_7981,N_7023);
and U8501 (N_8501,N_7537,N_7936);
nand U8502 (N_8502,N_7897,N_7723);
nand U8503 (N_8503,N_7380,N_7502);
and U8504 (N_8504,N_7708,N_7028);
xnor U8505 (N_8505,N_7357,N_7365);
or U8506 (N_8506,N_7373,N_7446);
nand U8507 (N_8507,N_7975,N_7813);
nand U8508 (N_8508,N_7981,N_7176);
nor U8509 (N_8509,N_7522,N_7459);
or U8510 (N_8510,N_7980,N_7487);
nor U8511 (N_8511,N_7890,N_7056);
nor U8512 (N_8512,N_7771,N_7199);
or U8513 (N_8513,N_7715,N_7559);
or U8514 (N_8514,N_7777,N_7448);
xor U8515 (N_8515,N_7167,N_7388);
and U8516 (N_8516,N_7594,N_7168);
nor U8517 (N_8517,N_7121,N_7461);
or U8518 (N_8518,N_7399,N_7265);
nand U8519 (N_8519,N_7885,N_7144);
or U8520 (N_8520,N_7739,N_7182);
nand U8521 (N_8521,N_7037,N_7411);
xor U8522 (N_8522,N_7674,N_7590);
nor U8523 (N_8523,N_7918,N_7250);
nor U8524 (N_8524,N_7989,N_7350);
nor U8525 (N_8525,N_7774,N_7213);
nor U8526 (N_8526,N_7947,N_7578);
or U8527 (N_8527,N_7400,N_7270);
nand U8528 (N_8528,N_7741,N_7501);
or U8529 (N_8529,N_7850,N_7857);
nor U8530 (N_8530,N_7776,N_7589);
nand U8531 (N_8531,N_7934,N_7344);
nor U8532 (N_8532,N_7870,N_7036);
nor U8533 (N_8533,N_7586,N_7753);
xor U8534 (N_8534,N_7965,N_7334);
nor U8535 (N_8535,N_7917,N_7963);
or U8536 (N_8536,N_7997,N_7855);
and U8537 (N_8537,N_7600,N_7400);
xor U8538 (N_8538,N_7303,N_7733);
nor U8539 (N_8539,N_7894,N_7657);
xor U8540 (N_8540,N_7888,N_7859);
nor U8541 (N_8541,N_7506,N_7880);
and U8542 (N_8542,N_7028,N_7698);
xnor U8543 (N_8543,N_7424,N_7319);
nand U8544 (N_8544,N_7158,N_7972);
nand U8545 (N_8545,N_7326,N_7228);
or U8546 (N_8546,N_7601,N_7165);
nand U8547 (N_8547,N_7508,N_7709);
or U8548 (N_8548,N_7158,N_7876);
nor U8549 (N_8549,N_7307,N_7737);
nand U8550 (N_8550,N_7996,N_7151);
and U8551 (N_8551,N_7081,N_7799);
or U8552 (N_8552,N_7122,N_7273);
nor U8553 (N_8553,N_7185,N_7332);
nor U8554 (N_8554,N_7134,N_7967);
nor U8555 (N_8555,N_7907,N_7289);
xor U8556 (N_8556,N_7741,N_7054);
nand U8557 (N_8557,N_7008,N_7418);
nor U8558 (N_8558,N_7518,N_7176);
xor U8559 (N_8559,N_7375,N_7627);
nand U8560 (N_8560,N_7767,N_7928);
nand U8561 (N_8561,N_7829,N_7933);
nand U8562 (N_8562,N_7691,N_7871);
or U8563 (N_8563,N_7996,N_7901);
xor U8564 (N_8564,N_7792,N_7280);
or U8565 (N_8565,N_7689,N_7599);
nand U8566 (N_8566,N_7512,N_7596);
and U8567 (N_8567,N_7482,N_7274);
or U8568 (N_8568,N_7438,N_7498);
and U8569 (N_8569,N_7905,N_7708);
nor U8570 (N_8570,N_7024,N_7734);
nand U8571 (N_8571,N_7298,N_7137);
or U8572 (N_8572,N_7118,N_7135);
and U8573 (N_8573,N_7059,N_7885);
or U8574 (N_8574,N_7381,N_7457);
or U8575 (N_8575,N_7938,N_7377);
or U8576 (N_8576,N_7974,N_7706);
and U8577 (N_8577,N_7440,N_7496);
and U8578 (N_8578,N_7311,N_7285);
xor U8579 (N_8579,N_7127,N_7674);
xnor U8580 (N_8580,N_7712,N_7166);
and U8581 (N_8581,N_7374,N_7774);
and U8582 (N_8582,N_7661,N_7769);
or U8583 (N_8583,N_7245,N_7728);
nor U8584 (N_8584,N_7917,N_7451);
xor U8585 (N_8585,N_7745,N_7201);
nand U8586 (N_8586,N_7234,N_7437);
and U8587 (N_8587,N_7453,N_7227);
nand U8588 (N_8588,N_7519,N_7993);
nand U8589 (N_8589,N_7866,N_7371);
nor U8590 (N_8590,N_7593,N_7647);
nor U8591 (N_8591,N_7843,N_7382);
xnor U8592 (N_8592,N_7227,N_7440);
xnor U8593 (N_8593,N_7014,N_7434);
nand U8594 (N_8594,N_7988,N_7643);
xor U8595 (N_8595,N_7742,N_7784);
nand U8596 (N_8596,N_7636,N_7218);
nor U8597 (N_8597,N_7423,N_7330);
nor U8598 (N_8598,N_7365,N_7060);
nor U8599 (N_8599,N_7052,N_7455);
nor U8600 (N_8600,N_7512,N_7772);
nor U8601 (N_8601,N_7397,N_7008);
and U8602 (N_8602,N_7735,N_7543);
and U8603 (N_8603,N_7446,N_7346);
xor U8604 (N_8604,N_7967,N_7807);
and U8605 (N_8605,N_7635,N_7716);
nand U8606 (N_8606,N_7272,N_7052);
and U8607 (N_8607,N_7564,N_7542);
or U8608 (N_8608,N_7048,N_7953);
nor U8609 (N_8609,N_7026,N_7448);
and U8610 (N_8610,N_7615,N_7480);
xor U8611 (N_8611,N_7396,N_7016);
xnor U8612 (N_8612,N_7061,N_7089);
and U8613 (N_8613,N_7899,N_7021);
nor U8614 (N_8614,N_7197,N_7944);
and U8615 (N_8615,N_7178,N_7807);
xor U8616 (N_8616,N_7783,N_7946);
xnor U8617 (N_8617,N_7038,N_7414);
nand U8618 (N_8618,N_7839,N_7362);
and U8619 (N_8619,N_7955,N_7503);
or U8620 (N_8620,N_7390,N_7582);
nand U8621 (N_8621,N_7639,N_7080);
and U8622 (N_8622,N_7701,N_7182);
nor U8623 (N_8623,N_7169,N_7249);
nand U8624 (N_8624,N_7461,N_7610);
xor U8625 (N_8625,N_7175,N_7786);
or U8626 (N_8626,N_7562,N_7632);
xnor U8627 (N_8627,N_7565,N_7399);
xor U8628 (N_8628,N_7523,N_7966);
and U8629 (N_8629,N_7678,N_7213);
nor U8630 (N_8630,N_7199,N_7406);
or U8631 (N_8631,N_7835,N_7244);
nor U8632 (N_8632,N_7008,N_7984);
and U8633 (N_8633,N_7732,N_7375);
and U8634 (N_8634,N_7640,N_7532);
xnor U8635 (N_8635,N_7555,N_7885);
nand U8636 (N_8636,N_7584,N_7716);
nor U8637 (N_8637,N_7067,N_7666);
nor U8638 (N_8638,N_7113,N_7149);
and U8639 (N_8639,N_7551,N_7977);
nor U8640 (N_8640,N_7763,N_7439);
nor U8641 (N_8641,N_7571,N_7355);
and U8642 (N_8642,N_7623,N_7642);
nand U8643 (N_8643,N_7807,N_7673);
nor U8644 (N_8644,N_7299,N_7097);
nand U8645 (N_8645,N_7108,N_7584);
or U8646 (N_8646,N_7750,N_7588);
nor U8647 (N_8647,N_7069,N_7064);
nand U8648 (N_8648,N_7696,N_7978);
or U8649 (N_8649,N_7363,N_7501);
nor U8650 (N_8650,N_7298,N_7450);
or U8651 (N_8651,N_7461,N_7012);
xor U8652 (N_8652,N_7804,N_7910);
nor U8653 (N_8653,N_7735,N_7250);
or U8654 (N_8654,N_7805,N_7560);
nor U8655 (N_8655,N_7453,N_7637);
or U8656 (N_8656,N_7463,N_7905);
nand U8657 (N_8657,N_7862,N_7907);
nor U8658 (N_8658,N_7608,N_7814);
nor U8659 (N_8659,N_7744,N_7472);
xnor U8660 (N_8660,N_7520,N_7147);
or U8661 (N_8661,N_7287,N_7067);
and U8662 (N_8662,N_7282,N_7671);
nand U8663 (N_8663,N_7328,N_7392);
or U8664 (N_8664,N_7983,N_7104);
or U8665 (N_8665,N_7594,N_7711);
xor U8666 (N_8666,N_7938,N_7556);
xnor U8667 (N_8667,N_7535,N_7559);
and U8668 (N_8668,N_7753,N_7184);
nor U8669 (N_8669,N_7690,N_7429);
xnor U8670 (N_8670,N_7214,N_7624);
nand U8671 (N_8671,N_7116,N_7144);
nor U8672 (N_8672,N_7847,N_7620);
xor U8673 (N_8673,N_7440,N_7354);
and U8674 (N_8674,N_7629,N_7090);
nor U8675 (N_8675,N_7481,N_7300);
xnor U8676 (N_8676,N_7900,N_7733);
or U8677 (N_8677,N_7732,N_7284);
nor U8678 (N_8678,N_7299,N_7754);
and U8679 (N_8679,N_7382,N_7809);
nand U8680 (N_8680,N_7375,N_7001);
xnor U8681 (N_8681,N_7701,N_7896);
nor U8682 (N_8682,N_7084,N_7684);
nor U8683 (N_8683,N_7570,N_7349);
xor U8684 (N_8684,N_7057,N_7024);
nand U8685 (N_8685,N_7888,N_7719);
nor U8686 (N_8686,N_7888,N_7122);
xor U8687 (N_8687,N_7336,N_7471);
nor U8688 (N_8688,N_7844,N_7424);
or U8689 (N_8689,N_7847,N_7445);
and U8690 (N_8690,N_7543,N_7534);
nand U8691 (N_8691,N_7656,N_7741);
nand U8692 (N_8692,N_7995,N_7445);
or U8693 (N_8693,N_7347,N_7579);
nor U8694 (N_8694,N_7794,N_7848);
nor U8695 (N_8695,N_7981,N_7314);
and U8696 (N_8696,N_7394,N_7504);
nand U8697 (N_8697,N_7618,N_7860);
and U8698 (N_8698,N_7477,N_7900);
and U8699 (N_8699,N_7423,N_7421);
nor U8700 (N_8700,N_7248,N_7998);
or U8701 (N_8701,N_7615,N_7118);
or U8702 (N_8702,N_7557,N_7203);
nor U8703 (N_8703,N_7652,N_7267);
xnor U8704 (N_8704,N_7255,N_7512);
nor U8705 (N_8705,N_7408,N_7271);
nor U8706 (N_8706,N_7499,N_7293);
nor U8707 (N_8707,N_7254,N_7248);
nand U8708 (N_8708,N_7349,N_7171);
xor U8709 (N_8709,N_7725,N_7636);
nand U8710 (N_8710,N_7785,N_7272);
nor U8711 (N_8711,N_7029,N_7912);
and U8712 (N_8712,N_7260,N_7658);
nand U8713 (N_8713,N_7054,N_7651);
xnor U8714 (N_8714,N_7582,N_7230);
xnor U8715 (N_8715,N_7664,N_7364);
and U8716 (N_8716,N_7710,N_7471);
and U8717 (N_8717,N_7290,N_7125);
xnor U8718 (N_8718,N_7167,N_7833);
nor U8719 (N_8719,N_7797,N_7023);
or U8720 (N_8720,N_7823,N_7205);
nand U8721 (N_8721,N_7586,N_7012);
xor U8722 (N_8722,N_7488,N_7692);
nor U8723 (N_8723,N_7278,N_7656);
xnor U8724 (N_8724,N_7696,N_7558);
xnor U8725 (N_8725,N_7271,N_7342);
and U8726 (N_8726,N_7245,N_7678);
and U8727 (N_8727,N_7817,N_7947);
xor U8728 (N_8728,N_7083,N_7990);
and U8729 (N_8729,N_7786,N_7418);
or U8730 (N_8730,N_7752,N_7696);
nor U8731 (N_8731,N_7932,N_7526);
nor U8732 (N_8732,N_7256,N_7444);
nor U8733 (N_8733,N_7888,N_7032);
and U8734 (N_8734,N_7372,N_7293);
nor U8735 (N_8735,N_7513,N_7111);
nand U8736 (N_8736,N_7787,N_7562);
nor U8737 (N_8737,N_7201,N_7216);
nand U8738 (N_8738,N_7335,N_7911);
nand U8739 (N_8739,N_7718,N_7673);
xnor U8740 (N_8740,N_7956,N_7358);
nor U8741 (N_8741,N_7970,N_7323);
or U8742 (N_8742,N_7837,N_7953);
or U8743 (N_8743,N_7156,N_7727);
nand U8744 (N_8744,N_7582,N_7401);
xnor U8745 (N_8745,N_7068,N_7737);
or U8746 (N_8746,N_7056,N_7274);
nand U8747 (N_8747,N_7742,N_7681);
xnor U8748 (N_8748,N_7701,N_7352);
nor U8749 (N_8749,N_7952,N_7561);
or U8750 (N_8750,N_7339,N_7199);
nor U8751 (N_8751,N_7857,N_7662);
xnor U8752 (N_8752,N_7496,N_7534);
nor U8753 (N_8753,N_7069,N_7086);
or U8754 (N_8754,N_7909,N_7019);
nor U8755 (N_8755,N_7692,N_7626);
nor U8756 (N_8756,N_7704,N_7146);
xor U8757 (N_8757,N_7027,N_7729);
xnor U8758 (N_8758,N_7189,N_7993);
nand U8759 (N_8759,N_7755,N_7654);
nand U8760 (N_8760,N_7935,N_7467);
nor U8761 (N_8761,N_7303,N_7795);
and U8762 (N_8762,N_7950,N_7110);
or U8763 (N_8763,N_7518,N_7103);
and U8764 (N_8764,N_7161,N_7369);
xnor U8765 (N_8765,N_7726,N_7587);
or U8766 (N_8766,N_7927,N_7261);
nand U8767 (N_8767,N_7744,N_7996);
nor U8768 (N_8768,N_7607,N_7294);
nand U8769 (N_8769,N_7705,N_7255);
or U8770 (N_8770,N_7348,N_7032);
and U8771 (N_8771,N_7474,N_7195);
and U8772 (N_8772,N_7693,N_7256);
nor U8773 (N_8773,N_7468,N_7116);
nand U8774 (N_8774,N_7813,N_7690);
xor U8775 (N_8775,N_7930,N_7966);
nor U8776 (N_8776,N_7992,N_7020);
or U8777 (N_8777,N_7350,N_7091);
or U8778 (N_8778,N_7840,N_7960);
nor U8779 (N_8779,N_7800,N_7675);
or U8780 (N_8780,N_7407,N_7502);
nand U8781 (N_8781,N_7805,N_7706);
nand U8782 (N_8782,N_7516,N_7425);
xor U8783 (N_8783,N_7996,N_7560);
xnor U8784 (N_8784,N_7742,N_7267);
and U8785 (N_8785,N_7783,N_7155);
nor U8786 (N_8786,N_7920,N_7250);
xor U8787 (N_8787,N_7073,N_7360);
and U8788 (N_8788,N_7552,N_7532);
nand U8789 (N_8789,N_7979,N_7440);
or U8790 (N_8790,N_7841,N_7409);
nand U8791 (N_8791,N_7229,N_7247);
nor U8792 (N_8792,N_7742,N_7228);
nor U8793 (N_8793,N_7457,N_7569);
and U8794 (N_8794,N_7178,N_7951);
xor U8795 (N_8795,N_7128,N_7626);
and U8796 (N_8796,N_7020,N_7166);
nor U8797 (N_8797,N_7031,N_7266);
or U8798 (N_8798,N_7059,N_7870);
nor U8799 (N_8799,N_7699,N_7360);
xor U8800 (N_8800,N_7175,N_7617);
nor U8801 (N_8801,N_7819,N_7684);
and U8802 (N_8802,N_7344,N_7286);
or U8803 (N_8803,N_7438,N_7131);
nor U8804 (N_8804,N_7507,N_7210);
nor U8805 (N_8805,N_7682,N_7193);
xor U8806 (N_8806,N_7143,N_7313);
and U8807 (N_8807,N_7675,N_7876);
and U8808 (N_8808,N_7152,N_7315);
or U8809 (N_8809,N_7530,N_7391);
or U8810 (N_8810,N_7008,N_7920);
nand U8811 (N_8811,N_7824,N_7097);
nand U8812 (N_8812,N_7101,N_7183);
xnor U8813 (N_8813,N_7368,N_7106);
nand U8814 (N_8814,N_7772,N_7114);
nor U8815 (N_8815,N_7106,N_7547);
xnor U8816 (N_8816,N_7706,N_7025);
xor U8817 (N_8817,N_7174,N_7758);
xor U8818 (N_8818,N_7692,N_7717);
nor U8819 (N_8819,N_7491,N_7057);
and U8820 (N_8820,N_7580,N_7189);
nor U8821 (N_8821,N_7253,N_7693);
and U8822 (N_8822,N_7836,N_7853);
nor U8823 (N_8823,N_7389,N_7050);
and U8824 (N_8824,N_7654,N_7750);
or U8825 (N_8825,N_7157,N_7888);
nor U8826 (N_8826,N_7261,N_7051);
nor U8827 (N_8827,N_7024,N_7132);
or U8828 (N_8828,N_7632,N_7810);
nand U8829 (N_8829,N_7134,N_7160);
xnor U8830 (N_8830,N_7699,N_7767);
nand U8831 (N_8831,N_7337,N_7871);
nand U8832 (N_8832,N_7864,N_7317);
and U8833 (N_8833,N_7101,N_7361);
and U8834 (N_8834,N_7381,N_7760);
and U8835 (N_8835,N_7331,N_7805);
and U8836 (N_8836,N_7634,N_7512);
and U8837 (N_8837,N_7929,N_7814);
nor U8838 (N_8838,N_7718,N_7453);
nand U8839 (N_8839,N_7958,N_7754);
and U8840 (N_8840,N_7515,N_7090);
nor U8841 (N_8841,N_7298,N_7886);
and U8842 (N_8842,N_7829,N_7731);
xor U8843 (N_8843,N_7434,N_7097);
and U8844 (N_8844,N_7558,N_7756);
nor U8845 (N_8845,N_7575,N_7821);
and U8846 (N_8846,N_7058,N_7390);
and U8847 (N_8847,N_7468,N_7264);
or U8848 (N_8848,N_7500,N_7446);
nand U8849 (N_8849,N_7015,N_7813);
or U8850 (N_8850,N_7421,N_7349);
and U8851 (N_8851,N_7689,N_7763);
nor U8852 (N_8852,N_7998,N_7177);
or U8853 (N_8853,N_7317,N_7246);
nand U8854 (N_8854,N_7064,N_7089);
or U8855 (N_8855,N_7871,N_7463);
and U8856 (N_8856,N_7539,N_7106);
xnor U8857 (N_8857,N_7501,N_7452);
nand U8858 (N_8858,N_7885,N_7985);
nor U8859 (N_8859,N_7117,N_7936);
and U8860 (N_8860,N_7655,N_7442);
nor U8861 (N_8861,N_7645,N_7768);
and U8862 (N_8862,N_7875,N_7452);
nor U8863 (N_8863,N_7535,N_7809);
nand U8864 (N_8864,N_7508,N_7586);
xor U8865 (N_8865,N_7203,N_7485);
nand U8866 (N_8866,N_7686,N_7497);
nand U8867 (N_8867,N_7512,N_7438);
nor U8868 (N_8868,N_7780,N_7263);
xnor U8869 (N_8869,N_7308,N_7615);
or U8870 (N_8870,N_7576,N_7904);
nand U8871 (N_8871,N_7096,N_7193);
xor U8872 (N_8872,N_7603,N_7978);
xor U8873 (N_8873,N_7802,N_7588);
or U8874 (N_8874,N_7138,N_7785);
nor U8875 (N_8875,N_7278,N_7794);
or U8876 (N_8876,N_7055,N_7274);
nand U8877 (N_8877,N_7517,N_7024);
nor U8878 (N_8878,N_7314,N_7943);
xor U8879 (N_8879,N_7641,N_7274);
nand U8880 (N_8880,N_7142,N_7700);
or U8881 (N_8881,N_7285,N_7450);
nor U8882 (N_8882,N_7338,N_7219);
xnor U8883 (N_8883,N_7147,N_7201);
nand U8884 (N_8884,N_7540,N_7542);
nand U8885 (N_8885,N_7723,N_7176);
and U8886 (N_8886,N_7281,N_7818);
or U8887 (N_8887,N_7706,N_7612);
nand U8888 (N_8888,N_7333,N_7928);
xor U8889 (N_8889,N_7608,N_7539);
and U8890 (N_8890,N_7636,N_7411);
nand U8891 (N_8891,N_7968,N_7617);
nor U8892 (N_8892,N_7588,N_7377);
nor U8893 (N_8893,N_7503,N_7157);
and U8894 (N_8894,N_7354,N_7091);
nor U8895 (N_8895,N_7629,N_7285);
or U8896 (N_8896,N_7110,N_7137);
or U8897 (N_8897,N_7491,N_7433);
xor U8898 (N_8898,N_7011,N_7831);
nor U8899 (N_8899,N_7100,N_7005);
nand U8900 (N_8900,N_7371,N_7050);
xor U8901 (N_8901,N_7796,N_7077);
nor U8902 (N_8902,N_7230,N_7193);
xor U8903 (N_8903,N_7329,N_7528);
or U8904 (N_8904,N_7443,N_7576);
or U8905 (N_8905,N_7783,N_7406);
or U8906 (N_8906,N_7640,N_7630);
nand U8907 (N_8907,N_7246,N_7725);
nor U8908 (N_8908,N_7180,N_7396);
or U8909 (N_8909,N_7537,N_7008);
and U8910 (N_8910,N_7209,N_7359);
nand U8911 (N_8911,N_7156,N_7377);
nor U8912 (N_8912,N_7042,N_7128);
nand U8913 (N_8913,N_7603,N_7221);
xnor U8914 (N_8914,N_7803,N_7847);
xor U8915 (N_8915,N_7980,N_7164);
nand U8916 (N_8916,N_7109,N_7862);
and U8917 (N_8917,N_7158,N_7841);
or U8918 (N_8918,N_7502,N_7782);
xor U8919 (N_8919,N_7280,N_7878);
nor U8920 (N_8920,N_7994,N_7862);
and U8921 (N_8921,N_7354,N_7001);
or U8922 (N_8922,N_7271,N_7494);
and U8923 (N_8923,N_7359,N_7814);
nand U8924 (N_8924,N_7885,N_7139);
and U8925 (N_8925,N_7474,N_7042);
or U8926 (N_8926,N_7881,N_7137);
nor U8927 (N_8927,N_7938,N_7422);
nand U8928 (N_8928,N_7099,N_7284);
or U8929 (N_8929,N_7505,N_7392);
nand U8930 (N_8930,N_7141,N_7296);
xor U8931 (N_8931,N_7415,N_7361);
nor U8932 (N_8932,N_7314,N_7557);
nand U8933 (N_8933,N_7806,N_7064);
or U8934 (N_8934,N_7088,N_7358);
nor U8935 (N_8935,N_7679,N_7093);
nor U8936 (N_8936,N_7411,N_7686);
and U8937 (N_8937,N_7669,N_7733);
xnor U8938 (N_8938,N_7299,N_7653);
or U8939 (N_8939,N_7353,N_7811);
nor U8940 (N_8940,N_7816,N_7017);
xnor U8941 (N_8941,N_7960,N_7272);
and U8942 (N_8942,N_7834,N_7581);
nand U8943 (N_8943,N_7982,N_7905);
or U8944 (N_8944,N_7476,N_7675);
xnor U8945 (N_8945,N_7718,N_7128);
or U8946 (N_8946,N_7204,N_7753);
xnor U8947 (N_8947,N_7384,N_7232);
xor U8948 (N_8948,N_7812,N_7566);
nor U8949 (N_8949,N_7181,N_7729);
or U8950 (N_8950,N_7898,N_7791);
xor U8951 (N_8951,N_7134,N_7643);
xnor U8952 (N_8952,N_7514,N_7457);
nand U8953 (N_8953,N_7817,N_7246);
or U8954 (N_8954,N_7600,N_7191);
or U8955 (N_8955,N_7870,N_7191);
and U8956 (N_8956,N_7702,N_7440);
nor U8957 (N_8957,N_7623,N_7321);
nand U8958 (N_8958,N_7769,N_7766);
nor U8959 (N_8959,N_7770,N_7825);
xor U8960 (N_8960,N_7116,N_7189);
or U8961 (N_8961,N_7442,N_7224);
nor U8962 (N_8962,N_7267,N_7988);
xnor U8963 (N_8963,N_7968,N_7812);
or U8964 (N_8964,N_7041,N_7964);
or U8965 (N_8965,N_7613,N_7650);
xor U8966 (N_8966,N_7509,N_7294);
xor U8967 (N_8967,N_7874,N_7219);
or U8968 (N_8968,N_7881,N_7976);
and U8969 (N_8969,N_7776,N_7518);
and U8970 (N_8970,N_7832,N_7745);
nor U8971 (N_8971,N_7343,N_7439);
nand U8972 (N_8972,N_7774,N_7770);
nand U8973 (N_8973,N_7578,N_7701);
xor U8974 (N_8974,N_7435,N_7698);
xor U8975 (N_8975,N_7762,N_7151);
nand U8976 (N_8976,N_7906,N_7689);
nor U8977 (N_8977,N_7815,N_7786);
or U8978 (N_8978,N_7015,N_7091);
nand U8979 (N_8979,N_7906,N_7285);
xnor U8980 (N_8980,N_7565,N_7296);
nand U8981 (N_8981,N_7485,N_7484);
nand U8982 (N_8982,N_7322,N_7218);
or U8983 (N_8983,N_7768,N_7436);
nand U8984 (N_8984,N_7011,N_7707);
nand U8985 (N_8985,N_7615,N_7868);
nor U8986 (N_8986,N_7722,N_7703);
nand U8987 (N_8987,N_7145,N_7122);
xor U8988 (N_8988,N_7025,N_7210);
or U8989 (N_8989,N_7622,N_7798);
xnor U8990 (N_8990,N_7738,N_7606);
or U8991 (N_8991,N_7581,N_7772);
nand U8992 (N_8992,N_7809,N_7830);
xor U8993 (N_8993,N_7497,N_7098);
or U8994 (N_8994,N_7103,N_7727);
and U8995 (N_8995,N_7386,N_7843);
xor U8996 (N_8996,N_7243,N_7186);
or U8997 (N_8997,N_7892,N_7819);
nand U8998 (N_8998,N_7823,N_7487);
and U8999 (N_8999,N_7006,N_7340);
xor U9000 (N_9000,N_8054,N_8549);
nor U9001 (N_9001,N_8184,N_8430);
or U9002 (N_9002,N_8472,N_8438);
or U9003 (N_9003,N_8590,N_8098);
nand U9004 (N_9004,N_8761,N_8219);
xnor U9005 (N_9005,N_8035,N_8767);
nand U9006 (N_9006,N_8018,N_8450);
or U9007 (N_9007,N_8027,N_8447);
nand U9008 (N_9008,N_8819,N_8903);
nand U9009 (N_9009,N_8280,N_8000);
nor U9010 (N_9010,N_8374,N_8569);
and U9011 (N_9011,N_8502,N_8608);
or U9012 (N_9012,N_8799,N_8473);
and U9013 (N_9013,N_8227,N_8983);
or U9014 (N_9014,N_8157,N_8544);
and U9015 (N_9015,N_8200,N_8644);
xnor U9016 (N_9016,N_8727,N_8876);
nand U9017 (N_9017,N_8183,N_8164);
nand U9018 (N_9018,N_8631,N_8313);
nor U9019 (N_9019,N_8861,N_8193);
nor U9020 (N_9020,N_8724,N_8477);
nand U9021 (N_9021,N_8241,N_8225);
nand U9022 (N_9022,N_8902,N_8088);
nor U9023 (N_9023,N_8960,N_8664);
or U9024 (N_9024,N_8505,N_8422);
xnor U9025 (N_9025,N_8912,N_8776);
xnor U9026 (N_9026,N_8476,N_8714);
nand U9027 (N_9027,N_8595,N_8543);
nand U9028 (N_9028,N_8362,N_8316);
nor U9029 (N_9029,N_8262,N_8406);
and U9030 (N_9030,N_8479,N_8467);
nor U9031 (N_9031,N_8222,N_8182);
xnor U9032 (N_9032,N_8272,N_8626);
and U9033 (N_9033,N_8594,N_8787);
or U9034 (N_9034,N_8348,N_8548);
or U9035 (N_9035,N_8943,N_8809);
xor U9036 (N_9036,N_8329,N_8984);
and U9037 (N_9037,N_8743,N_8516);
xnor U9038 (N_9038,N_8640,N_8715);
and U9039 (N_9039,N_8305,N_8656);
nand U9040 (N_9040,N_8342,N_8730);
xnor U9041 (N_9041,N_8307,N_8791);
nor U9042 (N_9042,N_8519,N_8710);
nor U9043 (N_9043,N_8336,N_8042);
xnor U9044 (N_9044,N_8913,N_8132);
nand U9045 (N_9045,N_8366,N_8251);
nor U9046 (N_9046,N_8674,N_8199);
nor U9047 (N_9047,N_8794,N_8257);
xor U9048 (N_9048,N_8378,N_8442);
xnor U9049 (N_9049,N_8083,N_8289);
xnor U9050 (N_9050,N_8462,N_8385);
xnor U9051 (N_9051,N_8567,N_8056);
xnor U9052 (N_9052,N_8433,N_8793);
nor U9053 (N_9053,N_8552,N_8321);
or U9054 (N_9054,N_8732,N_8753);
nor U9055 (N_9055,N_8405,N_8437);
and U9056 (N_9056,N_8811,N_8972);
nor U9057 (N_9057,N_8883,N_8116);
and U9058 (N_9058,N_8250,N_8109);
and U9059 (N_9059,N_8151,N_8139);
and U9060 (N_9060,N_8512,N_8536);
nand U9061 (N_9061,N_8044,N_8330);
nor U9062 (N_9062,N_8518,N_8175);
and U9063 (N_9063,N_8621,N_8315);
nand U9064 (N_9064,N_8868,N_8103);
or U9065 (N_9065,N_8822,N_8360);
nor U9066 (N_9066,N_8739,N_8161);
xnor U9067 (N_9067,N_8844,N_8299);
and U9068 (N_9068,N_8154,N_8888);
nor U9069 (N_9069,N_8603,N_8410);
nor U9070 (N_9070,N_8852,N_8275);
nand U9071 (N_9071,N_8750,N_8345);
or U9072 (N_9072,N_8551,N_8005);
xnor U9073 (N_9073,N_8854,N_8185);
nand U9074 (N_9074,N_8741,N_8760);
nand U9075 (N_9075,N_8891,N_8464);
nand U9076 (N_9076,N_8547,N_8639);
and U9077 (N_9077,N_8525,N_8804);
nor U9078 (N_9078,N_8927,N_8441);
xor U9079 (N_9079,N_8818,N_8142);
or U9080 (N_9080,N_8038,N_8858);
and U9081 (N_9081,N_8504,N_8019);
and U9082 (N_9082,N_8254,N_8165);
xor U9083 (N_9083,N_8230,N_8465);
xor U9084 (N_9084,N_8559,N_8685);
or U9085 (N_9085,N_8343,N_8245);
nor U9086 (N_9086,N_8681,N_8720);
or U9087 (N_9087,N_8389,N_8179);
nand U9088 (N_9088,N_8436,N_8102);
and U9089 (N_9089,N_8700,N_8747);
and U9090 (N_9090,N_8783,N_8981);
and U9091 (N_9091,N_8218,N_8484);
or U9092 (N_9092,N_8381,N_8763);
nand U9093 (N_9093,N_8388,N_8428);
xnor U9094 (N_9094,N_8932,N_8668);
nand U9095 (N_9095,N_8082,N_8400);
xnor U9096 (N_9096,N_8453,N_8826);
or U9097 (N_9097,N_8337,N_8982);
and U9098 (N_9098,N_8662,N_8770);
xor U9099 (N_9099,N_8420,N_8751);
nor U9100 (N_9100,N_8106,N_8025);
nand U9101 (N_9101,N_8006,N_8539);
and U9102 (N_9102,N_8297,N_8521);
or U9103 (N_9103,N_8955,N_8276);
and U9104 (N_9104,N_8373,N_8119);
xor U9105 (N_9105,N_8703,N_8969);
or U9106 (N_9106,N_8115,N_8862);
or U9107 (N_9107,N_8253,N_8252);
xnor U9108 (N_9108,N_8424,N_8034);
nand U9109 (N_9109,N_8013,N_8153);
nand U9110 (N_9110,N_8769,N_8701);
nor U9111 (N_9111,N_8623,N_8234);
and U9112 (N_9112,N_8684,N_8789);
nor U9113 (N_9113,N_8050,N_8634);
nor U9114 (N_9114,N_8563,N_8650);
or U9115 (N_9115,N_8538,N_8093);
nor U9116 (N_9116,N_8863,N_8036);
nand U9117 (N_9117,N_8580,N_8210);
and U9118 (N_9118,N_8509,N_8152);
nor U9119 (N_9119,N_8768,N_8449);
and U9120 (N_9120,N_8470,N_8146);
and U9121 (N_9121,N_8849,N_8033);
xnor U9122 (N_9122,N_8215,N_8461);
xnor U9123 (N_9123,N_8775,N_8745);
nand U9124 (N_9124,N_8187,N_8718);
nor U9125 (N_9125,N_8244,N_8530);
nor U9126 (N_9126,N_8655,N_8945);
and U9127 (N_9127,N_8734,N_8797);
xor U9128 (N_9128,N_8211,N_8659);
nand U9129 (N_9129,N_8243,N_8309);
nor U9130 (N_9130,N_8810,N_8756);
or U9131 (N_9131,N_8398,N_8204);
nand U9132 (N_9132,N_8850,N_8779);
xnor U9133 (N_9133,N_8665,N_8875);
and U9134 (N_9134,N_8079,N_8369);
xnor U9135 (N_9135,N_8529,N_8326);
or U9136 (N_9136,N_8189,N_8292);
or U9137 (N_9137,N_8371,N_8113);
nand U9138 (N_9138,N_8556,N_8736);
xor U9139 (N_9139,N_8508,N_8300);
and U9140 (N_9140,N_8722,N_8795);
and U9141 (N_9141,N_8302,N_8625);
nor U9142 (N_9142,N_8452,N_8133);
and U9143 (N_9143,N_8125,N_8499);
nor U9144 (N_9144,N_8705,N_8843);
or U9145 (N_9145,N_8660,N_8416);
nor U9146 (N_9146,N_8711,N_8894);
xor U9147 (N_9147,N_8323,N_8361);
nand U9148 (N_9148,N_8490,N_8985);
and U9149 (N_9149,N_8459,N_8045);
xor U9150 (N_9150,N_8733,N_8240);
nor U9151 (N_9151,N_8568,N_8956);
and U9152 (N_9152,N_8906,N_8749);
and U9153 (N_9153,N_8387,N_8584);
or U9154 (N_9154,N_8706,N_8535);
nor U9155 (N_9155,N_8216,N_8319);
nor U9156 (N_9156,N_8936,N_8480);
nand U9157 (N_9157,N_8393,N_8010);
nand U9158 (N_9158,N_8454,N_8364);
and U9159 (N_9159,N_8952,N_8037);
and U9160 (N_9160,N_8628,N_8596);
nor U9161 (N_9161,N_8483,N_8865);
or U9162 (N_9162,N_8950,N_8589);
and U9163 (N_9163,N_8808,N_8448);
nand U9164 (N_9164,N_8399,N_8575);
or U9165 (N_9165,N_8560,N_8629);
nor U9166 (N_9166,N_8383,N_8231);
or U9167 (N_9167,N_8869,N_8758);
xnor U9168 (N_9168,N_8310,N_8021);
nor U9169 (N_9169,N_8764,N_8898);
nor U9170 (N_9170,N_8635,N_8813);
and U9171 (N_9171,N_8429,N_8517);
nand U9172 (N_9172,N_8900,N_8143);
xnor U9173 (N_9173,N_8110,N_8555);
and U9174 (N_9174,N_8682,N_8344);
or U9175 (N_9175,N_8221,N_8148);
and U9176 (N_9176,N_8944,N_8641);
nor U9177 (N_9177,N_8506,N_8412);
xnor U9178 (N_9178,N_8986,N_8408);
xor U9179 (N_9179,N_8100,N_8318);
nand U9180 (N_9180,N_8638,N_8007);
nor U9181 (N_9181,N_8637,N_8683);
nor U9182 (N_9182,N_8047,N_8306);
xor U9183 (N_9183,N_8778,N_8661);
nand U9184 (N_9184,N_8729,N_8600);
xor U9185 (N_9185,N_8966,N_8482);
and U9186 (N_9186,N_8991,N_8123);
and U9187 (N_9187,N_8238,N_8087);
nor U9188 (N_9188,N_8114,N_8150);
xnor U9189 (N_9189,N_8574,N_8823);
and U9190 (N_9190,N_8968,N_8213);
nor U9191 (N_9191,N_8877,N_8101);
xor U9192 (N_9192,N_8643,N_8825);
or U9193 (N_9193,N_8554,N_8848);
or U9194 (N_9194,N_8978,N_8909);
and U9195 (N_9195,N_8076,N_8582);
nand U9196 (N_9196,N_8857,N_8851);
or U9197 (N_9197,N_8766,N_8678);
nand U9198 (N_9198,N_8149,N_8120);
and U9199 (N_9199,N_8921,N_8587);
nor U9200 (N_9200,N_8949,N_8624);
nand U9201 (N_9201,N_8015,N_8919);
and U9202 (N_9202,N_8828,N_8558);
nor U9203 (N_9203,N_8691,N_8127);
nand U9204 (N_9204,N_8415,N_8217);
nand U9205 (N_9205,N_8759,N_8145);
and U9206 (N_9206,N_8016,N_8856);
or U9207 (N_9207,N_8256,N_8118);
nand U9208 (N_9208,N_8170,N_8014);
and U9209 (N_9209,N_8261,N_8924);
nor U9210 (N_9210,N_8180,N_8439);
xnor U9211 (N_9211,N_8553,N_8485);
and U9212 (N_9212,N_8277,N_8572);
nand U9213 (N_9213,N_8541,N_8062);
or U9214 (N_9214,N_8202,N_8896);
nor U9215 (N_9215,N_8395,N_8576);
nor U9216 (N_9216,N_8041,N_8586);
nand U9217 (N_9217,N_8820,N_8561);
or U9218 (N_9218,N_8488,N_8391);
xor U9219 (N_9219,N_8402,N_8377);
or U9220 (N_9220,N_8026,N_8993);
xor U9221 (N_9221,N_8455,N_8673);
or U9222 (N_9222,N_8012,N_8612);
nand U9223 (N_9223,N_8958,N_8075);
nand U9224 (N_9224,N_8686,N_8353);
nand U9225 (N_9225,N_8354,N_8957);
xnor U9226 (N_9226,N_8588,N_8288);
nor U9227 (N_9227,N_8141,N_8579);
xor U9228 (N_9228,N_8899,N_8872);
xor U9229 (N_9229,N_8676,N_8107);
and U9230 (N_9230,N_8397,N_8744);
nand U9231 (N_9231,N_8737,N_8039);
nand U9232 (N_9232,N_8649,N_8081);
and U9233 (N_9233,N_8959,N_8270);
and U9234 (N_9234,N_8267,N_8557);
nand U9235 (N_9235,N_8011,N_8937);
or U9236 (N_9236,N_8363,N_8847);
or U9237 (N_9237,N_8281,N_8071);
nand U9238 (N_9238,N_8537,N_8996);
nand U9239 (N_9239,N_8803,N_8597);
and U9240 (N_9240,N_8992,N_8265);
nor U9241 (N_9241,N_8610,N_8973);
or U9242 (N_9242,N_8717,N_8291);
xnor U9243 (N_9243,N_8178,N_8347);
and U9244 (N_9244,N_8435,N_8696);
and U9245 (N_9245,N_8740,N_8812);
xor U9246 (N_9246,N_8111,N_8266);
xnor U9247 (N_9247,N_8980,N_8024);
nor U9248 (N_9248,N_8147,N_8827);
or U9249 (N_9249,N_8162,N_8177);
nor U9250 (N_9250,N_8918,N_8772);
nand U9251 (N_9251,N_8156,N_8497);
nand U9252 (N_9252,N_8708,N_8492);
xor U9253 (N_9253,N_8104,N_8976);
nor U9254 (N_9254,N_8667,N_8771);
nor U9255 (N_9255,N_8995,N_8773);
nor U9256 (N_9256,N_8196,N_8534);
or U9257 (N_9257,N_8507,N_8786);
nand U9258 (N_9258,N_8694,N_8155);
or U9259 (N_9259,N_8494,N_8570);
and U9260 (N_9260,N_8846,N_8585);
or U9261 (N_9261,N_8020,N_8814);
nand U9262 (N_9262,N_8049,N_8721);
nand U9263 (N_9263,N_8379,N_8317);
nand U9264 (N_9264,N_8229,N_8889);
or U9265 (N_9265,N_8112,N_8444);
xnor U9266 (N_9266,N_8802,N_8839);
xor U9267 (N_9267,N_8788,N_8940);
nor U9268 (N_9268,N_8214,N_8524);
xor U9269 (N_9269,N_8648,N_8738);
xor U9270 (N_9270,N_8731,N_8800);
nor U9271 (N_9271,N_8440,N_8320);
or U9272 (N_9272,N_8333,N_8390);
nor U9273 (N_9273,N_8340,N_8432);
xor U9274 (N_9274,N_8908,N_8312);
or U9275 (N_9275,N_8458,N_8404);
nor U9276 (N_9276,N_8191,N_8293);
xnor U9277 (N_9277,N_8427,N_8475);
and U9278 (N_9278,N_8971,N_8785);
xnor U9279 (N_9279,N_8532,N_8201);
or U9280 (N_9280,N_8573,N_8815);
xor U9281 (N_9281,N_8942,N_8816);
xnor U9282 (N_9282,N_8346,N_8871);
or U9283 (N_9283,N_8070,N_8614);
nand U9284 (N_9284,N_8413,N_8606);
nand U9285 (N_9285,N_8097,N_8136);
or U9286 (N_9286,N_8953,N_8784);
xnor U9287 (N_9287,N_8002,N_8917);
or U9288 (N_9288,N_8206,N_8652);
nand U9289 (N_9289,N_8925,N_8471);
nor U9290 (N_9290,N_8247,N_8599);
xnor U9291 (N_9291,N_8613,N_8807);
nor U9292 (N_9292,N_8190,N_8571);
xor U9293 (N_9293,N_8181,N_8298);
or U9294 (N_9294,N_8274,N_8593);
and U9295 (N_9295,N_8618,N_8421);
nand U9296 (N_9296,N_8646,N_8542);
nand U9297 (N_9297,N_8294,N_8798);
xnor U9298 (N_9298,N_8121,N_8258);
nand U9299 (N_9299,N_8058,N_8495);
xnor U9300 (N_9300,N_8089,N_8284);
xor U9301 (N_9301,N_8457,N_8417);
nor U9302 (N_9302,N_8926,N_8840);
nor U9303 (N_9303,N_8975,N_8411);
xnor U9304 (N_9304,N_8583,N_8355);
and U9305 (N_9305,N_8263,N_8053);
and U9306 (N_9306,N_8642,N_8658);
xnor U9307 (N_9307,N_8987,N_8688);
nor U9308 (N_9308,N_8550,N_8084);
xnor U9309 (N_9309,N_8134,N_8609);
nand U9310 (N_9310,N_8777,N_8468);
nor U9311 (N_9311,N_8689,N_8365);
nand U9312 (N_9312,N_8707,N_8735);
nand U9313 (N_9313,N_8463,N_8370);
nand U9314 (N_9314,N_8237,N_8781);
nor U9315 (N_9315,N_8223,N_8994);
and U9316 (N_9316,N_8334,N_8564);
nand U9317 (N_9317,N_8273,N_8043);
nor U9318 (N_9318,N_8748,N_8260);
and U9319 (N_9319,N_8964,N_8286);
nand U9320 (N_9320,N_8954,N_8630);
or U9321 (N_9321,N_8419,N_8842);
nor U9322 (N_9322,N_8086,N_8030);
nand U9323 (N_9323,N_8526,N_8545);
or U9324 (N_9324,N_8515,N_8128);
nand U9325 (N_9325,N_8914,N_8726);
nor U9326 (N_9326,N_8126,N_8746);
or U9327 (N_9327,N_8922,N_8094);
nor U9328 (N_9328,N_8672,N_8870);
or U9329 (N_9329,N_8878,N_8817);
xor U9330 (N_9330,N_8832,N_8999);
and U9331 (N_9331,N_8893,N_8308);
nor U9332 (N_9332,N_8144,N_8742);
and U9333 (N_9333,N_8931,N_8752);
or U9334 (N_9334,N_8008,N_8375);
nor U9335 (N_9335,N_8176,N_8066);
nand U9336 (N_9336,N_8915,N_8009);
nand U9337 (N_9337,N_8709,N_8074);
nand U9338 (N_9338,N_8531,N_8301);
and U9339 (N_9339,N_8311,N_8616);
or U9340 (N_9340,N_8208,N_8853);
nor U9341 (N_9341,N_8137,N_8693);
nand U9342 (N_9342,N_8910,N_8834);
nor U9343 (N_9343,N_8657,N_8687);
or U9344 (N_9344,N_8224,N_8394);
nor U9345 (N_9345,N_8129,N_8500);
or U9346 (N_9346,N_8063,N_8998);
xnor U9347 (N_9347,N_8017,N_8117);
xor U9348 (N_9348,N_8061,N_8423);
or U9349 (N_9349,N_8029,N_8278);
or U9350 (N_9350,N_8099,N_8496);
nand U9351 (N_9351,N_8431,N_8407);
and U9352 (N_9352,N_8974,N_8633);
nor U9353 (N_9353,N_8255,N_8719);
xnor U9354 (N_9354,N_8615,N_8796);
xor U9355 (N_9355,N_8203,N_8287);
xnor U9356 (N_9356,N_8669,N_8904);
or U9357 (N_9357,N_8474,N_8867);
nand U9358 (N_9358,N_8085,N_8124);
and U9359 (N_9359,N_8031,N_8384);
nand U9360 (N_9360,N_8282,N_8907);
or U9361 (N_9361,N_8935,N_8269);
nand U9362 (N_9362,N_8328,N_8692);
and U9363 (N_9363,N_8057,N_8478);
nand U9364 (N_9364,N_8723,N_8386);
and U9365 (N_9365,N_8122,N_8528);
nand U9366 (N_9366,N_8946,N_8205);
or U9367 (N_9367,N_8220,N_8283);
nand U9368 (N_9368,N_8514,N_8882);
nor U9369 (N_9369,N_8414,N_8533);
and U9370 (N_9370,N_8947,N_8911);
xor U9371 (N_9371,N_8879,N_8716);
and U9372 (N_9372,N_8977,N_8829);
nand U9373 (N_9373,N_8704,N_8249);
nand U9374 (N_9374,N_8651,N_8138);
xor U9375 (N_9375,N_8171,N_8671);
xnor U9376 (N_9376,N_8068,N_8067);
xnor U9377 (N_9377,N_8501,N_8352);
and U9378 (N_9378,N_8460,N_8698);
and U9379 (N_9379,N_8916,N_8236);
and U9380 (N_9380,N_8527,N_8513);
nand U9381 (N_9381,N_8368,N_8358);
and U9382 (N_9382,N_8697,N_8591);
or U9383 (N_9383,N_8197,N_8690);
and U9384 (N_9384,N_8860,N_8351);
and U9385 (N_9385,N_8290,N_8451);
or U9386 (N_9386,N_8108,N_8059);
or U9387 (N_9387,N_8491,N_8754);
nand U9388 (N_9388,N_8755,N_8774);
xnor U9389 (N_9389,N_8679,N_8356);
and U9390 (N_9390,N_8617,N_8792);
and U9391 (N_9391,N_8886,N_8418);
nand U9392 (N_9392,N_8065,N_8699);
and U9393 (N_9393,N_8670,N_8930);
nor U9394 (N_9394,N_8077,N_8443);
nand U9395 (N_9395,N_8228,N_8166);
nor U9396 (N_9396,N_8824,N_8341);
nand U9397 (N_9397,N_8855,N_8296);
nor U9398 (N_9398,N_8434,N_8578);
xnor U9399 (N_9399,N_8096,N_8801);
nor U9400 (N_9400,N_8131,N_8967);
xor U9401 (N_9401,N_8695,N_8663);
and U9402 (N_9402,N_8173,N_8169);
and U9403 (N_9403,N_8680,N_8090);
and U9404 (N_9404,N_8226,N_8324);
nor U9405 (N_9405,N_8051,N_8592);
xnor U9406 (N_9406,N_8446,N_8622);
nor U9407 (N_9407,N_8890,N_8577);
nand U9408 (N_9408,N_8604,N_8990);
xor U9409 (N_9409,N_8350,N_8487);
xor U9410 (N_9410,N_8757,N_8607);
xnor U9411 (N_9411,N_8004,N_8052);
xor U9412 (N_9412,N_8396,N_8831);
nor U9413 (N_9413,N_8409,N_8881);
nor U9414 (N_9414,N_8163,N_8359);
nand U9415 (N_9415,N_8702,N_8259);
and U9416 (N_9416,N_8264,N_8080);
and U9417 (N_9417,N_8445,N_8835);
xor U9418 (N_9418,N_8546,N_8962);
and U9419 (N_9419,N_8928,N_8765);
xnor U9420 (N_9420,N_8022,N_8489);
or U9421 (N_9421,N_8158,N_8327);
nor U9422 (N_9422,N_8195,N_8790);
nand U9423 (N_9423,N_8837,N_8522);
and U9424 (N_9424,N_8920,N_8885);
or U9425 (N_9425,N_8929,N_8905);
nand U9426 (N_9426,N_8939,N_8469);
xor U9427 (N_9427,N_8965,N_8520);
and U9428 (N_9428,N_8105,N_8897);
nand U9429 (N_9429,N_8160,N_8988);
or U9430 (N_9430,N_8159,N_8271);
or U9431 (N_9431,N_8069,N_8239);
xnor U9432 (N_9432,N_8503,N_8979);
or U9433 (N_9433,N_8295,N_8841);
nand U9434 (N_9434,N_8232,N_8782);
and U9435 (N_9435,N_8647,N_8540);
nor U9436 (N_9436,N_8095,N_8493);
or U9437 (N_9437,N_8620,N_8268);
xnor U9438 (N_9438,N_8078,N_8401);
nor U9439 (N_9439,N_8632,N_8023);
nor U9440 (N_9440,N_8498,N_8970);
xor U9441 (N_9441,N_8725,N_8285);
nand U9442 (N_9442,N_8892,N_8140);
or U9443 (N_9443,N_8713,N_8895);
nand U9444 (N_9444,N_8923,N_8997);
or U9445 (N_9445,N_8174,N_8339);
xnor U9446 (N_9446,N_8880,N_8188);
or U9447 (N_9447,N_8873,N_8963);
xnor U9448 (N_9448,N_8866,N_8510);
or U9449 (N_9449,N_8581,N_8332);
nand U9450 (N_9450,N_8091,N_8933);
or U9451 (N_9451,N_8887,N_8060);
and U9452 (N_9452,N_8314,N_8864);
nand U9453 (N_9453,N_8601,N_8565);
xnor U9454 (N_9454,N_8349,N_8675);
and U9455 (N_9455,N_8335,N_8466);
and U9456 (N_9456,N_8961,N_8192);
xnor U9457 (N_9457,N_8938,N_8653);
or U9458 (N_9458,N_8279,N_8073);
nor U9459 (N_9459,N_8627,N_8304);
nand U9460 (N_9460,N_8830,N_8836);
xor U9461 (N_9461,N_8248,N_8845);
nand U9462 (N_9462,N_8130,N_8805);
and U9463 (N_9463,N_8762,N_8046);
and U9464 (N_9464,N_8666,N_8380);
nand U9465 (N_9465,N_8948,N_8611);
nand U9466 (N_9466,N_8048,N_8001);
nor U9467 (N_9467,N_8194,N_8357);
nor U9468 (N_9468,N_8951,N_8092);
nor U9469 (N_9469,N_8322,N_8989);
xnor U9470 (N_9470,N_8456,N_8172);
nand U9471 (N_9471,N_8198,N_8135);
nand U9472 (N_9472,N_8806,N_8403);
nand U9473 (N_9473,N_8003,N_8654);
nand U9474 (N_9474,N_8712,N_8833);
and U9475 (N_9475,N_8246,N_8376);
and U9476 (N_9476,N_8367,N_8838);
nor U9477 (N_9477,N_8168,N_8372);
xor U9478 (N_9478,N_8032,N_8392);
xnor U9479 (N_9479,N_8055,N_8859);
nor U9480 (N_9480,N_8728,N_8821);
nand U9481 (N_9481,N_8207,N_8934);
or U9482 (N_9482,N_8064,N_8481);
and U9483 (N_9483,N_8209,N_8780);
nor U9484 (N_9484,N_8235,N_8598);
nor U9485 (N_9485,N_8486,N_8212);
nor U9486 (N_9486,N_8874,N_8242);
xnor U9487 (N_9487,N_8426,N_8425);
nand U9488 (N_9488,N_8186,N_8325);
nand U9489 (N_9489,N_8040,N_8382);
nor U9490 (N_9490,N_8901,N_8167);
xor U9491 (N_9491,N_8619,N_8511);
or U9492 (N_9492,N_8028,N_8941);
xnor U9493 (N_9493,N_8233,N_8677);
nor U9494 (N_9494,N_8303,N_8884);
nand U9495 (N_9495,N_8338,N_8523);
nand U9496 (N_9496,N_8566,N_8605);
or U9497 (N_9497,N_8331,N_8072);
xor U9498 (N_9498,N_8636,N_8645);
nor U9499 (N_9499,N_8562,N_8602);
nand U9500 (N_9500,N_8983,N_8330);
or U9501 (N_9501,N_8770,N_8645);
xor U9502 (N_9502,N_8849,N_8858);
and U9503 (N_9503,N_8989,N_8710);
and U9504 (N_9504,N_8421,N_8265);
nand U9505 (N_9505,N_8493,N_8818);
and U9506 (N_9506,N_8335,N_8319);
nand U9507 (N_9507,N_8107,N_8197);
xnor U9508 (N_9508,N_8282,N_8567);
nor U9509 (N_9509,N_8535,N_8420);
nand U9510 (N_9510,N_8873,N_8502);
xnor U9511 (N_9511,N_8866,N_8749);
or U9512 (N_9512,N_8696,N_8910);
and U9513 (N_9513,N_8102,N_8035);
and U9514 (N_9514,N_8393,N_8470);
nor U9515 (N_9515,N_8675,N_8405);
xor U9516 (N_9516,N_8443,N_8843);
and U9517 (N_9517,N_8030,N_8777);
nor U9518 (N_9518,N_8436,N_8953);
or U9519 (N_9519,N_8988,N_8803);
nand U9520 (N_9520,N_8345,N_8344);
nor U9521 (N_9521,N_8656,N_8261);
and U9522 (N_9522,N_8819,N_8915);
or U9523 (N_9523,N_8520,N_8769);
or U9524 (N_9524,N_8396,N_8176);
or U9525 (N_9525,N_8899,N_8333);
xor U9526 (N_9526,N_8362,N_8645);
xnor U9527 (N_9527,N_8706,N_8024);
and U9528 (N_9528,N_8966,N_8524);
nand U9529 (N_9529,N_8820,N_8276);
nand U9530 (N_9530,N_8732,N_8943);
nand U9531 (N_9531,N_8296,N_8896);
xor U9532 (N_9532,N_8030,N_8478);
xnor U9533 (N_9533,N_8091,N_8887);
nor U9534 (N_9534,N_8830,N_8866);
nand U9535 (N_9535,N_8278,N_8314);
nand U9536 (N_9536,N_8614,N_8252);
nand U9537 (N_9537,N_8604,N_8912);
nand U9538 (N_9538,N_8662,N_8489);
or U9539 (N_9539,N_8262,N_8145);
and U9540 (N_9540,N_8262,N_8479);
nor U9541 (N_9541,N_8521,N_8731);
nor U9542 (N_9542,N_8616,N_8410);
or U9543 (N_9543,N_8234,N_8576);
xnor U9544 (N_9544,N_8636,N_8245);
xor U9545 (N_9545,N_8491,N_8123);
xnor U9546 (N_9546,N_8112,N_8925);
xor U9547 (N_9547,N_8291,N_8310);
xor U9548 (N_9548,N_8834,N_8866);
and U9549 (N_9549,N_8361,N_8647);
or U9550 (N_9550,N_8211,N_8144);
or U9551 (N_9551,N_8535,N_8875);
nand U9552 (N_9552,N_8528,N_8704);
and U9553 (N_9553,N_8823,N_8798);
nor U9554 (N_9554,N_8633,N_8049);
and U9555 (N_9555,N_8609,N_8012);
xor U9556 (N_9556,N_8674,N_8645);
or U9557 (N_9557,N_8208,N_8358);
nor U9558 (N_9558,N_8345,N_8999);
and U9559 (N_9559,N_8725,N_8850);
or U9560 (N_9560,N_8315,N_8302);
or U9561 (N_9561,N_8964,N_8425);
and U9562 (N_9562,N_8028,N_8691);
and U9563 (N_9563,N_8515,N_8576);
or U9564 (N_9564,N_8697,N_8133);
or U9565 (N_9565,N_8438,N_8582);
xnor U9566 (N_9566,N_8291,N_8777);
nand U9567 (N_9567,N_8401,N_8597);
nand U9568 (N_9568,N_8925,N_8150);
xnor U9569 (N_9569,N_8424,N_8554);
and U9570 (N_9570,N_8487,N_8231);
and U9571 (N_9571,N_8028,N_8207);
xnor U9572 (N_9572,N_8691,N_8918);
nor U9573 (N_9573,N_8368,N_8040);
xnor U9574 (N_9574,N_8833,N_8308);
xor U9575 (N_9575,N_8039,N_8719);
and U9576 (N_9576,N_8202,N_8545);
nand U9577 (N_9577,N_8919,N_8428);
xor U9578 (N_9578,N_8591,N_8174);
and U9579 (N_9579,N_8841,N_8153);
and U9580 (N_9580,N_8930,N_8362);
and U9581 (N_9581,N_8105,N_8860);
and U9582 (N_9582,N_8229,N_8004);
or U9583 (N_9583,N_8049,N_8941);
and U9584 (N_9584,N_8257,N_8159);
nor U9585 (N_9585,N_8553,N_8410);
nand U9586 (N_9586,N_8488,N_8829);
xor U9587 (N_9587,N_8316,N_8997);
and U9588 (N_9588,N_8390,N_8373);
and U9589 (N_9589,N_8636,N_8196);
xor U9590 (N_9590,N_8354,N_8881);
or U9591 (N_9591,N_8312,N_8893);
and U9592 (N_9592,N_8595,N_8420);
xnor U9593 (N_9593,N_8845,N_8559);
and U9594 (N_9594,N_8209,N_8394);
xor U9595 (N_9595,N_8809,N_8915);
or U9596 (N_9596,N_8392,N_8257);
xnor U9597 (N_9597,N_8671,N_8861);
nand U9598 (N_9598,N_8095,N_8695);
and U9599 (N_9599,N_8566,N_8986);
or U9600 (N_9600,N_8077,N_8464);
xnor U9601 (N_9601,N_8035,N_8489);
or U9602 (N_9602,N_8466,N_8733);
and U9603 (N_9603,N_8880,N_8146);
nor U9604 (N_9604,N_8575,N_8545);
and U9605 (N_9605,N_8724,N_8727);
nor U9606 (N_9606,N_8441,N_8503);
xor U9607 (N_9607,N_8773,N_8523);
and U9608 (N_9608,N_8589,N_8404);
nand U9609 (N_9609,N_8609,N_8081);
nand U9610 (N_9610,N_8671,N_8062);
nand U9611 (N_9611,N_8803,N_8593);
or U9612 (N_9612,N_8274,N_8336);
or U9613 (N_9613,N_8359,N_8219);
nor U9614 (N_9614,N_8294,N_8996);
nor U9615 (N_9615,N_8959,N_8374);
and U9616 (N_9616,N_8504,N_8124);
nand U9617 (N_9617,N_8193,N_8063);
nand U9618 (N_9618,N_8514,N_8153);
and U9619 (N_9619,N_8351,N_8996);
xor U9620 (N_9620,N_8870,N_8509);
nand U9621 (N_9621,N_8882,N_8533);
nor U9622 (N_9622,N_8760,N_8410);
and U9623 (N_9623,N_8899,N_8127);
nor U9624 (N_9624,N_8502,N_8719);
xnor U9625 (N_9625,N_8998,N_8567);
and U9626 (N_9626,N_8947,N_8985);
xor U9627 (N_9627,N_8843,N_8342);
nand U9628 (N_9628,N_8867,N_8824);
and U9629 (N_9629,N_8828,N_8365);
and U9630 (N_9630,N_8941,N_8414);
and U9631 (N_9631,N_8760,N_8744);
and U9632 (N_9632,N_8520,N_8423);
xor U9633 (N_9633,N_8086,N_8385);
or U9634 (N_9634,N_8771,N_8022);
nor U9635 (N_9635,N_8571,N_8530);
nor U9636 (N_9636,N_8312,N_8225);
nor U9637 (N_9637,N_8204,N_8702);
xor U9638 (N_9638,N_8738,N_8271);
nand U9639 (N_9639,N_8513,N_8975);
nor U9640 (N_9640,N_8593,N_8586);
or U9641 (N_9641,N_8374,N_8876);
and U9642 (N_9642,N_8859,N_8594);
and U9643 (N_9643,N_8695,N_8949);
xor U9644 (N_9644,N_8939,N_8401);
and U9645 (N_9645,N_8180,N_8912);
nor U9646 (N_9646,N_8176,N_8514);
nor U9647 (N_9647,N_8625,N_8479);
nand U9648 (N_9648,N_8406,N_8067);
nand U9649 (N_9649,N_8812,N_8832);
xor U9650 (N_9650,N_8376,N_8558);
xor U9651 (N_9651,N_8458,N_8494);
and U9652 (N_9652,N_8346,N_8587);
xor U9653 (N_9653,N_8469,N_8758);
nand U9654 (N_9654,N_8111,N_8056);
nor U9655 (N_9655,N_8076,N_8267);
nor U9656 (N_9656,N_8730,N_8007);
and U9657 (N_9657,N_8683,N_8983);
xor U9658 (N_9658,N_8177,N_8105);
nand U9659 (N_9659,N_8179,N_8758);
and U9660 (N_9660,N_8328,N_8225);
or U9661 (N_9661,N_8304,N_8470);
or U9662 (N_9662,N_8587,N_8113);
nor U9663 (N_9663,N_8396,N_8156);
xor U9664 (N_9664,N_8252,N_8800);
nor U9665 (N_9665,N_8813,N_8801);
xor U9666 (N_9666,N_8706,N_8680);
or U9667 (N_9667,N_8264,N_8705);
nor U9668 (N_9668,N_8977,N_8444);
xor U9669 (N_9669,N_8368,N_8975);
xnor U9670 (N_9670,N_8902,N_8184);
and U9671 (N_9671,N_8392,N_8536);
and U9672 (N_9672,N_8206,N_8927);
nand U9673 (N_9673,N_8672,N_8583);
or U9674 (N_9674,N_8257,N_8372);
or U9675 (N_9675,N_8127,N_8362);
nor U9676 (N_9676,N_8027,N_8669);
xnor U9677 (N_9677,N_8722,N_8753);
nand U9678 (N_9678,N_8479,N_8350);
nor U9679 (N_9679,N_8263,N_8573);
nand U9680 (N_9680,N_8936,N_8727);
or U9681 (N_9681,N_8888,N_8624);
nor U9682 (N_9682,N_8944,N_8032);
or U9683 (N_9683,N_8054,N_8434);
nor U9684 (N_9684,N_8222,N_8066);
or U9685 (N_9685,N_8167,N_8083);
or U9686 (N_9686,N_8568,N_8271);
nor U9687 (N_9687,N_8332,N_8707);
nand U9688 (N_9688,N_8348,N_8158);
nand U9689 (N_9689,N_8735,N_8250);
nor U9690 (N_9690,N_8024,N_8729);
or U9691 (N_9691,N_8822,N_8217);
and U9692 (N_9692,N_8043,N_8172);
xor U9693 (N_9693,N_8391,N_8147);
nor U9694 (N_9694,N_8053,N_8682);
and U9695 (N_9695,N_8490,N_8262);
or U9696 (N_9696,N_8819,N_8561);
nand U9697 (N_9697,N_8199,N_8450);
xor U9698 (N_9698,N_8835,N_8130);
xor U9699 (N_9699,N_8208,N_8304);
xnor U9700 (N_9700,N_8333,N_8645);
or U9701 (N_9701,N_8384,N_8296);
nand U9702 (N_9702,N_8538,N_8428);
xnor U9703 (N_9703,N_8264,N_8357);
and U9704 (N_9704,N_8978,N_8754);
xnor U9705 (N_9705,N_8598,N_8385);
nand U9706 (N_9706,N_8436,N_8447);
nand U9707 (N_9707,N_8672,N_8692);
xor U9708 (N_9708,N_8729,N_8581);
nor U9709 (N_9709,N_8814,N_8164);
or U9710 (N_9710,N_8479,N_8937);
nand U9711 (N_9711,N_8292,N_8856);
nand U9712 (N_9712,N_8657,N_8511);
nand U9713 (N_9713,N_8516,N_8707);
nand U9714 (N_9714,N_8151,N_8788);
nand U9715 (N_9715,N_8388,N_8913);
and U9716 (N_9716,N_8020,N_8112);
or U9717 (N_9717,N_8372,N_8665);
or U9718 (N_9718,N_8971,N_8243);
or U9719 (N_9719,N_8869,N_8914);
nand U9720 (N_9720,N_8957,N_8664);
xor U9721 (N_9721,N_8555,N_8128);
or U9722 (N_9722,N_8234,N_8705);
nand U9723 (N_9723,N_8790,N_8939);
xor U9724 (N_9724,N_8910,N_8479);
and U9725 (N_9725,N_8153,N_8336);
nor U9726 (N_9726,N_8544,N_8976);
and U9727 (N_9727,N_8229,N_8907);
nand U9728 (N_9728,N_8385,N_8542);
xor U9729 (N_9729,N_8566,N_8827);
and U9730 (N_9730,N_8703,N_8779);
or U9731 (N_9731,N_8630,N_8162);
nand U9732 (N_9732,N_8779,N_8795);
nand U9733 (N_9733,N_8741,N_8461);
nand U9734 (N_9734,N_8752,N_8337);
nand U9735 (N_9735,N_8322,N_8236);
or U9736 (N_9736,N_8458,N_8479);
and U9737 (N_9737,N_8515,N_8531);
nor U9738 (N_9738,N_8221,N_8561);
nand U9739 (N_9739,N_8197,N_8353);
nand U9740 (N_9740,N_8327,N_8624);
nor U9741 (N_9741,N_8582,N_8412);
nand U9742 (N_9742,N_8608,N_8655);
or U9743 (N_9743,N_8554,N_8761);
or U9744 (N_9744,N_8824,N_8513);
or U9745 (N_9745,N_8206,N_8960);
or U9746 (N_9746,N_8808,N_8421);
nand U9747 (N_9747,N_8587,N_8633);
xnor U9748 (N_9748,N_8701,N_8616);
xnor U9749 (N_9749,N_8498,N_8060);
xor U9750 (N_9750,N_8213,N_8440);
xnor U9751 (N_9751,N_8768,N_8706);
xor U9752 (N_9752,N_8851,N_8764);
nor U9753 (N_9753,N_8192,N_8924);
nand U9754 (N_9754,N_8966,N_8509);
xor U9755 (N_9755,N_8042,N_8977);
nand U9756 (N_9756,N_8048,N_8310);
and U9757 (N_9757,N_8456,N_8318);
and U9758 (N_9758,N_8319,N_8842);
or U9759 (N_9759,N_8767,N_8223);
nor U9760 (N_9760,N_8341,N_8587);
nand U9761 (N_9761,N_8619,N_8236);
or U9762 (N_9762,N_8560,N_8988);
nor U9763 (N_9763,N_8861,N_8867);
nand U9764 (N_9764,N_8059,N_8237);
nand U9765 (N_9765,N_8128,N_8361);
nand U9766 (N_9766,N_8941,N_8320);
xnor U9767 (N_9767,N_8189,N_8758);
or U9768 (N_9768,N_8228,N_8021);
and U9769 (N_9769,N_8049,N_8013);
or U9770 (N_9770,N_8419,N_8467);
or U9771 (N_9771,N_8592,N_8244);
and U9772 (N_9772,N_8275,N_8499);
xor U9773 (N_9773,N_8883,N_8595);
and U9774 (N_9774,N_8438,N_8731);
or U9775 (N_9775,N_8226,N_8700);
xnor U9776 (N_9776,N_8241,N_8129);
xnor U9777 (N_9777,N_8608,N_8864);
or U9778 (N_9778,N_8736,N_8933);
xor U9779 (N_9779,N_8062,N_8046);
xnor U9780 (N_9780,N_8272,N_8329);
and U9781 (N_9781,N_8563,N_8679);
or U9782 (N_9782,N_8228,N_8698);
nand U9783 (N_9783,N_8403,N_8027);
or U9784 (N_9784,N_8297,N_8114);
and U9785 (N_9785,N_8898,N_8399);
nand U9786 (N_9786,N_8348,N_8855);
and U9787 (N_9787,N_8489,N_8877);
nor U9788 (N_9788,N_8688,N_8239);
nand U9789 (N_9789,N_8559,N_8474);
or U9790 (N_9790,N_8639,N_8984);
nand U9791 (N_9791,N_8670,N_8897);
xnor U9792 (N_9792,N_8718,N_8684);
xor U9793 (N_9793,N_8321,N_8967);
xor U9794 (N_9794,N_8371,N_8046);
and U9795 (N_9795,N_8138,N_8029);
nand U9796 (N_9796,N_8108,N_8136);
xor U9797 (N_9797,N_8856,N_8148);
xor U9798 (N_9798,N_8126,N_8464);
xor U9799 (N_9799,N_8056,N_8160);
or U9800 (N_9800,N_8803,N_8418);
and U9801 (N_9801,N_8637,N_8621);
xor U9802 (N_9802,N_8010,N_8570);
and U9803 (N_9803,N_8768,N_8095);
nor U9804 (N_9804,N_8127,N_8651);
xor U9805 (N_9805,N_8894,N_8544);
nor U9806 (N_9806,N_8070,N_8837);
and U9807 (N_9807,N_8821,N_8844);
and U9808 (N_9808,N_8182,N_8808);
nand U9809 (N_9809,N_8770,N_8632);
and U9810 (N_9810,N_8783,N_8825);
nand U9811 (N_9811,N_8582,N_8777);
or U9812 (N_9812,N_8109,N_8768);
xnor U9813 (N_9813,N_8899,N_8513);
or U9814 (N_9814,N_8954,N_8224);
xnor U9815 (N_9815,N_8968,N_8664);
xnor U9816 (N_9816,N_8245,N_8762);
or U9817 (N_9817,N_8886,N_8901);
or U9818 (N_9818,N_8854,N_8955);
or U9819 (N_9819,N_8569,N_8121);
nor U9820 (N_9820,N_8817,N_8094);
nor U9821 (N_9821,N_8910,N_8308);
nand U9822 (N_9822,N_8082,N_8486);
or U9823 (N_9823,N_8952,N_8824);
or U9824 (N_9824,N_8156,N_8645);
or U9825 (N_9825,N_8760,N_8222);
nor U9826 (N_9826,N_8661,N_8914);
nor U9827 (N_9827,N_8515,N_8481);
and U9828 (N_9828,N_8484,N_8516);
nand U9829 (N_9829,N_8563,N_8097);
and U9830 (N_9830,N_8481,N_8462);
xor U9831 (N_9831,N_8980,N_8676);
or U9832 (N_9832,N_8011,N_8108);
and U9833 (N_9833,N_8158,N_8393);
or U9834 (N_9834,N_8075,N_8336);
nand U9835 (N_9835,N_8544,N_8535);
nor U9836 (N_9836,N_8790,N_8012);
and U9837 (N_9837,N_8341,N_8633);
or U9838 (N_9838,N_8359,N_8871);
nand U9839 (N_9839,N_8775,N_8485);
nor U9840 (N_9840,N_8874,N_8296);
nand U9841 (N_9841,N_8026,N_8173);
nor U9842 (N_9842,N_8463,N_8339);
and U9843 (N_9843,N_8657,N_8002);
or U9844 (N_9844,N_8986,N_8765);
nand U9845 (N_9845,N_8223,N_8124);
or U9846 (N_9846,N_8853,N_8392);
and U9847 (N_9847,N_8322,N_8894);
xor U9848 (N_9848,N_8424,N_8233);
nand U9849 (N_9849,N_8496,N_8633);
xnor U9850 (N_9850,N_8907,N_8414);
and U9851 (N_9851,N_8655,N_8752);
and U9852 (N_9852,N_8948,N_8396);
and U9853 (N_9853,N_8367,N_8217);
and U9854 (N_9854,N_8739,N_8703);
nor U9855 (N_9855,N_8288,N_8495);
nand U9856 (N_9856,N_8054,N_8550);
xor U9857 (N_9857,N_8341,N_8577);
nor U9858 (N_9858,N_8001,N_8155);
nand U9859 (N_9859,N_8119,N_8104);
or U9860 (N_9860,N_8621,N_8178);
nor U9861 (N_9861,N_8470,N_8058);
and U9862 (N_9862,N_8778,N_8479);
nand U9863 (N_9863,N_8966,N_8512);
and U9864 (N_9864,N_8730,N_8286);
nor U9865 (N_9865,N_8134,N_8914);
and U9866 (N_9866,N_8040,N_8524);
xor U9867 (N_9867,N_8113,N_8473);
xnor U9868 (N_9868,N_8657,N_8421);
nor U9869 (N_9869,N_8878,N_8668);
nand U9870 (N_9870,N_8402,N_8626);
nor U9871 (N_9871,N_8752,N_8528);
nand U9872 (N_9872,N_8956,N_8903);
nand U9873 (N_9873,N_8267,N_8648);
nand U9874 (N_9874,N_8399,N_8049);
nand U9875 (N_9875,N_8466,N_8610);
nand U9876 (N_9876,N_8719,N_8636);
nand U9877 (N_9877,N_8637,N_8012);
nand U9878 (N_9878,N_8522,N_8732);
nor U9879 (N_9879,N_8240,N_8159);
or U9880 (N_9880,N_8022,N_8937);
and U9881 (N_9881,N_8144,N_8953);
nor U9882 (N_9882,N_8042,N_8724);
or U9883 (N_9883,N_8297,N_8794);
nor U9884 (N_9884,N_8722,N_8446);
nor U9885 (N_9885,N_8877,N_8370);
and U9886 (N_9886,N_8808,N_8298);
nand U9887 (N_9887,N_8495,N_8878);
or U9888 (N_9888,N_8236,N_8029);
xnor U9889 (N_9889,N_8657,N_8374);
xnor U9890 (N_9890,N_8330,N_8012);
or U9891 (N_9891,N_8410,N_8402);
xnor U9892 (N_9892,N_8746,N_8904);
and U9893 (N_9893,N_8274,N_8418);
and U9894 (N_9894,N_8585,N_8633);
nand U9895 (N_9895,N_8034,N_8129);
and U9896 (N_9896,N_8233,N_8415);
nand U9897 (N_9897,N_8782,N_8071);
or U9898 (N_9898,N_8846,N_8899);
nand U9899 (N_9899,N_8321,N_8896);
nand U9900 (N_9900,N_8166,N_8908);
nand U9901 (N_9901,N_8057,N_8304);
nor U9902 (N_9902,N_8564,N_8873);
or U9903 (N_9903,N_8209,N_8971);
nand U9904 (N_9904,N_8627,N_8858);
nand U9905 (N_9905,N_8588,N_8233);
nor U9906 (N_9906,N_8785,N_8375);
xnor U9907 (N_9907,N_8192,N_8271);
or U9908 (N_9908,N_8693,N_8184);
xnor U9909 (N_9909,N_8737,N_8989);
and U9910 (N_9910,N_8955,N_8424);
xnor U9911 (N_9911,N_8754,N_8171);
or U9912 (N_9912,N_8119,N_8963);
nor U9913 (N_9913,N_8634,N_8883);
nand U9914 (N_9914,N_8135,N_8599);
or U9915 (N_9915,N_8549,N_8230);
xor U9916 (N_9916,N_8735,N_8458);
and U9917 (N_9917,N_8754,N_8929);
or U9918 (N_9918,N_8881,N_8121);
nor U9919 (N_9919,N_8683,N_8636);
and U9920 (N_9920,N_8705,N_8629);
and U9921 (N_9921,N_8932,N_8793);
xnor U9922 (N_9922,N_8696,N_8092);
xnor U9923 (N_9923,N_8144,N_8209);
xnor U9924 (N_9924,N_8793,N_8388);
nor U9925 (N_9925,N_8441,N_8163);
xor U9926 (N_9926,N_8272,N_8712);
xnor U9927 (N_9927,N_8429,N_8422);
nor U9928 (N_9928,N_8807,N_8836);
and U9929 (N_9929,N_8552,N_8075);
or U9930 (N_9930,N_8700,N_8478);
nand U9931 (N_9931,N_8839,N_8560);
nor U9932 (N_9932,N_8755,N_8907);
xor U9933 (N_9933,N_8886,N_8008);
or U9934 (N_9934,N_8825,N_8353);
or U9935 (N_9935,N_8192,N_8114);
nand U9936 (N_9936,N_8651,N_8620);
xor U9937 (N_9937,N_8941,N_8486);
xor U9938 (N_9938,N_8666,N_8850);
nand U9939 (N_9939,N_8379,N_8037);
nand U9940 (N_9940,N_8849,N_8242);
nor U9941 (N_9941,N_8712,N_8576);
or U9942 (N_9942,N_8355,N_8053);
or U9943 (N_9943,N_8848,N_8113);
nand U9944 (N_9944,N_8486,N_8007);
or U9945 (N_9945,N_8920,N_8495);
xnor U9946 (N_9946,N_8171,N_8892);
xnor U9947 (N_9947,N_8984,N_8751);
xor U9948 (N_9948,N_8351,N_8978);
and U9949 (N_9949,N_8920,N_8157);
and U9950 (N_9950,N_8093,N_8895);
xor U9951 (N_9951,N_8469,N_8298);
nand U9952 (N_9952,N_8653,N_8532);
or U9953 (N_9953,N_8324,N_8819);
or U9954 (N_9954,N_8816,N_8115);
xnor U9955 (N_9955,N_8950,N_8914);
nor U9956 (N_9956,N_8103,N_8630);
or U9957 (N_9957,N_8807,N_8203);
nand U9958 (N_9958,N_8405,N_8162);
nor U9959 (N_9959,N_8592,N_8479);
nand U9960 (N_9960,N_8660,N_8630);
nor U9961 (N_9961,N_8874,N_8442);
xor U9962 (N_9962,N_8276,N_8332);
xor U9963 (N_9963,N_8663,N_8736);
nor U9964 (N_9964,N_8227,N_8743);
and U9965 (N_9965,N_8449,N_8394);
xor U9966 (N_9966,N_8095,N_8866);
or U9967 (N_9967,N_8013,N_8209);
nand U9968 (N_9968,N_8034,N_8057);
nand U9969 (N_9969,N_8210,N_8951);
or U9970 (N_9970,N_8215,N_8207);
nand U9971 (N_9971,N_8791,N_8609);
xor U9972 (N_9972,N_8858,N_8618);
nor U9973 (N_9973,N_8344,N_8214);
xor U9974 (N_9974,N_8896,N_8291);
xnor U9975 (N_9975,N_8490,N_8808);
and U9976 (N_9976,N_8312,N_8528);
or U9977 (N_9977,N_8004,N_8834);
xor U9978 (N_9978,N_8357,N_8280);
or U9979 (N_9979,N_8690,N_8060);
and U9980 (N_9980,N_8434,N_8777);
nand U9981 (N_9981,N_8370,N_8867);
xor U9982 (N_9982,N_8063,N_8431);
nor U9983 (N_9983,N_8204,N_8517);
or U9984 (N_9984,N_8752,N_8316);
and U9985 (N_9985,N_8964,N_8837);
xnor U9986 (N_9986,N_8119,N_8588);
nor U9987 (N_9987,N_8500,N_8269);
xnor U9988 (N_9988,N_8408,N_8521);
and U9989 (N_9989,N_8829,N_8349);
xor U9990 (N_9990,N_8407,N_8600);
and U9991 (N_9991,N_8673,N_8314);
or U9992 (N_9992,N_8620,N_8639);
or U9993 (N_9993,N_8091,N_8341);
nor U9994 (N_9994,N_8284,N_8815);
xor U9995 (N_9995,N_8319,N_8322);
and U9996 (N_9996,N_8745,N_8510);
or U9997 (N_9997,N_8067,N_8686);
or U9998 (N_9998,N_8507,N_8502);
and U9999 (N_9999,N_8217,N_8938);
and U10000 (N_10000,N_9292,N_9805);
or U10001 (N_10001,N_9372,N_9670);
or U10002 (N_10002,N_9435,N_9912);
nand U10003 (N_10003,N_9310,N_9527);
nand U10004 (N_10004,N_9413,N_9125);
nor U10005 (N_10005,N_9215,N_9083);
or U10006 (N_10006,N_9356,N_9890);
nor U10007 (N_10007,N_9687,N_9332);
nand U10008 (N_10008,N_9661,N_9023);
xnor U10009 (N_10009,N_9090,N_9876);
and U10010 (N_10010,N_9505,N_9592);
and U10011 (N_10011,N_9093,N_9766);
or U10012 (N_10012,N_9722,N_9241);
nor U10013 (N_10013,N_9422,N_9938);
xor U10014 (N_10014,N_9149,N_9638);
and U10015 (N_10015,N_9644,N_9052);
nor U10016 (N_10016,N_9784,N_9642);
nor U10017 (N_10017,N_9965,N_9764);
and U10018 (N_10018,N_9289,N_9309);
and U10019 (N_10019,N_9221,N_9866);
nor U10020 (N_10020,N_9769,N_9913);
and U10021 (N_10021,N_9955,N_9130);
and U10022 (N_10022,N_9377,N_9516);
nand U10023 (N_10023,N_9059,N_9346);
and U10024 (N_10024,N_9544,N_9240);
xor U10025 (N_10025,N_9019,N_9629);
and U10026 (N_10026,N_9392,N_9852);
nor U10027 (N_10027,N_9131,N_9094);
xnor U10028 (N_10028,N_9345,N_9326);
nand U10029 (N_10029,N_9024,N_9791);
and U10030 (N_10030,N_9248,N_9760);
or U10031 (N_10031,N_9018,N_9998);
nor U10032 (N_10032,N_9983,N_9757);
nand U10033 (N_10033,N_9821,N_9899);
and U10034 (N_10034,N_9300,N_9777);
xor U10035 (N_10035,N_9584,N_9370);
or U10036 (N_10036,N_9956,N_9279);
nor U10037 (N_10037,N_9324,N_9573);
xor U10038 (N_10038,N_9686,N_9773);
xor U10039 (N_10039,N_9949,N_9972);
xnor U10040 (N_10040,N_9917,N_9306);
nand U10041 (N_10041,N_9713,N_9541);
xnor U10042 (N_10042,N_9271,N_9257);
and U10043 (N_10043,N_9099,N_9837);
or U10044 (N_10044,N_9462,N_9360);
and U10045 (N_10045,N_9880,N_9648);
xnor U10046 (N_10046,N_9609,N_9311);
and U10047 (N_10047,N_9296,N_9261);
nand U10048 (N_10048,N_9961,N_9349);
nand U10049 (N_10049,N_9655,N_9603);
nand U10050 (N_10050,N_9555,N_9733);
nand U10051 (N_10051,N_9028,N_9148);
and U10052 (N_10052,N_9634,N_9513);
and U10053 (N_10053,N_9350,N_9438);
and U10054 (N_10054,N_9230,N_9994);
nand U10055 (N_10055,N_9159,N_9104);
nand U10056 (N_10056,N_9814,N_9385);
xnor U10057 (N_10057,N_9539,N_9204);
nor U10058 (N_10058,N_9782,N_9278);
xnor U10059 (N_10059,N_9667,N_9185);
or U10060 (N_10060,N_9981,N_9651);
or U10061 (N_10061,N_9613,N_9500);
nor U10062 (N_10062,N_9726,N_9160);
and U10063 (N_10063,N_9080,N_9245);
nor U10064 (N_10064,N_9266,N_9973);
or U10065 (N_10065,N_9016,N_9220);
xor U10066 (N_10066,N_9277,N_9953);
nand U10067 (N_10067,N_9902,N_9748);
or U10068 (N_10068,N_9276,N_9809);
and U10069 (N_10069,N_9563,N_9728);
nor U10070 (N_10070,N_9354,N_9301);
nand U10071 (N_10071,N_9931,N_9719);
or U10072 (N_10072,N_9041,N_9247);
xor U10073 (N_10073,N_9308,N_9113);
nor U10074 (N_10074,N_9872,N_9258);
xor U10075 (N_10075,N_9906,N_9910);
xnor U10076 (N_10076,N_9151,N_9492);
and U10077 (N_10077,N_9526,N_9206);
nand U10078 (N_10078,N_9101,N_9810);
and U10079 (N_10079,N_9829,N_9293);
nor U10080 (N_10080,N_9022,N_9677);
nand U10081 (N_10081,N_9854,N_9272);
nor U10082 (N_10082,N_9891,N_9237);
nand U10083 (N_10083,N_9923,N_9589);
xnor U10084 (N_10084,N_9624,N_9193);
nand U10085 (N_10085,N_9768,N_9534);
nor U10086 (N_10086,N_9055,N_9205);
nor U10087 (N_10087,N_9280,N_9542);
nand U10088 (N_10088,N_9176,N_9834);
nor U10089 (N_10089,N_9739,N_9254);
xor U10090 (N_10090,N_9063,N_9868);
nor U10091 (N_10091,N_9408,N_9781);
nor U10092 (N_10092,N_9611,N_9825);
nor U10093 (N_10093,N_9456,N_9997);
xnor U10094 (N_10094,N_9968,N_9143);
nor U10095 (N_10095,N_9776,N_9366);
nand U10096 (N_10096,N_9340,N_9894);
nor U10097 (N_10097,N_9479,N_9331);
xor U10098 (N_10098,N_9136,N_9317);
and U10099 (N_10099,N_9683,N_9610);
xnor U10100 (N_10100,N_9971,N_9323);
xor U10101 (N_10101,N_9086,N_9951);
nor U10102 (N_10102,N_9081,N_9915);
nand U10103 (N_10103,N_9993,N_9069);
xor U10104 (N_10104,N_9368,N_9364);
xnor U10105 (N_10105,N_9696,N_9316);
and U10106 (N_10106,N_9407,N_9515);
nor U10107 (N_10107,N_9133,N_9657);
xnor U10108 (N_10108,N_9823,N_9598);
nand U10109 (N_10109,N_9144,N_9811);
nor U10110 (N_10110,N_9464,N_9622);
xor U10111 (N_10111,N_9625,N_9399);
nor U10112 (N_10112,N_9882,N_9509);
nor U10113 (N_10113,N_9989,N_9889);
and U10114 (N_10114,N_9905,N_9991);
xor U10115 (N_10115,N_9156,N_9379);
and U10116 (N_10116,N_9750,N_9295);
or U10117 (N_10117,N_9494,N_9886);
nor U10118 (N_10118,N_9153,N_9618);
nor U10119 (N_10119,N_9561,N_9680);
xnor U10120 (N_10120,N_9134,N_9431);
and U10121 (N_10121,N_9627,N_9383);
nand U10122 (N_10122,N_9608,N_9294);
or U10123 (N_10123,N_9192,N_9304);
nand U10124 (N_10124,N_9984,N_9146);
and U10125 (N_10125,N_9362,N_9694);
nand U10126 (N_10126,N_9535,N_9470);
nor U10127 (N_10127,N_9703,N_9646);
or U10128 (N_10128,N_9112,N_9877);
nor U10129 (N_10129,N_9954,N_9730);
and U10130 (N_10130,N_9478,N_9168);
xnor U10131 (N_10131,N_9663,N_9074);
nand U10132 (N_10132,N_9723,N_9214);
nor U10133 (N_10133,N_9329,N_9297);
nand U10134 (N_10134,N_9046,N_9283);
nand U10135 (N_10135,N_9284,N_9091);
or U10136 (N_10136,N_9166,N_9458);
nand U10137 (N_10137,N_9386,N_9529);
nand U10138 (N_10138,N_9108,N_9344);
nand U10139 (N_10139,N_9171,N_9441);
and U10140 (N_10140,N_9562,N_9615);
xor U10141 (N_10141,N_9126,N_9471);
nand U10142 (N_10142,N_9732,N_9058);
nand U10143 (N_10143,N_9884,N_9161);
xnor U10144 (N_10144,N_9957,N_9740);
and U10145 (N_10145,N_9314,N_9384);
or U10146 (N_10146,N_9477,N_9574);
nor U10147 (N_10147,N_9941,N_9273);
nand U10148 (N_10148,N_9845,N_9832);
nand U10149 (N_10149,N_9184,N_9469);
nor U10150 (N_10150,N_9073,N_9461);
or U10151 (N_10151,N_9619,N_9715);
nand U10152 (N_10152,N_9096,N_9869);
nand U10153 (N_10153,N_9140,N_9669);
nand U10154 (N_10154,N_9786,N_9565);
xor U10155 (N_10155,N_9787,N_9229);
nor U10156 (N_10156,N_9506,N_9616);
nand U10157 (N_10157,N_9194,N_9933);
and U10158 (N_10158,N_9556,N_9975);
nor U10159 (N_10159,N_9859,N_9499);
and U10160 (N_10160,N_9958,N_9075);
nor U10161 (N_10161,N_9010,N_9577);
and U10162 (N_10162,N_9327,N_9780);
and U10163 (N_10163,N_9879,N_9996);
and U10164 (N_10164,N_9762,N_9508);
nand U10165 (N_10165,N_9631,N_9633);
and U10166 (N_10166,N_9927,N_9078);
and U10167 (N_10167,N_9200,N_9313);
or U10168 (N_10168,N_9801,N_9636);
nor U10169 (N_10169,N_9793,N_9488);
and U10170 (N_10170,N_9475,N_9390);
xor U10171 (N_10171,N_9495,N_9480);
and U10172 (N_10172,N_9034,N_9579);
or U10173 (N_10173,N_9639,N_9107);
nor U10174 (N_10174,N_9436,N_9575);
and U10175 (N_10175,N_9216,N_9770);
nand U10176 (N_10176,N_9348,N_9967);
nand U10177 (N_10177,N_9207,N_9745);
nor U10178 (N_10178,N_9549,N_9881);
or U10179 (N_10179,N_9738,N_9448);
nor U10180 (N_10180,N_9921,N_9578);
nor U10181 (N_10181,N_9371,N_9959);
and U10182 (N_10182,N_9459,N_9596);
xor U10183 (N_10183,N_9536,N_9567);
or U10184 (N_10184,N_9571,N_9342);
and U10185 (N_10185,N_9928,N_9822);
nor U10186 (N_10186,N_9789,N_9040);
or U10187 (N_10187,N_9922,N_9424);
and U10188 (N_10188,N_9946,N_9901);
nand U10189 (N_10189,N_9520,N_9446);
nand U10190 (N_10190,N_9824,N_9674);
xor U10191 (N_10191,N_9219,N_9602);
and U10192 (N_10192,N_9060,N_9201);
and U10193 (N_10193,N_9485,N_9502);
xnor U10194 (N_10194,N_9916,N_9400);
nand U10195 (N_10195,N_9919,N_9813);
xnor U10196 (N_10196,N_9759,N_9256);
nor U10197 (N_10197,N_9275,N_9152);
nand U10198 (N_10198,N_9614,N_9650);
xnor U10199 (N_10199,N_9576,N_9640);
xor U10200 (N_10200,N_9878,N_9393);
and U10201 (N_10201,N_9550,N_9758);
xor U10202 (N_10202,N_9196,N_9365);
nor U10203 (N_10203,N_9451,N_9678);
nand U10204 (N_10204,N_9681,N_9818);
xor U10205 (N_10205,N_9162,N_9027);
nor U10206 (N_10206,N_9566,N_9718);
or U10207 (N_10207,N_9597,N_9654);
and U10208 (N_10208,N_9483,N_9026);
or U10209 (N_10209,N_9966,N_9425);
and U10210 (N_10210,N_9778,N_9582);
xor U10211 (N_10211,N_9009,N_9269);
nand U10212 (N_10212,N_9706,N_9198);
xor U10213 (N_10213,N_9173,N_9065);
nor U10214 (N_10214,N_9716,N_9858);
nor U10215 (N_10215,N_9714,N_9432);
or U10216 (N_10216,N_9208,N_9755);
and U10217 (N_10217,N_9203,N_9337);
xnor U10218 (N_10218,N_9511,N_9320);
or U10219 (N_10219,N_9406,N_9830);
and U10220 (N_10220,N_9637,N_9044);
nand U10221 (N_10221,N_9465,N_9066);
and U10222 (N_10222,N_9684,N_9600);
xor U10223 (N_10223,N_9903,N_9045);
or U10224 (N_10224,N_9969,N_9803);
nand U10225 (N_10225,N_9021,N_9986);
nand U10226 (N_10226,N_9850,N_9274);
or U10227 (N_10227,N_9088,N_9007);
xor U10228 (N_10228,N_9222,N_9501);
nor U10229 (N_10229,N_9068,N_9202);
or U10230 (N_10230,N_9569,N_9754);
or U10231 (N_10231,N_9976,N_9265);
xor U10232 (N_10232,N_9417,N_9098);
nor U10233 (N_10233,N_9699,N_9286);
nand U10234 (N_10234,N_9774,N_9530);
nor U10235 (N_10235,N_9802,N_9403);
and U10236 (N_10236,N_9033,N_9887);
nand U10237 (N_10237,N_9111,N_9163);
xor U10238 (N_10238,N_9712,N_9930);
xor U10239 (N_10239,N_9893,N_9623);
and U10240 (N_10240,N_9717,N_9382);
and U10241 (N_10241,N_9226,N_9253);
and U10242 (N_10242,N_9792,N_9860);
xnor U10243 (N_10243,N_9689,N_9076);
xor U10244 (N_10244,N_9302,N_9808);
xnor U10245 (N_10245,N_9118,N_9775);
xnor U10246 (N_10246,N_9645,N_9123);
xnor U10247 (N_10247,N_9333,N_9165);
xor U10248 (N_10248,N_9135,N_9334);
xor U10249 (N_10249,N_9486,N_9217);
or U10250 (N_10250,N_9260,N_9794);
or U10251 (N_10251,N_9238,N_9389);
or U10252 (N_10252,N_9085,N_9433);
nand U10253 (N_10253,N_9591,N_9559);
nand U10254 (N_10254,N_9831,N_9347);
and U10255 (N_10255,N_9940,N_9155);
nor U10256 (N_10256,N_9585,N_9799);
or U10257 (N_10257,N_9401,N_9896);
xnor U10258 (N_10258,N_9932,N_9514);
and U10259 (N_10259,N_9992,N_9262);
nand U10260 (N_10260,N_9067,N_9231);
xor U10261 (N_10261,N_9593,N_9416);
nand U10262 (N_10262,N_9412,N_9978);
nor U10263 (N_10263,N_9013,N_9572);
nor U10264 (N_10264,N_9030,N_9374);
nand U10265 (N_10265,N_9054,N_9990);
and U10266 (N_10266,N_9988,N_9632);
or U10267 (N_10267,N_9628,N_9867);
nand U10268 (N_10268,N_9798,N_9761);
nand U10269 (N_10269,N_9741,N_9711);
and U10270 (N_10270,N_9756,N_9698);
or U10271 (N_10271,N_9132,N_9409);
xor U10272 (N_10272,N_9251,N_9195);
xnor U10273 (N_10273,N_9476,N_9395);
nand U10274 (N_10274,N_9147,N_9797);
xor U10275 (N_10275,N_9191,N_9396);
and U10276 (N_10276,N_9736,N_9355);
nor U10277 (N_10277,N_9128,N_9418);
nand U10278 (N_10278,N_9381,N_9002);
and U10279 (N_10279,N_9167,N_9865);
and U10280 (N_10280,N_9692,N_9102);
nand U10281 (N_10281,N_9904,N_9169);
nand U10282 (N_10282,N_9322,N_9907);
or U10283 (N_10283,N_9707,N_9870);
xnor U10284 (N_10284,N_9325,N_9528);
nor U10285 (N_10285,N_9227,N_9188);
and U10286 (N_10286,N_9507,N_9255);
xnor U10287 (N_10287,N_9186,N_9339);
nand U10288 (N_10288,N_9020,N_9551);
nand U10289 (N_10289,N_9950,N_9537);
and U10290 (N_10290,N_9553,N_9116);
xnor U10291 (N_10291,N_9763,N_9082);
nor U10292 (N_10292,N_9744,N_9664);
or U10293 (N_10293,N_9474,N_9735);
and U10294 (N_10294,N_9795,N_9343);
and U10295 (N_10295,N_9659,N_9137);
and U10296 (N_10296,N_9359,N_9017);
and U10297 (N_10297,N_9570,N_9452);
nand U10298 (N_10298,N_9328,N_9557);
xnor U10299 (N_10299,N_9532,N_9228);
xnor U10300 (N_10300,N_9855,N_9982);
nand U10301 (N_10301,N_9110,N_9234);
or U10302 (N_10302,N_9242,N_9223);
nor U10303 (N_10303,N_9607,N_9545);
and U10304 (N_10304,N_9935,N_9897);
xor U10305 (N_10305,N_9807,N_9012);
and U10306 (N_10306,N_9232,N_9145);
xnor U10307 (N_10307,N_9341,N_9072);
xor U10308 (N_10308,N_9236,N_9211);
xnor U10309 (N_10309,N_9693,N_9742);
xor U10310 (N_10310,N_9658,N_9164);
nand U10311 (N_10311,N_9487,N_9482);
or U10312 (N_10312,N_9106,N_9977);
nor U10313 (N_10313,N_9943,N_9839);
or U10314 (N_10314,N_9697,N_9178);
nand U10315 (N_10315,N_9036,N_9496);
and U10316 (N_10316,N_9043,N_9743);
and U10317 (N_10317,N_9042,N_9468);
and U10318 (N_10318,N_9109,N_9129);
and U10319 (N_10319,N_9049,N_9691);
nand U10320 (N_10320,N_9213,N_9397);
nor U10321 (N_10321,N_9523,N_9533);
nor U10322 (N_10322,N_9734,N_9626);
xnor U10323 (N_10323,N_9838,N_9911);
or U10324 (N_10324,N_9490,N_9358);
nand U10325 (N_10325,N_9233,N_9857);
or U10326 (N_10326,N_9444,N_9856);
nor U10327 (N_10327,N_9369,N_9114);
and U10328 (N_10328,N_9209,N_9252);
nor U10329 (N_10329,N_9586,N_9804);
nor U10330 (N_10330,N_9538,N_9620);
nand U10331 (N_10331,N_9548,N_9048);
nor U10332 (N_10332,N_9641,N_9330);
nand U10333 (N_10333,N_9427,N_9727);
nand U10334 (N_10334,N_9970,N_9440);
nor U10335 (N_10335,N_9851,N_9580);
xnor U10336 (N_10336,N_9449,N_9197);
xnor U10337 (N_10337,N_9785,N_9394);
nor U10338 (N_10338,N_9095,N_9092);
nand U10339 (N_10339,N_9939,N_9335);
nor U10340 (N_10340,N_9051,N_9087);
and U10341 (N_10341,N_9695,N_9429);
nand U10342 (N_10342,N_9029,N_9053);
xor U10343 (N_10343,N_9244,N_9652);
or U10344 (N_10344,N_9914,N_9702);
nor U10345 (N_10345,N_9466,N_9885);
and U10346 (N_10346,N_9373,N_9601);
or U10347 (N_10347,N_9025,N_9840);
xor U10348 (N_10348,N_9863,N_9239);
or U10349 (N_10349,N_9675,N_9710);
or U10350 (N_10350,N_9120,N_9319);
xnor U10351 (N_10351,N_9455,N_9387);
nor U10352 (N_10352,N_9378,N_9250);
xor U10353 (N_10353,N_9588,N_9685);
nand U10354 (N_10354,N_9182,N_9015);
and U10355 (N_10355,N_9158,N_9900);
and U10356 (N_10356,N_9122,N_9790);
nor U10357 (N_10357,N_9463,N_9725);
nand U10358 (N_10358,N_9558,N_9150);
or U10359 (N_10359,N_9709,N_9415);
or U10360 (N_10360,N_9828,N_9127);
or U10361 (N_10361,N_9376,N_9874);
xnor U10362 (N_10362,N_9942,N_9351);
nor U10363 (N_10363,N_9835,N_9014);
nand U10364 (N_10364,N_9985,N_9924);
and U10365 (N_10365,N_9268,N_9679);
or U10366 (N_10366,N_9826,N_9353);
or U10367 (N_10367,N_9606,N_9518);
nand U10368 (N_10368,N_9497,N_9605);
nand U10369 (N_10369,N_9510,N_9414);
nand U10370 (N_10370,N_9945,N_9056);
nand U10371 (N_10371,N_9139,N_9751);
or U10372 (N_10372,N_9987,N_9000);
nor U10373 (N_10373,N_9307,N_9212);
and U10374 (N_10374,N_9656,N_9243);
xnor U10375 (N_10375,N_9061,N_9543);
and U10376 (N_10376,N_9445,N_9357);
xor U10377 (N_10377,N_9746,N_9047);
or U10378 (N_10378,N_9649,N_9181);
or U10379 (N_10379,N_9361,N_9453);
and U10380 (N_10380,N_9079,N_9428);
and U10381 (N_10381,N_9170,N_9175);
xor U10382 (N_10382,N_9174,N_9848);
nor U10383 (N_10383,N_9404,N_9682);
or U10384 (N_10384,N_9815,N_9898);
nand U10385 (N_10385,N_9419,N_9721);
nor U10386 (N_10386,N_9443,N_9594);
and U10387 (N_10387,N_9920,N_9673);
nor U10388 (N_10388,N_9752,N_9522);
xor U10389 (N_10389,N_9587,N_9581);
nor U10390 (N_10390,N_9617,N_9484);
or U10391 (N_10391,N_9908,N_9157);
and U10392 (N_10392,N_9398,N_9225);
nand U10393 (N_10393,N_9704,N_9299);
or U10394 (N_10394,N_9963,N_9367);
or U10395 (N_10395,N_9783,N_9929);
nor U10396 (N_10396,N_9454,N_9962);
nand U10397 (N_10397,N_9918,N_9590);
or U10398 (N_10398,N_9481,N_9560);
or U10399 (N_10399,N_9298,N_9621);
and U10400 (N_10400,N_9948,N_9105);
and U10401 (N_10401,N_9062,N_9352);
or U10402 (N_10402,N_9363,N_9011);
nor U10403 (N_10403,N_9430,N_9979);
or U10404 (N_10404,N_9312,N_9554);
and U10405 (N_10405,N_9547,N_9934);
xnor U10406 (N_10406,N_9517,N_9039);
and U10407 (N_10407,N_9071,N_9599);
nand U10408 (N_10408,N_9421,N_9552);
and U10409 (N_10409,N_9003,N_9117);
nor U10410 (N_10410,N_9779,N_9006);
xnor U10411 (N_10411,N_9729,N_9800);
and U10412 (N_10412,N_9224,N_9875);
and U10413 (N_10413,N_9100,N_9853);
xnor U10414 (N_10414,N_9883,N_9318);
or U10415 (N_10415,N_9862,N_9287);
xnor U10416 (N_10416,N_9391,N_9190);
nand U10417 (N_10417,N_9138,N_9546);
xor U10418 (N_10418,N_9564,N_9926);
or U10419 (N_10419,N_9812,N_9057);
xnor U10420 (N_10420,N_9701,N_9662);
or U10421 (N_10421,N_9861,N_9183);
nand U10422 (N_10422,N_9583,N_9647);
nand U10423 (N_10423,N_9630,N_9964);
or U10424 (N_10424,N_9844,N_9525);
and U10425 (N_10425,N_9816,N_9124);
nor U10426 (N_10426,N_9305,N_9064);
or U10427 (N_10427,N_9491,N_9411);
and U10428 (N_10428,N_9154,N_9442);
xnor U10429 (N_10429,N_9199,N_9771);
xor U10430 (N_10430,N_9489,N_9888);
or U10431 (N_10431,N_9303,N_9434);
or U10432 (N_10432,N_9842,N_9708);
nand U10433 (N_10433,N_9005,N_9388);
or U10434 (N_10434,N_9503,N_9871);
xnor U10435 (N_10435,N_9288,N_9032);
nor U10436 (N_10436,N_9338,N_9660);
nor U10437 (N_10437,N_9285,N_9653);
xor U10438 (N_10438,N_9688,N_9282);
and U10439 (N_10439,N_9568,N_9259);
and U10440 (N_10440,N_9604,N_9038);
nand U10441 (N_10441,N_9249,N_9439);
nor U10442 (N_10442,N_9405,N_9512);
and U10443 (N_10443,N_9974,N_9747);
or U10444 (N_10444,N_9089,N_9947);
nor U10445 (N_10445,N_9724,N_9291);
or U10446 (N_10446,N_9031,N_9402);
or U10447 (N_10447,N_9410,N_9450);
xnor U10448 (N_10448,N_9960,N_9270);
nand U10449 (N_10449,N_9864,N_9457);
nor U10450 (N_10450,N_9690,N_9849);
and U10451 (N_10451,N_9423,N_9460);
nor U10452 (N_10452,N_9037,N_9179);
nor U10453 (N_10453,N_9035,N_9172);
xnor U10454 (N_10454,N_9519,N_9473);
or U10455 (N_10455,N_9375,N_9720);
nand U10456 (N_10456,N_9936,N_9420);
xor U10457 (N_10457,N_9315,N_9290);
xor U10458 (N_10458,N_9892,N_9246);
nand U10459 (N_10459,N_9187,N_9498);
nor U10460 (N_10460,N_9737,N_9531);
nor U10461 (N_10461,N_9008,N_9944);
xnor U10462 (N_10462,N_9142,N_9671);
and U10463 (N_10463,N_9846,N_9426);
or U10464 (N_10464,N_9827,N_9873);
nor U10465 (N_10465,N_9666,N_9820);
nor U10466 (N_10466,N_9817,N_9141);
xor U10467 (N_10467,N_9767,N_9321);
xor U10468 (N_10468,N_9235,N_9788);
nand U10469 (N_10469,N_9833,N_9925);
and U10470 (N_10470,N_9281,N_9676);
nand U10471 (N_10471,N_9847,N_9180);
nor U10472 (N_10472,N_9731,N_9210);
nand U10473 (N_10473,N_9004,N_9467);
xor U10474 (N_10474,N_9665,N_9705);
or U10475 (N_10475,N_9119,N_9612);
xnor U10476 (N_10476,N_9263,N_9937);
nor U10477 (N_10477,N_9103,N_9668);
xor U10478 (N_10478,N_9264,N_9995);
or U10479 (N_10479,N_9001,N_9980);
or U10480 (N_10480,N_9218,N_9084);
nand U10481 (N_10481,N_9753,N_9189);
and U10482 (N_10482,N_9643,N_9097);
nor U10483 (N_10483,N_9540,N_9336);
xnor U10484 (N_10484,N_9909,N_9472);
nand U10485 (N_10485,N_9635,N_9595);
and U10486 (N_10486,N_9796,N_9437);
and U10487 (N_10487,N_9765,N_9952);
nand U10488 (N_10488,N_9115,N_9843);
nand U10489 (N_10489,N_9700,N_9672);
xnor U10490 (N_10490,N_9836,N_9524);
xor U10491 (N_10491,N_9447,N_9493);
nand U10492 (N_10492,N_9521,N_9895);
and U10493 (N_10493,N_9504,N_9177);
and U10494 (N_10494,N_9749,N_9070);
xnor U10495 (N_10495,N_9806,N_9077);
nand U10496 (N_10496,N_9267,N_9841);
xor U10497 (N_10497,N_9380,N_9999);
xnor U10498 (N_10498,N_9121,N_9050);
and U10499 (N_10499,N_9772,N_9819);
nand U10500 (N_10500,N_9361,N_9075);
xnor U10501 (N_10501,N_9691,N_9901);
xor U10502 (N_10502,N_9346,N_9756);
xnor U10503 (N_10503,N_9020,N_9479);
xnor U10504 (N_10504,N_9737,N_9418);
or U10505 (N_10505,N_9912,N_9415);
and U10506 (N_10506,N_9830,N_9018);
nor U10507 (N_10507,N_9754,N_9079);
xor U10508 (N_10508,N_9263,N_9385);
nor U10509 (N_10509,N_9206,N_9521);
nand U10510 (N_10510,N_9836,N_9164);
nand U10511 (N_10511,N_9092,N_9105);
nand U10512 (N_10512,N_9350,N_9038);
or U10513 (N_10513,N_9944,N_9796);
nand U10514 (N_10514,N_9120,N_9043);
nand U10515 (N_10515,N_9935,N_9853);
xnor U10516 (N_10516,N_9952,N_9844);
nor U10517 (N_10517,N_9454,N_9460);
nor U10518 (N_10518,N_9736,N_9619);
nor U10519 (N_10519,N_9129,N_9504);
xnor U10520 (N_10520,N_9978,N_9152);
nor U10521 (N_10521,N_9269,N_9951);
nor U10522 (N_10522,N_9277,N_9816);
nand U10523 (N_10523,N_9083,N_9928);
and U10524 (N_10524,N_9214,N_9711);
nand U10525 (N_10525,N_9989,N_9137);
nor U10526 (N_10526,N_9528,N_9039);
or U10527 (N_10527,N_9482,N_9483);
or U10528 (N_10528,N_9111,N_9846);
nor U10529 (N_10529,N_9640,N_9497);
nor U10530 (N_10530,N_9681,N_9823);
nor U10531 (N_10531,N_9047,N_9413);
xnor U10532 (N_10532,N_9750,N_9826);
nor U10533 (N_10533,N_9425,N_9062);
xor U10534 (N_10534,N_9737,N_9144);
and U10535 (N_10535,N_9428,N_9678);
nor U10536 (N_10536,N_9998,N_9946);
and U10537 (N_10537,N_9957,N_9173);
xor U10538 (N_10538,N_9854,N_9683);
xnor U10539 (N_10539,N_9508,N_9161);
nand U10540 (N_10540,N_9334,N_9221);
nand U10541 (N_10541,N_9024,N_9318);
xnor U10542 (N_10542,N_9131,N_9085);
nand U10543 (N_10543,N_9024,N_9260);
or U10544 (N_10544,N_9492,N_9526);
nor U10545 (N_10545,N_9886,N_9617);
nand U10546 (N_10546,N_9655,N_9509);
nor U10547 (N_10547,N_9274,N_9444);
nand U10548 (N_10548,N_9325,N_9581);
xnor U10549 (N_10549,N_9388,N_9141);
nor U10550 (N_10550,N_9762,N_9163);
nand U10551 (N_10551,N_9351,N_9771);
nand U10552 (N_10552,N_9386,N_9842);
or U10553 (N_10553,N_9308,N_9427);
xnor U10554 (N_10554,N_9167,N_9797);
nand U10555 (N_10555,N_9224,N_9677);
xnor U10556 (N_10556,N_9273,N_9973);
xor U10557 (N_10557,N_9384,N_9986);
nand U10558 (N_10558,N_9962,N_9988);
nor U10559 (N_10559,N_9132,N_9046);
nand U10560 (N_10560,N_9918,N_9280);
xor U10561 (N_10561,N_9632,N_9195);
and U10562 (N_10562,N_9148,N_9222);
nand U10563 (N_10563,N_9600,N_9441);
and U10564 (N_10564,N_9201,N_9356);
xnor U10565 (N_10565,N_9281,N_9430);
and U10566 (N_10566,N_9427,N_9721);
or U10567 (N_10567,N_9044,N_9885);
nand U10568 (N_10568,N_9510,N_9185);
nor U10569 (N_10569,N_9863,N_9385);
nor U10570 (N_10570,N_9336,N_9387);
nand U10571 (N_10571,N_9162,N_9691);
or U10572 (N_10572,N_9615,N_9876);
xnor U10573 (N_10573,N_9358,N_9467);
nand U10574 (N_10574,N_9546,N_9135);
and U10575 (N_10575,N_9308,N_9702);
nand U10576 (N_10576,N_9784,N_9148);
nor U10577 (N_10577,N_9510,N_9378);
nand U10578 (N_10578,N_9247,N_9691);
and U10579 (N_10579,N_9132,N_9752);
nand U10580 (N_10580,N_9888,N_9671);
and U10581 (N_10581,N_9429,N_9843);
or U10582 (N_10582,N_9871,N_9372);
and U10583 (N_10583,N_9802,N_9317);
nand U10584 (N_10584,N_9017,N_9678);
or U10585 (N_10585,N_9055,N_9248);
nand U10586 (N_10586,N_9827,N_9322);
or U10587 (N_10587,N_9580,N_9098);
nand U10588 (N_10588,N_9389,N_9646);
nand U10589 (N_10589,N_9242,N_9628);
xnor U10590 (N_10590,N_9377,N_9652);
nor U10591 (N_10591,N_9344,N_9346);
or U10592 (N_10592,N_9908,N_9837);
nand U10593 (N_10593,N_9028,N_9597);
nand U10594 (N_10594,N_9315,N_9964);
nor U10595 (N_10595,N_9331,N_9646);
and U10596 (N_10596,N_9334,N_9977);
or U10597 (N_10597,N_9573,N_9068);
nor U10598 (N_10598,N_9367,N_9368);
xnor U10599 (N_10599,N_9242,N_9033);
and U10600 (N_10600,N_9739,N_9751);
xor U10601 (N_10601,N_9735,N_9649);
nor U10602 (N_10602,N_9786,N_9130);
and U10603 (N_10603,N_9990,N_9951);
and U10604 (N_10604,N_9508,N_9849);
and U10605 (N_10605,N_9899,N_9953);
nand U10606 (N_10606,N_9118,N_9860);
nand U10607 (N_10607,N_9646,N_9364);
nand U10608 (N_10608,N_9797,N_9700);
or U10609 (N_10609,N_9859,N_9191);
nand U10610 (N_10610,N_9373,N_9592);
or U10611 (N_10611,N_9202,N_9560);
nand U10612 (N_10612,N_9115,N_9836);
nand U10613 (N_10613,N_9614,N_9906);
and U10614 (N_10614,N_9945,N_9389);
nand U10615 (N_10615,N_9849,N_9166);
nand U10616 (N_10616,N_9191,N_9376);
and U10617 (N_10617,N_9835,N_9643);
xnor U10618 (N_10618,N_9415,N_9042);
and U10619 (N_10619,N_9077,N_9023);
nand U10620 (N_10620,N_9007,N_9172);
and U10621 (N_10621,N_9092,N_9913);
or U10622 (N_10622,N_9240,N_9691);
and U10623 (N_10623,N_9611,N_9163);
or U10624 (N_10624,N_9712,N_9595);
nor U10625 (N_10625,N_9890,N_9008);
and U10626 (N_10626,N_9514,N_9854);
nand U10627 (N_10627,N_9127,N_9323);
and U10628 (N_10628,N_9309,N_9780);
nand U10629 (N_10629,N_9815,N_9190);
or U10630 (N_10630,N_9154,N_9199);
and U10631 (N_10631,N_9146,N_9321);
nor U10632 (N_10632,N_9127,N_9369);
and U10633 (N_10633,N_9335,N_9544);
or U10634 (N_10634,N_9023,N_9601);
nand U10635 (N_10635,N_9468,N_9137);
nand U10636 (N_10636,N_9711,N_9750);
or U10637 (N_10637,N_9611,N_9455);
nand U10638 (N_10638,N_9624,N_9417);
or U10639 (N_10639,N_9161,N_9904);
and U10640 (N_10640,N_9791,N_9224);
and U10641 (N_10641,N_9110,N_9790);
xnor U10642 (N_10642,N_9205,N_9779);
nor U10643 (N_10643,N_9218,N_9669);
and U10644 (N_10644,N_9787,N_9725);
nor U10645 (N_10645,N_9083,N_9626);
and U10646 (N_10646,N_9294,N_9121);
or U10647 (N_10647,N_9665,N_9957);
nand U10648 (N_10648,N_9244,N_9886);
nor U10649 (N_10649,N_9849,N_9899);
nand U10650 (N_10650,N_9644,N_9392);
xor U10651 (N_10651,N_9446,N_9140);
or U10652 (N_10652,N_9135,N_9999);
xnor U10653 (N_10653,N_9614,N_9170);
and U10654 (N_10654,N_9177,N_9941);
nand U10655 (N_10655,N_9483,N_9522);
xnor U10656 (N_10656,N_9243,N_9556);
nor U10657 (N_10657,N_9267,N_9865);
or U10658 (N_10658,N_9038,N_9055);
nor U10659 (N_10659,N_9389,N_9186);
or U10660 (N_10660,N_9225,N_9785);
or U10661 (N_10661,N_9797,N_9517);
nand U10662 (N_10662,N_9516,N_9992);
xor U10663 (N_10663,N_9395,N_9874);
or U10664 (N_10664,N_9215,N_9225);
nand U10665 (N_10665,N_9258,N_9085);
xnor U10666 (N_10666,N_9784,N_9949);
or U10667 (N_10667,N_9561,N_9697);
xnor U10668 (N_10668,N_9790,N_9385);
nand U10669 (N_10669,N_9209,N_9134);
xor U10670 (N_10670,N_9766,N_9900);
and U10671 (N_10671,N_9233,N_9769);
or U10672 (N_10672,N_9598,N_9480);
or U10673 (N_10673,N_9563,N_9966);
or U10674 (N_10674,N_9480,N_9748);
nor U10675 (N_10675,N_9835,N_9445);
nor U10676 (N_10676,N_9671,N_9622);
nor U10677 (N_10677,N_9068,N_9194);
and U10678 (N_10678,N_9954,N_9531);
and U10679 (N_10679,N_9782,N_9703);
xor U10680 (N_10680,N_9234,N_9992);
nor U10681 (N_10681,N_9385,N_9499);
xnor U10682 (N_10682,N_9974,N_9885);
xnor U10683 (N_10683,N_9005,N_9369);
and U10684 (N_10684,N_9472,N_9301);
xnor U10685 (N_10685,N_9425,N_9600);
and U10686 (N_10686,N_9951,N_9642);
nor U10687 (N_10687,N_9823,N_9756);
nor U10688 (N_10688,N_9972,N_9654);
or U10689 (N_10689,N_9963,N_9354);
nand U10690 (N_10690,N_9599,N_9250);
or U10691 (N_10691,N_9218,N_9974);
xnor U10692 (N_10692,N_9783,N_9994);
or U10693 (N_10693,N_9969,N_9334);
and U10694 (N_10694,N_9338,N_9494);
nand U10695 (N_10695,N_9138,N_9587);
and U10696 (N_10696,N_9920,N_9947);
xor U10697 (N_10697,N_9939,N_9114);
and U10698 (N_10698,N_9570,N_9306);
nand U10699 (N_10699,N_9598,N_9806);
or U10700 (N_10700,N_9381,N_9218);
or U10701 (N_10701,N_9346,N_9115);
xnor U10702 (N_10702,N_9633,N_9923);
nand U10703 (N_10703,N_9280,N_9773);
xor U10704 (N_10704,N_9952,N_9337);
nand U10705 (N_10705,N_9504,N_9918);
or U10706 (N_10706,N_9544,N_9864);
or U10707 (N_10707,N_9856,N_9370);
xor U10708 (N_10708,N_9321,N_9317);
nand U10709 (N_10709,N_9418,N_9202);
xnor U10710 (N_10710,N_9656,N_9961);
and U10711 (N_10711,N_9922,N_9801);
xnor U10712 (N_10712,N_9962,N_9205);
nor U10713 (N_10713,N_9418,N_9855);
xnor U10714 (N_10714,N_9135,N_9159);
nand U10715 (N_10715,N_9699,N_9860);
and U10716 (N_10716,N_9381,N_9528);
xor U10717 (N_10717,N_9708,N_9671);
nand U10718 (N_10718,N_9811,N_9084);
nand U10719 (N_10719,N_9534,N_9252);
nor U10720 (N_10720,N_9326,N_9359);
xor U10721 (N_10721,N_9726,N_9913);
nor U10722 (N_10722,N_9361,N_9182);
xor U10723 (N_10723,N_9430,N_9121);
nand U10724 (N_10724,N_9496,N_9122);
nand U10725 (N_10725,N_9150,N_9802);
nor U10726 (N_10726,N_9328,N_9389);
nand U10727 (N_10727,N_9657,N_9194);
or U10728 (N_10728,N_9841,N_9062);
xnor U10729 (N_10729,N_9742,N_9306);
and U10730 (N_10730,N_9939,N_9916);
xor U10731 (N_10731,N_9227,N_9775);
and U10732 (N_10732,N_9390,N_9228);
xnor U10733 (N_10733,N_9366,N_9234);
xnor U10734 (N_10734,N_9396,N_9959);
nand U10735 (N_10735,N_9827,N_9895);
or U10736 (N_10736,N_9163,N_9085);
nand U10737 (N_10737,N_9978,N_9969);
or U10738 (N_10738,N_9245,N_9998);
nor U10739 (N_10739,N_9855,N_9511);
xor U10740 (N_10740,N_9766,N_9286);
nand U10741 (N_10741,N_9241,N_9308);
or U10742 (N_10742,N_9091,N_9117);
and U10743 (N_10743,N_9163,N_9195);
and U10744 (N_10744,N_9750,N_9268);
nand U10745 (N_10745,N_9944,N_9915);
xor U10746 (N_10746,N_9737,N_9983);
nor U10747 (N_10747,N_9693,N_9302);
nand U10748 (N_10748,N_9351,N_9021);
xnor U10749 (N_10749,N_9887,N_9137);
or U10750 (N_10750,N_9583,N_9609);
and U10751 (N_10751,N_9154,N_9603);
or U10752 (N_10752,N_9531,N_9253);
or U10753 (N_10753,N_9634,N_9615);
nor U10754 (N_10754,N_9432,N_9234);
nor U10755 (N_10755,N_9423,N_9554);
nor U10756 (N_10756,N_9451,N_9479);
xnor U10757 (N_10757,N_9001,N_9421);
or U10758 (N_10758,N_9774,N_9244);
and U10759 (N_10759,N_9546,N_9805);
xnor U10760 (N_10760,N_9195,N_9147);
and U10761 (N_10761,N_9699,N_9146);
xnor U10762 (N_10762,N_9690,N_9816);
or U10763 (N_10763,N_9983,N_9696);
nand U10764 (N_10764,N_9872,N_9038);
nand U10765 (N_10765,N_9323,N_9123);
nand U10766 (N_10766,N_9011,N_9054);
xnor U10767 (N_10767,N_9072,N_9854);
nand U10768 (N_10768,N_9622,N_9142);
nand U10769 (N_10769,N_9251,N_9316);
nor U10770 (N_10770,N_9484,N_9901);
nor U10771 (N_10771,N_9096,N_9130);
or U10772 (N_10772,N_9903,N_9731);
xnor U10773 (N_10773,N_9279,N_9903);
and U10774 (N_10774,N_9646,N_9091);
nand U10775 (N_10775,N_9302,N_9023);
nor U10776 (N_10776,N_9211,N_9391);
and U10777 (N_10777,N_9254,N_9632);
xnor U10778 (N_10778,N_9614,N_9889);
xor U10779 (N_10779,N_9830,N_9567);
or U10780 (N_10780,N_9497,N_9255);
nand U10781 (N_10781,N_9016,N_9168);
nor U10782 (N_10782,N_9793,N_9886);
or U10783 (N_10783,N_9303,N_9773);
nand U10784 (N_10784,N_9546,N_9308);
or U10785 (N_10785,N_9231,N_9880);
xor U10786 (N_10786,N_9567,N_9328);
or U10787 (N_10787,N_9846,N_9033);
nor U10788 (N_10788,N_9095,N_9536);
nand U10789 (N_10789,N_9724,N_9116);
xor U10790 (N_10790,N_9645,N_9367);
and U10791 (N_10791,N_9305,N_9002);
or U10792 (N_10792,N_9430,N_9404);
and U10793 (N_10793,N_9609,N_9691);
xor U10794 (N_10794,N_9536,N_9407);
nor U10795 (N_10795,N_9370,N_9412);
nand U10796 (N_10796,N_9345,N_9708);
nand U10797 (N_10797,N_9698,N_9138);
nand U10798 (N_10798,N_9563,N_9370);
nand U10799 (N_10799,N_9670,N_9025);
nor U10800 (N_10800,N_9808,N_9556);
nor U10801 (N_10801,N_9265,N_9786);
nand U10802 (N_10802,N_9109,N_9744);
nor U10803 (N_10803,N_9650,N_9082);
and U10804 (N_10804,N_9070,N_9527);
xnor U10805 (N_10805,N_9292,N_9831);
and U10806 (N_10806,N_9462,N_9309);
or U10807 (N_10807,N_9486,N_9615);
nand U10808 (N_10808,N_9459,N_9628);
nor U10809 (N_10809,N_9700,N_9903);
nand U10810 (N_10810,N_9721,N_9502);
nand U10811 (N_10811,N_9056,N_9978);
xor U10812 (N_10812,N_9222,N_9172);
or U10813 (N_10813,N_9644,N_9327);
or U10814 (N_10814,N_9406,N_9733);
nor U10815 (N_10815,N_9851,N_9457);
xnor U10816 (N_10816,N_9444,N_9097);
xor U10817 (N_10817,N_9935,N_9031);
xnor U10818 (N_10818,N_9688,N_9769);
nand U10819 (N_10819,N_9897,N_9318);
nand U10820 (N_10820,N_9000,N_9026);
nand U10821 (N_10821,N_9782,N_9025);
xnor U10822 (N_10822,N_9141,N_9208);
or U10823 (N_10823,N_9753,N_9871);
nor U10824 (N_10824,N_9002,N_9476);
nor U10825 (N_10825,N_9328,N_9867);
or U10826 (N_10826,N_9667,N_9700);
and U10827 (N_10827,N_9615,N_9169);
or U10828 (N_10828,N_9587,N_9285);
nor U10829 (N_10829,N_9416,N_9738);
or U10830 (N_10830,N_9621,N_9642);
and U10831 (N_10831,N_9016,N_9543);
or U10832 (N_10832,N_9819,N_9773);
xnor U10833 (N_10833,N_9584,N_9038);
nor U10834 (N_10834,N_9380,N_9298);
and U10835 (N_10835,N_9881,N_9571);
xnor U10836 (N_10836,N_9253,N_9782);
nor U10837 (N_10837,N_9963,N_9484);
and U10838 (N_10838,N_9143,N_9603);
nand U10839 (N_10839,N_9993,N_9700);
nand U10840 (N_10840,N_9153,N_9224);
nand U10841 (N_10841,N_9794,N_9153);
nand U10842 (N_10842,N_9460,N_9807);
nand U10843 (N_10843,N_9152,N_9660);
nor U10844 (N_10844,N_9651,N_9394);
or U10845 (N_10845,N_9896,N_9194);
or U10846 (N_10846,N_9417,N_9026);
and U10847 (N_10847,N_9552,N_9771);
xnor U10848 (N_10848,N_9667,N_9637);
xnor U10849 (N_10849,N_9740,N_9670);
nand U10850 (N_10850,N_9495,N_9149);
nor U10851 (N_10851,N_9747,N_9102);
nor U10852 (N_10852,N_9465,N_9076);
nand U10853 (N_10853,N_9389,N_9236);
nand U10854 (N_10854,N_9723,N_9478);
xnor U10855 (N_10855,N_9303,N_9013);
nor U10856 (N_10856,N_9356,N_9521);
nor U10857 (N_10857,N_9533,N_9230);
nand U10858 (N_10858,N_9502,N_9354);
nor U10859 (N_10859,N_9229,N_9752);
nand U10860 (N_10860,N_9777,N_9326);
or U10861 (N_10861,N_9379,N_9347);
and U10862 (N_10862,N_9890,N_9729);
nor U10863 (N_10863,N_9771,N_9349);
and U10864 (N_10864,N_9631,N_9046);
and U10865 (N_10865,N_9045,N_9007);
nand U10866 (N_10866,N_9940,N_9259);
nand U10867 (N_10867,N_9134,N_9585);
or U10868 (N_10868,N_9028,N_9421);
nand U10869 (N_10869,N_9707,N_9162);
nand U10870 (N_10870,N_9223,N_9826);
or U10871 (N_10871,N_9984,N_9325);
or U10872 (N_10872,N_9627,N_9208);
nand U10873 (N_10873,N_9677,N_9469);
or U10874 (N_10874,N_9849,N_9200);
nand U10875 (N_10875,N_9610,N_9532);
nor U10876 (N_10876,N_9360,N_9066);
nor U10877 (N_10877,N_9833,N_9514);
xnor U10878 (N_10878,N_9920,N_9519);
and U10879 (N_10879,N_9389,N_9230);
nor U10880 (N_10880,N_9558,N_9657);
xor U10881 (N_10881,N_9767,N_9901);
nor U10882 (N_10882,N_9514,N_9953);
and U10883 (N_10883,N_9454,N_9753);
xnor U10884 (N_10884,N_9254,N_9806);
xor U10885 (N_10885,N_9290,N_9670);
nor U10886 (N_10886,N_9465,N_9674);
nand U10887 (N_10887,N_9548,N_9539);
nand U10888 (N_10888,N_9058,N_9538);
nor U10889 (N_10889,N_9825,N_9331);
nor U10890 (N_10890,N_9631,N_9948);
or U10891 (N_10891,N_9322,N_9099);
nand U10892 (N_10892,N_9762,N_9487);
and U10893 (N_10893,N_9886,N_9772);
or U10894 (N_10894,N_9943,N_9741);
xnor U10895 (N_10895,N_9535,N_9258);
nor U10896 (N_10896,N_9839,N_9078);
nand U10897 (N_10897,N_9509,N_9454);
xor U10898 (N_10898,N_9749,N_9648);
and U10899 (N_10899,N_9657,N_9515);
or U10900 (N_10900,N_9221,N_9520);
xnor U10901 (N_10901,N_9235,N_9104);
and U10902 (N_10902,N_9741,N_9009);
and U10903 (N_10903,N_9687,N_9999);
nand U10904 (N_10904,N_9189,N_9584);
nand U10905 (N_10905,N_9836,N_9242);
or U10906 (N_10906,N_9767,N_9421);
or U10907 (N_10907,N_9298,N_9031);
or U10908 (N_10908,N_9738,N_9222);
xnor U10909 (N_10909,N_9214,N_9824);
xor U10910 (N_10910,N_9221,N_9997);
and U10911 (N_10911,N_9250,N_9135);
xnor U10912 (N_10912,N_9352,N_9872);
nor U10913 (N_10913,N_9160,N_9159);
xnor U10914 (N_10914,N_9209,N_9346);
nand U10915 (N_10915,N_9839,N_9320);
nor U10916 (N_10916,N_9044,N_9260);
xnor U10917 (N_10917,N_9510,N_9828);
nand U10918 (N_10918,N_9331,N_9934);
nor U10919 (N_10919,N_9994,N_9298);
nor U10920 (N_10920,N_9590,N_9741);
nand U10921 (N_10921,N_9477,N_9568);
and U10922 (N_10922,N_9024,N_9795);
xnor U10923 (N_10923,N_9502,N_9789);
nand U10924 (N_10924,N_9214,N_9922);
nor U10925 (N_10925,N_9429,N_9327);
xnor U10926 (N_10926,N_9289,N_9541);
and U10927 (N_10927,N_9014,N_9861);
and U10928 (N_10928,N_9309,N_9669);
or U10929 (N_10929,N_9171,N_9341);
nand U10930 (N_10930,N_9290,N_9456);
xor U10931 (N_10931,N_9126,N_9735);
nand U10932 (N_10932,N_9006,N_9894);
nor U10933 (N_10933,N_9573,N_9082);
xnor U10934 (N_10934,N_9129,N_9205);
nor U10935 (N_10935,N_9306,N_9831);
nand U10936 (N_10936,N_9220,N_9722);
nand U10937 (N_10937,N_9972,N_9315);
nand U10938 (N_10938,N_9076,N_9729);
or U10939 (N_10939,N_9522,N_9535);
or U10940 (N_10940,N_9889,N_9564);
or U10941 (N_10941,N_9698,N_9561);
nand U10942 (N_10942,N_9923,N_9065);
xnor U10943 (N_10943,N_9253,N_9698);
or U10944 (N_10944,N_9484,N_9798);
or U10945 (N_10945,N_9416,N_9107);
nor U10946 (N_10946,N_9068,N_9381);
or U10947 (N_10947,N_9089,N_9553);
and U10948 (N_10948,N_9551,N_9876);
and U10949 (N_10949,N_9720,N_9261);
or U10950 (N_10950,N_9790,N_9225);
xnor U10951 (N_10951,N_9590,N_9907);
nand U10952 (N_10952,N_9140,N_9806);
and U10953 (N_10953,N_9860,N_9473);
and U10954 (N_10954,N_9766,N_9512);
xnor U10955 (N_10955,N_9282,N_9850);
nand U10956 (N_10956,N_9392,N_9443);
and U10957 (N_10957,N_9943,N_9082);
and U10958 (N_10958,N_9285,N_9436);
xor U10959 (N_10959,N_9967,N_9713);
and U10960 (N_10960,N_9969,N_9463);
or U10961 (N_10961,N_9665,N_9089);
nand U10962 (N_10962,N_9241,N_9150);
xnor U10963 (N_10963,N_9624,N_9440);
xnor U10964 (N_10964,N_9717,N_9568);
nor U10965 (N_10965,N_9815,N_9699);
or U10966 (N_10966,N_9945,N_9254);
and U10967 (N_10967,N_9739,N_9177);
nor U10968 (N_10968,N_9598,N_9158);
or U10969 (N_10969,N_9429,N_9598);
and U10970 (N_10970,N_9494,N_9484);
nand U10971 (N_10971,N_9741,N_9364);
nor U10972 (N_10972,N_9783,N_9875);
or U10973 (N_10973,N_9359,N_9871);
xnor U10974 (N_10974,N_9944,N_9635);
and U10975 (N_10975,N_9927,N_9093);
nand U10976 (N_10976,N_9360,N_9646);
nor U10977 (N_10977,N_9310,N_9330);
nor U10978 (N_10978,N_9543,N_9730);
xor U10979 (N_10979,N_9498,N_9966);
nand U10980 (N_10980,N_9896,N_9154);
xor U10981 (N_10981,N_9370,N_9752);
nand U10982 (N_10982,N_9148,N_9524);
nand U10983 (N_10983,N_9325,N_9950);
or U10984 (N_10984,N_9289,N_9252);
nor U10985 (N_10985,N_9144,N_9233);
or U10986 (N_10986,N_9478,N_9364);
nand U10987 (N_10987,N_9667,N_9840);
nand U10988 (N_10988,N_9631,N_9785);
nor U10989 (N_10989,N_9893,N_9101);
and U10990 (N_10990,N_9829,N_9732);
xor U10991 (N_10991,N_9496,N_9856);
nand U10992 (N_10992,N_9811,N_9309);
xnor U10993 (N_10993,N_9940,N_9556);
and U10994 (N_10994,N_9343,N_9450);
xor U10995 (N_10995,N_9369,N_9700);
xnor U10996 (N_10996,N_9813,N_9884);
nor U10997 (N_10997,N_9404,N_9779);
and U10998 (N_10998,N_9400,N_9283);
nand U10999 (N_10999,N_9326,N_9384);
xor U11000 (N_11000,N_10770,N_10574);
xnor U11001 (N_11001,N_10436,N_10157);
and U11002 (N_11002,N_10365,N_10227);
or U11003 (N_11003,N_10091,N_10177);
and U11004 (N_11004,N_10487,N_10355);
or U11005 (N_11005,N_10404,N_10794);
or U11006 (N_11006,N_10951,N_10644);
nand U11007 (N_11007,N_10788,N_10041);
and U11008 (N_11008,N_10996,N_10843);
and U11009 (N_11009,N_10350,N_10403);
and U11010 (N_11010,N_10988,N_10978);
nand U11011 (N_11011,N_10182,N_10834);
nand U11012 (N_11012,N_10952,N_10336);
nor U11013 (N_11013,N_10603,N_10594);
nand U11014 (N_11014,N_10322,N_10194);
nand U11015 (N_11015,N_10765,N_10946);
nor U11016 (N_11016,N_10650,N_10107);
and U11017 (N_11017,N_10887,N_10238);
xor U11018 (N_11018,N_10721,N_10888);
xor U11019 (N_11019,N_10954,N_10400);
and U11020 (N_11020,N_10936,N_10640);
xor U11021 (N_11021,N_10993,N_10595);
xor U11022 (N_11022,N_10375,N_10851);
nand U11023 (N_11023,N_10009,N_10926);
nand U11024 (N_11024,N_10327,N_10195);
nand U11025 (N_11025,N_10933,N_10221);
nand U11026 (N_11026,N_10256,N_10529);
nor U11027 (N_11027,N_10781,N_10496);
nand U11028 (N_11028,N_10492,N_10373);
nor U11029 (N_11029,N_10903,N_10695);
nand U11030 (N_11030,N_10393,N_10074);
xnor U11031 (N_11031,N_10534,N_10729);
nor U11032 (N_11032,N_10555,N_10663);
xnor U11033 (N_11033,N_10583,N_10390);
nand U11034 (N_11034,N_10550,N_10176);
and U11035 (N_11035,N_10518,N_10384);
nand U11036 (N_11036,N_10615,N_10066);
nand U11037 (N_11037,N_10179,N_10522);
nor U11038 (N_11038,N_10573,N_10808);
xor U11039 (N_11039,N_10323,N_10697);
nand U11040 (N_11040,N_10245,N_10764);
nand U11041 (N_11041,N_10995,N_10832);
xor U11042 (N_11042,N_10304,N_10798);
nand U11043 (N_11043,N_10532,N_10280);
nor U11044 (N_11044,N_10171,N_10253);
and U11045 (N_11045,N_10067,N_10088);
xor U11046 (N_11046,N_10859,N_10466);
nor U11047 (N_11047,N_10477,N_10810);
nand U11048 (N_11048,N_10866,N_10144);
or U11049 (N_11049,N_10514,N_10479);
and U11050 (N_11050,N_10448,N_10818);
nor U11051 (N_11051,N_10052,N_10830);
or U11052 (N_11052,N_10209,N_10192);
or U11053 (N_11053,N_10269,N_10688);
and U11054 (N_11054,N_10505,N_10848);
nor U11055 (N_11055,N_10320,N_10910);
nor U11056 (N_11056,N_10478,N_10472);
and U11057 (N_11057,N_10005,N_10498);
xor U11058 (N_11058,N_10298,N_10000);
or U11059 (N_11059,N_10608,N_10367);
or U11060 (N_11060,N_10998,N_10060);
xnor U11061 (N_11061,N_10878,N_10019);
nor U11062 (N_11062,N_10733,N_10230);
nor U11063 (N_11063,N_10699,N_10755);
and U11064 (N_11064,N_10839,N_10405);
nor U11065 (N_11065,N_10175,N_10307);
and U11066 (N_11066,N_10124,N_10528);
nand U11067 (N_11067,N_10321,N_10677);
nor U11068 (N_11068,N_10345,N_10912);
xor U11069 (N_11069,N_10348,N_10070);
or U11070 (N_11070,N_10357,N_10485);
and U11071 (N_11071,N_10480,N_10940);
xor U11072 (N_11072,N_10205,N_10189);
or U11073 (N_11073,N_10835,N_10117);
nand U11074 (N_11074,N_10805,N_10791);
nand U11075 (N_11075,N_10215,N_10605);
xor U11076 (N_11076,N_10491,N_10914);
or U11077 (N_11077,N_10017,N_10763);
nor U11078 (N_11078,N_10658,N_10310);
xnor U11079 (N_11079,N_10389,N_10619);
nand U11080 (N_11080,N_10982,N_10539);
nor U11081 (N_11081,N_10642,N_10265);
or U11082 (N_11082,N_10493,N_10531);
nand U11083 (N_11083,N_10795,N_10294);
and U11084 (N_11084,N_10451,N_10266);
or U11085 (N_11085,N_10533,N_10001);
xnor U11086 (N_11086,N_10787,N_10628);
or U11087 (N_11087,N_10409,N_10879);
nand U11088 (N_11088,N_10128,N_10186);
and U11089 (N_11089,N_10447,N_10981);
or U11090 (N_11090,N_10726,N_10458);
xor U11091 (N_11091,N_10031,N_10443);
nand U11092 (N_11092,N_10698,N_10500);
nor U11093 (N_11093,N_10849,N_10377);
nor U11094 (N_11094,N_10140,N_10928);
nand U11095 (N_11095,N_10095,N_10228);
xnor U11096 (N_11096,N_10752,N_10735);
or U11097 (N_11097,N_10356,N_10481);
nor U11098 (N_11098,N_10246,N_10809);
nand U11099 (N_11099,N_10609,N_10692);
xnor U11100 (N_11100,N_10068,N_10984);
nor U11101 (N_11101,N_10340,N_10065);
nand U11102 (N_11102,N_10651,N_10652);
xnor U11103 (N_11103,N_10872,N_10180);
xor U11104 (N_11104,N_10217,N_10613);
or U11105 (N_11105,N_10351,N_10199);
or U11106 (N_11106,N_10836,N_10793);
nand U11107 (N_11107,N_10643,N_10754);
xor U11108 (N_11108,N_10125,N_10890);
nand U11109 (N_11109,N_10801,N_10164);
and U11110 (N_11110,N_10596,N_10856);
nor U11111 (N_11111,N_10722,N_10100);
or U11112 (N_11112,N_10827,N_10459);
nor U11113 (N_11113,N_10414,N_10271);
xor U11114 (N_11114,N_10693,N_10673);
nand U11115 (N_11115,N_10967,N_10150);
or U11116 (N_11116,N_10681,N_10667);
nand U11117 (N_11117,N_10371,N_10965);
xor U11118 (N_11118,N_10482,N_10274);
nor U11119 (N_11119,N_10049,N_10937);
xnor U11120 (N_11120,N_10899,N_10994);
nand U11121 (N_11121,N_10167,N_10366);
nand U11122 (N_11122,N_10840,N_10876);
nand U11123 (N_11123,N_10886,N_10495);
nor U11124 (N_11124,N_10076,N_10907);
or U11125 (N_11125,N_10331,N_10904);
nand U11126 (N_11126,N_10063,N_10947);
nor U11127 (N_11127,N_10625,N_10523);
xor U11128 (N_11128,N_10465,N_10762);
nand U11129 (N_11129,N_10515,N_10376);
or U11130 (N_11130,N_10551,N_10425);
xnor U11131 (N_11131,N_10489,N_10773);
nand U11132 (N_11132,N_10558,N_10397);
or U11133 (N_11133,N_10338,N_10790);
and U11134 (N_11134,N_10272,N_10044);
nor U11135 (N_11135,N_10509,N_10062);
xnor U11136 (N_11136,N_10567,N_10169);
or U11137 (N_11137,N_10724,N_10694);
and U11138 (N_11138,N_10637,N_10882);
or U11139 (N_11139,N_10889,N_10126);
xnor U11140 (N_11140,N_10446,N_10138);
xor U11141 (N_11141,N_10742,N_10906);
and U11142 (N_11142,N_10873,N_10418);
or U11143 (N_11143,N_10391,N_10855);
or U11144 (N_11144,N_10083,N_10399);
and U11145 (N_11145,N_10109,N_10602);
or U11146 (N_11146,N_10584,N_10864);
xnor U11147 (N_11147,N_10197,N_10792);
nor U11148 (N_11148,N_10557,N_10381);
xor U11149 (N_11149,N_10814,N_10885);
and U11150 (N_11150,N_10168,N_10290);
xnor U11151 (N_11151,N_10131,N_10641);
and U11152 (N_11152,N_10507,N_10449);
and U11153 (N_11153,N_10213,N_10181);
nor U11154 (N_11154,N_10368,N_10302);
and U11155 (N_11155,N_10282,N_10714);
xnor U11156 (N_11156,N_10284,N_10084);
nor U11157 (N_11157,N_10353,N_10428);
or U11158 (N_11158,N_10212,N_10015);
or U11159 (N_11159,N_10438,N_10080);
nand U11160 (N_11160,N_10612,N_10162);
xnor U11161 (N_11161,N_10717,N_10004);
xor U11162 (N_11162,N_10313,N_10276);
or U11163 (N_11163,N_10342,N_10690);
nor U11164 (N_11164,N_10318,N_10917);
nand U11165 (N_11165,N_10631,N_10121);
and U11166 (N_11166,N_10536,N_10160);
xnor U11167 (N_11167,N_10308,N_10152);
and U11168 (N_11168,N_10564,N_10614);
and U11169 (N_11169,N_10582,N_10785);
nand U11170 (N_11170,N_10561,N_10032);
nand U11171 (N_11171,N_10546,N_10270);
nand U11172 (N_11172,N_10905,N_10789);
xnor U11173 (N_11173,N_10746,N_10920);
xor U11174 (N_11174,N_10737,N_10516);
and U11175 (N_11175,N_10973,N_10254);
or U11176 (N_11176,N_10782,N_10151);
nand U11177 (N_11177,N_10863,N_10277);
and U11178 (N_11178,N_10589,N_10155);
and U11179 (N_11179,N_10286,N_10330);
nand U11180 (N_11180,N_10211,N_10382);
or U11181 (N_11181,N_10016,N_10847);
nand U11182 (N_11182,N_10780,N_10841);
nor U11183 (N_11183,N_10300,N_10547);
xnor U11184 (N_11184,N_10328,N_10966);
nand U11185 (N_11185,N_10442,N_10105);
nand U11186 (N_11186,N_10666,N_10706);
nor U11187 (N_11187,N_10526,N_10172);
or U11188 (N_11188,N_10343,N_10895);
and U11189 (N_11189,N_10852,N_10020);
nor U11190 (N_11190,N_10646,N_10476);
nand U11191 (N_11191,N_10241,N_10196);
and U11192 (N_11192,N_10548,N_10985);
nand U11193 (N_11193,N_10587,N_10796);
or U11194 (N_11194,N_10440,N_10960);
and U11195 (N_11195,N_10829,N_10048);
nand U11196 (N_11196,N_10456,N_10970);
and U11197 (N_11197,N_10054,N_10287);
nor U11198 (N_11198,N_10311,N_10623);
and U11199 (N_11199,N_10053,N_10090);
xnor U11200 (N_11200,N_10296,N_10850);
and U11201 (N_11201,N_10111,N_10305);
xnor U11202 (N_11202,N_10352,N_10103);
nor U11203 (N_11203,N_10725,N_10606);
and U11204 (N_11204,N_10379,N_10112);
or U11205 (N_11205,N_10624,N_10831);
or U11206 (N_11206,N_10134,N_10204);
nand U11207 (N_11207,N_10736,N_10193);
nor U11208 (N_11208,N_10158,N_10362);
xor U11209 (N_11209,N_10648,N_10133);
or U11210 (N_11210,N_10122,N_10378);
xor U11211 (N_11211,N_10950,N_10671);
xnor U11212 (N_11212,N_10082,N_10747);
xor U11213 (N_11213,N_10453,N_10219);
and U11214 (N_11214,N_10075,N_10408);
nor U11215 (N_11215,N_10233,N_10325);
nand U11216 (N_11216,N_10249,N_10638);
or U11217 (N_11217,N_10139,N_10943);
nor U11218 (N_11218,N_10335,N_10388);
and U11219 (N_11219,N_10099,N_10702);
or U11220 (N_11220,N_10113,N_10187);
xnor U11221 (N_11221,N_10712,N_10517);
nor U11222 (N_11222,N_10751,N_10439);
nor U11223 (N_11223,N_10469,N_10415);
nand U11224 (N_11224,N_10042,N_10653);
nand U11225 (N_11225,N_10844,N_10929);
and U11226 (N_11226,N_10329,N_10444);
xor U11227 (N_11227,N_10045,N_10865);
and U11228 (N_11228,N_10869,N_10347);
nor U11229 (N_11229,N_10108,N_10087);
and U11230 (N_11230,N_10069,N_10279);
or U11231 (N_11231,N_10046,N_10508);
xnor U11232 (N_11232,N_10437,N_10288);
xor U11233 (N_11233,N_10813,N_10190);
nor U11234 (N_11234,N_10527,N_10760);
nor U11235 (N_11235,N_10301,N_10815);
nand U11236 (N_11236,N_10749,N_10064);
and U11237 (N_11237,N_10766,N_10986);
and U11238 (N_11238,N_10894,N_10433);
and U11239 (N_11239,N_10260,N_10774);
nor U11240 (N_11240,N_10344,N_10104);
nor U11241 (N_11241,N_10661,N_10445);
nand U11242 (N_11242,N_10394,N_10188);
nand U11243 (N_11243,N_10333,N_10545);
nand U11244 (N_11244,N_10756,N_10707);
xnor U11245 (N_11245,N_10452,N_10251);
xor U11246 (N_11246,N_10314,N_10918);
nor U11247 (N_11247,N_10559,N_10079);
xor U11248 (N_11248,N_10908,N_10038);
nor U11249 (N_11249,N_10685,N_10392);
nor U11250 (N_11250,N_10833,N_10842);
xnor U11251 (N_11251,N_10426,N_10891);
nand U11252 (N_11252,N_10524,N_10374);
and U11253 (N_11253,N_10326,N_10925);
nand U11254 (N_11254,N_10040,N_10012);
or U11255 (N_11255,N_10097,N_10145);
xor U11256 (N_11256,N_10923,N_10556);
or U11257 (N_11257,N_10183,N_10096);
nor U11258 (N_11258,N_10576,N_10184);
nand U11259 (N_11259,N_10002,N_10924);
xor U11260 (N_11260,N_10569,N_10964);
and U11261 (N_11261,N_10291,N_10146);
nand U11262 (N_11262,N_10473,N_10784);
and U11263 (N_11263,N_10817,N_10043);
or U11264 (N_11264,N_10728,N_10474);
or U11265 (N_11265,N_10022,N_10137);
nand U11266 (N_11266,N_10039,N_10106);
nand U11267 (N_11267,N_10922,N_10475);
or U11268 (N_11268,N_10421,N_10319);
xnor U11269 (N_11269,N_10216,N_10123);
and U11270 (N_11270,N_10115,N_10092);
or U11271 (N_11271,N_10191,N_10708);
nand U11272 (N_11272,N_10881,N_10220);
nor U11273 (N_11273,N_10285,N_10262);
nor U11274 (N_11274,N_10570,N_10972);
xor U11275 (N_11275,N_10141,N_10315);
nor U11276 (N_11276,N_10396,N_10597);
or U11277 (N_11277,N_10114,N_10825);
and U11278 (N_11278,N_10130,N_10501);
and U11279 (N_11279,N_10208,N_10713);
xnor U11280 (N_11280,N_10530,N_10292);
nand U11281 (N_11281,N_10316,N_10143);
nor U11282 (N_11282,N_10739,N_10525);
or U11283 (N_11283,N_10948,N_10059);
and U11284 (N_11284,N_10240,N_10727);
or U11285 (N_11285,N_10976,N_10156);
and U11286 (N_11286,N_10237,N_10701);
xor U11287 (N_11287,N_10730,N_10147);
nand U11288 (N_11288,N_10035,N_10281);
nand U11289 (N_11289,N_10731,N_10880);
or U11290 (N_11290,N_10497,N_10716);
and U11291 (N_11291,N_10222,N_10243);
or U11292 (N_11292,N_10011,N_10503);
nor U11293 (N_11293,N_10600,N_10334);
xnor U11294 (N_11294,N_10369,N_10013);
nand U11295 (N_11295,N_10461,N_10575);
xor U11296 (N_11296,N_10588,N_10098);
and U11297 (N_11297,N_10586,N_10771);
and U11298 (N_11298,N_10242,N_10629);
xor U11299 (N_11299,N_10684,N_10902);
and U11300 (N_11300,N_10683,N_10682);
xor U11301 (N_11301,N_10380,N_10846);
xnor U11302 (N_11302,N_10753,N_10413);
nor U11303 (N_11303,N_10838,N_10610);
or U11304 (N_11304,N_10089,N_10457);
xor U11305 (N_11305,N_10185,N_10868);
or U11306 (N_11306,N_10293,N_10704);
nand U11307 (N_11307,N_10938,N_10406);
nand U11308 (N_11308,N_10268,N_10900);
xor U11309 (N_11309,N_10823,N_10423);
xor U11310 (N_11310,N_10029,N_10626);
or U11311 (N_11311,N_10153,N_10883);
xor U11312 (N_11312,N_10662,N_10630);
nand U11313 (N_11313,N_10897,N_10971);
and U11314 (N_11314,N_10974,N_10871);
and U11315 (N_11315,N_10968,N_10804);
xor U11316 (N_11316,N_10420,N_10454);
xnor U11317 (N_11317,N_10927,N_10299);
nor U11318 (N_11318,N_10675,N_10161);
nand U11319 (N_11319,N_10259,N_10455);
xnor U11320 (N_11320,N_10854,N_10027);
or U11321 (N_11321,N_10520,N_10008);
nor U11322 (N_11322,N_10306,N_10511);
and U11323 (N_11323,N_10398,N_10734);
nand U11324 (N_11324,N_10828,N_10257);
xor U11325 (N_11325,N_10030,N_10655);
or U11326 (N_11326,N_10538,N_10510);
or U11327 (N_11327,N_10935,N_10003);
nor U11328 (N_11328,N_10119,N_10349);
xnor U11329 (N_11329,N_10488,N_10429);
nand U11330 (N_11330,N_10802,N_10148);
nor U11331 (N_11331,N_10687,N_10544);
nor U11332 (N_11332,N_10990,N_10401);
xnor U11333 (N_11333,N_10358,N_10077);
nor U11334 (N_11334,N_10991,N_10512);
xor U11335 (N_11335,N_10467,N_10963);
and U11336 (N_11336,N_10800,N_10593);
nor U11337 (N_11337,N_10709,N_10740);
nor U11338 (N_11338,N_10416,N_10225);
nand U11339 (N_11339,N_10072,N_10235);
nor U11340 (N_11340,N_10598,N_10361);
xnor U11341 (N_11341,N_10686,N_10419);
or U11342 (N_11342,N_10432,N_10541);
and U11343 (N_11343,N_10332,N_10585);
xnor U11344 (N_11344,N_10395,N_10961);
xnor U11345 (N_11345,N_10464,N_10247);
and U11346 (N_11346,N_10231,N_10135);
xnor U11347 (N_11347,N_10580,N_10599);
nand U11348 (N_11348,N_10620,N_10711);
nand U11349 (N_11349,N_10255,N_10198);
and U11350 (N_11350,N_10086,N_10261);
nor U11351 (N_11351,N_10672,N_10424);
nand U11352 (N_11352,N_10056,N_10434);
nand U11353 (N_11353,N_10867,N_10860);
nor U11354 (N_11354,N_10218,N_10521);
and U11355 (N_11355,N_10581,N_10207);
xnor U11356 (N_11356,N_10962,N_10163);
xor U11357 (N_11357,N_10519,N_10178);
or U11358 (N_11358,N_10861,N_10006);
xnor U11359 (N_11359,N_10337,N_10719);
xor U11360 (N_11360,N_10223,N_10411);
or U11361 (N_11361,N_10635,N_10942);
and U11362 (N_11362,N_10647,N_10670);
or U11363 (N_11363,N_10370,N_10010);
nand U11364 (N_11364,N_10656,N_10870);
nand U11365 (N_11365,N_10921,N_10543);
nand U11366 (N_11366,N_10824,N_10094);
nor U11367 (N_11367,N_10592,N_10776);
and U11368 (N_11368,N_10214,N_10892);
xnor U11369 (N_11369,N_10422,N_10295);
nor U11370 (N_11370,N_10578,N_10346);
or U11371 (N_11371,N_10779,N_10050);
and U11372 (N_11372,N_10992,N_10483);
and U11373 (N_11373,N_10470,N_10901);
nand U11374 (N_11374,N_10412,N_10387);
or U11375 (N_11375,N_10120,N_10034);
or U11376 (N_11376,N_10654,N_10462);
or U11377 (N_11377,N_10427,N_10226);
xnor U11378 (N_11378,N_10816,N_10590);
or U11379 (N_11379,N_10649,N_10939);
xor U11380 (N_11380,N_10775,N_10980);
and U11381 (N_11381,N_10837,N_10759);
and U11382 (N_11382,N_10786,N_10136);
or U11383 (N_11383,N_10149,N_10761);
or U11384 (N_11384,N_10468,N_10577);
xnor U11385 (N_11385,N_10664,N_10263);
and U11386 (N_11386,N_10499,N_10118);
xor U11387 (N_11387,N_10073,N_10748);
nand U11388 (N_11388,N_10165,N_10407);
nor U11389 (N_11389,N_10772,N_10679);
nor U11390 (N_11390,N_10689,N_10875);
xnor U11391 (N_11391,N_10504,N_10078);
and U11392 (N_11392,N_10660,N_10058);
and U11393 (N_11393,N_10057,N_10142);
xor U11394 (N_11394,N_10055,N_10081);
nand U11395 (N_11395,N_10705,N_10821);
and U11396 (N_11396,N_10363,N_10537);
nor U11397 (N_11397,N_10668,N_10819);
xnor U11398 (N_11398,N_10025,N_10703);
nor U11399 (N_11399,N_10680,N_10506);
xor U11400 (N_11400,N_10979,N_10745);
nand U11401 (N_11401,N_10502,N_10639);
xor U11402 (N_11402,N_10958,N_10258);
xor U11403 (N_11403,N_10460,N_10777);
xnor U11404 (N_11404,N_10959,N_10845);
xor U11405 (N_11405,N_10633,N_10732);
and U11406 (N_11406,N_10718,N_10093);
xor U11407 (N_11407,N_10715,N_10758);
and U11408 (N_11408,N_10159,N_10601);
nor U11409 (N_11409,N_10811,N_10036);
nand U11410 (N_11410,N_10743,N_10486);
nor U11411 (N_11411,N_10206,N_10239);
nor U11412 (N_11412,N_10007,N_10252);
and U11413 (N_11413,N_10862,N_10248);
nand U11414 (N_11414,N_10132,N_10553);
xnor U11415 (N_11415,N_10385,N_10303);
and U11416 (N_11416,N_10028,N_10566);
or U11417 (N_11417,N_10540,N_10441);
or U11418 (N_11418,N_10744,N_10750);
or U11419 (N_11419,N_10858,N_10450);
and U11420 (N_11420,N_10023,N_10560);
or U11421 (N_11421,N_10607,N_10312);
and U11422 (N_11422,N_10604,N_10676);
nand U11423 (N_11423,N_10826,N_10154);
xnor U11424 (N_11424,N_10033,N_10278);
nor U11425 (N_11425,N_10579,N_10571);
and U11426 (N_11426,N_10360,N_10987);
nand U11427 (N_11427,N_10757,N_10977);
xor U11428 (N_11428,N_10955,N_10621);
xor U11429 (N_11429,N_10021,N_10919);
xor U11430 (N_11430,N_10909,N_10014);
and U11431 (N_11431,N_10953,N_10224);
xor U11432 (N_11432,N_10250,N_10769);
and U11433 (N_11433,N_10949,N_10202);
xor U11434 (N_11434,N_10024,N_10657);
xnor U11435 (N_11435,N_10616,N_10116);
xnor U11436 (N_11436,N_10803,N_10691);
or U11437 (N_11437,N_10916,N_10174);
and U11438 (N_11438,N_10431,N_10203);
and U11439 (N_11439,N_10513,N_10857);
and U11440 (N_11440,N_10723,N_10047);
nor U11441 (N_11441,N_10562,N_10463);
or U11442 (N_11442,N_10309,N_10283);
and U11443 (N_11443,N_10234,N_10244);
nand U11444 (N_11444,N_10359,N_10110);
or U11445 (N_11445,N_10768,N_10129);
nor U11446 (N_11446,N_10201,N_10051);
xor U11447 (N_11447,N_10417,N_10710);
and U11448 (N_11448,N_10572,N_10778);
and U11449 (N_11449,N_10364,N_10822);
and U11450 (N_11450,N_10934,N_10273);
xnor U11451 (N_11451,N_10893,N_10275);
and U11452 (N_11452,N_10799,N_10037);
and U11453 (N_11453,N_10200,N_10535);
or U11454 (N_11454,N_10665,N_10669);
nor U11455 (N_11455,N_10071,N_10944);
nor U11456 (N_11456,N_10645,N_10884);
nand U11457 (N_11457,N_10568,N_10264);
nor U11458 (N_11458,N_10552,N_10297);
and U11459 (N_11459,N_10170,N_10941);
nor U11460 (N_11460,N_10591,N_10983);
nor U11461 (N_11461,N_10173,N_10783);
nor U11462 (N_11462,N_10678,N_10435);
xor U11463 (N_11463,N_10896,N_10324);
nand U11464 (N_11464,N_10957,N_10611);
nand U11465 (N_11465,N_10915,N_10026);
and U11466 (N_11466,N_10969,N_10738);
nor U11467 (N_11467,N_10565,N_10101);
nor U11468 (N_11468,N_10636,N_10807);
nor U11469 (N_11469,N_10989,N_10632);
nor U11470 (N_11470,N_10853,N_10797);
or U11471 (N_11471,N_10618,N_10806);
nand U11472 (N_11472,N_10563,N_10236);
nand U11473 (N_11473,N_10354,N_10490);
xnor U11474 (N_11474,N_10554,N_10471);
or U11475 (N_11475,N_10430,N_10874);
xnor U11476 (N_11476,N_10767,N_10627);
and U11477 (N_11477,N_10341,N_10267);
xor U11478 (N_11478,N_10210,N_10911);
xor U11479 (N_11479,N_10931,N_10339);
nor U11480 (N_11480,N_10085,N_10930);
nor U11481 (N_11481,N_10956,N_10542);
and U11482 (N_11482,N_10317,N_10700);
and U11483 (N_11483,N_10127,N_10674);
or U11484 (N_11484,N_10386,N_10877);
nor U11485 (N_11485,N_10820,N_10289);
and U11486 (N_11486,N_10372,N_10484);
or U11487 (N_11487,N_10997,N_10232);
nand U11488 (N_11488,N_10494,N_10812);
or U11489 (N_11489,N_10549,N_10018);
and U11490 (N_11490,N_10898,N_10402);
xnor U11491 (N_11491,N_10061,N_10229);
or U11492 (N_11492,N_10383,N_10696);
and U11493 (N_11493,N_10932,N_10720);
nand U11494 (N_11494,N_10634,N_10975);
nand U11495 (N_11495,N_10410,N_10913);
nand U11496 (N_11496,N_10617,N_10945);
xnor U11497 (N_11497,N_10102,N_10741);
or U11498 (N_11498,N_10622,N_10166);
xor U11499 (N_11499,N_10999,N_10659);
nand U11500 (N_11500,N_10778,N_10611);
nor U11501 (N_11501,N_10200,N_10500);
nand U11502 (N_11502,N_10247,N_10015);
nor U11503 (N_11503,N_10742,N_10189);
nand U11504 (N_11504,N_10310,N_10674);
xor U11505 (N_11505,N_10462,N_10894);
or U11506 (N_11506,N_10003,N_10419);
and U11507 (N_11507,N_10118,N_10356);
or U11508 (N_11508,N_10533,N_10017);
xor U11509 (N_11509,N_10492,N_10708);
nand U11510 (N_11510,N_10684,N_10876);
or U11511 (N_11511,N_10654,N_10989);
or U11512 (N_11512,N_10058,N_10348);
nand U11513 (N_11513,N_10776,N_10867);
and U11514 (N_11514,N_10579,N_10785);
nor U11515 (N_11515,N_10483,N_10897);
nor U11516 (N_11516,N_10878,N_10766);
or U11517 (N_11517,N_10400,N_10130);
nand U11518 (N_11518,N_10036,N_10869);
nor U11519 (N_11519,N_10370,N_10850);
nand U11520 (N_11520,N_10368,N_10715);
nor U11521 (N_11521,N_10714,N_10018);
nand U11522 (N_11522,N_10057,N_10996);
xor U11523 (N_11523,N_10297,N_10788);
and U11524 (N_11524,N_10207,N_10505);
nor U11525 (N_11525,N_10845,N_10514);
nor U11526 (N_11526,N_10884,N_10035);
xnor U11527 (N_11527,N_10128,N_10173);
xor U11528 (N_11528,N_10567,N_10991);
nand U11529 (N_11529,N_10897,N_10315);
xnor U11530 (N_11530,N_10640,N_10495);
xor U11531 (N_11531,N_10344,N_10132);
and U11532 (N_11532,N_10677,N_10864);
xnor U11533 (N_11533,N_10875,N_10853);
nor U11534 (N_11534,N_10516,N_10098);
and U11535 (N_11535,N_10281,N_10983);
or U11536 (N_11536,N_10891,N_10885);
nor U11537 (N_11537,N_10971,N_10547);
xnor U11538 (N_11538,N_10294,N_10041);
and U11539 (N_11539,N_10667,N_10848);
xnor U11540 (N_11540,N_10266,N_10090);
or U11541 (N_11541,N_10298,N_10784);
and U11542 (N_11542,N_10892,N_10655);
nand U11543 (N_11543,N_10819,N_10973);
xor U11544 (N_11544,N_10215,N_10648);
and U11545 (N_11545,N_10040,N_10573);
or U11546 (N_11546,N_10512,N_10340);
or U11547 (N_11547,N_10914,N_10689);
or U11548 (N_11548,N_10081,N_10532);
nand U11549 (N_11549,N_10825,N_10099);
xor U11550 (N_11550,N_10826,N_10867);
nor U11551 (N_11551,N_10807,N_10128);
nor U11552 (N_11552,N_10447,N_10889);
or U11553 (N_11553,N_10354,N_10047);
or U11554 (N_11554,N_10076,N_10142);
nor U11555 (N_11555,N_10962,N_10032);
and U11556 (N_11556,N_10055,N_10059);
xor U11557 (N_11557,N_10944,N_10676);
and U11558 (N_11558,N_10046,N_10918);
and U11559 (N_11559,N_10676,N_10678);
nand U11560 (N_11560,N_10726,N_10736);
or U11561 (N_11561,N_10053,N_10852);
and U11562 (N_11562,N_10958,N_10396);
and U11563 (N_11563,N_10233,N_10098);
xnor U11564 (N_11564,N_10003,N_10784);
xor U11565 (N_11565,N_10734,N_10505);
xor U11566 (N_11566,N_10736,N_10212);
and U11567 (N_11567,N_10888,N_10693);
nor U11568 (N_11568,N_10203,N_10510);
or U11569 (N_11569,N_10553,N_10628);
or U11570 (N_11570,N_10698,N_10988);
xnor U11571 (N_11571,N_10355,N_10526);
and U11572 (N_11572,N_10537,N_10882);
nand U11573 (N_11573,N_10097,N_10047);
or U11574 (N_11574,N_10480,N_10316);
nand U11575 (N_11575,N_10602,N_10220);
and U11576 (N_11576,N_10411,N_10456);
and U11577 (N_11577,N_10981,N_10432);
xor U11578 (N_11578,N_10684,N_10225);
and U11579 (N_11579,N_10677,N_10495);
xnor U11580 (N_11580,N_10910,N_10453);
and U11581 (N_11581,N_10959,N_10691);
xor U11582 (N_11582,N_10321,N_10073);
or U11583 (N_11583,N_10437,N_10147);
and U11584 (N_11584,N_10385,N_10309);
and U11585 (N_11585,N_10319,N_10241);
or U11586 (N_11586,N_10946,N_10858);
nor U11587 (N_11587,N_10224,N_10603);
and U11588 (N_11588,N_10225,N_10170);
and U11589 (N_11589,N_10387,N_10193);
nor U11590 (N_11590,N_10945,N_10616);
or U11591 (N_11591,N_10401,N_10527);
and U11592 (N_11592,N_10302,N_10734);
or U11593 (N_11593,N_10769,N_10357);
or U11594 (N_11594,N_10607,N_10139);
or U11595 (N_11595,N_10213,N_10305);
or U11596 (N_11596,N_10903,N_10966);
nand U11597 (N_11597,N_10182,N_10537);
and U11598 (N_11598,N_10890,N_10700);
xor U11599 (N_11599,N_10527,N_10512);
nand U11600 (N_11600,N_10879,N_10391);
nand U11601 (N_11601,N_10612,N_10029);
nand U11602 (N_11602,N_10652,N_10315);
nor U11603 (N_11603,N_10137,N_10825);
and U11604 (N_11604,N_10231,N_10182);
nor U11605 (N_11605,N_10326,N_10613);
and U11606 (N_11606,N_10238,N_10821);
nand U11607 (N_11607,N_10553,N_10258);
nor U11608 (N_11608,N_10144,N_10423);
or U11609 (N_11609,N_10005,N_10952);
nand U11610 (N_11610,N_10411,N_10856);
nand U11611 (N_11611,N_10817,N_10368);
nor U11612 (N_11612,N_10127,N_10361);
nand U11613 (N_11613,N_10675,N_10736);
xor U11614 (N_11614,N_10381,N_10220);
and U11615 (N_11615,N_10104,N_10793);
or U11616 (N_11616,N_10211,N_10622);
or U11617 (N_11617,N_10071,N_10697);
nor U11618 (N_11618,N_10929,N_10792);
xnor U11619 (N_11619,N_10392,N_10053);
nor U11620 (N_11620,N_10733,N_10402);
nor U11621 (N_11621,N_10280,N_10862);
xor U11622 (N_11622,N_10654,N_10511);
or U11623 (N_11623,N_10283,N_10024);
or U11624 (N_11624,N_10618,N_10529);
xor U11625 (N_11625,N_10874,N_10644);
and U11626 (N_11626,N_10380,N_10610);
nand U11627 (N_11627,N_10778,N_10273);
or U11628 (N_11628,N_10343,N_10034);
xor U11629 (N_11629,N_10675,N_10615);
nor U11630 (N_11630,N_10499,N_10560);
nor U11631 (N_11631,N_10698,N_10723);
nand U11632 (N_11632,N_10683,N_10989);
nand U11633 (N_11633,N_10748,N_10012);
and U11634 (N_11634,N_10282,N_10591);
or U11635 (N_11635,N_10985,N_10317);
or U11636 (N_11636,N_10218,N_10281);
xor U11637 (N_11637,N_10123,N_10555);
xnor U11638 (N_11638,N_10233,N_10456);
and U11639 (N_11639,N_10485,N_10052);
nor U11640 (N_11640,N_10299,N_10101);
nor U11641 (N_11641,N_10160,N_10183);
nor U11642 (N_11642,N_10639,N_10662);
nor U11643 (N_11643,N_10915,N_10922);
nand U11644 (N_11644,N_10895,N_10223);
or U11645 (N_11645,N_10611,N_10793);
xnor U11646 (N_11646,N_10082,N_10127);
nand U11647 (N_11647,N_10383,N_10794);
and U11648 (N_11648,N_10649,N_10681);
xor U11649 (N_11649,N_10785,N_10353);
or U11650 (N_11650,N_10368,N_10226);
and U11651 (N_11651,N_10621,N_10970);
and U11652 (N_11652,N_10521,N_10679);
xnor U11653 (N_11653,N_10229,N_10082);
and U11654 (N_11654,N_10380,N_10211);
nor U11655 (N_11655,N_10198,N_10923);
and U11656 (N_11656,N_10729,N_10736);
or U11657 (N_11657,N_10923,N_10803);
nand U11658 (N_11658,N_10194,N_10116);
nor U11659 (N_11659,N_10803,N_10200);
xor U11660 (N_11660,N_10509,N_10598);
nor U11661 (N_11661,N_10888,N_10655);
xnor U11662 (N_11662,N_10137,N_10724);
or U11663 (N_11663,N_10539,N_10658);
xnor U11664 (N_11664,N_10824,N_10946);
nor U11665 (N_11665,N_10145,N_10387);
xor U11666 (N_11666,N_10207,N_10715);
nand U11667 (N_11667,N_10983,N_10056);
or U11668 (N_11668,N_10518,N_10164);
xor U11669 (N_11669,N_10668,N_10921);
xor U11670 (N_11670,N_10002,N_10221);
xnor U11671 (N_11671,N_10455,N_10364);
xor U11672 (N_11672,N_10284,N_10402);
and U11673 (N_11673,N_10720,N_10949);
nand U11674 (N_11674,N_10274,N_10316);
or U11675 (N_11675,N_10370,N_10715);
xor U11676 (N_11676,N_10595,N_10453);
or U11677 (N_11677,N_10244,N_10957);
or U11678 (N_11678,N_10049,N_10901);
or U11679 (N_11679,N_10318,N_10128);
nor U11680 (N_11680,N_10469,N_10245);
nand U11681 (N_11681,N_10347,N_10790);
or U11682 (N_11682,N_10156,N_10159);
or U11683 (N_11683,N_10886,N_10342);
or U11684 (N_11684,N_10684,N_10933);
nand U11685 (N_11685,N_10867,N_10749);
nand U11686 (N_11686,N_10519,N_10775);
xor U11687 (N_11687,N_10320,N_10928);
nor U11688 (N_11688,N_10691,N_10203);
nor U11689 (N_11689,N_10874,N_10010);
nor U11690 (N_11690,N_10860,N_10708);
or U11691 (N_11691,N_10043,N_10846);
xnor U11692 (N_11692,N_10720,N_10675);
or U11693 (N_11693,N_10344,N_10668);
and U11694 (N_11694,N_10042,N_10625);
xnor U11695 (N_11695,N_10362,N_10459);
or U11696 (N_11696,N_10936,N_10486);
xor U11697 (N_11697,N_10940,N_10922);
xnor U11698 (N_11698,N_10657,N_10059);
nand U11699 (N_11699,N_10857,N_10492);
or U11700 (N_11700,N_10025,N_10760);
nor U11701 (N_11701,N_10747,N_10884);
or U11702 (N_11702,N_10928,N_10156);
nor U11703 (N_11703,N_10466,N_10691);
nand U11704 (N_11704,N_10127,N_10915);
nor U11705 (N_11705,N_10732,N_10651);
and U11706 (N_11706,N_10668,N_10587);
or U11707 (N_11707,N_10056,N_10663);
nor U11708 (N_11708,N_10165,N_10171);
nand U11709 (N_11709,N_10712,N_10895);
or U11710 (N_11710,N_10815,N_10970);
or U11711 (N_11711,N_10819,N_10537);
and U11712 (N_11712,N_10863,N_10758);
nor U11713 (N_11713,N_10124,N_10240);
nand U11714 (N_11714,N_10649,N_10699);
nor U11715 (N_11715,N_10424,N_10927);
nor U11716 (N_11716,N_10717,N_10765);
xnor U11717 (N_11717,N_10041,N_10288);
and U11718 (N_11718,N_10696,N_10112);
nand U11719 (N_11719,N_10815,N_10160);
nand U11720 (N_11720,N_10209,N_10469);
xor U11721 (N_11721,N_10083,N_10912);
and U11722 (N_11722,N_10103,N_10622);
or U11723 (N_11723,N_10033,N_10089);
and U11724 (N_11724,N_10749,N_10192);
xnor U11725 (N_11725,N_10921,N_10207);
xnor U11726 (N_11726,N_10353,N_10550);
xor U11727 (N_11727,N_10749,N_10358);
nand U11728 (N_11728,N_10560,N_10438);
or U11729 (N_11729,N_10330,N_10457);
nor U11730 (N_11730,N_10249,N_10788);
and U11731 (N_11731,N_10462,N_10429);
nor U11732 (N_11732,N_10682,N_10485);
or U11733 (N_11733,N_10982,N_10571);
and U11734 (N_11734,N_10369,N_10768);
or U11735 (N_11735,N_10835,N_10144);
nand U11736 (N_11736,N_10003,N_10522);
and U11737 (N_11737,N_10280,N_10283);
xnor U11738 (N_11738,N_10562,N_10903);
and U11739 (N_11739,N_10989,N_10440);
and U11740 (N_11740,N_10788,N_10166);
xnor U11741 (N_11741,N_10275,N_10699);
xor U11742 (N_11742,N_10465,N_10601);
xor U11743 (N_11743,N_10600,N_10582);
xnor U11744 (N_11744,N_10802,N_10210);
nor U11745 (N_11745,N_10115,N_10487);
and U11746 (N_11746,N_10735,N_10926);
xor U11747 (N_11747,N_10581,N_10164);
or U11748 (N_11748,N_10730,N_10135);
nand U11749 (N_11749,N_10832,N_10176);
nand U11750 (N_11750,N_10453,N_10408);
and U11751 (N_11751,N_10675,N_10614);
nor U11752 (N_11752,N_10195,N_10377);
nor U11753 (N_11753,N_10200,N_10808);
and U11754 (N_11754,N_10909,N_10494);
or U11755 (N_11755,N_10465,N_10028);
or U11756 (N_11756,N_10268,N_10958);
or U11757 (N_11757,N_10882,N_10511);
nor U11758 (N_11758,N_10617,N_10032);
nand U11759 (N_11759,N_10569,N_10232);
nand U11760 (N_11760,N_10461,N_10252);
or U11761 (N_11761,N_10125,N_10848);
nand U11762 (N_11762,N_10494,N_10195);
and U11763 (N_11763,N_10824,N_10133);
and U11764 (N_11764,N_10186,N_10068);
xnor U11765 (N_11765,N_10821,N_10558);
nor U11766 (N_11766,N_10665,N_10466);
and U11767 (N_11767,N_10752,N_10237);
nor U11768 (N_11768,N_10779,N_10188);
xor U11769 (N_11769,N_10121,N_10661);
nand U11770 (N_11770,N_10992,N_10296);
nor U11771 (N_11771,N_10493,N_10651);
or U11772 (N_11772,N_10352,N_10367);
and U11773 (N_11773,N_10876,N_10393);
nor U11774 (N_11774,N_10260,N_10178);
or U11775 (N_11775,N_10472,N_10411);
nor U11776 (N_11776,N_10514,N_10106);
xnor U11777 (N_11777,N_10837,N_10964);
and U11778 (N_11778,N_10364,N_10814);
nand U11779 (N_11779,N_10500,N_10352);
nand U11780 (N_11780,N_10584,N_10794);
nor U11781 (N_11781,N_10249,N_10389);
nand U11782 (N_11782,N_10501,N_10020);
nand U11783 (N_11783,N_10658,N_10212);
or U11784 (N_11784,N_10822,N_10839);
nand U11785 (N_11785,N_10799,N_10683);
nor U11786 (N_11786,N_10963,N_10813);
xor U11787 (N_11787,N_10527,N_10429);
nor U11788 (N_11788,N_10531,N_10137);
and U11789 (N_11789,N_10791,N_10517);
nand U11790 (N_11790,N_10811,N_10555);
nand U11791 (N_11791,N_10379,N_10384);
nor U11792 (N_11792,N_10514,N_10978);
nor U11793 (N_11793,N_10942,N_10200);
xnor U11794 (N_11794,N_10554,N_10428);
or U11795 (N_11795,N_10207,N_10835);
and U11796 (N_11796,N_10951,N_10625);
nand U11797 (N_11797,N_10780,N_10954);
nand U11798 (N_11798,N_10947,N_10528);
or U11799 (N_11799,N_10848,N_10198);
nand U11800 (N_11800,N_10725,N_10273);
or U11801 (N_11801,N_10270,N_10471);
nand U11802 (N_11802,N_10321,N_10041);
and U11803 (N_11803,N_10447,N_10354);
and U11804 (N_11804,N_10445,N_10582);
xor U11805 (N_11805,N_10665,N_10990);
xnor U11806 (N_11806,N_10774,N_10795);
nand U11807 (N_11807,N_10154,N_10975);
or U11808 (N_11808,N_10313,N_10090);
xnor U11809 (N_11809,N_10265,N_10980);
or U11810 (N_11810,N_10627,N_10261);
and U11811 (N_11811,N_10497,N_10717);
and U11812 (N_11812,N_10374,N_10336);
or U11813 (N_11813,N_10493,N_10813);
nand U11814 (N_11814,N_10682,N_10049);
nand U11815 (N_11815,N_10880,N_10668);
or U11816 (N_11816,N_10556,N_10921);
xnor U11817 (N_11817,N_10925,N_10145);
xor U11818 (N_11818,N_10505,N_10794);
nand U11819 (N_11819,N_10014,N_10157);
xor U11820 (N_11820,N_10141,N_10132);
or U11821 (N_11821,N_10798,N_10815);
and U11822 (N_11822,N_10318,N_10560);
nand U11823 (N_11823,N_10945,N_10098);
xor U11824 (N_11824,N_10557,N_10753);
or U11825 (N_11825,N_10869,N_10365);
and U11826 (N_11826,N_10996,N_10294);
xnor U11827 (N_11827,N_10640,N_10612);
xnor U11828 (N_11828,N_10856,N_10423);
nor U11829 (N_11829,N_10284,N_10975);
or U11830 (N_11830,N_10614,N_10015);
xor U11831 (N_11831,N_10708,N_10511);
nand U11832 (N_11832,N_10508,N_10782);
xor U11833 (N_11833,N_10608,N_10511);
or U11834 (N_11834,N_10981,N_10292);
and U11835 (N_11835,N_10571,N_10619);
or U11836 (N_11836,N_10880,N_10245);
and U11837 (N_11837,N_10430,N_10399);
and U11838 (N_11838,N_10282,N_10626);
xnor U11839 (N_11839,N_10789,N_10744);
xnor U11840 (N_11840,N_10865,N_10050);
and U11841 (N_11841,N_10231,N_10684);
xor U11842 (N_11842,N_10548,N_10800);
xnor U11843 (N_11843,N_10121,N_10083);
or U11844 (N_11844,N_10752,N_10367);
or U11845 (N_11845,N_10670,N_10790);
and U11846 (N_11846,N_10626,N_10469);
nand U11847 (N_11847,N_10507,N_10769);
xor U11848 (N_11848,N_10242,N_10418);
nand U11849 (N_11849,N_10854,N_10073);
or U11850 (N_11850,N_10266,N_10911);
or U11851 (N_11851,N_10009,N_10471);
nand U11852 (N_11852,N_10098,N_10383);
or U11853 (N_11853,N_10783,N_10425);
nand U11854 (N_11854,N_10318,N_10978);
nor U11855 (N_11855,N_10829,N_10663);
and U11856 (N_11856,N_10746,N_10822);
nand U11857 (N_11857,N_10418,N_10910);
or U11858 (N_11858,N_10875,N_10940);
or U11859 (N_11859,N_10158,N_10783);
xor U11860 (N_11860,N_10818,N_10385);
nor U11861 (N_11861,N_10845,N_10836);
nor U11862 (N_11862,N_10638,N_10826);
nand U11863 (N_11863,N_10303,N_10456);
xnor U11864 (N_11864,N_10367,N_10414);
nor U11865 (N_11865,N_10601,N_10576);
and U11866 (N_11866,N_10737,N_10224);
nand U11867 (N_11867,N_10127,N_10622);
nor U11868 (N_11868,N_10261,N_10511);
and U11869 (N_11869,N_10597,N_10319);
xor U11870 (N_11870,N_10909,N_10941);
or U11871 (N_11871,N_10500,N_10882);
and U11872 (N_11872,N_10065,N_10239);
and U11873 (N_11873,N_10960,N_10981);
xnor U11874 (N_11874,N_10031,N_10474);
xor U11875 (N_11875,N_10414,N_10904);
nor U11876 (N_11876,N_10136,N_10063);
or U11877 (N_11877,N_10511,N_10564);
xnor U11878 (N_11878,N_10188,N_10892);
nor U11879 (N_11879,N_10625,N_10694);
and U11880 (N_11880,N_10563,N_10409);
nor U11881 (N_11881,N_10835,N_10631);
nand U11882 (N_11882,N_10160,N_10132);
nand U11883 (N_11883,N_10116,N_10151);
and U11884 (N_11884,N_10153,N_10698);
and U11885 (N_11885,N_10856,N_10951);
or U11886 (N_11886,N_10608,N_10636);
xnor U11887 (N_11887,N_10297,N_10718);
or U11888 (N_11888,N_10378,N_10928);
nor U11889 (N_11889,N_10096,N_10452);
nand U11890 (N_11890,N_10951,N_10010);
or U11891 (N_11891,N_10152,N_10161);
and U11892 (N_11892,N_10541,N_10147);
and U11893 (N_11893,N_10285,N_10974);
nor U11894 (N_11894,N_10563,N_10602);
or U11895 (N_11895,N_10749,N_10224);
xnor U11896 (N_11896,N_10600,N_10803);
or U11897 (N_11897,N_10450,N_10095);
nor U11898 (N_11898,N_10929,N_10268);
or U11899 (N_11899,N_10360,N_10988);
xor U11900 (N_11900,N_10276,N_10409);
xnor U11901 (N_11901,N_10710,N_10209);
and U11902 (N_11902,N_10260,N_10951);
and U11903 (N_11903,N_10042,N_10305);
nor U11904 (N_11904,N_10029,N_10691);
or U11905 (N_11905,N_10167,N_10480);
nand U11906 (N_11906,N_10043,N_10035);
nand U11907 (N_11907,N_10746,N_10520);
xnor U11908 (N_11908,N_10290,N_10936);
nand U11909 (N_11909,N_10643,N_10497);
nor U11910 (N_11910,N_10612,N_10916);
nand U11911 (N_11911,N_10738,N_10134);
nand U11912 (N_11912,N_10542,N_10692);
or U11913 (N_11913,N_10384,N_10132);
nand U11914 (N_11914,N_10819,N_10295);
xor U11915 (N_11915,N_10316,N_10191);
and U11916 (N_11916,N_10922,N_10072);
xnor U11917 (N_11917,N_10979,N_10686);
or U11918 (N_11918,N_10006,N_10566);
or U11919 (N_11919,N_10031,N_10078);
xnor U11920 (N_11920,N_10539,N_10554);
xnor U11921 (N_11921,N_10263,N_10912);
nor U11922 (N_11922,N_10696,N_10153);
nor U11923 (N_11923,N_10763,N_10044);
nand U11924 (N_11924,N_10659,N_10728);
xnor U11925 (N_11925,N_10937,N_10943);
xor U11926 (N_11926,N_10876,N_10506);
nand U11927 (N_11927,N_10660,N_10093);
and U11928 (N_11928,N_10778,N_10295);
and U11929 (N_11929,N_10130,N_10909);
nand U11930 (N_11930,N_10184,N_10595);
or U11931 (N_11931,N_10934,N_10763);
xnor U11932 (N_11932,N_10576,N_10826);
xor U11933 (N_11933,N_10573,N_10570);
and U11934 (N_11934,N_10262,N_10287);
xor U11935 (N_11935,N_10298,N_10628);
nand U11936 (N_11936,N_10331,N_10221);
xor U11937 (N_11937,N_10160,N_10584);
and U11938 (N_11938,N_10112,N_10023);
or U11939 (N_11939,N_10310,N_10390);
nand U11940 (N_11940,N_10075,N_10176);
or U11941 (N_11941,N_10843,N_10956);
nand U11942 (N_11942,N_10165,N_10056);
or U11943 (N_11943,N_10611,N_10627);
or U11944 (N_11944,N_10351,N_10919);
xnor U11945 (N_11945,N_10272,N_10119);
or U11946 (N_11946,N_10870,N_10459);
nand U11947 (N_11947,N_10063,N_10081);
or U11948 (N_11948,N_10101,N_10697);
and U11949 (N_11949,N_10306,N_10406);
xnor U11950 (N_11950,N_10962,N_10528);
nand U11951 (N_11951,N_10849,N_10531);
nor U11952 (N_11952,N_10884,N_10609);
or U11953 (N_11953,N_10296,N_10836);
and U11954 (N_11954,N_10363,N_10755);
nor U11955 (N_11955,N_10056,N_10274);
or U11956 (N_11956,N_10783,N_10542);
nor U11957 (N_11957,N_10566,N_10087);
and U11958 (N_11958,N_10384,N_10504);
and U11959 (N_11959,N_10251,N_10909);
and U11960 (N_11960,N_10231,N_10764);
or U11961 (N_11961,N_10076,N_10055);
xnor U11962 (N_11962,N_10896,N_10628);
xor U11963 (N_11963,N_10613,N_10263);
nand U11964 (N_11964,N_10128,N_10544);
nand U11965 (N_11965,N_10917,N_10257);
and U11966 (N_11966,N_10358,N_10769);
or U11967 (N_11967,N_10372,N_10900);
or U11968 (N_11968,N_10134,N_10564);
nor U11969 (N_11969,N_10195,N_10906);
nor U11970 (N_11970,N_10783,N_10983);
or U11971 (N_11971,N_10123,N_10469);
or U11972 (N_11972,N_10238,N_10977);
and U11973 (N_11973,N_10024,N_10091);
xnor U11974 (N_11974,N_10115,N_10177);
nor U11975 (N_11975,N_10741,N_10629);
nand U11976 (N_11976,N_10021,N_10875);
xnor U11977 (N_11977,N_10531,N_10662);
and U11978 (N_11978,N_10334,N_10953);
nor U11979 (N_11979,N_10122,N_10446);
nor U11980 (N_11980,N_10150,N_10518);
xnor U11981 (N_11981,N_10392,N_10616);
xnor U11982 (N_11982,N_10655,N_10137);
nand U11983 (N_11983,N_10251,N_10063);
and U11984 (N_11984,N_10515,N_10937);
nor U11985 (N_11985,N_10454,N_10074);
or U11986 (N_11986,N_10622,N_10602);
or U11987 (N_11987,N_10673,N_10162);
and U11988 (N_11988,N_10095,N_10387);
and U11989 (N_11989,N_10753,N_10924);
or U11990 (N_11990,N_10434,N_10398);
nor U11991 (N_11991,N_10055,N_10825);
nand U11992 (N_11992,N_10187,N_10011);
and U11993 (N_11993,N_10096,N_10028);
nand U11994 (N_11994,N_10865,N_10876);
nand U11995 (N_11995,N_10986,N_10386);
xor U11996 (N_11996,N_10835,N_10796);
nand U11997 (N_11997,N_10107,N_10002);
or U11998 (N_11998,N_10332,N_10180);
and U11999 (N_11999,N_10193,N_10055);
nand U12000 (N_12000,N_11883,N_11499);
nand U12001 (N_12001,N_11031,N_11486);
and U12002 (N_12002,N_11145,N_11452);
nand U12003 (N_12003,N_11964,N_11591);
nor U12004 (N_12004,N_11411,N_11703);
nor U12005 (N_12005,N_11331,N_11852);
nand U12006 (N_12006,N_11969,N_11825);
or U12007 (N_12007,N_11754,N_11455);
nand U12008 (N_12008,N_11888,N_11010);
or U12009 (N_12009,N_11677,N_11404);
or U12010 (N_12010,N_11831,N_11971);
or U12011 (N_12011,N_11718,N_11166);
and U12012 (N_12012,N_11976,N_11779);
or U12013 (N_12013,N_11472,N_11725);
nand U12014 (N_12014,N_11350,N_11337);
or U12015 (N_12015,N_11817,N_11321);
nor U12016 (N_12016,N_11663,N_11657);
xnor U12017 (N_12017,N_11672,N_11605);
nor U12018 (N_12018,N_11340,N_11383);
and U12019 (N_12019,N_11083,N_11592);
and U12020 (N_12020,N_11866,N_11271);
and U12021 (N_12021,N_11051,N_11181);
nor U12022 (N_12022,N_11930,N_11717);
nor U12023 (N_12023,N_11542,N_11105);
and U12024 (N_12024,N_11550,N_11264);
xnor U12025 (N_12025,N_11508,N_11222);
xor U12026 (N_12026,N_11034,N_11562);
nor U12027 (N_12027,N_11483,N_11143);
nand U12028 (N_12028,N_11133,N_11458);
nor U12029 (N_12029,N_11644,N_11116);
and U12030 (N_12030,N_11630,N_11967);
or U12031 (N_12031,N_11119,N_11233);
nor U12032 (N_12032,N_11566,N_11739);
and U12033 (N_12033,N_11152,N_11648);
or U12034 (N_12034,N_11540,N_11281);
and U12035 (N_12035,N_11859,N_11001);
and U12036 (N_12036,N_11393,N_11307);
xor U12037 (N_12037,N_11737,N_11865);
nand U12038 (N_12038,N_11423,N_11492);
nand U12039 (N_12039,N_11583,N_11033);
or U12040 (N_12040,N_11706,N_11169);
nand U12041 (N_12041,N_11952,N_11005);
and U12042 (N_12042,N_11374,N_11827);
nand U12043 (N_12043,N_11646,N_11114);
nor U12044 (N_12044,N_11256,N_11816);
xor U12045 (N_12045,N_11137,N_11571);
nand U12046 (N_12046,N_11667,N_11514);
or U12047 (N_12047,N_11359,N_11622);
or U12048 (N_12048,N_11266,N_11398);
and U12049 (N_12049,N_11498,N_11786);
nor U12050 (N_12050,N_11532,N_11559);
xor U12051 (N_12051,N_11178,N_11280);
and U12052 (N_12052,N_11796,N_11288);
xnor U12053 (N_12053,N_11387,N_11129);
or U12054 (N_12054,N_11733,N_11229);
or U12055 (N_12055,N_11585,N_11531);
nand U12056 (N_12056,N_11135,N_11056);
nor U12057 (N_12057,N_11029,N_11927);
nor U12058 (N_12058,N_11028,N_11875);
nand U12059 (N_12059,N_11521,N_11830);
xor U12060 (N_12060,N_11651,N_11579);
nor U12061 (N_12061,N_11656,N_11209);
xnor U12062 (N_12062,N_11738,N_11343);
and U12063 (N_12063,N_11985,N_11197);
and U12064 (N_12064,N_11287,N_11609);
nand U12065 (N_12065,N_11090,N_11120);
and U12066 (N_12066,N_11047,N_11035);
or U12067 (N_12067,N_11496,N_11490);
nand U12068 (N_12068,N_11019,N_11603);
nor U12069 (N_12069,N_11075,N_11467);
and U12070 (N_12070,N_11273,N_11303);
nor U12071 (N_12071,N_11749,N_11970);
and U12072 (N_12072,N_11654,N_11440);
xnor U12073 (N_12073,N_11153,N_11957);
xnor U12074 (N_12074,N_11727,N_11743);
nand U12075 (N_12075,N_11040,N_11820);
nor U12076 (N_12076,N_11054,N_11772);
xor U12077 (N_12077,N_11876,N_11442);
xnor U12078 (N_12078,N_11501,N_11430);
or U12079 (N_12079,N_11134,N_11803);
nand U12080 (N_12080,N_11941,N_11977);
or U12081 (N_12081,N_11915,N_11728);
nor U12082 (N_12082,N_11380,N_11860);
or U12083 (N_12083,N_11513,N_11841);
or U12084 (N_12084,N_11889,N_11077);
nor U12085 (N_12085,N_11230,N_11880);
nand U12086 (N_12086,N_11024,N_11372);
or U12087 (N_12087,N_11184,N_11381);
nor U12088 (N_12088,N_11881,N_11551);
and U12089 (N_12089,N_11580,N_11587);
nand U12090 (N_12090,N_11260,N_11155);
and U12091 (N_12091,N_11891,N_11265);
nor U12092 (N_12092,N_11910,N_11601);
xnor U12093 (N_12093,N_11182,N_11569);
xor U12094 (N_12094,N_11436,N_11267);
xor U12095 (N_12095,N_11544,N_11529);
or U12096 (N_12096,N_11702,N_11638);
nor U12097 (N_12097,N_11762,N_11548);
xnor U12098 (N_12098,N_11300,N_11424);
nor U12099 (N_12099,N_11560,N_11225);
nand U12100 (N_12100,N_11022,N_11946);
nand U12101 (N_12101,N_11636,N_11805);
and U12102 (N_12102,N_11572,N_11610);
nor U12103 (N_12103,N_11854,N_11568);
xnor U12104 (N_12104,N_11797,N_11641);
nor U12105 (N_12105,N_11744,N_11892);
and U12106 (N_12106,N_11216,N_11798);
xnor U12107 (N_12107,N_11647,N_11355);
nor U12108 (N_12108,N_11917,N_11819);
and U12109 (N_12109,N_11305,N_11027);
nor U12110 (N_12110,N_11956,N_11959);
or U12111 (N_12111,N_11773,N_11503);
or U12112 (N_12112,N_11870,N_11414);
nand U12113 (N_12113,N_11050,N_11484);
nor U12114 (N_12114,N_11058,N_11761);
nand U12115 (N_12115,N_11422,N_11962);
and U12116 (N_12116,N_11417,N_11682);
xnor U12117 (N_12117,N_11815,N_11687);
nand U12118 (N_12118,N_11136,N_11722);
nand U12119 (N_12119,N_11185,N_11335);
or U12120 (N_12120,N_11386,N_11533);
and U12121 (N_12121,N_11038,N_11071);
or U12122 (N_12122,N_11555,N_11205);
and U12123 (N_12123,N_11148,N_11836);
or U12124 (N_12124,N_11893,N_11319);
xor U12125 (N_12125,N_11026,N_11212);
or U12126 (N_12126,N_11416,N_11839);
xor U12127 (N_12127,N_11103,N_11294);
nor U12128 (N_12128,N_11669,N_11057);
nor U12129 (N_12129,N_11905,N_11629);
or U12130 (N_12130,N_11925,N_11916);
xnor U12131 (N_12131,N_11724,N_11624);
xnor U12132 (N_12132,N_11074,N_11278);
nor U12133 (N_12133,N_11125,N_11705);
nor U12134 (N_12134,N_11901,N_11558);
nand U12135 (N_12135,N_11882,N_11988);
or U12136 (N_12136,N_11258,N_11245);
and U12137 (N_12137,N_11014,N_11661);
or U12138 (N_12138,N_11244,N_11284);
xor U12139 (N_12139,N_11409,N_11588);
and U12140 (N_12140,N_11076,N_11365);
nor U12141 (N_12141,N_11360,N_11344);
nand U12142 (N_12142,N_11060,N_11862);
nor U12143 (N_12143,N_11481,N_11736);
xnor U12144 (N_12144,N_11223,N_11361);
xor U12145 (N_12145,N_11561,N_11594);
xor U12146 (N_12146,N_11263,N_11784);
xnor U12147 (N_12147,N_11429,N_11131);
nor U12148 (N_12148,N_11945,N_11720);
nand U12149 (N_12149,N_11109,N_11793);
nand U12150 (N_12150,N_11085,N_11206);
nor U12151 (N_12151,N_11584,N_11975);
xor U12152 (N_12152,N_11752,N_11457);
xor U12153 (N_12153,N_11164,N_11375);
xnor U12154 (N_12154,N_11464,N_11237);
xnor U12155 (N_12155,N_11673,N_11810);
nand U12156 (N_12156,N_11502,N_11494);
or U12157 (N_12157,N_11576,N_11991);
nor U12158 (N_12158,N_11312,N_11402);
and U12159 (N_12159,N_11989,N_11998);
xnor U12160 (N_12160,N_11236,N_11138);
and U12161 (N_12161,N_11747,N_11140);
nor U12162 (N_12162,N_11482,N_11275);
xnor U12163 (N_12163,N_11593,N_11239);
xnor U12164 (N_12164,N_11723,N_11879);
nor U12165 (N_12165,N_11814,N_11167);
nor U12166 (N_12166,N_11834,N_11929);
xor U12167 (N_12167,N_11535,N_11208);
nor U12168 (N_12168,N_11388,N_11589);
nand U12169 (N_12169,N_11771,N_11403);
nand U12170 (N_12170,N_11689,N_11397);
xnor U12171 (N_12171,N_11679,N_11290);
and U12172 (N_12172,N_11221,N_11084);
nand U12173 (N_12173,N_11401,N_11680);
xor U12174 (N_12174,N_11463,N_11701);
xnor U12175 (N_12175,N_11867,N_11317);
nor U12176 (N_12176,N_11745,N_11384);
and U12177 (N_12177,N_11141,N_11575);
or U12178 (N_12178,N_11768,N_11520);
nand U12179 (N_12179,N_11684,N_11213);
nand U12180 (N_12180,N_11011,N_11619);
nand U12181 (N_12181,N_11104,N_11983);
nor U12182 (N_12182,N_11899,N_11269);
nand U12183 (N_12183,N_11537,N_11246);
and U12184 (N_12184,N_11394,N_11543);
nand U12185 (N_12185,N_11459,N_11844);
nand U12186 (N_12186,N_11923,N_11352);
and U12187 (N_12187,N_11306,N_11719);
nand U12188 (N_12188,N_11214,N_11470);
and U12189 (N_12189,N_11309,N_11110);
nor U12190 (N_12190,N_11694,N_11695);
and U12191 (N_12191,N_11362,N_11163);
xor U12192 (N_12192,N_11347,N_11730);
nor U12193 (N_12193,N_11480,N_11396);
and U12194 (N_12194,N_11091,N_11864);
nand U12195 (N_12195,N_11783,N_11493);
nand U12196 (N_12196,N_11378,N_11690);
nor U12197 (N_12197,N_11190,N_11323);
and U12198 (N_12198,N_11293,N_11504);
or U12199 (N_12199,N_11189,N_11757);
xor U12200 (N_12200,N_11444,N_11358);
xor U12201 (N_12201,N_11982,N_11021);
and U12202 (N_12202,N_11960,N_11226);
xor U12203 (N_12203,N_11794,N_11753);
or U12204 (N_12204,N_11241,N_11848);
xor U12205 (N_12205,N_11080,N_11299);
and U12206 (N_12206,N_11519,N_11295);
and U12207 (N_12207,N_11150,N_11740);
xor U12208 (N_12208,N_11356,N_11215);
nand U12209 (N_12209,N_11978,N_11391);
and U12210 (N_12210,N_11688,N_11894);
xnor U12211 (N_12211,N_11660,N_11811);
xnor U12212 (N_12212,N_11055,N_11297);
nor U12213 (N_12213,N_11774,N_11869);
xnor U12214 (N_12214,N_11025,N_11611);
or U12215 (N_12215,N_11926,N_11564);
nor U12216 (N_12216,N_11523,N_11554);
nor U12217 (N_12217,N_11479,N_11721);
nor U12218 (N_12218,N_11577,N_11782);
and U12219 (N_12219,N_11495,N_11913);
xor U12220 (N_12220,N_11345,N_11389);
and U12221 (N_12221,N_11686,N_11052);
nor U12222 (N_12222,N_11268,N_11835);
or U12223 (N_12223,N_11900,N_11346);
xnor U12224 (N_12224,N_11064,N_11990);
xnor U12225 (N_12225,N_11943,N_11107);
nor U12226 (N_12226,N_11565,N_11325);
xor U12227 (N_12227,N_11813,N_11234);
and U12228 (N_12228,N_11668,N_11262);
nand U12229 (N_12229,N_11139,N_11043);
nand U12230 (N_12230,N_11581,N_11068);
xor U12231 (N_12231,N_11007,N_11364);
nand U12232 (N_12232,N_11949,N_11853);
and U12233 (N_12233,N_11008,N_11183);
or U12234 (N_12234,N_11311,N_11858);
nor U12235 (N_12235,N_11981,N_11921);
nor U12236 (N_12236,N_11338,N_11549);
xnor U12237 (N_12237,N_11456,N_11600);
and U12238 (N_12238,N_11354,N_11478);
nor U12239 (N_12239,N_11951,N_11407);
nor U12240 (N_12240,N_11062,N_11106);
or U12241 (N_12241,N_11902,N_11015);
nor U12242 (N_12242,N_11912,N_11868);
nand U12243 (N_12243,N_11332,N_11965);
or U12244 (N_12244,N_11098,N_11557);
xnor U12245 (N_12245,N_11086,N_11691);
nor U12246 (N_12246,N_11218,N_11210);
nand U12247 (N_12247,N_11979,N_11821);
nor U12248 (N_12248,N_11349,N_11063);
nor U12249 (N_12249,N_11872,N_11897);
nand U12250 (N_12250,N_11995,N_11170);
and U12251 (N_12251,N_11539,N_11379);
and U12252 (N_12252,N_11896,N_11732);
nor U12253 (N_12253,N_11441,N_11826);
nand U12254 (N_12254,N_11298,N_11069);
or U12255 (N_12255,N_11595,N_11530);
nor U12256 (N_12256,N_11645,N_11147);
xor U12257 (N_12257,N_11002,N_11670);
xnor U12258 (N_12258,N_11639,N_11200);
nor U12259 (N_12259,N_11289,N_11809);
and U12260 (N_12260,N_11607,N_11987);
nand U12261 (N_12261,N_11469,N_11751);
or U12262 (N_12262,N_11179,N_11746);
nor U12263 (N_12263,N_11671,N_11474);
or U12264 (N_12264,N_11612,N_11996);
nor U12265 (N_12265,N_11685,N_11427);
xor U12266 (N_12266,N_11412,N_11270);
and U12267 (N_12267,N_11111,N_11192);
nand U12268 (N_12268,N_11997,N_11828);
and U12269 (N_12269,N_11369,N_11257);
nand U12270 (N_12270,N_11570,N_11808);
and U12271 (N_12271,N_11909,N_11681);
nand U12272 (N_12272,N_11666,N_11082);
or U12273 (N_12273,N_11092,N_11528);
nand U12274 (N_12274,N_11408,N_11065);
or U12275 (N_12275,N_11276,N_11177);
nor U12276 (N_12276,N_11445,N_11204);
nor U12277 (N_12277,N_11122,N_11908);
and U12278 (N_12278,N_11487,N_11596);
or U12279 (N_12279,N_11541,N_11628);
and U12280 (N_12280,N_11778,N_11972);
nor U12281 (N_12281,N_11861,N_11342);
xnor U12282 (N_12282,N_11196,N_11121);
nor U12283 (N_12283,N_11446,N_11709);
and U12284 (N_12284,N_11253,N_11400);
nor U12285 (N_12285,N_11093,N_11371);
nor U12286 (N_12286,N_11497,N_11986);
nand U12287 (N_12287,N_11180,N_11471);
xnor U12288 (N_12288,N_11635,N_11302);
nand U12289 (N_12289,N_11567,N_11741);
or U12290 (N_12290,N_11842,N_11696);
nor U12291 (N_12291,N_11327,N_11715);
or U12292 (N_12292,N_11078,N_11785);
nor U12293 (N_12293,N_11066,N_11443);
nor U12294 (N_12294,N_11451,N_11904);
or U12295 (N_12295,N_11895,N_11553);
nand U12296 (N_12296,N_11873,N_11525);
and U12297 (N_12297,N_11020,N_11755);
nand U12298 (N_12298,N_11961,N_11462);
and U12299 (N_12299,N_11582,N_11032);
or U12300 (N_12300,N_11632,N_11087);
or U12301 (N_12301,N_11454,N_11292);
xor U12302 (N_12302,N_11348,N_11716);
or U12303 (N_12303,N_11489,N_11079);
and U12304 (N_12304,N_11162,N_11194);
nand U12305 (N_12305,N_11439,N_11413);
and U12306 (N_12306,N_11099,N_11248);
or U12307 (N_12307,N_11992,N_11791);
nor U12308 (N_12308,N_11748,N_11833);
and U12309 (N_12309,N_11220,N_11676);
nor U12310 (N_12310,N_11198,N_11334);
xor U12311 (N_12311,N_11390,N_11088);
nand U12312 (N_12312,N_11320,N_11665);
and U12313 (N_12313,N_11505,N_11186);
nor U12314 (N_12314,N_11818,N_11219);
xor U12315 (N_12315,N_11405,N_11799);
nand U12316 (N_12316,N_11634,N_11763);
or U12317 (N_12317,N_11420,N_11448);
nand U12318 (N_12318,N_11775,N_11048);
nand U12319 (N_12319,N_11759,N_11285);
nor U12320 (N_12320,N_11252,N_11769);
or U12321 (N_12321,N_11855,N_11507);
xor U12322 (N_12322,N_11385,N_11787);
xor U12323 (N_12323,N_11061,N_11536);
nand U12324 (N_12324,N_11602,N_11884);
or U12325 (N_12325,N_11795,N_11261);
xnor U12326 (N_12326,N_11527,N_11937);
nand U12327 (N_12327,N_11151,N_11758);
or U12328 (N_12328,N_11518,N_11620);
and U12329 (N_12329,N_11765,N_11675);
and U12330 (N_12330,N_11806,N_11538);
nor U12331 (N_12331,N_11942,N_11291);
or U12332 (N_12332,N_11512,N_11286);
nor U12333 (N_12333,N_11046,N_11447);
or U12334 (N_12334,N_11449,N_11655);
and U12335 (N_12335,N_11004,N_11191);
nand U12336 (N_12336,N_11142,N_11108);
xor U12337 (N_12337,N_11802,N_11936);
or U12338 (N_12338,N_11041,N_11053);
or U12339 (N_12339,N_11726,N_11800);
and U12340 (N_12340,N_11829,N_11003);
xor U12341 (N_12341,N_11914,N_11789);
or U12342 (N_12342,N_11938,N_11130);
xnor U12343 (N_12343,N_11161,N_11973);
nand U12344 (N_12344,N_11376,N_11419);
and U12345 (N_12345,N_11433,N_11096);
xnor U12346 (N_12346,N_11249,N_11154);
xnor U12347 (N_12347,N_11175,N_11247);
xnor U12348 (N_12348,N_11734,N_11918);
xnor U12349 (N_12349,N_11511,N_11195);
nand U12350 (N_12350,N_11188,N_11059);
nor U12351 (N_12351,N_11425,N_11102);
xnor U12352 (N_12352,N_11878,N_11199);
or U12353 (N_12353,N_11940,N_11168);
and U12354 (N_12354,N_11203,N_11165);
or U12355 (N_12355,N_11009,N_11933);
nor U12356 (N_12356,N_11729,N_11468);
nand U12357 (N_12357,N_11613,N_11708);
nand U12358 (N_12358,N_11640,N_11710);
or U12359 (N_12359,N_11231,N_11906);
and U12360 (N_12360,N_11903,N_11823);
xor U12361 (N_12361,N_11950,N_11845);
nor U12362 (N_12362,N_11159,N_11556);
and U12363 (N_12363,N_11012,N_11112);
nor U12364 (N_12364,N_11650,N_11857);
and U12365 (N_12365,N_11693,N_11172);
and U12366 (N_12366,N_11958,N_11993);
xnor U12367 (N_12367,N_11030,N_11790);
and U12368 (N_12368,N_11627,N_11118);
nand U12369 (N_12369,N_11485,N_11526);
nand U12370 (N_12370,N_11313,N_11849);
nor U12371 (N_12371,N_11308,N_11597);
and U12372 (N_12372,N_11767,N_11392);
and U12373 (N_12373,N_11649,N_11461);
nand U12374 (N_12374,N_11115,N_11211);
or U12375 (N_12375,N_11368,N_11545);
or U12376 (N_12376,N_11421,N_11149);
xor U12377 (N_12377,N_11932,N_11843);
nand U12378 (N_12378,N_11201,N_11517);
xnor U12379 (N_12379,N_11310,N_11089);
and U12380 (N_12380,N_11984,N_11316);
and U12381 (N_12381,N_11251,N_11399);
nand U12382 (N_12382,N_11434,N_11804);
nand U12383 (N_12383,N_11473,N_11522);
nor U12384 (N_12384,N_11546,N_11766);
xnor U12385 (N_12385,N_11006,N_11304);
and U12386 (N_12386,N_11101,N_11227);
nand U12387 (N_12387,N_11922,N_11621);
xor U12388 (N_12388,N_11377,N_11847);
and U12389 (N_12389,N_11160,N_11944);
and U12390 (N_12390,N_11658,N_11370);
or U12391 (N_12391,N_11509,N_11238);
and U12392 (N_12392,N_11367,N_11885);
or U12393 (N_12393,N_11081,N_11711);
nor U12394 (N_12394,N_11477,N_11157);
or U12395 (N_12395,N_11935,N_11919);
or U12396 (N_12396,N_11637,N_11626);
nand U12397 (N_12397,N_11678,N_11840);
xor U12398 (N_12398,N_11770,N_11475);
xnor U12399 (N_12399,N_11506,N_11254);
nand U12400 (N_12400,N_11272,N_11333);
or U12401 (N_12401,N_11623,N_11018);
nand U12402 (N_12402,N_11948,N_11874);
xor U12403 (N_12403,N_11049,N_11516);
and U12404 (N_12404,N_11939,N_11491);
xor U12405 (N_12405,N_11132,N_11617);
or U12406 (N_12406,N_11760,N_11097);
and U12407 (N_12407,N_11590,N_11598);
nor U12408 (N_12408,N_11683,N_11171);
and U12409 (N_12409,N_11563,N_11822);
xor U12410 (N_12410,N_11837,N_11606);
and U12411 (N_12411,N_11395,N_11954);
nand U12412 (N_12412,N_11714,N_11341);
and U12413 (N_12413,N_11037,N_11756);
and U12414 (N_12414,N_11232,N_11336);
and U12415 (N_12415,N_11277,N_11807);
and U12416 (N_12416,N_11931,N_11328);
nand U12417 (N_12417,N_11039,N_11968);
or U12418 (N_12418,N_11534,N_11788);
nor U12419 (N_12419,N_11146,N_11731);
xor U12420 (N_12420,N_11406,N_11966);
and U12421 (N_12421,N_11604,N_11144);
and U12422 (N_12422,N_11699,N_11016);
xor U12423 (N_12423,N_11450,N_11460);
and U12424 (N_12424,N_11315,N_11735);
or U12425 (N_12425,N_11123,N_11887);
and U12426 (N_12426,N_11776,N_11780);
xor U12427 (N_12427,N_11279,N_11642);
xor U12428 (N_12428,N_11283,N_11633);
nand U12429 (N_12429,N_11073,N_11924);
or U12430 (N_12430,N_11124,N_11934);
xnor U12431 (N_12431,N_11158,N_11242);
nand U12432 (N_12432,N_11070,N_11428);
and U12433 (N_12433,N_11067,N_11578);
nor U12434 (N_12434,N_11777,N_11326);
nand U12435 (N_12435,N_11353,N_11044);
nor U12436 (N_12436,N_11095,N_11500);
and U12437 (N_12437,N_11653,N_11692);
nor U12438 (N_12438,N_11643,N_11000);
or U12439 (N_12439,N_11697,N_11907);
and U12440 (N_12440,N_11547,N_11156);
nand U12441 (N_12441,N_11351,N_11259);
xor U12442 (N_12442,N_11674,N_11928);
nor U12443 (N_12443,N_11126,N_11339);
nor U12444 (N_12444,N_11042,N_11838);
or U12445 (N_12445,N_11599,N_11324);
and U12446 (N_12446,N_11296,N_11476);
nand U12447 (N_12447,N_11574,N_11255);
and U12448 (N_12448,N_11877,N_11432);
or U12449 (N_12449,N_11850,N_11330);
and U12450 (N_12450,N_11357,N_11127);
or U12451 (N_12451,N_11824,N_11437);
nand U12452 (N_12452,N_11953,N_11366);
or U12453 (N_12453,N_11488,N_11466);
nor U12454 (N_12454,N_11573,N_11128);
and U12455 (N_12455,N_11217,N_11453);
xor U12456 (N_12456,N_11250,N_11781);
nor U12457 (N_12457,N_11329,N_11618);
and U12458 (N_12458,N_11426,N_11045);
nand U12459 (N_12459,N_11898,N_11801);
nand U12460 (N_12460,N_11524,N_11890);
xnor U12461 (N_12461,N_11418,N_11193);
nand U12462 (N_12462,N_11174,N_11431);
or U12463 (N_12463,N_11980,N_11955);
nand U12464 (N_12464,N_11886,N_11552);
nor U12465 (N_12465,N_11631,N_11282);
or U12466 (N_12466,N_11713,N_11625);
nand U12467 (N_12467,N_11100,N_11318);
xor U12468 (N_12468,N_11871,N_11920);
nor U12469 (N_12469,N_11832,N_11363);
and U12470 (N_12470,N_11228,N_11187);
nand U12471 (N_12471,N_11072,N_11224);
nand U12472 (N_12472,N_11911,N_11415);
nand U12473 (N_12473,N_11176,N_11846);
nand U12474 (N_12474,N_11017,N_11202);
nor U12475 (N_12475,N_11614,N_11207);
or U12476 (N_12476,N_11750,N_11707);
or U12477 (N_12477,N_11994,N_11792);
and U12478 (N_12478,N_11036,N_11947);
nand U12479 (N_12479,N_11382,N_11117);
and U12480 (N_12480,N_11515,N_11438);
and U12481 (N_12481,N_11240,N_11742);
nor U12482 (N_12482,N_11023,N_11856);
nor U12483 (N_12483,N_11322,N_11664);
nand U12484 (N_12484,N_11235,N_11373);
xor U12485 (N_12485,N_11999,N_11704);
xor U12486 (N_12486,N_11863,N_11616);
xnor U12487 (N_12487,N_11652,N_11465);
or U12488 (N_12488,N_11510,N_11698);
and U12489 (N_12489,N_11410,N_11963);
or U12490 (N_12490,N_11608,N_11013);
nand U12491 (N_12491,N_11094,N_11851);
nand U12492 (N_12492,N_11243,N_11974);
xor U12493 (N_12493,N_11274,N_11435);
or U12494 (N_12494,N_11764,N_11113);
nand U12495 (N_12495,N_11314,N_11659);
nand U12496 (N_12496,N_11615,N_11586);
xor U12497 (N_12497,N_11812,N_11662);
or U12498 (N_12498,N_11712,N_11173);
nand U12499 (N_12499,N_11700,N_11301);
and U12500 (N_12500,N_11242,N_11849);
and U12501 (N_12501,N_11774,N_11427);
and U12502 (N_12502,N_11806,N_11234);
nand U12503 (N_12503,N_11767,N_11309);
nor U12504 (N_12504,N_11897,N_11881);
or U12505 (N_12505,N_11992,N_11637);
nand U12506 (N_12506,N_11356,N_11401);
nand U12507 (N_12507,N_11902,N_11033);
nand U12508 (N_12508,N_11288,N_11641);
or U12509 (N_12509,N_11590,N_11011);
xnor U12510 (N_12510,N_11011,N_11239);
xor U12511 (N_12511,N_11525,N_11810);
and U12512 (N_12512,N_11668,N_11917);
and U12513 (N_12513,N_11863,N_11821);
nor U12514 (N_12514,N_11739,N_11061);
nand U12515 (N_12515,N_11407,N_11102);
xor U12516 (N_12516,N_11785,N_11208);
nor U12517 (N_12517,N_11183,N_11728);
or U12518 (N_12518,N_11239,N_11272);
or U12519 (N_12519,N_11216,N_11689);
nand U12520 (N_12520,N_11513,N_11492);
or U12521 (N_12521,N_11912,N_11580);
nand U12522 (N_12522,N_11211,N_11646);
or U12523 (N_12523,N_11531,N_11902);
xor U12524 (N_12524,N_11541,N_11287);
nor U12525 (N_12525,N_11204,N_11554);
nor U12526 (N_12526,N_11724,N_11874);
nor U12527 (N_12527,N_11301,N_11076);
or U12528 (N_12528,N_11165,N_11116);
or U12529 (N_12529,N_11388,N_11082);
xor U12530 (N_12530,N_11937,N_11726);
xnor U12531 (N_12531,N_11622,N_11358);
nand U12532 (N_12532,N_11933,N_11118);
nor U12533 (N_12533,N_11048,N_11879);
and U12534 (N_12534,N_11459,N_11863);
or U12535 (N_12535,N_11271,N_11212);
or U12536 (N_12536,N_11245,N_11754);
nor U12537 (N_12537,N_11047,N_11725);
nor U12538 (N_12538,N_11265,N_11422);
or U12539 (N_12539,N_11273,N_11117);
xnor U12540 (N_12540,N_11896,N_11362);
and U12541 (N_12541,N_11064,N_11989);
nor U12542 (N_12542,N_11429,N_11928);
nor U12543 (N_12543,N_11572,N_11260);
nand U12544 (N_12544,N_11271,N_11566);
nand U12545 (N_12545,N_11196,N_11328);
or U12546 (N_12546,N_11800,N_11794);
or U12547 (N_12547,N_11887,N_11450);
or U12548 (N_12548,N_11801,N_11559);
xnor U12549 (N_12549,N_11095,N_11327);
and U12550 (N_12550,N_11775,N_11350);
and U12551 (N_12551,N_11189,N_11955);
nand U12552 (N_12552,N_11916,N_11904);
and U12553 (N_12553,N_11692,N_11951);
xnor U12554 (N_12554,N_11297,N_11983);
or U12555 (N_12555,N_11344,N_11522);
and U12556 (N_12556,N_11970,N_11212);
or U12557 (N_12557,N_11719,N_11759);
and U12558 (N_12558,N_11587,N_11750);
nand U12559 (N_12559,N_11619,N_11198);
or U12560 (N_12560,N_11092,N_11478);
xor U12561 (N_12561,N_11850,N_11159);
nand U12562 (N_12562,N_11532,N_11312);
nor U12563 (N_12563,N_11985,N_11869);
nor U12564 (N_12564,N_11514,N_11367);
xor U12565 (N_12565,N_11267,N_11215);
or U12566 (N_12566,N_11877,N_11611);
xor U12567 (N_12567,N_11887,N_11463);
or U12568 (N_12568,N_11119,N_11616);
and U12569 (N_12569,N_11740,N_11089);
nand U12570 (N_12570,N_11094,N_11537);
or U12571 (N_12571,N_11130,N_11341);
nor U12572 (N_12572,N_11096,N_11322);
or U12573 (N_12573,N_11951,N_11071);
xor U12574 (N_12574,N_11624,N_11953);
nand U12575 (N_12575,N_11899,N_11878);
xnor U12576 (N_12576,N_11842,N_11051);
nand U12577 (N_12577,N_11401,N_11854);
nand U12578 (N_12578,N_11926,N_11076);
nor U12579 (N_12579,N_11807,N_11211);
nor U12580 (N_12580,N_11262,N_11032);
or U12581 (N_12581,N_11489,N_11383);
nand U12582 (N_12582,N_11079,N_11024);
and U12583 (N_12583,N_11660,N_11541);
xnor U12584 (N_12584,N_11644,N_11926);
and U12585 (N_12585,N_11725,N_11710);
and U12586 (N_12586,N_11714,N_11871);
nor U12587 (N_12587,N_11236,N_11842);
nor U12588 (N_12588,N_11766,N_11512);
and U12589 (N_12589,N_11337,N_11805);
nand U12590 (N_12590,N_11888,N_11626);
xor U12591 (N_12591,N_11213,N_11195);
xnor U12592 (N_12592,N_11108,N_11445);
nand U12593 (N_12593,N_11355,N_11430);
or U12594 (N_12594,N_11214,N_11991);
nand U12595 (N_12595,N_11526,N_11098);
xor U12596 (N_12596,N_11295,N_11391);
or U12597 (N_12597,N_11029,N_11235);
or U12598 (N_12598,N_11610,N_11571);
and U12599 (N_12599,N_11946,N_11506);
nor U12600 (N_12600,N_11102,N_11513);
xor U12601 (N_12601,N_11640,N_11178);
nor U12602 (N_12602,N_11534,N_11898);
nand U12603 (N_12603,N_11974,N_11633);
and U12604 (N_12604,N_11400,N_11823);
xnor U12605 (N_12605,N_11980,N_11682);
nor U12606 (N_12606,N_11394,N_11829);
and U12607 (N_12607,N_11754,N_11392);
nand U12608 (N_12608,N_11504,N_11429);
or U12609 (N_12609,N_11126,N_11446);
nand U12610 (N_12610,N_11740,N_11363);
and U12611 (N_12611,N_11820,N_11252);
and U12612 (N_12612,N_11339,N_11670);
nor U12613 (N_12613,N_11889,N_11255);
or U12614 (N_12614,N_11605,N_11623);
or U12615 (N_12615,N_11908,N_11669);
nand U12616 (N_12616,N_11882,N_11543);
and U12617 (N_12617,N_11779,N_11382);
and U12618 (N_12618,N_11629,N_11928);
nand U12619 (N_12619,N_11508,N_11432);
nor U12620 (N_12620,N_11479,N_11942);
xnor U12621 (N_12621,N_11723,N_11055);
nor U12622 (N_12622,N_11787,N_11330);
and U12623 (N_12623,N_11786,N_11539);
or U12624 (N_12624,N_11802,N_11017);
or U12625 (N_12625,N_11436,N_11531);
nor U12626 (N_12626,N_11224,N_11296);
and U12627 (N_12627,N_11874,N_11158);
and U12628 (N_12628,N_11673,N_11069);
nor U12629 (N_12629,N_11182,N_11516);
or U12630 (N_12630,N_11510,N_11922);
nand U12631 (N_12631,N_11768,N_11703);
nor U12632 (N_12632,N_11612,N_11445);
nand U12633 (N_12633,N_11336,N_11909);
nor U12634 (N_12634,N_11209,N_11017);
or U12635 (N_12635,N_11400,N_11190);
and U12636 (N_12636,N_11453,N_11900);
nor U12637 (N_12637,N_11740,N_11781);
and U12638 (N_12638,N_11569,N_11774);
nor U12639 (N_12639,N_11990,N_11155);
nand U12640 (N_12640,N_11016,N_11100);
nand U12641 (N_12641,N_11876,N_11747);
and U12642 (N_12642,N_11994,N_11942);
nand U12643 (N_12643,N_11659,N_11061);
and U12644 (N_12644,N_11276,N_11450);
and U12645 (N_12645,N_11257,N_11150);
xor U12646 (N_12646,N_11447,N_11510);
or U12647 (N_12647,N_11792,N_11294);
xnor U12648 (N_12648,N_11393,N_11024);
or U12649 (N_12649,N_11922,N_11631);
nor U12650 (N_12650,N_11497,N_11552);
nor U12651 (N_12651,N_11678,N_11833);
or U12652 (N_12652,N_11363,N_11400);
and U12653 (N_12653,N_11131,N_11077);
xnor U12654 (N_12654,N_11172,N_11554);
and U12655 (N_12655,N_11797,N_11522);
or U12656 (N_12656,N_11823,N_11442);
nand U12657 (N_12657,N_11644,N_11862);
xor U12658 (N_12658,N_11164,N_11539);
nand U12659 (N_12659,N_11859,N_11158);
or U12660 (N_12660,N_11571,N_11692);
and U12661 (N_12661,N_11400,N_11053);
nor U12662 (N_12662,N_11675,N_11119);
nor U12663 (N_12663,N_11506,N_11332);
or U12664 (N_12664,N_11282,N_11031);
and U12665 (N_12665,N_11158,N_11308);
and U12666 (N_12666,N_11513,N_11496);
nor U12667 (N_12667,N_11523,N_11220);
or U12668 (N_12668,N_11437,N_11659);
and U12669 (N_12669,N_11066,N_11839);
nor U12670 (N_12670,N_11777,N_11490);
nand U12671 (N_12671,N_11754,N_11687);
and U12672 (N_12672,N_11230,N_11898);
and U12673 (N_12673,N_11976,N_11543);
and U12674 (N_12674,N_11865,N_11710);
and U12675 (N_12675,N_11001,N_11806);
nor U12676 (N_12676,N_11269,N_11456);
or U12677 (N_12677,N_11351,N_11700);
xor U12678 (N_12678,N_11228,N_11171);
xnor U12679 (N_12679,N_11478,N_11127);
xor U12680 (N_12680,N_11521,N_11589);
nor U12681 (N_12681,N_11233,N_11754);
and U12682 (N_12682,N_11655,N_11835);
or U12683 (N_12683,N_11471,N_11203);
nor U12684 (N_12684,N_11127,N_11186);
nor U12685 (N_12685,N_11310,N_11581);
and U12686 (N_12686,N_11803,N_11194);
nor U12687 (N_12687,N_11522,N_11251);
and U12688 (N_12688,N_11307,N_11141);
xnor U12689 (N_12689,N_11079,N_11203);
and U12690 (N_12690,N_11013,N_11776);
or U12691 (N_12691,N_11637,N_11439);
nor U12692 (N_12692,N_11909,N_11747);
and U12693 (N_12693,N_11757,N_11505);
or U12694 (N_12694,N_11370,N_11651);
xnor U12695 (N_12695,N_11255,N_11093);
or U12696 (N_12696,N_11475,N_11141);
or U12697 (N_12697,N_11861,N_11259);
xnor U12698 (N_12698,N_11052,N_11253);
nor U12699 (N_12699,N_11696,N_11659);
or U12700 (N_12700,N_11739,N_11998);
nand U12701 (N_12701,N_11544,N_11716);
nor U12702 (N_12702,N_11384,N_11724);
xnor U12703 (N_12703,N_11780,N_11699);
nand U12704 (N_12704,N_11754,N_11223);
xnor U12705 (N_12705,N_11547,N_11284);
xor U12706 (N_12706,N_11823,N_11879);
nor U12707 (N_12707,N_11877,N_11939);
or U12708 (N_12708,N_11769,N_11385);
nor U12709 (N_12709,N_11733,N_11737);
or U12710 (N_12710,N_11140,N_11744);
and U12711 (N_12711,N_11248,N_11588);
nor U12712 (N_12712,N_11107,N_11239);
nand U12713 (N_12713,N_11784,N_11075);
nor U12714 (N_12714,N_11390,N_11646);
or U12715 (N_12715,N_11925,N_11530);
nand U12716 (N_12716,N_11027,N_11896);
and U12717 (N_12717,N_11618,N_11301);
nand U12718 (N_12718,N_11607,N_11775);
xnor U12719 (N_12719,N_11754,N_11671);
nand U12720 (N_12720,N_11904,N_11522);
nand U12721 (N_12721,N_11003,N_11732);
xor U12722 (N_12722,N_11382,N_11375);
or U12723 (N_12723,N_11629,N_11080);
and U12724 (N_12724,N_11943,N_11744);
xnor U12725 (N_12725,N_11383,N_11939);
and U12726 (N_12726,N_11541,N_11882);
xnor U12727 (N_12727,N_11630,N_11373);
nand U12728 (N_12728,N_11788,N_11352);
xnor U12729 (N_12729,N_11753,N_11151);
xor U12730 (N_12730,N_11121,N_11438);
xor U12731 (N_12731,N_11003,N_11432);
xnor U12732 (N_12732,N_11529,N_11226);
or U12733 (N_12733,N_11577,N_11606);
nor U12734 (N_12734,N_11052,N_11637);
or U12735 (N_12735,N_11317,N_11495);
nand U12736 (N_12736,N_11842,N_11633);
nand U12737 (N_12737,N_11963,N_11054);
or U12738 (N_12738,N_11987,N_11719);
and U12739 (N_12739,N_11548,N_11025);
or U12740 (N_12740,N_11909,N_11553);
and U12741 (N_12741,N_11770,N_11869);
nand U12742 (N_12742,N_11695,N_11577);
xor U12743 (N_12743,N_11222,N_11711);
and U12744 (N_12744,N_11444,N_11475);
or U12745 (N_12745,N_11116,N_11638);
xor U12746 (N_12746,N_11495,N_11313);
nand U12747 (N_12747,N_11359,N_11048);
nor U12748 (N_12748,N_11031,N_11811);
xor U12749 (N_12749,N_11632,N_11530);
nor U12750 (N_12750,N_11831,N_11840);
nor U12751 (N_12751,N_11762,N_11004);
nor U12752 (N_12752,N_11657,N_11392);
or U12753 (N_12753,N_11811,N_11675);
or U12754 (N_12754,N_11264,N_11640);
nor U12755 (N_12755,N_11312,N_11681);
or U12756 (N_12756,N_11600,N_11945);
nand U12757 (N_12757,N_11957,N_11247);
nand U12758 (N_12758,N_11031,N_11757);
and U12759 (N_12759,N_11130,N_11279);
nor U12760 (N_12760,N_11564,N_11017);
or U12761 (N_12761,N_11330,N_11009);
xor U12762 (N_12762,N_11182,N_11105);
nor U12763 (N_12763,N_11173,N_11647);
xnor U12764 (N_12764,N_11060,N_11050);
xnor U12765 (N_12765,N_11279,N_11142);
or U12766 (N_12766,N_11445,N_11696);
nor U12767 (N_12767,N_11856,N_11721);
nand U12768 (N_12768,N_11925,N_11860);
xor U12769 (N_12769,N_11045,N_11706);
nor U12770 (N_12770,N_11320,N_11819);
or U12771 (N_12771,N_11420,N_11354);
and U12772 (N_12772,N_11161,N_11235);
or U12773 (N_12773,N_11969,N_11977);
or U12774 (N_12774,N_11456,N_11761);
or U12775 (N_12775,N_11512,N_11984);
or U12776 (N_12776,N_11313,N_11386);
xnor U12777 (N_12777,N_11055,N_11565);
nor U12778 (N_12778,N_11801,N_11505);
or U12779 (N_12779,N_11910,N_11905);
or U12780 (N_12780,N_11931,N_11936);
nand U12781 (N_12781,N_11773,N_11727);
or U12782 (N_12782,N_11615,N_11134);
nor U12783 (N_12783,N_11056,N_11699);
nand U12784 (N_12784,N_11060,N_11665);
xor U12785 (N_12785,N_11155,N_11969);
and U12786 (N_12786,N_11759,N_11479);
nand U12787 (N_12787,N_11839,N_11842);
xor U12788 (N_12788,N_11339,N_11287);
nor U12789 (N_12789,N_11101,N_11499);
nor U12790 (N_12790,N_11825,N_11086);
xnor U12791 (N_12791,N_11082,N_11506);
or U12792 (N_12792,N_11321,N_11636);
xnor U12793 (N_12793,N_11072,N_11478);
or U12794 (N_12794,N_11292,N_11251);
nand U12795 (N_12795,N_11277,N_11189);
nor U12796 (N_12796,N_11873,N_11814);
nor U12797 (N_12797,N_11752,N_11108);
nand U12798 (N_12798,N_11369,N_11266);
nor U12799 (N_12799,N_11207,N_11425);
nor U12800 (N_12800,N_11483,N_11388);
and U12801 (N_12801,N_11576,N_11335);
nor U12802 (N_12802,N_11308,N_11077);
or U12803 (N_12803,N_11258,N_11038);
or U12804 (N_12804,N_11818,N_11881);
nor U12805 (N_12805,N_11183,N_11461);
nand U12806 (N_12806,N_11074,N_11775);
and U12807 (N_12807,N_11724,N_11216);
nand U12808 (N_12808,N_11783,N_11890);
nand U12809 (N_12809,N_11208,N_11506);
and U12810 (N_12810,N_11816,N_11510);
nor U12811 (N_12811,N_11059,N_11018);
nand U12812 (N_12812,N_11174,N_11392);
or U12813 (N_12813,N_11323,N_11186);
and U12814 (N_12814,N_11894,N_11936);
nand U12815 (N_12815,N_11558,N_11560);
or U12816 (N_12816,N_11304,N_11184);
nand U12817 (N_12817,N_11111,N_11777);
nor U12818 (N_12818,N_11070,N_11779);
or U12819 (N_12819,N_11772,N_11393);
nand U12820 (N_12820,N_11348,N_11244);
and U12821 (N_12821,N_11455,N_11873);
nand U12822 (N_12822,N_11114,N_11604);
xor U12823 (N_12823,N_11309,N_11406);
xor U12824 (N_12824,N_11933,N_11184);
nor U12825 (N_12825,N_11065,N_11229);
and U12826 (N_12826,N_11568,N_11312);
xor U12827 (N_12827,N_11110,N_11873);
or U12828 (N_12828,N_11348,N_11674);
nor U12829 (N_12829,N_11489,N_11326);
nor U12830 (N_12830,N_11851,N_11558);
nor U12831 (N_12831,N_11335,N_11552);
and U12832 (N_12832,N_11331,N_11385);
and U12833 (N_12833,N_11616,N_11974);
and U12834 (N_12834,N_11475,N_11693);
or U12835 (N_12835,N_11102,N_11811);
or U12836 (N_12836,N_11287,N_11511);
xnor U12837 (N_12837,N_11904,N_11724);
and U12838 (N_12838,N_11005,N_11028);
xnor U12839 (N_12839,N_11419,N_11631);
nor U12840 (N_12840,N_11129,N_11748);
nand U12841 (N_12841,N_11041,N_11341);
nand U12842 (N_12842,N_11100,N_11964);
or U12843 (N_12843,N_11404,N_11177);
nor U12844 (N_12844,N_11470,N_11077);
xnor U12845 (N_12845,N_11454,N_11961);
or U12846 (N_12846,N_11242,N_11336);
and U12847 (N_12847,N_11645,N_11744);
nand U12848 (N_12848,N_11773,N_11647);
nor U12849 (N_12849,N_11587,N_11280);
nor U12850 (N_12850,N_11141,N_11673);
xor U12851 (N_12851,N_11075,N_11795);
or U12852 (N_12852,N_11478,N_11338);
or U12853 (N_12853,N_11210,N_11746);
xnor U12854 (N_12854,N_11206,N_11193);
or U12855 (N_12855,N_11672,N_11369);
xnor U12856 (N_12856,N_11311,N_11232);
or U12857 (N_12857,N_11821,N_11545);
nand U12858 (N_12858,N_11337,N_11148);
xor U12859 (N_12859,N_11267,N_11245);
and U12860 (N_12860,N_11657,N_11931);
or U12861 (N_12861,N_11461,N_11221);
xnor U12862 (N_12862,N_11181,N_11433);
or U12863 (N_12863,N_11311,N_11279);
xnor U12864 (N_12864,N_11181,N_11664);
nand U12865 (N_12865,N_11383,N_11771);
and U12866 (N_12866,N_11022,N_11186);
nor U12867 (N_12867,N_11241,N_11856);
nor U12868 (N_12868,N_11972,N_11351);
and U12869 (N_12869,N_11962,N_11352);
and U12870 (N_12870,N_11742,N_11890);
nor U12871 (N_12871,N_11902,N_11154);
xor U12872 (N_12872,N_11882,N_11111);
xor U12873 (N_12873,N_11074,N_11385);
and U12874 (N_12874,N_11070,N_11985);
and U12875 (N_12875,N_11362,N_11321);
and U12876 (N_12876,N_11328,N_11062);
nand U12877 (N_12877,N_11246,N_11325);
or U12878 (N_12878,N_11697,N_11079);
xor U12879 (N_12879,N_11915,N_11863);
nor U12880 (N_12880,N_11184,N_11288);
nor U12881 (N_12881,N_11995,N_11279);
xor U12882 (N_12882,N_11983,N_11905);
nor U12883 (N_12883,N_11271,N_11569);
xnor U12884 (N_12884,N_11672,N_11150);
or U12885 (N_12885,N_11402,N_11168);
nor U12886 (N_12886,N_11508,N_11713);
or U12887 (N_12887,N_11701,N_11627);
xor U12888 (N_12888,N_11151,N_11083);
nor U12889 (N_12889,N_11720,N_11175);
nor U12890 (N_12890,N_11834,N_11134);
xor U12891 (N_12891,N_11733,N_11411);
xor U12892 (N_12892,N_11670,N_11538);
nor U12893 (N_12893,N_11966,N_11811);
xnor U12894 (N_12894,N_11030,N_11514);
xnor U12895 (N_12895,N_11573,N_11264);
nor U12896 (N_12896,N_11277,N_11634);
xor U12897 (N_12897,N_11911,N_11582);
or U12898 (N_12898,N_11036,N_11524);
nand U12899 (N_12899,N_11533,N_11206);
or U12900 (N_12900,N_11515,N_11299);
nand U12901 (N_12901,N_11272,N_11911);
and U12902 (N_12902,N_11517,N_11541);
nand U12903 (N_12903,N_11742,N_11434);
and U12904 (N_12904,N_11891,N_11953);
nand U12905 (N_12905,N_11865,N_11522);
xor U12906 (N_12906,N_11303,N_11610);
or U12907 (N_12907,N_11069,N_11053);
nand U12908 (N_12908,N_11768,N_11117);
xnor U12909 (N_12909,N_11307,N_11137);
nand U12910 (N_12910,N_11985,N_11630);
nand U12911 (N_12911,N_11127,N_11937);
nor U12912 (N_12912,N_11136,N_11774);
xor U12913 (N_12913,N_11095,N_11428);
xnor U12914 (N_12914,N_11978,N_11540);
and U12915 (N_12915,N_11962,N_11252);
nand U12916 (N_12916,N_11991,N_11043);
nor U12917 (N_12917,N_11589,N_11721);
or U12918 (N_12918,N_11119,N_11590);
and U12919 (N_12919,N_11357,N_11612);
nand U12920 (N_12920,N_11073,N_11806);
nor U12921 (N_12921,N_11980,N_11746);
and U12922 (N_12922,N_11000,N_11946);
or U12923 (N_12923,N_11996,N_11150);
nand U12924 (N_12924,N_11474,N_11898);
nor U12925 (N_12925,N_11657,N_11914);
and U12926 (N_12926,N_11122,N_11681);
xnor U12927 (N_12927,N_11067,N_11761);
nand U12928 (N_12928,N_11684,N_11978);
nor U12929 (N_12929,N_11994,N_11345);
nand U12930 (N_12930,N_11290,N_11811);
xnor U12931 (N_12931,N_11424,N_11675);
or U12932 (N_12932,N_11077,N_11404);
or U12933 (N_12933,N_11919,N_11397);
or U12934 (N_12934,N_11004,N_11315);
or U12935 (N_12935,N_11071,N_11074);
nand U12936 (N_12936,N_11644,N_11261);
nor U12937 (N_12937,N_11380,N_11708);
xor U12938 (N_12938,N_11299,N_11413);
or U12939 (N_12939,N_11844,N_11848);
and U12940 (N_12940,N_11917,N_11389);
xnor U12941 (N_12941,N_11934,N_11114);
and U12942 (N_12942,N_11196,N_11719);
or U12943 (N_12943,N_11900,N_11835);
nor U12944 (N_12944,N_11013,N_11475);
nand U12945 (N_12945,N_11584,N_11437);
or U12946 (N_12946,N_11700,N_11682);
or U12947 (N_12947,N_11553,N_11929);
nor U12948 (N_12948,N_11726,N_11061);
nor U12949 (N_12949,N_11869,N_11904);
or U12950 (N_12950,N_11460,N_11245);
nor U12951 (N_12951,N_11094,N_11585);
nand U12952 (N_12952,N_11851,N_11169);
nor U12953 (N_12953,N_11088,N_11107);
nor U12954 (N_12954,N_11176,N_11003);
xor U12955 (N_12955,N_11912,N_11837);
nor U12956 (N_12956,N_11433,N_11564);
xnor U12957 (N_12957,N_11874,N_11585);
nand U12958 (N_12958,N_11400,N_11531);
xor U12959 (N_12959,N_11216,N_11743);
xnor U12960 (N_12960,N_11381,N_11494);
xnor U12961 (N_12961,N_11974,N_11625);
or U12962 (N_12962,N_11165,N_11962);
nor U12963 (N_12963,N_11337,N_11098);
xor U12964 (N_12964,N_11728,N_11417);
xnor U12965 (N_12965,N_11756,N_11675);
nor U12966 (N_12966,N_11949,N_11047);
and U12967 (N_12967,N_11967,N_11106);
or U12968 (N_12968,N_11642,N_11218);
or U12969 (N_12969,N_11712,N_11057);
xnor U12970 (N_12970,N_11179,N_11031);
or U12971 (N_12971,N_11728,N_11332);
xnor U12972 (N_12972,N_11905,N_11935);
or U12973 (N_12973,N_11743,N_11591);
nor U12974 (N_12974,N_11199,N_11699);
nand U12975 (N_12975,N_11472,N_11398);
nor U12976 (N_12976,N_11510,N_11400);
or U12977 (N_12977,N_11240,N_11911);
xor U12978 (N_12978,N_11188,N_11527);
xnor U12979 (N_12979,N_11816,N_11809);
nand U12980 (N_12980,N_11421,N_11909);
xor U12981 (N_12981,N_11741,N_11596);
nand U12982 (N_12982,N_11115,N_11976);
xor U12983 (N_12983,N_11366,N_11428);
or U12984 (N_12984,N_11520,N_11697);
xnor U12985 (N_12985,N_11344,N_11761);
and U12986 (N_12986,N_11691,N_11381);
xor U12987 (N_12987,N_11557,N_11757);
nand U12988 (N_12988,N_11593,N_11477);
or U12989 (N_12989,N_11299,N_11961);
nand U12990 (N_12990,N_11188,N_11534);
and U12991 (N_12991,N_11972,N_11650);
nor U12992 (N_12992,N_11914,N_11728);
or U12993 (N_12993,N_11197,N_11740);
or U12994 (N_12994,N_11815,N_11018);
nand U12995 (N_12995,N_11501,N_11467);
xnor U12996 (N_12996,N_11845,N_11500);
or U12997 (N_12997,N_11206,N_11643);
xor U12998 (N_12998,N_11208,N_11367);
nor U12999 (N_12999,N_11562,N_11608);
xnor U13000 (N_13000,N_12448,N_12478);
nand U13001 (N_13001,N_12468,N_12158);
or U13002 (N_13002,N_12852,N_12427);
nand U13003 (N_13003,N_12167,N_12419);
xor U13004 (N_13004,N_12637,N_12494);
nand U13005 (N_13005,N_12923,N_12596);
nor U13006 (N_13006,N_12324,N_12995);
nand U13007 (N_13007,N_12517,N_12997);
nand U13008 (N_13008,N_12524,N_12193);
and U13009 (N_13009,N_12213,N_12134);
or U13010 (N_13010,N_12713,N_12571);
nor U13011 (N_13011,N_12679,N_12576);
nand U13012 (N_13012,N_12646,N_12858);
or U13013 (N_13013,N_12741,N_12699);
nor U13014 (N_13014,N_12509,N_12957);
nor U13015 (N_13015,N_12212,N_12444);
and U13016 (N_13016,N_12023,N_12716);
or U13017 (N_13017,N_12674,N_12166);
nor U13018 (N_13018,N_12283,N_12927);
or U13019 (N_13019,N_12019,N_12221);
and U13020 (N_13020,N_12278,N_12626);
or U13021 (N_13021,N_12085,N_12941);
or U13022 (N_13022,N_12835,N_12895);
or U13023 (N_13023,N_12773,N_12216);
or U13024 (N_13024,N_12628,N_12723);
nand U13025 (N_13025,N_12779,N_12873);
nor U13026 (N_13026,N_12218,N_12263);
or U13027 (N_13027,N_12132,N_12017);
or U13028 (N_13028,N_12762,N_12799);
and U13029 (N_13029,N_12244,N_12705);
nand U13030 (N_13030,N_12093,N_12590);
or U13031 (N_13031,N_12230,N_12503);
or U13032 (N_13032,N_12714,N_12630);
or U13033 (N_13033,N_12165,N_12528);
nor U13034 (N_13034,N_12840,N_12574);
nor U13035 (N_13035,N_12903,N_12098);
nand U13036 (N_13036,N_12789,N_12354);
xor U13037 (N_13037,N_12822,N_12851);
xor U13038 (N_13038,N_12692,N_12560);
nand U13039 (N_13039,N_12638,N_12855);
nand U13040 (N_13040,N_12090,N_12872);
or U13041 (N_13041,N_12422,N_12170);
nand U13042 (N_13042,N_12141,N_12575);
nand U13043 (N_13043,N_12512,N_12377);
nand U13044 (N_13044,N_12437,N_12355);
and U13045 (N_13045,N_12272,N_12916);
nor U13046 (N_13046,N_12235,N_12197);
and U13047 (N_13047,N_12340,N_12955);
xnor U13048 (N_13048,N_12857,N_12209);
nor U13049 (N_13049,N_12959,N_12695);
nor U13050 (N_13050,N_12759,N_12388);
or U13051 (N_13051,N_12318,N_12189);
nand U13052 (N_13052,N_12529,N_12942);
nand U13053 (N_13053,N_12373,N_12070);
nand U13054 (N_13054,N_12492,N_12949);
or U13055 (N_13055,N_12884,N_12499);
and U13056 (N_13056,N_12184,N_12636);
or U13057 (N_13057,N_12936,N_12386);
and U13058 (N_13058,N_12076,N_12527);
xor U13059 (N_13059,N_12930,N_12645);
xor U13060 (N_13060,N_12135,N_12103);
xnor U13061 (N_13061,N_12801,N_12832);
nand U13062 (N_13062,N_12069,N_12876);
xnor U13063 (N_13063,N_12077,N_12378);
xnor U13064 (N_13064,N_12042,N_12776);
nand U13065 (N_13065,N_12068,N_12680);
nand U13066 (N_13066,N_12345,N_12127);
xor U13067 (N_13067,N_12697,N_12176);
xnor U13068 (N_13068,N_12627,N_12972);
nor U13069 (N_13069,N_12234,N_12183);
and U13070 (N_13070,N_12612,N_12943);
or U13071 (N_13071,N_12486,N_12353);
or U13072 (N_13072,N_12225,N_12771);
nand U13073 (N_13073,N_12429,N_12635);
xnor U13074 (N_13074,N_12298,N_12276);
xor U13075 (N_13075,N_12553,N_12702);
xnor U13076 (N_13076,N_12660,N_12744);
nor U13077 (N_13077,N_12124,N_12530);
or U13078 (N_13078,N_12296,N_12459);
nand U13079 (N_13079,N_12672,N_12721);
or U13080 (N_13080,N_12161,N_12010);
nand U13081 (N_13081,N_12048,N_12902);
xor U13082 (N_13082,N_12964,N_12177);
xor U13083 (N_13083,N_12515,N_12411);
or U13084 (N_13084,N_12506,N_12752);
nand U13085 (N_13085,N_12226,N_12201);
and U13086 (N_13086,N_12996,N_12531);
and U13087 (N_13087,N_12266,N_12642);
xnor U13088 (N_13088,N_12569,N_12675);
and U13089 (N_13089,N_12656,N_12446);
nand U13090 (N_13090,N_12152,N_12875);
or U13091 (N_13091,N_12814,N_12215);
nand U13092 (N_13092,N_12862,N_12271);
nand U13093 (N_13093,N_12089,N_12322);
xnor U13094 (N_13094,N_12368,N_12262);
and U13095 (N_13095,N_12175,N_12409);
nor U13096 (N_13096,N_12921,N_12479);
nand U13097 (N_13097,N_12319,N_12313);
nand U13098 (N_13098,N_12620,N_12148);
or U13099 (N_13099,N_12982,N_12097);
or U13100 (N_13100,N_12860,N_12570);
or U13101 (N_13101,N_12102,N_12761);
xnor U13102 (N_13102,N_12687,N_12920);
nor U13103 (N_13103,N_12611,N_12182);
xnor U13104 (N_13104,N_12131,N_12844);
nor U13105 (N_13105,N_12770,N_12990);
xnor U13106 (N_13106,N_12362,N_12836);
xor U13107 (N_13107,N_12772,N_12281);
and U13108 (N_13108,N_12797,N_12550);
or U13109 (N_13109,N_12588,N_12008);
nor U13110 (N_13110,N_12979,N_12586);
and U13111 (N_13111,N_12824,N_12028);
xor U13112 (N_13112,N_12798,N_12168);
nand U13113 (N_13113,N_12109,N_12379);
and U13114 (N_13114,N_12350,N_12326);
nor U13115 (N_13115,N_12467,N_12243);
or U13116 (N_13116,N_12154,N_12540);
nand U13117 (N_13117,N_12328,N_12986);
or U13118 (N_13118,N_12677,N_12587);
xor U13119 (N_13119,N_12060,N_12147);
xnor U13120 (N_13120,N_12805,N_12537);
nor U13121 (N_13121,N_12732,N_12595);
xor U13122 (N_13122,N_12849,N_12399);
xnor U13123 (N_13123,N_12347,N_12589);
nand U13124 (N_13124,N_12274,N_12864);
and U13125 (N_13125,N_12025,N_12129);
and U13126 (N_13126,N_12160,N_12380);
xor U13127 (N_13127,N_12623,N_12480);
and U13128 (N_13128,N_12790,N_12662);
nand U13129 (N_13129,N_12178,N_12251);
nand U13130 (N_13130,N_12375,N_12180);
nand U13131 (N_13131,N_12254,N_12412);
and U13132 (N_13132,N_12162,N_12036);
nor U13133 (N_13133,N_12848,N_12004);
and U13134 (N_13134,N_12746,N_12603);
xor U13135 (N_13135,N_12066,N_12397);
xor U13136 (N_13136,N_12498,N_12335);
xor U13137 (N_13137,N_12892,N_12100);
nor U13138 (N_13138,N_12608,N_12303);
nor U13139 (N_13139,N_12634,N_12242);
or U13140 (N_13140,N_12426,N_12227);
or U13141 (N_13141,N_12079,N_12461);
or U13142 (N_13142,N_12548,N_12153);
xor U13143 (N_13143,N_12150,N_12998);
and U13144 (N_13144,N_12317,N_12974);
and U13145 (N_13145,N_12658,N_12250);
xnor U13146 (N_13146,N_12223,N_12821);
or U13147 (N_13147,N_12554,N_12406);
xnor U13148 (N_13148,N_12035,N_12891);
nor U13149 (N_13149,N_12051,N_12403);
and U13150 (N_13150,N_12074,N_12791);
xnor U13151 (N_13151,N_12592,N_12126);
xnor U13152 (N_13152,N_12806,N_12453);
or U13153 (N_13153,N_12146,N_12958);
nor U13154 (N_13154,N_12113,N_12624);
nand U13155 (N_13155,N_12044,N_12925);
and U13156 (N_13156,N_12615,N_12885);
xor U13157 (N_13157,N_12745,N_12879);
and U13158 (N_13158,N_12014,N_12483);
xor U13159 (N_13159,N_12039,N_12617);
nand U13160 (N_13160,N_12470,N_12447);
nor U13161 (N_13161,N_12064,N_12522);
or U13162 (N_13162,N_12749,N_12676);
nand U13163 (N_13163,N_12555,N_12561);
nor U13164 (N_13164,N_12632,N_12142);
and U13165 (N_13165,N_12577,N_12484);
and U13166 (N_13166,N_12562,N_12719);
or U13167 (N_13167,N_12402,N_12265);
or U13168 (N_13168,N_12727,N_12031);
xnor U13169 (N_13169,N_12246,N_12295);
and U13170 (N_13170,N_12502,N_12698);
nor U13171 (N_13171,N_12393,N_12880);
xor U13172 (N_13172,N_12214,N_12984);
nor U13173 (N_13173,N_12735,N_12711);
nand U13174 (N_13174,N_12939,N_12725);
nand U13175 (N_13175,N_12482,N_12953);
or U13176 (N_13176,N_12471,N_12788);
or U13177 (N_13177,N_12659,N_12436);
and U13178 (N_13178,N_12785,N_12123);
nor U13179 (N_13179,N_12294,N_12720);
or U13180 (N_13180,N_12544,N_12121);
nand U13181 (N_13181,N_12424,N_12080);
or U13182 (N_13182,N_12906,N_12975);
and U13183 (N_13183,N_12803,N_12756);
and U13184 (N_13184,N_12690,N_12384);
nor U13185 (N_13185,N_12137,N_12673);
or U13186 (N_13186,N_12534,N_12866);
xnor U13187 (N_13187,N_12049,N_12703);
nand U13188 (N_13188,N_12606,N_12889);
or U13189 (N_13189,N_12715,N_12289);
xnor U13190 (N_13190,N_12466,N_12253);
nand U13191 (N_13191,N_12099,N_12978);
nand U13192 (N_13192,N_12918,N_12348);
or U13193 (N_13193,N_12087,N_12839);
xnor U13194 (N_13194,N_12969,N_12913);
nor U13195 (N_13195,N_12107,N_12582);
nand U13196 (N_13196,N_12143,N_12363);
and U13197 (N_13197,N_12516,N_12956);
and U13198 (N_13198,N_12033,N_12372);
or U13199 (N_13199,N_12259,N_12869);
or U13200 (N_13200,N_12245,N_12417);
xnor U13201 (N_13201,N_12490,N_12547);
nand U13202 (N_13202,N_12346,N_12613);
nor U13203 (N_13203,N_12401,N_12452);
and U13204 (N_13204,N_12757,N_12204);
and U13205 (N_13205,N_12344,N_12256);
and U13206 (N_13206,N_12130,N_12546);
xor U13207 (N_13207,N_12750,N_12261);
nand U13208 (N_13208,N_12946,N_12200);
nand U13209 (N_13209,N_12738,N_12106);
or U13210 (N_13210,N_12600,N_12886);
nand U13211 (N_13211,N_12011,N_12774);
and U13212 (N_13212,N_12022,N_12542);
or U13213 (N_13213,N_12641,N_12138);
or U13214 (N_13214,N_12309,N_12240);
xnor U13215 (N_13215,N_12700,N_12172);
or U13216 (N_13216,N_12445,N_12909);
nor U13217 (N_13217,N_12981,N_12139);
xor U13218 (N_13218,N_12451,N_12668);
or U13219 (N_13219,N_12888,N_12707);
nand U13220 (N_13220,N_12464,N_12859);
xor U13221 (N_13221,N_12140,N_12144);
and U13222 (N_13222,N_12476,N_12911);
xor U13223 (N_13223,N_12601,N_12977);
nand U13224 (N_13224,N_12754,N_12369);
nor U13225 (N_13225,N_12329,N_12360);
xnor U13226 (N_13226,N_12057,N_12118);
or U13227 (N_13227,N_12210,N_12654);
xor U13228 (N_13228,N_12398,N_12222);
nand U13229 (N_13229,N_12050,N_12032);
nand U13230 (N_13230,N_12951,N_12430);
nor U13231 (N_13231,N_12067,N_12096);
and U13232 (N_13232,N_12151,N_12812);
nor U13233 (N_13233,N_12449,N_12105);
or U13234 (N_13234,N_12894,N_12332);
or U13235 (N_13235,N_12046,N_12633);
nand U13236 (N_13236,N_12693,N_12462);
nand U13237 (N_13237,N_12370,N_12922);
nand U13238 (N_13238,N_12198,N_12709);
and U13239 (N_13239,N_12813,N_12683);
and U13240 (N_13240,N_12513,N_12287);
nand U13241 (N_13241,N_12463,N_12030);
and U13242 (N_13242,N_12568,N_12962);
nand U13243 (N_13243,N_12685,N_12795);
or U13244 (N_13244,N_12382,N_12435);
xnor U13245 (N_13245,N_12258,N_12686);
nand U13246 (N_13246,N_12907,N_12514);
nand U13247 (N_13247,N_12657,N_12358);
nor U13248 (N_13248,N_12432,N_12604);
nand U13249 (N_13249,N_12357,N_12924);
or U13250 (N_13250,N_12441,N_12965);
nor U13251 (N_13251,N_12865,N_12063);
nand U13252 (N_13252,N_12861,N_12914);
nor U13253 (N_13253,N_12456,N_12999);
and U13254 (N_13254,N_12784,N_12396);
or U13255 (N_13255,N_12766,N_12820);
nor U13256 (N_13256,N_12301,N_12901);
and U13257 (N_13257,N_12199,N_12117);
xnor U13258 (N_13258,N_12739,N_12081);
nand U13259 (N_13259,N_12352,N_12248);
and U13260 (N_13260,N_12616,N_12334);
or U13261 (N_13261,N_12431,N_12605);
nand U13262 (N_13262,N_12648,N_12538);
nor U13263 (N_13263,N_12418,N_12159);
nor U13264 (N_13264,N_12898,N_12233);
xor U13265 (N_13265,N_12663,N_12194);
nand U13266 (N_13266,N_12325,N_12708);
or U13267 (N_13267,N_12056,N_12807);
or U13268 (N_13268,N_12917,N_12778);
and U13269 (N_13269,N_12652,N_12163);
nor U13270 (N_13270,N_12853,N_12751);
and U13271 (N_13271,N_12012,N_12543);
nand U13272 (N_13272,N_12169,N_12566);
nand U13273 (N_13273,N_12491,N_12238);
nor U13274 (N_13274,N_12868,N_12818);
nand U13275 (N_13275,N_12496,N_12816);
nor U13276 (N_13276,N_12838,N_12960);
nor U13277 (N_13277,N_12661,N_12190);
xor U13278 (N_13278,N_12434,N_12521);
nor U13279 (N_13279,N_12000,N_12239);
nand U13280 (N_13280,N_12366,N_12205);
nand U13281 (N_13281,N_12228,N_12217);
and U13282 (N_13282,N_12810,N_12501);
or U13283 (N_13283,N_12450,N_12910);
and U13284 (N_13284,N_12800,N_12195);
nand U13285 (N_13285,N_12224,N_12336);
or U13286 (N_13286,N_12564,N_12730);
xor U13287 (N_13287,N_12830,N_12967);
xor U13288 (N_13288,N_12045,N_12072);
nor U13289 (N_13289,N_12013,N_12185);
nor U13290 (N_13290,N_12084,N_12856);
and U13291 (N_13291,N_12696,N_12394);
nor U13292 (N_13292,N_12473,N_12095);
and U13293 (N_13293,N_12614,N_12966);
xor U13294 (N_13294,N_12061,N_12594);
and U13295 (N_13295,N_12487,N_12833);
and U13296 (N_13296,N_12780,N_12877);
or U13297 (N_13297,N_12112,N_12665);
and U13298 (N_13298,N_12310,N_12742);
xnor U13299 (N_13299,N_12383,N_12871);
nand U13300 (N_13300,N_12992,N_12987);
or U13301 (N_13301,N_12622,N_12088);
nand U13302 (N_13302,N_12405,N_12015);
or U13303 (N_13303,N_12120,N_12125);
nand U13304 (N_13304,N_12629,N_12481);
and U13305 (N_13305,N_12580,N_12994);
and U13306 (N_13306,N_12808,N_12187);
nand U13307 (N_13307,N_12255,N_12058);
and U13308 (N_13308,N_12518,N_12883);
xor U13309 (N_13309,N_12179,N_12082);
and U13310 (N_13310,N_12433,N_12331);
nand U13311 (N_13311,N_12947,N_12395);
or U13312 (N_13312,N_12333,N_12438);
xor U13313 (N_13313,N_12414,N_12108);
or U13314 (N_13314,N_12653,N_12579);
nor U13315 (N_13315,N_12071,N_12323);
xnor U13316 (N_13316,N_12937,N_12706);
xor U13317 (N_13317,N_12710,N_12915);
nor U13318 (N_13318,N_12110,N_12878);
nor U13319 (N_13319,N_12508,N_12954);
nand U13320 (N_13320,N_12989,N_12796);
and U13321 (N_13321,N_12489,N_12122);
or U13322 (N_13322,N_12610,N_12507);
and U13323 (N_13323,N_12863,N_12038);
nand U13324 (N_13324,N_12231,N_12578);
nand U13325 (N_13325,N_12728,N_12269);
nand U13326 (N_13326,N_12339,N_12841);
and U13327 (N_13327,N_12005,N_12306);
nor U13328 (N_13328,N_12171,N_12743);
and U13329 (N_13329,N_12273,N_12619);
nor U13330 (N_13330,N_12241,N_12704);
nand U13331 (N_13331,N_12961,N_12767);
xnor U13332 (N_13332,N_12155,N_12850);
xor U13333 (N_13333,N_12493,N_12500);
nor U13334 (N_13334,N_12181,N_12037);
or U13335 (N_13335,N_12196,N_12440);
nand U13336 (N_13336,N_12647,N_12689);
xor U13337 (N_13337,N_12718,N_12279);
nor U13338 (N_13338,N_12760,N_12607);
or U13339 (N_13339,N_12991,N_12504);
xor U13340 (N_13340,N_12034,N_12938);
nand U13341 (N_13341,N_12469,N_12302);
or U13342 (N_13342,N_12712,N_12391);
nand U13343 (N_13343,N_12264,N_12374);
and U13344 (N_13344,N_12367,N_12428);
and U13345 (N_13345,N_12284,N_12202);
or U13346 (N_13346,N_12091,N_12308);
and U13347 (N_13347,N_12305,N_12846);
nand U13348 (N_13348,N_12236,N_12455);
and U13349 (N_13349,N_12136,N_12041);
nor U13350 (N_13350,N_12421,N_12678);
nand U13351 (N_13351,N_12003,N_12342);
or U13352 (N_13352,N_12511,N_12389);
xor U13353 (N_13353,N_12387,N_12655);
xnor U13354 (N_13354,N_12315,N_12926);
and U13355 (N_13355,N_12985,N_12343);
and U13356 (N_13356,N_12040,N_12018);
and U13357 (N_13357,N_12945,N_12485);
xnor U13358 (N_13358,N_12585,N_12940);
or U13359 (N_13359,N_12400,N_12581);
xnor U13360 (N_13360,N_12726,N_12359);
or U13361 (N_13361,N_12731,N_12073);
and U13362 (N_13362,N_12599,N_12206);
and U13363 (N_13363,N_12312,N_12474);
nor U13364 (N_13364,N_12293,N_12684);
nand U13365 (N_13365,N_12912,N_12993);
or U13366 (N_13366,N_12845,N_12442);
nand U13367 (N_13367,N_12327,N_12029);
xnor U13368 (N_13368,N_12618,N_12681);
nand U13369 (N_13369,N_12001,N_12829);
nand U13370 (N_13370,N_12104,N_12908);
nand U13371 (N_13371,N_12270,N_12817);
and U13372 (N_13372,N_12968,N_12052);
xor U13373 (N_13373,N_12827,N_12247);
xnor U13374 (N_13374,N_12900,N_12783);
nand U13375 (N_13375,N_12532,N_12598);
and U13376 (N_13376,N_12458,N_12988);
nand U13377 (N_13377,N_12929,N_12682);
nand U13378 (N_13378,N_12219,N_12465);
xor U13379 (N_13379,N_12823,N_12016);
and U13380 (N_13380,N_12371,N_12802);
and U13381 (N_13381,N_12551,N_12556);
and U13382 (N_13382,N_12288,N_12831);
and U13383 (N_13383,N_12828,N_12971);
or U13384 (N_13384,N_12316,N_12083);
nor U13385 (N_13385,N_12425,N_12874);
nor U13386 (N_13386,N_12497,N_12392);
and U13387 (N_13387,N_12330,N_12007);
nor U13388 (N_13388,N_12567,N_12268);
nand U13389 (N_13389,N_12541,N_12980);
xnor U13390 (N_13390,N_12837,N_12186);
nand U13391 (N_13391,N_12758,N_12047);
nand U13392 (N_13392,N_12252,N_12948);
nor U13393 (N_13393,N_12249,N_12149);
xor U13394 (N_13394,N_12285,N_12775);
nand U13395 (N_13395,N_12893,N_12671);
and U13396 (N_13396,N_12002,N_12644);
and U13397 (N_13397,N_12237,N_12794);
or U13398 (N_13398,N_12128,N_12549);
nor U13399 (N_13399,N_12811,N_12280);
or U13400 (N_13400,N_12737,N_12021);
xor U13401 (N_13401,N_12826,N_12413);
xnor U13402 (N_13402,N_12390,N_12075);
and U13403 (N_13403,N_12809,N_12055);
and U13404 (N_13404,N_12651,N_12834);
nand U13405 (N_13405,N_12404,N_12086);
xor U13406 (N_13406,N_12510,N_12934);
nor U13407 (N_13407,N_12882,N_12232);
nand U13408 (N_13408,N_12691,N_12558);
xor U13409 (N_13409,N_12173,N_12609);
nand U13410 (N_13410,N_12952,N_12059);
xor U13411 (N_13411,N_12351,N_12299);
and U13412 (N_13412,N_12174,N_12364);
xnor U13413 (N_13413,N_12539,N_12026);
nand U13414 (N_13414,N_12804,N_12722);
xnor U13415 (N_13415,N_12854,N_12415);
nand U13416 (N_13416,N_12423,N_12769);
nand U13417 (N_13417,N_12733,N_12825);
and U13418 (N_13418,N_12282,N_12734);
and U13419 (N_13419,N_12208,N_12457);
nor U13420 (N_13420,N_12053,N_12747);
and U13421 (N_13421,N_12454,N_12290);
nor U13422 (N_13422,N_12420,N_12009);
nor U13423 (N_13423,N_12024,N_12593);
and U13424 (N_13424,N_12519,N_12890);
xor U13425 (N_13425,N_12572,N_12062);
xnor U13426 (N_13426,N_12094,N_12533);
nand U13427 (N_13427,N_12740,N_12027);
nand U13428 (N_13428,N_12729,N_12597);
and U13429 (N_13429,N_12763,N_12667);
or U13430 (N_13430,N_12145,N_12191);
nand U13431 (N_13431,N_12286,N_12664);
nand U13432 (N_13432,N_12649,N_12764);
or U13433 (N_13433,N_12748,N_12408);
or U13434 (N_13434,N_12116,N_12843);
or U13435 (N_13435,N_12133,N_12314);
nor U13436 (N_13436,N_12292,N_12361);
and U13437 (N_13437,N_12950,N_12559);
xnor U13438 (N_13438,N_12291,N_12565);
and U13439 (N_13439,N_12944,N_12792);
or U13440 (N_13440,N_12870,N_12591);
and U13441 (N_13441,N_12460,N_12092);
nor U13442 (N_13442,N_12321,N_12933);
nor U13443 (N_13443,N_12111,N_12337);
nand U13444 (N_13444,N_12341,N_12356);
nand U13445 (N_13445,N_12505,N_12552);
xor U13446 (N_13446,N_12584,N_12897);
or U13447 (N_13447,N_12320,N_12765);
or U13448 (N_13448,N_12203,N_12973);
nor U13449 (N_13449,N_12385,N_12526);
xor U13450 (N_13450,N_12896,N_12407);
xor U13451 (N_13451,N_12899,N_12439);
nand U13452 (N_13452,N_12786,N_12300);
and U13453 (N_13453,N_12904,N_12338);
nor U13454 (N_13454,N_12631,N_12815);
nor U13455 (N_13455,N_12275,N_12114);
and U13456 (N_13456,N_12931,N_12583);
xnor U13457 (N_13457,N_12311,N_12349);
nand U13458 (N_13458,N_12257,N_12905);
nor U13459 (N_13459,N_12477,N_12694);
nand U13460 (N_13460,N_12192,N_12304);
nor U13461 (N_13461,N_12669,N_12736);
nor U13462 (N_13462,N_12643,N_12782);
nand U13463 (N_13463,N_12777,N_12666);
xnor U13464 (N_13464,N_12842,N_12847);
nor U13465 (N_13465,N_12207,N_12416);
or U13466 (N_13466,N_12755,N_12887);
xor U13467 (N_13467,N_12078,N_12495);
xnor U13468 (N_13468,N_12525,N_12119);
nor U13469 (N_13469,N_12881,N_12932);
xor U13470 (N_13470,N_12229,N_12472);
nand U13471 (N_13471,N_12983,N_12557);
nor U13472 (N_13472,N_12277,N_12211);
xnor U13473 (N_13473,N_12602,N_12963);
or U13474 (N_13474,N_12781,N_12164);
or U13475 (N_13475,N_12717,N_12488);
nand U13476 (N_13476,N_12523,N_12639);
and U13477 (N_13477,N_12545,N_12307);
and U13478 (N_13478,N_12650,N_12115);
nor U13479 (N_13479,N_12381,N_12670);
nor U13480 (N_13480,N_12260,N_12297);
nor U13481 (N_13481,N_12573,N_12410);
nor U13482 (N_13482,N_12793,N_12006);
xor U13483 (N_13483,N_12724,N_12701);
and U13484 (N_13484,N_12443,N_12156);
nand U13485 (N_13485,N_12819,N_12867);
and U13486 (N_13486,N_12563,N_12188);
xor U13487 (N_13487,N_12935,N_12535);
xnor U13488 (N_13488,N_12928,N_12376);
and U13489 (N_13489,N_12267,N_12520);
nor U13490 (N_13490,N_12536,N_12688);
or U13491 (N_13491,N_12625,N_12640);
nand U13492 (N_13492,N_12054,N_12065);
and U13493 (N_13493,N_12365,N_12621);
nand U13494 (N_13494,N_12101,N_12787);
or U13495 (N_13495,N_12768,N_12753);
and U13496 (N_13496,N_12157,N_12976);
or U13497 (N_13497,N_12220,N_12043);
and U13498 (N_13498,N_12475,N_12020);
nor U13499 (N_13499,N_12970,N_12919);
and U13500 (N_13500,N_12593,N_12746);
nor U13501 (N_13501,N_12084,N_12224);
nor U13502 (N_13502,N_12917,N_12766);
or U13503 (N_13503,N_12032,N_12717);
and U13504 (N_13504,N_12764,N_12028);
and U13505 (N_13505,N_12170,N_12816);
and U13506 (N_13506,N_12866,N_12142);
nand U13507 (N_13507,N_12779,N_12473);
and U13508 (N_13508,N_12071,N_12105);
nor U13509 (N_13509,N_12001,N_12343);
and U13510 (N_13510,N_12967,N_12562);
or U13511 (N_13511,N_12508,N_12778);
nand U13512 (N_13512,N_12240,N_12576);
nor U13513 (N_13513,N_12432,N_12504);
and U13514 (N_13514,N_12133,N_12325);
and U13515 (N_13515,N_12913,N_12344);
nor U13516 (N_13516,N_12574,N_12279);
or U13517 (N_13517,N_12401,N_12392);
nor U13518 (N_13518,N_12555,N_12500);
or U13519 (N_13519,N_12731,N_12460);
and U13520 (N_13520,N_12850,N_12778);
and U13521 (N_13521,N_12037,N_12083);
or U13522 (N_13522,N_12854,N_12908);
xor U13523 (N_13523,N_12808,N_12768);
xnor U13524 (N_13524,N_12406,N_12278);
or U13525 (N_13525,N_12315,N_12636);
nand U13526 (N_13526,N_12981,N_12517);
xnor U13527 (N_13527,N_12800,N_12606);
and U13528 (N_13528,N_12034,N_12422);
or U13529 (N_13529,N_12323,N_12534);
xor U13530 (N_13530,N_12811,N_12511);
and U13531 (N_13531,N_12116,N_12104);
nand U13532 (N_13532,N_12842,N_12298);
nor U13533 (N_13533,N_12143,N_12734);
and U13534 (N_13534,N_12502,N_12762);
nor U13535 (N_13535,N_12175,N_12308);
nand U13536 (N_13536,N_12672,N_12434);
and U13537 (N_13537,N_12854,N_12056);
and U13538 (N_13538,N_12108,N_12687);
nor U13539 (N_13539,N_12658,N_12229);
nand U13540 (N_13540,N_12298,N_12683);
nor U13541 (N_13541,N_12479,N_12050);
nand U13542 (N_13542,N_12573,N_12767);
xnor U13543 (N_13543,N_12661,N_12464);
nor U13544 (N_13544,N_12548,N_12086);
nor U13545 (N_13545,N_12900,N_12116);
nand U13546 (N_13546,N_12009,N_12144);
and U13547 (N_13547,N_12559,N_12709);
nand U13548 (N_13548,N_12786,N_12393);
and U13549 (N_13549,N_12639,N_12798);
or U13550 (N_13550,N_12845,N_12013);
or U13551 (N_13551,N_12413,N_12773);
or U13552 (N_13552,N_12837,N_12875);
xor U13553 (N_13553,N_12944,N_12563);
xnor U13554 (N_13554,N_12745,N_12395);
and U13555 (N_13555,N_12862,N_12478);
nand U13556 (N_13556,N_12636,N_12329);
xnor U13557 (N_13557,N_12854,N_12645);
nand U13558 (N_13558,N_12947,N_12572);
xor U13559 (N_13559,N_12583,N_12733);
xor U13560 (N_13560,N_12281,N_12482);
xor U13561 (N_13561,N_12999,N_12412);
and U13562 (N_13562,N_12124,N_12375);
nand U13563 (N_13563,N_12022,N_12235);
nor U13564 (N_13564,N_12338,N_12595);
xnor U13565 (N_13565,N_12648,N_12286);
xnor U13566 (N_13566,N_12297,N_12437);
xnor U13567 (N_13567,N_12067,N_12073);
or U13568 (N_13568,N_12849,N_12401);
xnor U13569 (N_13569,N_12556,N_12920);
nand U13570 (N_13570,N_12262,N_12069);
or U13571 (N_13571,N_12430,N_12886);
and U13572 (N_13572,N_12762,N_12558);
or U13573 (N_13573,N_12804,N_12876);
or U13574 (N_13574,N_12422,N_12244);
nor U13575 (N_13575,N_12335,N_12716);
or U13576 (N_13576,N_12484,N_12336);
xor U13577 (N_13577,N_12075,N_12010);
nand U13578 (N_13578,N_12667,N_12135);
and U13579 (N_13579,N_12638,N_12707);
or U13580 (N_13580,N_12048,N_12518);
xnor U13581 (N_13581,N_12160,N_12465);
xor U13582 (N_13582,N_12494,N_12846);
nand U13583 (N_13583,N_12414,N_12643);
and U13584 (N_13584,N_12367,N_12300);
and U13585 (N_13585,N_12619,N_12851);
nor U13586 (N_13586,N_12095,N_12371);
or U13587 (N_13587,N_12244,N_12829);
nor U13588 (N_13588,N_12058,N_12083);
and U13589 (N_13589,N_12630,N_12465);
nand U13590 (N_13590,N_12926,N_12658);
nand U13591 (N_13591,N_12146,N_12705);
and U13592 (N_13592,N_12010,N_12369);
nor U13593 (N_13593,N_12034,N_12610);
nand U13594 (N_13594,N_12511,N_12633);
nand U13595 (N_13595,N_12056,N_12618);
and U13596 (N_13596,N_12498,N_12024);
nand U13597 (N_13597,N_12966,N_12586);
or U13598 (N_13598,N_12285,N_12276);
and U13599 (N_13599,N_12798,N_12184);
or U13600 (N_13600,N_12800,N_12378);
nor U13601 (N_13601,N_12939,N_12643);
and U13602 (N_13602,N_12888,N_12703);
nor U13603 (N_13603,N_12578,N_12400);
xor U13604 (N_13604,N_12220,N_12426);
xor U13605 (N_13605,N_12484,N_12601);
nand U13606 (N_13606,N_12894,N_12849);
nand U13607 (N_13607,N_12809,N_12906);
nand U13608 (N_13608,N_12428,N_12045);
nand U13609 (N_13609,N_12360,N_12023);
or U13610 (N_13610,N_12805,N_12038);
and U13611 (N_13611,N_12423,N_12741);
xnor U13612 (N_13612,N_12956,N_12688);
and U13613 (N_13613,N_12865,N_12448);
nand U13614 (N_13614,N_12092,N_12725);
xnor U13615 (N_13615,N_12134,N_12603);
nor U13616 (N_13616,N_12567,N_12721);
and U13617 (N_13617,N_12024,N_12565);
xor U13618 (N_13618,N_12663,N_12703);
nand U13619 (N_13619,N_12754,N_12110);
nor U13620 (N_13620,N_12543,N_12546);
xnor U13621 (N_13621,N_12037,N_12575);
nor U13622 (N_13622,N_12079,N_12903);
nor U13623 (N_13623,N_12267,N_12314);
nand U13624 (N_13624,N_12355,N_12165);
nor U13625 (N_13625,N_12106,N_12793);
and U13626 (N_13626,N_12692,N_12857);
and U13627 (N_13627,N_12842,N_12767);
nor U13628 (N_13628,N_12674,N_12859);
nor U13629 (N_13629,N_12948,N_12644);
xnor U13630 (N_13630,N_12068,N_12770);
xor U13631 (N_13631,N_12181,N_12178);
nand U13632 (N_13632,N_12049,N_12663);
nor U13633 (N_13633,N_12185,N_12871);
nor U13634 (N_13634,N_12237,N_12979);
or U13635 (N_13635,N_12041,N_12678);
nor U13636 (N_13636,N_12065,N_12797);
xor U13637 (N_13637,N_12772,N_12960);
nor U13638 (N_13638,N_12218,N_12337);
xor U13639 (N_13639,N_12487,N_12644);
nand U13640 (N_13640,N_12248,N_12002);
and U13641 (N_13641,N_12123,N_12928);
nor U13642 (N_13642,N_12135,N_12320);
nor U13643 (N_13643,N_12763,N_12666);
nor U13644 (N_13644,N_12349,N_12375);
or U13645 (N_13645,N_12144,N_12810);
and U13646 (N_13646,N_12145,N_12889);
or U13647 (N_13647,N_12545,N_12223);
and U13648 (N_13648,N_12272,N_12028);
nor U13649 (N_13649,N_12383,N_12574);
and U13650 (N_13650,N_12047,N_12597);
nor U13651 (N_13651,N_12992,N_12002);
or U13652 (N_13652,N_12933,N_12110);
and U13653 (N_13653,N_12393,N_12559);
xor U13654 (N_13654,N_12044,N_12393);
xor U13655 (N_13655,N_12733,N_12599);
nand U13656 (N_13656,N_12763,N_12460);
nor U13657 (N_13657,N_12315,N_12264);
nor U13658 (N_13658,N_12156,N_12499);
nor U13659 (N_13659,N_12058,N_12615);
or U13660 (N_13660,N_12263,N_12524);
xor U13661 (N_13661,N_12575,N_12965);
nand U13662 (N_13662,N_12606,N_12157);
or U13663 (N_13663,N_12391,N_12936);
nand U13664 (N_13664,N_12093,N_12875);
or U13665 (N_13665,N_12747,N_12162);
nor U13666 (N_13666,N_12348,N_12128);
and U13667 (N_13667,N_12967,N_12932);
nand U13668 (N_13668,N_12732,N_12272);
and U13669 (N_13669,N_12481,N_12138);
xor U13670 (N_13670,N_12779,N_12486);
and U13671 (N_13671,N_12531,N_12393);
nand U13672 (N_13672,N_12840,N_12381);
nand U13673 (N_13673,N_12574,N_12381);
or U13674 (N_13674,N_12284,N_12808);
nor U13675 (N_13675,N_12218,N_12735);
nand U13676 (N_13676,N_12901,N_12344);
and U13677 (N_13677,N_12351,N_12978);
nand U13678 (N_13678,N_12926,N_12691);
nand U13679 (N_13679,N_12231,N_12779);
nor U13680 (N_13680,N_12669,N_12761);
or U13681 (N_13681,N_12123,N_12514);
and U13682 (N_13682,N_12049,N_12183);
nor U13683 (N_13683,N_12528,N_12199);
or U13684 (N_13684,N_12295,N_12331);
nand U13685 (N_13685,N_12341,N_12737);
xnor U13686 (N_13686,N_12325,N_12050);
and U13687 (N_13687,N_12652,N_12424);
nand U13688 (N_13688,N_12814,N_12910);
nand U13689 (N_13689,N_12023,N_12286);
xnor U13690 (N_13690,N_12334,N_12402);
xor U13691 (N_13691,N_12334,N_12740);
nor U13692 (N_13692,N_12859,N_12028);
nor U13693 (N_13693,N_12732,N_12253);
xor U13694 (N_13694,N_12956,N_12614);
or U13695 (N_13695,N_12685,N_12251);
and U13696 (N_13696,N_12575,N_12317);
and U13697 (N_13697,N_12704,N_12001);
nand U13698 (N_13698,N_12528,N_12359);
nand U13699 (N_13699,N_12400,N_12641);
xor U13700 (N_13700,N_12247,N_12394);
or U13701 (N_13701,N_12564,N_12385);
xnor U13702 (N_13702,N_12537,N_12292);
or U13703 (N_13703,N_12516,N_12584);
nor U13704 (N_13704,N_12829,N_12205);
nand U13705 (N_13705,N_12190,N_12836);
nor U13706 (N_13706,N_12232,N_12984);
xnor U13707 (N_13707,N_12743,N_12854);
and U13708 (N_13708,N_12132,N_12028);
xnor U13709 (N_13709,N_12589,N_12952);
nor U13710 (N_13710,N_12354,N_12399);
nor U13711 (N_13711,N_12437,N_12144);
nor U13712 (N_13712,N_12315,N_12113);
nor U13713 (N_13713,N_12989,N_12841);
or U13714 (N_13714,N_12543,N_12129);
xor U13715 (N_13715,N_12083,N_12555);
xnor U13716 (N_13716,N_12692,N_12108);
xnor U13717 (N_13717,N_12142,N_12589);
nor U13718 (N_13718,N_12119,N_12825);
and U13719 (N_13719,N_12983,N_12893);
nand U13720 (N_13720,N_12491,N_12992);
or U13721 (N_13721,N_12666,N_12235);
nand U13722 (N_13722,N_12900,N_12719);
xor U13723 (N_13723,N_12026,N_12405);
and U13724 (N_13724,N_12630,N_12494);
or U13725 (N_13725,N_12948,N_12766);
xor U13726 (N_13726,N_12796,N_12115);
nor U13727 (N_13727,N_12541,N_12003);
xnor U13728 (N_13728,N_12094,N_12526);
and U13729 (N_13729,N_12577,N_12172);
nand U13730 (N_13730,N_12524,N_12990);
xor U13731 (N_13731,N_12905,N_12220);
nor U13732 (N_13732,N_12195,N_12542);
and U13733 (N_13733,N_12469,N_12145);
or U13734 (N_13734,N_12542,N_12132);
nor U13735 (N_13735,N_12474,N_12267);
xnor U13736 (N_13736,N_12909,N_12668);
nand U13737 (N_13737,N_12092,N_12260);
and U13738 (N_13738,N_12974,N_12894);
or U13739 (N_13739,N_12614,N_12171);
and U13740 (N_13740,N_12133,N_12937);
or U13741 (N_13741,N_12999,N_12957);
and U13742 (N_13742,N_12035,N_12136);
or U13743 (N_13743,N_12042,N_12841);
nor U13744 (N_13744,N_12325,N_12436);
nand U13745 (N_13745,N_12636,N_12648);
nand U13746 (N_13746,N_12209,N_12013);
xnor U13747 (N_13747,N_12387,N_12677);
and U13748 (N_13748,N_12977,N_12956);
nand U13749 (N_13749,N_12227,N_12246);
nor U13750 (N_13750,N_12369,N_12954);
nand U13751 (N_13751,N_12043,N_12856);
and U13752 (N_13752,N_12006,N_12151);
xnor U13753 (N_13753,N_12712,N_12185);
xnor U13754 (N_13754,N_12050,N_12000);
or U13755 (N_13755,N_12126,N_12108);
nor U13756 (N_13756,N_12359,N_12678);
nand U13757 (N_13757,N_12134,N_12060);
nor U13758 (N_13758,N_12285,N_12736);
or U13759 (N_13759,N_12849,N_12621);
or U13760 (N_13760,N_12690,N_12088);
nand U13761 (N_13761,N_12377,N_12785);
or U13762 (N_13762,N_12103,N_12324);
nand U13763 (N_13763,N_12359,N_12249);
nand U13764 (N_13764,N_12069,N_12033);
or U13765 (N_13765,N_12129,N_12900);
xor U13766 (N_13766,N_12353,N_12256);
nand U13767 (N_13767,N_12109,N_12722);
nand U13768 (N_13768,N_12398,N_12099);
nor U13769 (N_13769,N_12780,N_12320);
and U13770 (N_13770,N_12040,N_12833);
nor U13771 (N_13771,N_12559,N_12819);
nor U13772 (N_13772,N_12861,N_12311);
xor U13773 (N_13773,N_12312,N_12724);
nor U13774 (N_13774,N_12720,N_12693);
nand U13775 (N_13775,N_12389,N_12193);
nand U13776 (N_13776,N_12084,N_12534);
and U13777 (N_13777,N_12217,N_12868);
and U13778 (N_13778,N_12912,N_12278);
xor U13779 (N_13779,N_12569,N_12742);
nor U13780 (N_13780,N_12053,N_12026);
or U13781 (N_13781,N_12014,N_12257);
nor U13782 (N_13782,N_12478,N_12922);
xor U13783 (N_13783,N_12529,N_12640);
and U13784 (N_13784,N_12291,N_12601);
or U13785 (N_13785,N_12274,N_12163);
and U13786 (N_13786,N_12924,N_12119);
xnor U13787 (N_13787,N_12196,N_12784);
nand U13788 (N_13788,N_12193,N_12785);
and U13789 (N_13789,N_12310,N_12468);
xnor U13790 (N_13790,N_12511,N_12461);
nor U13791 (N_13791,N_12955,N_12624);
nor U13792 (N_13792,N_12551,N_12823);
xnor U13793 (N_13793,N_12895,N_12288);
nor U13794 (N_13794,N_12986,N_12902);
xor U13795 (N_13795,N_12208,N_12511);
xor U13796 (N_13796,N_12460,N_12961);
nand U13797 (N_13797,N_12611,N_12685);
or U13798 (N_13798,N_12115,N_12018);
nand U13799 (N_13799,N_12062,N_12063);
or U13800 (N_13800,N_12890,N_12221);
nand U13801 (N_13801,N_12789,N_12503);
nand U13802 (N_13802,N_12568,N_12390);
nor U13803 (N_13803,N_12348,N_12041);
nor U13804 (N_13804,N_12484,N_12016);
nor U13805 (N_13805,N_12360,N_12016);
or U13806 (N_13806,N_12633,N_12075);
nor U13807 (N_13807,N_12960,N_12443);
nand U13808 (N_13808,N_12528,N_12953);
or U13809 (N_13809,N_12445,N_12603);
xnor U13810 (N_13810,N_12044,N_12469);
nand U13811 (N_13811,N_12777,N_12655);
nor U13812 (N_13812,N_12175,N_12568);
or U13813 (N_13813,N_12951,N_12343);
nand U13814 (N_13814,N_12819,N_12110);
nor U13815 (N_13815,N_12097,N_12955);
nand U13816 (N_13816,N_12347,N_12546);
nor U13817 (N_13817,N_12067,N_12769);
or U13818 (N_13818,N_12587,N_12853);
nand U13819 (N_13819,N_12922,N_12767);
and U13820 (N_13820,N_12375,N_12609);
nor U13821 (N_13821,N_12048,N_12808);
nand U13822 (N_13822,N_12198,N_12181);
nor U13823 (N_13823,N_12241,N_12287);
and U13824 (N_13824,N_12235,N_12268);
nand U13825 (N_13825,N_12303,N_12493);
or U13826 (N_13826,N_12343,N_12809);
xor U13827 (N_13827,N_12566,N_12407);
nand U13828 (N_13828,N_12287,N_12135);
xnor U13829 (N_13829,N_12137,N_12503);
or U13830 (N_13830,N_12945,N_12739);
nor U13831 (N_13831,N_12316,N_12439);
and U13832 (N_13832,N_12723,N_12799);
and U13833 (N_13833,N_12834,N_12447);
and U13834 (N_13834,N_12425,N_12327);
nand U13835 (N_13835,N_12916,N_12312);
xnor U13836 (N_13836,N_12856,N_12485);
xnor U13837 (N_13837,N_12481,N_12975);
nor U13838 (N_13838,N_12466,N_12567);
nor U13839 (N_13839,N_12793,N_12552);
nor U13840 (N_13840,N_12481,N_12414);
nor U13841 (N_13841,N_12528,N_12654);
nor U13842 (N_13842,N_12840,N_12590);
xnor U13843 (N_13843,N_12245,N_12230);
nor U13844 (N_13844,N_12151,N_12866);
nor U13845 (N_13845,N_12733,N_12093);
and U13846 (N_13846,N_12009,N_12014);
or U13847 (N_13847,N_12005,N_12857);
or U13848 (N_13848,N_12379,N_12879);
or U13849 (N_13849,N_12528,N_12464);
xnor U13850 (N_13850,N_12333,N_12914);
nor U13851 (N_13851,N_12870,N_12884);
and U13852 (N_13852,N_12433,N_12875);
nor U13853 (N_13853,N_12957,N_12570);
xor U13854 (N_13854,N_12946,N_12256);
nor U13855 (N_13855,N_12658,N_12422);
and U13856 (N_13856,N_12113,N_12064);
nor U13857 (N_13857,N_12450,N_12548);
or U13858 (N_13858,N_12900,N_12759);
nor U13859 (N_13859,N_12190,N_12789);
or U13860 (N_13860,N_12083,N_12397);
and U13861 (N_13861,N_12600,N_12046);
nand U13862 (N_13862,N_12402,N_12932);
nor U13863 (N_13863,N_12418,N_12104);
and U13864 (N_13864,N_12589,N_12157);
or U13865 (N_13865,N_12029,N_12336);
and U13866 (N_13866,N_12559,N_12883);
nor U13867 (N_13867,N_12800,N_12818);
nand U13868 (N_13868,N_12474,N_12333);
xor U13869 (N_13869,N_12881,N_12383);
nand U13870 (N_13870,N_12836,N_12764);
nand U13871 (N_13871,N_12380,N_12372);
or U13872 (N_13872,N_12871,N_12513);
nor U13873 (N_13873,N_12072,N_12947);
xor U13874 (N_13874,N_12413,N_12070);
or U13875 (N_13875,N_12945,N_12588);
xnor U13876 (N_13876,N_12555,N_12655);
or U13877 (N_13877,N_12602,N_12698);
nand U13878 (N_13878,N_12322,N_12644);
and U13879 (N_13879,N_12226,N_12731);
and U13880 (N_13880,N_12382,N_12559);
and U13881 (N_13881,N_12477,N_12883);
xor U13882 (N_13882,N_12866,N_12924);
nand U13883 (N_13883,N_12816,N_12847);
nor U13884 (N_13884,N_12317,N_12875);
and U13885 (N_13885,N_12258,N_12400);
or U13886 (N_13886,N_12620,N_12904);
xnor U13887 (N_13887,N_12033,N_12238);
nand U13888 (N_13888,N_12226,N_12108);
xnor U13889 (N_13889,N_12447,N_12247);
nor U13890 (N_13890,N_12292,N_12968);
xnor U13891 (N_13891,N_12155,N_12701);
xnor U13892 (N_13892,N_12712,N_12130);
nor U13893 (N_13893,N_12142,N_12598);
or U13894 (N_13894,N_12464,N_12249);
or U13895 (N_13895,N_12362,N_12110);
and U13896 (N_13896,N_12453,N_12560);
or U13897 (N_13897,N_12327,N_12379);
nor U13898 (N_13898,N_12029,N_12664);
or U13899 (N_13899,N_12861,N_12255);
or U13900 (N_13900,N_12071,N_12747);
and U13901 (N_13901,N_12956,N_12444);
xor U13902 (N_13902,N_12102,N_12578);
and U13903 (N_13903,N_12671,N_12062);
nand U13904 (N_13904,N_12427,N_12186);
xor U13905 (N_13905,N_12159,N_12016);
xnor U13906 (N_13906,N_12281,N_12296);
and U13907 (N_13907,N_12451,N_12959);
or U13908 (N_13908,N_12304,N_12136);
or U13909 (N_13909,N_12614,N_12248);
nor U13910 (N_13910,N_12818,N_12156);
nor U13911 (N_13911,N_12786,N_12931);
nor U13912 (N_13912,N_12881,N_12592);
nor U13913 (N_13913,N_12378,N_12833);
nand U13914 (N_13914,N_12498,N_12833);
nand U13915 (N_13915,N_12801,N_12473);
or U13916 (N_13916,N_12848,N_12455);
or U13917 (N_13917,N_12248,N_12875);
nor U13918 (N_13918,N_12573,N_12908);
or U13919 (N_13919,N_12495,N_12883);
or U13920 (N_13920,N_12918,N_12811);
nor U13921 (N_13921,N_12795,N_12920);
and U13922 (N_13922,N_12232,N_12896);
or U13923 (N_13923,N_12742,N_12849);
xnor U13924 (N_13924,N_12655,N_12685);
and U13925 (N_13925,N_12005,N_12783);
nand U13926 (N_13926,N_12437,N_12942);
nor U13927 (N_13927,N_12884,N_12504);
nand U13928 (N_13928,N_12843,N_12367);
nor U13929 (N_13929,N_12921,N_12159);
and U13930 (N_13930,N_12870,N_12869);
and U13931 (N_13931,N_12023,N_12630);
or U13932 (N_13932,N_12486,N_12165);
or U13933 (N_13933,N_12268,N_12860);
and U13934 (N_13934,N_12948,N_12927);
nand U13935 (N_13935,N_12566,N_12355);
nor U13936 (N_13936,N_12158,N_12899);
nor U13937 (N_13937,N_12162,N_12619);
and U13938 (N_13938,N_12582,N_12558);
and U13939 (N_13939,N_12378,N_12158);
and U13940 (N_13940,N_12352,N_12224);
xor U13941 (N_13941,N_12044,N_12514);
or U13942 (N_13942,N_12106,N_12495);
nor U13943 (N_13943,N_12768,N_12258);
nor U13944 (N_13944,N_12208,N_12223);
nand U13945 (N_13945,N_12531,N_12475);
nor U13946 (N_13946,N_12183,N_12797);
nand U13947 (N_13947,N_12135,N_12322);
and U13948 (N_13948,N_12285,N_12067);
and U13949 (N_13949,N_12592,N_12164);
nor U13950 (N_13950,N_12973,N_12966);
xor U13951 (N_13951,N_12084,N_12286);
nor U13952 (N_13952,N_12887,N_12960);
nor U13953 (N_13953,N_12758,N_12305);
nand U13954 (N_13954,N_12383,N_12806);
xor U13955 (N_13955,N_12361,N_12704);
or U13956 (N_13956,N_12677,N_12870);
nand U13957 (N_13957,N_12037,N_12362);
or U13958 (N_13958,N_12984,N_12770);
xnor U13959 (N_13959,N_12031,N_12133);
nor U13960 (N_13960,N_12266,N_12472);
or U13961 (N_13961,N_12204,N_12591);
and U13962 (N_13962,N_12792,N_12759);
xor U13963 (N_13963,N_12737,N_12198);
or U13964 (N_13964,N_12011,N_12792);
xnor U13965 (N_13965,N_12715,N_12732);
xnor U13966 (N_13966,N_12079,N_12650);
xor U13967 (N_13967,N_12913,N_12935);
xor U13968 (N_13968,N_12760,N_12602);
nor U13969 (N_13969,N_12096,N_12649);
nor U13970 (N_13970,N_12576,N_12935);
or U13971 (N_13971,N_12691,N_12348);
and U13972 (N_13972,N_12350,N_12928);
xor U13973 (N_13973,N_12952,N_12673);
and U13974 (N_13974,N_12856,N_12393);
nor U13975 (N_13975,N_12728,N_12614);
and U13976 (N_13976,N_12095,N_12405);
and U13977 (N_13977,N_12125,N_12189);
and U13978 (N_13978,N_12766,N_12352);
or U13979 (N_13979,N_12425,N_12475);
xor U13980 (N_13980,N_12182,N_12008);
nor U13981 (N_13981,N_12932,N_12975);
or U13982 (N_13982,N_12836,N_12097);
nor U13983 (N_13983,N_12957,N_12689);
xnor U13984 (N_13984,N_12338,N_12705);
xnor U13985 (N_13985,N_12421,N_12948);
nor U13986 (N_13986,N_12324,N_12700);
nand U13987 (N_13987,N_12405,N_12166);
nand U13988 (N_13988,N_12867,N_12608);
or U13989 (N_13989,N_12940,N_12539);
nor U13990 (N_13990,N_12007,N_12912);
or U13991 (N_13991,N_12565,N_12750);
nand U13992 (N_13992,N_12041,N_12032);
and U13993 (N_13993,N_12498,N_12880);
nor U13994 (N_13994,N_12942,N_12628);
xnor U13995 (N_13995,N_12331,N_12461);
xor U13996 (N_13996,N_12633,N_12439);
nand U13997 (N_13997,N_12309,N_12776);
nand U13998 (N_13998,N_12967,N_12442);
nor U13999 (N_13999,N_12115,N_12779);
and U14000 (N_14000,N_13681,N_13364);
or U14001 (N_14001,N_13697,N_13657);
and U14002 (N_14002,N_13580,N_13721);
nand U14003 (N_14003,N_13074,N_13779);
and U14004 (N_14004,N_13861,N_13476);
nand U14005 (N_14005,N_13761,N_13178);
nor U14006 (N_14006,N_13749,N_13979);
nand U14007 (N_14007,N_13716,N_13319);
or U14008 (N_14008,N_13582,N_13013);
or U14009 (N_14009,N_13269,N_13594);
xnor U14010 (N_14010,N_13526,N_13070);
xor U14011 (N_14011,N_13992,N_13939);
nor U14012 (N_14012,N_13741,N_13324);
xor U14013 (N_14013,N_13776,N_13957);
and U14014 (N_14014,N_13161,N_13362);
and U14015 (N_14015,N_13900,N_13558);
nor U14016 (N_14016,N_13607,N_13296);
nand U14017 (N_14017,N_13018,N_13763);
nor U14018 (N_14018,N_13952,N_13856);
or U14019 (N_14019,N_13329,N_13976);
xnor U14020 (N_14020,N_13165,N_13214);
or U14021 (N_14021,N_13670,N_13980);
nor U14022 (N_14022,N_13897,N_13148);
or U14023 (N_14023,N_13340,N_13770);
nor U14024 (N_14024,N_13750,N_13474);
or U14025 (N_14025,N_13602,N_13513);
nor U14026 (N_14026,N_13511,N_13932);
xnor U14027 (N_14027,N_13091,N_13821);
and U14028 (N_14028,N_13272,N_13688);
and U14029 (N_14029,N_13442,N_13617);
nor U14030 (N_14030,N_13244,N_13533);
or U14031 (N_14031,N_13408,N_13982);
xnor U14032 (N_14032,N_13230,N_13392);
or U14033 (N_14033,N_13867,N_13792);
and U14034 (N_14034,N_13702,N_13133);
or U14035 (N_14035,N_13940,N_13562);
nor U14036 (N_14036,N_13935,N_13410);
xor U14037 (N_14037,N_13446,N_13514);
or U14038 (N_14038,N_13916,N_13263);
xnor U14039 (N_14039,N_13655,N_13368);
nor U14040 (N_14040,N_13960,N_13304);
nor U14041 (N_14041,N_13172,N_13220);
xnor U14042 (N_14042,N_13774,N_13287);
xor U14043 (N_14043,N_13372,N_13841);
or U14044 (N_14044,N_13644,N_13208);
and U14045 (N_14045,N_13301,N_13934);
and U14046 (N_14046,N_13496,N_13241);
xnor U14047 (N_14047,N_13394,N_13783);
and U14048 (N_14048,N_13120,N_13805);
nor U14049 (N_14049,N_13577,N_13807);
nand U14050 (N_14050,N_13699,N_13246);
xnor U14051 (N_14051,N_13522,N_13370);
nor U14052 (N_14052,N_13682,N_13633);
or U14053 (N_14053,N_13024,N_13309);
and U14054 (N_14054,N_13045,N_13405);
nand U14055 (N_14055,N_13796,N_13691);
nor U14056 (N_14056,N_13573,N_13436);
xnor U14057 (N_14057,N_13556,N_13615);
nor U14058 (N_14058,N_13316,N_13549);
nor U14059 (N_14059,N_13205,N_13618);
and U14060 (N_14060,N_13327,N_13102);
and U14061 (N_14061,N_13217,N_13253);
and U14062 (N_14062,N_13273,N_13321);
xor U14063 (N_14063,N_13833,N_13355);
nor U14064 (N_14064,N_13396,N_13781);
nand U14065 (N_14065,N_13495,N_13747);
or U14066 (N_14066,N_13733,N_13828);
nand U14067 (N_14067,N_13004,N_13970);
nand U14068 (N_14068,N_13482,N_13994);
and U14069 (N_14069,N_13213,N_13595);
or U14070 (N_14070,N_13125,N_13181);
nand U14071 (N_14071,N_13698,N_13068);
and U14072 (N_14072,N_13778,N_13515);
or U14073 (N_14073,N_13433,N_13009);
nand U14074 (N_14074,N_13664,N_13251);
and U14075 (N_14075,N_13645,N_13658);
nor U14076 (N_14076,N_13569,N_13270);
nor U14077 (N_14077,N_13059,N_13634);
and U14078 (N_14078,N_13113,N_13787);
and U14079 (N_14079,N_13249,N_13237);
xor U14080 (N_14080,N_13334,N_13744);
xnor U14081 (N_14081,N_13153,N_13336);
nand U14082 (N_14082,N_13966,N_13956);
nor U14083 (N_14083,N_13075,N_13444);
and U14084 (N_14084,N_13012,N_13837);
and U14085 (N_14085,N_13060,N_13069);
nor U14086 (N_14086,N_13568,N_13669);
nand U14087 (N_14087,N_13654,N_13748);
nand U14088 (N_14088,N_13460,N_13855);
nor U14089 (N_14089,N_13641,N_13608);
xnor U14090 (N_14090,N_13083,N_13795);
nor U14091 (N_14091,N_13583,N_13167);
xnor U14092 (N_14092,N_13693,N_13646);
xor U14093 (N_14093,N_13825,N_13192);
nand U14094 (N_14094,N_13518,N_13404);
nor U14095 (N_14095,N_13660,N_13988);
and U14096 (N_14096,N_13938,N_13008);
xor U14097 (N_14097,N_13930,N_13754);
nand U14098 (N_14098,N_13739,N_13708);
nor U14099 (N_14099,N_13772,N_13676);
and U14100 (N_14100,N_13285,N_13160);
nand U14101 (N_14101,N_13530,N_13485);
xnor U14102 (N_14102,N_13414,N_13824);
or U14103 (N_14103,N_13677,N_13949);
and U14104 (N_14104,N_13435,N_13337);
nor U14105 (N_14105,N_13948,N_13943);
or U14106 (N_14106,N_13159,N_13672);
or U14107 (N_14107,N_13603,N_13374);
xor U14108 (N_14108,N_13995,N_13508);
nand U14109 (N_14109,N_13894,N_13944);
and U14110 (N_14110,N_13310,N_13308);
nand U14111 (N_14111,N_13490,N_13042);
nand U14112 (N_14112,N_13541,N_13713);
or U14113 (N_14113,N_13211,N_13001);
nor U14114 (N_14114,N_13542,N_13601);
or U14115 (N_14115,N_13517,N_13202);
nor U14116 (N_14116,N_13844,N_13576);
or U14117 (N_14117,N_13946,N_13107);
nand U14118 (N_14118,N_13984,N_13111);
xor U14119 (N_14119,N_13743,N_13061);
nor U14120 (N_14120,N_13348,N_13563);
nand U14121 (N_14121,N_13371,N_13027);
xor U14122 (N_14122,N_13328,N_13432);
nor U14123 (N_14123,N_13416,N_13357);
xnor U14124 (N_14124,N_13135,N_13604);
and U14125 (N_14125,N_13891,N_13250);
xor U14126 (N_14126,N_13302,N_13020);
nor U14127 (N_14127,N_13499,N_13006);
nand U14128 (N_14128,N_13144,N_13265);
nand U14129 (N_14129,N_13430,N_13489);
and U14130 (N_14130,N_13959,N_13598);
nor U14131 (N_14131,N_13458,N_13768);
xnor U14132 (N_14132,N_13406,N_13315);
nor U14133 (N_14133,N_13890,N_13011);
nand U14134 (N_14134,N_13806,N_13369);
or U14135 (N_14135,N_13906,N_13917);
xor U14136 (N_14136,N_13876,N_13740);
or U14137 (N_14137,N_13142,N_13239);
and U14138 (N_14138,N_13438,N_13375);
nor U14139 (N_14139,N_13636,N_13794);
nand U14140 (N_14140,N_13479,N_13629);
xor U14141 (N_14141,N_13424,N_13464);
or U14142 (N_14142,N_13929,N_13950);
nor U14143 (N_14143,N_13170,N_13437);
xor U14144 (N_14144,N_13227,N_13997);
nor U14145 (N_14145,N_13579,N_13343);
and U14146 (N_14146,N_13784,N_13145);
xnor U14147 (N_14147,N_13463,N_13745);
xnor U14148 (N_14148,N_13073,N_13233);
and U14149 (N_14149,N_13502,N_13650);
nand U14150 (N_14150,N_13860,N_13863);
nand U14151 (N_14151,N_13840,N_13986);
xnor U14152 (N_14152,N_13184,N_13290);
and U14153 (N_14153,N_13643,N_13961);
nor U14154 (N_14154,N_13467,N_13168);
xor U14155 (N_14155,N_13095,N_13921);
nor U14156 (N_14156,N_13468,N_13183);
xor U14157 (N_14157,N_13570,N_13387);
or U14158 (N_14158,N_13667,N_13880);
or U14159 (N_14159,N_13690,N_13581);
nand U14160 (N_14160,N_13675,N_13225);
and U14161 (N_14161,N_13236,N_13320);
nand U14162 (N_14162,N_13852,N_13235);
or U14163 (N_14163,N_13866,N_13695);
nor U14164 (N_14164,N_13257,N_13622);
nand U14165 (N_14165,N_13928,N_13299);
nor U14166 (N_14166,N_13140,N_13311);
xnor U14167 (N_14167,N_13947,N_13462);
nand U14168 (N_14168,N_13922,N_13864);
nor U14169 (N_14169,N_13481,N_13788);
and U14170 (N_14170,N_13051,N_13187);
nor U14171 (N_14171,N_13103,N_13224);
and U14172 (N_14172,N_13497,N_13516);
and U14173 (N_14173,N_13112,N_13456);
nor U14174 (N_14174,N_13386,N_13560);
nand U14175 (N_14175,N_13535,N_13030);
nor U14176 (N_14176,N_13726,N_13358);
xnor U14177 (N_14177,N_13108,N_13593);
or U14178 (N_14178,N_13157,N_13600);
and U14179 (N_14179,N_13751,N_13494);
nand U14180 (N_14180,N_13710,N_13123);
and U14181 (N_14181,N_13247,N_13663);
or U14182 (N_14182,N_13367,N_13899);
and U14183 (N_14183,N_13131,N_13684);
and U14184 (N_14184,N_13293,N_13962);
or U14185 (N_14185,N_13245,N_13313);
xnor U14186 (N_14186,N_13835,N_13912);
and U14187 (N_14187,N_13551,N_13908);
and U14188 (N_14188,N_13647,N_13762);
xnor U14189 (N_14189,N_13727,N_13640);
or U14190 (N_14190,N_13557,N_13289);
and U14191 (N_14191,N_13326,N_13126);
xor U14192 (N_14192,N_13847,N_13548);
and U14193 (N_14193,N_13280,N_13810);
nor U14194 (N_14194,N_13441,N_13661);
nor U14195 (N_14195,N_13440,N_13286);
or U14196 (N_14196,N_13469,N_13094);
nand U14197 (N_14197,N_13816,N_13127);
or U14198 (N_14198,N_13390,N_13067);
xnor U14199 (N_14199,N_13082,N_13883);
nand U14200 (N_14200,N_13199,N_13719);
and U14201 (N_14201,N_13377,N_13903);
nor U14202 (N_14202,N_13789,N_13814);
or U14203 (N_14203,N_13339,N_13700);
xor U14204 (N_14204,N_13656,N_13936);
or U14205 (N_14205,N_13543,N_13968);
nand U14206 (N_14206,N_13746,N_13879);
and U14207 (N_14207,N_13521,N_13905);
nor U14208 (N_14208,N_13483,N_13283);
xor U14209 (N_14209,N_13064,N_13201);
nand U14210 (N_14210,N_13207,N_13473);
xnor U14211 (N_14211,N_13854,N_13033);
nor U14212 (N_14212,N_13356,N_13753);
and U14213 (N_14213,N_13063,N_13717);
xnor U14214 (N_14214,N_13491,N_13705);
nand U14215 (N_14215,N_13252,N_13799);
nor U14216 (N_14216,N_13775,N_13758);
xnor U14217 (N_14217,N_13453,N_13134);
or U14218 (N_14218,N_13179,N_13981);
nor U14219 (N_14219,N_13016,N_13868);
xor U14220 (N_14220,N_13609,N_13545);
and U14221 (N_14221,N_13232,N_13571);
nor U14222 (N_14222,N_13097,N_13062);
nand U14223 (N_14223,N_13901,N_13418);
and U14224 (N_14224,N_13862,N_13305);
nor U14225 (N_14225,N_13941,N_13403);
xnor U14226 (N_14226,N_13471,N_13005);
and U14227 (N_14227,N_13534,N_13226);
and U14228 (N_14228,N_13706,N_13026);
and U14229 (N_14229,N_13826,N_13029);
xor U14230 (N_14230,N_13843,N_13216);
or U14231 (N_14231,N_13838,N_13010);
and U14232 (N_14232,N_13271,N_13884);
nor U14233 (N_14233,N_13223,N_13877);
and U14234 (N_14234,N_13079,N_13072);
xnor U14235 (N_14235,N_13998,N_13492);
xnor U14236 (N_14236,N_13136,N_13307);
nand U14237 (N_14237,N_13084,N_13592);
and U14238 (N_14238,N_13197,N_13722);
or U14239 (N_14239,N_13034,N_13673);
nand U14240 (N_14240,N_13365,N_13507);
nor U14241 (N_14241,N_13527,N_13605);
and U14242 (N_14242,N_13780,N_13718);
nor U14243 (N_14243,N_13574,N_13735);
or U14244 (N_14244,N_13823,N_13623);
nor U14245 (N_14245,N_13455,N_13448);
nor U14246 (N_14246,N_13206,N_13146);
and U14247 (N_14247,N_13037,N_13049);
xnor U14248 (N_14248,N_13300,N_13175);
and U14249 (N_14249,N_13459,N_13915);
or U14250 (N_14250,N_13965,N_13204);
nand U14251 (N_14251,N_13023,N_13039);
nand U14252 (N_14252,N_13141,N_13588);
xor U14253 (N_14253,N_13351,N_13550);
or U14254 (N_14254,N_13347,N_13978);
and U14255 (N_14255,N_13544,N_13873);
nor U14256 (N_14256,N_13397,N_13798);
nor U14257 (N_14257,N_13100,N_13415);
and U14258 (N_14258,N_13128,N_13532);
and U14259 (N_14259,N_13048,N_13114);
xor U14260 (N_14260,N_13118,N_13509);
or U14261 (N_14261,N_13674,N_13158);
and U14262 (N_14262,N_13383,N_13756);
nor U14263 (N_14263,N_13869,N_13282);
xnor U14264 (N_14264,N_13911,N_13830);
xnor U14265 (N_14265,N_13914,N_13683);
and U14266 (N_14266,N_13231,N_13686);
or U14267 (N_14267,N_13987,N_13931);
and U14268 (N_14268,N_13769,N_13056);
nand U14269 (N_14269,N_13427,N_13477);
and U14270 (N_14270,N_13389,N_13346);
nor U14271 (N_14271,N_13610,N_13338);
and U14272 (N_14272,N_13597,N_13065);
or U14273 (N_14273,N_13590,N_13186);
or U14274 (N_14274,N_13709,N_13361);
nor U14275 (N_14275,N_13025,N_13274);
nand U14276 (N_14276,N_13124,N_13760);
nor U14277 (N_14277,N_13606,N_13925);
nand U14278 (N_14278,N_13553,N_13344);
and U14279 (N_14279,N_13510,N_13815);
nor U14280 (N_14280,N_13439,N_13689);
and U14281 (N_14281,N_13000,N_13166);
nor U14282 (N_14282,N_13639,N_13896);
nand U14283 (N_14283,N_13564,N_13189);
and U14284 (N_14284,N_13506,N_13395);
xor U14285 (N_14285,N_13500,N_13626);
xor U14286 (N_14286,N_13391,N_13973);
nand U14287 (N_14287,N_13243,N_13625);
and U14288 (N_14288,N_13523,N_13193);
nor U14289 (N_14289,N_13555,N_13953);
nand U14290 (N_14290,N_13450,N_13993);
xnor U14291 (N_14291,N_13540,N_13528);
nor U14292 (N_14292,N_13898,N_13261);
or U14293 (N_14293,N_13017,N_13723);
or U14294 (N_14294,N_13052,N_13859);
nor U14295 (N_14295,N_13729,N_13110);
nand U14296 (N_14296,N_13565,N_13054);
and U14297 (N_14297,N_13196,N_13332);
nand U14298 (N_14298,N_13200,N_13919);
and U14299 (N_14299,N_13194,N_13714);
xnor U14300 (N_14300,N_13801,N_13417);
nor U14301 (N_14301,N_13022,N_13820);
or U14302 (N_14302,N_13384,N_13665);
nor U14303 (N_14303,N_13635,N_13266);
nor U14304 (N_14304,N_13028,N_13470);
nor U14305 (N_14305,N_13180,N_13793);
or U14306 (N_14306,N_13732,N_13771);
or U14307 (N_14307,N_13561,N_13724);
nand U14308 (N_14308,N_13267,N_13631);
nor U14309 (N_14309,N_13893,N_13933);
xnor U14310 (N_14310,N_13087,N_13923);
nand U14311 (N_14311,N_13865,N_13578);
nand U14312 (N_14312,N_13104,N_13376);
nor U14313 (N_14313,N_13611,N_13325);
nor U14314 (N_14314,N_13849,N_13425);
xnor U14315 (N_14315,N_13137,N_13198);
xor U14316 (N_14316,N_13076,N_13752);
xor U14317 (N_14317,N_13885,N_13874);
nand U14318 (N_14318,N_13501,N_13215);
and U14319 (N_14319,N_13203,N_13519);
nor U14320 (N_14320,N_13738,N_13306);
or U14321 (N_14321,N_13969,N_13575);
and U14322 (N_14322,N_13851,N_13909);
xor U14323 (N_14323,N_13057,N_13790);
nor U14324 (N_14324,N_13850,N_13164);
nand U14325 (N_14325,N_13262,N_13552);
nor U14326 (N_14326,N_13529,N_13105);
xnor U14327 (N_14327,N_13138,N_13803);
nor U14328 (N_14328,N_13407,N_13926);
and U14329 (N_14329,N_13503,N_13401);
xor U14330 (N_14330,N_13696,N_13021);
xnor U14331 (N_14331,N_13151,N_13651);
and U14332 (N_14332,N_13954,N_13971);
xnor U14333 (N_14333,N_13385,N_13685);
or U14334 (N_14334,N_13659,N_13229);
or U14335 (N_14335,N_13388,N_13451);
and U14336 (N_14336,N_13349,N_13080);
nand U14337 (N_14337,N_13742,N_13149);
or U14338 (N_14338,N_13991,N_13419);
nand U14339 (N_14339,N_13904,N_13871);
nor U14340 (N_14340,N_13380,N_13046);
and U14341 (N_14341,N_13895,N_13078);
and U14342 (N_14342,N_13572,N_13466);
and U14343 (N_14343,N_13053,N_13312);
and U14344 (N_14344,N_13791,N_13587);
nand U14345 (N_14345,N_13119,N_13209);
xnor U14346 (N_14346,N_13152,N_13295);
nand U14347 (N_14347,N_13480,N_13712);
nand U14348 (N_14348,N_13147,N_13536);
or U14349 (N_14349,N_13832,N_13129);
xnor U14350 (N_14350,N_13155,N_13730);
or U14351 (N_14351,N_13212,N_13275);
xnor U14352 (N_14352,N_13139,N_13679);
xor U14353 (N_14353,N_13122,N_13853);
or U14354 (N_14354,N_13411,N_13294);
nand U14355 (N_14355,N_13964,N_13443);
nor U14356 (N_14356,N_13447,N_13942);
nand U14357 (N_14357,N_13888,N_13003);
xor U14358 (N_14358,N_13547,N_13619);
or U14359 (N_14359,N_13802,N_13191);
and U14360 (N_14360,N_13566,N_13808);
nand U14361 (N_14361,N_13218,N_13701);
or U14362 (N_14362,N_13279,N_13678);
and U14363 (N_14363,N_13945,N_13258);
nand U14364 (N_14364,N_13278,N_13345);
and U14365 (N_14365,N_13628,N_13081);
nand U14366 (N_14366,N_13096,N_13694);
nor U14367 (N_14367,N_13627,N_13354);
and U14368 (N_14368,N_13043,N_13412);
nand U14369 (N_14369,N_13967,N_13014);
nand U14370 (N_14370,N_13333,N_13620);
or U14371 (N_14371,N_13538,N_13323);
nor U14372 (N_14372,N_13420,N_13413);
xnor U14373 (N_14373,N_13546,N_13379);
xnor U14374 (N_14374,N_13638,N_13363);
and U14375 (N_14375,N_13298,N_13586);
and U14376 (N_14376,N_13019,N_13238);
nor U14377 (N_14377,N_13101,N_13445);
nand U14378 (N_14378,N_13281,N_13058);
and U14379 (N_14379,N_13234,N_13381);
nor U14380 (N_14380,N_13845,N_13870);
nor U14381 (N_14381,N_13350,N_13613);
and U14382 (N_14382,N_13366,N_13098);
nor U14383 (N_14383,N_13154,N_13666);
xnor U14384 (N_14384,N_13143,N_13591);
nor U14385 (N_14385,N_13637,N_13648);
and U14386 (N_14386,N_13132,N_13822);
nor U14387 (N_14387,N_13818,N_13819);
and U14388 (N_14388,N_13887,N_13150);
xor U14389 (N_14389,N_13817,N_13985);
nor U14390 (N_14390,N_13927,N_13484);
or U14391 (N_14391,N_13955,N_13452);
nand U14392 (N_14392,N_13537,N_13937);
or U14393 (N_14393,N_13121,N_13041);
nand U14394 (N_14394,N_13055,N_13878);
xor U14395 (N_14395,N_13268,N_13882);
nand U14396 (N_14396,N_13848,N_13242);
nand U14397 (N_14397,N_13765,N_13185);
or U14398 (N_14398,N_13210,N_13668);
xor U14399 (N_14399,N_13255,N_13429);
xor U14400 (N_14400,N_13800,N_13488);
or U14401 (N_14401,N_13759,N_13035);
nand U14402 (N_14402,N_13704,N_13291);
or U14403 (N_14403,N_13047,N_13090);
nor U14404 (N_14404,N_13924,N_13359);
xor U14405 (N_14405,N_13115,N_13498);
or U14406 (N_14406,N_13812,N_13222);
and U14407 (N_14407,N_13428,N_13116);
xnor U14408 (N_14408,N_13335,N_13773);
xnor U14409 (N_14409,N_13292,N_13195);
and U14410 (N_14410,N_13907,N_13260);
nor U14411 (N_14411,N_13525,N_13834);
nor U14412 (N_14412,N_13378,N_13475);
and U14413 (N_14413,N_13431,N_13177);
nand U14414 (N_14414,N_13653,N_13842);
nand U14415 (N_14415,N_13734,N_13958);
and U14416 (N_14416,N_13248,N_13512);
nand U14417 (N_14417,N_13839,N_13240);
nand U14418 (N_14418,N_13176,N_13277);
nor U14419 (N_14419,N_13093,N_13764);
nand U14420 (N_14420,N_13117,N_13188);
and U14421 (N_14421,N_13804,N_13589);
or U14422 (N_14422,N_13831,N_13303);
xnor U14423 (N_14423,N_13886,N_13813);
xnor U14424 (N_14424,N_13171,N_13989);
xnor U14425 (N_14425,N_13162,N_13652);
or U14426 (N_14426,N_13465,N_13872);
or U14427 (N_14427,N_13322,N_13777);
nand U14428 (N_14428,N_13106,N_13786);
nand U14429 (N_14429,N_13190,N_13330);
nand U14430 (N_14430,N_13554,N_13007);
nand U14431 (N_14431,N_13846,N_13360);
or U14432 (N_14432,N_13766,N_13461);
and U14433 (N_14433,N_13130,N_13757);
xor U14434 (N_14434,N_13725,N_13520);
nand U14435 (N_14435,N_13680,N_13109);
xnor U14436 (N_14436,N_13975,N_13254);
and U14437 (N_14437,N_13983,N_13472);
nor U14438 (N_14438,N_13173,N_13409);
xor U14439 (N_14439,N_13423,N_13797);
and U14440 (N_14440,N_13085,N_13297);
or U14441 (N_14441,N_13314,N_13038);
nor U14442 (N_14442,N_13918,N_13259);
or U14443 (N_14443,N_13398,N_13015);
and U14444 (N_14444,N_13221,N_13454);
nor U14445 (N_14445,N_13071,N_13858);
nor U14446 (N_14446,N_13457,N_13382);
and U14447 (N_14447,N_13531,N_13284);
nand U14448 (N_14448,N_13505,N_13352);
nor U14449 (N_14449,N_13099,N_13393);
and U14450 (N_14450,N_13827,N_13434);
nand U14451 (N_14451,N_13044,N_13031);
nand U14452 (N_14452,N_13642,N_13977);
xnor U14453 (N_14453,N_13720,N_13809);
nand U14454 (N_14454,N_13621,N_13707);
xnor U14455 (N_14455,N_13182,N_13703);
or U14456 (N_14456,N_13288,N_13077);
nand U14457 (N_14457,N_13174,N_13892);
nand U14458 (N_14458,N_13341,N_13692);
xnor U14459 (N_14459,N_13630,N_13857);
and U14460 (N_14460,N_13156,N_13228);
and U14461 (N_14461,N_13889,N_13400);
or U14462 (N_14462,N_13951,N_13920);
nor U14463 (N_14463,N_13737,N_13567);
or U14464 (N_14464,N_13317,N_13066);
xnor U14465 (N_14465,N_13486,N_13219);
nor U14466 (N_14466,N_13649,N_13032);
or U14467 (N_14467,N_13089,N_13487);
or U14468 (N_14468,N_13399,N_13913);
nor U14469 (N_14469,N_13996,N_13264);
and U14470 (N_14470,N_13002,N_13671);
xor U14471 (N_14471,N_13875,N_13811);
or U14472 (N_14472,N_13086,N_13163);
or U14473 (N_14473,N_13353,N_13999);
and U14474 (N_14474,N_13881,N_13040);
and U14475 (N_14475,N_13632,N_13599);
nor U14476 (N_14476,N_13782,N_13990);
xnor U14477 (N_14477,N_13711,N_13974);
nand U14478 (N_14478,N_13504,N_13715);
nand U14479 (N_14479,N_13836,N_13276);
or U14480 (N_14480,N_13736,N_13624);
or U14481 (N_14481,N_13421,N_13585);
nor U14482 (N_14482,N_13972,N_13036);
xor U14483 (N_14483,N_13402,N_13256);
and U14484 (N_14484,N_13614,N_13088);
and U14485 (N_14485,N_13169,N_13342);
nand U14486 (N_14486,N_13785,N_13331);
nand U14487 (N_14487,N_13092,N_13584);
nor U14488 (N_14488,N_13596,N_13373);
xnor U14489 (N_14489,N_13687,N_13616);
xor U14490 (N_14490,N_13612,N_13910);
and U14491 (N_14491,N_13829,N_13728);
and U14492 (N_14492,N_13662,N_13539);
nand U14493 (N_14493,N_13449,N_13755);
xor U14494 (N_14494,N_13478,N_13902);
or U14495 (N_14495,N_13559,N_13422);
or U14496 (N_14496,N_13050,N_13731);
and U14497 (N_14497,N_13767,N_13493);
xor U14498 (N_14498,N_13524,N_13426);
nor U14499 (N_14499,N_13963,N_13318);
xnor U14500 (N_14500,N_13114,N_13625);
and U14501 (N_14501,N_13350,N_13379);
and U14502 (N_14502,N_13984,N_13411);
xor U14503 (N_14503,N_13760,N_13221);
and U14504 (N_14504,N_13784,N_13760);
xor U14505 (N_14505,N_13672,N_13468);
xnor U14506 (N_14506,N_13915,N_13439);
nand U14507 (N_14507,N_13681,N_13853);
or U14508 (N_14508,N_13764,N_13611);
xor U14509 (N_14509,N_13983,N_13032);
nand U14510 (N_14510,N_13020,N_13632);
nand U14511 (N_14511,N_13486,N_13547);
or U14512 (N_14512,N_13435,N_13265);
nor U14513 (N_14513,N_13977,N_13589);
nor U14514 (N_14514,N_13722,N_13764);
nand U14515 (N_14515,N_13909,N_13306);
nor U14516 (N_14516,N_13021,N_13748);
and U14517 (N_14517,N_13028,N_13787);
and U14518 (N_14518,N_13519,N_13431);
and U14519 (N_14519,N_13420,N_13968);
nor U14520 (N_14520,N_13377,N_13467);
and U14521 (N_14521,N_13049,N_13096);
nand U14522 (N_14522,N_13361,N_13676);
nor U14523 (N_14523,N_13148,N_13758);
nand U14524 (N_14524,N_13639,N_13727);
nand U14525 (N_14525,N_13153,N_13371);
nand U14526 (N_14526,N_13384,N_13972);
nor U14527 (N_14527,N_13584,N_13028);
or U14528 (N_14528,N_13955,N_13580);
or U14529 (N_14529,N_13478,N_13477);
or U14530 (N_14530,N_13819,N_13319);
nor U14531 (N_14531,N_13498,N_13655);
or U14532 (N_14532,N_13447,N_13070);
nand U14533 (N_14533,N_13897,N_13687);
nand U14534 (N_14534,N_13240,N_13822);
or U14535 (N_14535,N_13091,N_13038);
xnor U14536 (N_14536,N_13630,N_13984);
nand U14537 (N_14537,N_13145,N_13901);
and U14538 (N_14538,N_13302,N_13099);
nand U14539 (N_14539,N_13045,N_13572);
nand U14540 (N_14540,N_13435,N_13002);
nand U14541 (N_14541,N_13582,N_13489);
nand U14542 (N_14542,N_13040,N_13279);
or U14543 (N_14543,N_13120,N_13737);
nand U14544 (N_14544,N_13768,N_13386);
xor U14545 (N_14545,N_13819,N_13045);
or U14546 (N_14546,N_13875,N_13442);
nand U14547 (N_14547,N_13781,N_13355);
or U14548 (N_14548,N_13585,N_13244);
xor U14549 (N_14549,N_13502,N_13125);
nand U14550 (N_14550,N_13577,N_13186);
xnor U14551 (N_14551,N_13955,N_13045);
and U14552 (N_14552,N_13417,N_13883);
and U14553 (N_14553,N_13210,N_13671);
xor U14554 (N_14554,N_13190,N_13179);
xnor U14555 (N_14555,N_13409,N_13784);
or U14556 (N_14556,N_13612,N_13191);
or U14557 (N_14557,N_13172,N_13542);
nand U14558 (N_14558,N_13654,N_13589);
xor U14559 (N_14559,N_13027,N_13394);
nor U14560 (N_14560,N_13936,N_13323);
or U14561 (N_14561,N_13798,N_13550);
nor U14562 (N_14562,N_13101,N_13184);
and U14563 (N_14563,N_13649,N_13534);
and U14564 (N_14564,N_13011,N_13019);
xor U14565 (N_14565,N_13395,N_13891);
nor U14566 (N_14566,N_13569,N_13614);
nor U14567 (N_14567,N_13802,N_13761);
or U14568 (N_14568,N_13313,N_13744);
xnor U14569 (N_14569,N_13568,N_13187);
nand U14570 (N_14570,N_13097,N_13411);
or U14571 (N_14571,N_13302,N_13376);
or U14572 (N_14572,N_13182,N_13908);
or U14573 (N_14573,N_13413,N_13801);
nand U14574 (N_14574,N_13191,N_13609);
nand U14575 (N_14575,N_13957,N_13964);
and U14576 (N_14576,N_13708,N_13157);
or U14577 (N_14577,N_13485,N_13170);
xnor U14578 (N_14578,N_13474,N_13964);
nor U14579 (N_14579,N_13416,N_13022);
nand U14580 (N_14580,N_13524,N_13333);
and U14581 (N_14581,N_13900,N_13966);
xnor U14582 (N_14582,N_13764,N_13059);
nor U14583 (N_14583,N_13279,N_13372);
nand U14584 (N_14584,N_13475,N_13500);
nand U14585 (N_14585,N_13938,N_13529);
nor U14586 (N_14586,N_13893,N_13021);
nor U14587 (N_14587,N_13627,N_13986);
xor U14588 (N_14588,N_13627,N_13237);
nand U14589 (N_14589,N_13964,N_13256);
xor U14590 (N_14590,N_13502,N_13386);
xnor U14591 (N_14591,N_13657,N_13016);
xnor U14592 (N_14592,N_13159,N_13480);
xnor U14593 (N_14593,N_13709,N_13820);
and U14594 (N_14594,N_13989,N_13219);
and U14595 (N_14595,N_13351,N_13609);
and U14596 (N_14596,N_13195,N_13009);
and U14597 (N_14597,N_13600,N_13501);
nand U14598 (N_14598,N_13254,N_13517);
or U14599 (N_14599,N_13855,N_13674);
and U14600 (N_14600,N_13405,N_13376);
xnor U14601 (N_14601,N_13025,N_13769);
xnor U14602 (N_14602,N_13568,N_13896);
xor U14603 (N_14603,N_13428,N_13427);
xnor U14604 (N_14604,N_13506,N_13375);
and U14605 (N_14605,N_13603,N_13036);
and U14606 (N_14606,N_13428,N_13102);
nand U14607 (N_14607,N_13882,N_13346);
or U14608 (N_14608,N_13104,N_13934);
or U14609 (N_14609,N_13230,N_13273);
nor U14610 (N_14610,N_13452,N_13483);
and U14611 (N_14611,N_13141,N_13571);
or U14612 (N_14612,N_13958,N_13783);
and U14613 (N_14613,N_13264,N_13520);
xnor U14614 (N_14614,N_13440,N_13815);
nand U14615 (N_14615,N_13187,N_13057);
nand U14616 (N_14616,N_13318,N_13841);
or U14617 (N_14617,N_13226,N_13190);
nor U14618 (N_14618,N_13200,N_13041);
and U14619 (N_14619,N_13670,N_13950);
or U14620 (N_14620,N_13864,N_13067);
and U14621 (N_14621,N_13972,N_13469);
and U14622 (N_14622,N_13366,N_13407);
or U14623 (N_14623,N_13880,N_13209);
and U14624 (N_14624,N_13553,N_13708);
nand U14625 (N_14625,N_13687,N_13969);
and U14626 (N_14626,N_13806,N_13414);
or U14627 (N_14627,N_13423,N_13326);
nor U14628 (N_14628,N_13928,N_13051);
xor U14629 (N_14629,N_13244,N_13973);
nor U14630 (N_14630,N_13104,N_13281);
nor U14631 (N_14631,N_13716,N_13793);
xor U14632 (N_14632,N_13560,N_13211);
nor U14633 (N_14633,N_13628,N_13928);
nor U14634 (N_14634,N_13403,N_13389);
nor U14635 (N_14635,N_13224,N_13523);
nand U14636 (N_14636,N_13948,N_13274);
nand U14637 (N_14637,N_13156,N_13587);
nor U14638 (N_14638,N_13922,N_13091);
xnor U14639 (N_14639,N_13215,N_13811);
xor U14640 (N_14640,N_13858,N_13705);
nor U14641 (N_14641,N_13735,N_13856);
nand U14642 (N_14642,N_13879,N_13685);
xor U14643 (N_14643,N_13954,N_13177);
nor U14644 (N_14644,N_13181,N_13001);
nand U14645 (N_14645,N_13588,N_13761);
or U14646 (N_14646,N_13436,N_13599);
or U14647 (N_14647,N_13792,N_13143);
nand U14648 (N_14648,N_13805,N_13802);
xnor U14649 (N_14649,N_13433,N_13761);
nor U14650 (N_14650,N_13584,N_13876);
or U14651 (N_14651,N_13355,N_13621);
xor U14652 (N_14652,N_13515,N_13110);
and U14653 (N_14653,N_13922,N_13441);
nand U14654 (N_14654,N_13414,N_13989);
xnor U14655 (N_14655,N_13884,N_13622);
nor U14656 (N_14656,N_13036,N_13013);
or U14657 (N_14657,N_13522,N_13789);
nor U14658 (N_14658,N_13497,N_13606);
nor U14659 (N_14659,N_13481,N_13462);
or U14660 (N_14660,N_13945,N_13787);
or U14661 (N_14661,N_13822,N_13074);
xnor U14662 (N_14662,N_13245,N_13502);
xor U14663 (N_14663,N_13340,N_13260);
xor U14664 (N_14664,N_13367,N_13221);
and U14665 (N_14665,N_13043,N_13341);
xor U14666 (N_14666,N_13433,N_13743);
xor U14667 (N_14667,N_13188,N_13266);
xnor U14668 (N_14668,N_13422,N_13451);
and U14669 (N_14669,N_13628,N_13033);
xor U14670 (N_14670,N_13221,N_13109);
xor U14671 (N_14671,N_13378,N_13608);
or U14672 (N_14672,N_13232,N_13777);
and U14673 (N_14673,N_13596,N_13362);
nor U14674 (N_14674,N_13278,N_13040);
nor U14675 (N_14675,N_13815,N_13385);
or U14676 (N_14676,N_13884,N_13985);
or U14677 (N_14677,N_13528,N_13747);
nand U14678 (N_14678,N_13041,N_13227);
or U14679 (N_14679,N_13695,N_13966);
nor U14680 (N_14680,N_13673,N_13263);
and U14681 (N_14681,N_13328,N_13146);
nor U14682 (N_14682,N_13542,N_13224);
xnor U14683 (N_14683,N_13081,N_13070);
nand U14684 (N_14684,N_13256,N_13026);
nor U14685 (N_14685,N_13904,N_13842);
nor U14686 (N_14686,N_13452,N_13438);
xor U14687 (N_14687,N_13531,N_13397);
nand U14688 (N_14688,N_13790,N_13301);
xor U14689 (N_14689,N_13583,N_13655);
or U14690 (N_14690,N_13808,N_13624);
and U14691 (N_14691,N_13748,N_13888);
xnor U14692 (N_14692,N_13175,N_13630);
or U14693 (N_14693,N_13292,N_13413);
or U14694 (N_14694,N_13042,N_13710);
nand U14695 (N_14695,N_13442,N_13613);
or U14696 (N_14696,N_13187,N_13807);
or U14697 (N_14697,N_13286,N_13351);
nand U14698 (N_14698,N_13780,N_13409);
and U14699 (N_14699,N_13501,N_13971);
nand U14700 (N_14700,N_13838,N_13854);
nand U14701 (N_14701,N_13418,N_13931);
nor U14702 (N_14702,N_13803,N_13395);
and U14703 (N_14703,N_13777,N_13898);
nor U14704 (N_14704,N_13219,N_13967);
nor U14705 (N_14705,N_13032,N_13953);
and U14706 (N_14706,N_13192,N_13545);
xor U14707 (N_14707,N_13590,N_13965);
or U14708 (N_14708,N_13814,N_13616);
or U14709 (N_14709,N_13190,N_13273);
nor U14710 (N_14710,N_13094,N_13428);
and U14711 (N_14711,N_13769,N_13380);
nand U14712 (N_14712,N_13040,N_13628);
or U14713 (N_14713,N_13008,N_13985);
or U14714 (N_14714,N_13273,N_13508);
nor U14715 (N_14715,N_13790,N_13330);
nor U14716 (N_14716,N_13129,N_13379);
nand U14717 (N_14717,N_13096,N_13223);
xnor U14718 (N_14718,N_13494,N_13067);
and U14719 (N_14719,N_13943,N_13265);
and U14720 (N_14720,N_13921,N_13609);
nand U14721 (N_14721,N_13365,N_13125);
xnor U14722 (N_14722,N_13250,N_13642);
xor U14723 (N_14723,N_13282,N_13280);
nand U14724 (N_14724,N_13120,N_13960);
nor U14725 (N_14725,N_13973,N_13591);
and U14726 (N_14726,N_13186,N_13474);
nor U14727 (N_14727,N_13751,N_13756);
nand U14728 (N_14728,N_13637,N_13346);
and U14729 (N_14729,N_13031,N_13902);
or U14730 (N_14730,N_13135,N_13579);
xor U14731 (N_14731,N_13247,N_13240);
and U14732 (N_14732,N_13513,N_13710);
nand U14733 (N_14733,N_13460,N_13287);
and U14734 (N_14734,N_13664,N_13794);
xor U14735 (N_14735,N_13647,N_13627);
nor U14736 (N_14736,N_13422,N_13828);
or U14737 (N_14737,N_13904,N_13224);
xnor U14738 (N_14738,N_13792,N_13650);
nand U14739 (N_14739,N_13657,N_13653);
nor U14740 (N_14740,N_13340,N_13885);
or U14741 (N_14741,N_13784,N_13371);
xor U14742 (N_14742,N_13819,N_13513);
nand U14743 (N_14743,N_13254,N_13799);
nor U14744 (N_14744,N_13733,N_13168);
nand U14745 (N_14745,N_13632,N_13988);
nand U14746 (N_14746,N_13405,N_13921);
or U14747 (N_14747,N_13573,N_13113);
and U14748 (N_14748,N_13457,N_13298);
and U14749 (N_14749,N_13698,N_13035);
xnor U14750 (N_14750,N_13061,N_13116);
nor U14751 (N_14751,N_13646,N_13732);
xor U14752 (N_14752,N_13330,N_13442);
nor U14753 (N_14753,N_13212,N_13568);
nor U14754 (N_14754,N_13398,N_13996);
xor U14755 (N_14755,N_13749,N_13477);
or U14756 (N_14756,N_13382,N_13647);
and U14757 (N_14757,N_13922,N_13901);
or U14758 (N_14758,N_13015,N_13984);
xnor U14759 (N_14759,N_13045,N_13118);
nor U14760 (N_14760,N_13314,N_13568);
xnor U14761 (N_14761,N_13872,N_13518);
and U14762 (N_14762,N_13658,N_13177);
or U14763 (N_14763,N_13498,N_13693);
nand U14764 (N_14764,N_13376,N_13721);
nor U14765 (N_14765,N_13533,N_13549);
and U14766 (N_14766,N_13309,N_13930);
or U14767 (N_14767,N_13074,N_13166);
or U14768 (N_14768,N_13986,N_13527);
xor U14769 (N_14769,N_13750,N_13387);
nor U14770 (N_14770,N_13954,N_13175);
nor U14771 (N_14771,N_13243,N_13179);
or U14772 (N_14772,N_13327,N_13716);
or U14773 (N_14773,N_13370,N_13628);
nor U14774 (N_14774,N_13746,N_13905);
xnor U14775 (N_14775,N_13754,N_13640);
nor U14776 (N_14776,N_13922,N_13382);
nand U14777 (N_14777,N_13900,N_13945);
nand U14778 (N_14778,N_13476,N_13770);
nand U14779 (N_14779,N_13813,N_13562);
xnor U14780 (N_14780,N_13042,N_13944);
nor U14781 (N_14781,N_13454,N_13355);
nor U14782 (N_14782,N_13178,N_13344);
nor U14783 (N_14783,N_13885,N_13272);
or U14784 (N_14784,N_13593,N_13853);
xor U14785 (N_14785,N_13157,N_13968);
or U14786 (N_14786,N_13064,N_13249);
and U14787 (N_14787,N_13010,N_13065);
and U14788 (N_14788,N_13156,N_13012);
or U14789 (N_14789,N_13426,N_13091);
nand U14790 (N_14790,N_13941,N_13772);
nand U14791 (N_14791,N_13179,N_13438);
nor U14792 (N_14792,N_13181,N_13857);
or U14793 (N_14793,N_13465,N_13900);
and U14794 (N_14794,N_13548,N_13578);
nand U14795 (N_14795,N_13868,N_13784);
nor U14796 (N_14796,N_13881,N_13235);
nand U14797 (N_14797,N_13788,N_13930);
and U14798 (N_14798,N_13602,N_13229);
and U14799 (N_14799,N_13629,N_13110);
xor U14800 (N_14800,N_13382,N_13591);
or U14801 (N_14801,N_13384,N_13372);
nor U14802 (N_14802,N_13772,N_13041);
and U14803 (N_14803,N_13811,N_13830);
nand U14804 (N_14804,N_13561,N_13621);
and U14805 (N_14805,N_13607,N_13331);
xnor U14806 (N_14806,N_13324,N_13880);
or U14807 (N_14807,N_13360,N_13487);
or U14808 (N_14808,N_13361,N_13722);
and U14809 (N_14809,N_13942,N_13768);
xor U14810 (N_14810,N_13441,N_13572);
xor U14811 (N_14811,N_13738,N_13762);
or U14812 (N_14812,N_13054,N_13733);
and U14813 (N_14813,N_13513,N_13497);
and U14814 (N_14814,N_13362,N_13599);
nand U14815 (N_14815,N_13324,N_13350);
or U14816 (N_14816,N_13944,N_13723);
and U14817 (N_14817,N_13791,N_13999);
and U14818 (N_14818,N_13458,N_13598);
nand U14819 (N_14819,N_13658,N_13689);
and U14820 (N_14820,N_13169,N_13459);
nand U14821 (N_14821,N_13529,N_13881);
or U14822 (N_14822,N_13871,N_13974);
nor U14823 (N_14823,N_13560,N_13126);
or U14824 (N_14824,N_13917,N_13766);
nor U14825 (N_14825,N_13039,N_13667);
xor U14826 (N_14826,N_13195,N_13244);
nand U14827 (N_14827,N_13507,N_13513);
nor U14828 (N_14828,N_13536,N_13273);
and U14829 (N_14829,N_13258,N_13972);
nand U14830 (N_14830,N_13463,N_13139);
xnor U14831 (N_14831,N_13624,N_13651);
nand U14832 (N_14832,N_13481,N_13400);
or U14833 (N_14833,N_13529,N_13277);
nor U14834 (N_14834,N_13669,N_13072);
nor U14835 (N_14835,N_13549,N_13433);
xnor U14836 (N_14836,N_13079,N_13161);
nand U14837 (N_14837,N_13319,N_13028);
nor U14838 (N_14838,N_13345,N_13690);
and U14839 (N_14839,N_13903,N_13942);
and U14840 (N_14840,N_13444,N_13456);
nand U14841 (N_14841,N_13071,N_13651);
nor U14842 (N_14842,N_13476,N_13376);
and U14843 (N_14843,N_13315,N_13252);
and U14844 (N_14844,N_13006,N_13081);
or U14845 (N_14845,N_13733,N_13429);
and U14846 (N_14846,N_13046,N_13437);
nand U14847 (N_14847,N_13761,N_13022);
xnor U14848 (N_14848,N_13799,N_13186);
and U14849 (N_14849,N_13678,N_13253);
and U14850 (N_14850,N_13659,N_13601);
and U14851 (N_14851,N_13460,N_13522);
xnor U14852 (N_14852,N_13215,N_13543);
and U14853 (N_14853,N_13842,N_13767);
or U14854 (N_14854,N_13632,N_13184);
and U14855 (N_14855,N_13624,N_13372);
nand U14856 (N_14856,N_13479,N_13304);
and U14857 (N_14857,N_13419,N_13001);
nor U14858 (N_14858,N_13796,N_13576);
nand U14859 (N_14859,N_13203,N_13848);
xnor U14860 (N_14860,N_13462,N_13930);
nor U14861 (N_14861,N_13051,N_13799);
or U14862 (N_14862,N_13569,N_13829);
or U14863 (N_14863,N_13124,N_13940);
nor U14864 (N_14864,N_13612,N_13801);
xor U14865 (N_14865,N_13565,N_13696);
or U14866 (N_14866,N_13907,N_13595);
nor U14867 (N_14867,N_13335,N_13233);
nor U14868 (N_14868,N_13490,N_13692);
and U14869 (N_14869,N_13691,N_13523);
or U14870 (N_14870,N_13646,N_13538);
and U14871 (N_14871,N_13569,N_13361);
or U14872 (N_14872,N_13876,N_13382);
nor U14873 (N_14873,N_13206,N_13937);
or U14874 (N_14874,N_13631,N_13061);
nor U14875 (N_14875,N_13735,N_13118);
nor U14876 (N_14876,N_13488,N_13154);
nor U14877 (N_14877,N_13534,N_13291);
xor U14878 (N_14878,N_13623,N_13201);
or U14879 (N_14879,N_13444,N_13678);
xnor U14880 (N_14880,N_13870,N_13899);
and U14881 (N_14881,N_13764,N_13489);
xnor U14882 (N_14882,N_13463,N_13415);
nor U14883 (N_14883,N_13329,N_13786);
and U14884 (N_14884,N_13496,N_13949);
nand U14885 (N_14885,N_13059,N_13452);
xor U14886 (N_14886,N_13923,N_13020);
xor U14887 (N_14887,N_13751,N_13053);
and U14888 (N_14888,N_13892,N_13169);
or U14889 (N_14889,N_13413,N_13782);
xor U14890 (N_14890,N_13780,N_13481);
nor U14891 (N_14891,N_13781,N_13120);
and U14892 (N_14892,N_13119,N_13297);
nor U14893 (N_14893,N_13000,N_13822);
or U14894 (N_14894,N_13810,N_13797);
nand U14895 (N_14895,N_13494,N_13846);
nand U14896 (N_14896,N_13434,N_13886);
nand U14897 (N_14897,N_13266,N_13199);
nor U14898 (N_14898,N_13643,N_13813);
xnor U14899 (N_14899,N_13558,N_13601);
nand U14900 (N_14900,N_13588,N_13954);
xnor U14901 (N_14901,N_13234,N_13470);
nor U14902 (N_14902,N_13690,N_13314);
and U14903 (N_14903,N_13607,N_13565);
nor U14904 (N_14904,N_13849,N_13365);
nand U14905 (N_14905,N_13744,N_13232);
nand U14906 (N_14906,N_13279,N_13461);
xor U14907 (N_14907,N_13814,N_13107);
and U14908 (N_14908,N_13462,N_13103);
or U14909 (N_14909,N_13795,N_13715);
nand U14910 (N_14910,N_13152,N_13652);
nand U14911 (N_14911,N_13313,N_13435);
nor U14912 (N_14912,N_13516,N_13308);
nor U14913 (N_14913,N_13614,N_13489);
or U14914 (N_14914,N_13472,N_13227);
or U14915 (N_14915,N_13844,N_13123);
or U14916 (N_14916,N_13443,N_13884);
nand U14917 (N_14917,N_13182,N_13108);
nor U14918 (N_14918,N_13858,N_13996);
or U14919 (N_14919,N_13365,N_13613);
and U14920 (N_14920,N_13103,N_13130);
nand U14921 (N_14921,N_13103,N_13229);
or U14922 (N_14922,N_13412,N_13233);
and U14923 (N_14923,N_13360,N_13807);
and U14924 (N_14924,N_13614,N_13450);
or U14925 (N_14925,N_13664,N_13153);
nand U14926 (N_14926,N_13449,N_13734);
or U14927 (N_14927,N_13404,N_13268);
nand U14928 (N_14928,N_13239,N_13703);
or U14929 (N_14929,N_13041,N_13837);
and U14930 (N_14930,N_13092,N_13095);
xnor U14931 (N_14931,N_13297,N_13947);
nand U14932 (N_14932,N_13892,N_13419);
xor U14933 (N_14933,N_13130,N_13152);
nand U14934 (N_14934,N_13619,N_13458);
xor U14935 (N_14935,N_13206,N_13774);
or U14936 (N_14936,N_13600,N_13085);
nand U14937 (N_14937,N_13759,N_13441);
nand U14938 (N_14938,N_13840,N_13913);
nor U14939 (N_14939,N_13040,N_13726);
nor U14940 (N_14940,N_13746,N_13459);
and U14941 (N_14941,N_13495,N_13988);
and U14942 (N_14942,N_13058,N_13347);
nand U14943 (N_14943,N_13853,N_13094);
nor U14944 (N_14944,N_13863,N_13423);
xor U14945 (N_14945,N_13708,N_13656);
and U14946 (N_14946,N_13802,N_13243);
nor U14947 (N_14947,N_13559,N_13460);
and U14948 (N_14948,N_13217,N_13701);
or U14949 (N_14949,N_13757,N_13103);
or U14950 (N_14950,N_13599,N_13193);
and U14951 (N_14951,N_13243,N_13091);
nand U14952 (N_14952,N_13406,N_13385);
and U14953 (N_14953,N_13663,N_13302);
nand U14954 (N_14954,N_13718,N_13617);
or U14955 (N_14955,N_13189,N_13431);
xor U14956 (N_14956,N_13986,N_13688);
and U14957 (N_14957,N_13299,N_13767);
and U14958 (N_14958,N_13359,N_13116);
xnor U14959 (N_14959,N_13283,N_13414);
or U14960 (N_14960,N_13477,N_13603);
xor U14961 (N_14961,N_13947,N_13920);
nand U14962 (N_14962,N_13900,N_13432);
or U14963 (N_14963,N_13865,N_13231);
or U14964 (N_14964,N_13843,N_13361);
nand U14965 (N_14965,N_13981,N_13584);
nor U14966 (N_14966,N_13269,N_13921);
and U14967 (N_14967,N_13202,N_13288);
and U14968 (N_14968,N_13330,N_13019);
xnor U14969 (N_14969,N_13339,N_13830);
nand U14970 (N_14970,N_13719,N_13642);
xor U14971 (N_14971,N_13912,N_13174);
nand U14972 (N_14972,N_13100,N_13880);
xor U14973 (N_14973,N_13020,N_13171);
nor U14974 (N_14974,N_13007,N_13351);
nor U14975 (N_14975,N_13396,N_13663);
xnor U14976 (N_14976,N_13981,N_13839);
or U14977 (N_14977,N_13775,N_13818);
nor U14978 (N_14978,N_13989,N_13842);
nand U14979 (N_14979,N_13541,N_13316);
nand U14980 (N_14980,N_13315,N_13203);
xnor U14981 (N_14981,N_13877,N_13365);
nor U14982 (N_14982,N_13602,N_13630);
nand U14983 (N_14983,N_13128,N_13116);
and U14984 (N_14984,N_13391,N_13881);
xor U14985 (N_14985,N_13079,N_13694);
xnor U14986 (N_14986,N_13668,N_13563);
or U14987 (N_14987,N_13964,N_13456);
or U14988 (N_14988,N_13337,N_13389);
nor U14989 (N_14989,N_13478,N_13667);
xor U14990 (N_14990,N_13136,N_13745);
and U14991 (N_14991,N_13826,N_13085);
nor U14992 (N_14992,N_13105,N_13776);
and U14993 (N_14993,N_13988,N_13331);
nor U14994 (N_14994,N_13381,N_13210);
or U14995 (N_14995,N_13782,N_13346);
or U14996 (N_14996,N_13717,N_13012);
nor U14997 (N_14997,N_13516,N_13833);
or U14998 (N_14998,N_13800,N_13937);
xnor U14999 (N_14999,N_13333,N_13556);
or U15000 (N_15000,N_14969,N_14940);
xor U15001 (N_15001,N_14056,N_14182);
or U15002 (N_15002,N_14154,N_14738);
nor U15003 (N_15003,N_14540,N_14436);
xor U15004 (N_15004,N_14227,N_14753);
nor U15005 (N_15005,N_14390,N_14083);
xor U15006 (N_15006,N_14462,N_14243);
xor U15007 (N_15007,N_14952,N_14121);
nand U15008 (N_15008,N_14471,N_14675);
xor U15009 (N_15009,N_14316,N_14449);
or U15010 (N_15010,N_14160,N_14334);
xnor U15011 (N_15011,N_14102,N_14809);
nor U15012 (N_15012,N_14852,N_14130);
and U15013 (N_15013,N_14114,N_14556);
and U15014 (N_15014,N_14444,N_14304);
nor U15015 (N_15015,N_14187,N_14501);
and U15016 (N_15016,N_14564,N_14917);
xor U15017 (N_15017,N_14957,N_14399);
nand U15018 (N_15018,N_14290,N_14080);
or U15019 (N_15019,N_14499,N_14126);
nand U15020 (N_15020,N_14301,N_14885);
nand U15021 (N_15021,N_14202,N_14495);
nand U15022 (N_15022,N_14104,N_14192);
nor U15023 (N_15023,N_14335,N_14826);
and U15024 (N_15024,N_14589,N_14156);
nor U15025 (N_15025,N_14461,N_14504);
and U15026 (N_15026,N_14568,N_14300);
nand U15027 (N_15027,N_14094,N_14140);
nor U15028 (N_15028,N_14904,N_14880);
nor U15029 (N_15029,N_14167,N_14332);
nand U15030 (N_15030,N_14420,N_14312);
nor U15031 (N_15031,N_14092,N_14820);
xor U15032 (N_15032,N_14124,N_14109);
nor U15033 (N_15033,N_14922,N_14855);
or U15034 (N_15034,N_14977,N_14728);
and U15035 (N_15035,N_14769,N_14649);
nor U15036 (N_15036,N_14624,N_14910);
xnor U15037 (N_15037,N_14660,N_14017);
nor U15038 (N_15038,N_14741,N_14849);
xnor U15039 (N_15039,N_14196,N_14981);
xor U15040 (N_15040,N_14199,N_14630);
nand U15041 (N_15041,N_14889,N_14451);
xnor U15042 (N_15042,N_14309,N_14257);
nand U15043 (N_15043,N_14232,N_14413);
nor U15044 (N_15044,N_14747,N_14744);
and U15045 (N_15045,N_14680,N_14275);
and U15046 (N_15046,N_14547,N_14064);
xor U15047 (N_15047,N_14185,N_14356);
or U15048 (N_15048,N_14678,N_14530);
nor U15049 (N_15049,N_14091,N_14598);
nor U15050 (N_15050,N_14293,N_14037);
and U15051 (N_15051,N_14523,N_14086);
or U15052 (N_15052,N_14022,N_14221);
xnor U15053 (N_15053,N_14596,N_14672);
or U15054 (N_15054,N_14584,N_14563);
and U15055 (N_15055,N_14827,N_14722);
or U15056 (N_15056,N_14638,N_14016);
nand U15057 (N_15057,N_14143,N_14176);
or U15058 (N_15058,N_14215,N_14318);
and U15059 (N_15059,N_14695,N_14245);
xnor U15060 (N_15060,N_14162,N_14305);
or U15061 (N_15061,N_14492,N_14720);
nor U15062 (N_15062,N_14347,N_14433);
xor U15063 (N_15063,N_14098,N_14805);
and U15064 (N_15064,N_14198,N_14005);
xnor U15065 (N_15065,N_14682,N_14049);
or U15066 (N_15066,N_14396,N_14980);
nand U15067 (N_15067,N_14363,N_14976);
nor U15068 (N_15068,N_14455,N_14766);
or U15069 (N_15069,N_14476,N_14752);
nor U15070 (N_15070,N_14352,N_14844);
nor U15071 (N_15071,N_14522,N_14090);
nand U15072 (N_15072,N_14319,N_14018);
nand U15073 (N_15073,N_14466,N_14155);
xor U15074 (N_15074,N_14015,N_14958);
xor U15075 (N_15075,N_14440,N_14963);
or U15076 (N_15076,N_14600,N_14919);
or U15077 (N_15077,N_14531,N_14566);
nand U15078 (N_15078,N_14573,N_14705);
xor U15079 (N_15079,N_14250,N_14613);
nor U15080 (N_15080,N_14979,N_14278);
nand U15081 (N_15081,N_14608,N_14190);
and U15082 (N_15082,N_14913,N_14314);
or U15083 (N_15083,N_14838,N_14380);
nand U15084 (N_15084,N_14972,N_14004);
or U15085 (N_15085,N_14467,N_14191);
and U15086 (N_15086,N_14555,N_14830);
nor U15087 (N_15087,N_14279,N_14967);
nor U15088 (N_15088,N_14469,N_14841);
and U15089 (N_15089,N_14120,N_14439);
xor U15090 (N_15090,N_14585,N_14175);
nand U15091 (N_15091,N_14475,N_14622);
and U15092 (N_15092,N_14169,N_14510);
or U15093 (N_15093,N_14951,N_14829);
xnor U15094 (N_15094,N_14842,N_14450);
or U15095 (N_15095,N_14822,N_14403);
nor U15096 (N_15096,N_14365,N_14428);
nor U15097 (N_15097,N_14020,N_14574);
nor U15098 (N_15098,N_14170,N_14821);
nor U15099 (N_15099,N_14000,N_14061);
and U15100 (N_15100,N_14087,N_14375);
and U15101 (N_15101,N_14535,N_14276);
or U15102 (N_15102,N_14549,N_14161);
xnor U15103 (N_15103,N_14871,N_14545);
xnor U15104 (N_15104,N_14548,N_14872);
xnor U15105 (N_15105,N_14478,N_14618);
and U15106 (N_15106,N_14453,N_14108);
xnor U15107 (N_15107,N_14737,N_14485);
and U15108 (N_15108,N_14780,N_14788);
or U15109 (N_15109,N_14659,N_14890);
nor U15110 (N_15110,N_14359,N_14012);
xor U15111 (N_15111,N_14427,N_14664);
nor U15112 (N_15112,N_14599,N_14645);
xnor U15113 (N_15113,N_14321,N_14813);
and U15114 (N_15114,N_14745,N_14074);
nand U15115 (N_15115,N_14797,N_14222);
or U15116 (N_15116,N_14315,N_14764);
or U15117 (N_15117,N_14149,N_14799);
or U15118 (N_15118,N_14477,N_14908);
nor U15119 (N_15119,N_14690,N_14106);
xor U15120 (N_15120,N_14357,N_14336);
or U15121 (N_15121,N_14644,N_14537);
xnor U15122 (N_15122,N_14372,N_14570);
nor U15123 (N_15123,N_14238,N_14718);
and U15124 (N_15124,N_14544,N_14325);
xnor U15125 (N_15125,N_14247,N_14947);
and U15126 (N_15126,N_14837,N_14039);
or U15127 (N_15127,N_14425,N_14786);
and U15128 (N_15128,N_14628,N_14629);
nand U15129 (N_15129,N_14873,N_14714);
xor U15130 (N_15130,N_14231,N_14704);
nor U15131 (N_15131,N_14463,N_14429);
nand U15132 (N_15132,N_14076,N_14740);
xnor U15133 (N_15133,N_14691,N_14137);
xor U15134 (N_15134,N_14804,N_14223);
nand U15135 (N_15135,N_14962,N_14857);
and U15136 (N_15136,N_14875,N_14408);
or U15137 (N_15137,N_14409,N_14938);
xnor U15138 (N_15138,N_14671,N_14729);
nand U15139 (N_15139,N_14369,N_14755);
xor U15140 (N_15140,N_14031,N_14028);
or U15141 (N_15141,N_14320,N_14441);
or U15142 (N_15142,N_14684,N_14867);
xnor U15143 (N_15143,N_14734,N_14946);
nor U15144 (N_15144,N_14557,N_14953);
xnor U15145 (N_15145,N_14751,N_14870);
nor U15146 (N_15146,N_14254,N_14990);
nor U15147 (N_15147,N_14996,N_14330);
nor U15148 (N_15148,N_14151,N_14225);
nand U15149 (N_15149,N_14736,N_14586);
and U15150 (N_15150,N_14267,N_14932);
or U15151 (N_15151,N_14302,N_14412);
nor U15152 (N_15152,N_14416,N_14378);
or U15153 (N_15153,N_14253,N_14771);
xor U15154 (N_15154,N_14667,N_14533);
and U15155 (N_15155,N_14240,N_14043);
and U15156 (N_15156,N_14139,N_14653);
nand U15157 (N_15157,N_14159,N_14526);
nor U15158 (N_15158,N_14132,N_14474);
nand U15159 (N_15159,N_14717,N_14411);
xnor U15160 (N_15160,N_14107,N_14343);
and U15161 (N_15161,N_14702,N_14306);
and U15162 (N_15162,N_14577,N_14341);
nand U15163 (N_15163,N_14134,N_14295);
and U15164 (N_15164,N_14327,N_14975);
nand U15165 (N_15165,N_14898,N_14479);
xnor U15166 (N_15166,N_14065,N_14933);
nor U15167 (N_15167,N_14970,N_14235);
xor U15168 (N_15168,N_14739,N_14559);
xor U15169 (N_15169,N_14950,N_14034);
or U15170 (N_15170,N_14846,N_14512);
nor U15171 (N_15171,N_14633,N_14955);
or U15172 (N_15172,N_14208,N_14835);
xnor U15173 (N_15173,N_14165,N_14541);
xor U15174 (N_15174,N_14597,N_14284);
and U15175 (N_15175,N_14850,N_14438);
nand U15176 (N_15176,N_14219,N_14572);
nor U15177 (N_15177,N_14640,N_14171);
or U15178 (N_15178,N_14986,N_14650);
xor U15179 (N_15179,N_14553,N_14355);
nand U15180 (N_15180,N_14988,N_14576);
nor U15181 (N_15181,N_14242,N_14693);
nand U15182 (N_15182,N_14795,N_14839);
nand U15183 (N_15183,N_14311,N_14026);
and U15184 (N_15184,N_14882,N_14903);
nand U15185 (N_15185,N_14349,N_14603);
or U15186 (N_15186,N_14317,N_14847);
or U15187 (N_15187,N_14041,N_14796);
and U15188 (N_15188,N_14733,N_14960);
or U15189 (N_15189,N_14538,N_14498);
or U15190 (N_15190,N_14296,N_14234);
nand U15191 (N_15191,N_14641,N_14899);
xnor U15192 (N_15192,N_14674,N_14552);
nor U15193 (N_15193,N_14760,N_14272);
or U15194 (N_15194,N_14496,N_14178);
nor U15195 (N_15195,N_14135,N_14900);
xor U15196 (N_15196,N_14874,N_14848);
or U15197 (N_15197,N_14731,N_14619);
nor U15198 (N_15198,N_14735,N_14112);
and U15199 (N_15199,N_14713,N_14019);
or U15200 (N_15200,N_14285,N_14689);
nand U15201 (N_15201,N_14511,N_14730);
and U15202 (N_15202,N_14150,N_14864);
or U15203 (N_15203,N_14994,N_14186);
xnor U15204 (N_15204,N_14604,N_14807);
nor U15205 (N_15205,N_14033,N_14582);
and U15206 (N_15206,N_14237,N_14129);
xnor U15207 (N_15207,N_14626,N_14878);
and U15208 (N_15208,N_14832,N_14609);
or U15209 (N_15209,N_14534,N_14010);
nand U15210 (N_15210,N_14153,N_14793);
or U15211 (N_15211,N_14881,N_14710);
xnor U15212 (N_15212,N_14201,N_14400);
xor U15213 (N_15213,N_14648,N_14580);
xnor U15214 (N_15214,N_14269,N_14063);
xor U15215 (N_15215,N_14434,N_14959);
xor U15216 (N_15216,N_14442,N_14457);
or U15217 (N_15217,N_14014,N_14754);
and U15218 (N_15218,N_14184,N_14520);
nand U15219 (N_15219,N_14048,N_14152);
nand U15220 (N_15220,N_14519,N_14070);
nor U15221 (N_15221,N_14507,N_14289);
xnor U15222 (N_15222,N_14658,N_14044);
nand U15223 (N_15223,N_14765,N_14971);
or U15224 (N_15224,N_14924,N_14926);
nand U15225 (N_15225,N_14998,N_14265);
xor U15226 (N_15226,N_14213,N_14949);
xor U15227 (N_15227,N_14773,N_14274);
nor U15228 (N_15228,N_14709,N_14188);
or U15229 (N_15229,N_14775,N_14113);
or U15230 (N_15230,N_14100,N_14164);
or U15231 (N_15231,N_14383,N_14078);
nor U15232 (N_15232,N_14757,N_14790);
nor U15233 (N_15233,N_14825,N_14006);
nor U15234 (N_15234,N_14637,N_14244);
or U15235 (N_15235,N_14703,N_14402);
xnor U15236 (N_15236,N_14550,N_14360);
nor U15237 (N_15237,N_14561,N_14183);
nand U15238 (N_15238,N_14258,N_14344);
nand U15239 (N_15239,N_14816,N_14942);
nand U15240 (N_15240,N_14895,N_14869);
and U15241 (N_15241,N_14252,N_14647);
xnor U15242 (N_15242,N_14656,N_14923);
nand U15243 (N_15243,N_14029,N_14927);
nor U15244 (N_15244,N_14590,N_14491);
and U15245 (N_15245,N_14575,N_14662);
nor U15246 (N_15246,N_14866,N_14761);
xor U15247 (N_15247,N_14264,N_14639);
nor U15248 (N_15248,N_14886,N_14569);
xnor U15249 (N_15249,N_14912,N_14824);
xnor U15250 (N_15250,N_14785,N_14914);
or U15251 (N_15251,N_14116,N_14391);
or U15252 (N_15252,N_14494,N_14532);
nor U15253 (N_15253,N_14283,N_14207);
and U15254 (N_15254,N_14003,N_14101);
nor U15255 (N_15255,N_14750,N_14459);
and U15256 (N_15256,N_14422,N_14725);
nand U15257 (N_15257,N_14040,N_14055);
nand U15258 (N_15258,N_14211,N_14419);
xnor U15259 (N_15259,N_14509,N_14398);
and U15260 (N_15260,N_14758,N_14127);
nor U15261 (N_15261,N_14085,N_14936);
xor U15262 (N_15262,N_14468,N_14670);
nand U15263 (N_15263,N_14205,N_14935);
nor U15264 (N_15264,N_14606,N_14350);
nor U15265 (N_15265,N_14683,N_14431);
or U15266 (N_15266,N_14249,N_14214);
and U15267 (N_15267,N_14011,N_14669);
nor U15268 (N_15268,N_14934,N_14929);
and U15269 (N_15269,N_14464,N_14435);
and U15270 (N_15270,N_14546,N_14068);
nand U15271 (N_15271,N_14925,N_14261);
xnor U15272 (N_15272,N_14620,N_14862);
xnor U15273 (N_15273,N_14298,N_14907);
and U15274 (N_15274,N_14819,N_14587);
or U15275 (N_15275,N_14665,N_14726);
xnor U15276 (N_15276,N_14027,N_14749);
xnor U15277 (N_15277,N_14239,N_14337);
xnor U15278 (N_15278,N_14497,N_14397);
or U15279 (N_15279,N_14602,N_14681);
nor U15280 (N_15280,N_14798,N_14883);
xor U15281 (N_15281,N_14008,N_14338);
or U15282 (N_15282,N_14340,N_14921);
xnor U15283 (N_15283,N_14224,N_14173);
or U15284 (N_15284,N_14172,N_14262);
xnor U15285 (N_15285,N_14163,N_14291);
and U15286 (N_15286,N_14840,N_14313);
or U15287 (N_15287,N_14447,N_14787);
or U15288 (N_15288,N_14893,N_14905);
or U15289 (N_15289,N_14964,N_14777);
or U15290 (N_15290,N_14617,N_14456);
nand U15291 (N_15291,N_14808,N_14488);
xor U15292 (N_15292,N_14259,N_14646);
and U15293 (N_15293,N_14845,N_14333);
xor U15294 (N_15294,N_14013,N_14077);
xor U15295 (N_15295,N_14482,N_14723);
nand U15296 (N_15296,N_14452,N_14634);
nand U15297 (N_15297,N_14918,N_14487);
xnor U15298 (N_15298,N_14915,N_14268);
nand U15299 (N_15299,N_14260,N_14310);
nor U15300 (N_15300,N_14525,N_14217);
xnor U15301 (N_15301,N_14489,N_14030);
or U15302 (N_15302,N_14248,N_14288);
and U15303 (N_15303,N_14368,N_14147);
nand U15304 (N_15304,N_14303,N_14668);
xor U15305 (N_15305,N_14700,N_14414);
and U15306 (N_15306,N_14483,N_14328);
or U15307 (N_15307,N_14782,N_14685);
nor U15308 (N_15308,N_14698,N_14742);
xor U15309 (N_15309,N_14607,N_14326);
or U15310 (N_15310,N_14983,N_14542);
or U15311 (N_15311,N_14677,N_14993);
xnor U15312 (N_15312,N_14073,N_14810);
xor U15313 (N_15313,N_14323,N_14601);
nor U15314 (N_15314,N_14432,N_14251);
nand U15315 (N_15315,N_14888,N_14508);
nor U15316 (N_15316,N_14776,N_14699);
and U15317 (N_15317,N_14118,N_14529);
and U15318 (N_15318,N_14802,N_14756);
and U15319 (N_15319,N_14273,N_14715);
or U15320 (N_15320,N_14811,N_14407);
and U15321 (N_15321,N_14666,N_14067);
or U15322 (N_15322,N_14241,N_14516);
nand U15323 (N_15323,N_14036,N_14374);
nor U15324 (N_15324,N_14896,N_14768);
or U15325 (N_15325,N_14299,N_14930);
and U15326 (N_15326,N_14446,N_14505);
nand U15327 (N_15327,N_14592,N_14954);
and U15328 (N_15328,N_14351,N_14676);
nand U15329 (N_15329,N_14616,N_14581);
xor U15330 (N_15330,N_14051,N_14696);
xor U15331 (N_15331,N_14707,N_14853);
nand U15332 (N_15332,N_14901,N_14465);
nor U15333 (N_15333,N_14528,N_14806);
or U15334 (N_15334,N_14075,N_14943);
nor U15335 (N_15335,N_14122,N_14518);
xor U15336 (N_15336,N_14458,N_14995);
nand U15337 (N_15337,N_14454,N_14884);
or U15338 (N_15338,N_14643,N_14057);
xnor U15339 (N_15339,N_14803,N_14748);
or U15340 (N_15340,N_14687,N_14712);
xor U15341 (N_15341,N_14387,N_14554);
nand U15342 (N_15342,N_14181,N_14473);
and U15343 (N_15343,N_14145,N_14021);
nor U15344 (N_15344,N_14189,N_14042);
nor U15345 (N_15345,N_14636,N_14931);
nand U15346 (N_15346,N_14833,N_14423);
nor U15347 (N_15347,N_14887,N_14117);
and U15348 (N_15348,N_14082,N_14079);
or U15349 (N_15349,N_14370,N_14767);
or U15350 (N_15350,N_14783,N_14331);
and U15351 (N_15351,N_14916,N_14103);
nor U15352 (N_15352,N_14610,N_14035);
nor U15353 (N_15353,N_14791,N_14131);
or U15354 (N_15354,N_14395,N_14421);
nor U15355 (N_15355,N_14719,N_14345);
xor U15356 (N_15356,N_14158,N_14578);
xor U15357 (N_15357,N_14920,N_14448);
and U15358 (N_15358,N_14831,N_14472);
xor U15359 (N_15359,N_14136,N_14324);
or U15360 (N_15360,N_14418,N_14818);
nand U15361 (N_15361,N_14047,N_14661);
xnor U15362 (N_15362,N_14346,N_14937);
nand U15363 (N_15363,N_14814,N_14524);
or U15364 (N_15364,N_14892,N_14594);
nor U15365 (N_15365,N_14513,N_14210);
nand U15366 (N_15366,N_14774,N_14406);
nand U15367 (N_15367,N_14386,N_14342);
nor U15368 (N_15368,N_14792,N_14263);
nand U15369 (N_15369,N_14385,N_14093);
nor U15370 (N_15370,N_14377,N_14789);
and U15371 (N_15371,N_14911,N_14125);
nand U15372 (N_15372,N_14111,N_14974);
and U15373 (N_15373,N_14843,N_14817);
or U15374 (N_15374,N_14194,N_14379);
xnor U15375 (N_15375,N_14503,N_14373);
nand U15376 (N_15376,N_14579,N_14195);
nand U15377 (N_15377,N_14174,N_14621);
or U15378 (N_15378,N_14329,N_14404);
nand U15379 (N_15379,N_14024,N_14536);
nor U15380 (N_15380,N_14743,N_14066);
nor U15381 (N_15381,N_14657,N_14612);
or U15382 (N_15382,N_14627,N_14623);
nor U15383 (N_15383,N_14812,N_14128);
xnor U15384 (N_15384,N_14277,N_14220);
or U15385 (N_15385,N_14025,N_14692);
nor U15386 (N_15386,N_14706,N_14212);
and U15387 (N_15387,N_14828,N_14384);
nand U15388 (N_15388,N_14281,N_14746);
nor U15389 (N_15389,N_14292,N_14591);
nand U15390 (N_15390,N_14944,N_14089);
nor U15391 (N_15391,N_14157,N_14226);
or U15392 (N_15392,N_14961,N_14965);
nor U15393 (N_15393,N_14146,N_14486);
nor U15394 (N_15394,N_14851,N_14652);
nor U15395 (N_15395,N_14141,N_14339);
or U15396 (N_15396,N_14023,N_14354);
xnor U15397 (N_15397,N_14879,N_14415);
and U15398 (N_15398,N_14180,N_14115);
and U15399 (N_15399,N_14985,N_14361);
nand U15400 (N_15400,N_14992,N_14308);
nor U15401 (N_15401,N_14297,N_14228);
nand U15402 (N_15402,N_14437,N_14565);
and U15403 (N_15403,N_14539,N_14991);
nor U15404 (N_15404,N_14119,N_14987);
nand U15405 (N_15405,N_14956,N_14426);
and U15406 (N_15406,N_14778,N_14928);
and U15407 (N_15407,N_14209,N_14856);
nand U15408 (N_15408,N_14697,N_14865);
nand U15409 (N_15409,N_14654,N_14502);
xnor U15410 (N_15410,N_14514,N_14168);
nor U15411 (N_15411,N_14999,N_14280);
nand U15412 (N_15412,N_14894,N_14759);
and U15413 (N_15413,N_14688,N_14836);
or U15414 (N_15414,N_14562,N_14727);
and U15415 (N_15415,N_14142,N_14781);
nand U15416 (N_15416,N_14716,N_14506);
nand U15417 (N_15417,N_14001,N_14770);
nor U15418 (N_15418,N_14410,N_14353);
or U15419 (N_15419,N_14984,N_14470);
nand U15420 (N_15420,N_14294,N_14138);
xor U15421 (N_15421,N_14480,N_14651);
nand U15422 (N_15422,N_14054,N_14854);
nand U15423 (N_15423,N_14891,N_14784);
and U15424 (N_15424,N_14701,N_14038);
or U15425 (N_15425,N_14800,N_14200);
xnor U15426 (N_15426,N_14405,N_14877);
nand U15427 (N_15427,N_14417,N_14233);
nor U15428 (N_15428,N_14997,N_14179);
nand U15429 (N_15429,N_14246,N_14203);
nor U15430 (N_15430,N_14358,N_14148);
or U15431 (N_15431,N_14625,N_14968);
nand U15432 (N_15432,N_14307,N_14801);
nand U15433 (N_15433,N_14144,N_14364);
nor U15434 (N_15434,N_14567,N_14095);
nor U15435 (N_15435,N_14255,N_14543);
and U15436 (N_15436,N_14197,N_14271);
or U15437 (N_15437,N_14945,N_14517);
xnor U15438 (N_15438,N_14493,N_14206);
nor U15439 (N_15439,N_14071,N_14002);
xnor U15440 (N_15440,N_14939,N_14794);
and U15441 (N_15441,N_14348,N_14218);
nand U15442 (N_15442,N_14096,N_14445);
nand U15443 (N_15443,N_14069,N_14388);
nand U15444 (N_15444,N_14443,N_14941);
nor U15445 (N_15445,N_14763,N_14859);
xor U15446 (N_15446,N_14823,N_14389);
nor U15447 (N_15447,N_14088,N_14270);
xor U15448 (N_15448,N_14815,N_14460);
or U15449 (N_15449,N_14635,N_14858);
or U15450 (N_15450,N_14424,N_14050);
or U15451 (N_15451,N_14694,N_14834);
or U15452 (N_15452,N_14362,N_14382);
nor U15453 (N_15453,N_14322,N_14133);
or U15454 (N_15454,N_14058,N_14060);
xnor U15455 (N_15455,N_14721,N_14072);
nand U15456 (N_15456,N_14583,N_14724);
or U15457 (N_15457,N_14366,N_14266);
or U15458 (N_15458,N_14062,N_14177);
or U15459 (N_15459,N_14216,N_14863);
and U15460 (N_15460,N_14571,N_14558);
or U15461 (N_15461,N_14876,N_14595);
or U15462 (N_15462,N_14732,N_14632);
nor U15463 (N_15463,N_14394,N_14097);
or U15464 (N_15464,N_14105,N_14376);
nor U15465 (N_15465,N_14906,N_14673);
nand U15466 (N_15466,N_14401,N_14500);
nor U15467 (N_15467,N_14642,N_14663);
nand U15468 (N_15468,N_14204,N_14099);
xor U15469 (N_15469,N_14282,N_14430);
xor U15470 (N_15470,N_14711,N_14032);
and U15471 (N_15471,N_14236,N_14588);
or U15472 (N_15472,N_14081,N_14481);
nor U15473 (N_15473,N_14686,N_14084);
nand U15474 (N_15474,N_14593,N_14861);
nand U15475 (N_15475,N_14614,N_14521);
nor U15476 (N_15476,N_14897,N_14779);
xor U15477 (N_15477,N_14392,N_14978);
and U15478 (N_15478,N_14551,N_14909);
xor U15479 (N_15479,N_14560,N_14527);
xnor U15480 (N_15480,N_14966,N_14045);
or U15481 (N_15481,N_14868,N_14229);
xor U15482 (N_15482,N_14393,N_14052);
nand U15483 (N_15483,N_14287,N_14902);
and U15484 (N_15484,N_14059,N_14772);
xnor U15485 (N_15485,N_14989,N_14708);
xnor U15486 (N_15486,N_14973,N_14053);
and U15487 (N_15487,N_14948,N_14166);
nand U15488 (N_15488,N_14007,N_14367);
nand U15489 (N_15489,N_14230,N_14123);
nand U15490 (N_15490,N_14982,N_14631);
nor U15491 (N_15491,N_14371,N_14611);
or U15492 (N_15492,N_14286,N_14615);
xnor U15493 (N_15493,N_14490,N_14110);
or U15494 (N_15494,N_14605,N_14046);
nor U15495 (N_15495,N_14484,N_14515);
nand U15496 (N_15496,N_14655,N_14679);
nand U15497 (N_15497,N_14762,N_14860);
nor U15498 (N_15498,N_14009,N_14193);
xnor U15499 (N_15499,N_14381,N_14256);
or U15500 (N_15500,N_14880,N_14960);
nand U15501 (N_15501,N_14325,N_14761);
xor U15502 (N_15502,N_14888,N_14683);
nand U15503 (N_15503,N_14314,N_14657);
and U15504 (N_15504,N_14607,N_14541);
nor U15505 (N_15505,N_14112,N_14868);
xor U15506 (N_15506,N_14648,N_14431);
or U15507 (N_15507,N_14541,N_14220);
nand U15508 (N_15508,N_14988,N_14510);
and U15509 (N_15509,N_14133,N_14059);
or U15510 (N_15510,N_14929,N_14166);
or U15511 (N_15511,N_14309,N_14141);
or U15512 (N_15512,N_14268,N_14101);
or U15513 (N_15513,N_14342,N_14920);
or U15514 (N_15514,N_14858,N_14660);
xor U15515 (N_15515,N_14150,N_14461);
or U15516 (N_15516,N_14531,N_14743);
xnor U15517 (N_15517,N_14863,N_14620);
xnor U15518 (N_15518,N_14904,N_14483);
and U15519 (N_15519,N_14820,N_14267);
or U15520 (N_15520,N_14258,N_14607);
nand U15521 (N_15521,N_14157,N_14636);
nand U15522 (N_15522,N_14175,N_14917);
xnor U15523 (N_15523,N_14095,N_14501);
xor U15524 (N_15524,N_14702,N_14458);
nor U15525 (N_15525,N_14084,N_14719);
or U15526 (N_15526,N_14929,N_14827);
xor U15527 (N_15527,N_14490,N_14477);
or U15528 (N_15528,N_14403,N_14586);
or U15529 (N_15529,N_14840,N_14734);
nand U15530 (N_15530,N_14082,N_14912);
nand U15531 (N_15531,N_14471,N_14155);
and U15532 (N_15532,N_14824,N_14685);
nor U15533 (N_15533,N_14742,N_14947);
and U15534 (N_15534,N_14397,N_14879);
or U15535 (N_15535,N_14225,N_14472);
or U15536 (N_15536,N_14602,N_14041);
or U15537 (N_15537,N_14617,N_14295);
xor U15538 (N_15538,N_14913,N_14766);
nand U15539 (N_15539,N_14898,N_14661);
and U15540 (N_15540,N_14130,N_14926);
or U15541 (N_15541,N_14150,N_14312);
xor U15542 (N_15542,N_14117,N_14007);
nor U15543 (N_15543,N_14137,N_14966);
nand U15544 (N_15544,N_14066,N_14357);
nor U15545 (N_15545,N_14666,N_14902);
and U15546 (N_15546,N_14649,N_14815);
or U15547 (N_15547,N_14403,N_14721);
nor U15548 (N_15548,N_14912,N_14971);
xor U15549 (N_15549,N_14840,N_14381);
or U15550 (N_15550,N_14265,N_14878);
nor U15551 (N_15551,N_14601,N_14549);
or U15552 (N_15552,N_14327,N_14665);
or U15553 (N_15553,N_14658,N_14795);
xor U15554 (N_15554,N_14630,N_14216);
nor U15555 (N_15555,N_14076,N_14131);
nand U15556 (N_15556,N_14067,N_14330);
and U15557 (N_15557,N_14366,N_14448);
nor U15558 (N_15558,N_14254,N_14957);
nor U15559 (N_15559,N_14147,N_14042);
and U15560 (N_15560,N_14114,N_14560);
xnor U15561 (N_15561,N_14077,N_14786);
xor U15562 (N_15562,N_14486,N_14848);
nor U15563 (N_15563,N_14763,N_14409);
and U15564 (N_15564,N_14091,N_14191);
nand U15565 (N_15565,N_14927,N_14816);
nor U15566 (N_15566,N_14062,N_14021);
xor U15567 (N_15567,N_14309,N_14759);
or U15568 (N_15568,N_14168,N_14754);
or U15569 (N_15569,N_14714,N_14171);
xor U15570 (N_15570,N_14151,N_14740);
and U15571 (N_15571,N_14835,N_14802);
xnor U15572 (N_15572,N_14858,N_14963);
xnor U15573 (N_15573,N_14183,N_14714);
and U15574 (N_15574,N_14435,N_14568);
or U15575 (N_15575,N_14877,N_14769);
or U15576 (N_15576,N_14759,N_14298);
nand U15577 (N_15577,N_14997,N_14721);
and U15578 (N_15578,N_14847,N_14606);
and U15579 (N_15579,N_14863,N_14254);
nor U15580 (N_15580,N_14216,N_14506);
and U15581 (N_15581,N_14884,N_14380);
and U15582 (N_15582,N_14948,N_14687);
xor U15583 (N_15583,N_14500,N_14966);
nand U15584 (N_15584,N_14157,N_14970);
nand U15585 (N_15585,N_14381,N_14004);
and U15586 (N_15586,N_14782,N_14871);
xor U15587 (N_15587,N_14008,N_14825);
or U15588 (N_15588,N_14426,N_14748);
nand U15589 (N_15589,N_14632,N_14908);
xor U15590 (N_15590,N_14190,N_14287);
xnor U15591 (N_15591,N_14509,N_14442);
nor U15592 (N_15592,N_14490,N_14880);
nand U15593 (N_15593,N_14190,N_14035);
nand U15594 (N_15594,N_14197,N_14505);
and U15595 (N_15595,N_14895,N_14570);
xor U15596 (N_15596,N_14113,N_14558);
xor U15597 (N_15597,N_14633,N_14802);
and U15598 (N_15598,N_14256,N_14957);
and U15599 (N_15599,N_14584,N_14822);
and U15600 (N_15600,N_14790,N_14387);
and U15601 (N_15601,N_14966,N_14782);
or U15602 (N_15602,N_14433,N_14046);
and U15603 (N_15603,N_14755,N_14288);
nor U15604 (N_15604,N_14257,N_14928);
and U15605 (N_15605,N_14393,N_14941);
nor U15606 (N_15606,N_14091,N_14251);
nor U15607 (N_15607,N_14501,N_14408);
nor U15608 (N_15608,N_14882,N_14272);
or U15609 (N_15609,N_14515,N_14715);
or U15610 (N_15610,N_14227,N_14697);
and U15611 (N_15611,N_14755,N_14645);
nor U15612 (N_15612,N_14576,N_14932);
and U15613 (N_15613,N_14677,N_14728);
and U15614 (N_15614,N_14609,N_14559);
and U15615 (N_15615,N_14418,N_14554);
or U15616 (N_15616,N_14659,N_14654);
and U15617 (N_15617,N_14237,N_14604);
or U15618 (N_15618,N_14782,N_14026);
nand U15619 (N_15619,N_14954,N_14935);
or U15620 (N_15620,N_14052,N_14398);
or U15621 (N_15621,N_14794,N_14632);
nand U15622 (N_15622,N_14304,N_14191);
nand U15623 (N_15623,N_14967,N_14256);
or U15624 (N_15624,N_14658,N_14763);
nor U15625 (N_15625,N_14110,N_14070);
xor U15626 (N_15626,N_14300,N_14766);
and U15627 (N_15627,N_14269,N_14127);
or U15628 (N_15628,N_14107,N_14264);
or U15629 (N_15629,N_14245,N_14835);
and U15630 (N_15630,N_14570,N_14569);
and U15631 (N_15631,N_14336,N_14241);
or U15632 (N_15632,N_14014,N_14641);
and U15633 (N_15633,N_14840,N_14317);
nor U15634 (N_15634,N_14843,N_14245);
and U15635 (N_15635,N_14111,N_14237);
nand U15636 (N_15636,N_14603,N_14383);
nor U15637 (N_15637,N_14203,N_14416);
nand U15638 (N_15638,N_14121,N_14575);
nor U15639 (N_15639,N_14143,N_14698);
nand U15640 (N_15640,N_14598,N_14875);
nor U15641 (N_15641,N_14526,N_14458);
or U15642 (N_15642,N_14179,N_14024);
and U15643 (N_15643,N_14359,N_14569);
and U15644 (N_15644,N_14972,N_14138);
nor U15645 (N_15645,N_14457,N_14052);
nor U15646 (N_15646,N_14465,N_14633);
nor U15647 (N_15647,N_14029,N_14375);
nor U15648 (N_15648,N_14272,N_14128);
nand U15649 (N_15649,N_14815,N_14091);
nand U15650 (N_15650,N_14634,N_14740);
xor U15651 (N_15651,N_14371,N_14225);
xor U15652 (N_15652,N_14501,N_14684);
nand U15653 (N_15653,N_14361,N_14276);
nor U15654 (N_15654,N_14492,N_14647);
nor U15655 (N_15655,N_14221,N_14157);
or U15656 (N_15656,N_14459,N_14696);
and U15657 (N_15657,N_14627,N_14821);
nand U15658 (N_15658,N_14275,N_14597);
xor U15659 (N_15659,N_14712,N_14992);
or U15660 (N_15660,N_14420,N_14509);
nor U15661 (N_15661,N_14083,N_14623);
or U15662 (N_15662,N_14439,N_14313);
or U15663 (N_15663,N_14067,N_14006);
nand U15664 (N_15664,N_14755,N_14629);
xnor U15665 (N_15665,N_14733,N_14008);
or U15666 (N_15666,N_14226,N_14466);
nor U15667 (N_15667,N_14248,N_14182);
xnor U15668 (N_15668,N_14850,N_14191);
and U15669 (N_15669,N_14754,N_14817);
and U15670 (N_15670,N_14508,N_14168);
nand U15671 (N_15671,N_14734,N_14894);
nor U15672 (N_15672,N_14355,N_14778);
or U15673 (N_15673,N_14424,N_14005);
xnor U15674 (N_15674,N_14579,N_14783);
or U15675 (N_15675,N_14869,N_14349);
or U15676 (N_15676,N_14371,N_14485);
or U15677 (N_15677,N_14374,N_14228);
nor U15678 (N_15678,N_14837,N_14198);
nand U15679 (N_15679,N_14272,N_14254);
xor U15680 (N_15680,N_14182,N_14151);
or U15681 (N_15681,N_14254,N_14019);
or U15682 (N_15682,N_14014,N_14438);
or U15683 (N_15683,N_14182,N_14527);
nor U15684 (N_15684,N_14710,N_14791);
nand U15685 (N_15685,N_14455,N_14291);
xor U15686 (N_15686,N_14866,N_14727);
and U15687 (N_15687,N_14538,N_14937);
nor U15688 (N_15688,N_14093,N_14744);
xor U15689 (N_15689,N_14178,N_14944);
xnor U15690 (N_15690,N_14688,N_14425);
nand U15691 (N_15691,N_14394,N_14269);
xor U15692 (N_15692,N_14043,N_14284);
or U15693 (N_15693,N_14638,N_14826);
or U15694 (N_15694,N_14544,N_14684);
and U15695 (N_15695,N_14432,N_14106);
nand U15696 (N_15696,N_14535,N_14172);
nor U15697 (N_15697,N_14028,N_14172);
nor U15698 (N_15698,N_14350,N_14507);
and U15699 (N_15699,N_14240,N_14793);
and U15700 (N_15700,N_14122,N_14265);
xnor U15701 (N_15701,N_14215,N_14943);
nor U15702 (N_15702,N_14251,N_14680);
and U15703 (N_15703,N_14490,N_14879);
and U15704 (N_15704,N_14337,N_14054);
nand U15705 (N_15705,N_14908,N_14359);
and U15706 (N_15706,N_14820,N_14198);
nor U15707 (N_15707,N_14331,N_14113);
nor U15708 (N_15708,N_14990,N_14454);
or U15709 (N_15709,N_14354,N_14041);
nand U15710 (N_15710,N_14684,N_14051);
or U15711 (N_15711,N_14839,N_14785);
nand U15712 (N_15712,N_14665,N_14918);
xnor U15713 (N_15713,N_14830,N_14509);
and U15714 (N_15714,N_14820,N_14177);
xor U15715 (N_15715,N_14852,N_14389);
or U15716 (N_15716,N_14737,N_14788);
xnor U15717 (N_15717,N_14819,N_14859);
nand U15718 (N_15718,N_14635,N_14696);
nand U15719 (N_15719,N_14101,N_14339);
and U15720 (N_15720,N_14377,N_14000);
or U15721 (N_15721,N_14653,N_14096);
nand U15722 (N_15722,N_14432,N_14894);
or U15723 (N_15723,N_14073,N_14930);
xnor U15724 (N_15724,N_14181,N_14623);
and U15725 (N_15725,N_14558,N_14798);
nor U15726 (N_15726,N_14391,N_14831);
or U15727 (N_15727,N_14941,N_14158);
nor U15728 (N_15728,N_14198,N_14155);
or U15729 (N_15729,N_14328,N_14503);
nor U15730 (N_15730,N_14775,N_14257);
or U15731 (N_15731,N_14013,N_14912);
xor U15732 (N_15732,N_14884,N_14004);
xor U15733 (N_15733,N_14916,N_14948);
or U15734 (N_15734,N_14288,N_14757);
xor U15735 (N_15735,N_14320,N_14122);
and U15736 (N_15736,N_14226,N_14519);
nand U15737 (N_15737,N_14269,N_14743);
or U15738 (N_15738,N_14454,N_14039);
and U15739 (N_15739,N_14038,N_14985);
and U15740 (N_15740,N_14249,N_14577);
nand U15741 (N_15741,N_14265,N_14511);
nand U15742 (N_15742,N_14231,N_14578);
nand U15743 (N_15743,N_14305,N_14126);
nor U15744 (N_15744,N_14796,N_14088);
or U15745 (N_15745,N_14557,N_14272);
or U15746 (N_15746,N_14367,N_14317);
nand U15747 (N_15747,N_14120,N_14898);
and U15748 (N_15748,N_14407,N_14436);
xor U15749 (N_15749,N_14126,N_14537);
and U15750 (N_15750,N_14074,N_14006);
and U15751 (N_15751,N_14162,N_14667);
or U15752 (N_15752,N_14962,N_14259);
or U15753 (N_15753,N_14647,N_14546);
nor U15754 (N_15754,N_14774,N_14623);
or U15755 (N_15755,N_14668,N_14273);
xor U15756 (N_15756,N_14228,N_14749);
nand U15757 (N_15757,N_14326,N_14463);
and U15758 (N_15758,N_14634,N_14172);
or U15759 (N_15759,N_14552,N_14547);
and U15760 (N_15760,N_14068,N_14011);
and U15761 (N_15761,N_14268,N_14727);
nor U15762 (N_15762,N_14486,N_14337);
nand U15763 (N_15763,N_14151,N_14835);
nor U15764 (N_15764,N_14150,N_14145);
nor U15765 (N_15765,N_14425,N_14514);
nand U15766 (N_15766,N_14011,N_14136);
or U15767 (N_15767,N_14657,N_14428);
xor U15768 (N_15768,N_14585,N_14894);
or U15769 (N_15769,N_14202,N_14286);
nand U15770 (N_15770,N_14682,N_14865);
nand U15771 (N_15771,N_14191,N_14567);
xnor U15772 (N_15772,N_14681,N_14367);
nand U15773 (N_15773,N_14044,N_14156);
xnor U15774 (N_15774,N_14424,N_14631);
or U15775 (N_15775,N_14315,N_14944);
and U15776 (N_15776,N_14843,N_14818);
nor U15777 (N_15777,N_14750,N_14637);
nor U15778 (N_15778,N_14303,N_14240);
nand U15779 (N_15779,N_14897,N_14896);
xnor U15780 (N_15780,N_14589,N_14242);
nor U15781 (N_15781,N_14728,N_14393);
and U15782 (N_15782,N_14873,N_14246);
nor U15783 (N_15783,N_14333,N_14156);
nand U15784 (N_15784,N_14066,N_14911);
or U15785 (N_15785,N_14597,N_14702);
xnor U15786 (N_15786,N_14216,N_14055);
and U15787 (N_15787,N_14388,N_14818);
and U15788 (N_15788,N_14825,N_14894);
nand U15789 (N_15789,N_14878,N_14770);
nand U15790 (N_15790,N_14167,N_14739);
xor U15791 (N_15791,N_14332,N_14736);
and U15792 (N_15792,N_14844,N_14650);
nand U15793 (N_15793,N_14699,N_14589);
nand U15794 (N_15794,N_14315,N_14591);
nor U15795 (N_15795,N_14425,N_14694);
xnor U15796 (N_15796,N_14338,N_14738);
nand U15797 (N_15797,N_14222,N_14834);
nand U15798 (N_15798,N_14742,N_14121);
nand U15799 (N_15799,N_14938,N_14087);
nor U15800 (N_15800,N_14224,N_14753);
nor U15801 (N_15801,N_14778,N_14342);
nor U15802 (N_15802,N_14711,N_14920);
nor U15803 (N_15803,N_14620,N_14652);
or U15804 (N_15804,N_14440,N_14040);
and U15805 (N_15805,N_14640,N_14444);
xor U15806 (N_15806,N_14321,N_14844);
xor U15807 (N_15807,N_14519,N_14197);
nor U15808 (N_15808,N_14330,N_14287);
xor U15809 (N_15809,N_14913,N_14551);
nand U15810 (N_15810,N_14993,N_14035);
nand U15811 (N_15811,N_14686,N_14585);
or U15812 (N_15812,N_14720,N_14791);
nand U15813 (N_15813,N_14201,N_14315);
nor U15814 (N_15814,N_14073,N_14105);
nand U15815 (N_15815,N_14796,N_14797);
nand U15816 (N_15816,N_14480,N_14997);
nand U15817 (N_15817,N_14666,N_14740);
xnor U15818 (N_15818,N_14879,N_14486);
and U15819 (N_15819,N_14132,N_14356);
nor U15820 (N_15820,N_14183,N_14530);
nor U15821 (N_15821,N_14907,N_14337);
or U15822 (N_15822,N_14154,N_14135);
nor U15823 (N_15823,N_14615,N_14058);
xor U15824 (N_15824,N_14280,N_14655);
or U15825 (N_15825,N_14441,N_14252);
nor U15826 (N_15826,N_14378,N_14556);
nor U15827 (N_15827,N_14502,N_14159);
nor U15828 (N_15828,N_14837,N_14862);
nor U15829 (N_15829,N_14543,N_14813);
and U15830 (N_15830,N_14972,N_14564);
or U15831 (N_15831,N_14739,N_14684);
or U15832 (N_15832,N_14484,N_14216);
nor U15833 (N_15833,N_14897,N_14389);
xor U15834 (N_15834,N_14989,N_14106);
nor U15835 (N_15835,N_14258,N_14912);
nor U15836 (N_15836,N_14871,N_14074);
or U15837 (N_15837,N_14701,N_14860);
nor U15838 (N_15838,N_14913,N_14851);
and U15839 (N_15839,N_14353,N_14506);
and U15840 (N_15840,N_14247,N_14188);
nand U15841 (N_15841,N_14891,N_14643);
and U15842 (N_15842,N_14289,N_14655);
or U15843 (N_15843,N_14474,N_14946);
and U15844 (N_15844,N_14304,N_14523);
nor U15845 (N_15845,N_14351,N_14381);
nand U15846 (N_15846,N_14274,N_14579);
nor U15847 (N_15847,N_14265,N_14039);
nand U15848 (N_15848,N_14454,N_14059);
nor U15849 (N_15849,N_14260,N_14975);
nor U15850 (N_15850,N_14027,N_14886);
nand U15851 (N_15851,N_14506,N_14905);
and U15852 (N_15852,N_14096,N_14195);
xnor U15853 (N_15853,N_14273,N_14803);
or U15854 (N_15854,N_14350,N_14479);
nand U15855 (N_15855,N_14489,N_14140);
or U15856 (N_15856,N_14374,N_14338);
or U15857 (N_15857,N_14866,N_14995);
xnor U15858 (N_15858,N_14834,N_14182);
and U15859 (N_15859,N_14099,N_14260);
xor U15860 (N_15860,N_14560,N_14397);
and U15861 (N_15861,N_14304,N_14364);
or U15862 (N_15862,N_14255,N_14772);
nor U15863 (N_15863,N_14109,N_14405);
xor U15864 (N_15864,N_14712,N_14034);
xnor U15865 (N_15865,N_14872,N_14930);
or U15866 (N_15866,N_14533,N_14406);
and U15867 (N_15867,N_14489,N_14580);
or U15868 (N_15868,N_14697,N_14921);
nand U15869 (N_15869,N_14726,N_14317);
xor U15870 (N_15870,N_14281,N_14841);
xor U15871 (N_15871,N_14618,N_14378);
xor U15872 (N_15872,N_14019,N_14078);
xor U15873 (N_15873,N_14791,N_14594);
and U15874 (N_15874,N_14024,N_14375);
xor U15875 (N_15875,N_14446,N_14125);
and U15876 (N_15876,N_14271,N_14955);
and U15877 (N_15877,N_14590,N_14209);
nor U15878 (N_15878,N_14962,N_14835);
and U15879 (N_15879,N_14258,N_14019);
xnor U15880 (N_15880,N_14120,N_14069);
xor U15881 (N_15881,N_14179,N_14610);
and U15882 (N_15882,N_14750,N_14357);
nor U15883 (N_15883,N_14655,N_14972);
or U15884 (N_15884,N_14169,N_14793);
nand U15885 (N_15885,N_14306,N_14948);
or U15886 (N_15886,N_14977,N_14625);
or U15887 (N_15887,N_14218,N_14593);
nor U15888 (N_15888,N_14893,N_14147);
or U15889 (N_15889,N_14227,N_14470);
nor U15890 (N_15890,N_14593,N_14940);
and U15891 (N_15891,N_14362,N_14261);
and U15892 (N_15892,N_14322,N_14260);
nor U15893 (N_15893,N_14910,N_14816);
or U15894 (N_15894,N_14539,N_14242);
xor U15895 (N_15895,N_14274,N_14120);
and U15896 (N_15896,N_14711,N_14727);
or U15897 (N_15897,N_14100,N_14214);
nor U15898 (N_15898,N_14271,N_14861);
xnor U15899 (N_15899,N_14575,N_14728);
and U15900 (N_15900,N_14800,N_14003);
nand U15901 (N_15901,N_14672,N_14248);
xor U15902 (N_15902,N_14093,N_14671);
or U15903 (N_15903,N_14112,N_14079);
or U15904 (N_15904,N_14333,N_14502);
and U15905 (N_15905,N_14972,N_14606);
xor U15906 (N_15906,N_14638,N_14410);
or U15907 (N_15907,N_14701,N_14511);
and U15908 (N_15908,N_14356,N_14075);
nor U15909 (N_15909,N_14287,N_14118);
nand U15910 (N_15910,N_14876,N_14529);
and U15911 (N_15911,N_14912,N_14231);
and U15912 (N_15912,N_14983,N_14528);
nand U15913 (N_15913,N_14440,N_14917);
nor U15914 (N_15914,N_14935,N_14381);
or U15915 (N_15915,N_14928,N_14191);
nor U15916 (N_15916,N_14400,N_14634);
or U15917 (N_15917,N_14215,N_14156);
or U15918 (N_15918,N_14279,N_14886);
and U15919 (N_15919,N_14676,N_14379);
or U15920 (N_15920,N_14868,N_14441);
or U15921 (N_15921,N_14401,N_14030);
and U15922 (N_15922,N_14997,N_14127);
nand U15923 (N_15923,N_14908,N_14311);
nor U15924 (N_15924,N_14321,N_14663);
or U15925 (N_15925,N_14281,N_14667);
xor U15926 (N_15926,N_14433,N_14922);
nand U15927 (N_15927,N_14642,N_14137);
nand U15928 (N_15928,N_14013,N_14178);
nand U15929 (N_15929,N_14749,N_14085);
xor U15930 (N_15930,N_14772,N_14317);
xor U15931 (N_15931,N_14864,N_14048);
nand U15932 (N_15932,N_14432,N_14697);
or U15933 (N_15933,N_14927,N_14433);
and U15934 (N_15934,N_14530,N_14366);
or U15935 (N_15935,N_14228,N_14798);
or U15936 (N_15936,N_14910,N_14581);
and U15937 (N_15937,N_14840,N_14862);
xor U15938 (N_15938,N_14941,N_14587);
and U15939 (N_15939,N_14017,N_14126);
xor U15940 (N_15940,N_14996,N_14196);
nor U15941 (N_15941,N_14156,N_14541);
and U15942 (N_15942,N_14544,N_14657);
nor U15943 (N_15943,N_14400,N_14877);
or U15944 (N_15944,N_14505,N_14714);
nand U15945 (N_15945,N_14750,N_14109);
nand U15946 (N_15946,N_14761,N_14906);
or U15947 (N_15947,N_14119,N_14734);
xnor U15948 (N_15948,N_14519,N_14906);
nor U15949 (N_15949,N_14873,N_14255);
and U15950 (N_15950,N_14780,N_14190);
and U15951 (N_15951,N_14228,N_14676);
and U15952 (N_15952,N_14533,N_14384);
and U15953 (N_15953,N_14743,N_14082);
nor U15954 (N_15954,N_14052,N_14005);
nor U15955 (N_15955,N_14244,N_14461);
or U15956 (N_15956,N_14999,N_14128);
nor U15957 (N_15957,N_14270,N_14243);
nand U15958 (N_15958,N_14547,N_14003);
xor U15959 (N_15959,N_14239,N_14500);
nor U15960 (N_15960,N_14183,N_14138);
xor U15961 (N_15961,N_14518,N_14804);
nand U15962 (N_15962,N_14110,N_14539);
xor U15963 (N_15963,N_14183,N_14348);
nand U15964 (N_15964,N_14755,N_14786);
nor U15965 (N_15965,N_14718,N_14834);
and U15966 (N_15966,N_14654,N_14128);
xor U15967 (N_15967,N_14360,N_14293);
nand U15968 (N_15968,N_14907,N_14047);
nand U15969 (N_15969,N_14122,N_14108);
or U15970 (N_15970,N_14155,N_14200);
nor U15971 (N_15971,N_14123,N_14652);
xor U15972 (N_15972,N_14651,N_14027);
nor U15973 (N_15973,N_14976,N_14135);
or U15974 (N_15974,N_14249,N_14632);
nand U15975 (N_15975,N_14923,N_14233);
or U15976 (N_15976,N_14730,N_14780);
nand U15977 (N_15977,N_14373,N_14638);
and U15978 (N_15978,N_14184,N_14230);
nand U15979 (N_15979,N_14427,N_14405);
nand U15980 (N_15980,N_14451,N_14684);
and U15981 (N_15981,N_14320,N_14801);
or U15982 (N_15982,N_14919,N_14802);
or U15983 (N_15983,N_14889,N_14700);
or U15984 (N_15984,N_14205,N_14713);
xnor U15985 (N_15985,N_14403,N_14471);
xor U15986 (N_15986,N_14989,N_14121);
nand U15987 (N_15987,N_14870,N_14339);
and U15988 (N_15988,N_14466,N_14937);
and U15989 (N_15989,N_14730,N_14323);
nand U15990 (N_15990,N_14036,N_14762);
or U15991 (N_15991,N_14324,N_14620);
nor U15992 (N_15992,N_14170,N_14890);
or U15993 (N_15993,N_14523,N_14020);
nand U15994 (N_15994,N_14368,N_14383);
nor U15995 (N_15995,N_14085,N_14091);
or U15996 (N_15996,N_14686,N_14457);
and U15997 (N_15997,N_14111,N_14838);
xnor U15998 (N_15998,N_14336,N_14862);
and U15999 (N_15999,N_14573,N_14799);
or U16000 (N_16000,N_15258,N_15753);
and U16001 (N_16001,N_15348,N_15901);
and U16002 (N_16002,N_15519,N_15131);
and U16003 (N_16003,N_15745,N_15398);
and U16004 (N_16004,N_15953,N_15528);
and U16005 (N_16005,N_15313,N_15473);
nand U16006 (N_16006,N_15713,N_15161);
xor U16007 (N_16007,N_15707,N_15891);
and U16008 (N_16008,N_15344,N_15459);
xor U16009 (N_16009,N_15168,N_15098);
or U16010 (N_16010,N_15133,N_15309);
xor U16011 (N_16011,N_15379,N_15107);
xnor U16012 (N_16012,N_15765,N_15173);
xor U16013 (N_16013,N_15251,N_15302);
or U16014 (N_16014,N_15439,N_15125);
and U16015 (N_16015,N_15254,N_15896);
nand U16016 (N_16016,N_15962,N_15598);
nand U16017 (N_16017,N_15867,N_15204);
and U16018 (N_16018,N_15362,N_15038);
xnor U16019 (N_16019,N_15829,N_15921);
xnor U16020 (N_16020,N_15400,N_15821);
and U16021 (N_16021,N_15672,N_15194);
nor U16022 (N_16022,N_15925,N_15682);
and U16023 (N_16023,N_15832,N_15044);
nor U16024 (N_16024,N_15620,N_15421);
nor U16025 (N_16025,N_15551,N_15010);
xor U16026 (N_16026,N_15074,N_15675);
or U16027 (N_16027,N_15640,N_15630);
or U16028 (N_16028,N_15319,N_15604);
nand U16029 (N_16029,N_15082,N_15160);
xor U16030 (N_16030,N_15422,N_15142);
nand U16031 (N_16031,N_15690,N_15474);
xnor U16032 (N_16032,N_15547,N_15288);
nand U16033 (N_16033,N_15000,N_15294);
nor U16034 (N_16034,N_15565,N_15138);
nand U16035 (N_16035,N_15412,N_15004);
nand U16036 (N_16036,N_15226,N_15911);
and U16037 (N_16037,N_15240,N_15648);
xnor U16038 (N_16038,N_15023,N_15156);
xnor U16039 (N_16039,N_15043,N_15747);
or U16040 (N_16040,N_15453,N_15637);
nand U16041 (N_16041,N_15740,N_15213);
and U16042 (N_16042,N_15202,N_15402);
nor U16043 (N_16043,N_15314,N_15008);
xnor U16044 (N_16044,N_15979,N_15242);
nand U16045 (N_16045,N_15900,N_15777);
or U16046 (N_16046,N_15817,N_15292);
xnor U16047 (N_16047,N_15636,N_15062);
and U16048 (N_16048,N_15550,N_15358);
nor U16049 (N_16049,N_15255,N_15115);
nor U16050 (N_16050,N_15933,N_15522);
and U16051 (N_16051,N_15558,N_15337);
nor U16052 (N_16052,N_15529,N_15413);
xnor U16053 (N_16053,N_15723,N_15660);
and U16054 (N_16054,N_15375,N_15606);
nor U16055 (N_16055,N_15846,N_15795);
or U16056 (N_16056,N_15643,N_15757);
xor U16057 (N_16057,N_15289,N_15336);
or U16058 (N_16058,N_15789,N_15866);
nor U16059 (N_16059,N_15657,N_15322);
nand U16060 (N_16060,N_15340,N_15241);
and U16061 (N_16061,N_15441,N_15615);
nor U16062 (N_16062,N_15356,N_15075);
nor U16063 (N_16063,N_15404,N_15720);
xnor U16064 (N_16064,N_15633,N_15596);
xnor U16065 (N_16065,N_15500,N_15345);
and U16066 (N_16066,N_15080,N_15124);
or U16067 (N_16067,N_15097,N_15834);
and U16068 (N_16068,N_15256,N_15739);
or U16069 (N_16069,N_15151,N_15121);
nor U16070 (N_16070,N_15079,N_15912);
and U16071 (N_16071,N_15452,N_15868);
nand U16072 (N_16072,N_15715,N_15166);
nand U16073 (N_16073,N_15048,N_15132);
xor U16074 (N_16074,N_15666,N_15238);
and U16075 (N_16075,N_15839,N_15188);
xnor U16076 (N_16076,N_15355,N_15897);
or U16077 (N_16077,N_15792,N_15683);
nor U16078 (N_16078,N_15399,N_15759);
nand U16079 (N_16079,N_15786,N_15481);
xnor U16080 (N_16080,N_15686,N_15949);
xnor U16081 (N_16081,N_15510,N_15197);
or U16082 (N_16082,N_15857,N_15754);
xnor U16083 (N_16083,N_15814,N_15272);
and U16084 (N_16084,N_15673,N_15874);
xor U16085 (N_16085,N_15719,N_15527);
nand U16086 (N_16086,N_15969,N_15093);
nor U16087 (N_16087,N_15141,N_15948);
nor U16088 (N_16088,N_15028,N_15489);
and U16089 (N_16089,N_15600,N_15128);
or U16090 (N_16090,N_15718,N_15437);
or U16091 (N_16091,N_15454,N_15626);
nor U16092 (N_16092,N_15996,N_15982);
nand U16093 (N_16093,N_15011,N_15172);
or U16094 (N_16094,N_15861,N_15582);
xor U16095 (N_16095,N_15350,N_15416);
xor U16096 (N_16096,N_15650,N_15271);
xor U16097 (N_16097,N_15099,N_15091);
nand U16098 (N_16098,N_15518,N_15105);
and U16099 (N_16099,N_15317,N_15877);
nor U16100 (N_16100,N_15257,N_15072);
nand U16101 (N_16101,N_15705,N_15931);
or U16102 (N_16102,N_15059,N_15954);
nand U16103 (N_16103,N_15543,N_15102);
nand U16104 (N_16104,N_15248,N_15684);
xnor U16105 (N_16105,N_15590,N_15076);
nand U16106 (N_16106,N_15656,N_15065);
and U16107 (N_16107,N_15864,N_15957);
nor U16108 (N_16108,N_15992,N_15120);
xnor U16109 (N_16109,N_15273,N_15746);
and U16110 (N_16110,N_15343,N_15774);
nor U16111 (N_16111,N_15070,N_15902);
xor U16112 (N_16112,N_15117,N_15246);
nand U16113 (N_16113,N_15499,N_15155);
nor U16114 (N_16114,N_15333,N_15185);
nor U16115 (N_16115,N_15895,N_15200);
nor U16116 (N_16116,N_15974,N_15503);
nand U16117 (N_16117,N_15595,N_15649);
or U16118 (N_16118,N_15995,N_15784);
nor U16119 (N_16119,N_15041,N_15735);
nor U16120 (N_16120,N_15951,N_15351);
xnor U16121 (N_16121,N_15881,N_15009);
and U16122 (N_16122,N_15150,N_15145);
nor U16123 (N_16123,N_15870,N_15616);
nand U16124 (N_16124,N_15234,N_15052);
nand U16125 (N_16125,N_15377,N_15799);
xnor U16126 (N_16126,N_15963,N_15619);
and U16127 (N_16127,N_15396,N_15614);
xor U16128 (N_16128,N_15629,N_15808);
and U16129 (N_16129,N_15081,N_15129);
nand U16130 (N_16130,N_15899,N_15100);
nor U16131 (N_16131,N_15894,N_15661);
or U16132 (N_16132,N_15594,N_15118);
or U16133 (N_16133,N_15553,N_15176);
or U16134 (N_16134,N_15110,N_15077);
or U16135 (N_16135,N_15512,N_15823);
xnor U16136 (N_16136,N_15915,N_15893);
nor U16137 (N_16137,N_15884,N_15712);
nand U16138 (N_16138,N_15687,N_15970);
nand U16139 (N_16139,N_15461,N_15094);
or U16140 (N_16140,N_15722,N_15019);
or U16141 (N_16141,N_15483,N_15736);
nand U16142 (N_16142,N_15042,N_15169);
and U16143 (N_16143,N_15670,N_15793);
nor U16144 (N_16144,N_15725,N_15303);
xor U16145 (N_16145,N_15269,N_15212);
and U16146 (N_16146,N_15390,N_15385);
nand U16147 (N_16147,N_15498,N_15549);
xnor U16148 (N_16148,N_15423,N_15794);
or U16149 (N_16149,N_15732,N_15270);
nor U16150 (N_16150,N_15488,N_15451);
xnor U16151 (N_16151,N_15365,N_15984);
or U16152 (N_16152,N_15395,N_15943);
nand U16153 (N_16153,N_15930,N_15628);
and U16154 (N_16154,N_15205,N_15658);
and U16155 (N_16155,N_15146,N_15627);
nor U16156 (N_16156,N_15490,N_15371);
nor U16157 (N_16157,N_15993,N_15905);
and U16158 (N_16158,N_15986,N_15575);
or U16159 (N_16159,N_15158,N_15665);
and U16160 (N_16160,N_15852,N_15985);
xnor U16161 (N_16161,N_15427,N_15015);
and U16162 (N_16162,N_15659,N_15181);
nand U16163 (N_16163,N_15991,N_15280);
nor U16164 (N_16164,N_15177,N_15261);
xnor U16165 (N_16165,N_15007,N_15856);
xor U16166 (N_16166,N_15126,N_15298);
nand U16167 (N_16167,N_15005,N_15484);
nand U16168 (N_16168,N_15946,N_15468);
or U16169 (N_16169,N_15316,N_15406);
and U16170 (N_16170,N_15112,N_15137);
nand U16171 (N_16171,N_15171,N_15444);
nor U16172 (N_16172,N_15806,N_15493);
xnor U16173 (N_16173,N_15039,N_15278);
xnor U16174 (N_16174,N_15609,N_15655);
nand U16175 (N_16175,N_15539,N_15123);
or U16176 (N_16176,N_15116,N_15165);
and U16177 (N_16177,N_15699,N_15342);
nand U16178 (N_16178,N_15618,N_15942);
nor U16179 (N_16179,N_15597,N_15378);
nor U16180 (N_16180,N_15728,N_15347);
xnor U16181 (N_16181,N_15223,N_15192);
nor U16182 (N_16182,N_15443,N_15083);
xor U16183 (N_16183,N_15321,N_15469);
nand U16184 (N_16184,N_15583,N_15762);
and U16185 (N_16185,N_15002,N_15357);
or U16186 (N_16186,N_15608,N_15859);
nor U16187 (N_16187,N_15782,N_15387);
nand U16188 (N_16188,N_15230,N_15965);
or U16189 (N_16189,N_15642,N_15935);
nand U16190 (N_16190,N_15601,N_15369);
or U16191 (N_16191,N_15036,N_15758);
xor U16192 (N_16192,N_15103,N_15460);
xnor U16193 (N_16193,N_15523,N_15353);
nand U16194 (N_16194,N_15940,N_15632);
nor U16195 (N_16195,N_15383,N_15865);
xor U16196 (N_16196,N_15752,N_15088);
nand U16197 (N_16197,N_15729,N_15652);
nor U16198 (N_16198,N_15694,N_15875);
nor U16199 (N_16199,N_15981,N_15361);
and U16200 (N_16200,N_15624,N_15898);
nor U16201 (N_16201,N_15195,N_15730);
or U16202 (N_16202,N_15664,N_15878);
xnor U16203 (N_16203,N_15513,N_15825);
nor U16204 (N_16204,N_15214,N_15971);
and U16205 (N_16205,N_15307,N_15959);
nand U16206 (N_16206,N_15190,N_15928);
xnor U16207 (N_16207,N_15136,N_15738);
or U16208 (N_16208,N_15464,N_15880);
and U16209 (N_16209,N_15446,N_15085);
nor U16210 (N_16210,N_15833,N_15061);
nor U16211 (N_16211,N_15693,N_15811);
nor U16212 (N_16212,N_15046,N_15462);
nor U16213 (N_16213,N_15668,N_15134);
and U16214 (N_16214,N_15162,N_15850);
or U16215 (N_16215,N_15836,N_15678);
and U16216 (N_16216,N_15835,N_15231);
nor U16217 (N_16217,N_15170,N_15574);
and U16218 (N_16218,N_15847,N_15026);
nor U16219 (N_16219,N_15457,N_15717);
nand U16220 (N_16220,N_15635,N_15411);
nor U16221 (N_16221,N_15521,N_15324);
nor U16222 (N_16222,N_15841,N_15370);
and U16223 (N_16223,N_15610,N_15696);
and U16224 (N_16224,N_15977,N_15653);
xor U16225 (N_16225,N_15560,N_15175);
and U16226 (N_16226,N_15003,N_15688);
and U16227 (N_16227,N_15929,N_15767);
xnor U16228 (N_16228,N_15561,N_15702);
and U16229 (N_16229,N_15709,N_15714);
or U16230 (N_16230,N_15537,N_15056);
xnor U16231 (N_16231,N_15584,N_15703);
or U16232 (N_16232,N_15389,N_15785);
xor U16233 (N_16233,N_15871,N_15196);
xnor U16234 (N_16234,N_15631,N_15566);
or U16235 (N_16235,N_15926,N_15382);
and U16236 (N_16236,N_15955,N_15997);
and U16237 (N_16237,N_15320,N_15944);
nor U16238 (N_16238,N_15546,N_15140);
xnor U16239 (N_16239,N_15809,N_15851);
nand U16240 (N_16240,N_15266,N_15711);
nand U16241 (N_16241,N_15299,N_15221);
xor U16242 (N_16242,N_15191,N_15305);
nor U16243 (N_16243,N_15024,N_15679);
nor U16244 (N_16244,N_15477,N_15989);
nand U16245 (N_16245,N_15526,N_15647);
or U16246 (N_16246,N_15069,N_15936);
nor U16247 (N_16247,N_15207,N_15958);
or U16248 (N_16248,N_15047,N_15506);
or U16249 (N_16249,N_15780,N_15826);
or U16250 (N_16250,N_15491,N_15232);
xor U16251 (N_16251,N_15586,N_15667);
and U16252 (N_16252,N_15611,N_15397);
nand U16253 (N_16253,N_15530,N_15224);
xnor U16254 (N_16254,N_15095,N_15332);
and U16255 (N_16255,N_15950,N_15496);
nand U16256 (N_16256,N_15433,N_15922);
nand U16257 (N_16257,N_15927,N_15127);
nand U16258 (N_16258,N_15710,N_15695);
nor U16259 (N_16259,N_15068,N_15978);
nor U16260 (N_16260,N_15564,N_15029);
and U16261 (N_16261,N_15148,N_15589);
and U16262 (N_16262,N_15700,N_15578);
nor U16263 (N_16263,N_15910,N_15143);
nor U16264 (N_16264,N_15612,N_15532);
xnor U16265 (N_16265,N_15265,N_15691);
and U16266 (N_16266,N_15426,N_15677);
and U16267 (N_16267,N_15050,N_15516);
and U16268 (N_16268,N_15287,N_15308);
or U16269 (N_16269,N_15135,N_15297);
and U16270 (N_16270,N_15438,N_15435);
and U16271 (N_16271,N_15517,N_15791);
nand U16272 (N_16272,N_15034,N_15286);
and U16273 (N_16273,N_15554,N_15227);
xnor U16274 (N_16274,N_15078,N_15108);
or U16275 (N_16275,N_15283,N_15854);
nor U16276 (N_16276,N_15961,N_15244);
xor U16277 (N_16277,N_15450,N_15934);
nand U16278 (N_16278,N_15327,N_15312);
nand U16279 (N_16279,N_15486,N_15639);
or U16280 (N_16280,N_15372,N_15101);
and U16281 (N_16281,N_15281,N_15033);
or U16282 (N_16282,N_15781,N_15704);
nand U16283 (N_16283,N_15556,N_15674);
or U16284 (N_16284,N_15054,N_15159);
nor U16285 (N_16285,N_15084,N_15276);
or U16286 (N_16286,N_15359,N_15284);
or U16287 (N_16287,N_15907,N_15051);
or U16288 (N_16288,N_15300,N_15587);
xor U16289 (N_16289,N_15018,N_15139);
xnor U16290 (N_16290,N_15764,N_15178);
xor U16291 (N_16291,N_15755,N_15634);
or U16292 (N_16292,N_15701,N_15275);
or U16293 (N_16293,N_15206,N_15844);
nand U16294 (N_16294,N_15726,N_15027);
xor U16295 (N_16295,N_15778,N_15455);
nor U16296 (N_16296,N_15769,N_15032);
and U16297 (N_16297,N_15838,N_15417);
or U16298 (N_16298,N_15163,N_15973);
xnor U16299 (N_16299,N_15576,N_15721);
nor U16300 (N_16300,N_15964,N_15538);
or U16301 (N_16301,N_15064,N_15233);
nand U16302 (N_16302,N_15603,N_15222);
and U16303 (N_16303,N_15827,N_15282);
nor U16304 (N_16304,N_15779,N_15274);
and U16305 (N_16305,N_15917,N_15685);
xnor U16306 (N_16306,N_15149,N_15198);
xor U16307 (N_16307,N_15890,N_15252);
or U16308 (N_16308,N_15906,N_15253);
nor U16309 (N_16309,N_15339,N_15025);
or U16310 (N_16310,N_15733,N_15815);
nand U16311 (N_16311,N_15239,N_15772);
nand U16312 (N_16312,N_15579,N_15330);
or U16313 (N_16313,N_15057,N_15520);
nand U16314 (N_16314,N_15210,N_15662);
and U16315 (N_16315,N_15405,N_15296);
or U16316 (N_16316,N_15430,N_15315);
nor U16317 (N_16317,N_15756,N_15267);
nor U16318 (N_16318,N_15066,N_15904);
nor U16319 (N_16319,N_15326,N_15998);
and U16320 (N_16320,N_15568,N_15259);
and U16321 (N_16321,N_15956,N_15067);
nor U16322 (N_16322,N_15323,N_15511);
xnor U16323 (N_16323,N_15947,N_15883);
and U16324 (N_16324,N_15053,N_15237);
and U16325 (N_16325,N_15428,N_15663);
or U16326 (N_16326,N_15449,N_15541);
nand U16327 (N_16327,N_15775,N_15623);
nor U16328 (N_16328,N_15731,N_15157);
or U16329 (N_16329,N_15812,N_15373);
nor U16330 (N_16330,N_15972,N_15216);
and U16331 (N_16331,N_15860,N_15787);
and U16332 (N_16332,N_15360,N_15983);
or U16333 (N_16333,N_15408,N_15228);
and U16334 (N_16334,N_15751,N_15090);
and U16335 (N_16335,N_15030,N_15525);
xor U16336 (N_16336,N_15152,N_15475);
or U16337 (N_16337,N_15031,N_15909);
or U16338 (N_16338,N_15220,N_15535);
nor U16339 (N_16339,N_15388,N_15923);
and U16340 (N_16340,N_15804,N_15837);
nand U16341 (N_16341,N_15960,N_15882);
or U16342 (N_16342,N_15279,N_15555);
or U16343 (N_16343,N_15831,N_15037);
nor U16344 (N_16344,N_15536,N_15892);
or U16345 (N_16345,N_15310,N_15419);
or U16346 (N_16346,N_15293,N_15467);
and U16347 (N_16347,N_15698,N_15607);
and U16348 (N_16348,N_15651,N_15329);
or U16349 (N_16349,N_15201,N_15040);
or U16350 (N_16350,N_15096,N_15807);
nor U16351 (N_16351,N_15515,N_15916);
nor U16352 (N_16352,N_15060,N_15463);
or U16353 (N_16353,N_15773,N_15391);
or U16354 (N_16354,N_15876,N_15264);
or U16355 (N_16355,N_15012,N_15017);
or U16356 (N_16356,N_15750,N_15445);
xnor U16357 (N_16357,N_15681,N_15432);
nor U16358 (N_16358,N_15487,N_15122);
nor U16359 (N_16359,N_15366,N_15581);
nand U16360 (N_16360,N_15796,N_15215);
nor U16361 (N_16361,N_15987,N_15585);
nand U16362 (N_16362,N_15013,N_15466);
nand U16363 (N_16363,N_15479,N_15908);
xor U16364 (N_16364,N_15819,N_15384);
and U16365 (N_16365,N_15671,N_15501);
xnor U16366 (N_16366,N_15113,N_15798);
xnor U16367 (N_16367,N_15941,N_15544);
nand U16368 (N_16368,N_15676,N_15872);
nand U16369 (N_16369,N_15092,N_15914);
nor U16370 (N_16370,N_15144,N_15209);
or U16371 (N_16371,N_15830,N_15669);
nand U16372 (N_16372,N_15106,N_15820);
nor U16373 (N_16373,N_15545,N_15291);
xor U16374 (N_16374,N_15980,N_15020);
or U16375 (N_16375,N_15285,N_15803);
or U16376 (N_16376,N_15431,N_15505);
nand U16377 (N_16377,N_15420,N_15447);
nor U16378 (N_16378,N_15976,N_15247);
and U16379 (N_16379,N_15494,N_15104);
nand U16380 (N_16380,N_15073,N_15593);
or U16381 (N_16381,N_15187,N_15429);
nand U16382 (N_16382,N_15167,N_15087);
and U16383 (N_16383,N_15572,N_15354);
and U16384 (N_16384,N_15644,N_15381);
xor U16385 (N_16385,N_15071,N_15016);
xnor U16386 (N_16386,N_15021,N_15734);
or U16387 (N_16387,N_15824,N_15622);
nand U16388 (N_16388,N_15863,N_15334);
and U16389 (N_16389,N_15802,N_15591);
or U16390 (N_16390,N_15508,N_15374);
or U16391 (N_16391,N_15199,N_15822);
or U16392 (N_16392,N_15885,N_15770);
nor U16393 (N_16393,N_15049,N_15203);
nand U16394 (N_16394,N_15621,N_15999);
nor U16395 (N_16395,N_15328,N_15879);
or U16396 (N_16396,N_15235,N_15504);
and U16397 (N_16397,N_15843,N_15887);
nand U16398 (N_16398,N_15086,N_15456);
nor U16399 (N_16399,N_15692,N_15918);
nand U16400 (N_16400,N_15055,N_15306);
nor U16401 (N_16401,N_15768,N_15540);
nor U16402 (N_16402,N_15742,N_15741);
nor U16403 (N_16403,N_15886,N_15236);
nor U16404 (N_16404,N_15559,N_15842);
nor U16405 (N_16405,N_15063,N_15045);
nor U16406 (N_16406,N_15849,N_15563);
nor U16407 (N_16407,N_15352,N_15425);
xor U16408 (N_16408,N_15338,N_15262);
nor U16409 (N_16409,N_15760,N_15179);
nor U16410 (N_16410,N_15966,N_15888);
or U16411 (N_16411,N_15478,N_15577);
xor U16412 (N_16412,N_15617,N_15243);
nor U16413 (N_16413,N_15418,N_15208);
xor U16414 (N_16414,N_15364,N_15407);
nor U16415 (N_16415,N_15783,N_15828);
or U16416 (N_16416,N_15727,N_15245);
nand U16417 (N_16417,N_15014,N_15724);
nor U16418 (N_16418,N_15349,N_15939);
nand U16419 (N_16419,N_15848,N_15376);
or U16420 (N_16420,N_15335,N_15471);
nand U16421 (N_16421,N_15763,N_15625);
nand U16422 (N_16422,N_15788,N_15588);
or U16423 (N_16423,N_15557,N_15229);
nand U16424 (N_16424,N_15638,N_15465);
xnor U16425 (N_16425,N_15641,N_15654);
nor U16426 (N_16426,N_15800,N_15776);
and U16427 (N_16427,N_15706,N_15552);
or U16428 (N_16428,N_15853,N_15301);
or U16429 (N_16429,N_15840,N_15937);
xnor U16430 (N_16430,N_15436,N_15813);
or U16431 (N_16431,N_15035,N_15415);
nand U16432 (N_16432,N_15250,N_15311);
xnor U16433 (N_16433,N_15903,N_15182);
and U16434 (N_16434,N_15862,N_15502);
nand U16435 (N_16435,N_15805,N_15304);
nor U16436 (N_16436,N_15845,N_15570);
nand U16437 (N_16437,N_15737,N_15119);
and U16438 (N_16438,N_15346,N_15485);
nor U16439 (N_16439,N_15403,N_15534);
xor U16440 (N_16440,N_15748,N_15410);
and U16441 (N_16441,N_15211,N_15472);
nor U16442 (N_16442,N_15533,N_15368);
nor U16443 (N_16443,N_15495,N_15924);
nor U16444 (N_16444,N_15480,N_15363);
nand U16445 (N_16445,N_15147,N_15386);
or U16446 (N_16446,N_15689,N_15797);
nor U16447 (N_16447,N_15613,N_15394);
or U16448 (N_16448,N_15967,N_15761);
or U16449 (N_16449,N_15524,N_15645);
and U16450 (N_16450,N_15114,N_15749);
or U16451 (N_16451,N_15602,N_15186);
and U16452 (N_16452,N_15153,N_15509);
nor U16453 (N_16453,N_15766,N_15855);
nand U16454 (N_16454,N_15130,N_15771);
and U16455 (N_16455,N_15006,N_15217);
nor U16456 (N_16456,N_15249,N_15109);
nor U16457 (N_16457,N_15531,N_15154);
nor U16458 (N_16458,N_15919,N_15189);
nor U16459 (N_16459,N_15680,N_15743);
or U16460 (N_16460,N_15988,N_15001);
and U16461 (N_16461,N_15599,N_15994);
nor U16462 (N_16462,N_15440,N_15514);
nor U16463 (N_16463,N_15393,N_15542);
xor U16464 (N_16464,N_15810,N_15180);
xor U16465 (N_16465,N_15424,N_15318);
xnor U16466 (N_16466,N_15990,N_15858);
nand U16467 (N_16467,N_15414,N_15164);
or U16468 (N_16468,N_15058,N_15562);
and U16469 (N_16469,N_15869,N_15174);
xor U16470 (N_16470,N_15401,N_15470);
and U16471 (N_16471,N_15367,N_15938);
and U16472 (N_16472,N_15458,N_15295);
nand U16473 (N_16473,N_15022,N_15818);
nor U16474 (N_16474,N_15920,N_15790);
or U16475 (N_16475,N_15913,N_15507);
nor U16476 (N_16476,N_15968,N_15708);
nor U16477 (N_16477,N_15263,N_15945);
and U16478 (N_16478,N_15646,N_15193);
or U16479 (N_16479,N_15816,N_15380);
nand U16480 (N_16480,N_15482,N_15392);
nor U16481 (N_16481,N_15932,N_15434);
or U16482 (N_16482,N_15218,N_15268);
xnor U16483 (N_16483,N_15497,N_15260);
and U16484 (N_16484,N_15580,N_15889);
xor U16485 (N_16485,N_15697,N_15448);
or U16486 (N_16486,N_15341,N_15567);
or U16487 (N_16487,N_15573,N_15225);
nor U16488 (N_16488,N_15569,N_15219);
nor U16489 (N_16489,N_15476,N_15290);
or U16490 (N_16490,N_15744,N_15442);
and U16491 (N_16491,N_15184,N_15801);
or U16492 (N_16492,N_15571,N_15331);
and U16493 (N_16493,N_15605,N_15592);
nand U16494 (N_16494,N_15409,N_15089);
nor U16495 (N_16495,N_15952,N_15548);
nand U16496 (N_16496,N_15111,N_15325);
and U16497 (N_16497,N_15183,N_15277);
nand U16498 (N_16498,N_15873,N_15716);
xor U16499 (N_16499,N_15492,N_15975);
or U16500 (N_16500,N_15631,N_15295);
nand U16501 (N_16501,N_15261,N_15031);
xnor U16502 (N_16502,N_15553,N_15368);
nand U16503 (N_16503,N_15192,N_15045);
or U16504 (N_16504,N_15019,N_15304);
or U16505 (N_16505,N_15382,N_15108);
nand U16506 (N_16506,N_15571,N_15752);
or U16507 (N_16507,N_15534,N_15011);
nand U16508 (N_16508,N_15659,N_15995);
nor U16509 (N_16509,N_15695,N_15999);
or U16510 (N_16510,N_15139,N_15730);
nand U16511 (N_16511,N_15394,N_15423);
xor U16512 (N_16512,N_15454,N_15021);
or U16513 (N_16513,N_15810,N_15588);
xnor U16514 (N_16514,N_15023,N_15241);
nor U16515 (N_16515,N_15684,N_15425);
xor U16516 (N_16516,N_15904,N_15385);
nor U16517 (N_16517,N_15521,N_15728);
nor U16518 (N_16518,N_15452,N_15641);
and U16519 (N_16519,N_15689,N_15158);
nand U16520 (N_16520,N_15802,N_15261);
or U16521 (N_16521,N_15687,N_15419);
nand U16522 (N_16522,N_15708,N_15021);
or U16523 (N_16523,N_15797,N_15508);
nor U16524 (N_16524,N_15752,N_15837);
nand U16525 (N_16525,N_15846,N_15252);
and U16526 (N_16526,N_15129,N_15630);
and U16527 (N_16527,N_15976,N_15736);
and U16528 (N_16528,N_15142,N_15149);
and U16529 (N_16529,N_15496,N_15121);
xnor U16530 (N_16530,N_15471,N_15764);
and U16531 (N_16531,N_15212,N_15337);
nor U16532 (N_16532,N_15804,N_15158);
and U16533 (N_16533,N_15975,N_15574);
and U16534 (N_16534,N_15477,N_15488);
or U16535 (N_16535,N_15940,N_15431);
or U16536 (N_16536,N_15031,N_15911);
or U16537 (N_16537,N_15203,N_15120);
xor U16538 (N_16538,N_15624,N_15434);
and U16539 (N_16539,N_15542,N_15341);
nand U16540 (N_16540,N_15496,N_15132);
nor U16541 (N_16541,N_15125,N_15077);
nand U16542 (N_16542,N_15898,N_15933);
or U16543 (N_16543,N_15266,N_15508);
and U16544 (N_16544,N_15384,N_15102);
nand U16545 (N_16545,N_15418,N_15580);
nand U16546 (N_16546,N_15880,N_15184);
xnor U16547 (N_16547,N_15119,N_15975);
xor U16548 (N_16548,N_15441,N_15628);
or U16549 (N_16549,N_15078,N_15569);
and U16550 (N_16550,N_15232,N_15885);
and U16551 (N_16551,N_15138,N_15298);
xor U16552 (N_16552,N_15931,N_15624);
and U16553 (N_16553,N_15239,N_15589);
xnor U16554 (N_16554,N_15909,N_15801);
nand U16555 (N_16555,N_15051,N_15334);
nand U16556 (N_16556,N_15700,N_15469);
nor U16557 (N_16557,N_15931,N_15868);
nand U16558 (N_16558,N_15054,N_15129);
xor U16559 (N_16559,N_15539,N_15638);
xor U16560 (N_16560,N_15701,N_15129);
nand U16561 (N_16561,N_15550,N_15734);
xnor U16562 (N_16562,N_15338,N_15460);
nand U16563 (N_16563,N_15545,N_15474);
xor U16564 (N_16564,N_15536,N_15094);
and U16565 (N_16565,N_15166,N_15838);
xor U16566 (N_16566,N_15256,N_15418);
xor U16567 (N_16567,N_15184,N_15964);
or U16568 (N_16568,N_15948,N_15134);
nand U16569 (N_16569,N_15903,N_15044);
nand U16570 (N_16570,N_15710,N_15581);
and U16571 (N_16571,N_15968,N_15041);
xnor U16572 (N_16572,N_15436,N_15050);
nor U16573 (N_16573,N_15182,N_15253);
nor U16574 (N_16574,N_15602,N_15352);
xor U16575 (N_16575,N_15744,N_15188);
and U16576 (N_16576,N_15253,N_15159);
and U16577 (N_16577,N_15335,N_15604);
xnor U16578 (N_16578,N_15258,N_15421);
and U16579 (N_16579,N_15475,N_15699);
nand U16580 (N_16580,N_15451,N_15788);
nor U16581 (N_16581,N_15092,N_15435);
or U16582 (N_16582,N_15952,N_15017);
nand U16583 (N_16583,N_15952,N_15465);
nand U16584 (N_16584,N_15822,N_15217);
nor U16585 (N_16585,N_15344,N_15962);
xnor U16586 (N_16586,N_15265,N_15890);
and U16587 (N_16587,N_15780,N_15161);
or U16588 (N_16588,N_15064,N_15881);
nor U16589 (N_16589,N_15394,N_15214);
nor U16590 (N_16590,N_15865,N_15236);
and U16591 (N_16591,N_15194,N_15642);
nand U16592 (N_16592,N_15709,N_15264);
xor U16593 (N_16593,N_15930,N_15827);
nor U16594 (N_16594,N_15990,N_15158);
nor U16595 (N_16595,N_15161,N_15098);
and U16596 (N_16596,N_15284,N_15741);
nand U16597 (N_16597,N_15653,N_15266);
or U16598 (N_16598,N_15285,N_15226);
or U16599 (N_16599,N_15073,N_15665);
or U16600 (N_16600,N_15662,N_15723);
xnor U16601 (N_16601,N_15210,N_15251);
nor U16602 (N_16602,N_15380,N_15747);
nand U16603 (N_16603,N_15927,N_15265);
and U16604 (N_16604,N_15324,N_15123);
nand U16605 (N_16605,N_15536,N_15476);
nand U16606 (N_16606,N_15649,N_15140);
or U16607 (N_16607,N_15815,N_15313);
xnor U16608 (N_16608,N_15246,N_15087);
nor U16609 (N_16609,N_15609,N_15237);
or U16610 (N_16610,N_15582,N_15674);
nand U16611 (N_16611,N_15310,N_15821);
and U16612 (N_16612,N_15927,N_15148);
xor U16613 (N_16613,N_15677,N_15862);
xor U16614 (N_16614,N_15974,N_15847);
or U16615 (N_16615,N_15427,N_15200);
nand U16616 (N_16616,N_15267,N_15076);
and U16617 (N_16617,N_15487,N_15026);
nand U16618 (N_16618,N_15647,N_15781);
xnor U16619 (N_16619,N_15548,N_15822);
or U16620 (N_16620,N_15708,N_15518);
or U16621 (N_16621,N_15137,N_15787);
and U16622 (N_16622,N_15054,N_15059);
or U16623 (N_16623,N_15228,N_15828);
nor U16624 (N_16624,N_15703,N_15373);
xnor U16625 (N_16625,N_15798,N_15545);
nand U16626 (N_16626,N_15600,N_15172);
or U16627 (N_16627,N_15612,N_15361);
xor U16628 (N_16628,N_15162,N_15906);
or U16629 (N_16629,N_15821,N_15820);
xor U16630 (N_16630,N_15904,N_15782);
or U16631 (N_16631,N_15197,N_15394);
or U16632 (N_16632,N_15498,N_15955);
and U16633 (N_16633,N_15531,N_15984);
or U16634 (N_16634,N_15139,N_15527);
and U16635 (N_16635,N_15615,N_15754);
nand U16636 (N_16636,N_15902,N_15272);
xnor U16637 (N_16637,N_15827,N_15432);
nand U16638 (N_16638,N_15564,N_15841);
and U16639 (N_16639,N_15181,N_15608);
and U16640 (N_16640,N_15791,N_15644);
xnor U16641 (N_16641,N_15669,N_15450);
xor U16642 (N_16642,N_15386,N_15930);
and U16643 (N_16643,N_15124,N_15634);
nand U16644 (N_16644,N_15370,N_15764);
xor U16645 (N_16645,N_15724,N_15039);
nor U16646 (N_16646,N_15711,N_15956);
or U16647 (N_16647,N_15372,N_15862);
nor U16648 (N_16648,N_15465,N_15020);
or U16649 (N_16649,N_15614,N_15853);
or U16650 (N_16650,N_15595,N_15935);
or U16651 (N_16651,N_15075,N_15503);
or U16652 (N_16652,N_15316,N_15872);
and U16653 (N_16653,N_15199,N_15737);
and U16654 (N_16654,N_15608,N_15416);
and U16655 (N_16655,N_15495,N_15774);
nor U16656 (N_16656,N_15843,N_15587);
nand U16657 (N_16657,N_15931,N_15249);
nand U16658 (N_16658,N_15617,N_15655);
xor U16659 (N_16659,N_15428,N_15699);
xor U16660 (N_16660,N_15911,N_15855);
nor U16661 (N_16661,N_15339,N_15246);
nor U16662 (N_16662,N_15565,N_15880);
or U16663 (N_16663,N_15768,N_15737);
or U16664 (N_16664,N_15079,N_15617);
and U16665 (N_16665,N_15124,N_15340);
nand U16666 (N_16666,N_15521,N_15238);
or U16667 (N_16667,N_15255,N_15539);
nor U16668 (N_16668,N_15036,N_15410);
nand U16669 (N_16669,N_15565,N_15330);
nor U16670 (N_16670,N_15404,N_15924);
or U16671 (N_16671,N_15927,N_15413);
or U16672 (N_16672,N_15601,N_15299);
or U16673 (N_16673,N_15657,N_15917);
and U16674 (N_16674,N_15265,N_15144);
and U16675 (N_16675,N_15678,N_15556);
and U16676 (N_16676,N_15213,N_15691);
and U16677 (N_16677,N_15178,N_15168);
nand U16678 (N_16678,N_15831,N_15969);
or U16679 (N_16679,N_15041,N_15138);
or U16680 (N_16680,N_15352,N_15778);
and U16681 (N_16681,N_15050,N_15818);
and U16682 (N_16682,N_15804,N_15201);
xnor U16683 (N_16683,N_15261,N_15058);
and U16684 (N_16684,N_15265,N_15710);
nand U16685 (N_16685,N_15588,N_15171);
xnor U16686 (N_16686,N_15241,N_15153);
xnor U16687 (N_16687,N_15963,N_15681);
or U16688 (N_16688,N_15395,N_15638);
xor U16689 (N_16689,N_15454,N_15453);
xnor U16690 (N_16690,N_15868,N_15664);
and U16691 (N_16691,N_15213,N_15311);
or U16692 (N_16692,N_15157,N_15588);
xnor U16693 (N_16693,N_15622,N_15916);
xnor U16694 (N_16694,N_15111,N_15313);
nand U16695 (N_16695,N_15839,N_15067);
or U16696 (N_16696,N_15848,N_15904);
and U16697 (N_16697,N_15097,N_15366);
or U16698 (N_16698,N_15216,N_15834);
and U16699 (N_16699,N_15872,N_15473);
xnor U16700 (N_16700,N_15605,N_15366);
nand U16701 (N_16701,N_15189,N_15159);
nor U16702 (N_16702,N_15342,N_15148);
xor U16703 (N_16703,N_15545,N_15193);
nand U16704 (N_16704,N_15713,N_15958);
nor U16705 (N_16705,N_15268,N_15020);
and U16706 (N_16706,N_15956,N_15289);
and U16707 (N_16707,N_15392,N_15123);
or U16708 (N_16708,N_15139,N_15442);
nor U16709 (N_16709,N_15503,N_15100);
or U16710 (N_16710,N_15904,N_15095);
xnor U16711 (N_16711,N_15810,N_15103);
nand U16712 (N_16712,N_15194,N_15084);
and U16713 (N_16713,N_15107,N_15436);
or U16714 (N_16714,N_15545,N_15717);
xnor U16715 (N_16715,N_15268,N_15289);
xor U16716 (N_16716,N_15967,N_15745);
or U16717 (N_16717,N_15342,N_15771);
nand U16718 (N_16718,N_15629,N_15141);
nor U16719 (N_16719,N_15587,N_15416);
and U16720 (N_16720,N_15387,N_15855);
nand U16721 (N_16721,N_15103,N_15813);
nand U16722 (N_16722,N_15210,N_15250);
nand U16723 (N_16723,N_15380,N_15186);
xor U16724 (N_16724,N_15997,N_15129);
or U16725 (N_16725,N_15502,N_15198);
xnor U16726 (N_16726,N_15328,N_15792);
nor U16727 (N_16727,N_15663,N_15987);
xnor U16728 (N_16728,N_15011,N_15200);
and U16729 (N_16729,N_15933,N_15138);
xnor U16730 (N_16730,N_15762,N_15863);
and U16731 (N_16731,N_15555,N_15262);
nor U16732 (N_16732,N_15677,N_15393);
and U16733 (N_16733,N_15740,N_15100);
xor U16734 (N_16734,N_15216,N_15801);
and U16735 (N_16735,N_15826,N_15671);
nand U16736 (N_16736,N_15313,N_15711);
and U16737 (N_16737,N_15641,N_15760);
or U16738 (N_16738,N_15068,N_15242);
nor U16739 (N_16739,N_15753,N_15087);
nor U16740 (N_16740,N_15948,N_15083);
xor U16741 (N_16741,N_15256,N_15839);
nand U16742 (N_16742,N_15462,N_15999);
nor U16743 (N_16743,N_15284,N_15710);
or U16744 (N_16744,N_15539,N_15456);
or U16745 (N_16745,N_15224,N_15297);
nand U16746 (N_16746,N_15798,N_15915);
nor U16747 (N_16747,N_15498,N_15459);
or U16748 (N_16748,N_15148,N_15969);
and U16749 (N_16749,N_15129,N_15797);
xor U16750 (N_16750,N_15758,N_15681);
xnor U16751 (N_16751,N_15446,N_15257);
xor U16752 (N_16752,N_15531,N_15936);
nor U16753 (N_16753,N_15759,N_15702);
nand U16754 (N_16754,N_15505,N_15675);
and U16755 (N_16755,N_15888,N_15481);
xor U16756 (N_16756,N_15794,N_15169);
and U16757 (N_16757,N_15786,N_15038);
nand U16758 (N_16758,N_15560,N_15758);
and U16759 (N_16759,N_15008,N_15339);
nand U16760 (N_16760,N_15559,N_15033);
nor U16761 (N_16761,N_15063,N_15524);
or U16762 (N_16762,N_15041,N_15247);
xor U16763 (N_16763,N_15027,N_15110);
and U16764 (N_16764,N_15297,N_15269);
xnor U16765 (N_16765,N_15345,N_15744);
or U16766 (N_16766,N_15392,N_15917);
or U16767 (N_16767,N_15422,N_15663);
nand U16768 (N_16768,N_15074,N_15186);
nor U16769 (N_16769,N_15163,N_15327);
and U16770 (N_16770,N_15248,N_15309);
nand U16771 (N_16771,N_15442,N_15065);
and U16772 (N_16772,N_15858,N_15944);
or U16773 (N_16773,N_15671,N_15348);
nor U16774 (N_16774,N_15589,N_15965);
nand U16775 (N_16775,N_15336,N_15110);
and U16776 (N_16776,N_15310,N_15858);
or U16777 (N_16777,N_15076,N_15646);
and U16778 (N_16778,N_15246,N_15337);
nor U16779 (N_16779,N_15531,N_15512);
nor U16780 (N_16780,N_15700,N_15883);
or U16781 (N_16781,N_15067,N_15240);
nor U16782 (N_16782,N_15690,N_15914);
nand U16783 (N_16783,N_15952,N_15904);
nand U16784 (N_16784,N_15896,N_15835);
or U16785 (N_16785,N_15214,N_15727);
and U16786 (N_16786,N_15340,N_15518);
nand U16787 (N_16787,N_15928,N_15885);
and U16788 (N_16788,N_15255,N_15494);
or U16789 (N_16789,N_15696,N_15299);
nor U16790 (N_16790,N_15252,N_15445);
and U16791 (N_16791,N_15569,N_15053);
and U16792 (N_16792,N_15709,N_15431);
nand U16793 (N_16793,N_15316,N_15794);
or U16794 (N_16794,N_15670,N_15530);
or U16795 (N_16795,N_15960,N_15300);
nand U16796 (N_16796,N_15598,N_15306);
or U16797 (N_16797,N_15836,N_15155);
nor U16798 (N_16798,N_15534,N_15359);
xor U16799 (N_16799,N_15127,N_15628);
nand U16800 (N_16800,N_15758,N_15261);
or U16801 (N_16801,N_15351,N_15841);
and U16802 (N_16802,N_15262,N_15615);
nor U16803 (N_16803,N_15225,N_15269);
and U16804 (N_16804,N_15726,N_15282);
nand U16805 (N_16805,N_15946,N_15091);
xor U16806 (N_16806,N_15220,N_15782);
xnor U16807 (N_16807,N_15493,N_15109);
xnor U16808 (N_16808,N_15102,N_15122);
nor U16809 (N_16809,N_15233,N_15770);
or U16810 (N_16810,N_15870,N_15965);
xor U16811 (N_16811,N_15220,N_15368);
xnor U16812 (N_16812,N_15995,N_15967);
nand U16813 (N_16813,N_15398,N_15259);
xnor U16814 (N_16814,N_15810,N_15225);
xnor U16815 (N_16815,N_15924,N_15089);
and U16816 (N_16816,N_15012,N_15392);
or U16817 (N_16817,N_15895,N_15839);
xnor U16818 (N_16818,N_15621,N_15026);
or U16819 (N_16819,N_15642,N_15529);
and U16820 (N_16820,N_15116,N_15780);
xor U16821 (N_16821,N_15640,N_15242);
and U16822 (N_16822,N_15485,N_15291);
xor U16823 (N_16823,N_15894,N_15804);
nor U16824 (N_16824,N_15272,N_15656);
nand U16825 (N_16825,N_15836,N_15216);
xor U16826 (N_16826,N_15750,N_15325);
nor U16827 (N_16827,N_15415,N_15006);
nor U16828 (N_16828,N_15786,N_15716);
nand U16829 (N_16829,N_15082,N_15173);
xor U16830 (N_16830,N_15625,N_15274);
and U16831 (N_16831,N_15458,N_15140);
and U16832 (N_16832,N_15250,N_15074);
and U16833 (N_16833,N_15451,N_15753);
or U16834 (N_16834,N_15238,N_15664);
nor U16835 (N_16835,N_15205,N_15600);
xor U16836 (N_16836,N_15750,N_15536);
nor U16837 (N_16837,N_15067,N_15147);
and U16838 (N_16838,N_15262,N_15370);
nor U16839 (N_16839,N_15421,N_15432);
nand U16840 (N_16840,N_15691,N_15546);
xnor U16841 (N_16841,N_15288,N_15507);
nand U16842 (N_16842,N_15219,N_15141);
nor U16843 (N_16843,N_15267,N_15030);
xnor U16844 (N_16844,N_15103,N_15556);
and U16845 (N_16845,N_15028,N_15914);
or U16846 (N_16846,N_15770,N_15836);
nand U16847 (N_16847,N_15511,N_15844);
and U16848 (N_16848,N_15853,N_15670);
or U16849 (N_16849,N_15605,N_15269);
nand U16850 (N_16850,N_15898,N_15090);
nand U16851 (N_16851,N_15612,N_15055);
xnor U16852 (N_16852,N_15057,N_15525);
xor U16853 (N_16853,N_15151,N_15771);
or U16854 (N_16854,N_15160,N_15294);
nand U16855 (N_16855,N_15089,N_15622);
nor U16856 (N_16856,N_15297,N_15074);
and U16857 (N_16857,N_15138,N_15277);
nand U16858 (N_16858,N_15127,N_15472);
and U16859 (N_16859,N_15607,N_15797);
xor U16860 (N_16860,N_15900,N_15603);
nand U16861 (N_16861,N_15513,N_15395);
nand U16862 (N_16862,N_15374,N_15531);
and U16863 (N_16863,N_15712,N_15470);
and U16864 (N_16864,N_15029,N_15844);
and U16865 (N_16865,N_15621,N_15446);
or U16866 (N_16866,N_15541,N_15125);
or U16867 (N_16867,N_15385,N_15838);
nand U16868 (N_16868,N_15182,N_15012);
nand U16869 (N_16869,N_15979,N_15592);
or U16870 (N_16870,N_15367,N_15314);
xor U16871 (N_16871,N_15805,N_15422);
xnor U16872 (N_16872,N_15117,N_15334);
nor U16873 (N_16873,N_15209,N_15682);
or U16874 (N_16874,N_15770,N_15054);
or U16875 (N_16875,N_15177,N_15572);
and U16876 (N_16876,N_15930,N_15244);
or U16877 (N_16877,N_15113,N_15602);
or U16878 (N_16878,N_15693,N_15057);
nand U16879 (N_16879,N_15640,N_15591);
nor U16880 (N_16880,N_15316,N_15777);
xor U16881 (N_16881,N_15143,N_15828);
nand U16882 (N_16882,N_15403,N_15552);
and U16883 (N_16883,N_15165,N_15858);
nand U16884 (N_16884,N_15871,N_15419);
nor U16885 (N_16885,N_15297,N_15260);
and U16886 (N_16886,N_15539,N_15838);
or U16887 (N_16887,N_15281,N_15050);
nand U16888 (N_16888,N_15042,N_15492);
nand U16889 (N_16889,N_15871,N_15797);
nand U16890 (N_16890,N_15566,N_15297);
nor U16891 (N_16891,N_15908,N_15415);
and U16892 (N_16892,N_15122,N_15289);
nand U16893 (N_16893,N_15476,N_15640);
nor U16894 (N_16894,N_15336,N_15069);
or U16895 (N_16895,N_15850,N_15387);
and U16896 (N_16896,N_15876,N_15514);
or U16897 (N_16897,N_15458,N_15451);
xor U16898 (N_16898,N_15297,N_15992);
nand U16899 (N_16899,N_15738,N_15801);
and U16900 (N_16900,N_15415,N_15463);
nand U16901 (N_16901,N_15832,N_15801);
and U16902 (N_16902,N_15831,N_15087);
and U16903 (N_16903,N_15189,N_15597);
and U16904 (N_16904,N_15797,N_15622);
or U16905 (N_16905,N_15759,N_15580);
xor U16906 (N_16906,N_15034,N_15884);
or U16907 (N_16907,N_15817,N_15791);
and U16908 (N_16908,N_15924,N_15663);
nor U16909 (N_16909,N_15128,N_15141);
nor U16910 (N_16910,N_15680,N_15790);
or U16911 (N_16911,N_15664,N_15601);
xnor U16912 (N_16912,N_15206,N_15065);
nor U16913 (N_16913,N_15280,N_15645);
or U16914 (N_16914,N_15646,N_15430);
or U16915 (N_16915,N_15988,N_15718);
nand U16916 (N_16916,N_15132,N_15921);
and U16917 (N_16917,N_15816,N_15844);
xnor U16918 (N_16918,N_15468,N_15298);
nand U16919 (N_16919,N_15113,N_15239);
xor U16920 (N_16920,N_15337,N_15851);
and U16921 (N_16921,N_15915,N_15515);
or U16922 (N_16922,N_15294,N_15076);
and U16923 (N_16923,N_15150,N_15006);
or U16924 (N_16924,N_15743,N_15247);
and U16925 (N_16925,N_15414,N_15606);
nor U16926 (N_16926,N_15244,N_15103);
nand U16927 (N_16927,N_15799,N_15307);
nor U16928 (N_16928,N_15384,N_15675);
xnor U16929 (N_16929,N_15645,N_15582);
or U16930 (N_16930,N_15213,N_15727);
nand U16931 (N_16931,N_15556,N_15390);
nor U16932 (N_16932,N_15204,N_15900);
nor U16933 (N_16933,N_15803,N_15479);
nand U16934 (N_16934,N_15127,N_15680);
and U16935 (N_16935,N_15686,N_15784);
nor U16936 (N_16936,N_15785,N_15032);
nand U16937 (N_16937,N_15489,N_15312);
nor U16938 (N_16938,N_15746,N_15107);
xnor U16939 (N_16939,N_15453,N_15868);
nand U16940 (N_16940,N_15415,N_15876);
nand U16941 (N_16941,N_15637,N_15132);
xnor U16942 (N_16942,N_15039,N_15255);
or U16943 (N_16943,N_15259,N_15721);
or U16944 (N_16944,N_15894,N_15072);
and U16945 (N_16945,N_15775,N_15598);
nor U16946 (N_16946,N_15592,N_15328);
and U16947 (N_16947,N_15381,N_15682);
nor U16948 (N_16948,N_15548,N_15978);
and U16949 (N_16949,N_15983,N_15111);
xor U16950 (N_16950,N_15463,N_15724);
and U16951 (N_16951,N_15113,N_15127);
and U16952 (N_16952,N_15368,N_15577);
or U16953 (N_16953,N_15448,N_15462);
xor U16954 (N_16954,N_15327,N_15981);
nor U16955 (N_16955,N_15564,N_15962);
xor U16956 (N_16956,N_15421,N_15521);
or U16957 (N_16957,N_15474,N_15320);
nand U16958 (N_16958,N_15670,N_15832);
or U16959 (N_16959,N_15145,N_15954);
or U16960 (N_16960,N_15601,N_15822);
nand U16961 (N_16961,N_15192,N_15052);
or U16962 (N_16962,N_15415,N_15369);
nor U16963 (N_16963,N_15755,N_15146);
and U16964 (N_16964,N_15222,N_15733);
xnor U16965 (N_16965,N_15075,N_15562);
or U16966 (N_16966,N_15473,N_15098);
or U16967 (N_16967,N_15904,N_15976);
or U16968 (N_16968,N_15990,N_15317);
or U16969 (N_16969,N_15232,N_15344);
nor U16970 (N_16970,N_15832,N_15308);
nor U16971 (N_16971,N_15093,N_15177);
xnor U16972 (N_16972,N_15462,N_15605);
nor U16973 (N_16973,N_15092,N_15289);
nor U16974 (N_16974,N_15598,N_15206);
and U16975 (N_16975,N_15679,N_15557);
and U16976 (N_16976,N_15433,N_15487);
or U16977 (N_16977,N_15981,N_15415);
nor U16978 (N_16978,N_15163,N_15161);
nor U16979 (N_16979,N_15574,N_15268);
nor U16980 (N_16980,N_15912,N_15578);
and U16981 (N_16981,N_15992,N_15931);
and U16982 (N_16982,N_15429,N_15922);
xnor U16983 (N_16983,N_15001,N_15800);
nor U16984 (N_16984,N_15921,N_15565);
nand U16985 (N_16985,N_15297,N_15185);
nor U16986 (N_16986,N_15996,N_15643);
or U16987 (N_16987,N_15133,N_15861);
xnor U16988 (N_16988,N_15543,N_15718);
or U16989 (N_16989,N_15236,N_15911);
nor U16990 (N_16990,N_15898,N_15089);
or U16991 (N_16991,N_15575,N_15610);
and U16992 (N_16992,N_15052,N_15368);
nand U16993 (N_16993,N_15619,N_15847);
nor U16994 (N_16994,N_15908,N_15937);
nand U16995 (N_16995,N_15239,N_15810);
nand U16996 (N_16996,N_15729,N_15239);
nand U16997 (N_16997,N_15736,N_15233);
and U16998 (N_16998,N_15202,N_15998);
nor U16999 (N_16999,N_15240,N_15477);
or U17000 (N_17000,N_16614,N_16912);
xor U17001 (N_17001,N_16256,N_16768);
nor U17002 (N_17002,N_16241,N_16441);
or U17003 (N_17003,N_16771,N_16871);
nand U17004 (N_17004,N_16608,N_16917);
nand U17005 (N_17005,N_16916,N_16514);
and U17006 (N_17006,N_16158,N_16326);
or U17007 (N_17007,N_16252,N_16755);
or U17008 (N_17008,N_16536,N_16601);
xnor U17009 (N_17009,N_16644,N_16167);
and U17010 (N_17010,N_16957,N_16224);
or U17011 (N_17011,N_16913,N_16584);
nand U17012 (N_17012,N_16604,N_16000);
or U17013 (N_17013,N_16367,N_16937);
and U17014 (N_17014,N_16515,N_16715);
nand U17015 (N_17015,N_16890,N_16829);
xnor U17016 (N_17016,N_16418,N_16749);
nand U17017 (N_17017,N_16783,N_16814);
nand U17018 (N_17018,N_16782,N_16131);
nand U17019 (N_17019,N_16493,N_16468);
or U17020 (N_17020,N_16853,N_16691);
nand U17021 (N_17021,N_16348,N_16803);
xnor U17022 (N_17022,N_16033,N_16234);
xor U17023 (N_17023,N_16636,N_16409);
nor U17024 (N_17024,N_16732,N_16927);
xor U17025 (N_17025,N_16322,N_16383);
xnor U17026 (N_17026,N_16382,N_16618);
nand U17027 (N_17027,N_16526,N_16754);
nor U17028 (N_17028,N_16545,N_16574);
xnor U17029 (N_17029,N_16101,N_16753);
and U17030 (N_17030,N_16053,N_16953);
and U17031 (N_17031,N_16959,N_16040);
or U17032 (N_17032,N_16787,N_16855);
xor U17033 (N_17033,N_16496,N_16664);
or U17034 (N_17034,N_16825,N_16698);
nand U17035 (N_17035,N_16541,N_16200);
or U17036 (N_17036,N_16936,N_16943);
or U17037 (N_17037,N_16102,N_16136);
and U17038 (N_17038,N_16891,N_16794);
nor U17039 (N_17039,N_16354,N_16907);
xor U17040 (N_17040,N_16027,N_16481);
and U17041 (N_17041,N_16193,N_16672);
xnor U17042 (N_17042,N_16061,N_16060);
xnor U17043 (N_17043,N_16870,N_16284);
nor U17044 (N_17044,N_16307,N_16702);
xnor U17045 (N_17045,N_16214,N_16550);
and U17046 (N_17046,N_16900,N_16110);
or U17047 (N_17047,N_16824,N_16652);
nor U17048 (N_17048,N_16126,N_16840);
or U17049 (N_17049,N_16296,N_16483);
nor U17050 (N_17050,N_16763,N_16598);
or U17051 (N_17051,N_16565,N_16162);
nor U17052 (N_17052,N_16624,N_16924);
nand U17053 (N_17053,N_16248,N_16124);
nor U17054 (N_17054,N_16222,N_16740);
and U17055 (N_17055,N_16457,N_16654);
and U17056 (N_17056,N_16616,N_16105);
nor U17057 (N_17057,N_16625,N_16517);
or U17058 (N_17058,N_16497,N_16716);
nand U17059 (N_17059,N_16251,N_16549);
nor U17060 (N_17060,N_16236,N_16095);
or U17061 (N_17061,N_16002,N_16998);
xor U17062 (N_17062,N_16933,N_16298);
xor U17063 (N_17063,N_16120,N_16888);
xnor U17064 (N_17064,N_16589,N_16190);
nor U17065 (N_17065,N_16649,N_16400);
nor U17066 (N_17066,N_16100,N_16967);
and U17067 (N_17067,N_16952,N_16440);
nor U17068 (N_17068,N_16524,N_16731);
nor U17069 (N_17069,N_16257,N_16336);
nor U17070 (N_17070,N_16311,N_16678);
nand U17071 (N_17071,N_16417,N_16914);
nand U17072 (N_17072,N_16387,N_16262);
or U17073 (N_17073,N_16792,N_16280);
nor U17074 (N_17074,N_16779,N_16041);
or U17075 (N_17075,N_16909,N_16466);
xnor U17076 (N_17076,N_16991,N_16321);
xnor U17077 (N_17077,N_16218,N_16020);
and U17078 (N_17078,N_16264,N_16301);
or U17079 (N_17079,N_16302,N_16266);
nor U17080 (N_17080,N_16064,N_16974);
and U17081 (N_17081,N_16031,N_16923);
nor U17082 (N_17082,N_16271,N_16004);
or U17083 (N_17083,N_16699,N_16137);
xnor U17084 (N_17084,N_16981,N_16237);
nor U17085 (N_17085,N_16227,N_16361);
or U17086 (N_17086,N_16419,N_16588);
xnor U17087 (N_17087,N_16893,N_16259);
xnor U17088 (N_17088,N_16747,N_16945);
nand U17089 (N_17089,N_16168,N_16939);
xnor U17090 (N_17090,N_16908,N_16976);
nand U17091 (N_17091,N_16926,N_16411);
xnor U17092 (N_17092,N_16895,N_16355);
nor U17093 (N_17093,N_16529,N_16484);
nor U17094 (N_17094,N_16290,N_16820);
and U17095 (N_17095,N_16425,N_16746);
or U17096 (N_17096,N_16019,N_16370);
nand U17097 (N_17097,N_16671,N_16198);
nor U17098 (N_17098,N_16465,N_16500);
and U17099 (N_17099,N_16947,N_16767);
and U17100 (N_17100,N_16076,N_16539);
or U17101 (N_17101,N_16569,N_16351);
or U17102 (N_17102,N_16899,N_16603);
nor U17103 (N_17103,N_16685,N_16179);
nand U17104 (N_17104,N_16217,N_16429);
nand U17105 (N_17105,N_16182,N_16445);
and U17106 (N_17106,N_16297,N_16192);
nand U17107 (N_17107,N_16204,N_16244);
xnor U17108 (N_17108,N_16170,N_16918);
or U17109 (N_17109,N_16003,N_16071);
and U17110 (N_17110,N_16159,N_16795);
and U17111 (N_17111,N_16316,N_16450);
and U17112 (N_17112,N_16130,N_16532);
nor U17113 (N_17113,N_16174,N_16530);
and U17114 (N_17114,N_16254,N_16555);
nand U17115 (N_17115,N_16379,N_16365);
xnor U17116 (N_17116,N_16531,N_16950);
nand U17117 (N_17117,N_16373,N_16276);
xnor U17118 (N_17118,N_16621,N_16760);
or U17119 (N_17119,N_16701,N_16811);
nor U17120 (N_17120,N_16097,N_16310);
xnor U17121 (N_17121,N_16312,N_16403);
nor U17122 (N_17122,N_16566,N_16941);
nor U17123 (N_17123,N_16665,N_16866);
xnor U17124 (N_17124,N_16593,N_16223);
and U17125 (N_17125,N_16576,N_16881);
xnor U17126 (N_17126,N_16764,N_16960);
and U17127 (N_17127,N_16303,N_16163);
xor U17128 (N_17128,N_16045,N_16595);
and U17129 (N_17129,N_16051,N_16435);
nand U17130 (N_17130,N_16535,N_16859);
and U17131 (N_17131,N_16925,N_16885);
nand U17132 (N_17132,N_16491,N_16821);
and U17133 (N_17133,N_16727,N_16743);
nor U17134 (N_17134,N_16988,N_16930);
and U17135 (N_17135,N_16381,N_16096);
nor U17136 (N_17136,N_16229,N_16323);
xor U17137 (N_17137,N_16453,N_16470);
or U17138 (N_17138,N_16836,N_16129);
nand U17139 (N_17139,N_16447,N_16340);
nand U17140 (N_17140,N_16639,N_16333);
nor U17141 (N_17141,N_16889,N_16971);
and U17142 (N_17142,N_16328,N_16875);
or U17143 (N_17143,N_16352,N_16730);
and U17144 (N_17144,N_16837,N_16751);
xnor U17145 (N_17145,N_16293,N_16294);
xnor U17146 (N_17146,N_16001,N_16809);
nand U17147 (N_17147,N_16852,N_16299);
nand U17148 (N_17148,N_16830,N_16581);
and U17149 (N_17149,N_16958,N_16434);
nand U17150 (N_17150,N_16479,N_16669);
nand U17151 (N_17151,N_16540,N_16023);
nand U17152 (N_17152,N_16670,N_16050);
and U17153 (N_17153,N_16117,N_16187);
and U17154 (N_17154,N_16029,N_16970);
nor U17155 (N_17155,N_16145,N_16700);
xor U17156 (N_17156,N_16788,N_16686);
and U17157 (N_17157,N_16647,N_16066);
or U17158 (N_17158,N_16552,N_16818);
nand U17159 (N_17159,N_16178,N_16165);
nand U17160 (N_17160,N_16490,N_16842);
nand U17161 (N_17161,N_16592,N_16068);
nand U17162 (N_17162,N_16920,N_16277);
xnor U17163 (N_17163,N_16774,N_16544);
or U17164 (N_17164,N_16494,N_16084);
xor U17165 (N_17165,N_16720,N_16006);
nor U17166 (N_17166,N_16646,N_16951);
nand U17167 (N_17167,N_16663,N_16523);
and U17168 (N_17168,N_16538,N_16346);
nor U17169 (N_17169,N_16590,N_16240);
and U17170 (N_17170,N_16693,N_16246);
or U17171 (N_17171,N_16688,N_16164);
and U17172 (N_17172,N_16074,N_16087);
nor U17173 (N_17173,N_16161,N_16209);
or U17174 (N_17174,N_16395,N_16780);
nand U17175 (N_17175,N_16273,N_16839);
and U17176 (N_17176,N_16123,N_16656);
nand U17177 (N_17177,N_16662,N_16687);
and U17178 (N_17178,N_16078,N_16106);
or U17179 (N_17179,N_16327,N_16047);
nand U17180 (N_17180,N_16350,N_16189);
or U17181 (N_17181,N_16210,N_16807);
or U17182 (N_17182,N_16609,N_16643);
nand U17183 (N_17183,N_16439,N_16808);
nand U17184 (N_17184,N_16784,N_16025);
nand U17185 (N_17185,N_16399,N_16832);
xor U17186 (N_17186,N_16680,N_16357);
xor U17187 (N_17187,N_16456,N_16631);
nor U17188 (N_17188,N_16378,N_16030);
nand U17189 (N_17189,N_16287,N_16330);
and U17190 (N_17190,N_16841,N_16342);
or U17191 (N_17191,N_16632,N_16949);
and U17192 (N_17192,N_16486,N_16557);
nor U17193 (N_17193,N_16738,N_16961);
xor U17194 (N_17194,N_16176,N_16079);
and U17195 (N_17195,N_16427,N_16542);
or U17196 (N_17196,N_16247,N_16083);
or U17197 (N_17197,N_16401,N_16903);
nor U17198 (N_17198,N_16709,N_16847);
nand U17199 (N_17199,N_16777,N_16673);
xnor U17200 (N_17200,N_16704,N_16519);
or U17201 (N_17201,N_16623,N_16243);
nor U17202 (N_17202,N_16010,N_16986);
or U17203 (N_17203,N_16172,N_16313);
and U17204 (N_17204,N_16320,N_16628);
nand U17205 (N_17205,N_16408,N_16442);
and U17206 (N_17206,N_16113,N_16392);
xor U17207 (N_17207,N_16469,N_16366);
and U17208 (N_17208,N_16461,N_16734);
xor U17209 (N_17209,N_16690,N_16140);
or U17210 (N_17210,N_16436,N_16577);
and U17211 (N_17211,N_16377,N_16478);
or U17212 (N_17212,N_16048,N_16773);
xor U17213 (N_17213,N_16054,N_16044);
nand U17214 (N_17214,N_16955,N_16769);
xor U17215 (N_17215,N_16547,N_16733);
and U17216 (N_17216,N_16127,N_16798);
or U17217 (N_17217,N_16558,N_16756);
or U17218 (N_17218,N_16444,N_16148);
or U17219 (N_17219,N_16509,N_16512);
nor U17220 (N_17220,N_16846,N_16992);
and U17221 (N_17221,N_16506,N_16677);
nand U17222 (N_17222,N_16719,N_16827);
or U17223 (N_17223,N_16089,N_16125);
or U17224 (N_17224,N_16093,N_16615);
xor U17225 (N_17225,N_16339,N_16188);
or U17226 (N_17226,N_16116,N_16527);
nor U17227 (N_17227,N_16085,N_16265);
nor U17228 (N_17228,N_16359,N_16586);
xnor U17229 (N_17229,N_16056,N_16850);
and U17230 (N_17230,N_16804,N_16281);
nor U17231 (N_17231,N_16356,N_16405);
nor U17232 (N_17232,N_16650,N_16398);
and U17233 (N_17233,N_16843,N_16729);
nor U17234 (N_17234,N_16848,N_16260);
and U17235 (N_17235,N_16407,N_16674);
and U17236 (N_17236,N_16906,N_16283);
nor U17237 (N_17237,N_16038,N_16215);
xnor U17238 (N_17238,N_16462,N_16208);
and U17239 (N_17239,N_16705,N_16965);
xor U17240 (N_17240,N_16122,N_16452);
and U17241 (N_17241,N_16666,N_16521);
nor U17242 (N_17242,N_16969,N_16424);
or U17243 (N_17243,N_16606,N_16714);
and U17244 (N_17244,N_16985,N_16343);
xor U17245 (N_17245,N_16617,N_16833);
nor U17246 (N_17246,N_16344,N_16869);
and U17247 (N_17247,N_16482,N_16360);
and U17248 (N_17248,N_16633,N_16799);
and U17249 (N_17249,N_16202,N_16009);
or U17250 (N_17250,N_16583,N_16725);
xnor U17251 (N_17251,N_16430,N_16384);
nand U17252 (N_17252,N_16416,N_16458);
xnor U17253 (N_17253,N_16088,N_16962);
nand U17254 (N_17254,N_16995,N_16393);
nor U17255 (N_17255,N_16718,N_16325);
nor U17256 (N_17256,N_16793,N_16203);
xnor U17257 (N_17257,N_16258,N_16362);
and U17258 (N_17258,N_16070,N_16928);
xnor U17259 (N_17259,N_16863,N_16683);
nand U17260 (N_17260,N_16472,N_16750);
nand U17261 (N_17261,N_16139,N_16942);
or U17262 (N_17262,N_16422,N_16684);
or U17263 (N_17263,N_16292,N_16641);
xnor U17264 (N_17264,N_16516,N_16910);
nand U17265 (N_17265,N_16249,N_16495);
nand U17266 (N_17266,N_16255,N_16706);
and U17267 (N_17267,N_16948,N_16619);
or U17268 (N_17268,N_16791,N_16114);
xnor U17269 (N_17269,N_16964,N_16790);
and U17270 (N_17270,N_16591,N_16011);
xor U17271 (N_17271,N_16039,N_16270);
xor U17272 (N_17272,N_16876,N_16554);
xnor U17273 (N_17273,N_16776,N_16502);
or U17274 (N_17274,N_16973,N_16402);
nor U17275 (N_17275,N_16710,N_16622);
and U17276 (N_17276,N_16533,N_16268);
nand U17277 (N_17277,N_16668,N_16508);
xor U17278 (N_17278,N_16872,N_16037);
and U17279 (N_17279,N_16826,N_16028);
and U17280 (N_17280,N_16874,N_16213);
nor U17281 (N_17281,N_16492,N_16388);
or U17282 (N_17282,N_16155,N_16058);
xnor U17283 (N_17283,N_16338,N_16815);
or U17284 (N_17284,N_16337,N_16786);
nor U17285 (N_17285,N_16012,N_16868);
nor U17286 (N_17286,N_16433,N_16475);
xnor U17287 (N_17287,N_16745,N_16956);
nor U17288 (N_17288,N_16655,N_16059);
and U17289 (N_17289,N_16762,N_16736);
nand U17290 (N_17290,N_16153,N_16865);
nor U17291 (N_17291,N_16696,N_16369);
and U17292 (N_17292,N_16658,N_16332);
or U17293 (N_17293,N_16175,N_16765);
xnor U17294 (N_17294,N_16504,N_16195);
and U17295 (N_17295,N_16659,N_16132);
and U17296 (N_17296,N_16713,N_16559);
nand U17297 (N_17297,N_16212,N_16349);
xnor U17298 (N_17298,N_16570,N_16073);
xnor U17299 (N_17299,N_16883,N_16897);
xnor U17300 (N_17300,N_16737,N_16488);
nand U17301 (N_17301,N_16568,N_16645);
xor U17302 (N_17302,N_16728,N_16415);
nor U17303 (N_17303,N_16315,N_16263);
and U17304 (N_17304,N_16564,N_16414);
or U17305 (N_17305,N_16744,N_16154);
or U17306 (N_17306,N_16186,N_16295);
xor U17307 (N_17307,N_16080,N_16477);
nor U17308 (N_17308,N_16977,N_16757);
nor U17309 (N_17309,N_16201,N_16703);
nand U17310 (N_17310,N_16391,N_16397);
or U17311 (N_17311,N_16109,N_16358);
nand U17312 (N_17312,N_16443,N_16055);
and U17313 (N_17313,N_16451,N_16235);
nand U17314 (N_17314,N_16230,N_16946);
xnor U17315 (N_17315,N_16726,N_16046);
or U17316 (N_17316,N_16640,N_16428);
or U17317 (N_17317,N_16341,N_16573);
nor U17318 (N_17318,N_16607,N_16057);
and U17319 (N_17319,N_16620,N_16390);
nand U17320 (N_17320,N_16752,N_16239);
nor U17321 (N_17321,N_16697,N_16485);
xnor U17322 (N_17322,N_16626,N_16594);
and U17323 (N_17323,N_16724,N_16579);
nor U17324 (N_17324,N_16982,N_16347);
nor U17325 (N_17325,N_16854,N_16021);
nor U17326 (N_17326,N_16972,N_16758);
and U17327 (N_17327,N_16413,N_16112);
or U17328 (N_17328,N_16610,N_16660);
or U17329 (N_17329,N_16968,N_16884);
or U17330 (N_17330,N_16371,N_16036);
nor U17331 (N_17331,N_16092,N_16835);
nor U17332 (N_17332,N_16963,N_16887);
or U17333 (N_17333,N_16169,N_16375);
nand U17334 (N_17334,N_16922,N_16374);
nor U17335 (N_17335,N_16759,N_16199);
nor U17336 (N_17336,N_16135,N_16845);
and U17337 (N_17337,N_16286,N_16134);
or U17338 (N_17338,N_16232,N_16994);
nand U17339 (N_17339,N_16785,N_16562);
nand U17340 (N_17340,N_16082,N_16886);
nor U17341 (N_17341,N_16308,N_16291);
or U17342 (N_17342,N_16880,N_16432);
or U17343 (N_17343,N_16858,N_16597);
nand U17344 (N_17344,N_16363,N_16548);
nand U17345 (N_17345,N_16676,N_16551);
xor U17346 (N_17346,N_16211,N_16525);
or U17347 (N_17347,N_16438,N_16386);
or U17348 (N_17348,N_16077,N_16142);
nand U17349 (N_17349,N_16449,N_16507);
nor U17350 (N_17350,N_16692,N_16708);
nand U17351 (N_17351,N_16675,N_16138);
nor U17352 (N_17352,N_16898,N_16410);
and U17353 (N_17353,N_16602,N_16471);
nor U17354 (N_17354,N_16630,N_16915);
or U17355 (N_17355,N_16599,N_16761);
nor U17356 (N_17356,N_16150,N_16860);
or U17357 (N_17357,N_16072,N_16722);
or U17358 (N_17358,N_16455,N_16838);
or U17359 (N_17359,N_16233,N_16999);
nand U17360 (N_17360,N_16274,N_16879);
and U17361 (N_17361,N_16166,N_16634);
nor U17362 (N_17362,N_16269,N_16935);
or U17363 (N_17363,N_16712,N_16099);
and U17364 (N_17364,N_16892,N_16086);
xor U17365 (N_17365,N_16775,N_16812);
xnor U17366 (N_17366,N_16667,N_16067);
and U17367 (N_17367,N_16331,N_16220);
and U17368 (N_17368,N_16062,N_16035);
or U17369 (N_17369,N_16103,N_16834);
or U17370 (N_17370,N_16335,N_16996);
xnor U17371 (N_17371,N_16796,N_16115);
or U17372 (N_17372,N_16934,N_16587);
nand U17373 (N_17373,N_16228,N_16772);
xor U17374 (N_17374,N_16707,N_16171);
nor U17375 (N_17375,N_16474,N_16987);
nor U17376 (N_17376,N_16431,N_16008);
nor U17377 (N_17377,N_16144,N_16278);
nor U17378 (N_17378,N_16467,N_16537);
and U17379 (N_17379,N_16627,N_16226);
nor U17380 (N_17380,N_16997,N_16238);
nor U17381 (N_17381,N_16575,N_16816);
and U17382 (N_17382,N_16689,N_16090);
nor U17383 (N_17383,N_16742,N_16141);
and U17384 (N_17384,N_16406,N_16463);
xnor U17385 (N_17385,N_16318,N_16454);
or U17386 (N_17386,N_16065,N_16196);
nor U17387 (N_17387,N_16931,N_16205);
xnor U17388 (N_17388,N_16648,N_16007);
and U17389 (N_17389,N_16851,N_16081);
xnor U17390 (N_17390,N_16543,N_16520);
and U17391 (N_17391,N_16563,N_16063);
and U17392 (N_17392,N_16111,N_16661);
nand U17393 (N_17393,N_16990,N_16878);
or U17394 (N_17394,N_16739,N_16143);
nand U17395 (N_17395,N_16993,N_16817);
and U17396 (N_17396,N_16919,N_16151);
nor U17397 (N_17397,N_16368,N_16806);
nor U17398 (N_17398,N_16789,N_16245);
nor U17399 (N_17399,N_16556,N_16197);
xnor U17400 (N_17400,N_16285,N_16194);
and U17401 (N_17401,N_16032,N_16075);
nor U17402 (N_17402,N_16364,N_16394);
or U17403 (N_17403,N_16306,N_16024);
and U17404 (N_17404,N_16324,N_16476);
nor U17405 (N_17405,N_16043,N_16282);
nor U17406 (N_17406,N_16844,N_16911);
xor U17407 (N_17407,N_16582,N_16412);
nand U17408 (N_17408,N_16721,N_16014);
nand U17409 (N_17409,N_16635,N_16108);
and U17410 (N_17410,N_16905,N_16423);
and U17411 (N_17411,N_16446,N_16638);
nor U17412 (N_17412,N_16857,N_16546);
nor U17413 (N_17413,N_16219,N_16448);
nand U17414 (N_17414,N_16978,N_16813);
nand U17415 (N_17415,N_16567,N_16156);
nor U17416 (N_17416,N_16651,N_16864);
nor U17417 (N_17417,N_16052,N_16018);
and U17418 (N_17418,N_16781,N_16420);
and U17419 (N_17419,N_16954,N_16221);
and U17420 (N_17420,N_16334,N_16637);
xor U17421 (N_17421,N_16894,N_16118);
nor U17422 (N_17422,N_16017,N_16612);
or U17423 (N_17423,N_16505,N_16572);
xor U17424 (N_17424,N_16944,N_16819);
nor U17425 (N_17425,N_16207,N_16571);
nand U17426 (N_17426,N_16437,N_16225);
and U17427 (N_17427,N_16250,N_16980);
nor U17428 (N_17428,N_16861,N_16133);
and U17429 (N_17429,N_16015,N_16578);
or U17430 (N_17430,N_16510,N_16938);
nand U17431 (N_17431,N_16989,N_16372);
or U17432 (N_17432,N_16711,N_16404);
and U17433 (N_17433,N_16717,N_16805);
and U17434 (N_17434,N_16319,N_16489);
xor U17435 (N_17435,N_16983,N_16766);
nor U17436 (N_17436,N_16191,N_16121);
nor U17437 (N_17437,N_16242,N_16042);
or U17438 (N_17438,N_16741,N_16146);
nor U17439 (N_17439,N_16682,N_16289);
and U17440 (N_17440,N_16314,N_16653);
xor U17441 (N_17441,N_16929,N_16498);
xor U17442 (N_17442,N_16511,N_16975);
nor U17443 (N_17443,N_16421,N_16480);
or U17444 (N_17444,N_16695,N_16152);
nand U17445 (N_17445,N_16694,N_16831);
xor U17446 (N_17446,N_16013,N_16580);
xor U17447 (N_17447,N_16157,N_16828);
nor U17448 (N_17448,N_16534,N_16091);
or U17449 (N_17449,N_16317,N_16288);
xor U17450 (N_17450,N_16501,N_16629);
or U17451 (N_17451,N_16005,N_16810);
nor U17452 (N_17452,N_16613,N_16770);
nand U17453 (N_17453,N_16098,N_16778);
or U17454 (N_17454,N_16657,N_16049);
nor U17455 (N_17455,N_16862,N_16503);
nand U17456 (N_17456,N_16173,N_16460);
or U17457 (N_17457,N_16518,N_16329);
or U17458 (N_17458,N_16932,N_16561);
xor U17459 (N_17459,N_16119,N_16600);
nor U17460 (N_17460,N_16797,N_16877);
and U17461 (N_17461,N_16309,N_16801);
nor U17462 (N_17462,N_16528,N_16679);
or U17463 (N_17463,N_16513,N_16016);
nor U17464 (N_17464,N_16380,N_16185);
or U17465 (N_17465,N_16735,N_16376);
or U17466 (N_17466,N_16823,N_16681);
or U17467 (N_17467,N_16305,N_16069);
and U17468 (N_17468,N_16585,N_16487);
nand U17469 (N_17469,N_16596,N_16940);
or U17470 (N_17470,N_16522,N_16553);
nor U17471 (N_17471,N_16800,N_16181);
nor U17472 (N_17472,N_16177,N_16896);
xnor U17473 (N_17473,N_16426,N_16183);
and U17474 (N_17474,N_16261,N_16499);
nand U17475 (N_17475,N_16748,N_16459);
or U17476 (N_17476,N_16231,N_16353);
or U17477 (N_17477,N_16034,N_16160);
nand U17478 (N_17478,N_16272,N_16802);
nand U17479 (N_17479,N_16304,N_16128);
or U17480 (N_17480,N_16022,N_16902);
nand U17481 (N_17481,N_16147,N_16873);
nor U17482 (N_17482,N_16275,N_16560);
nand U17483 (N_17483,N_16279,N_16822);
xor U17484 (N_17484,N_16253,N_16723);
and U17485 (N_17485,N_16267,N_16849);
nand U17486 (N_17486,N_16867,N_16180);
nor U17487 (N_17487,N_16216,N_16605);
nand U17488 (N_17488,N_16149,N_16389);
nand U17489 (N_17489,N_16026,N_16979);
nor U17490 (N_17490,N_16300,N_16904);
nand U17491 (N_17491,N_16921,N_16464);
xor U17492 (N_17492,N_16184,N_16611);
or U17493 (N_17493,N_16396,N_16856);
nand U17494 (N_17494,N_16206,N_16385);
and U17495 (N_17495,N_16966,N_16107);
and U17496 (N_17496,N_16984,N_16473);
and U17497 (N_17497,N_16642,N_16104);
nand U17498 (N_17498,N_16094,N_16901);
xor U17499 (N_17499,N_16345,N_16882);
nor U17500 (N_17500,N_16130,N_16627);
nor U17501 (N_17501,N_16203,N_16815);
xnor U17502 (N_17502,N_16767,N_16246);
and U17503 (N_17503,N_16013,N_16337);
or U17504 (N_17504,N_16865,N_16121);
xor U17505 (N_17505,N_16174,N_16092);
and U17506 (N_17506,N_16785,N_16619);
xnor U17507 (N_17507,N_16816,N_16114);
nor U17508 (N_17508,N_16021,N_16316);
or U17509 (N_17509,N_16573,N_16780);
nand U17510 (N_17510,N_16539,N_16260);
xor U17511 (N_17511,N_16821,N_16967);
and U17512 (N_17512,N_16340,N_16585);
nor U17513 (N_17513,N_16201,N_16812);
or U17514 (N_17514,N_16966,N_16901);
nor U17515 (N_17515,N_16283,N_16659);
nor U17516 (N_17516,N_16931,N_16075);
nor U17517 (N_17517,N_16593,N_16292);
nor U17518 (N_17518,N_16928,N_16199);
nor U17519 (N_17519,N_16420,N_16102);
nor U17520 (N_17520,N_16219,N_16942);
or U17521 (N_17521,N_16968,N_16406);
or U17522 (N_17522,N_16064,N_16340);
nor U17523 (N_17523,N_16075,N_16834);
nand U17524 (N_17524,N_16646,N_16201);
nand U17525 (N_17525,N_16775,N_16884);
nor U17526 (N_17526,N_16399,N_16913);
and U17527 (N_17527,N_16415,N_16045);
nor U17528 (N_17528,N_16956,N_16131);
nand U17529 (N_17529,N_16343,N_16976);
or U17530 (N_17530,N_16475,N_16270);
nor U17531 (N_17531,N_16989,N_16986);
or U17532 (N_17532,N_16856,N_16088);
or U17533 (N_17533,N_16693,N_16830);
nor U17534 (N_17534,N_16698,N_16900);
or U17535 (N_17535,N_16534,N_16895);
nor U17536 (N_17536,N_16112,N_16834);
nand U17537 (N_17537,N_16847,N_16076);
xnor U17538 (N_17538,N_16831,N_16405);
nand U17539 (N_17539,N_16352,N_16400);
nand U17540 (N_17540,N_16730,N_16236);
xnor U17541 (N_17541,N_16419,N_16306);
or U17542 (N_17542,N_16501,N_16108);
nand U17543 (N_17543,N_16932,N_16896);
xor U17544 (N_17544,N_16463,N_16013);
xnor U17545 (N_17545,N_16318,N_16613);
and U17546 (N_17546,N_16793,N_16121);
nand U17547 (N_17547,N_16472,N_16174);
xnor U17548 (N_17548,N_16088,N_16573);
nor U17549 (N_17549,N_16229,N_16232);
or U17550 (N_17550,N_16923,N_16233);
nand U17551 (N_17551,N_16301,N_16800);
or U17552 (N_17552,N_16456,N_16514);
or U17553 (N_17553,N_16292,N_16038);
xnor U17554 (N_17554,N_16782,N_16464);
and U17555 (N_17555,N_16384,N_16565);
or U17556 (N_17556,N_16199,N_16329);
xnor U17557 (N_17557,N_16833,N_16080);
nor U17558 (N_17558,N_16198,N_16508);
xnor U17559 (N_17559,N_16921,N_16724);
or U17560 (N_17560,N_16789,N_16682);
nor U17561 (N_17561,N_16317,N_16302);
or U17562 (N_17562,N_16744,N_16012);
nor U17563 (N_17563,N_16425,N_16643);
xor U17564 (N_17564,N_16642,N_16772);
or U17565 (N_17565,N_16033,N_16674);
nor U17566 (N_17566,N_16703,N_16256);
nand U17567 (N_17567,N_16572,N_16149);
or U17568 (N_17568,N_16826,N_16229);
and U17569 (N_17569,N_16855,N_16781);
xor U17570 (N_17570,N_16860,N_16086);
or U17571 (N_17571,N_16836,N_16432);
nand U17572 (N_17572,N_16809,N_16596);
nor U17573 (N_17573,N_16547,N_16621);
or U17574 (N_17574,N_16828,N_16517);
nand U17575 (N_17575,N_16322,N_16690);
nor U17576 (N_17576,N_16600,N_16488);
xnor U17577 (N_17577,N_16820,N_16519);
and U17578 (N_17578,N_16395,N_16235);
xor U17579 (N_17579,N_16231,N_16146);
nand U17580 (N_17580,N_16920,N_16043);
or U17581 (N_17581,N_16791,N_16695);
xnor U17582 (N_17582,N_16468,N_16787);
nor U17583 (N_17583,N_16465,N_16092);
xnor U17584 (N_17584,N_16075,N_16701);
nand U17585 (N_17585,N_16493,N_16646);
and U17586 (N_17586,N_16896,N_16921);
nand U17587 (N_17587,N_16024,N_16525);
and U17588 (N_17588,N_16213,N_16081);
xnor U17589 (N_17589,N_16681,N_16983);
or U17590 (N_17590,N_16856,N_16497);
and U17591 (N_17591,N_16497,N_16182);
nor U17592 (N_17592,N_16927,N_16514);
nor U17593 (N_17593,N_16935,N_16811);
or U17594 (N_17594,N_16483,N_16791);
or U17595 (N_17595,N_16306,N_16430);
nand U17596 (N_17596,N_16441,N_16233);
xor U17597 (N_17597,N_16406,N_16455);
nor U17598 (N_17598,N_16391,N_16105);
nor U17599 (N_17599,N_16574,N_16867);
nand U17600 (N_17600,N_16525,N_16808);
and U17601 (N_17601,N_16750,N_16792);
and U17602 (N_17602,N_16991,N_16162);
nor U17603 (N_17603,N_16318,N_16183);
nand U17604 (N_17604,N_16473,N_16718);
and U17605 (N_17605,N_16927,N_16873);
xnor U17606 (N_17606,N_16696,N_16773);
xnor U17607 (N_17607,N_16252,N_16573);
or U17608 (N_17608,N_16806,N_16491);
or U17609 (N_17609,N_16308,N_16591);
nand U17610 (N_17610,N_16182,N_16833);
nor U17611 (N_17611,N_16136,N_16956);
nand U17612 (N_17612,N_16602,N_16879);
nor U17613 (N_17613,N_16460,N_16198);
nor U17614 (N_17614,N_16331,N_16870);
and U17615 (N_17615,N_16254,N_16804);
nand U17616 (N_17616,N_16009,N_16749);
nor U17617 (N_17617,N_16099,N_16135);
nor U17618 (N_17618,N_16430,N_16414);
or U17619 (N_17619,N_16635,N_16557);
nor U17620 (N_17620,N_16328,N_16700);
nand U17621 (N_17621,N_16324,N_16339);
nand U17622 (N_17622,N_16395,N_16012);
xor U17623 (N_17623,N_16194,N_16638);
nand U17624 (N_17624,N_16792,N_16977);
nand U17625 (N_17625,N_16690,N_16460);
and U17626 (N_17626,N_16569,N_16871);
xor U17627 (N_17627,N_16189,N_16154);
nor U17628 (N_17628,N_16151,N_16969);
and U17629 (N_17629,N_16894,N_16257);
xnor U17630 (N_17630,N_16836,N_16843);
xor U17631 (N_17631,N_16732,N_16237);
or U17632 (N_17632,N_16158,N_16581);
nand U17633 (N_17633,N_16444,N_16554);
nor U17634 (N_17634,N_16090,N_16740);
nand U17635 (N_17635,N_16375,N_16916);
nand U17636 (N_17636,N_16841,N_16198);
nand U17637 (N_17637,N_16361,N_16143);
or U17638 (N_17638,N_16015,N_16254);
and U17639 (N_17639,N_16141,N_16579);
and U17640 (N_17640,N_16340,N_16391);
and U17641 (N_17641,N_16057,N_16107);
nor U17642 (N_17642,N_16292,N_16474);
nand U17643 (N_17643,N_16354,N_16149);
and U17644 (N_17644,N_16646,N_16596);
nor U17645 (N_17645,N_16762,N_16943);
and U17646 (N_17646,N_16304,N_16237);
xor U17647 (N_17647,N_16101,N_16920);
and U17648 (N_17648,N_16616,N_16360);
nand U17649 (N_17649,N_16545,N_16441);
nand U17650 (N_17650,N_16962,N_16307);
nor U17651 (N_17651,N_16206,N_16219);
nand U17652 (N_17652,N_16983,N_16764);
and U17653 (N_17653,N_16694,N_16019);
and U17654 (N_17654,N_16178,N_16399);
nand U17655 (N_17655,N_16607,N_16229);
xor U17656 (N_17656,N_16465,N_16991);
nor U17657 (N_17657,N_16518,N_16702);
or U17658 (N_17658,N_16980,N_16059);
nor U17659 (N_17659,N_16472,N_16688);
xor U17660 (N_17660,N_16009,N_16314);
nor U17661 (N_17661,N_16568,N_16786);
or U17662 (N_17662,N_16171,N_16321);
and U17663 (N_17663,N_16414,N_16041);
or U17664 (N_17664,N_16222,N_16737);
nand U17665 (N_17665,N_16075,N_16616);
nand U17666 (N_17666,N_16506,N_16860);
nand U17667 (N_17667,N_16983,N_16046);
nor U17668 (N_17668,N_16556,N_16050);
nor U17669 (N_17669,N_16554,N_16426);
nand U17670 (N_17670,N_16505,N_16234);
xor U17671 (N_17671,N_16145,N_16196);
nand U17672 (N_17672,N_16037,N_16544);
and U17673 (N_17673,N_16896,N_16616);
xor U17674 (N_17674,N_16518,N_16792);
nand U17675 (N_17675,N_16474,N_16434);
nand U17676 (N_17676,N_16824,N_16550);
nand U17677 (N_17677,N_16119,N_16969);
nand U17678 (N_17678,N_16069,N_16936);
nor U17679 (N_17679,N_16328,N_16924);
nand U17680 (N_17680,N_16795,N_16117);
and U17681 (N_17681,N_16939,N_16736);
or U17682 (N_17682,N_16529,N_16367);
xor U17683 (N_17683,N_16451,N_16317);
nand U17684 (N_17684,N_16768,N_16385);
nand U17685 (N_17685,N_16660,N_16000);
nand U17686 (N_17686,N_16209,N_16993);
nand U17687 (N_17687,N_16855,N_16779);
or U17688 (N_17688,N_16567,N_16735);
or U17689 (N_17689,N_16494,N_16726);
nor U17690 (N_17690,N_16560,N_16343);
or U17691 (N_17691,N_16080,N_16966);
nor U17692 (N_17692,N_16824,N_16789);
or U17693 (N_17693,N_16512,N_16901);
xor U17694 (N_17694,N_16777,N_16183);
nand U17695 (N_17695,N_16634,N_16290);
and U17696 (N_17696,N_16848,N_16010);
nand U17697 (N_17697,N_16095,N_16634);
nand U17698 (N_17698,N_16015,N_16150);
xor U17699 (N_17699,N_16382,N_16443);
nor U17700 (N_17700,N_16186,N_16885);
and U17701 (N_17701,N_16818,N_16257);
xor U17702 (N_17702,N_16560,N_16322);
xnor U17703 (N_17703,N_16595,N_16968);
nor U17704 (N_17704,N_16957,N_16351);
and U17705 (N_17705,N_16663,N_16021);
nand U17706 (N_17706,N_16925,N_16748);
nor U17707 (N_17707,N_16567,N_16063);
nor U17708 (N_17708,N_16010,N_16558);
xnor U17709 (N_17709,N_16819,N_16613);
and U17710 (N_17710,N_16485,N_16276);
or U17711 (N_17711,N_16777,N_16870);
xnor U17712 (N_17712,N_16765,N_16906);
nand U17713 (N_17713,N_16895,N_16563);
and U17714 (N_17714,N_16754,N_16710);
and U17715 (N_17715,N_16980,N_16684);
or U17716 (N_17716,N_16440,N_16986);
nand U17717 (N_17717,N_16023,N_16207);
or U17718 (N_17718,N_16223,N_16251);
or U17719 (N_17719,N_16426,N_16887);
or U17720 (N_17720,N_16364,N_16156);
nand U17721 (N_17721,N_16360,N_16096);
nor U17722 (N_17722,N_16714,N_16929);
nand U17723 (N_17723,N_16649,N_16802);
nor U17724 (N_17724,N_16518,N_16460);
and U17725 (N_17725,N_16630,N_16584);
xnor U17726 (N_17726,N_16747,N_16248);
or U17727 (N_17727,N_16719,N_16696);
nand U17728 (N_17728,N_16215,N_16081);
nor U17729 (N_17729,N_16572,N_16441);
and U17730 (N_17730,N_16885,N_16373);
and U17731 (N_17731,N_16055,N_16451);
nor U17732 (N_17732,N_16448,N_16013);
nand U17733 (N_17733,N_16041,N_16711);
nand U17734 (N_17734,N_16450,N_16248);
xnor U17735 (N_17735,N_16488,N_16847);
or U17736 (N_17736,N_16154,N_16074);
nand U17737 (N_17737,N_16052,N_16059);
and U17738 (N_17738,N_16116,N_16625);
or U17739 (N_17739,N_16394,N_16645);
nand U17740 (N_17740,N_16860,N_16603);
or U17741 (N_17741,N_16626,N_16811);
or U17742 (N_17742,N_16937,N_16880);
and U17743 (N_17743,N_16108,N_16517);
nand U17744 (N_17744,N_16473,N_16159);
and U17745 (N_17745,N_16393,N_16491);
nor U17746 (N_17746,N_16655,N_16323);
nand U17747 (N_17747,N_16119,N_16996);
or U17748 (N_17748,N_16218,N_16185);
xor U17749 (N_17749,N_16529,N_16293);
nand U17750 (N_17750,N_16310,N_16314);
and U17751 (N_17751,N_16967,N_16976);
nor U17752 (N_17752,N_16516,N_16271);
or U17753 (N_17753,N_16736,N_16774);
nand U17754 (N_17754,N_16767,N_16969);
and U17755 (N_17755,N_16490,N_16409);
xor U17756 (N_17756,N_16733,N_16794);
or U17757 (N_17757,N_16506,N_16901);
nand U17758 (N_17758,N_16128,N_16020);
and U17759 (N_17759,N_16143,N_16224);
nand U17760 (N_17760,N_16923,N_16063);
or U17761 (N_17761,N_16600,N_16113);
nand U17762 (N_17762,N_16153,N_16533);
and U17763 (N_17763,N_16378,N_16797);
nand U17764 (N_17764,N_16171,N_16081);
and U17765 (N_17765,N_16423,N_16585);
xor U17766 (N_17766,N_16256,N_16743);
nor U17767 (N_17767,N_16134,N_16438);
and U17768 (N_17768,N_16502,N_16751);
and U17769 (N_17769,N_16768,N_16839);
nor U17770 (N_17770,N_16952,N_16585);
xor U17771 (N_17771,N_16395,N_16677);
or U17772 (N_17772,N_16631,N_16062);
or U17773 (N_17773,N_16291,N_16490);
nand U17774 (N_17774,N_16352,N_16277);
nor U17775 (N_17775,N_16611,N_16681);
nor U17776 (N_17776,N_16924,N_16213);
nor U17777 (N_17777,N_16299,N_16005);
nor U17778 (N_17778,N_16812,N_16914);
xnor U17779 (N_17779,N_16549,N_16734);
xnor U17780 (N_17780,N_16913,N_16286);
or U17781 (N_17781,N_16570,N_16128);
nor U17782 (N_17782,N_16274,N_16104);
xor U17783 (N_17783,N_16490,N_16813);
nand U17784 (N_17784,N_16687,N_16578);
and U17785 (N_17785,N_16275,N_16979);
nand U17786 (N_17786,N_16714,N_16443);
nor U17787 (N_17787,N_16596,N_16935);
xor U17788 (N_17788,N_16321,N_16530);
xor U17789 (N_17789,N_16422,N_16276);
nand U17790 (N_17790,N_16806,N_16860);
nand U17791 (N_17791,N_16790,N_16267);
xor U17792 (N_17792,N_16333,N_16470);
or U17793 (N_17793,N_16651,N_16832);
xnor U17794 (N_17794,N_16074,N_16378);
or U17795 (N_17795,N_16388,N_16923);
xnor U17796 (N_17796,N_16240,N_16561);
nor U17797 (N_17797,N_16458,N_16564);
nand U17798 (N_17798,N_16543,N_16712);
or U17799 (N_17799,N_16408,N_16320);
nand U17800 (N_17800,N_16475,N_16259);
xor U17801 (N_17801,N_16243,N_16483);
nor U17802 (N_17802,N_16368,N_16198);
nor U17803 (N_17803,N_16054,N_16010);
or U17804 (N_17804,N_16689,N_16315);
or U17805 (N_17805,N_16725,N_16930);
nor U17806 (N_17806,N_16843,N_16299);
xor U17807 (N_17807,N_16142,N_16800);
xor U17808 (N_17808,N_16876,N_16117);
and U17809 (N_17809,N_16285,N_16704);
or U17810 (N_17810,N_16037,N_16296);
and U17811 (N_17811,N_16076,N_16180);
xor U17812 (N_17812,N_16719,N_16547);
xor U17813 (N_17813,N_16294,N_16616);
and U17814 (N_17814,N_16417,N_16352);
xor U17815 (N_17815,N_16072,N_16901);
nand U17816 (N_17816,N_16291,N_16607);
nor U17817 (N_17817,N_16303,N_16086);
xnor U17818 (N_17818,N_16476,N_16070);
nor U17819 (N_17819,N_16647,N_16432);
and U17820 (N_17820,N_16040,N_16558);
xnor U17821 (N_17821,N_16408,N_16838);
nor U17822 (N_17822,N_16089,N_16889);
and U17823 (N_17823,N_16039,N_16940);
or U17824 (N_17824,N_16310,N_16851);
nor U17825 (N_17825,N_16969,N_16291);
or U17826 (N_17826,N_16190,N_16694);
nor U17827 (N_17827,N_16741,N_16793);
nor U17828 (N_17828,N_16527,N_16928);
or U17829 (N_17829,N_16122,N_16312);
nand U17830 (N_17830,N_16787,N_16840);
and U17831 (N_17831,N_16768,N_16114);
nor U17832 (N_17832,N_16176,N_16359);
or U17833 (N_17833,N_16931,N_16164);
and U17834 (N_17834,N_16097,N_16032);
or U17835 (N_17835,N_16416,N_16105);
nand U17836 (N_17836,N_16601,N_16113);
nor U17837 (N_17837,N_16573,N_16595);
nand U17838 (N_17838,N_16396,N_16804);
or U17839 (N_17839,N_16451,N_16211);
xnor U17840 (N_17840,N_16156,N_16211);
or U17841 (N_17841,N_16530,N_16983);
and U17842 (N_17842,N_16417,N_16891);
xnor U17843 (N_17843,N_16341,N_16739);
xor U17844 (N_17844,N_16296,N_16166);
nor U17845 (N_17845,N_16434,N_16377);
and U17846 (N_17846,N_16632,N_16165);
or U17847 (N_17847,N_16339,N_16723);
nand U17848 (N_17848,N_16418,N_16531);
nand U17849 (N_17849,N_16120,N_16907);
and U17850 (N_17850,N_16674,N_16631);
nor U17851 (N_17851,N_16983,N_16370);
nand U17852 (N_17852,N_16571,N_16491);
or U17853 (N_17853,N_16583,N_16440);
or U17854 (N_17854,N_16218,N_16217);
and U17855 (N_17855,N_16335,N_16017);
and U17856 (N_17856,N_16905,N_16873);
nor U17857 (N_17857,N_16074,N_16016);
nor U17858 (N_17858,N_16929,N_16726);
xor U17859 (N_17859,N_16579,N_16184);
nor U17860 (N_17860,N_16008,N_16823);
nor U17861 (N_17861,N_16029,N_16330);
nand U17862 (N_17862,N_16744,N_16445);
and U17863 (N_17863,N_16249,N_16727);
or U17864 (N_17864,N_16378,N_16415);
or U17865 (N_17865,N_16701,N_16536);
nand U17866 (N_17866,N_16636,N_16020);
or U17867 (N_17867,N_16083,N_16983);
xor U17868 (N_17868,N_16715,N_16275);
nor U17869 (N_17869,N_16977,N_16362);
nor U17870 (N_17870,N_16903,N_16756);
or U17871 (N_17871,N_16418,N_16500);
and U17872 (N_17872,N_16980,N_16550);
and U17873 (N_17873,N_16727,N_16135);
xnor U17874 (N_17874,N_16963,N_16950);
and U17875 (N_17875,N_16479,N_16310);
nor U17876 (N_17876,N_16977,N_16723);
and U17877 (N_17877,N_16661,N_16365);
nand U17878 (N_17878,N_16921,N_16570);
or U17879 (N_17879,N_16843,N_16050);
or U17880 (N_17880,N_16445,N_16322);
nor U17881 (N_17881,N_16251,N_16562);
and U17882 (N_17882,N_16818,N_16745);
nand U17883 (N_17883,N_16548,N_16798);
xnor U17884 (N_17884,N_16783,N_16457);
or U17885 (N_17885,N_16361,N_16662);
or U17886 (N_17886,N_16515,N_16110);
nor U17887 (N_17887,N_16788,N_16520);
and U17888 (N_17888,N_16375,N_16653);
or U17889 (N_17889,N_16167,N_16796);
nor U17890 (N_17890,N_16745,N_16730);
xor U17891 (N_17891,N_16966,N_16968);
and U17892 (N_17892,N_16337,N_16259);
nand U17893 (N_17893,N_16612,N_16316);
nand U17894 (N_17894,N_16612,N_16597);
or U17895 (N_17895,N_16605,N_16545);
nand U17896 (N_17896,N_16022,N_16923);
or U17897 (N_17897,N_16139,N_16869);
nand U17898 (N_17898,N_16227,N_16162);
or U17899 (N_17899,N_16482,N_16346);
xor U17900 (N_17900,N_16651,N_16667);
xor U17901 (N_17901,N_16033,N_16463);
xnor U17902 (N_17902,N_16418,N_16065);
nand U17903 (N_17903,N_16843,N_16167);
or U17904 (N_17904,N_16604,N_16772);
nor U17905 (N_17905,N_16592,N_16104);
nand U17906 (N_17906,N_16770,N_16503);
xnor U17907 (N_17907,N_16061,N_16038);
and U17908 (N_17908,N_16426,N_16923);
or U17909 (N_17909,N_16138,N_16805);
nand U17910 (N_17910,N_16702,N_16473);
xnor U17911 (N_17911,N_16599,N_16849);
and U17912 (N_17912,N_16240,N_16442);
xnor U17913 (N_17913,N_16268,N_16196);
and U17914 (N_17914,N_16747,N_16227);
xor U17915 (N_17915,N_16300,N_16305);
nand U17916 (N_17916,N_16055,N_16525);
and U17917 (N_17917,N_16392,N_16400);
or U17918 (N_17918,N_16853,N_16416);
nor U17919 (N_17919,N_16446,N_16926);
xor U17920 (N_17920,N_16686,N_16560);
and U17921 (N_17921,N_16916,N_16548);
or U17922 (N_17922,N_16912,N_16249);
or U17923 (N_17923,N_16539,N_16532);
nor U17924 (N_17924,N_16611,N_16658);
nor U17925 (N_17925,N_16983,N_16213);
or U17926 (N_17926,N_16656,N_16310);
nand U17927 (N_17927,N_16542,N_16220);
nand U17928 (N_17928,N_16160,N_16215);
nand U17929 (N_17929,N_16887,N_16018);
nor U17930 (N_17930,N_16455,N_16461);
nor U17931 (N_17931,N_16937,N_16986);
or U17932 (N_17932,N_16974,N_16550);
nor U17933 (N_17933,N_16653,N_16250);
xnor U17934 (N_17934,N_16851,N_16898);
nor U17935 (N_17935,N_16133,N_16985);
nand U17936 (N_17936,N_16231,N_16591);
nor U17937 (N_17937,N_16639,N_16202);
xnor U17938 (N_17938,N_16600,N_16649);
and U17939 (N_17939,N_16616,N_16009);
or U17940 (N_17940,N_16652,N_16469);
and U17941 (N_17941,N_16936,N_16662);
and U17942 (N_17942,N_16368,N_16765);
nand U17943 (N_17943,N_16955,N_16066);
and U17944 (N_17944,N_16590,N_16582);
nand U17945 (N_17945,N_16742,N_16455);
nand U17946 (N_17946,N_16376,N_16557);
nor U17947 (N_17947,N_16696,N_16949);
nor U17948 (N_17948,N_16116,N_16725);
xnor U17949 (N_17949,N_16166,N_16206);
nor U17950 (N_17950,N_16301,N_16142);
and U17951 (N_17951,N_16876,N_16240);
nor U17952 (N_17952,N_16511,N_16866);
and U17953 (N_17953,N_16543,N_16986);
nand U17954 (N_17954,N_16076,N_16952);
nor U17955 (N_17955,N_16776,N_16823);
nor U17956 (N_17956,N_16077,N_16302);
or U17957 (N_17957,N_16577,N_16731);
xor U17958 (N_17958,N_16700,N_16099);
or U17959 (N_17959,N_16290,N_16885);
nand U17960 (N_17960,N_16242,N_16021);
nor U17961 (N_17961,N_16984,N_16309);
xnor U17962 (N_17962,N_16828,N_16294);
and U17963 (N_17963,N_16856,N_16612);
xnor U17964 (N_17964,N_16220,N_16335);
nor U17965 (N_17965,N_16957,N_16449);
nand U17966 (N_17966,N_16490,N_16861);
nor U17967 (N_17967,N_16237,N_16865);
and U17968 (N_17968,N_16331,N_16271);
nor U17969 (N_17969,N_16121,N_16973);
nand U17970 (N_17970,N_16232,N_16074);
and U17971 (N_17971,N_16016,N_16708);
xnor U17972 (N_17972,N_16661,N_16316);
nand U17973 (N_17973,N_16130,N_16211);
and U17974 (N_17974,N_16123,N_16173);
xor U17975 (N_17975,N_16619,N_16156);
xor U17976 (N_17976,N_16092,N_16384);
xor U17977 (N_17977,N_16108,N_16935);
xor U17978 (N_17978,N_16394,N_16477);
and U17979 (N_17979,N_16519,N_16686);
xnor U17980 (N_17980,N_16066,N_16742);
and U17981 (N_17981,N_16002,N_16094);
and U17982 (N_17982,N_16178,N_16753);
nor U17983 (N_17983,N_16490,N_16868);
nand U17984 (N_17984,N_16156,N_16275);
and U17985 (N_17985,N_16474,N_16674);
nand U17986 (N_17986,N_16834,N_16610);
nand U17987 (N_17987,N_16939,N_16214);
nand U17988 (N_17988,N_16403,N_16465);
xor U17989 (N_17989,N_16048,N_16158);
nand U17990 (N_17990,N_16208,N_16588);
xor U17991 (N_17991,N_16474,N_16572);
xnor U17992 (N_17992,N_16729,N_16282);
xnor U17993 (N_17993,N_16512,N_16773);
and U17994 (N_17994,N_16377,N_16808);
or U17995 (N_17995,N_16942,N_16598);
xnor U17996 (N_17996,N_16164,N_16209);
or U17997 (N_17997,N_16165,N_16618);
and U17998 (N_17998,N_16231,N_16475);
xor U17999 (N_17999,N_16202,N_16664);
and U18000 (N_18000,N_17011,N_17729);
or U18001 (N_18001,N_17322,N_17596);
or U18002 (N_18002,N_17382,N_17356);
or U18003 (N_18003,N_17180,N_17485);
or U18004 (N_18004,N_17962,N_17978);
xor U18005 (N_18005,N_17034,N_17611);
xor U18006 (N_18006,N_17927,N_17768);
or U18007 (N_18007,N_17987,N_17149);
and U18008 (N_18008,N_17994,N_17607);
and U18009 (N_18009,N_17215,N_17642);
nand U18010 (N_18010,N_17855,N_17067);
and U18011 (N_18011,N_17396,N_17459);
and U18012 (N_18012,N_17571,N_17648);
or U18013 (N_18013,N_17901,N_17033);
nand U18014 (N_18014,N_17995,N_17699);
or U18015 (N_18015,N_17989,N_17092);
or U18016 (N_18016,N_17095,N_17153);
xor U18017 (N_18017,N_17467,N_17991);
nand U18018 (N_18018,N_17531,N_17638);
nor U18019 (N_18019,N_17047,N_17845);
nand U18020 (N_18020,N_17246,N_17264);
and U18021 (N_18021,N_17281,N_17670);
xor U18022 (N_18022,N_17376,N_17713);
or U18023 (N_18023,N_17239,N_17885);
or U18024 (N_18024,N_17619,N_17694);
or U18025 (N_18025,N_17554,N_17380);
xor U18026 (N_18026,N_17850,N_17860);
and U18027 (N_18027,N_17450,N_17959);
nand U18028 (N_18028,N_17480,N_17803);
and U18029 (N_18029,N_17448,N_17552);
and U18030 (N_18030,N_17905,N_17392);
xnor U18031 (N_18031,N_17673,N_17411);
or U18032 (N_18032,N_17135,N_17661);
nor U18033 (N_18033,N_17216,N_17645);
or U18034 (N_18034,N_17605,N_17214);
xnor U18035 (N_18035,N_17224,N_17964);
nor U18036 (N_18036,N_17118,N_17290);
nand U18037 (N_18037,N_17443,N_17430);
and U18038 (N_18038,N_17347,N_17933);
or U18039 (N_18039,N_17136,N_17403);
and U18040 (N_18040,N_17444,N_17874);
nor U18041 (N_18041,N_17494,N_17117);
and U18042 (N_18042,N_17925,N_17379);
nor U18043 (N_18043,N_17078,N_17553);
xnor U18044 (N_18044,N_17132,N_17314);
nand U18045 (N_18045,N_17439,N_17414);
nor U18046 (N_18046,N_17102,N_17779);
nand U18047 (N_18047,N_17723,N_17664);
xnor U18048 (N_18048,N_17853,N_17339);
nor U18049 (N_18049,N_17865,N_17377);
nor U18050 (N_18050,N_17819,N_17837);
or U18051 (N_18051,N_17996,N_17836);
or U18052 (N_18052,N_17847,N_17676);
or U18053 (N_18053,N_17099,N_17076);
xnor U18054 (N_18054,N_17464,N_17911);
or U18055 (N_18055,N_17308,N_17919);
nor U18056 (N_18056,N_17624,N_17728);
and U18057 (N_18057,N_17540,N_17242);
xor U18058 (N_18058,N_17125,N_17882);
and U18059 (N_18059,N_17241,N_17810);
nor U18060 (N_18060,N_17397,N_17710);
nor U18061 (N_18061,N_17566,N_17757);
and U18062 (N_18062,N_17634,N_17975);
or U18063 (N_18063,N_17301,N_17643);
nand U18064 (N_18064,N_17835,N_17963);
nand U18065 (N_18065,N_17981,N_17427);
and U18066 (N_18066,N_17691,N_17876);
and U18067 (N_18067,N_17802,N_17086);
and U18068 (N_18068,N_17019,N_17781);
or U18069 (N_18069,N_17539,N_17415);
xor U18070 (N_18070,N_17830,N_17862);
nor U18071 (N_18071,N_17696,N_17869);
or U18072 (N_18072,N_17460,N_17232);
or U18073 (N_18073,N_17583,N_17159);
or U18074 (N_18074,N_17240,N_17692);
nand U18075 (N_18075,N_17725,N_17808);
xor U18076 (N_18076,N_17668,N_17529);
nand U18077 (N_18077,N_17682,N_17013);
or U18078 (N_18078,N_17533,N_17702);
xor U18079 (N_18079,N_17892,N_17689);
xnor U18080 (N_18080,N_17451,N_17362);
nor U18081 (N_18081,N_17526,N_17740);
and U18082 (N_18082,N_17253,N_17775);
and U18083 (N_18083,N_17857,N_17030);
and U18084 (N_18084,N_17353,N_17103);
xnor U18085 (N_18085,N_17859,N_17334);
nand U18086 (N_18086,N_17832,N_17755);
nand U18087 (N_18087,N_17207,N_17754);
xor U18088 (N_18088,N_17262,N_17982);
and U18089 (N_18089,N_17598,N_17325);
and U18090 (N_18090,N_17595,N_17312);
xor U18091 (N_18091,N_17647,N_17160);
nor U18092 (N_18092,N_17489,N_17897);
or U18093 (N_18093,N_17059,N_17337);
or U18094 (N_18094,N_17195,N_17867);
nor U18095 (N_18095,N_17690,N_17105);
xnor U18096 (N_18096,N_17273,N_17721);
xnor U18097 (N_18097,N_17880,N_17898);
xnor U18098 (N_18098,N_17852,N_17199);
and U18099 (N_18099,N_17499,N_17131);
nor U18100 (N_18100,N_17031,N_17577);
nor U18101 (N_18101,N_17589,N_17795);
or U18102 (N_18102,N_17868,N_17568);
and U18103 (N_18103,N_17493,N_17644);
and U18104 (N_18104,N_17509,N_17157);
xor U18105 (N_18105,N_17049,N_17525);
nor U18106 (N_18106,N_17085,N_17309);
nor U18107 (N_18107,N_17681,N_17208);
xnor U18108 (N_18108,N_17942,N_17594);
or U18109 (N_18109,N_17612,N_17820);
or U18110 (N_18110,N_17759,N_17021);
nand U18111 (N_18111,N_17821,N_17902);
nor U18112 (N_18112,N_17579,N_17999);
nor U18113 (N_18113,N_17413,N_17514);
or U18114 (N_18114,N_17502,N_17338);
or U18115 (N_18115,N_17045,N_17864);
and U18116 (N_18116,N_17395,N_17355);
nor U18117 (N_18117,N_17812,N_17090);
nand U18118 (N_18118,N_17035,N_17747);
xor U18119 (N_18119,N_17561,N_17550);
xnor U18120 (N_18120,N_17546,N_17177);
nor U18121 (N_18121,N_17667,N_17536);
xor U18122 (N_18122,N_17244,N_17635);
xnor U18123 (N_18123,N_17073,N_17712);
and U18124 (N_18124,N_17662,N_17584);
nand U18125 (N_18125,N_17791,N_17907);
nand U18126 (N_18126,N_17777,N_17744);
or U18127 (N_18127,N_17288,N_17703);
or U18128 (N_18128,N_17877,N_17774);
nor U18129 (N_18129,N_17390,N_17425);
nand U18130 (N_18130,N_17929,N_17751);
nand U18131 (N_18131,N_17112,N_17567);
nand U18132 (N_18132,N_17651,N_17471);
and U18133 (N_18133,N_17918,N_17341);
or U18134 (N_18134,N_17437,N_17599);
or U18135 (N_18135,N_17171,N_17766);
or U18136 (N_18136,N_17631,N_17772);
nand U18137 (N_18137,N_17029,N_17084);
and U18138 (N_18138,N_17372,N_17482);
nor U18139 (N_18139,N_17182,N_17655);
xor U18140 (N_18140,N_17449,N_17279);
xnor U18141 (N_18141,N_17063,N_17275);
xnor U18142 (N_18142,N_17993,N_17152);
or U18143 (N_18143,N_17145,N_17887);
xor U18144 (N_18144,N_17789,N_17446);
or U18145 (N_18145,N_17767,N_17894);
and U18146 (N_18146,N_17861,N_17604);
and U18147 (N_18147,N_17475,N_17278);
nand U18148 (N_18148,N_17510,N_17243);
nand U18149 (N_18149,N_17101,N_17018);
and U18150 (N_18150,N_17490,N_17495);
xnor U18151 (N_18151,N_17628,N_17248);
nor U18152 (N_18152,N_17683,N_17792);
or U18153 (N_18153,N_17983,N_17800);
or U18154 (N_18154,N_17373,N_17693);
or U18155 (N_18155,N_17423,N_17004);
nand U18156 (N_18156,N_17816,N_17298);
and U18157 (N_18157,N_17616,N_17293);
nor U18158 (N_18158,N_17824,N_17139);
or U18159 (N_18159,N_17829,N_17585);
and U18160 (N_18160,N_17931,N_17722);
xor U18161 (N_18161,N_17340,N_17948);
xnor U18162 (N_18162,N_17705,N_17187);
and U18163 (N_18163,N_17410,N_17051);
xor U18164 (N_18164,N_17038,N_17237);
nand U18165 (N_18165,N_17787,N_17671);
or U18166 (N_18166,N_17613,N_17303);
or U18167 (N_18167,N_17209,N_17100);
xnor U18168 (N_18168,N_17069,N_17197);
and U18169 (N_18169,N_17156,N_17833);
xor U18170 (N_18170,N_17269,N_17516);
and U18171 (N_18171,N_17822,N_17104);
xor U18172 (N_18172,N_17434,N_17746);
nor U18173 (N_18173,N_17972,N_17297);
nand U18174 (N_18174,N_17026,N_17633);
and U18175 (N_18175,N_17271,N_17923);
nand U18176 (N_18176,N_17809,N_17888);
xor U18177 (N_18177,N_17017,N_17870);
nand U18178 (N_18178,N_17147,N_17399);
and U18179 (N_18179,N_17486,N_17228);
nand U18180 (N_18180,N_17956,N_17827);
xnor U18181 (N_18181,N_17844,N_17198);
or U18182 (N_18182,N_17739,N_17438);
and U18183 (N_18183,N_17790,N_17474);
nor U18184 (N_18184,N_17088,N_17210);
and U18185 (N_18185,N_17071,N_17307);
nor U18186 (N_18186,N_17679,N_17010);
or U18187 (N_18187,N_17569,N_17649);
and U18188 (N_18188,N_17054,N_17386);
or U18189 (N_18189,N_17363,N_17422);
nand U18190 (N_18190,N_17274,N_17134);
nand U18191 (N_18191,N_17174,N_17375);
xnor U18192 (N_18192,N_17706,N_17487);
or U18193 (N_18193,N_17841,N_17517);
and U18194 (N_18194,N_17831,N_17771);
xor U18195 (N_18195,N_17762,N_17277);
xnor U18196 (N_18196,N_17154,N_17609);
xor U18197 (N_18197,N_17939,N_17917);
xnor U18198 (N_18198,N_17914,N_17632);
and U18199 (N_18199,N_17285,N_17732);
nand U18200 (N_18200,N_17249,N_17967);
xnor U18201 (N_18201,N_17416,N_17700);
xnor U18202 (N_18202,N_17626,N_17707);
and U18203 (N_18203,N_17534,N_17093);
nand U18204 (N_18204,N_17736,N_17627);
and U18205 (N_18205,N_17265,N_17150);
nand U18206 (N_18206,N_17137,N_17954);
nand U18207 (N_18207,N_17043,N_17184);
nand U18208 (N_18208,N_17424,N_17960);
nand U18209 (N_18209,N_17878,N_17400);
or U18210 (N_18210,N_17436,N_17476);
nor U18211 (N_18211,N_17223,N_17798);
nor U18212 (N_18212,N_17141,N_17564);
nand U18213 (N_18213,N_17801,N_17014);
nor U18214 (N_18214,N_17406,N_17440);
or U18215 (N_18215,N_17404,N_17606);
or U18216 (N_18216,N_17618,N_17333);
xor U18217 (N_18217,N_17022,N_17283);
or U18218 (N_18218,N_17231,N_17320);
xnor U18219 (N_18219,N_17497,N_17555);
xor U18220 (N_18220,N_17716,N_17167);
nand U18221 (N_18221,N_17973,N_17358);
nor U18222 (N_18222,N_17061,N_17955);
nor U18223 (N_18223,N_17976,N_17393);
xor U18224 (N_18224,N_17701,N_17037);
nand U18225 (N_18225,N_17941,N_17818);
and U18226 (N_18226,N_17122,N_17903);
and U18227 (N_18227,N_17462,N_17621);
or U18228 (N_18228,N_17080,N_17066);
nor U18229 (N_18229,N_17202,N_17773);
xnor U18230 (N_18230,N_17794,N_17254);
xor U18231 (N_18231,N_17922,N_17507);
or U18232 (N_18232,N_17343,N_17630);
nor U18233 (N_18233,N_17496,N_17908);
and U18234 (N_18234,N_17761,N_17221);
xor U18235 (N_18235,N_17985,N_17155);
and U18236 (N_18236,N_17688,N_17515);
xor U18237 (N_18237,N_17009,N_17114);
or U18238 (N_18238,N_17345,N_17201);
xor U18239 (N_18239,N_17335,N_17402);
nand U18240 (N_18240,N_17256,N_17506);
nor U18241 (N_18241,N_17165,N_17371);
nor U18242 (N_18242,N_17697,N_17834);
nand U18243 (N_18243,N_17977,N_17328);
nor U18244 (N_18244,N_17530,N_17558);
or U18245 (N_18245,N_17354,N_17367);
xor U18246 (N_18246,N_17944,N_17058);
and U18247 (N_18247,N_17814,N_17916);
xnor U18248 (N_18248,N_17551,N_17730);
xnor U18249 (N_18249,N_17943,N_17909);
and U18250 (N_18250,N_17512,N_17384);
nand U18251 (N_18251,N_17823,N_17669);
xor U18252 (N_18252,N_17513,N_17565);
and U18253 (N_18253,N_17806,N_17083);
xnor U18254 (N_18254,N_17368,N_17126);
and U18255 (N_18255,N_17257,N_17557);
nor U18256 (N_18256,N_17417,N_17263);
nand U18257 (N_18257,N_17023,N_17650);
xnor U18258 (N_18258,N_17646,N_17087);
and U18259 (N_18259,N_17191,N_17421);
or U18260 (N_18260,N_17468,N_17639);
or U18261 (N_18261,N_17842,N_17574);
nor U18262 (N_18262,N_17268,N_17704);
or U18263 (N_18263,N_17235,N_17484);
nand U18264 (N_18264,N_17350,N_17997);
or U18265 (N_18265,N_17666,N_17286);
and U18266 (N_18266,N_17176,N_17405);
nor U18267 (N_18267,N_17714,N_17840);
or U18268 (N_18268,N_17518,N_17206);
xor U18269 (N_18269,N_17653,N_17726);
nand U18270 (N_18270,N_17299,N_17289);
and U18271 (N_18271,N_17179,N_17111);
xnor U18272 (N_18272,N_17129,N_17096);
nor U18273 (N_18273,N_17734,N_17065);
nor U18274 (N_18274,N_17002,N_17158);
xor U18275 (N_18275,N_17674,N_17077);
and U18276 (N_18276,N_17107,N_17012);
nor U18277 (N_18277,N_17466,N_17280);
and U18278 (N_18278,N_17896,N_17050);
nand U18279 (N_18279,N_17441,N_17326);
nand U18280 (N_18280,N_17053,N_17970);
xor U18281 (N_18281,N_17477,N_17189);
nor U18282 (N_18282,N_17582,N_17252);
xnor U18283 (N_18283,N_17883,N_17979);
nor U18284 (N_18284,N_17151,N_17764);
xnor U18285 (N_18285,N_17799,N_17780);
nor U18286 (N_18286,N_17431,N_17116);
and U18287 (N_18287,N_17259,N_17162);
or U18288 (N_18288,N_17226,N_17057);
nand U18289 (N_18289,N_17270,N_17219);
xnor U18290 (N_18290,N_17005,N_17469);
nor U18291 (N_18291,N_17610,N_17573);
nand U18292 (N_18292,N_17735,N_17986);
nor U18293 (N_18293,N_17294,N_17166);
or U18294 (N_18294,N_17027,N_17586);
xor U18295 (N_18295,N_17200,N_17752);
nand U18296 (N_18296,N_17961,N_17899);
nor U18297 (N_18297,N_17893,N_17447);
xor U18298 (N_18298,N_17319,N_17348);
nand U18299 (N_18299,N_17708,N_17230);
or U18300 (N_18300,N_17760,N_17863);
xnor U18301 (N_18301,N_17081,N_17592);
nor U18302 (N_18302,N_17433,N_17854);
or U18303 (N_18303,N_17741,N_17370);
nand U18304 (N_18304,N_17327,N_17316);
xor U18305 (N_18305,N_17560,N_17074);
or U18306 (N_18306,N_17846,N_17588);
xor U18307 (N_18307,N_17990,N_17342);
xor U18308 (N_18308,N_17538,N_17935);
nand U18309 (N_18309,N_17542,N_17391);
nand U18310 (N_18310,N_17637,N_17520);
and U18311 (N_18311,N_17659,N_17889);
and U18312 (N_18312,N_17251,N_17234);
nor U18313 (N_18313,N_17064,N_17742);
xnor U18314 (N_18314,N_17284,N_17591);
nor U18315 (N_18315,N_17680,N_17938);
and U18316 (N_18316,N_17365,N_17904);
nand U18317 (N_18317,N_17387,N_17848);
or U18318 (N_18318,N_17055,N_17825);
nor U18319 (N_18319,N_17188,N_17937);
nand U18320 (N_18320,N_17305,N_17750);
xor U18321 (N_18321,N_17185,N_17695);
nor U18322 (N_18322,N_17140,N_17315);
nor U18323 (N_18323,N_17193,N_17532);
nor U18324 (N_18324,N_17936,N_17287);
xnor U18325 (N_18325,N_17615,N_17346);
nand U18326 (N_18326,N_17097,N_17389);
or U18327 (N_18327,N_17782,N_17603);
nor U18328 (N_18328,N_17600,N_17543);
and U18329 (N_18329,N_17549,N_17932);
and U18330 (N_18330,N_17212,N_17302);
nor U18331 (N_18331,N_17988,N_17336);
nor U18332 (N_18332,N_17304,N_17470);
nor U18333 (N_18333,N_17324,N_17217);
and U18334 (N_18334,N_17144,N_17119);
nand U18335 (N_18335,N_17590,N_17218);
nor U18336 (N_18336,N_17478,N_17608);
xnor U18337 (N_18337,N_17731,N_17170);
and U18338 (N_18338,N_17974,N_17146);
nor U18339 (N_18339,N_17082,N_17875);
nor U18340 (N_18340,N_17250,N_17547);
nor U18341 (N_18341,N_17383,N_17544);
and U18342 (N_18342,N_17980,N_17811);
nand U18343 (N_18343,N_17900,N_17044);
and U18344 (N_18344,N_17622,N_17205);
and U18345 (N_18345,N_17039,N_17587);
nand U18346 (N_18346,N_17120,N_17041);
nand U18347 (N_18347,N_17108,N_17138);
or U18348 (N_18348,N_17461,N_17310);
and U18349 (N_18349,N_17479,N_17965);
and U18350 (N_18350,N_17492,N_17169);
nor U18351 (N_18351,N_17295,N_17575);
nand U18352 (N_18352,N_17660,N_17665);
nor U18353 (N_18353,N_17472,N_17204);
nor U18354 (N_18354,N_17687,N_17306);
xor U18355 (N_18355,N_17620,N_17617);
and U18356 (N_18356,N_17719,N_17501);
xnor U18357 (N_18357,N_17508,N_17432);
xor U18358 (N_18358,N_17593,N_17048);
nand U18359 (N_18359,N_17717,N_17236);
or U18360 (N_18360,N_17194,N_17727);
and U18361 (N_18361,N_17738,N_17545);
nor U18362 (N_18362,N_17020,N_17419);
xor U18363 (N_18363,N_17656,N_17971);
xor U18364 (N_18364,N_17381,N_17229);
nor U18365 (N_18365,N_17718,N_17452);
and U18366 (N_18366,N_17164,N_17428);
xnor U18367 (N_18367,N_17748,N_17758);
and U18368 (N_18368,N_17890,N_17805);
and U18369 (N_18369,N_17323,N_17412);
nand U18370 (N_18370,N_17511,N_17463);
and U18371 (N_18371,N_17580,N_17527);
nand U18372 (N_18372,N_17886,N_17374);
nor U18373 (N_18373,N_17858,N_17032);
or U18374 (N_18374,N_17926,N_17951);
nor U18375 (N_18375,N_17070,N_17984);
or U18376 (N_18376,N_17351,N_17458);
nand U18377 (N_18377,N_17040,N_17260);
nor U18378 (N_18378,N_17548,N_17946);
nand U18379 (N_18379,N_17578,N_17958);
nor U18380 (N_18380,N_17094,N_17331);
nand U18381 (N_18381,N_17213,N_17756);
nor U18382 (N_18382,N_17839,N_17684);
xnor U18383 (N_18383,N_17124,N_17849);
and U18384 (N_18384,N_17175,N_17778);
and U18385 (N_18385,N_17091,N_17815);
and U18386 (N_18386,N_17016,N_17504);
and U18387 (N_18387,N_17769,N_17998);
and U18388 (N_18388,N_17968,N_17678);
xor U18389 (N_18389,N_17966,N_17245);
nand U18390 (N_18390,N_17969,N_17793);
and U18391 (N_18391,N_17581,N_17409);
or U18392 (N_18392,N_17001,N_17163);
nand U18393 (N_18393,N_17068,N_17359);
xor U18394 (N_18394,N_17025,N_17737);
nand U18395 (N_18395,N_17535,N_17357);
xnor U18396 (N_18396,N_17947,N_17420);
nand U18397 (N_18397,N_17724,N_17385);
and U18398 (N_18398,N_17765,N_17743);
xor U18399 (N_18399,N_17804,N_17042);
or U18400 (N_18400,N_17796,N_17602);
nand U18401 (N_18401,N_17528,N_17491);
nand U18402 (N_18402,N_17161,N_17227);
xnor U18403 (N_18403,N_17006,N_17930);
or U18404 (N_18404,N_17203,N_17953);
and U18405 (N_18405,N_17813,N_17838);
xnor U18406 (N_18406,N_17873,N_17233);
and U18407 (N_18407,N_17292,N_17329);
and U18408 (N_18408,N_17454,N_17675);
nand U18409 (N_18409,N_17106,N_17576);
nand U18410 (N_18410,N_17453,N_17435);
or U18411 (N_18411,N_17807,N_17401);
or U18412 (N_18412,N_17817,N_17465);
nor U18413 (N_18413,N_17503,N_17143);
nor U18414 (N_18414,N_17186,N_17788);
and U18415 (N_18415,N_17113,N_17225);
or U18416 (N_18416,N_17614,N_17949);
or U18417 (N_18417,N_17623,N_17522);
and U18418 (N_18418,N_17686,N_17123);
xnor U18419 (N_18419,N_17318,N_17196);
or U18420 (N_18420,N_17121,N_17473);
and U18421 (N_18421,N_17445,N_17168);
nand U18422 (N_18422,N_17028,N_17915);
nand U18423 (N_18423,N_17709,N_17928);
nand U18424 (N_18424,N_17784,N_17276);
nor U18425 (N_18425,N_17629,N_17426);
or U18426 (N_18426,N_17797,N_17785);
or U18427 (N_18427,N_17408,N_17418);
and U18428 (N_18428,N_17950,N_17313);
xor U18429 (N_18429,N_17776,N_17505);
nor U18430 (N_18430,N_17332,N_17429);
and U18431 (N_18431,N_17843,N_17879);
or U18432 (N_18432,N_17110,N_17183);
xor U18433 (N_18433,N_17211,N_17753);
and U18434 (N_18434,N_17523,N_17172);
and U18435 (N_18435,N_17062,N_17388);
nand U18436 (N_18436,N_17015,N_17181);
and U18437 (N_18437,N_17945,N_17261);
and U18438 (N_18438,N_17733,N_17828);
or U18439 (N_18439,N_17657,N_17992);
nand U18440 (N_18440,N_17321,N_17394);
nor U18441 (N_18441,N_17007,N_17024);
xor U18442 (N_18442,N_17258,N_17570);
nor U18443 (N_18443,N_17036,N_17749);
and U18444 (N_18444,N_17500,N_17524);
nand U18445 (N_18445,N_17130,N_17881);
nor U18446 (N_18446,N_17455,N_17222);
xnor U18447 (N_18447,N_17378,N_17952);
and U18448 (N_18448,N_17247,N_17056);
xnor U18449 (N_18449,N_17072,N_17089);
nand U18450 (N_18450,N_17003,N_17913);
nand U18451 (N_18451,N_17079,N_17672);
xnor U18452 (N_18452,N_17317,N_17488);
nand U18453 (N_18453,N_17763,N_17562);
or U18454 (N_18454,N_17360,N_17895);
nor U18455 (N_18455,N_17891,N_17563);
nand U18456 (N_18456,N_17173,N_17127);
nor U18457 (N_18457,N_17481,N_17745);
xnor U18458 (N_18458,N_17148,N_17349);
xor U18459 (N_18459,N_17000,N_17770);
nand U18460 (N_18460,N_17910,N_17654);
xnor U18461 (N_18461,N_17783,N_17625);
or U18462 (N_18462,N_17060,N_17924);
xor U18463 (N_18463,N_17192,N_17300);
or U18464 (N_18464,N_17920,N_17133);
nor U18465 (N_18465,N_17641,N_17128);
or U18466 (N_18466,N_17851,N_17658);
and U18467 (N_18467,N_17075,N_17685);
xor U18468 (N_18468,N_17912,N_17296);
or U18469 (N_18469,N_17872,N_17267);
and U18470 (N_18470,N_17498,N_17398);
nor U18471 (N_18471,N_17652,N_17330);
or U18472 (N_18472,N_17519,N_17541);
xor U18473 (N_18473,N_17456,N_17369);
or U18474 (N_18474,N_17698,N_17537);
nand U18475 (N_18475,N_17282,N_17407);
or U18476 (N_18476,N_17921,N_17866);
and U18477 (N_18477,N_17109,N_17597);
nand U18478 (N_18478,N_17178,N_17826);
nor U18479 (N_18479,N_17601,N_17715);
nor U18480 (N_18480,N_17640,N_17934);
or U18481 (N_18481,N_17115,N_17008);
xnor U18482 (N_18482,N_17457,N_17442);
or U18483 (N_18483,N_17291,N_17663);
nand U18484 (N_18484,N_17364,N_17521);
and U18485 (N_18485,N_17046,N_17957);
xnor U18486 (N_18486,N_17272,N_17711);
nor U18487 (N_18487,N_17677,N_17190);
nor U18488 (N_18488,N_17361,N_17266);
and U18489 (N_18489,N_17871,N_17142);
or U18490 (N_18490,N_17906,N_17856);
nor U18491 (N_18491,N_17366,N_17344);
nor U18492 (N_18492,N_17311,N_17255);
xor U18493 (N_18493,N_17884,N_17556);
xnor U18494 (N_18494,N_17940,N_17720);
xor U18495 (N_18495,N_17098,N_17572);
nand U18496 (N_18496,N_17238,N_17559);
or U18497 (N_18497,N_17483,N_17052);
nor U18498 (N_18498,N_17352,N_17636);
xnor U18499 (N_18499,N_17220,N_17786);
nand U18500 (N_18500,N_17909,N_17473);
or U18501 (N_18501,N_17299,N_17981);
nand U18502 (N_18502,N_17935,N_17479);
and U18503 (N_18503,N_17215,N_17588);
xnor U18504 (N_18504,N_17560,N_17385);
or U18505 (N_18505,N_17306,N_17417);
and U18506 (N_18506,N_17256,N_17696);
xor U18507 (N_18507,N_17952,N_17241);
or U18508 (N_18508,N_17277,N_17366);
xor U18509 (N_18509,N_17869,N_17511);
nand U18510 (N_18510,N_17441,N_17723);
nand U18511 (N_18511,N_17880,N_17989);
and U18512 (N_18512,N_17983,N_17311);
nor U18513 (N_18513,N_17452,N_17655);
nor U18514 (N_18514,N_17303,N_17604);
and U18515 (N_18515,N_17139,N_17601);
and U18516 (N_18516,N_17725,N_17728);
nand U18517 (N_18517,N_17952,N_17586);
nand U18518 (N_18518,N_17616,N_17122);
and U18519 (N_18519,N_17679,N_17127);
nand U18520 (N_18520,N_17315,N_17974);
and U18521 (N_18521,N_17736,N_17316);
xor U18522 (N_18522,N_17580,N_17686);
xnor U18523 (N_18523,N_17660,N_17146);
or U18524 (N_18524,N_17870,N_17288);
and U18525 (N_18525,N_17151,N_17835);
and U18526 (N_18526,N_17895,N_17054);
nor U18527 (N_18527,N_17828,N_17466);
nand U18528 (N_18528,N_17640,N_17842);
nor U18529 (N_18529,N_17976,N_17424);
nor U18530 (N_18530,N_17164,N_17070);
nor U18531 (N_18531,N_17647,N_17030);
and U18532 (N_18532,N_17250,N_17225);
or U18533 (N_18533,N_17964,N_17995);
nor U18534 (N_18534,N_17743,N_17119);
xnor U18535 (N_18535,N_17901,N_17497);
xnor U18536 (N_18536,N_17173,N_17653);
xor U18537 (N_18537,N_17457,N_17261);
or U18538 (N_18538,N_17768,N_17093);
nand U18539 (N_18539,N_17943,N_17916);
xnor U18540 (N_18540,N_17812,N_17270);
xnor U18541 (N_18541,N_17896,N_17286);
nor U18542 (N_18542,N_17166,N_17224);
or U18543 (N_18543,N_17355,N_17963);
and U18544 (N_18544,N_17972,N_17876);
nand U18545 (N_18545,N_17997,N_17305);
nor U18546 (N_18546,N_17808,N_17503);
nand U18547 (N_18547,N_17162,N_17532);
xor U18548 (N_18548,N_17594,N_17473);
and U18549 (N_18549,N_17683,N_17820);
or U18550 (N_18550,N_17284,N_17445);
nor U18551 (N_18551,N_17361,N_17924);
and U18552 (N_18552,N_17154,N_17545);
nor U18553 (N_18553,N_17283,N_17126);
nand U18554 (N_18554,N_17293,N_17549);
xnor U18555 (N_18555,N_17391,N_17071);
or U18556 (N_18556,N_17466,N_17737);
nor U18557 (N_18557,N_17469,N_17212);
or U18558 (N_18558,N_17752,N_17219);
and U18559 (N_18559,N_17414,N_17391);
nand U18560 (N_18560,N_17830,N_17122);
nor U18561 (N_18561,N_17301,N_17502);
or U18562 (N_18562,N_17439,N_17250);
and U18563 (N_18563,N_17140,N_17914);
xnor U18564 (N_18564,N_17855,N_17050);
nand U18565 (N_18565,N_17113,N_17039);
nor U18566 (N_18566,N_17246,N_17232);
nor U18567 (N_18567,N_17953,N_17775);
or U18568 (N_18568,N_17223,N_17679);
or U18569 (N_18569,N_17229,N_17989);
nand U18570 (N_18570,N_17398,N_17987);
xnor U18571 (N_18571,N_17128,N_17040);
nor U18572 (N_18572,N_17835,N_17494);
and U18573 (N_18573,N_17321,N_17412);
and U18574 (N_18574,N_17570,N_17646);
nand U18575 (N_18575,N_17244,N_17580);
nor U18576 (N_18576,N_17302,N_17209);
nand U18577 (N_18577,N_17499,N_17663);
nand U18578 (N_18578,N_17010,N_17557);
or U18579 (N_18579,N_17865,N_17581);
or U18580 (N_18580,N_17152,N_17140);
xnor U18581 (N_18581,N_17150,N_17988);
nand U18582 (N_18582,N_17119,N_17714);
xor U18583 (N_18583,N_17195,N_17234);
nor U18584 (N_18584,N_17658,N_17754);
nand U18585 (N_18585,N_17934,N_17288);
nor U18586 (N_18586,N_17286,N_17094);
nor U18587 (N_18587,N_17963,N_17228);
or U18588 (N_18588,N_17259,N_17760);
nand U18589 (N_18589,N_17540,N_17260);
nor U18590 (N_18590,N_17709,N_17252);
nor U18591 (N_18591,N_17722,N_17892);
and U18592 (N_18592,N_17180,N_17432);
nand U18593 (N_18593,N_17953,N_17114);
and U18594 (N_18594,N_17426,N_17614);
xor U18595 (N_18595,N_17554,N_17920);
xor U18596 (N_18596,N_17001,N_17523);
xnor U18597 (N_18597,N_17544,N_17220);
nor U18598 (N_18598,N_17185,N_17588);
nand U18599 (N_18599,N_17988,N_17971);
nor U18600 (N_18600,N_17060,N_17109);
xnor U18601 (N_18601,N_17983,N_17403);
nor U18602 (N_18602,N_17011,N_17717);
nor U18603 (N_18603,N_17576,N_17248);
or U18604 (N_18604,N_17518,N_17061);
and U18605 (N_18605,N_17148,N_17109);
xnor U18606 (N_18606,N_17249,N_17075);
or U18607 (N_18607,N_17310,N_17453);
or U18608 (N_18608,N_17651,N_17812);
and U18609 (N_18609,N_17488,N_17058);
xnor U18610 (N_18610,N_17889,N_17743);
nor U18611 (N_18611,N_17910,N_17012);
nor U18612 (N_18612,N_17593,N_17544);
or U18613 (N_18613,N_17280,N_17607);
or U18614 (N_18614,N_17397,N_17800);
nand U18615 (N_18615,N_17350,N_17456);
nand U18616 (N_18616,N_17330,N_17257);
or U18617 (N_18617,N_17064,N_17056);
nor U18618 (N_18618,N_17818,N_17862);
nand U18619 (N_18619,N_17280,N_17987);
nand U18620 (N_18620,N_17322,N_17250);
nor U18621 (N_18621,N_17967,N_17076);
nand U18622 (N_18622,N_17990,N_17589);
nor U18623 (N_18623,N_17900,N_17411);
nand U18624 (N_18624,N_17927,N_17046);
and U18625 (N_18625,N_17842,N_17554);
or U18626 (N_18626,N_17792,N_17681);
and U18627 (N_18627,N_17951,N_17458);
nand U18628 (N_18628,N_17283,N_17217);
or U18629 (N_18629,N_17153,N_17177);
xnor U18630 (N_18630,N_17563,N_17259);
nand U18631 (N_18631,N_17786,N_17707);
or U18632 (N_18632,N_17539,N_17690);
and U18633 (N_18633,N_17276,N_17873);
nor U18634 (N_18634,N_17757,N_17960);
xor U18635 (N_18635,N_17219,N_17073);
and U18636 (N_18636,N_17947,N_17850);
or U18637 (N_18637,N_17880,N_17126);
nor U18638 (N_18638,N_17926,N_17554);
and U18639 (N_18639,N_17258,N_17226);
or U18640 (N_18640,N_17165,N_17931);
nor U18641 (N_18641,N_17503,N_17110);
nor U18642 (N_18642,N_17676,N_17752);
and U18643 (N_18643,N_17819,N_17002);
nand U18644 (N_18644,N_17588,N_17136);
and U18645 (N_18645,N_17789,N_17083);
or U18646 (N_18646,N_17509,N_17405);
and U18647 (N_18647,N_17431,N_17017);
nor U18648 (N_18648,N_17671,N_17409);
nand U18649 (N_18649,N_17862,N_17605);
nand U18650 (N_18650,N_17475,N_17787);
or U18651 (N_18651,N_17071,N_17480);
and U18652 (N_18652,N_17905,N_17688);
nand U18653 (N_18653,N_17486,N_17741);
xnor U18654 (N_18654,N_17316,N_17776);
and U18655 (N_18655,N_17482,N_17481);
or U18656 (N_18656,N_17810,N_17048);
and U18657 (N_18657,N_17290,N_17937);
nand U18658 (N_18658,N_17810,N_17486);
and U18659 (N_18659,N_17435,N_17155);
nand U18660 (N_18660,N_17962,N_17380);
xor U18661 (N_18661,N_17174,N_17749);
xnor U18662 (N_18662,N_17627,N_17971);
nor U18663 (N_18663,N_17471,N_17503);
xnor U18664 (N_18664,N_17490,N_17535);
nand U18665 (N_18665,N_17912,N_17896);
nor U18666 (N_18666,N_17281,N_17065);
nand U18667 (N_18667,N_17427,N_17728);
nand U18668 (N_18668,N_17335,N_17458);
or U18669 (N_18669,N_17301,N_17893);
and U18670 (N_18670,N_17701,N_17421);
or U18671 (N_18671,N_17338,N_17495);
xor U18672 (N_18672,N_17619,N_17232);
or U18673 (N_18673,N_17134,N_17361);
or U18674 (N_18674,N_17725,N_17753);
or U18675 (N_18675,N_17843,N_17570);
and U18676 (N_18676,N_17060,N_17876);
or U18677 (N_18677,N_17529,N_17322);
xnor U18678 (N_18678,N_17693,N_17997);
xnor U18679 (N_18679,N_17856,N_17952);
nor U18680 (N_18680,N_17664,N_17347);
nand U18681 (N_18681,N_17584,N_17729);
nor U18682 (N_18682,N_17643,N_17175);
nand U18683 (N_18683,N_17500,N_17622);
nor U18684 (N_18684,N_17417,N_17832);
nand U18685 (N_18685,N_17534,N_17469);
and U18686 (N_18686,N_17328,N_17910);
or U18687 (N_18687,N_17659,N_17574);
nor U18688 (N_18688,N_17472,N_17186);
xnor U18689 (N_18689,N_17951,N_17994);
and U18690 (N_18690,N_17963,N_17149);
nand U18691 (N_18691,N_17593,N_17030);
or U18692 (N_18692,N_17473,N_17285);
nor U18693 (N_18693,N_17074,N_17873);
and U18694 (N_18694,N_17029,N_17930);
nor U18695 (N_18695,N_17304,N_17777);
or U18696 (N_18696,N_17246,N_17446);
or U18697 (N_18697,N_17930,N_17993);
nand U18698 (N_18698,N_17016,N_17863);
nor U18699 (N_18699,N_17093,N_17413);
nor U18700 (N_18700,N_17563,N_17572);
or U18701 (N_18701,N_17651,N_17693);
nand U18702 (N_18702,N_17576,N_17050);
nand U18703 (N_18703,N_17632,N_17511);
or U18704 (N_18704,N_17899,N_17906);
and U18705 (N_18705,N_17767,N_17552);
nor U18706 (N_18706,N_17304,N_17117);
nor U18707 (N_18707,N_17032,N_17296);
or U18708 (N_18708,N_17235,N_17222);
and U18709 (N_18709,N_17664,N_17547);
nand U18710 (N_18710,N_17357,N_17519);
xnor U18711 (N_18711,N_17166,N_17606);
xor U18712 (N_18712,N_17767,N_17328);
or U18713 (N_18713,N_17236,N_17828);
and U18714 (N_18714,N_17535,N_17590);
nor U18715 (N_18715,N_17673,N_17105);
xnor U18716 (N_18716,N_17892,N_17112);
nand U18717 (N_18717,N_17523,N_17430);
xor U18718 (N_18718,N_17099,N_17451);
xor U18719 (N_18719,N_17107,N_17286);
nor U18720 (N_18720,N_17835,N_17265);
nor U18721 (N_18721,N_17086,N_17580);
and U18722 (N_18722,N_17150,N_17645);
nand U18723 (N_18723,N_17002,N_17680);
xnor U18724 (N_18724,N_17251,N_17546);
and U18725 (N_18725,N_17049,N_17483);
xnor U18726 (N_18726,N_17376,N_17122);
xor U18727 (N_18727,N_17854,N_17806);
nor U18728 (N_18728,N_17489,N_17316);
xnor U18729 (N_18729,N_17290,N_17521);
nand U18730 (N_18730,N_17556,N_17071);
and U18731 (N_18731,N_17212,N_17829);
nand U18732 (N_18732,N_17304,N_17667);
xor U18733 (N_18733,N_17847,N_17732);
nand U18734 (N_18734,N_17998,N_17824);
nand U18735 (N_18735,N_17680,N_17796);
nor U18736 (N_18736,N_17089,N_17994);
nor U18737 (N_18737,N_17780,N_17654);
and U18738 (N_18738,N_17215,N_17958);
nand U18739 (N_18739,N_17986,N_17243);
nor U18740 (N_18740,N_17602,N_17165);
xnor U18741 (N_18741,N_17540,N_17149);
nor U18742 (N_18742,N_17504,N_17339);
or U18743 (N_18743,N_17952,N_17170);
nor U18744 (N_18744,N_17554,N_17718);
nand U18745 (N_18745,N_17831,N_17093);
and U18746 (N_18746,N_17928,N_17822);
and U18747 (N_18747,N_17526,N_17619);
nor U18748 (N_18748,N_17843,N_17061);
nor U18749 (N_18749,N_17907,N_17675);
xnor U18750 (N_18750,N_17213,N_17779);
xnor U18751 (N_18751,N_17943,N_17794);
nor U18752 (N_18752,N_17620,N_17112);
or U18753 (N_18753,N_17857,N_17373);
nor U18754 (N_18754,N_17923,N_17217);
or U18755 (N_18755,N_17478,N_17844);
or U18756 (N_18756,N_17978,N_17029);
or U18757 (N_18757,N_17251,N_17414);
xnor U18758 (N_18758,N_17810,N_17308);
or U18759 (N_18759,N_17612,N_17347);
nor U18760 (N_18760,N_17543,N_17840);
or U18761 (N_18761,N_17594,N_17589);
xor U18762 (N_18762,N_17572,N_17260);
or U18763 (N_18763,N_17771,N_17101);
nand U18764 (N_18764,N_17521,N_17717);
nand U18765 (N_18765,N_17637,N_17086);
xnor U18766 (N_18766,N_17326,N_17256);
xor U18767 (N_18767,N_17951,N_17264);
and U18768 (N_18768,N_17506,N_17831);
xnor U18769 (N_18769,N_17735,N_17288);
and U18770 (N_18770,N_17371,N_17063);
xor U18771 (N_18771,N_17133,N_17980);
nand U18772 (N_18772,N_17466,N_17888);
xnor U18773 (N_18773,N_17304,N_17223);
nor U18774 (N_18774,N_17420,N_17798);
nand U18775 (N_18775,N_17506,N_17317);
nand U18776 (N_18776,N_17666,N_17925);
nor U18777 (N_18777,N_17379,N_17817);
nor U18778 (N_18778,N_17553,N_17213);
nand U18779 (N_18779,N_17029,N_17812);
nor U18780 (N_18780,N_17809,N_17752);
and U18781 (N_18781,N_17241,N_17766);
nor U18782 (N_18782,N_17017,N_17370);
and U18783 (N_18783,N_17023,N_17099);
xnor U18784 (N_18784,N_17194,N_17939);
nand U18785 (N_18785,N_17190,N_17116);
xnor U18786 (N_18786,N_17911,N_17979);
nor U18787 (N_18787,N_17096,N_17371);
nand U18788 (N_18788,N_17245,N_17488);
and U18789 (N_18789,N_17399,N_17758);
nor U18790 (N_18790,N_17830,N_17838);
nor U18791 (N_18791,N_17211,N_17236);
and U18792 (N_18792,N_17086,N_17711);
and U18793 (N_18793,N_17228,N_17184);
nand U18794 (N_18794,N_17726,N_17306);
nor U18795 (N_18795,N_17553,N_17159);
or U18796 (N_18796,N_17571,N_17546);
and U18797 (N_18797,N_17672,N_17816);
xor U18798 (N_18798,N_17348,N_17861);
or U18799 (N_18799,N_17669,N_17517);
nand U18800 (N_18800,N_17922,N_17190);
or U18801 (N_18801,N_17006,N_17985);
xnor U18802 (N_18802,N_17854,N_17106);
nor U18803 (N_18803,N_17537,N_17337);
or U18804 (N_18804,N_17278,N_17405);
xnor U18805 (N_18805,N_17780,N_17204);
nand U18806 (N_18806,N_17322,N_17863);
and U18807 (N_18807,N_17619,N_17150);
nor U18808 (N_18808,N_17618,N_17700);
and U18809 (N_18809,N_17433,N_17813);
nor U18810 (N_18810,N_17795,N_17825);
nand U18811 (N_18811,N_17340,N_17598);
nor U18812 (N_18812,N_17713,N_17596);
nand U18813 (N_18813,N_17749,N_17492);
xor U18814 (N_18814,N_17811,N_17917);
and U18815 (N_18815,N_17768,N_17622);
nor U18816 (N_18816,N_17605,N_17341);
or U18817 (N_18817,N_17306,N_17289);
or U18818 (N_18818,N_17719,N_17098);
and U18819 (N_18819,N_17120,N_17978);
and U18820 (N_18820,N_17433,N_17081);
or U18821 (N_18821,N_17926,N_17831);
nor U18822 (N_18822,N_17238,N_17080);
or U18823 (N_18823,N_17615,N_17551);
xor U18824 (N_18824,N_17741,N_17363);
nand U18825 (N_18825,N_17385,N_17958);
nor U18826 (N_18826,N_17809,N_17801);
and U18827 (N_18827,N_17940,N_17642);
xor U18828 (N_18828,N_17522,N_17960);
or U18829 (N_18829,N_17881,N_17699);
xor U18830 (N_18830,N_17319,N_17905);
nor U18831 (N_18831,N_17771,N_17601);
nand U18832 (N_18832,N_17935,N_17986);
nor U18833 (N_18833,N_17947,N_17611);
and U18834 (N_18834,N_17194,N_17776);
xnor U18835 (N_18835,N_17221,N_17300);
and U18836 (N_18836,N_17850,N_17679);
or U18837 (N_18837,N_17357,N_17723);
nand U18838 (N_18838,N_17890,N_17311);
nand U18839 (N_18839,N_17721,N_17871);
or U18840 (N_18840,N_17418,N_17404);
xnor U18841 (N_18841,N_17722,N_17008);
or U18842 (N_18842,N_17759,N_17317);
and U18843 (N_18843,N_17593,N_17275);
and U18844 (N_18844,N_17711,N_17982);
or U18845 (N_18845,N_17070,N_17925);
xor U18846 (N_18846,N_17197,N_17329);
nor U18847 (N_18847,N_17453,N_17259);
and U18848 (N_18848,N_17935,N_17991);
nor U18849 (N_18849,N_17435,N_17717);
xor U18850 (N_18850,N_17313,N_17844);
and U18851 (N_18851,N_17445,N_17665);
xor U18852 (N_18852,N_17719,N_17616);
xor U18853 (N_18853,N_17502,N_17588);
nand U18854 (N_18854,N_17213,N_17338);
and U18855 (N_18855,N_17334,N_17258);
nand U18856 (N_18856,N_17971,N_17858);
nor U18857 (N_18857,N_17515,N_17854);
nand U18858 (N_18858,N_17248,N_17600);
nor U18859 (N_18859,N_17857,N_17485);
and U18860 (N_18860,N_17908,N_17012);
and U18861 (N_18861,N_17742,N_17399);
and U18862 (N_18862,N_17724,N_17239);
or U18863 (N_18863,N_17900,N_17905);
or U18864 (N_18864,N_17593,N_17872);
and U18865 (N_18865,N_17227,N_17000);
nand U18866 (N_18866,N_17510,N_17889);
nor U18867 (N_18867,N_17762,N_17966);
nand U18868 (N_18868,N_17202,N_17338);
nand U18869 (N_18869,N_17118,N_17505);
xnor U18870 (N_18870,N_17983,N_17454);
or U18871 (N_18871,N_17814,N_17069);
or U18872 (N_18872,N_17320,N_17245);
and U18873 (N_18873,N_17896,N_17391);
nor U18874 (N_18874,N_17736,N_17405);
or U18875 (N_18875,N_17383,N_17275);
nor U18876 (N_18876,N_17133,N_17178);
nor U18877 (N_18877,N_17632,N_17015);
or U18878 (N_18878,N_17720,N_17372);
nand U18879 (N_18879,N_17171,N_17623);
nor U18880 (N_18880,N_17916,N_17371);
xnor U18881 (N_18881,N_17586,N_17624);
or U18882 (N_18882,N_17609,N_17536);
xor U18883 (N_18883,N_17089,N_17660);
xor U18884 (N_18884,N_17290,N_17517);
and U18885 (N_18885,N_17212,N_17668);
and U18886 (N_18886,N_17789,N_17435);
xor U18887 (N_18887,N_17661,N_17032);
nor U18888 (N_18888,N_17422,N_17977);
nand U18889 (N_18889,N_17319,N_17914);
nor U18890 (N_18890,N_17310,N_17548);
xnor U18891 (N_18891,N_17395,N_17197);
and U18892 (N_18892,N_17603,N_17659);
or U18893 (N_18893,N_17769,N_17851);
nand U18894 (N_18894,N_17310,N_17184);
or U18895 (N_18895,N_17667,N_17423);
or U18896 (N_18896,N_17929,N_17809);
or U18897 (N_18897,N_17120,N_17307);
xor U18898 (N_18898,N_17900,N_17708);
and U18899 (N_18899,N_17994,N_17729);
or U18900 (N_18900,N_17891,N_17643);
or U18901 (N_18901,N_17813,N_17812);
nor U18902 (N_18902,N_17416,N_17797);
nand U18903 (N_18903,N_17765,N_17470);
xor U18904 (N_18904,N_17921,N_17870);
nand U18905 (N_18905,N_17698,N_17368);
nor U18906 (N_18906,N_17267,N_17905);
nand U18907 (N_18907,N_17528,N_17839);
nor U18908 (N_18908,N_17659,N_17346);
xnor U18909 (N_18909,N_17032,N_17287);
xor U18910 (N_18910,N_17579,N_17991);
nor U18911 (N_18911,N_17594,N_17669);
nor U18912 (N_18912,N_17591,N_17089);
nand U18913 (N_18913,N_17934,N_17950);
or U18914 (N_18914,N_17296,N_17231);
xor U18915 (N_18915,N_17055,N_17992);
and U18916 (N_18916,N_17398,N_17666);
xnor U18917 (N_18917,N_17855,N_17403);
xor U18918 (N_18918,N_17353,N_17681);
and U18919 (N_18919,N_17501,N_17088);
or U18920 (N_18920,N_17094,N_17129);
nand U18921 (N_18921,N_17916,N_17026);
and U18922 (N_18922,N_17302,N_17102);
and U18923 (N_18923,N_17910,N_17079);
nand U18924 (N_18924,N_17168,N_17646);
xor U18925 (N_18925,N_17344,N_17833);
nand U18926 (N_18926,N_17267,N_17083);
or U18927 (N_18927,N_17092,N_17990);
nand U18928 (N_18928,N_17861,N_17143);
nand U18929 (N_18929,N_17035,N_17120);
nor U18930 (N_18930,N_17946,N_17927);
or U18931 (N_18931,N_17095,N_17319);
nor U18932 (N_18932,N_17900,N_17307);
and U18933 (N_18933,N_17851,N_17674);
nand U18934 (N_18934,N_17729,N_17959);
xor U18935 (N_18935,N_17242,N_17924);
xnor U18936 (N_18936,N_17947,N_17070);
and U18937 (N_18937,N_17915,N_17606);
xnor U18938 (N_18938,N_17070,N_17894);
and U18939 (N_18939,N_17728,N_17046);
xnor U18940 (N_18940,N_17184,N_17351);
nor U18941 (N_18941,N_17858,N_17997);
nor U18942 (N_18942,N_17849,N_17063);
nor U18943 (N_18943,N_17530,N_17068);
and U18944 (N_18944,N_17163,N_17018);
xor U18945 (N_18945,N_17986,N_17833);
and U18946 (N_18946,N_17311,N_17304);
or U18947 (N_18947,N_17724,N_17335);
nor U18948 (N_18948,N_17923,N_17709);
or U18949 (N_18949,N_17594,N_17220);
xor U18950 (N_18950,N_17931,N_17694);
nand U18951 (N_18951,N_17297,N_17787);
nand U18952 (N_18952,N_17310,N_17918);
nand U18953 (N_18953,N_17003,N_17593);
or U18954 (N_18954,N_17816,N_17621);
and U18955 (N_18955,N_17003,N_17566);
nor U18956 (N_18956,N_17520,N_17630);
nor U18957 (N_18957,N_17824,N_17043);
nor U18958 (N_18958,N_17853,N_17239);
xor U18959 (N_18959,N_17794,N_17704);
xnor U18960 (N_18960,N_17157,N_17898);
xnor U18961 (N_18961,N_17759,N_17633);
nor U18962 (N_18962,N_17909,N_17985);
nand U18963 (N_18963,N_17391,N_17647);
nand U18964 (N_18964,N_17678,N_17835);
nand U18965 (N_18965,N_17254,N_17660);
xor U18966 (N_18966,N_17908,N_17073);
nor U18967 (N_18967,N_17689,N_17241);
and U18968 (N_18968,N_17712,N_17255);
nor U18969 (N_18969,N_17454,N_17640);
xor U18970 (N_18970,N_17711,N_17435);
and U18971 (N_18971,N_17018,N_17395);
and U18972 (N_18972,N_17479,N_17062);
nor U18973 (N_18973,N_17723,N_17030);
or U18974 (N_18974,N_17092,N_17579);
nand U18975 (N_18975,N_17308,N_17820);
or U18976 (N_18976,N_17445,N_17185);
nand U18977 (N_18977,N_17151,N_17765);
or U18978 (N_18978,N_17182,N_17288);
nor U18979 (N_18979,N_17542,N_17596);
nor U18980 (N_18980,N_17359,N_17159);
nor U18981 (N_18981,N_17820,N_17444);
nor U18982 (N_18982,N_17941,N_17882);
nand U18983 (N_18983,N_17116,N_17485);
xnor U18984 (N_18984,N_17697,N_17555);
and U18985 (N_18985,N_17817,N_17978);
or U18986 (N_18986,N_17724,N_17723);
xnor U18987 (N_18987,N_17311,N_17057);
xor U18988 (N_18988,N_17367,N_17961);
and U18989 (N_18989,N_17139,N_17003);
nor U18990 (N_18990,N_17689,N_17703);
or U18991 (N_18991,N_17251,N_17613);
nand U18992 (N_18992,N_17824,N_17124);
xor U18993 (N_18993,N_17366,N_17462);
nand U18994 (N_18994,N_17866,N_17955);
xor U18995 (N_18995,N_17464,N_17343);
or U18996 (N_18996,N_17086,N_17335);
or U18997 (N_18997,N_17460,N_17512);
nor U18998 (N_18998,N_17806,N_17200);
nand U18999 (N_18999,N_17105,N_17733);
nand U19000 (N_19000,N_18837,N_18066);
nand U19001 (N_19001,N_18899,N_18523);
and U19002 (N_19002,N_18862,N_18611);
xor U19003 (N_19003,N_18627,N_18392);
nor U19004 (N_19004,N_18120,N_18993);
or U19005 (N_19005,N_18635,N_18548);
nand U19006 (N_19006,N_18775,N_18579);
xnor U19007 (N_19007,N_18310,N_18081);
nand U19008 (N_19008,N_18337,N_18923);
xor U19009 (N_19009,N_18061,N_18686);
xor U19010 (N_19010,N_18535,N_18035);
and U19011 (N_19011,N_18164,N_18677);
and U19012 (N_19012,N_18400,N_18491);
xor U19013 (N_19013,N_18090,N_18986);
nand U19014 (N_19014,N_18209,N_18052);
nor U19015 (N_19015,N_18303,N_18435);
xnor U19016 (N_19016,N_18600,N_18177);
xor U19017 (N_19017,N_18628,N_18722);
xor U19018 (N_19018,N_18465,N_18846);
xor U19019 (N_19019,N_18985,N_18918);
and U19020 (N_19020,N_18625,N_18317);
and U19021 (N_19021,N_18786,N_18530);
and U19022 (N_19022,N_18049,N_18217);
nand U19023 (N_19023,N_18683,N_18972);
nor U19024 (N_19024,N_18716,N_18723);
nand U19025 (N_19025,N_18223,N_18495);
xnor U19026 (N_19026,N_18371,N_18352);
or U19027 (N_19027,N_18962,N_18332);
and U19028 (N_19028,N_18642,N_18030);
or U19029 (N_19029,N_18142,N_18037);
or U19030 (N_19030,N_18071,N_18069);
and U19031 (N_19031,N_18411,N_18025);
or U19032 (N_19032,N_18931,N_18092);
xor U19033 (N_19033,N_18898,N_18318);
or U19034 (N_19034,N_18018,N_18552);
or U19035 (N_19035,N_18678,N_18533);
xor U19036 (N_19036,N_18656,N_18793);
nor U19037 (N_19037,N_18199,N_18784);
nand U19038 (N_19038,N_18129,N_18612);
and U19039 (N_19039,N_18867,N_18155);
nand U19040 (N_19040,N_18850,N_18334);
xor U19041 (N_19041,N_18618,N_18203);
xnor U19042 (N_19042,N_18496,N_18950);
or U19043 (N_19043,N_18865,N_18198);
nor U19044 (N_19044,N_18944,N_18331);
nor U19045 (N_19045,N_18514,N_18562);
or U19046 (N_19046,N_18991,N_18373);
nand U19047 (N_19047,N_18802,N_18320);
and U19048 (N_19048,N_18606,N_18688);
or U19049 (N_19049,N_18104,N_18238);
xor U19050 (N_19050,N_18988,N_18106);
or U19051 (N_19051,N_18692,N_18345);
xor U19052 (N_19052,N_18679,N_18195);
xnor U19053 (N_19053,N_18834,N_18302);
nor U19054 (N_19054,N_18829,N_18489);
or U19055 (N_19055,N_18614,N_18433);
nor U19056 (N_19056,N_18509,N_18116);
nand U19057 (N_19057,N_18809,N_18580);
xnor U19058 (N_19058,N_18251,N_18445);
nand U19059 (N_19059,N_18304,N_18135);
and U19060 (N_19060,N_18560,N_18827);
nor U19061 (N_19061,N_18875,N_18715);
or U19062 (N_19062,N_18022,N_18570);
or U19063 (N_19063,N_18211,N_18202);
nor U19064 (N_19064,N_18836,N_18425);
or U19065 (N_19065,N_18736,N_18498);
and U19066 (N_19066,N_18443,N_18741);
xor U19067 (N_19067,N_18339,N_18000);
nor U19068 (N_19068,N_18272,N_18516);
nand U19069 (N_19069,N_18743,N_18316);
xor U19070 (N_19070,N_18055,N_18609);
nand U19071 (N_19071,N_18270,N_18946);
or U19072 (N_19072,N_18776,N_18146);
and U19073 (N_19073,N_18232,N_18349);
nand U19074 (N_19074,N_18161,N_18650);
nor U19075 (N_19075,N_18219,N_18529);
and U19076 (N_19076,N_18454,N_18595);
nor U19077 (N_19077,N_18541,N_18321);
and U19078 (N_19078,N_18814,N_18540);
nor U19079 (N_19079,N_18021,N_18015);
nand U19080 (N_19080,N_18093,N_18763);
nand U19081 (N_19081,N_18921,N_18453);
nand U19082 (N_19082,N_18156,N_18997);
or U19083 (N_19083,N_18102,N_18706);
nor U19084 (N_19084,N_18592,N_18010);
nand U19085 (N_19085,N_18521,N_18571);
and U19086 (N_19086,N_18978,N_18101);
nand U19087 (N_19087,N_18182,N_18306);
nor U19088 (N_19088,N_18404,N_18584);
and U19089 (N_19089,N_18911,N_18315);
or U19090 (N_19090,N_18075,N_18860);
and U19091 (N_19091,N_18599,N_18452);
or U19092 (N_19092,N_18705,N_18690);
xnor U19093 (N_19093,N_18577,N_18231);
nand U19094 (N_19094,N_18294,N_18328);
nor U19095 (N_19095,N_18805,N_18649);
xnor U19096 (N_19096,N_18630,N_18386);
xnor U19097 (N_19097,N_18131,N_18620);
xor U19098 (N_19098,N_18765,N_18589);
or U19099 (N_19099,N_18994,N_18651);
nand U19100 (N_19100,N_18242,N_18711);
and U19101 (N_19101,N_18534,N_18712);
nand U19102 (N_19102,N_18007,N_18419);
nor U19103 (N_19103,N_18138,N_18378);
and U19104 (N_19104,N_18522,N_18338);
or U19105 (N_19105,N_18812,N_18664);
or U19106 (N_19106,N_18346,N_18308);
and U19107 (N_19107,N_18740,N_18727);
xor U19108 (N_19108,N_18753,N_18429);
nor U19109 (N_19109,N_18890,N_18781);
nor U19110 (N_19110,N_18083,N_18681);
xor U19111 (N_19111,N_18633,N_18363);
or U19112 (N_19112,N_18808,N_18162);
xnor U19113 (N_19113,N_18250,N_18047);
or U19114 (N_19114,N_18665,N_18148);
xnor U19115 (N_19115,N_18257,N_18476);
nor U19116 (N_19116,N_18369,N_18983);
and U19117 (N_19117,N_18907,N_18732);
and U19118 (N_19118,N_18504,N_18224);
and U19119 (N_19119,N_18569,N_18210);
or U19120 (N_19120,N_18896,N_18894);
and U19121 (N_19121,N_18256,N_18414);
nand U19122 (N_19122,N_18998,N_18428);
xnor U19123 (N_19123,N_18141,N_18268);
or U19124 (N_19124,N_18544,N_18613);
nor U19125 (N_19125,N_18221,N_18641);
or U19126 (N_19126,N_18418,N_18309);
and U19127 (N_19127,N_18391,N_18745);
nand U19128 (N_19128,N_18032,N_18855);
and U19129 (N_19129,N_18974,N_18758);
xnor U19130 (N_19130,N_18943,N_18130);
nand U19131 (N_19131,N_18942,N_18228);
xor U19132 (N_19132,N_18960,N_18340);
nand U19133 (N_19133,N_18149,N_18167);
or U19134 (N_19134,N_18285,N_18700);
and U19135 (N_19135,N_18118,N_18995);
nand U19136 (N_19136,N_18551,N_18208);
nor U19137 (N_19137,N_18542,N_18575);
nor U19138 (N_19138,N_18872,N_18409);
or U19139 (N_19139,N_18536,N_18582);
or U19140 (N_19140,N_18401,N_18863);
nor U19141 (N_19141,N_18670,N_18799);
nor U19142 (N_19142,N_18241,N_18629);
xor U19143 (N_19143,N_18327,N_18263);
xnor U19144 (N_19144,N_18956,N_18725);
xnor U19145 (N_19145,N_18427,N_18234);
nand U19146 (N_19146,N_18961,N_18841);
and U19147 (N_19147,N_18832,N_18383);
nand U19148 (N_19148,N_18503,N_18751);
or U19149 (N_19149,N_18659,N_18920);
nor U19150 (N_19150,N_18204,N_18744);
nand U19151 (N_19151,N_18977,N_18755);
xnor U19152 (N_19152,N_18928,N_18869);
or U19153 (N_19153,N_18905,N_18280);
nor U19154 (N_19154,N_18157,N_18849);
xor U19155 (N_19155,N_18696,N_18798);
nand U19156 (N_19156,N_18379,N_18697);
nand U19157 (N_19157,N_18220,N_18792);
nand U19158 (N_19158,N_18201,N_18779);
nand U19159 (N_19159,N_18230,N_18734);
or U19160 (N_19160,N_18380,N_18353);
or U19161 (N_19161,N_18939,N_18399);
or U19162 (N_19162,N_18111,N_18191);
or U19163 (N_19163,N_18402,N_18660);
nor U19164 (N_19164,N_18347,N_18861);
nor U19165 (N_19165,N_18531,N_18174);
or U19166 (N_19166,N_18107,N_18051);
nor U19167 (N_19167,N_18212,N_18123);
xnor U19168 (N_19168,N_18227,N_18481);
nor U19169 (N_19169,N_18152,N_18494);
and U19170 (N_19170,N_18384,N_18970);
nor U19171 (N_19171,N_18901,N_18619);
nand U19172 (N_19172,N_18864,N_18298);
and U19173 (N_19173,N_18992,N_18447);
nor U19174 (N_19174,N_18462,N_18581);
nand U19175 (N_19175,N_18770,N_18237);
nand U19176 (N_19176,N_18532,N_18053);
or U19177 (N_19177,N_18255,N_18439);
nor U19178 (N_19178,N_18934,N_18281);
xnor U19179 (N_19179,N_18676,N_18830);
and U19180 (N_19180,N_18958,N_18024);
and U19181 (N_19181,N_18643,N_18880);
or U19182 (N_19182,N_18121,N_18076);
xor U19183 (N_19183,N_18311,N_18737);
or U19184 (N_19184,N_18615,N_18019);
xnor U19185 (N_19185,N_18068,N_18502);
nor U19186 (N_19186,N_18747,N_18617);
nor U19187 (N_19187,N_18012,N_18044);
nor U19188 (N_19188,N_18057,N_18205);
or U19189 (N_19189,N_18179,N_18370);
nand U19190 (N_19190,N_18296,N_18169);
nor U19191 (N_19191,N_18701,N_18766);
xnor U19192 (N_19192,N_18305,N_18001);
xnor U19193 (N_19193,N_18089,N_18671);
xor U19194 (N_19194,N_18543,N_18361);
nand U19195 (N_19195,N_18602,N_18440);
and U19196 (N_19196,N_18839,N_18858);
and U19197 (N_19197,N_18062,N_18906);
nor U19198 (N_19198,N_18936,N_18193);
and U19199 (N_19199,N_18276,N_18828);
xnor U19200 (N_19200,N_18871,N_18971);
and U19201 (N_19201,N_18546,N_18851);
xnor U19202 (N_19202,N_18325,N_18119);
nor U19203 (N_19203,N_18470,N_18594);
nor U19204 (N_19204,N_18002,N_18695);
and U19205 (N_19205,N_18576,N_18847);
nand U19206 (N_19206,N_18631,N_18054);
nor U19207 (N_19207,N_18393,N_18154);
xor U19208 (N_19208,N_18791,N_18785);
nand U19209 (N_19209,N_18730,N_18567);
nor U19210 (N_19210,N_18158,N_18020);
or U19211 (N_19211,N_18109,N_18039);
nand U19212 (N_19212,N_18413,N_18955);
or U19213 (N_19213,N_18598,N_18464);
and U19214 (N_19214,N_18490,N_18085);
xor U19215 (N_19215,N_18564,N_18915);
nand U19216 (N_19216,N_18166,N_18153);
or U19217 (N_19217,N_18222,N_18247);
and U19218 (N_19218,N_18291,N_18113);
nand U19219 (N_19219,N_18127,N_18810);
nand U19220 (N_19220,N_18181,N_18940);
or U19221 (N_19221,N_18508,N_18537);
or U19222 (N_19222,N_18246,N_18011);
and U19223 (N_19223,N_18329,N_18597);
and U19224 (N_19224,N_18213,N_18644);
nand U19225 (N_19225,N_18790,N_18450);
nor U19226 (N_19226,N_18163,N_18767);
nand U19227 (N_19227,N_18271,N_18634);
or U19228 (N_19228,N_18387,N_18870);
or U19229 (N_19229,N_18284,N_18937);
xnor U19230 (N_19230,N_18760,N_18831);
xnor U19231 (N_19231,N_18165,N_18382);
and U19232 (N_19232,N_18381,N_18590);
nand U19233 (N_19233,N_18930,N_18122);
xor U19234 (N_19234,N_18218,N_18507);
and U19235 (N_19235,N_18350,N_18804);
or U19236 (N_19236,N_18200,N_18789);
or U19237 (N_19237,N_18526,N_18330);
nand U19238 (N_19238,N_18859,N_18903);
nand U19239 (N_19239,N_18417,N_18762);
nor U19240 (N_19240,N_18434,N_18801);
nor U19241 (N_19241,N_18214,N_18095);
nand U19242 (N_19242,N_18922,N_18175);
and U19243 (N_19243,N_18726,N_18100);
and U19244 (N_19244,N_18515,N_18965);
and U19245 (N_19245,N_18500,N_18720);
or U19246 (N_19246,N_18886,N_18989);
or U19247 (N_19247,N_18151,N_18895);
nor U19248 (N_19248,N_18694,N_18684);
nand U19249 (N_19249,N_18455,N_18426);
or U19250 (N_19250,N_18446,N_18806);
xnor U19251 (N_19251,N_18484,N_18145);
nand U19252 (N_19252,N_18461,N_18261);
xnor U19253 (N_19253,N_18045,N_18638);
or U19254 (N_19254,N_18412,N_18358);
or U19255 (N_19255,N_18626,N_18714);
xnor U19256 (N_19256,N_18501,N_18279);
nand U19257 (N_19257,N_18188,N_18756);
nor U19258 (N_19258,N_18857,N_18463);
and U19259 (N_19259,N_18360,N_18290);
nand U19260 (N_19260,N_18084,N_18505);
nand U19261 (N_19261,N_18239,N_18835);
xnor U19262 (N_19262,N_18687,N_18004);
xnor U19263 (N_19263,N_18248,N_18033);
xor U19264 (N_19264,N_18368,N_18027);
and U19265 (N_19265,N_18953,N_18607);
xnor U19266 (N_19266,N_18112,N_18957);
nand U19267 (N_19267,N_18797,N_18608);
and U19268 (N_19268,N_18545,N_18881);
nor U19269 (N_19269,N_18672,N_18389);
xor U19270 (N_19270,N_18249,N_18245);
or U19271 (N_19271,N_18685,N_18823);
nand U19272 (N_19272,N_18207,N_18954);
and U19273 (N_19273,N_18448,N_18796);
nor U19274 (N_19274,N_18184,N_18818);
xnor U19275 (N_19275,N_18874,N_18528);
xor U19276 (N_19276,N_18674,N_18873);
nand U19277 (N_19277,N_18416,N_18487);
xor U19278 (N_19278,N_18794,N_18206);
xor U19279 (N_19279,N_18882,N_18194);
nor U19280 (N_19280,N_18663,N_18355);
and U19281 (N_19281,N_18739,N_18493);
nor U19282 (N_19282,N_18511,N_18233);
nor U19283 (N_19283,N_18574,N_18488);
nor U19284 (N_19284,N_18058,N_18553);
and U19285 (N_19285,N_18466,N_18326);
nand U19286 (N_19286,N_18034,N_18845);
nand U19287 (N_19287,N_18385,N_18229);
nor U19288 (N_19288,N_18623,N_18675);
nor U19289 (N_19289,N_18422,N_18645);
nor U19290 (N_19290,N_18398,N_18323);
or U19291 (N_19291,N_18260,N_18596);
and U19292 (N_19292,N_18506,N_18510);
xnor U19293 (N_19293,N_18023,N_18273);
nor U19294 (N_19294,N_18252,N_18764);
nor U19295 (N_19295,N_18717,N_18287);
xor U19296 (N_19296,N_18648,N_18666);
xor U19297 (N_19297,N_18622,N_18376);
nand U19298 (N_19298,N_18652,N_18825);
or U19299 (N_19299,N_18587,N_18319);
and U19300 (N_19300,N_18059,N_18550);
xor U19301 (N_19301,N_18253,N_18840);
nor U19302 (N_19302,N_18919,N_18431);
and U19303 (N_19303,N_18243,N_18816);
nand U19304 (N_19304,N_18041,N_18038);
nor U19305 (N_19305,N_18275,N_18877);
and U19306 (N_19306,N_18006,N_18254);
or U19307 (N_19307,N_18708,N_18952);
and U19308 (N_19308,N_18999,N_18110);
and U19309 (N_19309,N_18632,N_18539);
or U19310 (N_19310,N_18031,N_18354);
and U19311 (N_19311,N_18854,N_18593);
nand U19312 (N_19312,N_18140,N_18807);
and U19313 (N_19313,N_18314,N_18408);
and U19314 (N_19314,N_18657,N_18709);
and U19315 (N_19315,N_18975,N_18566);
and U19316 (N_19316,N_18702,N_18703);
nor U19317 (N_19317,N_18868,N_18026);
nor U19318 (N_19318,N_18554,N_18235);
and U19319 (N_19319,N_18884,N_18848);
nand U19320 (N_19320,N_18485,N_18458);
and U19321 (N_19321,N_18366,N_18719);
nor U19322 (N_19322,N_18588,N_18980);
xnor U19323 (N_19323,N_18265,N_18916);
nand U19324 (N_19324,N_18333,N_18172);
xor U19325 (N_19325,N_18056,N_18096);
nand U19326 (N_19326,N_18196,N_18927);
nand U19327 (N_19327,N_18173,N_18499);
nand U19328 (N_19328,N_18967,N_18844);
nor U19329 (N_19329,N_18074,N_18601);
xor U19330 (N_19330,N_18568,N_18342);
xnor U19331 (N_19331,N_18639,N_18178);
nand U19332 (N_19332,N_18236,N_18080);
and U19333 (N_19333,N_18713,N_18563);
nand U19334 (N_19334,N_18133,N_18143);
nand U19335 (N_19335,N_18357,N_18691);
xor U19336 (N_19336,N_18658,N_18750);
xnor U19337 (N_19337,N_18605,N_18017);
or U19338 (N_19338,N_18636,N_18555);
or U19339 (N_19339,N_18186,N_18929);
and U19340 (N_19340,N_18159,N_18761);
nor U19341 (N_19341,N_18407,N_18150);
or U19342 (N_19342,N_18438,N_18826);
and U19343 (N_19343,N_18996,N_18866);
nor U19344 (N_19344,N_18336,N_18187);
or U19345 (N_19345,N_18078,N_18699);
xor U19346 (N_19346,N_18099,N_18653);
xor U19347 (N_19347,N_18973,N_18374);
nand U19348 (N_19348,N_18673,N_18497);
nor U19349 (N_19349,N_18079,N_18094);
and U19350 (N_19350,N_18788,N_18561);
nor U19351 (N_19351,N_18707,N_18293);
and U19352 (N_19352,N_18520,N_18103);
nand U19353 (N_19353,N_18147,N_18073);
and U19354 (N_19354,N_18008,N_18815);
or U19355 (N_19355,N_18114,N_18969);
or U19356 (N_19356,N_18259,N_18479);
nor U19357 (N_19357,N_18324,N_18403);
and U19358 (N_19358,N_18917,N_18282);
nor U19359 (N_19359,N_18283,N_18050);
and U19360 (N_19360,N_18933,N_18949);
or U19361 (N_19361,N_18299,N_18689);
and U19362 (N_19362,N_18356,N_18449);
xnor U19363 (N_19363,N_18240,N_18359);
nand U19364 (N_19364,N_18394,N_18192);
nand U19365 (N_19365,N_18144,N_18538);
or U19366 (N_19366,N_18189,N_18396);
nand U19367 (N_19367,N_18469,N_18908);
or U19368 (N_19368,N_18979,N_18655);
or U19369 (N_19369,N_18573,N_18909);
xor U19370 (N_19370,N_18585,N_18170);
and U19371 (N_19371,N_18063,N_18432);
xnor U19372 (N_19372,N_18902,N_18215);
nand U19373 (N_19373,N_18897,N_18519);
nor U19374 (N_19374,N_18437,N_18932);
or U19375 (N_19375,N_18813,N_18410);
nor U19376 (N_19376,N_18735,N_18475);
nand U19377 (N_19377,N_18483,N_18941);
xnor U19378 (N_19378,N_18278,N_18473);
nor U19379 (N_19379,N_18527,N_18457);
and U19380 (N_19380,N_18262,N_18108);
and U19381 (N_19381,N_18128,N_18547);
nand U19382 (N_19382,N_18780,N_18040);
xor U19383 (N_19383,N_18388,N_18013);
xnor U19384 (N_19384,N_18976,N_18168);
xor U19385 (N_19385,N_18893,N_18300);
nand U19386 (N_19386,N_18264,N_18367);
nor U19387 (N_19387,N_18800,N_18925);
and U19388 (N_19388,N_18914,N_18746);
nor U19389 (N_19389,N_18724,N_18322);
nor U19390 (N_19390,N_18364,N_18183);
nand U19391 (N_19391,N_18981,N_18266);
and U19392 (N_19392,N_18086,N_18028);
and U19393 (N_19393,N_18517,N_18046);
nor U19394 (N_19394,N_18817,N_18754);
or U19395 (N_19395,N_18258,N_18693);
xnor U19396 (N_19396,N_18889,N_18787);
and U19397 (N_19397,N_18768,N_18297);
nor U19398 (N_19398,N_18729,N_18772);
nand U19399 (N_19399,N_18892,N_18343);
xnor U19400 (N_19400,N_18803,N_18966);
nand U19401 (N_19401,N_18087,N_18821);
nor U19402 (N_19402,N_18295,N_18048);
nor U19403 (N_19403,N_18938,N_18351);
and U19404 (N_19404,N_18710,N_18468);
xnor U19405 (N_19405,N_18984,N_18838);
nor U19406 (N_19406,N_18513,N_18405);
nor U19407 (N_19407,N_18795,N_18647);
nand U19408 (N_19408,N_18738,N_18226);
xnor U19409 (N_19409,N_18406,N_18459);
nor U19410 (N_19410,N_18312,N_18139);
and U19411 (N_19411,N_18365,N_18244);
nor U19412 (N_19412,N_18662,N_18190);
nand U19413 (N_19413,N_18126,N_18963);
nand U19414 (N_19414,N_18512,N_18879);
xnor U19415 (N_19415,N_18492,N_18269);
or U19416 (N_19416,N_18137,N_18668);
nand U19417 (N_19417,N_18372,N_18924);
xor U19418 (N_19418,N_18436,N_18637);
nor U19419 (N_19419,N_18824,N_18009);
or U19420 (N_19420,N_18124,N_18819);
or U19421 (N_19421,N_18042,N_18583);
nor U19422 (N_19422,N_18987,N_18748);
xor U19423 (N_19423,N_18171,N_18160);
and U19424 (N_19424,N_18572,N_18964);
and U19425 (N_19425,N_18395,N_18621);
nor U19426 (N_19426,N_18682,N_18876);
nand U19427 (N_19427,N_18091,N_18415);
nand U19428 (N_19428,N_18669,N_18524);
or U19429 (N_19429,N_18728,N_18016);
nand U19430 (N_19430,N_18752,N_18070);
or U19431 (N_19431,N_18288,N_18778);
nor U19432 (N_19432,N_18397,N_18610);
nand U19433 (N_19433,N_18640,N_18098);
xnor U19434 (N_19434,N_18197,N_18820);
and U19435 (N_19435,N_18777,N_18313);
xnor U19436 (N_19436,N_18586,N_18910);
and U19437 (N_19437,N_18518,N_18082);
xor U19438 (N_19438,N_18565,N_18891);
xnor U19439 (N_19439,N_18474,N_18467);
nand U19440 (N_19440,N_18180,N_18067);
and U19441 (N_19441,N_18900,N_18883);
nand U19442 (N_19442,N_18935,N_18654);
or U19443 (N_19443,N_18301,N_18292);
and U19444 (N_19444,N_18117,N_18856);
nor U19445 (N_19445,N_18742,N_18757);
nor U19446 (N_19446,N_18661,N_18134);
or U19447 (N_19447,N_18557,N_18132);
nand U19448 (N_19448,N_18556,N_18811);
nor U19449 (N_19449,N_18341,N_18646);
or U19450 (N_19450,N_18951,N_18307);
nor U19451 (N_19451,N_18176,N_18990);
xor U19452 (N_19452,N_18014,N_18852);
and U19453 (N_19453,N_18477,N_18375);
xnor U19454 (N_19454,N_18482,N_18486);
nor U19455 (N_19455,N_18344,N_18945);
nor U19456 (N_19456,N_18853,N_18667);
nor U19457 (N_19457,N_18769,N_18948);
nand U19458 (N_19458,N_18904,N_18783);
or U19459 (N_19459,N_18456,N_18005);
nand U19460 (N_19460,N_18926,N_18423);
nand U19461 (N_19461,N_18968,N_18472);
xnor U19462 (N_19462,N_18721,N_18913);
nand U19463 (N_19463,N_18286,N_18097);
nor U19464 (N_19464,N_18771,N_18430);
nor U19465 (N_19465,N_18616,N_18065);
and U19466 (N_19466,N_18731,N_18759);
xor U19467 (N_19467,N_18060,N_18105);
or U19468 (N_19468,N_18267,N_18277);
or U19469 (N_19469,N_18451,N_18833);
nand U19470 (N_19470,N_18603,N_18578);
and U19471 (N_19471,N_18680,N_18064);
or U19472 (N_19472,N_18773,N_18982);
nand U19473 (N_19473,N_18525,N_18274);
xor U19474 (N_19474,N_18885,N_18442);
xor U19475 (N_19475,N_18947,N_18843);
and U19476 (N_19476,N_18043,N_18072);
and U19477 (N_19477,N_18125,N_18077);
nor U19478 (N_19478,N_18471,N_18225);
nand U19479 (N_19479,N_18115,N_18782);
nand U19480 (N_19480,N_18558,N_18604);
or U19481 (N_19481,N_18424,N_18377);
or U19482 (N_19482,N_18480,N_18591);
xor U19483 (N_19483,N_18390,N_18441);
xnor U19484 (N_19484,N_18733,N_18878);
or U19485 (N_19485,N_18136,N_18959);
xor U19486 (N_19486,N_18348,N_18460);
nand U19487 (N_19487,N_18185,N_18444);
nor U19488 (N_19488,N_18289,N_18088);
and U19489 (N_19489,N_18704,N_18420);
and U19490 (N_19490,N_18888,N_18774);
or U19491 (N_19491,N_18029,N_18036);
or U19492 (N_19492,N_18421,N_18822);
nand U19493 (N_19493,N_18912,N_18842);
nand U19494 (N_19494,N_18698,N_18549);
nand U19495 (N_19495,N_18887,N_18362);
nand U19496 (N_19496,N_18559,N_18478);
or U19497 (N_19497,N_18003,N_18718);
and U19498 (N_19498,N_18335,N_18749);
nand U19499 (N_19499,N_18624,N_18216);
nor U19500 (N_19500,N_18280,N_18384);
or U19501 (N_19501,N_18101,N_18459);
and U19502 (N_19502,N_18922,N_18782);
or U19503 (N_19503,N_18990,N_18328);
nor U19504 (N_19504,N_18629,N_18881);
and U19505 (N_19505,N_18264,N_18678);
and U19506 (N_19506,N_18931,N_18171);
nand U19507 (N_19507,N_18641,N_18293);
or U19508 (N_19508,N_18071,N_18304);
nor U19509 (N_19509,N_18961,N_18460);
or U19510 (N_19510,N_18716,N_18238);
xor U19511 (N_19511,N_18030,N_18065);
and U19512 (N_19512,N_18115,N_18799);
nor U19513 (N_19513,N_18005,N_18321);
and U19514 (N_19514,N_18169,N_18686);
nand U19515 (N_19515,N_18760,N_18355);
or U19516 (N_19516,N_18789,N_18029);
nor U19517 (N_19517,N_18599,N_18468);
xor U19518 (N_19518,N_18058,N_18398);
nand U19519 (N_19519,N_18834,N_18228);
or U19520 (N_19520,N_18277,N_18314);
and U19521 (N_19521,N_18571,N_18170);
nor U19522 (N_19522,N_18947,N_18719);
or U19523 (N_19523,N_18766,N_18854);
xnor U19524 (N_19524,N_18896,N_18199);
xnor U19525 (N_19525,N_18246,N_18774);
and U19526 (N_19526,N_18041,N_18961);
nand U19527 (N_19527,N_18019,N_18025);
and U19528 (N_19528,N_18997,N_18828);
and U19529 (N_19529,N_18717,N_18147);
xnor U19530 (N_19530,N_18681,N_18521);
or U19531 (N_19531,N_18966,N_18101);
xor U19532 (N_19532,N_18766,N_18483);
or U19533 (N_19533,N_18823,N_18771);
and U19534 (N_19534,N_18409,N_18703);
and U19535 (N_19535,N_18891,N_18381);
xnor U19536 (N_19536,N_18472,N_18204);
or U19537 (N_19537,N_18830,N_18173);
or U19538 (N_19538,N_18881,N_18791);
xor U19539 (N_19539,N_18761,N_18634);
or U19540 (N_19540,N_18835,N_18773);
nand U19541 (N_19541,N_18643,N_18885);
nand U19542 (N_19542,N_18029,N_18157);
nand U19543 (N_19543,N_18528,N_18493);
and U19544 (N_19544,N_18354,N_18715);
nor U19545 (N_19545,N_18254,N_18201);
nand U19546 (N_19546,N_18604,N_18411);
nand U19547 (N_19547,N_18758,N_18685);
nor U19548 (N_19548,N_18710,N_18813);
xnor U19549 (N_19549,N_18861,N_18823);
and U19550 (N_19550,N_18602,N_18366);
nand U19551 (N_19551,N_18987,N_18623);
nand U19552 (N_19552,N_18840,N_18665);
nor U19553 (N_19553,N_18246,N_18271);
and U19554 (N_19554,N_18129,N_18403);
and U19555 (N_19555,N_18050,N_18354);
nor U19556 (N_19556,N_18865,N_18296);
nand U19557 (N_19557,N_18873,N_18048);
nor U19558 (N_19558,N_18438,N_18055);
nor U19559 (N_19559,N_18971,N_18472);
or U19560 (N_19560,N_18327,N_18824);
xnor U19561 (N_19561,N_18887,N_18738);
xnor U19562 (N_19562,N_18546,N_18970);
or U19563 (N_19563,N_18802,N_18302);
or U19564 (N_19564,N_18778,N_18798);
and U19565 (N_19565,N_18536,N_18510);
nand U19566 (N_19566,N_18680,N_18496);
nor U19567 (N_19567,N_18162,N_18777);
or U19568 (N_19568,N_18530,N_18408);
nor U19569 (N_19569,N_18757,N_18722);
nor U19570 (N_19570,N_18823,N_18637);
xor U19571 (N_19571,N_18626,N_18837);
nor U19572 (N_19572,N_18641,N_18831);
nand U19573 (N_19573,N_18923,N_18693);
nand U19574 (N_19574,N_18369,N_18110);
xor U19575 (N_19575,N_18501,N_18171);
nor U19576 (N_19576,N_18724,N_18096);
and U19577 (N_19577,N_18713,N_18362);
nor U19578 (N_19578,N_18152,N_18135);
or U19579 (N_19579,N_18036,N_18480);
or U19580 (N_19580,N_18856,N_18497);
and U19581 (N_19581,N_18746,N_18100);
nor U19582 (N_19582,N_18170,N_18338);
or U19583 (N_19583,N_18060,N_18458);
xor U19584 (N_19584,N_18347,N_18785);
nand U19585 (N_19585,N_18266,N_18885);
or U19586 (N_19586,N_18259,N_18694);
xnor U19587 (N_19587,N_18566,N_18838);
nor U19588 (N_19588,N_18787,N_18840);
nor U19589 (N_19589,N_18185,N_18976);
or U19590 (N_19590,N_18844,N_18914);
nand U19591 (N_19591,N_18424,N_18912);
nor U19592 (N_19592,N_18865,N_18864);
and U19593 (N_19593,N_18668,N_18244);
nor U19594 (N_19594,N_18105,N_18750);
or U19595 (N_19595,N_18697,N_18642);
and U19596 (N_19596,N_18279,N_18825);
nor U19597 (N_19597,N_18153,N_18971);
nand U19598 (N_19598,N_18029,N_18264);
and U19599 (N_19599,N_18525,N_18260);
nand U19600 (N_19600,N_18366,N_18626);
nor U19601 (N_19601,N_18814,N_18217);
nand U19602 (N_19602,N_18193,N_18132);
and U19603 (N_19603,N_18440,N_18000);
nor U19604 (N_19604,N_18694,N_18716);
nor U19605 (N_19605,N_18468,N_18512);
xor U19606 (N_19606,N_18551,N_18108);
and U19607 (N_19607,N_18745,N_18669);
and U19608 (N_19608,N_18698,N_18865);
and U19609 (N_19609,N_18331,N_18909);
nor U19610 (N_19610,N_18972,N_18954);
xnor U19611 (N_19611,N_18123,N_18845);
or U19612 (N_19612,N_18899,N_18755);
xor U19613 (N_19613,N_18235,N_18798);
nor U19614 (N_19614,N_18175,N_18143);
nand U19615 (N_19615,N_18228,N_18012);
and U19616 (N_19616,N_18511,N_18479);
and U19617 (N_19617,N_18051,N_18080);
or U19618 (N_19618,N_18139,N_18707);
nand U19619 (N_19619,N_18757,N_18645);
nand U19620 (N_19620,N_18611,N_18694);
nand U19621 (N_19621,N_18297,N_18945);
and U19622 (N_19622,N_18712,N_18957);
nand U19623 (N_19623,N_18925,N_18517);
or U19624 (N_19624,N_18254,N_18716);
and U19625 (N_19625,N_18590,N_18961);
nor U19626 (N_19626,N_18957,N_18326);
xor U19627 (N_19627,N_18603,N_18407);
xnor U19628 (N_19628,N_18992,N_18379);
nand U19629 (N_19629,N_18952,N_18428);
or U19630 (N_19630,N_18888,N_18213);
or U19631 (N_19631,N_18664,N_18432);
and U19632 (N_19632,N_18040,N_18238);
and U19633 (N_19633,N_18353,N_18406);
or U19634 (N_19634,N_18115,N_18867);
or U19635 (N_19635,N_18557,N_18971);
nor U19636 (N_19636,N_18247,N_18142);
xor U19637 (N_19637,N_18418,N_18816);
nand U19638 (N_19638,N_18294,N_18505);
or U19639 (N_19639,N_18951,N_18641);
or U19640 (N_19640,N_18848,N_18114);
xnor U19641 (N_19641,N_18535,N_18456);
and U19642 (N_19642,N_18345,N_18410);
nand U19643 (N_19643,N_18312,N_18047);
or U19644 (N_19644,N_18739,N_18190);
nand U19645 (N_19645,N_18114,N_18705);
nor U19646 (N_19646,N_18271,N_18036);
xnor U19647 (N_19647,N_18950,N_18982);
xnor U19648 (N_19648,N_18548,N_18852);
nor U19649 (N_19649,N_18522,N_18249);
nand U19650 (N_19650,N_18319,N_18795);
or U19651 (N_19651,N_18317,N_18470);
or U19652 (N_19652,N_18325,N_18288);
xor U19653 (N_19653,N_18752,N_18728);
nor U19654 (N_19654,N_18631,N_18721);
xor U19655 (N_19655,N_18470,N_18137);
xnor U19656 (N_19656,N_18869,N_18770);
xnor U19657 (N_19657,N_18475,N_18702);
nand U19658 (N_19658,N_18402,N_18913);
nand U19659 (N_19659,N_18795,N_18295);
xor U19660 (N_19660,N_18078,N_18362);
xor U19661 (N_19661,N_18698,N_18044);
and U19662 (N_19662,N_18018,N_18268);
nand U19663 (N_19663,N_18082,N_18344);
nand U19664 (N_19664,N_18611,N_18303);
xnor U19665 (N_19665,N_18553,N_18839);
and U19666 (N_19666,N_18397,N_18993);
xor U19667 (N_19667,N_18894,N_18746);
nand U19668 (N_19668,N_18227,N_18048);
nor U19669 (N_19669,N_18106,N_18009);
and U19670 (N_19670,N_18612,N_18954);
and U19671 (N_19671,N_18984,N_18005);
and U19672 (N_19672,N_18865,N_18143);
nand U19673 (N_19673,N_18658,N_18703);
nand U19674 (N_19674,N_18035,N_18232);
nand U19675 (N_19675,N_18436,N_18373);
or U19676 (N_19676,N_18778,N_18875);
or U19677 (N_19677,N_18473,N_18270);
nand U19678 (N_19678,N_18490,N_18156);
nor U19679 (N_19679,N_18273,N_18645);
nand U19680 (N_19680,N_18332,N_18453);
and U19681 (N_19681,N_18881,N_18753);
nor U19682 (N_19682,N_18674,N_18756);
nor U19683 (N_19683,N_18776,N_18027);
and U19684 (N_19684,N_18723,N_18357);
nor U19685 (N_19685,N_18123,N_18691);
nor U19686 (N_19686,N_18554,N_18603);
or U19687 (N_19687,N_18961,N_18297);
and U19688 (N_19688,N_18437,N_18951);
or U19689 (N_19689,N_18388,N_18425);
nand U19690 (N_19690,N_18837,N_18983);
and U19691 (N_19691,N_18429,N_18527);
or U19692 (N_19692,N_18838,N_18948);
xnor U19693 (N_19693,N_18076,N_18012);
nand U19694 (N_19694,N_18050,N_18015);
nand U19695 (N_19695,N_18282,N_18747);
or U19696 (N_19696,N_18652,N_18962);
nor U19697 (N_19697,N_18671,N_18696);
or U19698 (N_19698,N_18923,N_18995);
nand U19699 (N_19699,N_18064,N_18565);
nand U19700 (N_19700,N_18500,N_18707);
and U19701 (N_19701,N_18950,N_18118);
nor U19702 (N_19702,N_18381,N_18909);
and U19703 (N_19703,N_18727,N_18805);
nor U19704 (N_19704,N_18314,N_18885);
and U19705 (N_19705,N_18623,N_18887);
xnor U19706 (N_19706,N_18490,N_18946);
xor U19707 (N_19707,N_18364,N_18606);
nand U19708 (N_19708,N_18505,N_18840);
and U19709 (N_19709,N_18113,N_18901);
xor U19710 (N_19710,N_18289,N_18435);
nor U19711 (N_19711,N_18586,N_18960);
nand U19712 (N_19712,N_18000,N_18718);
or U19713 (N_19713,N_18217,N_18704);
nand U19714 (N_19714,N_18172,N_18331);
and U19715 (N_19715,N_18456,N_18395);
and U19716 (N_19716,N_18445,N_18360);
xnor U19717 (N_19717,N_18703,N_18914);
xnor U19718 (N_19718,N_18085,N_18890);
nand U19719 (N_19719,N_18527,N_18573);
nor U19720 (N_19720,N_18026,N_18312);
xor U19721 (N_19721,N_18558,N_18192);
and U19722 (N_19722,N_18470,N_18158);
nand U19723 (N_19723,N_18838,N_18603);
or U19724 (N_19724,N_18314,N_18946);
or U19725 (N_19725,N_18989,N_18399);
nand U19726 (N_19726,N_18667,N_18808);
xor U19727 (N_19727,N_18895,N_18302);
nor U19728 (N_19728,N_18679,N_18688);
xnor U19729 (N_19729,N_18237,N_18687);
and U19730 (N_19730,N_18136,N_18331);
xor U19731 (N_19731,N_18928,N_18186);
and U19732 (N_19732,N_18535,N_18622);
or U19733 (N_19733,N_18548,N_18673);
xor U19734 (N_19734,N_18150,N_18551);
and U19735 (N_19735,N_18946,N_18585);
xnor U19736 (N_19736,N_18206,N_18061);
xor U19737 (N_19737,N_18380,N_18337);
and U19738 (N_19738,N_18223,N_18463);
nand U19739 (N_19739,N_18270,N_18315);
and U19740 (N_19740,N_18436,N_18320);
xor U19741 (N_19741,N_18006,N_18644);
or U19742 (N_19742,N_18486,N_18862);
or U19743 (N_19743,N_18062,N_18510);
nand U19744 (N_19744,N_18706,N_18655);
nand U19745 (N_19745,N_18249,N_18311);
and U19746 (N_19746,N_18489,N_18603);
or U19747 (N_19747,N_18443,N_18149);
nand U19748 (N_19748,N_18460,N_18929);
and U19749 (N_19749,N_18141,N_18239);
and U19750 (N_19750,N_18231,N_18135);
or U19751 (N_19751,N_18777,N_18930);
nand U19752 (N_19752,N_18411,N_18263);
xnor U19753 (N_19753,N_18247,N_18174);
nand U19754 (N_19754,N_18796,N_18820);
and U19755 (N_19755,N_18270,N_18025);
xor U19756 (N_19756,N_18302,N_18070);
or U19757 (N_19757,N_18962,N_18248);
nand U19758 (N_19758,N_18016,N_18525);
nand U19759 (N_19759,N_18664,N_18018);
nor U19760 (N_19760,N_18580,N_18056);
nor U19761 (N_19761,N_18106,N_18785);
nor U19762 (N_19762,N_18841,N_18586);
or U19763 (N_19763,N_18151,N_18516);
xnor U19764 (N_19764,N_18708,N_18768);
and U19765 (N_19765,N_18750,N_18034);
or U19766 (N_19766,N_18218,N_18789);
nor U19767 (N_19767,N_18107,N_18313);
nand U19768 (N_19768,N_18987,N_18519);
xor U19769 (N_19769,N_18704,N_18233);
xor U19770 (N_19770,N_18946,N_18227);
or U19771 (N_19771,N_18661,N_18261);
or U19772 (N_19772,N_18144,N_18894);
nand U19773 (N_19773,N_18356,N_18234);
or U19774 (N_19774,N_18986,N_18728);
xnor U19775 (N_19775,N_18290,N_18915);
nor U19776 (N_19776,N_18862,N_18510);
and U19777 (N_19777,N_18808,N_18294);
nand U19778 (N_19778,N_18722,N_18503);
nand U19779 (N_19779,N_18491,N_18977);
nand U19780 (N_19780,N_18434,N_18749);
or U19781 (N_19781,N_18803,N_18101);
xor U19782 (N_19782,N_18232,N_18475);
nand U19783 (N_19783,N_18058,N_18633);
xor U19784 (N_19784,N_18058,N_18434);
or U19785 (N_19785,N_18674,N_18690);
nand U19786 (N_19786,N_18546,N_18442);
nand U19787 (N_19787,N_18100,N_18072);
or U19788 (N_19788,N_18459,N_18217);
or U19789 (N_19789,N_18511,N_18022);
and U19790 (N_19790,N_18077,N_18235);
nor U19791 (N_19791,N_18518,N_18585);
nand U19792 (N_19792,N_18274,N_18146);
xor U19793 (N_19793,N_18548,N_18306);
nand U19794 (N_19794,N_18578,N_18777);
xnor U19795 (N_19795,N_18932,N_18661);
nand U19796 (N_19796,N_18594,N_18537);
nor U19797 (N_19797,N_18104,N_18274);
or U19798 (N_19798,N_18470,N_18001);
nand U19799 (N_19799,N_18672,N_18100);
and U19800 (N_19800,N_18267,N_18093);
xor U19801 (N_19801,N_18502,N_18050);
xnor U19802 (N_19802,N_18552,N_18798);
and U19803 (N_19803,N_18729,N_18937);
or U19804 (N_19804,N_18642,N_18667);
xnor U19805 (N_19805,N_18142,N_18316);
or U19806 (N_19806,N_18355,N_18672);
nand U19807 (N_19807,N_18857,N_18881);
nand U19808 (N_19808,N_18804,N_18954);
and U19809 (N_19809,N_18793,N_18837);
and U19810 (N_19810,N_18265,N_18154);
nand U19811 (N_19811,N_18861,N_18827);
nor U19812 (N_19812,N_18588,N_18415);
or U19813 (N_19813,N_18864,N_18288);
nor U19814 (N_19814,N_18899,N_18692);
and U19815 (N_19815,N_18791,N_18685);
xor U19816 (N_19816,N_18720,N_18470);
or U19817 (N_19817,N_18761,N_18807);
and U19818 (N_19818,N_18763,N_18127);
nand U19819 (N_19819,N_18622,N_18776);
xor U19820 (N_19820,N_18392,N_18713);
or U19821 (N_19821,N_18086,N_18841);
nor U19822 (N_19822,N_18108,N_18805);
or U19823 (N_19823,N_18100,N_18386);
xnor U19824 (N_19824,N_18638,N_18068);
xor U19825 (N_19825,N_18840,N_18085);
nor U19826 (N_19826,N_18194,N_18445);
xnor U19827 (N_19827,N_18910,N_18555);
nor U19828 (N_19828,N_18764,N_18584);
or U19829 (N_19829,N_18691,N_18361);
xnor U19830 (N_19830,N_18008,N_18740);
or U19831 (N_19831,N_18011,N_18515);
nor U19832 (N_19832,N_18232,N_18240);
nor U19833 (N_19833,N_18231,N_18719);
or U19834 (N_19834,N_18754,N_18914);
xnor U19835 (N_19835,N_18529,N_18230);
nor U19836 (N_19836,N_18068,N_18618);
nor U19837 (N_19837,N_18689,N_18887);
or U19838 (N_19838,N_18138,N_18063);
nand U19839 (N_19839,N_18350,N_18237);
and U19840 (N_19840,N_18628,N_18863);
or U19841 (N_19841,N_18808,N_18483);
xor U19842 (N_19842,N_18440,N_18459);
and U19843 (N_19843,N_18775,N_18690);
nor U19844 (N_19844,N_18274,N_18931);
nand U19845 (N_19845,N_18381,N_18897);
xor U19846 (N_19846,N_18428,N_18827);
or U19847 (N_19847,N_18724,N_18704);
and U19848 (N_19848,N_18716,N_18728);
nor U19849 (N_19849,N_18887,N_18815);
xnor U19850 (N_19850,N_18459,N_18358);
nor U19851 (N_19851,N_18075,N_18032);
or U19852 (N_19852,N_18245,N_18995);
and U19853 (N_19853,N_18530,N_18927);
nand U19854 (N_19854,N_18971,N_18690);
nand U19855 (N_19855,N_18477,N_18459);
nand U19856 (N_19856,N_18041,N_18328);
and U19857 (N_19857,N_18341,N_18439);
nand U19858 (N_19858,N_18950,N_18169);
or U19859 (N_19859,N_18569,N_18264);
nand U19860 (N_19860,N_18086,N_18982);
nor U19861 (N_19861,N_18870,N_18750);
nand U19862 (N_19862,N_18300,N_18764);
xor U19863 (N_19863,N_18511,N_18590);
or U19864 (N_19864,N_18733,N_18672);
or U19865 (N_19865,N_18370,N_18235);
xor U19866 (N_19866,N_18269,N_18082);
nor U19867 (N_19867,N_18091,N_18012);
and U19868 (N_19868,N_18648,N_18036);
or U19869 (N_19869,N_18289,N_18237);
xnor U19870 (N_19870,N_18125,N_18615);
xor U19871 (N_19871,N_18514,N_18511);
xnor U19872 (N_19872,N_18066,N_18714);
and U19873 (N_19873,N_18126,N_18326);
xor U19874 (N_19874,N_18746,N_18915);
or U19875 (N_19875,N_18692,N_18032);
xnor U19876 (N_19876,N_18115,N_18234);
nand U19877 (N_19877,N_18234,N_18766);
nor U19878 (N_19878,N_18328,N_18370);
and U19879 (N_19879,N_18263,N_18136);
xor U19880 (N_19880,N_18115,N_18143);
or U19881 (N_19881,N_18008,N_18060);
or U19882 (N_19882,N_18866,N_18836);
and U19883 (N_19883,N_18643,N_18053);
nand U19884 (N_19884,N_18478,N_18536);
nor U19885 (N_19885,N_18868,N_18656);
or U19886 (N_19886,N_18592,N_18704);
nand U19887 (N_19887,N_18307,N_18927);
and U19888 (N_19888,N_18702,N_18040);
nor U19889 (N_19889,N_18676,N_18163);
or U19890 (N_19890,N_18459,N_18768);
nor U19891 (N_19891,N_18836,N_18864);
nand U19892 (N_19892,N_18231,N_18671);
and U19893 (N_19893,N_18059,N_18922);
nand U19894 (N_19894,N_18072,N_18825);
and U19895 (N_19895,N_18321,N_18547);
or U19896 (N_19896,N_18883,N_18458);
nand U19897 (N_19897,N_18561,N_18402);
nand U19898 (N_19898,N_18696,N_18191);
xnor U19899 (N_19899,N_18810,N_18608);
nand U19900 (N_19900,N_18337,N_18799);
nor U19901 (N_19901,N_18818,N_18680);
nand U19902 (N_19902,N_18980,N_18665);
nor U19903 (N_19903,N_18583,N_18684);
nor U19904 (N_19904,N_18525,N_18701);
nor U19905 (N_19905,N_18620,N_18278);
nand U19906 (N_19906,N_18521,N_18236);
xnor U19907 (N_19907,N_18350,N_18412);
or U19908 (N_19908,N_18249,N_18616);
xor U19909 (N_19909,N_18925,N_18043);
nor U19910 (N_19910,N_18241,N_18556);
nand U19911 (N_19911,N_18450,N_18156);
and U19912 (N_19912,N_18322,N_18666);
nand U19913 (N_19913,N_18112,N_18140);
nor U19914 (N_19914,N_18124,N_18964);
or U19915 (N_19915,N_18370,N_18623);
nand U19916 (N_19916,N_18793,N_18708);
or U19917 (N_19917,N_18460,N_18201);
xnor U19918 (N_19918,N_18725,N_18443);
and U19919 (N_19919,N_18395,N_18872);
xnor U19920 (N_19920,N_18918,N_18862);
or U19921 (N_19921,N_18275,N_18097);
nand U19922 (N_19922,N_18404,N_18663);
nand U19923 (N_19923,N_18621,N_18873);
and U19924 (N_19924,N_18070,N_18607);
nor U19925 (N_19925,N_18507,N_18153);
and U19926 (N_19926,N_18485,N_18621);
or U19927 (N_19927,N_18166,N_18407);
xnor U19928 (N_19928,N_18053,N_18727);
or U19929 (N_19929,N_18313,N_18631);
xor U19930 (N_19930,N_18005,N_18636);
nor U19931 (N_19931,N_18107,N_18293);
nand U19932 (N_19932,N_18121,N_18707);
xnor U19933 (N_19933,N_18162,N_18127);
or U19934 (N_19934,N_18126,N_18585);
xor U19935 (N_19935,N_18303,N_18095);
or U19936 (N_19936,N_18371,N_18338);
xnor U19937 (N_19937,N_18221,N_18108);
or U19938 (N_19938,N_18955,N_18706);
and U19939 (N_19939,N_18292,N_18598);
xor U19940 (N_19940,N_18707,N_18769);
or U19941 (N_19941,N_18742,N_18799);
nand U19942 (N_19942,N_18867,N_18227);
xor U19943 (N_19943,N_18082,N_18101);
nor U19944 (N_19944,N_18179,N_18151);
and U19945 (N_19945,N_18906,N_18353);
and U19946 (N_19946,N_18189,N_18154);
nand U19947 (N_19947,N_18254,N_18188);
or U19948 (N_19948,N_18779,N_18362);
and U19949 (N_19949,N_18938,N_18638);
xnor U19950 (N_19950,N_18912,N_18759);
nor U19951 (N_19951,N_18674,N_18820);
xnor U19952 (N_19952,N_18919,N_18466);
nand U19953 (N_19953,N_18088,N_18449);
and U19954 (N_19954,N_18704,N_18481);
nand U19955 (N_19955,N_18215,N_18571);
nor U19956 (N_19956,N_18064,N_18262);
and U19957 (N_19957,N_18323,N_18583);
nor U19958 (N_19958,N_18937,N_18588);
xor U19959 (N_19959,N_18521,N_18573);
and U19960 (N_19960,N_18481,N_18520);
nand U19961 (N_19961,N_18903,N_18502);
xnor U19962 (N_19962,N_18548,N_18117);
nand U19963 (N_19963,N_18830,N_18997);
or U19964 (N_19964,N_18232,N_18335);
and U19965 (N_19965,N_18700,N_18188);
or U19966 (N_19966,N_18064,N_18308);
or U19967 (N_19967,N_18743,N_18112);
nor U19968 (N_19968,N_18061,N_18001);
nor U19969 (N_19969,N_18294,N_18059);
nand U19970 (N_19970,N_18912,N_18749);
nor U19971 (N_19971,N_18559,N_18443);
and U19972 (N_19972,N_18498,N_18371);
and U19973 (N_19973,N_18693,N_18909);
nand U19974 (N_19974,N_18669,N_18866);
nand U19975 (N_19975,N_18995,N_18563);
or U19976 (N_19976,N_18615,N_18560);
or U19977 (N_19977,N_18242,N_18666);
nand U19978 (N_19978,N_18160,N_18550);
and U19979 (N_19979,N_18678,N_18253);
xnor U19980 (N_19980,N_18557,N_18920);
nand U19981 (N_19981,N_18813,N_18584);
and U19982 (N_19982,N_18299,N_18010);
or U19983 (N_19983,N_18650,N_18483);
nor U19984 (N_19984,N_18367,N_18104);
nand U19985 (N_19985,N_18954,N_18608);
or U19986 (N_19986,N_18218,N_18637);
nor U19987 (N_19987,N_18414,N_18844);
or U19988 (N_19988,N_18706,N_18880);
xor U19989 (N_19989,N_18043,N_18803);
or U19990 (N_19990,N_18231,N_18466);
and U19991 (N_19991,N_18714,N_18267);
nor U19992 (N_19992,N_18916,N_18793);
or U19993 (N_19993,N_18260,N_18644);
nor U19994 (N_19994,N_18906,N_18044);
nand U19995 (N_19995,N_18624,N_18283);
nor U19996 (N_19996,N_18726,N_18453);
xor U19997 (N_19997,N_18472,N_18489);
and U19998 (N_19998,N_18922,N_18912);
nor U19999 (N_19999,N_18978,N_18077);
or U20000 (N_20000,N_19664,N_19018);
nand U20001 (N_20001,N_19537,N_19007);
xnor U20002 (N_20002,N_19413,N_19347);
nor U20003 (N_20003,N_19375,N_19732);
nand U20004 (N_20004,N_19709,N_19948);
nor U20005 (N_20005,N_19695,N_19051);
xor U20006 (N_20006,N_19860,N_19882);
and U20007 (N_20007,N_19898,N_19974);
xor U20008 (N_20008,N_19570,N_19735);
nor U20009 (N_20009,N_19660,N_19901);
xor U20010 (N_20010,N_19779,N_19435);
and U20011 (N_20011,N_19543,N_19834);
xnor U20012 (N_20012,N_19149,N_19061);
or U20013 (N_20013,N_19278,N_19135);
nor U20014 (N_20014,N_19497,N_19981);
and U20015 (N_20015,N_19717,N_19388);
nand U20016 (N_20016,N_19158,N_19801);
or U20017 (N_20017,N_19271,N_19701);
or U20018 (N_20018,N_19270,N_19358);
and U20019 (N_20019,N_19304,N_19799);
or U20020 (N_20020,N_19085,N_19219);
nand U20021 (N_20021,N_19505,N_19551);
xor U20022 (N_20022,N_19708,N_19392);
nor U20023 (N_20023,N_19019,N_19675);
and U20024 (N_20024,N_19218,N_19386);
xor U20025 (N_20025,N_19819,N_19476);
xor U20026 (N_20026,N_19595,N_19105);
or U20027 (N_20027,N_19596,N_19716);
nand U20028 (N_20028,N_19071,N_19142);
nand U20029 (N_20029,N_19953,N_19743);
or U20030 (N_20030,N_19482,N_19858);
xnor U20031 (N_20031,N_19054,N_19305);
nor U20032 (N_20032,N_19024,N_19616);
nor U20033 (N_20033,N_19780,N_19557);
nand U20034 (N_20034,N_19726,N_19609);
or U20035 (N_20035,N_19035,N_19066);
or U20036 (N_20036,N_19839,N_19907);
and U20037 (N_20037,N_19844,N_19873);
xnor U20038 (N_20038,N_19196,N_19913);
or U20039 (N_20039,N_19324,N_19266);
nor U20040 (N_20040,N_19074,N_19892);
xnor U20041 (N_20041,N_19242,N_19564);
nor U20042 (N_20042,N_19666,N_19849);
nand U20043 (N_20043,N_19740,N_19669);
xnor U20044 (N_20044,N_19684,N_19925);
and U20045 (N_20045,N_19467,N_19513);
nor U20046 (N_20046,N_19836,N_19311);
or U20047 (N_20047,N_19191,N_19177);
nand U20048 (N_20048,N_19460,N_19725);
and U20049 (N_20049,N_19759,N_19887);
xor U20050 (N_20050,N_19453,N_19996);
xor U20051 (N_20051,N_19113,N_19472);
and U20052 (N_20052,N_19417,N_19714);
and U20053 (N_20053,N_19079,N_19976);
nand U20054 (N_20054,N_19603,N_19293);
nor U20055 (N_20055,N_19313,N_19621);
and U20056 (N_20056,N_19397,N_19106);
nand U20057 (N_20057,N_19475,N_19802);
nor U20058 (N_20058,N_19440,N_19060);
nand U20059 (N_20059,N_19832,N_19081);
or U20060 (N_20060,N_19093,N_19524);
nor U20061 (N_20061,N_19639,N_19622);
nor U20062 (N_20062,N_19984,N_19457);
nor U20063 (N_20063,N_19938,N_19906);
nand U20064 (N_20064,N_19282,N_19585);
xnor U20065 (N_20065,N_19252,N_19367);
nor U20066 (N_20066,N_19021,N_19471);
nand U20067 (N_20067,N_19674,N_19031);
or U20068 (N_20068,N_19575,N_19944);
or U20069 (N_20069,N_19957,N_19541);
xnor U20070 (N_20070,N_19403,N_19080);
nor U20071 (N_20071,N_19438,N_19661);
nand U20072 (N_20072,N_19560,N_19805);
and U20073 (N_20073,N_19056,N_19798);
or U20074 (N_20074,N_19939,N_19045);
xnor U20075 (N_20075,N_19722,N_19934);
xnor U20076 (N_20076,N_19193,N_19126);
nor U20077 (N_20077,N_19419,N_19785);
nand U20078 (N_20078,N_19226,N_19001);
nor U20079 (N_20079,N_19961,N_19846);
xnor U20080 (N_20080,N_19151,N_19869);
or U20081 (N_20081,N_19364,N_19628);
xnor U20082 (N_20082,N_19992,N_19366);
xor U20083 (N_20083,N_19235,N_19721);
and U20084 (N_20084,N_19778,N_19147);
and U20085 (N_20085,N_19284,N_19421);
nand U20086 (N_20086,N_19496,N_19724);
nand U20087 (N_20087,N_19775,N_19583);
nor U20088 (N_20088,N_19723,N_19265);
and U20089 (N_20089,N_19122,N_19225);
nand U20090 (N_20090,N_19715,N_19355);
and U20091 (N_20091,N_19296,N_19243);
and U20092 (N_20092,N_19787,N_19258);
xnor U20093 (N_20093,N_19544,N_19167);
or U20094 (N_20094,N_19014,N_19977);
and U20095 (N_20095,N_19529,N_19084);
xor U20096 (N_20096,N_19433,N_19700);
nand U20097 (N_20097,N_19997,N_19444);
nand U20098 (N_20098,N_19838,N_19261);
xnor U20099 (N_20099,N_19229,N_19458);
and U20100 (N_20100,N_19890,N_19768);
and U20101 (N_20101,N_19201,N_19755);
and U20102 (N_20102,N_19437,N_19881);
nand U20103 (N_20103,N_19910,N_19631);
xnor U20104 (N_20104,N_19276,N_19222);
xnor U20105 (N_20105,N_19988,N_19871);
and U20106 (N_20106,N_19038,N_19062);
or U20107 (N_20107,N_19155,N_19809);
xnor U20108 (N_20108,N_19259,N_19966);
nor U20109 (N_20109,N_19416,N_19975);
and U20110 (N_20110,N_19315,N_19519);
and U20111 (N_20111,N_19777,N_19922);
xor U20112 (N_20112,N_19835,N_19582);
xor U20113 (N_20113,N_19445,N_19558);
and U20114 (N_20114,N_19088,N_19637);
nand U20115 (N_20115,N_19000,N_19587);
or U20116 (N_20116,N_19752,N_19788);
xnor U20117 (N_20117,N_19859,N_19268);
and U20118 (N_20118,N_19668,N_19929);
nand U20119 (N_20119,N_19746,N_19624);
xor U20120 (N_20120,N_19867,N_19810);
or U20121 (N_20121,N_19439,N_19868);
or U20122 (N_20122,N_19159,N_19144);
or U20123 (N_20123,N_19333,N_19174);
and U20124 (N_20124,N_19508,N_19211);
nor U20125 (N_20125,N_19659,N_19565);
nand U20126 (N_20126,N_19842,N_19964);
nor U20127 (N_20127,N_19783,N_19359);
xor U20128 (N_20128,N_19843,N_19442);
xor U20129 (N_20129,N_19916,N_19327);
xor U20130 (N_20130,N_19454,N_19418);
nor U20131 (N_20131,N_19663,N_19727);
nand U20132 (N_20132,N_19606,N_19904);
nor U20133 (N_20133,N_19391,N_19128);
and U20134 (N_20134,N_19223,N_19203);
xnor U20135 (N_20135,N_19401,N_19369);
nor U20136 (N_20136,N_19804,N_19200);
and U20137 (N_20137,N_19145,N_19792);
nor U20138 (N_20138,N_19772,N_19841);
and U20139 (N_20139,N_19169,N_19063);
or U20140 (N_20140,N_19094,N_19958);
and U20141 (N_20141,N_19370,N_19930);
or U20142 (N_20142,N_19591,N_19068);
and U20143 (N_20143,N_19815,N_19047);
nand U20144 (N_20144,N_19525,N_19067);
nor U20145 (N_20145,N_19954,N_19605);
nand U20146 (N_20146,N_19323,N_19116);
nand U20147 (N_20147,N_19368,N_19828);
and U20148 (N_20148,N_19963,N_19765);
xor U20149 (N_20149,N_19250,N_19016);
nand U20150 (N_20150,N_19993,N_19059);
or U20151 (N_20151,N_19255,N_19168);
nand U20152 (N_20152,N_19202,N_19353);
or U20153 (N_20153,N_19753,N_19314);
or U20154 (N_20154,N_19850,N_19481);
and U20155 (N_20155,N_19645,N_19334);
nand U20156 (N_20156,N_19990,N_19875);
nand U20157 (N_20157,N_19170,N_19443);
xnor U20158 (N_20158,N_19199,N_19900);
nand U20159 (N_20159,N_19322,N_19339);
nor U20160 (N_20160,N_19640,N_19190);
xnor U20161 (N_20161,N_19549,N_19090);
nor U20162 (N_20162,N_19279,N_19742);
or U20163 (N_20163,N_19461,N_19620);
nand U20164 (N_20164,N_19361,N_19406);
xor U20165 (N_20165,N_19216,N_19617);
xor U20166 (N_20166,N_19076,N_19536);
xor U20167 (N_20167,N_19487,N_19613);
or U20168 (N_20168,N_19580,N_19188);
and U20169 (N_20169,N_19987,N_19394);
nand U20170 (N_20170,N_19288,N_19414);
nand U20171 (N_20171,N_19123,N_19705);
xor U20172 (N_20172,N_19491,N_19604);
nand U20173 (N_20173,N_19632,N_19950);
nor U20174 (N_20174,N_19267,N_19118);
xnor U20175 (N_20175,N_19220,N_19477);
nor U20176 (N_20176,N_19703,N_19297);
or U20177 (N_20177,N_19247,N_19198);
xor U20178 (N_20178,N_19132,N_19986);
nor U20179 (N_20179,N_19100,N_19069);
nand U20180 (N_20180,N_19256,N_19166);
xnor U20181 (N_20181,N_19214,N_19326);
nand U20182 (N_20182,N_19824,N_19207);
and U20183 (N_20183,N_19646,N_19534);
nor U20184 (N_20184,N_19589,N_19729);
or U20185 (N_20185,N_19649,N_19806);
xor U20186 (N_20186,N_19510,N_19281);
and U20187 (N_20187,N_19527,N_19395);
or U20188 (N_20188,N_19559,N_19572);
nand U20189 (N_20189,N_19257,N_19023);
xnor U20190 (N_20190,N_19763,N_19340);
nor U20191 (N_20191,N_19163,N_19012);
xor U20192 (N_20192,N_19127,N_19152);
or U20193 (N_20193,N_19593,N_19171);
xor U20194 (N_20194,N_19754,N_19381);
xnor U20195 (N_20195,N_19160,N_19230);
nor U20196 (N_20196,N_19295,N_19547);
nor U20197 (N_20197,N_19474,N_19670);
nor U20198 (N_20198,N_19736,N_19463);
nand U20199 (N_20199,N_19466,N_19399);
xor U20200 (N_20200,N_19398,N_19921);
nand U20201 (N_20201,N_19514,N_19937);
xnor U20202 (N_20202,N_19498,N_19427);
nand U20203 (N_20203,N_19928,N_19518);
xnor U20204 (N_20204,N_19283,N_19586);
or U20205 (N_20205,N_19134,N_19485);
nand U20206 (N_20206,N_19577,N_19522);
nand U20207 (N_20207,N_19855,N_19822);
and U20208 (N_20208,N_19330,N_19215);
xnor U20209 (N_20209,N_19897,N_19351);
and U20210 (N_20210,N_19600,N_19486);
nand U20211 (N_20211,N_19206,N_19112);
nand U20212 (N_20212,N_19253,N_19277);
or U20213 (N_20213,N_19566,N_19346);
nor U20214 (N_20214,N_19512,N_19209);
xor U20215 (N_20215,N_19647,N_19136);
and U20216 (N_20216,N_19782,N_19852);
nand U20217 (N_20217,N_19478,N_19390);
or U20218 (N_20218,N_19376,N_19015);
or U20219 (N_20219,N_19556,N_19013);
nor U20220 (N_20220,N_19175,N_19107);
xnor U20221 (N_20221,N_19156,N_19415);
xor U20222 (N_20222,N_19793,N_19683);
and U20223 (N_20223,N_19681,N_19465);
and U20224 (N_20224,N_19241,N_19164);
nand U20225 (N_20225,N_19133,N_19773);
nor U20226 (N_20226,N_19656,N_19280);
xor U20227 (N_20227,N_19396,N_19452);
xnor U20228 (N_20228,N_19373,N_19037);
xor U20229 (N_20229,N_19292,N_19960);
xnor U20230 (N_20230,N_19503,N_19825);
nand U20231 (N_20231,N_19111,N_19706);
and U20232 (N_20232,N_19610,N_19973);
xor U20233 (N_20233,N_19404,N_19687);
nand U20234 (N_20234,N_19099,N_19576);
nand U20235 (N_20235,N_19821,N_19316);
nor U20236 (N_20236,N_19077,N_19959);
nor U20237 (N_20237,N_19232,N_19495);
and U20238 (N_20238,N_19146,N_19371);
nor U20239 (N_20239,N_19905,N_19446);
xor U20240 (N_20240,N_19648,N_19862);
or U20241 (N_20241,N_19644,N_19848);
and U20242 (N_20242,N_19927,N_19464);
xnor U20243 (N_20243,N_19856,N_19671);
and U20244 (N_20244,N_19034,N_19303);
or U20245 (N_20245,N_19702,N_19289);
xnor U20246 (N_20246,N_19618,N_19539);
nand U20247 (N_20247,N_19623,N_19429);
xor U20248 (N_20248,N_19228,N_19985);
and U20249 (N_20249,N_19883,N_19830);
xor U20250 (N_20250,N_19642,N_19363);
nand U20251 (N_20251,N_19161,N_19389);
xor U20252 (N_20252,N_19803,N_19238);
and U20253 (N_20253,N_19248,N_19291);
xnor U20254 (N_20254,N_19699,N_19026);
nand U20255 (N_20255,N_19713,N_19678);
nor U20256 (N_20256,N_19140,N_19273);
or U20257 (N_20257,N_19331,N_19006);
xor U20258 (N_20258,N_19573,N_19294);
and U20259 (N_20259,N_19075,N_19744);
and U20260 (N_20260,N_19057,N_19043);
nand U20261 (N_20261,N_19635,N_19823);
nand U20262 (N_20262,N_19837,N_19749);
nand U20263 (N_20263,N_19886,N_19712);
or U20264 (N_20264,N_19441,N_19506);
nand U20265 (N_20265,N_19634,N_19212);
or U20266 (N_20266,N_19857,N_19704);
xor U20267 (N_20267,N_19183,N_19626);
nor U20268 (N_20268,N_19816,N_19377);
or U20269 (N_20269,N_19138,N_19526);
and U20270 (N_20270,N_19182,N_19980);
or U20271 (N_20271,N_19968,N_19050);
nand U20272 (N_20272,N_19808,N_19629);
nor U20273 (N_20273,N_19833,N_19951);
and U20274 (N_20274,N_19840,N_19854);
or U20275 (N_20275,N_19731,N_19194);
and U20276 (N_20276,N_19468,N_19885);
nand U20277 (N_20277,N_19548,N_19563);
nand U20278 (N_20278,N_19535,N_19499);
nor U20279 (N_20279,N_19949,N_19747);
and U20280 (N_20280,N_19451,N_19470);
or U20281 (N_20281,N_19571,N_19919);
and U20282 (N_20282,N_19236,N_19638);
and U20283 (N_20283,N_19237,N_19383);
nand U20284 (N_20284,N_19745,N_19991);
or U20285 (N_20285,N_19989,N_19272);
and U20286 (N_20286,N_19172,N_19909);
nand U20287 (N_20287,N_19818,N_19335);
nor U20288 (N_20288,N_19298,N_19847);
xor U20289 (N_20289,N_19148,N_19597);
and U20290 (N_20290,N_19578,N_19790);
nand U20291 (N_20291,N_19052,N_19379);
nor U20292 (N_20292,N_19137,N_19899);
or U20293 (N_20293,N_19696,N_19387);
nand U20294 (N_20294,N_19728,N_19124);
nand U20295 (N_20295,N_19302,N_19933);
and U20296 (N_20296,N_19197,N_19042);
and U20297 (N_20297,N_19003,N_19679);
and U20298 (N_20298,N_19320,N_19515);
or U20299 (N_20299,N_19889,N_19378);
nand U20300 (N_20300,N_19480,N_19611);
nand U20301 (N_20301,N_19180,N_19408);
nor U20302 (N_20302,N_19365,N_19109);
nand U20303 (N_20303,N_19337,N_19309);
and U20304 (N_20304,N_19115,N_19129);
or U20305 (N_20305,N_19500,N_19762);
nand U20306 (N_20306,N_19254,N_19332);
nor U20307 (N_20307,N_19098,N_19103);
nand U20308 (N_20308,N_19956,N_19285);
nand U20309 (N_20309,N_19185,N_19150);
nand U20310 (N_20310,N_19509,N_19092);
nor U20311 (N_20311,N_19983,N_19627);
nand U20312 (N_20312,N_19943,N_19234);
nor U20313 (N_20313,N_19511,N_19430);
and U20314 (N_20314,N_19044,N_19579);
or U20315 (N_20315,N_19523,N_19336);
and U20316 (N_20316,N_19455,N_19952);
or U20317 (N_20317,N_19872,N_19581);
nor U20318 (N_20318,N_19532,N_19748);
xnor U20319 (N_20319,N_19025,N_19040);
nor U20320 (N_20320,N_19967,N_19733);
nor U20321 (N_20321,N_19010,N_19865);
xnor U20322 (N_20322,N_19459,N_19970);
nand U20323 (N_20323,N_19338,N_19665);
nand U20324 (N_20324,N_19962,N_19407);
nand U20325 (N_20325,N_19184,N_19130);
and U20326 (N_20326,N_19426,N_19650);
and U20327 (N_20327,N_19866,N_19384);
and U20328 (N_20328,N_19244,N_19791);
or U20329 (N_20329,N_19813,N_19374);
nand U20330 (N_20330,N_19004,N_19520);
nor U20331 (N_20331,N_19312,N_19870);
or U20332 (N_20332,N_19501,N_19318);
and U20333 (N_20333,N_19342,N_19795);
xnor U20334 (N_20334,N_19730,N_19619);
and U20335 (N_20335,N_19456,N_19345);
nor U20336 (N_20336,N_19800,N_19555);
nor U20337 (N_20337,N_19694,N_19676);
nand U20338 (N_20338,N_19811,N_19319);
nor U20339 (N_20339,N_19750,N_19658);
or U20340 (N_20340,N_19574,N_19208);
or U20341 (N_20341,N_19385,N_19915);
and U20342 (N_20342,N_19902,N_19654);
xor U20343 (N_20343,N_19058,N_19796);
nor U20344 (N_20344,N_19891,N_19502);
nor U20345 (N_20345,N_19751,N_19507);
xor U20346 (N_20346,N_19231,N_19097);
xnor U20347 (N_20347,N_19033,N_19690);
or U20348 (N_20348,N_19643,N_19820);
and U20349 (N_20349,N_19766,N_19531);
and U20350 (N_20350,N_19493,N_19362);
or U20351 (N_20351,N_19274,N_19344);
nand U20352 (N_20352,N_19139,N_19667);
nor U20353 (N_20353,N_19357,N_19425);
and U20354 (N_20354,N_19863,N_19269);
nor U20355 (N_20355,N_19720,N_19781);
xor U20356 (N_20356,N_19633,N_19769);
nor U20357 (N_20357,N_19546,N_19213);
or U20358 (N_20358,N_19349,N_19741);
or U20359 (N_20359,N_19776,N_19568);
and U20360 (N_20360,N_19924,N_19614);
nor U20361 (N_20361,N_19947,N_19758);
or U20362 (N_20362,N_19903,N_19423);
and U20363 (N_20363,N_19245,N_19176);
xnor U20364 (N_20364,N_19771,N_19221);
xnor U20365 (N_20365,N_19141,N_19114);
nand U20366 (N_20366,N_19249,N_19562);
xor U20367 (N_20367,N_19356,N_19517);
nand U20368 (N_20368,N_19002,N_19912);
nand U20369 (N_20369,N_19923,N_19926);
and U20370 (N_20370,N_19607,N_19096);
xnor U20371 (N_20371,N_19450,N_19698);
nor U20372 (N_20372,N_19757,N_19382);
xnor U20373 (N_20373,N_19055,N_19239);
and U20374 (N_20374,N_19405,N_19567);
xor U20375 (N_20375,N_19117,N_19095);
nor U20376 (N_20376,N_19343,N_19492);
or U20377 (N_20377,N_19784,N_19693);
and U20378 (N_20378,N_19469,N_19131);
nand U20379 (N_20379,N_19734,N_19041);
xor U20380 (N_20380,N_19995,N_19789);
xor U20381 (N_20381,N_19942,N_19260);
and U20382 (N_20382,N_19287,N_19530);
nor U20383 (N_20383,N_19488,N_19641);
and U20384 (N_20384,N_19601,N_19032);
xor U20385 (N_20385,N_19087,N_19422);
nand U20386 (N_20386,N_19205,N_19972);
and U20387 (N_20387,N_19301,N_19102);
nand U20388 (N_20388,N_19978,N_19911);
nor U20389 (N_20389,N_19707,N_19027);
nand U20390 (N_20390,N_19625,N_19125);
nor U20391 (N_20391,N_19048,N_19908);
nand U20392 (N_20392,N_19086,N_19738);
nand U20393 (N_20393,N_19300,N_19760);
or U20394 (N_20394,N_19286,N_19874);
nor U20395 (N_20395,N_19479,N_19774);
or U20396 (N_20396,N_19584,N_19447);
nor U20397 (N_20397,N_19089,N_19686);
or U20398 (N_20398,N_19072,N_19192);
or U20399 (N_20399,N_19263,N_19845);
xor U20400 (N_20400,N_19350,N_19070);
and U20401 (N_20401,N_19920,N_19814);
xor U20402 (N_20402,N_19317,N_19360);
nand U20403 (N_20403,N_19969,N_19264);
xor U20404 (N_20404,N_19651,N_19653);
or U20405 (N_20405,N_19153,N_19189);
and U20406 (N_20406,N_19186,N_19599);
and U20407 (N_20407,N_19677,N_19936);
or U20408 (N_20408,N_19590,N_19494);
or U20409 (N_20409,N_19955,N_19940);
or U20410 (N_20410,N_19410,N_19462);
nor U20411 (N_20411,N_19178,N_19680);
or U20412 (N_20412,N_19431,N_19380);
xnor U20413 (N_20413,N_19817,N_19030);
and U20414 (N_20414,N_19538,N_19473);
nor U20415 (N_20415,N_19227,N_19533);
and U20416 (N_20416,N_19420,N_19290);
xor U20417 (N_20417,N_19082,N_19348);
and U20418 (N_20418,N_19307,N_19341);
nor U20419 (N_20419,N_19308,N_19764);
xnor U20420 (N_20420,N_19434,N_19306);
and U20421 (N_20421,N_19554,N_19770);
nor U20422 (N_20422,N_19946,N_19372);
nor U20423 (N_20423,N_19449,N_19612);
nor U20424 (N_20424,N_19436,N_19894);
xor U20425 (N_20425,N_19608,N_19945);
nand U20426 (N_20426,N_19157,N_19210);
and U20427 (N_20427,N_19876,N_19829);
and U20428 (N_20428,N_19895,N_19009);
or U20429 (N_20429,N_19299,N_19917);
and U20430 (N_20430,N_19941,N_19028);
xor U20431 (N_20431,N_19119,N_19262);
xnor U20432 (N_20432,N_19979,N_19826);
nor U20433 (N_20433,N_19233,N_19321);
and U20434 (N_20434,N_19685,N_19251);
or U20435 (N_20435,N_19162,N_19101);
and U20436 (N_20436,N_19878,N_19393);
and U20437 (N_20437,N_19046,N_19246);
nor U20438 (N_20438,N_19154,N_19179);
and U20439 (N_20439,N_19329,N_19692);
xor U20440 (N_20440,N_19807,N_19008);
and U20441 (N_20441,N_19786,N_19691);
or U20442 (N_20442,N_19615,N_19932);
nor U20443 (N_20443,N_19689,N_19794);
nand U20444 (N_20444,N_19592,N_19711);
nor U20445 (N_20445,N_19036,N_19411);
or U20446 (N_20446,N_19861,N_19965);
nor U20447 (N_20447,N_19049,N_19412);
nand U20448 (N_20448,N_19598,N_19424);
xor U20449 (N_20449,N_19652,N_19719);
nand U20450 (N_20450,N_19521,N_19588);
nand U20451 (N_20451,N_19275,N_19053);
and U20452 (N_20452,N_19864,N_19971);
or U20453 (N_20453,N_19484,N_19400);
nand U20454 (N_20454,N_19065,N_19402);
nand U20455 (N_20455,N_19594,N_19195);
and U20456 (N_20456,N_19662,N_19310);
xnor U20457 (N_20457,N_19354,N_19879);
or U20458 (N_20458,N_19636,N_19552);
or U20459 (N_20459,N_19039,N_19204);
nand U20460 (N_20460,N_19224,N_19121);
nor U20461 (N_20461,N_19108,N_19064);
and U20462 (N_20462,N_19851,N_19017);
and U20463 (N_20463,N_19181,N_19673);
nor U20464 (N_20464,N_19737,N_19328);
xnor U20465 (N_20465,N_19240,N_19120);
nand U20466 (N_20466,N_19718,N_19569);
and U20467 (N_20467,N_19931,N_19409);
and U20468 (N_20468,N_19110,N_19682);
xor U20469 (N_20469,N_19767,N_19489);
xor U20470 (N_20470,N_19483,N_19553);
nand U20471 (N_20471,N_19143,N_19896);
or U20472 (N_20472,N_19710,N_19994);
nand U20473 (N_20473,N_19688,N_19797);
nor U20474 (N_20474,N_19550,N_19005);
nor U20475 (N_20475,N_19073,N_19880);
or U20476 (N_20476,N_19918,N_19078);
and U20477 (N_20477,N_19756,N_19011);
and U20478 (N_20478,N_19888,N_19999);
nor U20479 (N_20479,N_19831,N_19914);
or U20480 (N_20480,N_19893,N_19935);
nand U20481 (N_20481,N_19630,N_19561);
xnor U20482 (N_20482,N_19853,N_19165);
xor U20483 (N_20483,N_19545,N_19542);
xnor U20484 (N_20484,N_19083,N_19697);
xnor U20485 (N_20485,N_19352,N_19761);
and U20486 (N_20486,N_19432,N_19187);
nor U20487 (N_20487,N_19504,N_19528);
nand U20488 (N_20488,N_19877,N_19104);
and U20489 (N_20489,N_19325,N_19428);
nand U20490 (N_20490,N_19812,N_19022);
or U20491 (N_20491,N_19020,N_19602);
nor U20492 (N_20492,N_19982,N_19827);
and U20493 (N_20493,N_19173,N_19998);
nor U20494 (N_20494,N_19739,N_19672);
xnor U20495 (N_20495,N_19029,N_19217);
nand U20496 (N_20496,N_19490,N_19516);
and U20497 (N_20497,N_19655,N_19091);
and U20498 (N_20498,N_19657,N_19540);
or U20499 (N_20499,N_19884,N_19448);
xor U20500 (N_20500,N_19188,N_19558);
nor U20501 (N_20501,N_19685,N_19415);
xor U20502 (N_20502,N_19114,N_19632);
xor U20503 (N_20503,N_19854,N_19361);
and U20504 (N_20504,N_19937,N_19022);
nor U20505 (N_20505,N_19446,N_19930);
or U20506 (N_20506,N_19558,N_19720);
or U20507 (N_20507,N_19615,N_19418);
nand U20508 (N_20508,N_19540,N_19225);
xor U20509 (N_20509,N_19061,N_19320);
xnor U20510 (N_20510,N_19596,N_19416);
or U20511 (N_20511,N_19561,N_19969);
nor U20512 (N_20512,N_19695,N_19973);
and U20513 (N_20513,N_19842,N_19149);
and U20514 (N_20514,N_19971,N_19578);
xor U20515 (N_20515,N_19576,N_19798);
and U20516 (N_20516,N_19763,N_19038);
xnor U20517 (N_20517,N_19728,N_19110);
or U20518 (N_20518,N_19713,N_19599);
nand U20519 (N_20519,N_19708,N_19758);
nor U20520 (N_20520,N_19436,N_19572);
and U20521 (N_20521,N_19813,N_19250);
nand U20522 (N_20522,N_19755,N_19424);
or U20523 (N_20523,N_19400,N_19031);
xor U20524 (N_20524,N_19924,N_19047);
xor U20525 (N_20525,N_19559,N_19424);
and U20526 (N_20526,N_19616,N_19155);
and U20527 (N_20527,N_19285,N_19552);
nor U20528 (N_20528,N_19996,N_19155);
nand U20529 (N_20529,N_19000,N_19159);
xnor U20530 (N_20530,N_19294,N_19287);
or U20531 (N_20531,N_19198,N_19187);
and U20532 (N_20532,N_19585,N_19534);
and U20533 (N_20533,N_19459,N_19192);
xor U20534 (N_20534,N_19340,N_19549);
nand U20535 (N_20535,N_19185,N_19149);
nor U20536 (N_20536,N_19697,N_19492);
and U20537 (N_20537,N_19751,N_19441);
nor U20538 (N_20538,N_19874,N_19141);
xnor U20539 (N_20539,N_19899,N_19113);
or U20540 (N_20540,N_19636,N_19499);
nor U20541 (N_20541,N_19469,N_19277);
nor U20542 (N_20542,N_19101,N_19240);
or U20543 (N_20543,N_19550,N_19798);
and U20544 (N_20544,N_19314,N_19184);
nor U20545 (N_20545,N_19025,N_19444);
nand U20546 (N_20546,N_19969,N_19563);
xor U20547 (N_20547,N_19414,N_19421);
xor U20548 (N_20548,N_19991,N_19947);
xor U20549 (N_20549,N_19722,N_19751);
nand U20550 (N_20550,N_19265,N_19690);
or U20551 (N_20551,N_19617,N_19839);
and U20552 (N_20552,N_19504,N_19012);
nand U20553 (N_20553,N_19975,N_19535);
nand U20554 (N_20554,N_19292,N_19870);
or U20555 (N_20555,N_19350,N_19588);
or U20556 (N_20556,N_19793,N_19183);
xnor U20557 (N_20557,N_19427,N_19494);
nor U20558 (N_20558,N_19945,N_19079);
or U20559 (N_20559,N_19543,N_19275);
nor U20560 (N_20560,N_19897,N_19960);
nor U20561 (N_20561,N_19786,N_19530);
nor U20562 (N_20562,N_19489,N_19056);
nand U20563 (N_20563,N_19060,N_19538);
or U20564 (N_20564,N_19820,N_19185);
nor U20565 (N_20565,N_19487,N_19485);
and U20566 (N_20566,N_19789,N_19269);
or U20567 (N_20567,N_19964,N_19599);
and U20568 (N_20568,N_19901,N_19972);
and U20569 (N_20569,N_19336,N_19302);
nor U20570 (N_20570,N_19716,N_19742);
nand U20571 (N_20571,N_19203,N_19859);
nand U20572 (N_20572,N_19105,N_19640);
nor U20573 (N_20573,N_19301,N_19859);
nand U20574 (N_20574,N_19086,N_19456);
xor U20575 (N_20575,N_19592,N_19703);
nand U20576 (N_20576,N_19122,N_19603);
and U20577 (N_20577,N_19989,N_19186);
or U20578 (N_20578,N_19422,N_19394);
xnor U20579 (N_20579,N_19292,N_19326);
or U20580 (N_20580,N_19664,N_19685);
nor U20581 (N_20581,N_19375,N_19292);
and U20582 (N_20582,N_19391,N_19310);
or U20583 (N_20583,N_19811,N_19904);
xor U20584 (N_20584,N_19602,N_19996);
and U20585 (N_20585,N_19140,N_19008);
nand U20586 (N_20586,N_19154,N_19552);
xnor U20587 (N_20587,N_19841,N_19115);
or U20588 (N_20588,N_19291,N_19242);
and U20589 (N_20589,N_19505,N_19813);
nor U20590 (N_20590,N_19413,N_19248);
nand U20591 (N_20591,N_19628,N_19725);
or U20592 (N_20592,N_19565,N_19482);
xnor U20593 (N_20593,N_19355,N_19400);
nand U20594 (N_20594,N_19761,N_19567);
nand U20595 (N_20595,N_19344,N_19803);
or U20596 (N_20596,N_19366,N_19002);
xnor U20597 (N_20597,N_19484,N_19968);
nor U20598 (N_20598,N_19736,N_19777);
nand U20599 (N_20599,N_19027,N_19258);
xor U20600 (N_20600,N_19610,N_19569);
nor U20601 (N_20601,N_19128,N_19364);
and U20602 (N_20602,N_19607,N_19956);
and U20603 (N_20603,N_19968,N_19674);
nor U20604 (N_20604,N_19164,N_19005);
or U20605 (N_20605,N_19225,N_19669);
and U20606 (N_20606,N_19150,N_19318);
nand U20607 (N_20607,N_19909,N_19031);
and U20608 (N_20608,N_19980,N_19857);
nand U20609 (N_20609,N_19126,N_19545);
and U20610 (N_20610,N_19124,N_19267);
and U20611 (N_20611,N_19289,N_19045);
xor U20612 (N_20612,N_19448,N_19436);
or U20613 (N_20613,N_19535,N_19649);
xor U20614 (N_20614,N_19233,N_19414);
and U20615 (N_20615,N_19878,N_19562);
and U20616 (N_20616,N_19818,N_19977);
nor U20617 (N_20617,N_19567,N_19864);
nor U20618 (N_20618,N_19410,N_19234);
nand U20619 (N_20619,N_19281,N_19116);
nor U20620 (N_20620,N_19014,N_19137);
or U20621 (N_20621,N_19381,N_19074);
xnor U20622 (N_20622,N_19372,N_19497);
nor U20623 (N_20623,N_19487,N_19893);
and U20624 (N_20624,N_19617,N_19819);
and U20625 (N_20625,N_19102,N_19488);
xnor U20626 (N_20626,N_19482,N_19479);
or U20627 (N_20627,N_19881,N_19998);
nor U20628 (N_20628,N_19475,N_19357);
nand U20629 (N_20629,N_19959,N_19019);
nand U20630 (N_20630,N_19820,N_19553);
or U20631 (N_20631,N_19171,N_19174);
or U20632 (N_20632,N_19674,N_19927);
nand U20633 (N_20633,N_19795,N_19750);
nor U20634 (N_20634,N_19266,N_19325);
nand U20635 (N_20635,N_19140,N_19029);
xor U20636 (N_20636,N_19538,N_19292);
or U20637 (N_20637,N_19285,N_19360);
xor U20638 (N_20638,N_19745,N_19249);
nand U20639 (N_20639,N_19857,N_19074);
and U20640 (N_20640,N_19647,N_19250);
or U20641 (N_20641,N_19607,N_19253);
nand U20642 (N_20642,N_19399,N_19253);
or U20643 (N_20643,N_19105,N_19905);
or U20644 (N_20644,N_19651,N_19445);
nand U20645 (N_20645,N_19564,N_19977);
nand U20646 (N_20646,N_19115,N_19884);
xnor U20647 (N_20647,N_19462,N_19341);
and U20648 (N_20648,N_19063,N_19914);
or U20649 (N_20649,N_19818,N_19628);
xor U20650 (N_20650,N_19826,N_19069);
and U20651 (N_20651,N_19702,N_19048);
nor U20652 (N_20652,N_19977,N_19520);
xnor U20653 (N_20653,N_19943,N_19617);
or U20654 (N_20654,N_19170,N_19264);
nand U20655 (N_20655,N_19973,N_19036);
nand U20656 (N_20656,N_19514,N_19193);
nand U20657 (N_20657,N_19221,N_19508);
or U20658 (N_20658,N_19520,N_19455);
nor U20659 (N_20659,N_19346,N_19044);
xor U20660 (N_20660,N_19602,N_19961);
nand U20661 (N_20661,N_19823,N_19282);
and U20662 (N_20662,N_19452,N_19520);
xor U20663 (N_20663,N_19617,N_19487);
or U20664 (N_20664,N_19047,N_19238);
and U20665 (N_20665,N_19104,N_19943);
or U20666 (N_20666,N_19067,N_19338);
nor U20667 (N_20667,N_19764,N_19126);
nand U20668 (N_20668,N_19303,N_19135);
nand U20669 (N_20669,N_19465,N_19829);
nand U20670 (N_20670,N_19821,N_19460);
and U20671 (N_20671,N_19469,N_19314);
or U20672 (N_20672,N_19131,N_19440);
nand U20673 (N_20673,N_19783,N_19278);
nand U20674 (N_20674,N_19554,N_19679);
nand U20675 (N_20675,N_19591,N_19482);
nor U20676 (N_20676,N_19321,N_19655);
or U20677 (N_20677,N_19702,N_19511);
or U20678 (N_20678,N_19444,N_19799);
xor U20679 (N_20679,N_19449,N_19978);
nand U20680 (N_20680,N_19133,N_19050);
and U20681 (N_20681,N_19494,N_19789);
xnor U20682 (N_20682,N_19721,N_19645);
xor U20683 (N_20683,N_19782,N_19553);
or U20684 (N_20684,N_19417,N_19268);
or U20685 (N_20685,N_19651,N_19856);
and U20686 (N_20686,N_19638,N_19843);
nor U20687 (N_20687,N_19996,N_19128);
and U20688 (N_20688,N_19614,N_19572);
and U20689 (N_20689,N_19382,N_19599);
nor U20690 (N_20690,N_19730,N_19876);
nor U20691 (N_20691,N_19370,N_19422);
xnor U20692 (N_20692,N_19178,N_19424);
nor U20693 (N_20693,N_19312,N_19641);
and U20694 (N_20694,N_19799,N_19670);
nor U20695 (N_20695,N_19799,N_19650);
nand U20696 (N_20696,N_19948,N_19311);
and U20697 (N_20697,N_19993,N_19877);
nor U20698 (N_20698,N_19869,N_19437);
nand U20699 (N_20699,N_19634,N_19671);
xor U20700 (N_20700,N_19866,N_19744);
xnor U20701 (N_20701,N_19834,N_19425);
and U20702 (N_20702,N_19295,N_19591);
nand U20703 (N_20703,N_19317,N_19660);
nand U20704 (N_20704,N_19385,N_19573);
and U20705 (N_20705,N_19021,N_19889);
nand U20706 (N_20706,N_19288,N_19342);
nand U20707 (N_20707,N_19659,N_19532);
xnor U20708 (N_20708,N_19158,N_19508);
and U20709 (N_20709,N_19838,N_19473);
or U20710 (N_20710,N_19204,N_19394);
xnor U20711 (N_20711,N_19527,N_19970);
xor U20712 (N_20712,N_19745,N_19911);
nand U20713 (N_20713,N_19258,N_19245);
nor U20714 (N_20714,N_19336,N_19626);
nand U20715 (N_20715,N_19512,N_19398);
and U20716 (N_20716,N_19011,N_19082);
nand U20717 (N_20717,N_19993,N_19667);
nand U20718 (N_20718,N_19783,N_19054);
and U20719 (N_20719,N_19835,N_19781);
nor U20720 (N_20720,N_19673,N_19294);
and U20721 (N_20721,N_19715,N_19657);
nand U20722 (N_20722,N_19639,N_19075);
nand U20723 (N_20723,N_19512,N_19395);
nand U20724 (N_20724,N_19077,N_19082);
nand U20725 (N_20725,N_19370,N_19735);
nand U20726 (N_20726,N_19071,N_19742);
xnor U20727 (N_20727,N_19542,N_19571);
or U20728 (N_20728,N_19039,N_19688);
or U20729 (N_20729,N_19409,N_19510);
nand U20730 (N_20730,N_19049,N_19847);
nor U20731 (N_20731,N_19618,N_19829);
or U20732 (N_20732,N_19732,N_19158);
nor U20733 (N_20733,N_19973,N_19197);
xor U20734 (N_20734,N_19896,N_19925);
or U20735 (N_20735,N_19942,N_19816);
or U20736 (N_20736,N_19860,N_19272);
nor U20737 (N_20737,N_19103,N_19006);
and U20738 (N_20738,N_19574,N_19272);
or U20739 (N_20739,N_19561,N_19863);
nand U20740 (N_20740,N_19698,N_19893);
nand U20741 (N_20741,N_19233,N_19715);
nand U20742 (N_20742,N_19553,N_19075);
xnor U20743 (N_20743,N_19024,N_19098);
or U20744 (N_20744,N_19003,N_19785);
xnor U20745 (N_20745,N_19804,N_19370);
or U20746 (N_20746,N_19515,N_19808);
xor U20747 (N_20747,N_19376,N_19866);
and U20748 (N_20748,N_19064,N_19184);
xor U20749 (N_20749,N_19438,N_19324);
and U20750 (N_20750,N_19784,N_19871);
xor U20751 (N_20751,N_19059,N_19306);
or U20752 (N_20752,N_19005,N_19534);
and U20753 (N_20753,N_19444,N_19044);
nor U20754 (N_20754,N_19058,N_19531);
nand U20755 (N_20755,N_19180,N_19105);
nand U20756 (N_20756,N_19978,N_19753);
xnor U20757 (N_20757,N_19166,N_19896);
nand U20758 (N_20758,N_19424,N_19381);
nor U20759 (N_20759,N_19010,N_19547);
or U20760 (N_20760,N_19727,N_19022);
nor U20761 (N_20761,N_19166,N_19467);
xor U20762 (N_20762,N_19687,N_19704);
or U20763 (N_20763,N_19306,N_19199);
or U20764 (N_20764,N_19054,N_19457);
and U20765 (N_20765,N_19762,N_19137);
xnor U20766 (N_20766,N_19105,N_19977);
xnor U20767 (N_20767,N_19005,N_19360);
nand U20768 (N_20768,N_19523,N_19421);
xor U20769 (N_20769,N_19977,N_19529);
nand U20770 (N_20770,N_19764,N_19659);
nand U20771 (N_20771,N_19710,N_19528);
and U20772 (N_20772,N_19295,N_19234);
nor U20773 (N_20773,N_19429,N_19144);
and U20774 (N_20774,N_19546,N_19682);
or U20775 (N_20775,N_19163,N_19335);
nor U20776 (N_20776,N_19157,N_19152);
or U20777 (N_20777,N_19578,N_19407);
nor U20778 (N_20778,N_19390,N_19506);
or U20779 (N_20779,N_19405,N_19873);
xor U20780 (N_20780,N_19514,N_19828);
xnor U20781 (N_20781,N_19641,N_19048);
xnor U20782 (N_20782,N_19121,N_19156);
and U20783 (N_20783,N_19265,N_19176);
xor U20784 (N_20784,N_19784,N_19846);
or U20785 (N_20785,N_19719,N_19158);
and U20786 (N_20786,N_19982,N_19767);
xor U20787 (N_20787,N_19906,N_19992);
xor U20788 (N_20788,N_19167,N_19749);
and U20789 (N_20789,N_19816,N_19709);
nand U20790 (N_20790,N_19331,N_19631);
xnor U20791 (N_20791,N_19352,N_19212);
nor U20792 (N_20792,N_19022,N_19129);
nor U20793 (N_20793,N_19338,N_19129);
and U20794 (N_20794,N_19310,N_19947);
or U20795 (N_20795,N_19436,N_19950);
xor U20796 (N_20796,N_19490,N_19503);
xnor U20797 (N_20797,N_19964,N_19469);
and U20798 (N_20798,N_19983,N_19195);
and U20799 (N_20799,N_19958,N_19138);
xnor U20800 (N_20800,N_19164,N_19285);
nor U20801 (N_20801,N_19393,N_19863);
xor U20802 (N_20802,N_19948,N_19746);
nor U20803 (N_20803,N_19278,N_19434);
xor U20804 (N_20804,N_19254,N_19066);
or U20805 (N_20805,N_19940,N_19441);
nor U20806 (N_20806,N_19552,N_19120);
or U20807 (N_20807,N_19593,N_19478);
and U20808 (N_20808,N_19699,N_19629);
and U20809 (N_20809,N_19832,N_19448);
or U20810 (N_20810,N_19410,N_19131);
nand U20811 (N_20811,N_19972,N_19033);
xor U20812 (N_20812,N_19675,N_19876);
and U20813 (N_20813,N_19176,N_19740);
nand U20814 (N_20814,N_19051,N_19888);
xnor U20815 (N_20815,N_19769,N_19017);
nand U20816 (N_20816,N_19719,N_19084);
or U20817 (N_20817,N_19927,N_19870);
nand U20818 (N_20818,N_19753,N_19359);
or U20819 (N_20819,N_19822,N_19878);
nand U20820 (N_20820,N_19258,N_19869);
nor U20821 (N_20821,N_19432,N_19383);
nand U20822 (N_20822,N_19425,N_19517);
and U20823 (N_20823,N_19101,N_19844);
nor U20824 (N_20824,N_19639,N_19081);
nand U20825 (N_20825,N_19566,N_19011);
nor U20826 (N_20826,N_19932,N_19554);
nand U20827 (N_20827,N_19704,N_19916);
and U20828 (N_20828,N_19479,N_19509);
xnor U20829 (N_20829,N_19264,N_19097);
nand U20830 (N_20830,N_19230,N_19625);
and U20831 (N_20831,N_19426,N_19628);
nand U20832 (N_20832,N_19590,N_19446);
or U20833 (N_20833,N_19701,N_19826);
nor U20834 (N_20834,N_19261,N_19143);
xnor U20835 (N_20835,N_19128,N_19379);
or U20836 (N_20836,N_19913,N_19761);
nor U20837 (N_20837,N_19590,N_19513);
or U20838 (N_20838,N_19135,N_19871);
or U20839 (N_20839,N_19836,N_19571);
nand U20840 (N_20840,N_19343,N_19961);
nor U20841 (N_20841,N_19468,N_19016);
nor U20842 (N_20842,N_19357,N_19468);
xnor U20843 (N_20843,N_19563,N_19414);
xor U20844 (N_20844,N_19860,N_19369);
nand U20845 (N_20845,N_19076,N_19694);
nand U20846 (N_20846,N_19146,N_19915);
xor U20847 (N_20847,N_19565,N_19334);
nor U20848 (N_20848,N_19531,N_19573);
nor U20849 (N_20849,N_19392,N_19383);
nor U20850 (N_20850,N_19670,N_19772);
nor U20851 (N_20851,N_19969,N_19612);
nor U20852 (N_20852,N_19752,N_19649);
or U20853 (N_20853,N_19934,N_19845);
or U20854 (N_20854,N_19846,N_19288);
and U20855 (N_20855,N_19832,N_19406);
xor U20856 (N_20856,N_19365,N_19734);
nand U20857 (N_20857,N_19275,N_19986);
nor U20858 (N_20858,N_19270,N_19229);
nor U20859 (N_20859,N_19173,N_19280);
xor U20860 (N_20860,N_19825,N_19967);
and U20861 (N_20861,N_19452,N_19673);
nand U20862 (N_20862,N_19378,N_19077);
and U20863 (N_20863,N_19542,N_19895);
xnor U20864 (N_20864,N_19435,N_19549);
nor U20865 (N_20865,N_19941,N_19650);
nand U20866 (N_20866,N_19372,N_19994);
and U20867 (N_20867,N_19419,N_19174);
or U20868 (N_20868,N_19714,N_19173);
nor U20869 (N_20869,N_19005,N_19512);
nand U20870 (N_20870,N_19511,N_19411);
or U20871 (N_20871,N_19401,N_19463);
nor U20872 (N_20872,N_19180,N_19407);
nor U20873 (N_20873,N_19717,N_19471);
nand U20874 (N_20874,N_19452,N_19957);
nor U20875 (N_20875,N_19640,N_19506);
and U20876 (N_20876,N_19057,N_19206);
nor U20877 (N_20877,N_19125,N_19166);
nand U20878 (N_20878,N_19011,N_19873);
nor U20879 (N_20879,N_19262,N_19331);
and U20880 (N_20880,N_19474,N_19195);
nor U20881 (N_20881,N_19453,N_19636);
nor U20882 (N_20882,N_19109,N_19441);
nand U20883 (N_20883,N_19611,N_19270);
nor U20884 (N_20884,N_19806,N_19206);
nand U20885 (N_20885,N_19753,N_19723);
or U20886 (N_20886,N_19453,N_19890);
nand U20887 (N_20887,N_19345,N_19853);
or U20888 (N_20888,N_19847,N_19873);
or U20889 (N_20889,N_19901,N_19735);
and U20890 (N_20890,N_19731,N_19285);
or U20891 (N_20891,N_19062,N_19628);
or U20892 (N_20892,N_19711,N_19616);
nor U20893 (N_20893,N_19870,N_19148);
or U20894 (N_20894,N_19551,N_19632);
xor U20895 (N_20895,N_19641,N_19442);
xor U20896 (N_20896,N_19000,N_19177);
or U20897 (N_20897,N_19169,N_19904);
or U20898 (N_20898,N_19393,N_19352);
nor U20899 (N_20899,N_19715,N_19964);
and U20900 (N_20900,N_19481,N_19046);
nand U20901 (N_20901,N_19592,N_19051);
and U20902 (N_20902,N_19724,N_19631);
and U20903 (N_20903,N_19225,N_19898);
xnor U20904 (N_20904,N_19021,N_19851);
nor U20905 (N_20905,N_19768,N_19854);
nor U20906 (N_20906,N_19096,N_19310);
and U20907 (N_20907,N_19830,N_19360);
xor U20908 (N_20908,N_19538,N_19850);
and U20909 (N_20909,N_19094,N_19267);
and U20910 (N_20910,N_19779,N_19290);
or U20911 (N_20911,N_19076,N_19185);
xnor U20912 (N_20912,N_19901,N_19785);
xor U20913 (N_20913,N_19664,N_19120);
xnor U20914 (N_20914,N_19903,N_19682);
or U20915 (N_20915,N_19838,N_19082);
nor U20916 (N_20916,N_19526,N_19902);
xor U20917 (N_20917,N_19891,N_19954);
or U20918 (N_20918,N_19405,N_19691);
nor U20919 (N_20919,N_19902,N_19473);
nand U20920 (N_20920,N_19219,N_19525);
and U20921 (N_20921,N_19839,N_19364);
or U20922 (N_20922,N_19081,N_19833);
nand U20923 (N_20923,N_19604,N_19647);
and U20924 (N_20924,N_19834,N_19294);
nor U20925 (N_20925,N_19419,N_19230);
or U20926 (N_20926,N_19025,N_19023);
nand U20927 (N_20927,N_19413,N_19408);
nor U20928 (N_20928,N_19833,N_19717);
nand U20929 (N_20929,N_19811,N_19824);
nand U20930 (N_20930,N_19073,N_19527);
nor U20931 (N_20931,N_19059,N_19172);
or U20932 (N_20932,N_19251,N_19629);
and U20933 (N_20933,N_19084,N_19170);
nor U20934 (N_20934,N_19323,N_19111);
xor U20935 (N_20935,N_19209,N_19016);
xnor U20936 (N_20936,N_19839,N_19711);
nand U20937 (N_20937,N_19349,N_19251);
or U20938 (N_20938,N_19912,N_19132);
and U20939 (N_20939,N_19108,N_19627);
or U20940 (N_20940,N_19840,N_19548);
nand U20941 (N_20941,N_19058,N_19514);
or U20942 (N_20942,N_19426,N_19591);
nor U20943 (N_20943,N_19656,N_19685);
nor U20944 (N_20944,N_19274,N_19393);
or U20945 (N_20945,N_19465,N_19755);
or U20946 (N_20946,N_19204,N_19348);
nor U20947 (N_20947,N_19273,N_19455);
or U20948 (N_20948,N_19021,N_19075);
nor U20949 (N_20949,N_19174,N_19956);
nand U20950 (N_20950,N_19352,N_19131);
xor U20951 (N_20951,N_19034,N_19145);
nand U20952 (N_20952,N_19151,N_19998);
nand U20953 (N_20953,N_19555,N_19572);
or U20954 (N_20954,N_19355,N_19705);
and U20955 (N_20955,N_19636,N_19557);
and U20956 (N_20956,N_19614,N_19914);
nand U20957 (N_20957,N_19097,N_19130);
nand U20958 (N_20958,N_19665,N_19161);
and U20959 (N_20959,N_19576,N_19194);
nor U20960 (N_20960,N_19836,N_19896);
nand U20961 (N_20961,N_19771,N_19991);
nand U20962 (N_20962,N_19800,N_19135);
xor U20963 (N_20963,N_19008,N_19421);
and U20964 (N_20964,N_19396,N_19712);
nand U20965 (N_20965,N_19168,N_19292);
nor U20966 (N_20966,N_19565,N_19057);
xnor U20967 (N_20967,N_19304,N_19677);
nand U20968 (N_20968,N_19944,N_19235);
xor U20969 (N_20969,N_19932,N_19511);
xnor U20970 (N_20970,N_19973,N_19271);
xor U20971 (N_20971,N_19053,N_19210);
nor U20972 (N_20972,N_19506,N_19255);
nand U20973 (N_20973,N_19156,N_19036);
and U20974 (N_20974,N_19711,N_19314);
nor U20975 (N_20975,N_19029,N_19851);
nand U20976 (N_20976,N_19065,N_19684);
xnor U20977 (N_20977,N_19824,N_19122);
xnor U20978 (N_20978,N_19727,N_19762);
xor U20979 (N_20979,N_19457,N_19234);
nand U20980 (N_20980,N_19400,N_19402);
nor U20981 (N_20981,N_19886,N_19048);
xnor U20982 (N_20982,N_19498,N_19272);
nand U20983 (N_20983,N_19288,N_19038);
xor U20984 (N_20984,N_19925,N_19750);
nor U20985 (N_20985,N_19090,N_19813);
xnor U20986 (N_20986,N_19596,N_19335);
nor U20987 (N_20987,N_19442,N_19327);
and U20988 (N_20988,N_19923,N_19834);
and U20989 (N_20989,N_19370,N_19460);
nor U20990 (N_20990,N_19326,N_19120);
or U20991 (N_20991,N_19674,N_19051);
nor U20992 (N_20992,N_19165,N_19697);
xnor U20993 (N_20993,N_19950,N_19523);
or U20994 (N_20994,N_19613,N_19819);
and U20995 (N_20995,N_19642,N_19713);
and U20996 (N_20996,N_19785,N_19541);
xor U20997 (N_20997,N_19516,N_19079);
xnor U20998 (N_20998,N_19771,N_19917);
nand U20999 (N_20999,N_19310,N_19715);
nor U21000 (N_21000,N_20643,N_20217);
or U21001 (N_21001,N_20437,N_20762);
and U21002 (N_21002,N_20819,N_20603);
xnor U21003 (N_21003,N_20533,N_20035);
xor U21004 (N_21004,N_20172,N_20763);
or U21005 (N_21005,N_20992,N_20289);
and U21006 (N_21006,N_20135,N_20144);
and U21007 (N_21007,N_20474,N_20846);
xor U21008 (N_21008,N_20396,N_20337);
or U21009 (N_21009,N_20737,N_20063);
xnor U21010 (N_21010,N_20887,N_20752);
nand U21011 (N_21011,N_20236,N_20152);
nor U21012 (N_21012,N_20662,N_20939);
nor U21013 (N_21013,N_20299,N_20387);
nor U21014 (N_21014,N_20926,N_20410);
nor U21015 (N_21015,N_20491,N_20290);
nand U21016 (N_21016,N_20264,N_20528);
nor U21017 (N_21017,N_20599,N_20472);
or U21018 (N_21018,N_20419,N_20317);
xnor U21019 (N_21019,N_20739,N_20096);
xor U21020 (N_21020,N_20228,N_20732);
or U21021 (N_21021,N_20984,N_20072);
or U21022 (N_21022,N_20754,N_20532);
or U21023 (N_21023,N_20386,N_20067);
nand U21024 (N_21024,N_20481,N_20557);
or U21025 (N_21025,N_20915,N_20021);
or U21026 (N_21026,N_20475,N_20160);
nor U21027 (N_21027,N_20698,N_20354);
xnor U21028 (N_21028,N_20590,N_20831);
and U21029 (N_21029,N_20325,N_20143);
and U21030 (N_21030,N_20157,N_20880);
nor U21031 (N_21031,N_20666,N_20539);
xor U21032 (N_21032,N_20620,N_20190);
and U21033 (N_21033,N_20032,N_20787);
nand U21034 (N_21034,N_20448,N_20398);
or U21035 (N_21035,N_20037,N_20231);
and U21036 (N_21036,N_20150,N_20422);
and U21037 (N_21037,N_20045,N_20978);
and U21038 (N_21038,N_20324,N_20245);
or U21039 (N_21039,N_20464,N_20823);
or U21040 (N_21040,N_20937,N_20548);
and U21041 (N_21041,N_20495,N_20664);
and U21042 (N_21042,N_20073,N_20547);
and U21043 (N_21043,N_20965,N_20133);
nor U21044 (N_21044,N_20508,N_20641);
xor U21045 (N_21045,N_20404,N_20378);
nand U21046 (N_21046,N_20099,N_20468);
nor U21047 (N_21047,N_20928,N_20408);
xnor U21048 (N_21048,N_20027,N_20357);
nor U21049 (N_21049,N_20764,N_20889);
xor U21050 (N_21050,N_20569,N_20728);
xor U21051 (N_21051,N_20648,N_20794);
and U21052 (N_21052,N_20780,N_20991);
nor U21053 (N_21053,N_20974,N_20047);
or U21054 (N_21054,N_20114,N_20200);
nand U21055 (N_21055,N_20747,N_20761);
nor U21056 (N_21056,N_20594,N_20336);
nor U21057 (N_21057,N_20397,N_20130);
nand U21058 (N_21058,N_20403,N_20525);
nand U21059 (N_21059,N_20587,N_20914);
and U21060 (N_21060,N_20746,N_20815);
nand U21061 (N_21061,N_20103,N_20558);
or U21062 (N_21062,N_20733,N_20273);
and U21063 (N_21063,N_20729,N_20694);
xnor U21064 (N_21064,N_20607,N_20757);
xor U21065 (N_21065,N_20413,N_20486);
and U21066 (N_21066,N_20272,N_20003);
and U21067 (N_21067,N_20668,N_20283);
and U21068 (N_21068,N_20657,N_20162);
and U21069 (N_21069,N_20309,N_20682);
nand U21070 (N_21070,N_20421,N_20221);
nor U21071 (N_21071,N_20957,N_20089);
nand U21072 (N_21072,N_20541,N_20647);
nand U21073 (N_21073,N_20002,N_20189);
and U21074 (N_21074,N_20225,N_20683);
nand U21075 (N_21075,N_20675,N_20250);
xor U21076 (N_21076,N_20920,N_20768);
or U21077 (N_21077,N_20933,N_20559);
and U21078 (N_21078,N_20477,N_20756);
and U21079 (N_21079,N_20207,N_20621);
and U21080 (N_21080,N_20444,N_20543);
and U21081 (N_21081,N_20690,N_20406);
nand U21082 (N_21082,N_20750,N_20990);
xnor U21083 (N_21083,N_20791,N_20423);
nor U21084 (N_21084,N_20420,N_20490);
xnor U21085 (N_21085,N_20917,N_20237);
nand U21086 (N_21086,N_20848,N_20115);
nand U21087 (N_21087,N_20962,N_20902);
and U21088 (N_21088,N_20869,N_20196);
nor U21089 (N_21089,N_20342,N_20054);
nand U21090 (N_21090,N_20839,N_20948);
or U21091 (N_21091,N_20195,N_20348);
xor U21092 (N_21092,N_20083,N_20182);
nand U21093 (N_21093,N_20613,N_20667);
or U21094 (N_21094,N_20702,N_20604);
nor U21095 (N_21095,N_20308,N_20867);
or U21096 (N_21096,N_20463,N_20312);
and U21097 (N_21097,N_20676,N_20940);
xor U21098 (N_21098,N_20218,N_20923);
xor U21099 (N_21099,N_20895,N_20610);
nand U21100 (N_21100,N_20075,N_20986);
xnor U21101 (N_21101,N_20012,N_20435);
nor U21102 (N_21102,N_20011,N_20485);
nor U21103 (N_21103,N_20927,N_20596);
nor U21104 (N_21104,N_20153,N_20266);
nor U21105 (N_21105,N_20725,N_20802);
nand U21106 (N_21106,N_20088,N_20611);
and U21107 (N_21107,N_20456,N_20900);
and U21108 (N_21108,N_20629,N_20016);
or U21109 (N_21109,N_20222,N_20346);
nand U21110 (N_21110,N_20792,N_20241);
nor U21111 (N_21111,N_20767,N_20220);
and U21112 (N_21112,N_20110,N_20257);
nor U21113 (N_21113,N_20565,N_20977);
xor U21114 (N_21114,N_20595,N_20901);
or U21115 (N_21115,N_20051,N_20717);
nor U21116 (N_21116,N_20286,N_20042);
xor U21117 (N_21117,N_20805,N_20866);
or U21118 (N_21118,N_20136,N_20570);
nand U21119 (N_21119,N_20989,N_20310);
nor U21120 (N_21120,N_20068,N_20146);
or U21121 (N_21121,N_20947,N_20870);
xor U21122 (N_21122,N_20580,N_20740);
or U21123 (N_21123,N_20009,N_20918);
or U21124 (N_21124,N_20695,N_20686);
nand U21125 (N_21125,N_20797,N_20155);
or U21126 (N_21126,N_20279,N_20233);
xnor U21127 (N_21127,N_20632,N_20612);
and U21128 (N_21128,N_20693,N_20875);
or U21129 (N_21129,N_20362,N_20441);
nor U21130 (N_21130,N_20976,N_20333);
nor U21131 (N_21131,N_20425,N_20355);
nand U21132 (N_21132,N_20015,N_20637);
and U21133 (N_21133,N_20818,N_20820);
and U21134 (N_21134,N_20967,N_20811);
nor U21135 (N_21135,N_20727,N_20959);
nand U21136 (N_21136,N_20219,N_20391);
nor U21137 (N_21137,N_20276,N_20696);
xnor U21138 (N_21138,N_20874,N_20258);
or U21139 (N_21139,N_20714,N_20026);
or U21140 (N_21140,N_20000,N_20288);
and U21141 (N_21141,N_20365,N_20660);
xor U21142 (N_21142,N_20173,N_20784);
xor U21143 (N_21143,N_20673,N_20624);
nand U21144 (N_21144,N_20417,N_20679);
nand U21145 (N_21145,N_20092,N_20966);
and U21146 (N_21146,N_20879,N_20323);
xnor U21147 (N_21147,N_20770,N_20480);
nor U21148 (N_21148,N_20138,N_20462);
nor U21149 (N_21149,N_20007,N_20855);
or U21150 (N_21150,N_20023,N_20606);
or U21151 (N_21151,N_20314,N_20393);
xor U21152 (N_21152,N_20551,N_20809);
or U21153 (N_21153,N_20852,N_20706);
or U21154 (N_21154,N_20829,N_20185);
nand U21155 (N_21155,N_20251,N_20097);
and U21156 (N_21156,N_20450,N_20953);
and U21157 (N_21157,N_20426,N_20349);
xnor U21158 (N_21158,N_20644,N_20411);
nor U21159 (N_21159,N_20449,N_20469);
nor U21160 (N_21160,N_20996,N_20008);
or U21161 (N_21161,N_20036,N_20297);
xnor U21162 (N_21162,N_20758,N_20568);
xnor U21163 (N_21163,N_20001,N_20779);
and U21164 (N_21164,N_20566,N_20858);
and U21165 (N_21165,N_20424,N_20573);
or U21166 (N_21166,N_20141,N_20428);
nand U21167 (N_21167,N_20093,N_20341);
nand U21168 (N_21168,N_20843,N_20833);
nor U21169 (N_21169,N_20850,N_20107);
nand U21170 (N_21170,N_20244,N_20275);
or U21171 (N_21171,N_20951,N_20098);
nand U21172 (N_21172,N_20884,N_20260);
or U21173 (N_21173,N_20576,N_20102);
nand U21174 (N_21174,N_20871,N_20514);
and U21175 (N_21175,N_20512,N_20164);
nand U21176 (N_21176,N_20330,N_20210);
xnor U21177 (N_21177,N_20943,N_20363);
xor U21178 (N_21178,N_20821,N_20074);
or U21179 (N_21179,N_20436,N_20516);
or U21180 (N_21180,N_20734,N_20198);
nor U21181 (N_21181,N_20865,N_20626);
nand U21182 (N_21182,N_20513,N_20847);
nor U21183 (N_21183,N_20395,N_20432);
or U21184 (N_21184,N_20121,N_20674);
nand U21185 (N_21185,N_20502,N_20500);
xnor U21186 (N_21186,N_20771,N_20318);
nand U21187 (N_21187,N_20545,N_20139);
nor U21188 (N_21188,N_20546,N_20181);
xnor U21189 (N_21189,N_20505,N_20019);
nor U21190 (N_21190,N_20382,N_20639);
nor U21191 (N_21191,N_20375,N_20975);
xor U21192 (N_21192,N_20442,N_20439);
and U21193 (N_21193,N_20935,N_20519);
or U21194 (N_21194,N_20930,N_20520);
nor U21195 (N_21195,N_20118,N_20298);
and U21196 (N_21196,N_20854,N_20381);
and U21197 (N_21197,N_20824,N_20111);
or U21198 (N_21198,N_20095,N_20954);
or U21199 (N_21199,N_20646,N_20886);
xnor U21200 (N_21200,N_20368,N_20284);
nor U21201 (N_21201,N_20722,N_20452);
xor U21202 (N_21202,N_20161,N_20891);
and U21203 (N_21203,N_20583,N_20238);
or U21204 (N_21204,N_20535,N_20460);
nand U21205 (N_21205,N_20946,N_20215);
nor U21206 (N_21206,N_20890,N_20709);
nor U21207 (N_21207,N_20371,N_20373);
nor U21208 (N_21208,N_20229,N_20058);
nand U21209 (N_21209,N_20191,N_20904);
or U21210 (N_21210,N_20549,N_20531);
xor U21211 (N_21211,N_20090,N_20751);
or U21212 (N_21212,N_20881,N_20634);
nand U21213 (N_21213,N_20078,N_20430);
or U21214 (N_21214,N_20704,N_20744);
or U21215 (N_21215,N_20689,N_20473);
nand U21216 (N_21216,N_20672,N_20274);
xnor U21217 (N_21217,N_20384,N_20585);
nor U21218 (N_21218,N_20938,N_20394);
xnor U21219 (N_21219,N_20625,N_20159);
xnor U21220 (N_21220,N_20876,N_20069);
nor U21221 (N_21221,N_20331,N_20116);
nand U21222 (N_21222,N_20262,N_20730);
and U21223 (N_21223,N_20776,N_20555);
xnor U21224 (N_21224,N_20523,N_20239);
or U21225 (N_21225,N_20615,N_20017);
nor U21226 (N_21226,N_20801,N_20582);
and U21227 (N_21227,N_20995,N_20731);
xnor U21228 (N_21228,N_20993,N_20180);
nor U21229 (N_21229,N_20552,N_20994);
or U21230 (N_21230,N_20066,N_20235);
nor U21231 (N_21231,N_20781,N_20534);
and U21232 (N_21232,N_20131,N_20699);
or U21233 (N_21233,N_20872,N_20488);
or U21234 (N_21234,N_20489,N_20789);
and U21235 (N_21235,N_20353,N_20743);
or U21236 (N_21236,N_20671,N_20934);
nand U21237 (N_21237,N_20571,N_20705);
and U21238 (N_21238,N_20319,N_20223);
xnor U21239 (N_21239,N_20749,N_20504);
and U21240 (N_21240,N_20282,N_20214);
or U21241 (N_21241,N_20459,N_20106);
nor U21242 (N_21242,N_20014,N_20796);
or U21243 (N_21243,N_20822,N_20062);
and U21244 (N_21244,N_20484,N_20912);
xnor U21245 (N_21245,N_20574,N_20623);
or U21246 (N_21246,N_20405,N_20795);
xnor U21247 (N_21247,N_20906,N_20429);
xnor U21248 (N_21248,N_20482,N_20892);
nand U21249 (N_21249,N_20316,N_20041);
nand U21250 (N_21250,N_20772,N_20071);
nor U21251 (N_21251,N_20862,N_20140);
nand U21252 (N_21252,N_20670,N_20301);
and U21253 (N_21253,N_20203,N_20303);
or U21254 (N_21254,N_20838,N_20710);
xnor U21255 (N_21255,N_20285,N_20640);
xnor U21256 (N_21256,N_20808,N_20295);
nor U21257 (N_21257,N_20234,N_20483);
xnor U21258 (N_21258,N_20782,N_20572);
and U21259 (N_21259,N_20321,N_20005);
nor U21260 (N_21260,N_20457,N_20564);
or U21261 (N_21261,N_20493,N_20204);
xor U21262 (N_21262,N_20598,N_20038);
nand U21263 (N_21263,N_20379,N_20894);
nor U21264 (N_21264,N_20060,N_20389);
xor U21265 (N_21265,N_20911,N_20550);
nor U21266 (N_21266,N_20837,N_20560);
nand U21267 (N_21267,N_20618,N_20293);
or U21268 (N_21268,N_20878,N_20507);
nor U21269 (N_21269,N_20454,N_20307);
xnor U21270 (N_21270,N_20227,N_20803);
and U21271 (N_21271,N_20650,N_20112);
and U21272 (N_21272,N_20963,N_20170);
and U21273 (N_21273,N_20434,N_20633);
or U21274 (N_21274,N_20642,N_20628);
or U21275 (N_21275,N_20427,N_20487);
or U21276 (N_21276,N_20826,N_20703);
nand U21277 (N_21277,N_20581,N_20944);
or U21278 (N_21278,N_20154,N_20359);
xnor U21279 (N_21279,N_20498,N_20798);
or U21280 (N_21280,N_20562,N_20300);
or U21281 (N_21281,N_20151,N_20790);
nor U21282 (N_21282,N_20592,N_20137);
and U21283 (N_21283,N_20932,N_20908);
and U21284 (N_21284,N_20844,N_20941);
and U21285 (N_21285,N_20777,N_20882);
nand U21286 (N_21286,N_20503,N_20726);
nor U21287 (N_21287,N_20701,N_20385);
nor U21288 (N_21288,N_20885,N_20614);
nand U21289 (N_21289,N_20864,N_20540);
nand U21290 (N_21290,N_20294,N_20584);
or U21291 (N_21291,N_20267,N_20842);
nor U21292 (N_21292,N_20081,N_20561);
or U21293 (N_21293,N_20544,N_20313);
xnor U21294 (N_21294,N_20759,N_20192);
xnor U21295 (N_21295,N_20952,N_20329);
nand U21296 (N_21296,N_20208,N_20536);
xnor U21297 (N_21297,N_20748,N_20082);
or U21298 (N_21298,N_20471,N_20530);
nand U21299 (N_21299,N_20499,N_20388);
nand U21300 (N_21300,N_20194,N_20201);
xor U21301 (N_21301,N_20399,N_20020);
nand U21302 (N_21302,N_20183,N_20988);
nor U21303 (N_21303,N_20255,N_20120);
or U21304 (N_21304,N_20925,N_20806);
xor U21305 (N_21305,N_20997,N_20588);
nor U21306 (N_21306,N_20816,N_20972);
nor U21307 (N_21307,N_20835,N_20497);
and U21308 (N_21308,N_20352,N_20720);
or U21309 (N_21309,N_20445,N_20305);
or U21310 (N_21310,N_20999,N_20247);
or U21311 (N_21311,N_20188,N_20366);
or U21312 (N_21312,N_20440,N_20691);
and U21313 (N_21313,N_20707,N_20122);
nor U21314 (N_21314,N_20414,N_20367);
or U21315 (N_21315,N_20438,N_20268);
xor U21316 (N_21316,N_20537,N_20364);
nand U21317 (N_21317,N_20851,N_20807);
or U21318 (N_21318,N_20086,N_20246);
nor U21319 (N_21319,N_20376,N_20661);
and U21320 (N_21320,N_20609,N_20656);
and U21321 (N_21321,N_20700,N_20119);
nand U21322 (N_21322,N_20960,N_20416);
nand U21323 (N_21323,N_20360,N_20601);
nand U21324 (N_21324,N_20315,N_20374);
and U21325 (N_21325,N_20050,N_20109);
nand U21326 (N_21326,N_20226,N_20361);
xnor U21327 (N_21327,N_20248,N_20327);
or U21328 (N_21328,N_20013,N_20907);
xnor U21329 (N_21329,N_20971,N_20765);
nand U21330 (N_21330,N_20232,N_20358);
or U21331 (N_21331,N_20263,N_20048);
xor U21332 (N_21332,N_20883,N_20202);
or U21333 (N_21333,N_20921,N_20721);
xor U21334 (N_21334,N_20418,N_20024);
xnor U21335 (N_21335,N_20320,N_20735);
nand U21336 (N_21336,N_20857,N_20575);
and U21337 (N_21337,N_20335,N_20987);
and U21338 (N_21338,N_20649,N_20868);
or U21339 (N_21339,N_20903,N_20174);
and U21340 (N_21340,N_20753,N_20517);
nand U21341 (N_21341,N_20745,N_20859);
and U21342 (N_21342,N_20091,N_20949);
nand U21343 (N_21343,N_20973,N_20685);
nand U21344 (N_21344,N_20888,N_20980);
nor U21345 (N_21345,N_20893,N_20556);
or U21346 (N_21346,N_20080,N_20356);
nor U21347 (N_21347,N_20736,N_20455);
and U21348 (N_21348,N_20197,N_20981);
and U21349 (N_21349,N_20043,N_20128);
xor U21350 (N_21350,N_20810,N_20840);
xnor U21351 (N_21351,N_20783,N_20402);
or U21352 (N_21352,N_20149,N_20127);
nor U21353 (N_21353,N_20057,N_20719);
and U21354 (N_21354,N_20799,N_20898);
and U21355 (N_21355,N_20653,N_20025);
or U21356 (N_21356,N_20688,N_20018);
and U21357 (N_21357,N_20910,N_20065);
and U21358 (N_21358,N_20832,N_20304);
nor U21359 (N_21359,N_20351,N_20134);
nor U21360 (N_21360,N_20145,N_20243);
or U21361 (N_21361,N_20302,N_20800);
nor U21362 (N_21362,N_20774,N_20380);
nor U21363 (N_21363,N_20896,N_20899);
nand U21364 (N_21364,N_20863,N_20554);
and U21365 (N_21365,N_20079,N_20936);
or U21366 (N_21366,N_20028,N_20652);
xnor U21367 (N_21367,N_20982,N_20812);
or U21368 (N_21368,N_20669,N_20929);
xnor U21369 (N_21369,N_20254,N_20377);
nand U21370 (N_21370,N_20465,N_20919);
nor U21371 (N_21371,N_20958,N_20165);
nor U21372 (N_21372,N_20292,N_20658);
nor U21373 (N_21373,N_20269,N_20711);
nor U21374 (N_21374,N_20124,N_20602);
nand U21375 (N_21375,N_20775,N_20715);
nand U21376 (N_21376,N_20117,N_20281);
and U21377 (N_21377,N_20897,N_20760);
or U21378 (N_21378,N_20600,N_20004);
or U21379 (N_21379,N_20636,N_20148);
nand U21380 (N_21380,N_20061,N_20129);
xor U21381 (N_21381,N_20168,N_20296);
or U21382 (N_21382,N_20344,N_20006);
or U21383 (N_21383,N_20123,N_20586);
or U21384 (N_21384,N_20169,N_20877);
nor U21385 (N_21385,N_20224,N_20156);
or U21386 (N_21386,N_20040,N_20104);
nor U21387 (N_21387,N_20070,N_20506);
nor U21388 (N_21388,N_20950,N_20265);
nand U21389 (N_21389,N_20942,N_20212);
and U21390 (N_21390,N_20044,N_20501);
nand U21391 (N_21391,N_20521,N_20828);
nand U21392 (N_21392,N_20873,N_20338);
or U21393 (N_21393,N_20793,N_20741);
and U21394 (N_21394,N_20125,N_20627);
or U21395 (N_21395,N_20817,N_20467);
and U21396 (N_21396,N_20985,N_20479);
or U21397 (N_21397,N_20678,N_20849);
nor U21398 (N_21398,N_20446,N_20538);
and U21399 (N_21399,N_20087,N_20326);
and U21400 (N_21400,N_20515,N_20608);
nand U21401 (N_21401,N_20412,N_20022);
nand U21402 (N_21402,N_20825,N_20553);
or U21403 (N_21403,N_20055,N_20841);
and U21404 (N_21404,N_20968,N_20998);
nor U21405 (N_21405,N_20030,N_20578);
nor U21406 (N_21406,N_20913,N_20383);
nor U21407 (N_21407,N_20461,N_20617);
or U21408 (N_21408,N_20163,N_20291);
and U21409 (N_21409,N_20187,N_20814);
nor U21410 (N_21410,N_20579,N_20955);
and U21411 (N_21411,N_20659,N_20409);
xor U21412 (N_21412,N_20306,N_20259);
xnor U21413 (N_21413,N_20064,N_20242);
and U21414 (N_21414,N_20755,N_20924);
nand U21415 (N_21415,N_20970,N_20175);
or U21416 (N_21416,N_20665,N_20184);
and U21417 (N_21417,N_20813,N_20836);
nor U21418 (N_21418,N_20132,N_20638);
nor U21419 (N_21419,N_20687,N_20853);
or U21420 (N_21420,N_20094,N_20334);
xor U21421 (N_21421,N_20167,N_20697);
nand U21422 (N_21422,N_20077,N_20589);
and U21423 (N_21423,N_20723,N_20230);
and U21424 (N_21424,N_20046,N_20033);
or U21425 (N_21425,N_20769,N_20343);
and U21426 (N_21426,N_20392,N_20651);
nor U21427 (N_21427,N_20492,N_20635);
and U21428 (N_21428,N_20922,N_20252);
xnor U21429 (N_21429,N_20126,N_20773);
xor U21430 (N_21430,N_20179,N_20788);
xor U21431 (N_21431,N_20322,N_20085);
and U21432 (N_21432,N_20956,N_20390);
nand U21433 (N_21433,N_20084,N_20176);
and U21434 (N_21434,N_20655,N_20542);
nand U21435 (N_21435,N_20249,N_20861);
nor U21436 (N_21436,N_20622,N_20253);
nand U21437 (N_21437,N_20287,N_20645);
and U21438 (N_21438,N_20830,N_20328);
nor U21439 (N_21439,N_20372,N_20447);
or U21440 (N_21440,N_20415,N_20742);
and U21441 (N_21441,N_20654,N_20681);
nand U21442 (N_21442,N_20034,N_20476);
and U21443 (N_21443,N_20680,N_20478);
nor U21444 (N_21444,N_20186,N_20147);
nor U21445 (N_21445,N_20708,N_20510);
and U21446 (N_21446,N_20518,N_20010);
or U21447 (N_21447,N_20856,N_20206);
and U21448 (N_21448,N_20964,N_20280);
and U21449 (N_21449,N_20766,N_20470);
xnor U21450 (N_21450,N_20916,N_20407);
xor U21451 (N_21451,N_20270,N_20834);
nand U21452 (N_21452,N_20631,N_20527);
nand U21453 (N_21453,N_20677,N_20453);
or U21454 (N_21454,N_20433,N_20713);
xor U21455 (N_21455,N_20171,N_20577);
and U21456 (N_21456,N_20278,N_20108);
xor U21457 (N_21457,N_20692,N_20718);
and U21458 (N_21458,N_20211,N_20347);
nor U21459 (N_21459,N_20369,N_20969);
xnor U21460 (N_21460,N_20605,N_20786);
nand U21461 (N_21461,N_20804,N_20240);
nor U21462 (N_21462,N_20332,N_20261);
nor U21463 (N_21463,N_20663,N_20443);
or U21464 (N_21464,N_20738,N_20494);
xnor U21465 (N_21465,N_20039,N_20166);
xor U21466 (N_21466,N_20209,N_20716);
or U21467 (N_21467,N_20401,N_20905);
or U21468 (N_21468,N_20059,N_20961);
nor U21469 (N_21469,N_20193,N_20178);
nor U21470 (N_21470,N_20205,N_20860);
or U21471 (N_21471,N_20271,N_20076);
nor U21472 (N_21472,N_20451,N_20845);
nand U21473 (N_21473,N_20339,N_20619);
xnor U21474 (N_21474,N_20778,N_20524);
nand U21475 (N_21475,N_20256,N_20345);
or U21476 (N_21476,N_20597,N_20158);
xor U21477 (N_21477,N_20213,N_20785);
xnor U21478 (N_21478,N_20101,N_20049);
or U21479 (N_21479,N_20340,N_20522);
nor U21480 (N_21480,N_20142,N_20593);
nand U21481 (N_21481,N_20458,N_20177);
xnor U21482 (N_21482,N_20983,N_20909);
nand U21483 (N_21483,N_20056,N_20591);
nand U21484 (N_21484,N_20029,N_20526);
nor U21485 (N_21485,N_20216,N_20616);
nand U21486 (N_21486,N_20311,N_20400);
xnor U21487 (N_21487,N_20979,N_20496);
xor U21488 (N_21488,N_20724,N_20052);
or U21489 (N_21489,N_20567,N_20529);
xor U21490 (N_21490,N_20511,N_20630);
xor U21491 (N_21491,N_20945,N_20277);
nand U21492 (N_21492,N_20053,N_20509);
xor U21493 (N_21493,N_20931,N_20712);
nor U21494 (N_21494,N_20466,N_20827);
nand U21495 (N_21495,N_20370,N_20199);
and U21496 (N_21496,N_20684,N_20031);
nor U21497 (N_21497,N_20100,N_20563);
nand U21498 (N_21498,N_20105,N_20431);
or U21499 (N_21499,N_20350,N_20113);
xor U21500 (N_21500,N_20555,N_20434);
or U21501 (N_21501,N_20708,N_20857);
nand U21502 (N_21502,N_20114,N_20368);
nand U21503 (N_21503,N_20438,N_20500);
nand U21504 (N_21504,N_20329,N_20092);
or U21505 (N_21505,N_20309,N_20545);
xnor U21506 (N_21506,N_20199,N_20766);
nor U21507 (N_21507,N_20850,N_20717);
nand U21508 (N_21508,N_20970,N_20484);
nand U21509 (N_21509,N_20732,N_20328);
nand U21510 (N_21510,N_20453,N_20112);
xor U21511 (N_21511,N_20587,N_20903);
or U21512 (N_21512,N_20658,N_20073);
xnor U21513 (N_21513,N_20550,N_20471);
and U21514 (N_21514,N_20268,N_20828);
nor U21515 (N_21515,N_20022,N_20111);
or U21516 (N_21516,N_20552,N_20566);
and U21517 (N_21517,N_20418,N_20699);
nor U21518 (N_21518,N_20308,N_20520);
xor U21519 (N_21519,N_20920,N_20751);
nor U21520 (N_21520,N_20259,N_20804);
and U21521 (N_21521,N_20385,N_20110);
nor U21522 (N_21522,N_20280,N_20156);
nand U21523 (N_21523,N_20478,N_20178);
xnor U21524 (N_21524,N_20550,N_20708);
or U21525 (N_21525,N_20216,N_20502);
nor U21526 (N_21526,N_20138,N_20499);
nor U21527 (N_21527,N_20142,N_20336);
nor U21528 (N_21528,N_20738,N_20224);
or U21529 (N_21529,N_20321,N_20843);
or U21530 (N_21530,N_20265,N_20430);
nand U21531 (N_21531,N_20336,N_20373);
xor U21532 (N_21532,N_20630,N_20384);
xnor U21533 (N_21533,N_20602,N_20273);
or U21534 (N_21534,N_20772,N_20467);
nor U21535 (N_21535,N_20356,N_20769);
xor U21536 (N_21536,N_20707,N_20057);
xor U21537 (N_21537,N_20959,N_20990);
or U21538 (N_21538,N_20334,N_20936);
xnor U21539 (N_21539,N_20872,N_20990);
nand U21540 (N_21540,N_20862,N_20191);
nor U21541 (N_21541,N_20805,N_20520);
nand U21542 (N_21542,N_20843,N_20095);
nor U21543 (N_21543,N_20682,N_20768);
and U21544 (N_21544,N_20349,N_20060);
xor U21545 (N_21545,N_20142,N_20156);
xor U21546 (N_21546,N_20897,N_20912);
nor U21547 (N_21547,N_20990,N_20053);
nor U21548 (N_21548,N_20817,N_20873);
xor U21549 (N_21549,N_20871,N_20431);
nand U21550 (N_21550,N_20595,N_20854);
nand U21551 (N_21551,N_20653,N_20942);
nand U21552 (N_21552,N_20954,N_20044);
nand U21553 (N_21553,N_20926,N_20670);
or U21554 (N_21554,N_20946,N_20209);
nand U21555 (N_21555,N_20911,N_20032);
nor U21556 (N_21556,N_20059,N_20475);
nand U21557 (N_21557,N_20082,N_20352);
or U21558 (N_21558,N_20212,N_20449);
or U21559 (N_21559,N_20988,N_20244);
xnor U21560 (N_21560,N_20230,N_20867);
and U21561 (N_21561,N_20865,N_20934);
nor U21562 (N_21562,N_20865,N_20406);
nor U21563 (N_21563,N_20479,N_20422);
or U21564 (N_21564,N_20296,N_20442);
nor U21565 (N_21565,N_20823,N_20761);
nand U21566 (N_21566,N_20116,N_20447);
nor U21567 (N_21567,N_20703,N_20756);
nor U21568 (N_21568,N_20039,N_20177);
nor U21569 (N_21569,N_20578,N_20491);
nand U21570 (N_21570,N_20744,N_20573);
and U21571 (N_21571,N_20022,N_20024);
nor U21572 (N_21572,N_20740,N_20842);
nand U21573 (N_21573,N_20655,N_20427);
or U21574 (N_21574,N_20169,N_20498);
and U21575 (N_21575,N_20728,N_20072);
xnor U21576 (N_21576,N_20188,N_20282);
or U21577 (N_21577,N_20476,N_20012);
xor U21578 (N_21578,N_20124,N_20451);
nand U21579 (N_21579,N_20749,N_20323);
and U21580 (N_21580,N_20913,N_20993);
and U21581 (N_21581,N_20578,N_20659);
or U21582 (N_21582,N_20164,N_20222);
nor U21583 (N_21583,N_20323,N_20702);
nor U21584 (N_21584,N_20784,N_20688);
nand U21585 (N_21585,N_20899,N_20068);
xor U21586 (N_21586,N_20887,N_20129);
xnor U21587 (N_21587,N_20060,N_20877);
nor U21588 (N_21588,N_20418,N_20879);
nor U21589 (N_21589,N_20813,N_20585);
nand U21590 (N_21590,N_20269,N_20730);
nor U21591 (N_21591,N_20991,N_20082);
nor U21592 (N_21592,N_20816,N_20339);
or U21593 (N_21593,N_20108,N_20287);
nor U21594 (N_21594,N_20535,N_20137);
or U21595 (N_21595,N_20494,N_20035);
nor U21596 (N_21596,N_20574,N_20993);
nand U21597 (N_21597,N_20654,N_20497);
nor U21598 (N_21598,N_20485,N_20025);
nand U21599 (N_21599,N_20076,N_20504);
nand U21600 (N_21600,N_20408,N_20162);
and U21601 (N_21601,N_20314,N_20447);
nand U21602 (N_21602,N_20151,N_20651);
nand U21603 (N_21603,N_20837,N_20188);
or U21604 (N_21604,N_20906,N_20861);
and U21605 (N_21605,N_20487,N_20266);
or U21606 (N_21606,N_20687,N_20661);
and U21607 (N_21607,N_20516,N_20325);
nor U21608 (N_21608,N_20717,N_20320);
xnor U21609 (N_21609,N_20231,N_20368);
and U21610 (N_21610,N_20023,N_20625);
or U21611 (N_21611,N_20210,N_20322);
xor U21612 (N_21612,N_20073,N_20392);
xor U21613 (N_21613,N_20145,N_20052);
nor U21614 (N_21614,N_20284,N_20725);
nand U21615 (N_21615,N_20558,N_20675);
and U21616 (N_21616,N_20994,N_20194);
and U21617 (N_21617,N_20718,N_20211);
nor U21618 (N_21618,N_20484,N_20080);
nand U21619 (N_21619,N_20099,N_20679);
or U21620 (N_21620,N_20163,N_20174);
nand U21621 (N_21621,N_20302,N_20281);
nand U21622 (N_21622,N_20951,N_20136);
nand U21623 (N_21623,N_20021,N_20632);
xor U21624 (N_21624,N_20219,N_20564);
nand U21625 (N_21625,N_20062,N_20377);
xor U21626 (N_21626,N_20709,N_20086);
and U21627 (N_21627,N_20353,N_20345);
or U21628 (N_21628,N_20156,N_20194);
nor U21629 (N_21629,N_20813,N_20092);
and U21630 (N_21630,N_20105,N_20291);
or U21631 (N_21631,N_20276,N_20359);
nor U21632 (N_21632,N_20254,N_20810);
nor U21633 (N_21633,N_20349,N_20838);
nand U21634 (N_21634,N_20704,N_20745);
nand U21635 (N_21635,N_20417,N_20371);
and U21636 (N_21636,N_20782,N_20158);
nor U21637 (N_21637,N_20219,N_20624);
and U21638 (N_21638,N_20770,N_20203);
xnor U21639 (N_21639,N_20677,N_20779);
and U21640 (N_21640,N_20593,N_20087);
nor U21641 (N_21641,N_20165,N_20986);
or U21642 (N_21642,N_20076,N_20450);
xnor U21643 (N_21643,N_20783,N_20644);
or U21644 (N_21644,N_20114,N_20951);
and U21645 (N_21645,N_20449,N_20784);
or U21646 (N_21646,N_20626,N_20347);
xnor U21647 (N_21647,N_20467,N_20813);
nand U21648 (N_21648,N_20888,N_20335);
or U21649 (N_21649,N_20066,N_20044);
nor U21650 (N_21650,N_20843,N_20697);
or U21651 (N_21651,N_20523,N_20131);
and U21652 (N_21652,N_20072,N_20347);
nor U21653 (N_21653,N_20023,N_20457);
xor U21654 (N_21654,N_20918,N_20609);
xnor U21655 (N_21655,N_20728,N_20206);
xor U21656 (N_21656,N_20722,N_20790);
nor U21657 (N_21657,N_20618,N_20399);
xor U21658 (N_21658,N_20224,N_20986);
and U21659 (N_21659,N_20674,N_20521);
nand U21660 (N_21660,N_20325,N_20271);
or U21661 (N_21661,N_20844,N_20470);
and U21662 (N_21662,N_20432,N_20218);
and U21663 (N_21663,N_20866,N_20439);
nor U21664 (N_21664,N_20724,N_20642);
xor U21665 (N_21665,N_20333,N_20990);
and U21666 (N_21666,N_20012,N_20854);
or U21667 (N_21667,N_20510,N_20485);
xnor U21668 (N_21668,N_20425,N_20398);
xor U21669 (N_21669,N_20750,N_20442);
xnor U21670 (N_21670,N_20417,N_20680);
and U21671 (N_21671,N_20450,N_20865);
nand U21672 (N_21672,N_20702,N_20233);
nand U21673 (N_21673,N_20974,N_20433);
nand U21674 (N_21674,N_20416,N_20498);
xnor U21675 (N_21675,N_20343,N_20225);
nand U21676 (N_21676,N_20875,N_20393);
nand U21677 (N_21677,N_20238,N_20648);
xor U21678 (N_21678,N_20229,N_20700);
and U21679 (N_21679,N_20298,N_20996);
or U21680 (N_21680,N_20195,N_20120);
xnor U21681 (N_21681,N_20149,N_20080);
xor U21682 (N_21682,N_20594,N_20079);
xor U21683 (N_21683,N_20733,N_20403);
and U21684 (N_21684,N_20768,N_20379);
xor U21685 (N_21685,N_20037,N_20718);
nor U21686 (N_21686,N_20704,N_20054);
nand U21687 (N_21687,N_20374,N_20670);
nor U21688 (N_21688,N_20316,N_20889);
or U21689 (N_21689,N_20694,N_20481);
nor U21690 (N_21690,N_20259,N_20671);
nand U21691 (N_21691,N_20120,N_20135);
xor U21692 (N_21692,N_20631,N_20954);
and U21693 (N_21693,N_20418,N_20934);
xnor U21694 (N_21694,N_20052,N_20809);
or U21695 (N_21695,N_20517,N_20964);
nor U21696 (N_21696,N_20754,N_20868);
and U21697 (N_21697,N_20413,N_20741);
or U21698 (N_21698,N_20900,N_20489);
nor U21699 (N_21699,N_20502,N_20548);
nand U21700 (N_21700,N_20203,N_20953);
xnor U21701 (N_21701,N_20109,N_20591);
and U21702 (N_21702,N_20119,N_20948);
xor U21703 (N_21703,N_20083,N_20020);
nand U21704 (N_21704,N_20593,N_20667);
xnor U21705 (N_21705,N_20913,N_20409);
xnor U21706 (N_21706,N_20188,N_20182);
xor U21707 (N_21707,N_20090,N_20826);
xnor U21708 (N_21708,N_20488,N_20197);
or U21709 (N_21709,N_20719,N_20554);
nor U21710 (N_21710,N_20916,N_20243);
or U21711 (N_21711,N_20372,N_20195);
or U21712 (N_21712,N_20701,N_20451);
nand U21713 (N_21713,N_20612,N_20408);
nor U21714 (N_21714,N_20160,N_20348);
nor U21715 (N_21715,N_20328,N_20415);
and U21716 (N_21716,N_20904,N_20157);
nor U21717 (N_21717,N_20187,N_20092);
nor U21718 (N_21718,N_20089,N_20896);
and U21719 (N_21719,N_20293,N_20007);
or U21720 (N_21720,N_20468,N_20261);
and U21721 (N_21721,N_20500,N_20331);
and U21722 (N_21722,N_20097,N_20054);
and U21723 (N_21723,N_20433,N_20340);
nand U21724 (N_21724,N_20589,N_20773);
xor U21725 (N_21725,N_20283,N_20833);
or U21726 (N_21726,N_20372,N_20769);
and U21727 (N_21727,N_20129,N_20150);
nor U21728 (N_21728,N_20203,N_20830);
or U21729 (N_21729,N_20077,N_20491);
and U21730 (N_21730,N_20828,N_20210);
xnor U21731 (N_21731,N_20484,N_20800);
and U21732 (N_21732,N_20163,N_20376);
xor U21733 (N_21733,N_20662,N_20583);
nand U21734 (N_21734,N_20182,N_20611);
and U21735 (N_21735,N_20376,N_20850);
nor U21736 (N_21736,N_20042,N_20255);
nand U21737 (N_21737,N_20711,N_20041);
nor U21738 (N_21738,N_20839,N_20018);
nor U21739 (N_21739,N_20788,N_20562);
nand U21740 (N_21740,N_20834,N_20480);
xnor U21741 (N_21741,N_20335,N_20465);
nor U21742 (N_21742,N_20483,N_20159);
xor U21743 (N_21743,N_20180,N_20403);
nor U21744 (N_21744,N_20049,N_20010);
nand U21745 (N_21745,N_20951,N_20697);
nor U21746 (N_21746,N_20865,N_20727);
xor U21747 (N_21747,N_20358,N_20202);
or U21748 (N_21748,N_20929,N_20287);
nand U21749 (N_21749,N_20857,N_20970);
nor U21750 (N_21750,N_20340,N_20002);
or U21751 (N_21751,N_20910,N_20035);
nor U21752 (N_21752,N_20792,N_20658);
xor U21753 (N_21753,N_20410,N_20735);
and U21754 (N_21754,N_20146,N_20882);
or U21755 (N_21755,N_20166,N_20080);
and U21756 (N_21756,N_20034,N_20874);
and U21757 (N_21757,N_20792,N_20067);
and U21758 (N_21758,N_20889,N_20305);
nor U21759 (N_21759,N_20023,N_20143);
and U21760 (N_21760,N_20095,N_20036);
and U21761 (N_21761,N_20953,N_20693);
or U21762 (N_21762,N_20081,N_20696);
and U21763 (N_21763,N_20631,N_20328);
xnor U21764 (N_21764,N_20187,N_20481);
xnor U21765 (N_21765,N_20024,N_20122);
or U21766 (N_21766,N_20795,N_20934);
nor U21767 (N_21767,N_20500,N_20433);
nor U21768 (N_21768,N_20528,N_20883);
and U21769 (N_21769,N_20815,N_20759);
nand U21770 (N_21770,N_20095,N_20128);
nand U21771 (N_21771,N_20048,N_20165);
nand U21772 (N_21772,N_20394,N_20600);
nand U21773 (N_21773,N_20822,N_20922);
xor U21774 (N_21774,N_20502,N_20702);
xor U21775 (N_21775,N_20597,N_20870);
or U21776 (N_21776,N_20345,N_20596);
xor U21777 (N_21777,N_20714,N_20180);
nand U21778 (N_21778,N_20216,N_20170);
nor U21779 (N_21779,N_20650,N_20270);
xor U21780 (N_21780,N_20773,N_20377);
xnor U21781 (N_21781,N_20376,N_20269);
or U21782 (N_21782,N_20843,N_20999);
xor U21783 (N_21783,N_20684,N_20201);
nor U21784 (N_21784,N_20366,N_20617);
or U21785 (N_21785,N_20247,N_20321);
and U21786 (N_21786,N_20236,N_20862);
or U21787 (N_21787,N_20960,N_20327);
xor U21788 (N_21788,N_20293,N_20017);
nand U21789 (N_21789,N_20264,N_20466);
or U21790 (N_21790,N_20186,N_20038);
or U21791 (N_21791,N_20097,N_20480);
and U21792 (N_21792,N_20503,N_20297);
nand U21793 (N_21793,N_20731,N_20057);
xnor U21794 (N_21794,N_20540,N_20207);
and U21795 (N_21795,N_20818,N_20411);
nand U21796 (N_21796,N_20850,N_20613);
xnor U21797 (N_21797,N_20314,N_20619);
xor U21798 (N_21798,N_20613,N_20899);
and U21799 (N_21799,N_20744,N_20881);
xor U21800 (N_21800,N_20122,N_20520);
nor U21801 (N_21801,N_20392,N_20066);
nand U21802 (N_21802,N_20271,N_20061);
and U21803 (N_21803,N_20983,N_20046);
or U21804 (N_21804,N_20879,N_20517);
and U21805 (N_21805,N_20946,N_20431);
xnor U21806 (N_21806,N_20062,N_20234);
or U21807 (N_21807,N_20036,N_20141);
nand U21808 (N_21808,N_20935,N_20566);
and U21809 (N_21809,N_20079,N_20054);
nor U21810 (N_21810,N_20073,N_20526);
and U21811 (N_21811,N_20820,N_20941);
nor U21812 (N_21812,N_20962,N_20832);
nand U21813 (N_21813,N_20501,N_20839);
nand U21814 (N_21814,N_20985,N_20375);
or U21815 (N_21815,N_20493,N_20304);
nor U21816 (N_21816,N_20131,N_20748);
nand U21817 (N_21817,N_20226,N_20590);
xnor U21818 (N_21818,N_20914,N_20949);
or U21819 (N_21819,N_20488,N_20947);
xor U21820 (N_21820,N_20813,N_20665);
nand U21821 (N_21821,N_20055,N_20028);
and U21822 (N_21822,N_20053,N_20278);
xor U21823 (N_21823,N_20836,N_20211);
nand U21824 (N_21824,N_20062,N_20422);
nor U21825 (N_21825,N_20152,N_20101);
nand U21826 (N_21826,N_20742,N_20540);
nor U21827 (N_21827,N_20969,N_20640);
or U21828 (N_21828,N_20219,N_20061);
and U21829 (N_21829,N_20870,N_20004);
nand U21830 (N_21830,N_20687,N_20786);
xor U21831 (N_21831,N_20425,N_20782);
and U21832 (N_21832,N_20569,N_20578);
and U21833 (N_21833,N_20640,N_20172);
nand U21834 (N_21834,N_20896,N_20775);
xor U21835 (N_21835,N_20990,N_20408);
xor U21836 (N_21836,N_20768,N_20126);
nor U21837 (N_21837,N_20274,N_20964);
nor U21838 (N_21838,N_20795,N_20213);
or U21839 (N_21839,N_20633,N_20524);
nand U21840 (N_21840,N_20516,N_20209);
xnor U21841 (N_21841,N_20252,N_20626);
or U21842 (N_21842,N_20704,N_20614);
nor U21843 (N_21843,N_20526,N_20055);
nand U21844 (N_21844,N_20368,N_20522);
or U21845 (N_21845,N_20935,N_20989);
and U21846 (N_21846,N_20516,N_20173);
nor U21847 (N_21847,N_20557,N_20967);
and U21848 (N_21848,N_20194,N_20680);
and U21849 (N_21849,N_20828,N_20212);
nand U21850 (N_21850,N_20008,N_20897);
xor U21851 (N_21851,N_20788,N_20855);
nand U21852 (N_21852,N_20190,N_20057);
nor U21853 (N_21853,N_20745,N_20345);
xnor U21854 (N_21854,N_20747,N_20528);
and U21855 (N_21855,N_20741,N_20985);
nor U21856 (N_21856,N_20020,N_20445);
or U21857 (N_21857,N_20818,N_20341);
nor U21858 (N_21858,N_20479,N_20208);
and U21859 (N_21859,N_20501,N_20709);
nor U21860 (N_21860,N_20561,N_20583);
xor U21861 (N_21861,N_20140,N_20524);
or U21862 (N_21862,N_20754,N_20494);
nor U21863 (N_21863,N_20336,N_20239);
xor U21864 (N_21864,N_20543,N_20351);
xor U21865 (N_21865,N_20764,N_20839);
nand U21866 (N_21866,N_20023,N_20080);
xor U21867 (N_21867,N_20012,N_20656);
nand U21868 (N_21868,N_20267,N_20274);
nand U21869 (N_21869,N_20966,N_20768);
nand U21870 (N_21870,N_20058,N_20264);
xor U21871 (N_21871,N_20706,N_20202);
and U21872 (N_21872,N_20162,N_20968);
or U21873 (N_21873,N_20250,N_20498);
and U21874 (N_21874,N_20255,N_20691);
nand U21875 (N_21875,N_20149,N_20403);
nor U21876 (N_21876,N_20771,N_20944);
nor U21877 (N_21877,N_20976,N_20756);
and U21878 (N_21878,N_20767,N_20036);
or U21879 (N_21879,N_20803,N_20079);
xor U21880 (N_21880,N_20525,N_20548);
xor U21881 (N_21881,N_20618,N_20706);
nor U21882 (N_21882,N_20813,N_20732);
xor U21883 (N_21883,N_20191,N_20635);
nand U21884 (N_21884,N_20821,N_20152);
and U21885 (N_21885,N_20577,N_20187);
and U21886 (N_21886,N_20803,N_20109);
xnor U21887 (N_21887,N_20125,N_20099);
xor U21888 (N_21888,N_20602,N_20502);
nor U21889 (N_21889,N_20967,N_20029);
nand U21890 (N_21890,N_20755,N_20412);
or U21891 (N_21891,N_20337,N_20829);
xor U21892 (N_21892,N_20216,N_20619);
or U21893 (N_21893,N_20366,N_20068);
nand U21894 (N_21894,N_20197,N_20779);
or U21895 (N_21895,N_20114,N_20454);
nand U21896 (N_21896,N_20051,N_20023);
nand U21897 (N_21897,N_20150,N_20442);
or U21898 (N_21898,N_20302,N_20611);
or U21899 (N_21899,N_20850,N_20862);
nand U21900 (N_21900,N_20470,N_20997);
xnor U21901 (N_21901,N_20693,N_20498);
or U21902 (N_21902,N_20922,N_20063);
or U21903 (N_21903,N_20873,N_20936);
nor U21904 (N_21904,N_20365,N_20612);
or U21905 (N_21905,N_20498,N_20033);
xnor U21906 (N_21906,N_20388,N_20043);
and U21907 (N_21907,N_20228,N_20275);
nand U21908 (N_21908,N_20670,N_20392);
nor U21909 (N_21909,N_20787,N_20745);
nand U21910 (N_21910,N_20199,N_20795);
nand U21911 (N_21911,N_20265,N_20315);
nand U21912 (N_21912,N_20924,N_20226);
xor U21913 (N_21913,N_20711,N_20574);
xnor U21914 (N_21914,N_20800,N_20288);
or U21915 (N_21915,N_20947,N_20831);
or U21916 (N_21916,N_20680,N_20717);
and U21917 (N_21917,N_20513,N_20453);
xnor U21918 (N_21918,N_20416,N_20538);
nor U21919 (N_21919,N_20810,N_20279);
xor U21920 (N_21920,N_20024,N_20223);
or U21921 (N_21921,N_20784,N_20404);
nand U21922 (N_21922,N_20171,N_20536);
nand U21923 (N_21923,N_20546,N_20020);
and U21924 (N_21924,N_20371,N_20689);
nand U21925 (N_21925,N_20786,N_20530);
nor U21926 (N_21926,N_20627,N_20651);
xnor U21927 (N_21927,N_20579,N_20924);
xnor U21928 (N_21928,N_20180,N_20596);
and U21929 (N_21929,N_20982,N_20129);
and U21930 (N_21930,N_20885,N_20329);
and U21931 (N_21931,N_20061,N_20285);
xor U21932 (N_21932,N_20625,N_20821);
xor U21933 (N_21933,N_20428,N_20098);
xnor U21934 (N_21934,N_20320,N_20217);
and U21935 (N_21935,N_20699,N_20211);
or U21936 (N_21936,N_20373,N_20497);
nor U21937 (N_21937,N_20330,N_20003);
xor U21938 (N_21938,N_20590,N_20187);
nand U21939 (N_21939,N_20385,N_20418);
and U21940 (N_21940,N_20498,N_20708);
nor U21941 (N_21941,N_20618,N_20824);
and U21942 (N_21942,N_20982,N_20899);
or U21943 (N_21943,N_20760,N_20866);
xnor U21944 (N_21944,N_20383,N_20174);
and U21945 (N_21945,N_20714,N_20944);
nor U21946 (N_21946,N_20835,N_20331);
xnor U21947 (N_21947,N_20582,N_20533);
xor U21948 (N_21948,N_20645,N_20043);
nand U21949 (N_21949,N_20348,N_20018);
or U21950 (N_21950,N_20310,N_20939);
xnor U21951 (N_21951,N_20432,N_20104);
or U21952 (N_21952,N_20519,N_20871);
xor U21953 (N_21953,N_20616,N_20925);
or U21954 (N_21954,N_20928,N_20388);
and U21955 (N_21955,N_20696,N_20820);
or U21956 (N_21956,N_20115,N_20499);
and U21957 (N_21957,N_20901,N_20015);
and U21958 (N_21958,N_20186,N_20628);
nor U21959 (N_21959,N_20035,N_20848);
and U21960 (N_21960,N_20605,N_20780);
xor U21961 (N_21961,N_20454,N_20977);
nor U21962 (N_21962,N_20118,N_20281);
and U21963 (N_21963,N_20860,N_20714);
nand U21964 (N_21964,N_20513,N_20313);
xnor U21965 (N_21965,N_20111,N_20056);
or U21966 (N_21966,N_20392,N_20190);
and U21967 (N_21967,N_20202,N_20044);
xor U21968 (N_21968,N_20740,N_20599);
and U21969 (N_21969,N_20074,N_20023);
xor U21970 (N_21970,N_20228,N_20674);
or U21971 (N_21971,N_20307,N_20378);
nor U21972 (N_21972,N_20770,N_20412);
or U21973 (N_21973,N_20257,N_20938);
nand U21974 (N_21974,N_20342,N_20221);
nand U21975 (N_21975,N_20431,N_20962);
nand U21976 (N_21976,N_20176,N_20966);
nor U21977 (N_21977,N_20876,N_20681);
or U21978 (N_21978,N_20634,N_20783);
xnor U21979 (N_21979,N_20293,N_20208);
nand U21980 (N_21980,N_20641,N_20505);
or U21981 (N_21981,N_20558,N_20706);
or U21982 (N_21982,N_20032,N_20556);
or U21983 (N_21983,N_20748,N_20151);
xor U21984 (N_21984,N_20008,N_20851);
nor U21985 (N_21985,N_20995,N_20826);
nor U21986 (N_21986,N_20001,N_20176);
nor U21987 (N_21987,N_20970,N_20040);
xor U21988 (N_21988,N_20140,N_20184);
xor U21989 (N_21989,N_20844,N_20579);
nand U21990 (N_21990,N_20006,N_20355);
and U21991 (N_21991,N_20239,N_20377);
xor U21992 (N_21992,N_20888,N_20711);
or U21993 (N_21993,N_20169,N_20564);
nor U21994 (N_21994,N_20983,N_20332);
nand U21995 (N_21995,N_20173,N_20376);
xor U21996 (N_21996,N_20798,N_20379);
or U21997 (N_21997,N_20397,N_20515);
or U21998 (N_21998,N_20555,N_20439);
nand U21999 (N_21999,N_20307,N_20576);
or U22000 (N_22000,N_21143,N_21421);
nand U22001 (N_22001,N_21994,N_21564);
nand U22002 (N_22002,N_21612,N_21221);
nor U22003 (N_22003,N_21414,N_21529);
xor U22004 (N_22004,N_21418,N_21053);
and U22005 (N_22005,N_21307,N_21465);
nand U22006 (N_22006,N_21507,N_21736);
nand U22007 (N_22007,N_21352,N_21186);
xor U22008 (N_22008,N_21651,N_21625);
nand U22009 (N_22009,N_21109,N_21751);
xnor U22010 (N_22010,N_21572,N_21278);
or U22011 (N_22011,N_21754,N_21299);
nand U22012 (N_22012,N_21131,N_21142);
or U22013 (N_22013,N_21440,N_21865);
nor U22014 (N_22014,N_21846,N_21975);
nand U22015 (N_22015,N_21326,N_21513);
and U22016 (N_22016,N_21158,N_21796);
nor U22017 (N_22017,N_21079,N_21733);
xnor U22018 (N_22018,N_21954,N_21913);
and U22019 (N_22019,N_21303,N_21705);
xnor U22020 (N_22020,N_21607,N_21282);
nor U22021 (N_22021,N_21484,N_21939);
and U22022 (N_22022,N_21867,N_21104);
nand U22023 (N_22023,N_21187,N_21262);
and U22024 (N_22024,N_21858,N_21359);
nor U22025 (N_22025,N_21635,N_21049);
and U22026 (N_22026,N_21601,N_21811);
xor U22027 (N_22027,N_21230,N_21254);
nand U22028 (N_22028,N_21018,N_21242);
nand U22029 (N_22029,N_21401,N_21592);
and U22030 (N_22030,N_21770,N_21101);
and U22031 (N_22031,N_21068,N_21750);
or U22032 (N_22032,N_21188,N_21863);
and U22033 (N_22033,N_21845,N_21258);
xor U22034 (N_22034,N_21149,N_21100);
xor U22035 (N_22035,N_21439,N_21892);
nor U22036 (N_22036,N_21949,N_21089);
xor U22037 (N_22037,N_21585,N_21033);
or U22038 (N_22038,N_21611,N_21526);
and U22039 (N_22039,N_21971,N_21292);
nor U22040 (N_22040,N_21956,N_21017);
nor U22041 (N_22041,N_21606,N_21297);
xor U22042 (N_22042,N_21795,N_21061);
and U22043 (N_22043,N_21123,N_21725);
and U22044 (N_22044,N_21164,N_21854);
xnor U22045 (N_22045,N_21641,N_21983);
and U22046 (N_22046,N_21423,N_21191);
and U22047 (N_22047,N_21510,N_21261);
nand U22048 (N_22048,N_21807,N_21246);
xnor U22049 (N_22049,N_21429,N_21642);
nand U22050 (N_22050,N_21704,N_21316);
and U22051 (N_22051,N_21339,N_21662);
nor U22052 (N_22052,N_21509,N_21827);
and U22053 (N_22053,N_21748,N_21193);
and U22054 (N_22054,N_21372,N_21392);
xnor U22055 (N_22055,N_21095,N_21570);
nor U22056 (N_22056,N_21456,N_21235);
nand U22057 (N_22057,N_21639,N_21985);
nor U22058 (N_22058,N_21739,N_21692);
nand U22059 (N_22059,N_21217,N_21215);
or U22060 (N_22060,N_21400,N_21979);
nor U22061 (N_22061,N_21034,N_21594);
and U22062 (N_22062,N_21267,N_21765);
xor U22063 (N_22063,N_21668,N_21239);
nor U22064 (N_22064,N_21782,N_21532);
and U22065 (N_22065,N_21163,N_21669);
or U22066 (N_22066,N_21356,N_21379);
nor U22067 (N_22067,N_21703,N_21970);
or U22068 (N_22068,N_21523,N_21779);
or U22069 (N_22069,N_21296,N_21911);
and U22070 (N_22070,N_21499,N_21545);
nor U22071 (N_22071,N_21659,N_21286);
nor U22072 (N_22072,N_21551,N_21896);
or U22073 (N_22073,N_21432,N_21605);
nand U22074 (N_22074,N_21548,N_21721);
or U22075 (N_22075,N_21623,N_21218);
nor U22076 (N_22076,N_21730,N_21150);
nor U22077 (N_22077,N_21840,N_21402);
xnor U22078 (N_22078,N_21879,N_21318);
xnor U22079 (N_22079,N_21266,N_21619);
xor U22080 (N_22080,N_21055,N_21147);
or U22081 (N_22081,N_21534,N_21737);
nor U22082 (N_22082,N_21090,N_21773);
nand U22083 (N_22083,N_21944,N_21587);
nand U22084 (N_22084,N_21860,N_21153);
nor U22085 (N_22085,N_21505,N_21987);
and U22086 (N_22086,N_21032,N_21728);
or U22087 (N_22087,N_21080,N_21999);
nor U22088 (N_22088,N_21784,N_21767);
or U22089 (N_22089,N_21351,N_21675);
and U22090 (N_22090,N_21657,N_21760);
and U22091 (N_22091,N_21004,N_21341);
xnor U22092 (N_22092,N_21562,N_21916);
or U22093 (N_22093,N_21396,N_21152);
or U22094 (N_22094,N_21905,N_21161);
and U22095 (N_22095,N_21942,N_21146);
nand U22096 (N_22096,N_21539,N_21543);
or U22097 (N_22097,N_21769,N_21130);
or U22098 (N_22098,N_21009,N_21024);
nor U22099 (N_22099,N_21179,N_21696);
nand U22100 (N_22100,N_21986,N_21798);
and U22101 (N_22101,N_21457,N_21492);
and U22102 (N_22102,N_21604,N_21715);
and U22103 (N_22103,N_21415,N_21482);
and U22104 (N_22104,N_21577,N_21666);
and U22105 (N_22105,N_21849,N_21204);
or U22106 (N_22106,N_21554,N_21019);
xor U22107 (N_22107,N_21081,N_21445);
and U22108 (N_22108,N_21157,N_21788);
nand U22109 (N_22109,N_21023,N_21052);
nor U22110 (N_22110,N_21671,N_21155);
nand U22111 (N_22111,N_21225,N_21707);
or U22112 (N_22112,N_21870,N_21621);
or U22113 (N_22113,N_21294,N_21480);
and U22114 (N_22114,N_21808,N_21556);
and U22115 (N_22115,N_21399,N_21349);
or U22116 (N_22116,N_21244,N_21630);
nand U22117 (N_22117,N_21824,N_21832);
and U22118 (N_22118,N_21011,N_21139);
nand U22119 (N_22119,N_21148,N_21608);
or U22120 (N_22120,N_21342,N_21197);
or U22121 (N_22121,N_21709,N_21233);
nor U22122 (N_22122,N_21136,N_21054);
nand U22123 (N_22123,N_21462,N_21622);
or U22124 (N_22124,N_21506,N_21969);
nand U22125 (N_22125,N_21677,N_21514);
or U22126 (N_22126,N_21568,N_21794);
or U22127 (N_22127,N_21583,N_21664);
xnor U22128 (N_22128,N_21658,N_21394);
xnor U22129 (N_22129,N_21059,N_21672);
and U22130 (N_22130,N_21419,N_21466);
and U22131 (N_22131,N_21643,N_21236);
nor U22132 (N_22132,N_21243,N_21002);
and U22133 (N_22133,N_21744,N_21997);
or U22134 (N_22134,N_21718,N_21247);
nand U22135 (N_22135,N_21528,N_21648);
or U22136 (N_22136,N_21102,N_21412);
and U22137 (N_22137,N_21314,N_21459);
nor U22138 (N_22138,N_21822,N_21037);
nor U22139 (N_22139,N_21190,N_21256);
and U22140 (N_22140,N_21220,N_21135);
or U22141 (N_22141,N_21924,N_21008);
nor U22142 (N_22142,N_21404,N_21493);
nand U22143 (N_22143,N_21950,N_21159);
or U22144 (N_22144,N_21373,N_21409);
and U22145 (N_22145,N_21912,N_21154);
xor U22146 (N_22146,N_21407,N_21071);
nand U22147 (N_22147,N_21065,N_21354);
or U22148 (N_22148,N_21520,N_21460);
xor U22149 (N_22149,N_21093,N_21937);
nand U22150 (N_22150,N_21245,N_21497);
and U22151 (N_22151,N_21772,N_21042);
and U22152 (N_22152,N_21815,N_21702);
nor U22153 (N_22153,N_21603,N_21966);
and U22154 (N_22154,N_21617,N_21735);
or U22155 (N_22155,N_21681,N_21308);
xor U22156 (N_22156,N_21489,N_21477);
nor U22157 (N_22157,N_21005,N_21288);
and U22158 (N_22158,N_21108,N_21989);
nand U22159 (N_22159,N_21110,N_21063);
nor U22160 (N_22160,N_21335,N_21920);
nand U22161 (N_22161,N_21930,N_21590);
nand U22162 (N_22162,N_21348,N_21768);
or U22163 (N_22163,N_21934,N_21732);
nor U22164 (N_22164,N_21416,N_21806);
or U22165 (N_22165,N_21277,N_21380);
and U22166 (N_22166,N_21203,N_21700);
xnor U22167 (N_22167,N_21381,N_21519);
and U22168 (N_22168,N_21327,N_21302);
and U22169 (N_22169,N_21650,N_21540);
nand U22170 (N_22170,N_21250,N_21945);
nor U22171 (N_22171,N_21137,N_21022);
and U22172 (N_22172,N_21195,N_21836);
and U22173 (N_22173,N_21035,N_21649);
and U22174 (N_22174,N_21144,N_21804);
nor U22175 (N_22175,N_21676,N_21524);
nor U22176 (N_22176,N_21044,N_21763);
nand U22177 (N_22177,N_21038,N_21488);
and U22178 (N_22178,N_21813,N_21844);
xor U22179 (N_22179,N_21355,N_21084);
and U22180 (N_22180,N_21761,N_21263);
xor U22181 (N_22181,N_21753,N_21990);
or U22182 (N_22182,N_21869,N_21742);
xnor U22183 (N_22183,N_21511,N_21653);
or U22184 (N_22184,N_21550,N_21344);
or U22185 (N_22185,N_21428,N_21151);
nand U22186 (N_22186,N_21727,N_21322);
and U22187 (N_22187,N_21479,N_21178);
xnor U22188 (N_22188,N_21173,N_21198);
nand U22189 (N_22189,N_21338,N_21001);
or U22190 (N_22190,N_21450,N_21712);
or U22191 (N_22191,N_21443,N_21803);
and U22192 (N_22192,N_21336,N_21922);
and U22193 (N_22193,N_21516,N_21722);
nand U22194 (N_22194,N_21565,N_21853);
nor U22195 (N_22195,N_21695,N_21133);
nand U22196 (N_22196,N_21199,N_21817);
or U22197 (N_22197,N_21877,N_21938);
and U22198 (N_22198,N_21441,N_21571);
or U22199 (N_22199,N_21180,N_21688);
xor U22200 (N_22200,N_21743,N_21474);
nand U22201 (N_22201,N_21343,N_21051);
nor U22202 (N_22202,N_21117,N_21328);
or U22203 (N_22203,N_21376,N_21749);
nor U22204 (N_22204,N_21451,N_21923);
xnor U22205 (N_22205,N_21430,N_21114);
and U22206 (N_22206,N_21502,N_21932);
and U22207 (N_22207,N_21926,N_21325);
or U22208 (N_22208,N_21378,N_21780);
nor U22209 (N_22209,N_21775,N_21557);
and U22210 (N_22210,N_21786,N_21500);
nand U22211 (N_22211,N_21976,N_21881);
or U22212 (N_22212,N_21610,N_21495);
or U22213 (N_22213,N_21214,N_21483);
or U22214 (N_22214,N_21347,N_21275);
nand U22215 (N_22215,N_21957,N_21708);
nand U22216 (N_22216,N_21124,N_21972);
or U22217 (N_22217,N_21597,N_21251);
xor U22218 (N_22218,N_21633,N_21898);
nand U22219 (N_22219,N_21069,N_21216);
nand U22220 (N_22220,N_21961,N_21809);
nand U22221 (N_22221,N_21596,N_21627);
nand U22222 (N_22222,N_21998,N_21838);
nand U22223 (N_22223,N_21332,N_21362);
nor U22224 (N_22224,N_21876,N_21731);
nor U22225 (N_22225,N_21015,N_21016);
nor U22226 (N_22226,N_21036,N_21687);
nor U22227 (N_22227,N_21156,N_21778);
nand U22228 (N_22228,N_21360,N_21716);
or U22229 (N_22229,N_21312,N_21904);
xnor U22230 (N_22230,N_21943,N_21167);
and U22231 (N_22231,N_21050,N_21105);
or U22232 (N_22232,N_21678,N_21616);
xor U22233 (N_22233,N_21706,N_21444);
nor U22234 (N_22234,N_21914,N_21946);
and U22235 (N_22235,N_21843,N_21834);
nor U22236 (N_22236,N_21823,N_21435);
xnor U22237 (N_22237,N_21628,N_21802);
and U22238 (N_22238,N_21210,N_21206);
xor U22239 (N_22239,N_21382,N_21685);
and U22240 (N_22240,N_21406,N_21096);
or U22241 (N_22241,N_21291,N_21995);
nor U22242 (N_22242,N_21799,N_21097);
and U22243 (N_22243,N_21448,N_21007);
nor U22244 (N_22244,N_21030,N_21717);
nor U22245 (N_22245,N_21910,N_21464);
xnor U22246 (N_22246,N_21212,N_21284);
xor U22247 (N_22247,N_21965,N_21287);
nor U22248 (N_22248,N_21174,N_21257);
nand U22249 (N_22249,N_21469,N_21211);
nand U22250 (N_22250,N_21383,N_21991);
nand U22251 (N_22251,N_21968,N_21000);
nand U22252 (N_22252,N_21410,N_21313);
nor U22253 (N_22253,N_21561,N_21690);
xnor U22254 (N_22254,N_21674,N_21689);
or U22255 (N_22255,N_21405,N_21501);
or U22256 (N_22256,N_21756,N_21800);
or U22257 (N_22257,N_21933,N_21567);
and U22258 (N_22258,N_21856,N_21494);
nand U22259 (N_22259,N_21468,N_21279);
xnor U22260 (N_22260,N_21580,N_21830);
or U22261 (N_22261,N_21792,N_21029);
nor U22262 (N_22262,N_21184,N_21729);
or U22263 (N_22263,N_21334,N_21547);
and U22264 (N_22264,N_21241,N_21062);
and U22265 (N_22265,N_21602,N_21620);
nor U22266 (N_22266,N_21631,N_21390);
xor U22267 (N_22267,N_21091,N_21088);
xnor U22268 (N_22268,N_21487,N_21304);
or U22269 (N_22269,N_21172,N_21977);
nor U22270 (N_22270,N_21377,N_21569);
and U22271 (N_22271,N_21112,N_21213);
and U22272 (N_22272,N_21436,N_21848);
or U22273 (N_22273,N_21369,N_21533);
nor U22274 (N_22274,N_21544,N_21960);
and U22275 (N_22275,N_21085,N_21713);
and U22276 (N_22276,N_21560,N_21434);
nand U22277 (N_22277,N_21340,N_21886);
or U22278 (N_22278,N_21888,N_21039);
or U22279 (N_22279,N_21370,N_21320);
nor U22280 (N_22280,N_21598,N_21589);
xor U22281 (N_22281,N_21891,N_21535);
or U22282 (N_22282,N_21745,N_21363);
and U22283 (N_22283,N_21107,N_21542);
nand U22284 (N_22284,N_21652,N_21120);
nand U22285 (N_22285,N_21398,N_21295);
or U22286 (N_22286,N_21397,N_21697);
xor U22287 (N_22287,N_21227,N_21424);
nand U22288 (N_22288,N_21389,N_21058);
nand U22289 (N_22289,N_21973,N_21634);
or U22290 (N_22290,N_21422,N_21852);
xnor U22291 (N_22291,N_21259,N_21558);
nor U22292 (N_22292,N_21118,N_21070);
xor U22293 (N_22293,N_21723,N_21874);
nand U22294 (N_22294,N_21584,N_21300);
xor U22295 (N_22295,N_21955,N_21936);
and U22296 (N_22296,N_21740,N_21964);
nand U22297 (N_22297,N_21345,N_21385);
xor U22298 (N_22298,N_21637,N_21880);
nor U22299 (N_22299,N_21138,N_21305);
and U22300 (N_22300,N_21839,N_21862);
nand U22301 (N_22301,N_21981,N_21119);
or U22302 (N_22302,N_21726,N_21828);
xor U22303 (N_22303,N_21433,N_21271);
and U22304 (N_22304,N_21701,N_21208);
or U22305 (N_22305,N_21698,N_21006);
or U22306 (N_22306,N_21921,N_21940);
xnor U22307 (N_22307,N_21077,N_21546);
nand U22308 (N_22308,N_21873,N_21517);
and U22309 (N_22309,N_21591,N_21098);
or U22310 (N_22310,N_21498,N_21265);
and U22311 (N_22311,N_21762,N_21531);
or U22312 (N_22312,N_21887,N_21393);
and U22313 (N_22313,N_21982,N_21074);
nor U22314 (N_22314,N_21600,N_21319);
and U22315 (N_22315,N_21686,N_21980);
and U22316 (N_22316,N_21738,N_21638);
or U22317 (N_22317,N_21031,N_21645);
and U22318 (N_22318,N_21900,N_21951);
xor U22319 (N_22319,N_21490,N_21906);
xnor U22320 (N_22320,N_21872,N_21175);
nor U22321 (N_22321,N_21274,N_21764);
xor U22322 (N_22322,N_21057,N_21086);
xnor U22323 (N_22323,N_21826,N_21538);
xnor U22324 (N_22324,N_21272,N_21072);
xnor U22325 (N_22325,N_21895,N_21781);
xor U22326 (N_22326,N_21182,N_21614);
nor U22327 (N_22327,N_21115,N_21229);
or U22328 (N_22328,N_21021,N_21027);
and U22329 (N_22329,N_21249,N_21868);
xor U22330 (N_22330,N_21993,N_21066);
or U22331 (N_22331,N_21694,N_21812);
and U22332 (N_22332,N_21790,N_21064);
nand U22333 (N_22333,N_21927,N_21734);
nand U22334 (N_22334,N_21789,N_21438);
xnor U22335 (N_22335,N_21268,N_21446);
nand U22336 (N_22336,N_21576,N_21012);
xor U22337 (N_22337,N_21864,N_21953);
xor U22338 (N_22338,N_21329,N_21387);
nand U22339 (N_22339,N_21679,N_21646);
nor U22340 (N_22340,N_21128,N_21684);
xor U22341 (N_22341,N_21442,N_21301);
xor U22342 (N_22342,N_21427,N_21171);
nor U22343 (N_22343,N_21043,N_21842);
nand U22344 (N_22344,N_21525,N_21333);
or U22345 (N_22345,N_21908,N_21984);
nor U22346 (N_22346,N_21408,N_21388);
nand U22347 (N_22347,N_21169,N_21485);
nand U22348 (N_22348,N_21384,N_21783);
and U22349 (N_22349,N_21996,N_21632);
xor U22350 (N_22350,N_21145,N_21504);
nand U22351 (N_22351,N_21814,N_21766);
and U22352 (N_22352,N_21885,N_21831);
nand U22353 (N_22353,N_21192,N_21331);
nor U22354 (N_22354,N_21636,N_21067);
xnor U22355 (N_22355,N_21140,N_21508);
nor U22356 (N_22356,N_21231,N_21298);
nor U22357 (N_22357,N_21323,N_21897);
and U22358 (N_22358,N_21899,N_21682);
xnor U22359 (N_22359,N_21075,N_21974);
nor U22360 (N_22360,N_21890,N_21122);
xnor U22361 (N_22361,N_21988,N_21010);
and U22362 (N_22362,N_21771,N_21467);
and U22363 (N_22363,N_21094,N_21162);
xnor U22364 (N_22364,N_21805,N_21437);
xnor U22365 (N_22365,N_21575,N_21194);
nor U22366 (N_22366,N_21847,N_21087);
nand U22367 (N_22367,N_21941,N_21663);
and U22368 (N_22368,N_21473,N_21141);
and U22369 (N_22369,N_21078,N_21283);
and U22370 (N_22370,N_21395,N_21060);
xnor U22371 (N_22371,N_21720,N_21375);
and U22372 (N_22372,N_21200,N_21481);
and U22373 (N_22373,N_21579,N_21201);
xor U22374 (N_22374,N_21581,N_21586);
nor U22375 (N_22375,N_21917,N_21219);
xnor U22376 (N_22376,N_21470,N_21222);
or U22377 (N_22377,N_21290,N_21967);
nor U22378 (N_22378,N_21082,N_21458);
nand U22379 (N_22379,N_21593,N_21656);
or U22380 (N_22380,N_21963,N_21878);
nand U22381 (N_22381,N_21013,N_21699);
or U22382 (N_22382,N_21609,N_21209);
nand U22383 (N_22383,N_21915,N_21234);
and U22384 (N_22384,N_21819,N_21269);
or U22385 (N_22385,N_21264,N_21714);
xnor U22386 (N_22386,N_21431,N_21791);
or U22387 (N_22387,N_21624,N_21417);
nor U22388 (N_22388,N_21127,N_21820);
and U22389 (N_22389,N_21228,N_21240);
or U22390 (N_22390,N_21280,N_21889);
and U22391 (N_22391,N_21919,N_21574);
and U22392 (N_22392,N_21471,N_21588);
nand U22393 (N_22393,N_21541,N_21522);
nand U22394 (N_22394,N_21113,N_21857);
and U22395 (N_22395,N_21660,N_21476);
nand U22396 (N_22396,N_21902,N_21083);
nand U22397 (N_22397,N_21121,N_21613);
xor U22398 (N_22398,N_21238,N_21797);
nand U22399 (N_22399,N_21366,N_21324);
nand U22400 (N_22400,N_21045,N_21025);
xor U22401 (N_22401,N_21181,N_21909);
xor U22402 (N_22402,N_21825,N_21680);
or U22403 (N_22403,N_21403,N_21661);
nand U22404 (N_22404,N_21202,N_21183);
and U22405 (N_22405,N_21829,N_21654);
nor U22406 (N_22406,N_21670,N_21371);
xnor U22407 (N_22407,N_21177,N_21563);
and U22408 (N_22408,N_21129,N_21566);
nand U22409 (N_22409,N_21367,N_21273);
nand U22410 (N_22410,N_21665,N_21475);
nand U22411 (N_22411,N_21461,N_21205);
or U22412 (N_22412,N_21126,N_21894);
nand U22413 (N_22413,N_21170,N_21746);
or U22414 (N_22414,N_21929,N_21281);
nor U22415 (N_22415,N_21350,N_21992);
or U22416 (N_22416,N_21207,N_21306);
or U22417 (N_22417,N_21928,N_21353);
nand U22418 (N_22418,N_21472,N_21132);
nor U22419 (N_22419,N_21785,N_21232);
nand U22420 (N_22420,N_21866,N_21903);
and U22421 (N_22421,N_21463,N_21330);
or U22422 (N_22422,N_21599,N_21518);
nor U22423 (N_22423,N_21426,N_21116);
xnor U22424 (N_22424,N_21337,N_21758);
nand U22425 (N_22425,N_21673,N_21962);
or U22426 (N_22426,N_21391,N_21365);
or U22427 (N_22427,N_21253,N_21503);
nor U22428 (N_22428,N_21040,N_21189);
xor U22429 (N_22429,N_21835,N_21655);
nor U22430 (N_22430,N_21952,N_21125);
nand U22431 (N_22431,N_21449,N_21947);
xor U22432 (N_22432,N_21578,N_21226);
xor U22433 (N_22433,N_21310,N_21683);
nor U22434 (N_22434,N_21289,N_21046);
nand U22435 (N_22435,N_21752,N_21160);
and U22436 (N_22436,N_21047,N_21073);
and U22437 (N_22437,N_21901,N_21818);
xor U22438 (N_22438,N_21787,N_21759);
xnor U22439 (N_22439,N_21958,N_21048);
nand U22440 (N_22440,N_21747,N_21512);
nor U22441 (N_22441,N_21710,N_21724);
and U22442 (N_22442,N_21777,N_21014);
nand U22443 (N_22443,N_21255,N_21711);
and U22444 (N_22444,N_21134,N_21285);
and U22445 (N_22445,N_21755,N_21757);
nor U22446 (N_22446,N_21555,N_21176);
or U22447 (N_22447,N_21106,N_21931);
nand U22448 (N_22448,N_21185,N_21317);
nand U22449 (N_22449,N_21851,N_21076);
nand U22450 (N_22450,N_21311,N_21582);
or U22451 (N_22451,N_21223,N_21041);
and U22452 (N_22452,N_21358,N_21871);
xnor U22453 (N_22453,N_21850,N_21907);
or U22454 (N_22454,N_21455,N_21315);
nand U22455 (N_22455,N_21948,N_21413);
xor U22456 (N_22456,N_21276,N_21165);
nand U22457 (N_22457,N_21644,N_21893);
nand U22458 (N_22458,N_21420,N_21821);
or U22459 (N_22459,N_21810,N_21386);
xnor U22460 (N_22460,N_21361,N_21056);
xor U22461 (N_22461,N_21719,N_21452);
xnor U22462 (N_22462,N_21691,N_21270);
and U22463 (N_22463,N_21374,N_21693);
or U22464 (N_22464,N_21515,N_21553);
xor U22465 (N_22465,N_21527,N_21346);
nand U22466 (N_22466,N_21837,N_21252);
or U22467 (N_22467,N_21559,N_21092);
xor U22468 (N_22468,N_21491,N_21859);
and U22469 (N_22469,N_21959,N_21293);
xnor U22470 (N_22470,N_21486,N_21884);
xnor U22471 (N_22471,N_21935,N_21549);
xnor U22472 (N_22472,N_21168,N_21196);
or U22473 (N_22473,N_21425,N_21629);
nand U22474 (N_22474,N_21741,N_21615);
nand U22475 (N_22475,N_21595,N_21521);
xnor U22476 (N_22476,N_21793,N_21978);
nor U22477 (N_22477,N_21833,N_21855);
and U22478 (N_22478,N_21003,N_21099);
and U22479 (N_22479,N_21028,N_21454);
xor U22480 (N_22480,N_21536,N_21776);
xnor U22481 (N_22481,N_21667,N_21925);
xor U22482 (N_22482,N_21224,N_21260);
nor U22483 (N_22483,N_21411,N_21496);
nor U22484 (N_22484,N_21537,N_21573);
xor U22485 (N_22485,N_21861,N_21882);
or U22486 (N_22486,N_21364,N_21368);
or U22487 (N_22487,N_21453,N_21875);
or U22488 (N_22488,N_21626,N_21918);
nor U22489 (N_22489,N_21020,N_21103);
and U22490 (N_22490,N_21530,N_21237);
and U22491 (N_22491,N_21647,N_21309);
xor U22492 (N_22492,N_21321,N_21111);
and U22493 (N_22493,N_21841,N_21447);
or U22494 (N_22494,N_21618,N_21883);
nor U22495 (N_22495,N_21816,N_21026);
nor U22496 (N_22496,N_21640,N_21357);
xnor U22497 (N_22497,N_21552,N_21248);
nand U22498 (N_22498,N_21801,N_21478);
and U22499 (N_22499,N_21774,N_21166);
and U22500 (N_22500,N_21160,N_21083);
or U22501 (N_22501,N_21594,N_21483);
xor U22502 (N_22502,N_21749,N_21755);
xnor U22503 (N_22503,N_21960,N_21703);
nand U22504 (N_22504,N_21788,N_21155);
xnor U22505 (N_22505,N_21609,N_21073);
nand U22506 (N_22506,N_21133,N_21900);
and U22507 (N_22507,N_21276,N_21605);
and U22508 (N_22508,N_21383,N_21333);
or U22509 (N_22509,N_21261,N_21272);
nand U22510 (N_22510,N_21378,N_21801);
and U22511 (N_22511,N_21343,N_21079);
nor U22512 (N_22512,N_21469,N_21890);
or U22513 (N_22513,N_21303,N_21825);
and U22514 (N_22514,N_21785,N_21431);
and U22515 (N_22515,N_21533,N_21350);
or U22516 (N_22516,N_21594,N_21580);
nor U22517 (N_22517,N_21207,N_21215);
or U22518 (N_22518,N_21959,N_21681);
and U22519 (N_22519,N_21043,N_21071);
nor U22520 (N_22520,N_21871,N_21110);
or U22521 (N_22521,N_21124,N_21261);
nor U22522 (N_22522,N_21893,N_21823);
and U22523 (N_22523,N_21039,N_21559);
and U22524 (N_22524,N_21077,N_21213);
and U22525 (N_22525,N_21631,N_21286);
or U22526 (N_22526,N_21023,N_21376);
and U22527 (N_22527,N_21084,N_21406);
or U22528 (N_22528,N_21126,N_21747);
and U22529 (N_22529,N_21766,N_21630);
xnor U22530 (N_22530,N_21568,N_21326);
and U22531 (N_22531,N_21855,N_21066);
and U22532 (N_22532,N_21603,N_21362);
xor U22533 (N_22533,N_21321,N_21714);
xnor U22534 (N_22534,N_21183,N_21296);
nor U22535 (N_22535,N_21576,N_21685);
nand U22536 (N_22536,N_21857,N_21542);
xnor U22537 (N_22537,N_21794,N_21315);
nor U22538 (N_22538,N_21467,N_21750);
or U22539 (N_22539,N_21696,N_21207);
nor U22540 (N_22540,N_21744,N_21655);
and U22541 (N_22541,N_21472,N_21855);
nand U22542 (N_22542,N_21019,N_21216);
and U22543 (N_22543,N_21110,N_21244);
and U22544 (N_22544,N_21385,N_21605);
or U22545 (N_22545,N_21910,N_21586);
or U22546 (N_22546,N_21525,N_21942);
xor U22547 (N_22547,N_21716,N_21560);
or U22548 (N_22548,N_21407,N_21001);
nor U22549 (N_22549,N_21214,N_21519);
nor U22550 (N_22550,N_21738,N_21362);
and U22551 (N_22551,N_21219,N_21705);
and U22552 (N_22552,N_21973,N_21281);
nor U22553 (N_22553,N_21577,N_21429);
and U22554 (N_22554,N_21937,N_21297);
nor U22555 (N_22555,N_21590,N_21848);
and U22556 (N_22556,N_21911,N_21273);
nand U22557 (N_22557,N_21864,N_21520);
xor U22558 (N_22558,N_21761,N_21106);
and U22559 (N_22559,N_21443,N_21957);
nor U22560 (N_22560,N_21583,N_21980);
or U22561 (N_22561,N_21134,N_21471);
and U22562 (N_22562,N_21530,N_21075);
xnor U22563 (N_22563,N_21474,N_21043);
nand U22564 (N_22564,N_21040,N_21278);
or U22565 (N_22565,N_21708,N_21520);
xor U22566 (N_22566,N_21652,N_21803);
nand U22567 (N_22567,N_21575,N_21677);
nor U22568 (N_22568,N_21592,N_21354);
nand U22569 (N_22569,N_21693,N_21714);
and U22570 (N_22570,N_21654,N_21145);
nand U22571 (N_22571,N_21375,N_21235);
or U22572 (N_22572,N_21089,N_21935);
nand U22573 (N_22573,N_21212,N_21547);
nand U22574 (N_22574,N_21424,N_21548);
nor U22575 (N_22575,N_21677,N_21742);
and U22576 (N_22576,N_21302,N_21746);
nor U22577 (N_22577,N_21611,N_21402);
and U22578 (N_22578,N_21992,N_21035);
or U22579 (N_22579,N_21557,N_21385);
and U22580 (N_22580,N_21715,N_21118);
nand U22581 (N_22581,N_21855,N_21307);
nand U22582 (N_22582,N_21755,N_21189);
or U22583 (N_22583,N_21664,N_21515);
or U22584 (N_22584,N_21036,N_21701);
or U22585 (N_22585,N_21613,N_21658);
nor U22586 (N_22586,N_21683,N_21397);
or U22587 (N_22587,N_21185,N_21134);
nand U22588 (N_22588,N_21230,N_21389);
xor U22589 (N_22589,N_21751,N_21231);
nor U22590 (N_22590,N_21231,N_21040);
or U22591 (N_22591,N_21901,N_21042);
xnor U22592 (N_22592,N_21113,N_21462);
and U22593 (N_22593,N_21561,N_21093);
xnor U22594 (N_22594,N_21012,N_21175);
nand U22595 (N_22595,N_21524,N_21233);
nor U22596 (N_22596,N_21323,N_21887);
or U22597 (N_22597,N_21301,N_21910);
nand U22598 (N_22598,N_21924,N_21982);
xor U22599 (N_22599,N_21849,N_21569);
xor U22600 (N_22600,N_21235,N_21006);
nand U22601 (N_22601,N_21342,N_21708);
nand U22602 (N_22602,N_21756,N_21078);
and U22603 (N_22603,N_21307,N_21549);
and U22604 (N_22604,N_21450,N_21250);
nand U22605 (N_22605,N_21095,N_21524);
and U22606 (N_22606,N_21183,N_21335);
xnor U22607 (N_22607,N_21006,N_21818);
or U22608 (N_22608,N_21816,N_21566);
nand U22609 (N_22609,N_21238,N_21279);
nor U22610 (N_22610,N_21232,N_21047);
or U22611 (N_22611,N_21670,N_21896);
or U22612 (N_22612,N_21861,N_21092);
or U22613 (N_22613,N_21357,N_21124);
nor U22614 (N_22614,N_21997,N_21519);
nand U22615 (N_22615,N_21627,N_21426);
xnor U22616 (N_22616,N_21018,N_21465);
xnor U22617 (N_22617,N_21882,N_21033);
xor U22618 (N_22618,N_21302,N_21512);
and U22619 (N_22619,N_21502,N_21692);
xnor U22620 (N_22620,N_21788,N_21302);
xnor U22621 (N_22621,N_21585,N_21774);
and U22622 (N_22622,N_21227,N_21838);
or U22623 (N_22623,N_21805,N_21930);
or U22624 (N_22624,N_21074,N_21223);
or U22625 (N_22625,N_21242,N_21406);
and U22626 (N_22626,N_21120,N_21635);
nand U22627 (N_22627,N_21491,N_21431);
nand U22628 (N_22628,N_21559,N_21550);
nand U22629 (N_22629,N_21700,N_21696);
and U22630 (N_22630,N_21990,N_21335);
nor U22631 (N_22631,N_21511,N_21041);
nor U22632 (N_22632,N_21969,N_21806);
xnor U22633 (N_22633,N_21602,N_21107);
or U22634 (N_22634,N_21250,N_21464);
nand U22635 (N_22635,N_21018,N_21827);
and U22636 (N_22636,N_21836,N_21699);
nor U22637 (N_22637,N_21747,N_21023);
xor U22638 (N_22638,N_21422,N_21627);
xor U22639 (N_22639,N_21796,N_21551);
and U22640 (N_22640,N_21424,N_21312);
and U22641 (N_22641,N_21855,N_21270);
and U22642 (N_22642,N_21017,N_21229);
and U22643 (N_22643,N_21825,N_21089);
xor U22644 (N_22644,N_21653,N_21201);
or U22645 (N_22645,N_21701,N_21002);
xor U22646 (N_22646,N_21353,N_21002);
or U22647 (N_22647,N_21043,N_21112);
nor U22648 (N_22648,N_21619,N_21267);
xnor U22649 (N_22649,N_21801,N_21431);
nor U22650 (N_22650,N_21141,N_21073);
nor U22651 (N_22651,N_21377,N_21152);
or U22652 (N_22652,N_21197,N_21024);
and U22653 (N_22653,N_21433,N_21186);
nand U22654 (N_22654,N_21592,N_21788);
nor U22655 (N_22655,N_21366,N_21671);
nand U22656 (N_22656,N_21417,N_21070);
nand U22657 (N_22657,N_21103,N_21126);
nor U22658 (N_22658,N_21820,N_21148);
nand U22659 (N_22659,N_21910,N_21361);
nand U22660 (N_22660,N_21229,N_21716);
xor U22661 (N_22661,N_21640,N_21551);
nor U22662 (N_22662,N_21853,N_21650);
xor U22663 (N_22663,N_21064,N_21635);
nor U22664 (N_22664,N_21281,N_21467);
nor U22665 (N_22665,N_21166,N_21344);
and U22666 (N_22666,N_21701,N_21777);
nor U22667 (N_22667,N_21580,N_21826);
and U22668 (N_22668,N_21321,N_21592);
nor U22669 (N_22669,N_21489,N_21203);
nor U22670 (N_22670,N_21405,N_21155);
or U22671 (N_22671,N_21454,N_21366);
and U22672 (N_22672,N_21199,N_21835);
and U22673 (N_22673,N_21798,N_21839);
or U22674 (N_22674,N_21604,N_21921);
nor U22675 (N_22675,N_21617,N_21131);
xor U22676 (N_22676,N_21076,N_21992);
and U22677 (N_22677,N_21966,N_21419);
nand U22678 (N_22678,N_21365,N_21250);
or U22679 (N_22679,N_21899,N_21256);
nor U22680 (N_22680,N_21568,N_21331);
and U22681 (N_22681,N_21910,N_21102);
xnor U22682 (N_22682,N_21969,N_21523);
nand U22683 (N_22683,N_21461,N_21560);
and U22684 (N_22684,N_21745,N_21293);
xnor U22685 (N_22685,N_21778,N_21692);
or U22686 (N_22686,N_21485,N_21793);
nor U22687 (N_22687,N_21297,N_21958);
nand U22688 (N_22688,N_21763,N_21899);
nor U22689 (N_22689,N_21243,N_21506);
nand U22690 (N_22690,N_21364,N_21529);
nand U22691 (N_22691,N_21997,N_21238);
xor U22692 (N_22692,N_21109,N_21396);
xnor U22693 (N_22693,N_21331,N_21980);
and U22694 (N_22694,N_21918,N_21266);
xor U22695 (N_22695,N_21917,N_21956);
and U22696 (N_22696,N_21235,N_21088);
nand U22697 (N_22697,N_21306,N_21009);
nor U22698 (N_22698,N_21468,N_21845);
nor U22699 (N_22699,N_21450,N_21081);
and U22700 (N_22700,N_21379,N_21452);
nand U22701 (N_22701,N_21311,N_21574);
nor U22702 (N_22702,N_21850,N_21537);
nand U22703 (N_22703,N_21113,N_21720);
and U22704 (N_22704,N_21127,N_21437);
nand U22705 (N_22705,N_21799,N_21680);
nand U22706 (N_22706,N_21345,N_21021);
nand U22707 (N_22707,N_21232,N_21835);
or U22708 (N_22708,N_21507,N_21723);
or U22709 (N_22709,N_21882,N_21438);
nor U22710 (N_22710,N_21004,N_21822);
nor U22711 (N_22711,N_21348,N_21920);
and U22712 (N_22712,N_21105,N_21220);
xor U22713 (N_22713,N_21719,N_21522);
or U22714 (N_22714,N_21895,N_21837);
nand U22715 (N_22715,N_21146,N_21623);
or U22716 (N_22716,N_21404,N_21398);
or U22717 (N_22717,N_21710,N_21714);
and U22718 (N_22718,N_21612,N_21644);
nor U22719 (N_22719,N_21365,N_21774);
or U22720 (N_22720,N_21318,N_21104);
or U22721 (N_22721,N_21968,N_21048);
and U22722 (N_22722,N_21711,N_21798);
nand U22723 (N_22723,N_21175,N_21168);
nor U22724 (N_22724,N_21599,N_21306);
or U22725 (N_22725,N_21967,N_21276);
nand U22726 (N_22726,N_21907,N_21201);
or U22727 (N_22727,N_21018,N_21480);
nand U22728 (N_22728,N_21867,N_21926);
and U22729 (N_22729,N_21655,N_21910);
xnor U22730 (N_22730,N_21200,N_21864);
nor U22731 (N_22731,N_21223,N_21846);
xor U22732 (N_22732,N_21825,N_21176);
nand U22733 (N_22733,N_21540,N_21207);
nand U22734 (N_22734,N_21673,N_21718);
and U22735 (N_22735,N_21495,N_21784);
xor U22736 (N_22736,N_21625,N_21527);
xor U22737 (N_22737,N_21561,N_21040);
xnor U22738 (N_22738,N_21261,N_21447);
xor U22739 (N_22739,N_21965,N_21944);
nor U22740 (N_22740,N_21327,N_21890);
or U22741 (N_22741,N_21501,N_21813);
xnor U22742 (N_22742,N_21955,N_21398);
nand U22743 (N_22743,N_21078,N_21459);
or U22744 (N_22744,N_21256,N_21714);
xor U22745 (N_22745,N_21000,N_21903);
nand U22746 (N_22746,N_21226,N_21871);
nor U22747 (N_22747,N_21323,N_21941);
or U22748 (N_22748,N_21703,N_21627);
nor U22749 (N_22749,N_21081,N_21972);
nor U22750 (N_22750,N_21785,N_21111);
and U22751 (N_22751,N_21797,N_21652);
nor U22752 (N_22752,N_21772,N_21813);
nand U22753 (N_22753,N_21304,N_21183);
or U22754 (N_22754,N_21763,N_21828);
and U22755 (N_22755,N_21594,N_21957);
nand U22756 (N_22756,N_21849,N_21406);
nand U22757 (N_22757,N_21463,N_21601);
xnor U22758 (N_22758,N_21788,N_21446);
nor U22759 (N_22759,N_21629,N_21578);
or U22760 (N_22760,N_21240,N_21807);
nand U22761 (N_22761,N_21104,N_21426);
or U22762 (N_22762,N_21772,N_21368);
and U22763 (N_22763,N_21586,N_21129);
and U22764 (N_22764,N_21270,N_21075);
and U22765 (N_22765,N_21647,N_21728);
nand U22766 (N_22766,N_21365,N_21053);
xnor U22767 (N_22767,N_21249,N_21010);
nor U22768 (N_22768,N_21062,N_21150);
nand U22769 (N_22769,N_21556,N_21664);
nor U22770 (N_22770,N_21775,N_21357);
and U22771 (N_22771,N_21621,N_21540);
nand U22772 (N_22772,N_21632,N_21986);
nor U22773 (N_22773,N_21834,N_21659);
xor U22774 (N_22774,N_21527,N_21838);
or U22775 (N_22775,N_21336,N_21584);
and U22776 (N_22776,N_21671,N_21546);
nand U22777 (N_22777,N_21842,N_21275);
xnor U22778 (N_22778,N_21672,N_21292);
and U22779 (N_22779,N_21702,N_21092);
nor U22780 (N_22780,N_21610,N_21204);
and U22781 (N_22781,N_21462,N_21524);
or U22782 (N_22782,N_21921,N_21646);
xor U22783 (N_22783,N_21501,N_21578);
or U22784 (N_22784,N_21450,N_21749);
nand U22785 (N_22785,N_21733,N_21948);
or U22786 (N_22786,N_21936,N_21861);
and U22787 (N_22787,N_21725,N_21146);
xor U22788 (N_22788,N_21195,N_21025);
nor U22789 (N_22789,N_21517,N_21311);
and U22790 (N_22790,N_21570,N_21784);
nand U22791 (N_22791,N_21855,N_21777);
xor U22792 (N_22792,N_21403,N_21980);
and U22793 (N_22793,N_21266,N_21966);
and U22794 (N_22794,N_21681,N_21702);
nand U22795 (N_22795,N_21132,N_21077);
xnor U22796 (N_22796,N_21854,N_21146);
or U22797 (N_22797,N_21522,N_21331);
xnor U22798 (N_22798,N_21971,N_21377);
nand U22799 (N_22799,N_21956,N_21300);
nand U22800 (N_22800,N_21206,N_21041);
or U22801 (N_22801,N_21631,N_21237);
nor U22802 (N_22802,N_21587,N_21249);
or U22803 (N_22803,N_21873,N_21399);
xor U22804 (N_22804,N_21371,N_21859);
or U22805 (N_22805,N_21246,N_21255);
and U22806 (N_22806,N_21081,N_21953);
nand U22807 (N_22807,N_21697,N_21680);
nand U22808 (N_22808,N_21672,N_21567);
nor U22809 (N_22809,N_21368,N_21804);
xor U22810 (N_22810,N_21326,N_21108);
nor U22811 (N_22811,N_21924,N_21231);
nor U22812 (N_22812,N_21557,N_21034);
nand U22813 (N_22813,N_21437,N_21268);
xnor U22814 (N_22814,N_21214,N_21520);
or U22815 (N_22815,N_21519,N_21173);
and U22816 (N_22816,N_21968,N_21605);
or U22817 (N_22817,N_21576,N_21190);
nor U22818 (N_22818,N_21599,N_21989);
nor U22819 (N_22819,N_21665,N_21423);
xor U22820 (N_22820,N_21291,N_21568);
and U22821 (N_22821,N_21075,N_21291);
nand U22822 (N_22822,N_21966,N_21826);
or U22823 (N_22823,N_21056,N_21031);
and U22824 (N_22824,N_21274,N_21684);
xnor U22825 (N_22825,N_21947,N_21232);
and U22826 (N_22826,N_21787,N_21870);
and U22827 (N_22827,N_21464,N_21212);
nor U22828 (N_22828,N_21889,N_21705);
nand U22829 (N_22829,N_21101,N_21519);
xnor U22830 (N_22830,N_21791,N_21866);
or U22831 (N_22831,N_21746,N_21933);
xor U22832 (N_22832,N_21610,N_21003);
xor U22833 (N_22833,N_21935,N_21821);
nor U22834 (N_22834,N_21194,N_21111);
nor U22835 (N_22835,N_21957,N_21508);
nand U22836 (N_22836,N_21922,N_21605);
xor U22837 (N_22837,N_21513,N_21534);
xor U22838 (N_22838,N_21075,N_21090);
nand U22839 (N_22839,N_21486,N_21893);
and U22840 (N_22840,N_21652,N_21406);
nand U22841 (N_22841,N_21810,N_21966);
or U22842 (N_22842,N_21541,N_21233);
nor U22843 (N_22843,N_21348,N_21451);
nand U22844 (N_22844,N_21479,N_21844);
nor U22845 (N_22845,N_21137,N_21200);
or U22846 (N_22846,N_21072,N_21736);
and U22847 (N_22847,N_21345,N_21979);
nor U22848 (N_22848,N_21676,N_21686);
nor U22849 (N_22849,N_21309,N_21940);
and U22850 (N_22850,N_21011,N_21634);
or U22851 (N_22851,N_21029,N_21211);
nand U22852 (N_22852,N_21705,N_21594);
xnor U22853 (N_22853,N_21735,N_21248);
nand U22854 (N_22854,N_21829,N_21519);
and U22855 (N_22855,N_21950,N_21659);
nor U22856 (N_22856,N_21628,N_21201);
xnor U22857 (N_22857,N_21322,N_21464);
and U22858 (N_22858,N_21417,N_21540);
and U22859 (N_22859,N_21030,N_21673);
and U22860 (N_22860,N_21937,N_21732);
and U22861 (N_22861,N_21919,N_21928);
or U22862 (N_22862,N_21845,N_21058);
nand U22863 (N_22863,N_21637,N_21148);
nand U22864 (N_22864,N_21328,N_21963);
xnor U22865 (N_22865,N_21358,N_21779);
nor U22866 (N_22866,N_21252,N_21163);
nand U22867 (N_22867,N_21455,N_21486);
nand U22868 (N_22868,N_21958,N_21820);
xnor U22869 (N_22869,N_21949,N_21004);
or U22870 (N_22870,N_21177,N_21392);
xor U22871 (N_22871,N_21553,N_21749);
nor U22872 (N_22872,N_21415,N_21846);
nor U22873 (N_22873,N_21305,N_21805);
nand U22874 (N_22874,N_21922,N_21151);
or U22875 (N_22875,N_21770,N_21213);
nand U22876 (N_22876,N_21373,N_21712);
xor U22877 (N_22877,N_21460,N_21932);
nor U22878 (N_22878,N_21984,N_21902);
nor U22879 (N_22879,N_21867,N_21758);
xor U22880 (N_22880,N_21072,N_21448);
nor U22881 (N_22881,N_21655,N_21966);
nand U22882 (N_22882,N_21993,N_21947);
and U22883 (N_22883,N_21582,N_21942);
and U22884 (N_22884,N_21348,N_21656);
and U22885 (N_22885,N_21611,N_21270);
xnor U22886 (N_22886,N_21774,N_21035);
xor U22887 (N_22887,N_21175,N_21901);
nand U22888 (N_22888,N_21677,N_21367);
xor U22889 (N_22889,N_21543,N_21674);
nor U22890 (N_22890,N_21087,N_21426);
nand U22891 (N_22891,N_21704,N_21634);
or U22892 (N_22892,N_21982,N_21476);
or U22893 (N_22893,N_21626,N_21044);
xnor U22894 (N_22894,N_21877,N_21191);
nor U22895 (N_22895,N_21583,N_21696);
nand U22896 (N_22896,N_21146,N_21062);
or U22897 (N_22897,N_21054,N_21350);
or U22898 (N_22898,N_21903,N_21646);
or U22899 (N_22899,N_21061,N_21114);
nand U22900 (N_22900,N_21675,N_21894);
nand U22901 (N_22901,N_21816,N_21692);
nor U22902 (N_22902,N_21020,N_21779);
xnor U22903 (N_22903,N_21424,N_21380);
xor U22904 (N_22904,N_21920,N_21619);
nor U22905 (N_22905,N_21307,N_21361);
and U22906 (N_22906,N_21400,N_21449);
or U22907 (N_22907,N_21108,N_21273);
and U22908 (N_22908,N_21921,N_21398);
and U22909 (N_22909,N_21274,N_21717);
and U22910 (N_22910,N_21740,N_21647);
and U22911 (N_22911,N_21161,N_21402);
nand U22912 (N_22912,N_21011,N_21656);
xor U22913 (N_22913,N_21262,N_21459);
and U22914 (N_22914,N_21997,N_21677);
or U22915 (N_22915,N_21061,N_21621);
and U22916 (N_22916,N_21393,N_21611);
or U22917 (N_22917,N_21724,N_21259);
and U22918 (N_22918,N_21143,N_21402);
nand U22919 (N_22919,N_21218,N_21965);
nor U22920 (N_22920,N_21652,N_21798);
nor U22921 (N_22921,N_21114,N_21674);
or U22922 (N_22922,N_21589,N_21348);
nand U22923 (N_22923,N_21599,N_21750);
or U22924 (N_22924,N_21199,N_21485);
and U22925 (N_22925,N_21216,N_21374);
nand U22926 (N_22926,N_21927,N_21741);
nand U22927 (N_22927,N_21966,N_21931);
xnor U22928 (N_22928,N_21214,N_21547);
xor U22929 (N_22929,N_21001,N_21409);
nand U22930 (N_22930,N_21980,N_21036);
nor U22931 (N_22931,N_21862,N_21754);
xor U22932 (N_22932,N_21350,N_21843);
nand U22933 (N_22933,N_21910,N_21357);
and U22934 (N_22934,N_21100,N_21495);
or U22935 (N_22935,N_21083,N_21657);
or U22936 (N_22936,N_21472,N_21329);
xnor U22937 (N_22937,N_21065,N_21680);
nor U22938 (N_22938,N_21051,N_21454);
or U22939 (N_22939,N_21599,N_21670);
or U22940 (N_22940,N_21556,N_21923);
or U22941 (N_22941,N_21290,N_21180);
and U22942 (N_22942,N_21431,N_21617);
nor U22943 (N_22943,N_21084,N_21798);
xor U22944 (N_22944,N_21145,N_21768);
or U22945 (N_22945,N_21226,N_21213);
or U22946 (N_22946,N_21208,N_21255);
xnor U22947 (N_22947,N_21453,N_21202);
nand U22948 (N_22948,N_21841,N_21803);
nand U22949 (N_22949,N_21492,N_21626);
xnor U22950 (N_22950,N_21071,N_21408);
and U22951 (N_22951,N_21333,N_21255);
or U22952 (N_22952,N_21498,N_21760);
nor U22953 (N_22953,N_21926,N_21521);
nand U22954 (N_22954,N_21338,N_21253);
or U22955 (N_22955,N_21499,N_21025);
xor U22956 (N_22956,N_21855,N_21935);
nor U22957 (N_22957,N_21365,N_21045);
nand U22958 (N_22958,N_21031,N_21921);
nor U22959 (N_22959,N_21733,N_21810);
and U22960 (N_22960,N_21215,N_21965);
and U22961 (N_22961,N_21127,N_21791);
or U22962 (N_22962,N_21880,N_21337);
xor U22963 (N_22963,N_21090,N_21540);
or U22964 (N_22964,N_21557,N_21462);
nand U22965 (N_22965,N_21484,N_21566);
nor U22966 (N_22966,N_21859,N_21467);
xnor U22967 (N_22967,N_21489,N_21453);
nand U22968 (N_22968,N_21986,N_21831);
and U22969 (N_22969,N_21880,N_21175);
nand U22970 (N_22970,N_21662,N_21873);
nand U22971 (N_22971,N_21489,N_21743);
or U22972 (N_22972,N_21097,N_21994);
or U22973 (N_22973,N_21084,N_21936);
and U22974 (N_22974,N_21790,N_21438);
nand U22975 (N_22975,N_21326,N_21867);
nand U22976 (N_22976,N_21996,N_21283);
or U22977 (N_22977,N_21890,N_21781);
xor U22978 (N_22978,N_21452,N_21858);
and U22979 (N_22979,N_21369,N_21838);
xor U22980 (N_22980,N_21333,N_21474);
xnor U22981 (N_22981,N_21632,N_21660);
and U22982 (N_22982,N_21660,N_21408);
or U22983 (N_22983,N_21637,N_21371);
xnor U22984 (N_22984,N_21512,N_21242);
nor U22985 (N_22985,N_21254,N_21959);
and U22986 (N_22986,N_21927,N_21040);
and U22987 (N_22987,N_21275,N_21788);
nand U22988 (N_22988,N_21695,N_21664);
nor U22989 (N_22989,N_21185,N_21218);
and U22990 (N_22990,N_21931,N_21727);
nand U22991 (N_22991,N_21086,N_21205);
or U22992 (N_22992,N_21786,N_21884);
nand U22993 (N_22993,N_21606,N_21892);
nor U22994 (N_22994,N_21874,N_21603);
nor U22995 (N_22995,N_21104,N_21099);
nor U22996 (N_22996,N_21859,N_21416);
or U22997 (N_22997,N_21753,N_21739);
or U22998 (N_22998,N_21470,N_21460);
and U22999 (N_22999,N_21405,N_21164);
nand U23000 (N_23000,N_22224,N_22027);
or U23001 (N_23001,N_22333,N_22215);
xnor U23002 (N_23002,N_22855,N_22069);
and U23003 (N_23003,N_22595,N_22908);
nor U23004 (N_23004,N_22928,N_22718);
xor U23005 (N_23005,N_22948,N_22457);
xor U23006 (N_23006,N_22467,N_22829);
and U23007 (N_23007,N_22906,N_22754);
xor U23008 (N_23008,N_22346,N_22656);
and U23009 (N_23009,N_22678,N_22544);
xor U23010 (N_23010,N_22214,N_22440);
nor U23011 (N_23011,N_22784,N_22419);
nor U23012 (N_23012,N_22615,N_22771);
nand U23013 (N_23013,N_22063,N_22223);
or U23014 (N_23014,N_22597,N_22205);
or U23015 (N_23015,N_22587,N_22760);
or U23016 (N_23016,N_22222,N_22947);
nor U23017 (N_23017,N_22722,N_22283);
nand U23018 (N_23018,N_22688,N_22233);
or U23019 (N_23019,N_22669,N_22000);
nand U23020 (N_23020,N_22549,N_22163);
or U23021 (N_23021,N_22073,N_22972);
or U23022 (N_23022,N_22125,N_22823);
or U23023 (N_23023,N_22251,N_22909);
nand U23024 (N_23024,N_22904,N_22853);
nand U23025 (N_23025,N_22149,N_22141);
or U23026 (N_23026,N_22681,N_22262);
xor U23027 (N_23027,N_22422,N_22007);
and U23028 (N_23028,N_22323,N_22389);
xnor U23029 (N_23029,N_22401,N_22193);
nor U23030 (N_23030,N_22914,N_22324);
xnor U23031 (N_23031,N_22824,N_22484);
nor U23032 (N_23032,N_22242,N_22386);
or U23033 (N_23033,N_22311,N_22394);
xor U23034 (N_23034,N_22245,N_22710);
nand U23035 (N_23035,N_22835,N_22209);
nor U23036 (N_23036,N_22429,N_22685);
or U23037 (N_23037,N_22156,N_22028);
and U23038 (N_23038,N_22858,N_22620);
nand U23039 (N_23039,N_22190,N_22146);
nand U23040 (N_23040,N_22505,N_22658);
nand U23041 (N_23041,N_22815,N_22511);
xnor U23042 (N_23042,N_22319,N_22566);
nor U23043 (N_23043,N_22109,N_22409);
xnor U23044 (N_23044,N_22420,N_22257);
or U23045 (N_23045,N_22499,N_22139);
nand U23046 (N_23046,N_22961,N_22150);
nor U23047 (N_23047,N_22536,N_22955);
or U23048 (N_23048,N_22020,N_22956);
and U23049 (N_23049,N_22236,N_22160);
xor U23050 (N_23050,N_22811,N_22776);
and U23051 (N_23051,N_22520,N_22080);
nand U23052 (N_23052,N_22513,N_22260);
and U23053 (N_23053,N_22714,N_22134);
nor U23054 (N_23054,N_22300,N_22807);
or U23055 (N_23055,N_22765,N_22644);
and U23056 (N_23056,N_22833,N_22465);
xor U23057 (N_23057,N_22295,N_22808);
or U23058 (N_23058,N_22350,N_22062);
nand U23059 (N_23059,N_22294,N_22810);
and U23060 (N_23060,N_22702,N_22272);
nand U23061 (N_23061,N_22194,N_22869);
and U23062 (N_23062,N_22660,N_22453);
or U23063 (N_23063,N_22543,N_22009);
nor U23064 (N_23064,N_22426,N_22208);
and U23065 (N_23065,N_22524,N_22458);
or U23066 (N_23066,N_22200,N_22528);
nor U23067 (N_23067,N_22761,N_22100);
nand U23068 (N_23068,N_22753,N_22554);
nor U23069 (N_23069,N_22079,N_22423);
nand U23070 (N_23070,N_22362,N_22527);
xor U23071 (N_23071,N_22495,N_22220);
and U23072 (N_23072,N_22131,N_22707);
nand U23073 (N_23073,N_22946,N_22469);
nand U23074 (N_23074,N_22621,N_22694);
nor U23075 (N_23075,N_22567,N_22048);
or U23076 (N_23076,N_22535,N_22483);
or U23077 (N_23077,N_22992,N_22856);
and U23078 (N_23078,N_22332,N_22668);
or U23079 (N_23079,N_22170,N_22632);
xor U23080 (N_23080,N_22176,N_22530);
nand U23081 (N_23081,N_22274,N_22343);
nor U23082 (N_23082,N_22951,N_22548);
and U23083 (N_23083,N_22023,N_22894);
xor U23084 (N_23084,N_22296,N_22518);
or U23085 (N_23085,N_22128,N_22437);
nor U23086 (N_23086,N_22625,N_22025);
and U23087 (N_23087,N_22591,N_22608);
and U23088 (N_23088,N_22731,N_22960);
or U23089 (N_23089,N_22327,N_22845);
nand U23090 (N_23090,N_22634,N_22459);
xnor U23091 (N_23091,N_22110,N_22657);
xnor U23092 (N_23092,N_22162,N_22269);
nand U23093 (N_23093,N_22684,N_22144);
xor U23094 (N_23094,N_22305,N_22925);
and U23095 (N_23095,N_22261,N_22596);
and U23096 (N_23096,N_22979,N_22649);
nor U23097 (N_23097,N_22837,N_22574);
xnor U23098 (N_23098,N_22971,N_22341);
nor U23099 (N_23099,N_22339,N_22742);
and U23100 (N_23100,N_22034,N_22569);
or U23101 (N_23101,N_22646,N_22121);
nand U23102 (N_23102,N_22042,N_22123);
nor U23103 (N_23103,N_22801,N_22501);
and U23104 (N_23104,N_22576,N_22770);
or U23105 (N_23105,N_22817,N_22772);
and U23106 (N_23106,N_22637,N_22442);
nand U23107 (N_23107,N_22861,N_22425);
and U23108 (N_23108,N_22575,N_22699);
nand U23109 (N_23109,N_22828,N_22896);
nand U23110 (N_23110,N_22325,N_22840);
xor U23111 (N_23111,N_22502,N_22541);
and U23112 (N_23112,N_22822,N_22049);
xnor U23113 (N_23113,N_22174,N_22945);
nor U23114 (N_23114,N_22161,N_22439);
xor U23115 (N_23115,N_22151,N_22578);
nor U23116 (N_23116,N_22225,N_22903);
or U23117 (N_23117,N_22913,N_22201);
nand U23118 (N_23118,N_22169,N_22729);
nor U23119 (N_23119,N_22723,N_22304);
or U23120 (N_23120,N_22598,N_22240);
xnor U23121 (N_23121,N_22370,N_22766);
and U23122 (N_23122,N_22338,N_22683);
nor U23123 (N_23123,N_22806,N_22747);
and U23124 (N_23124,N_22187,N_22143);
nor U23125 (N_23125,N_22740,N_22147);
nand U23126 (N_23126,N_22171,N_22568);
or U23127 (N_23127,N_22538,N_22796);
and U23128 (N_23128,N_22210,N_22455);
and U23129 (N_23129,N_22302,N_22044);
nor U23130 (N_23130,N_22217,N_22583);
nand U23131 (N_23131,N_22291,N_22166);
xnor U23132 (N_23132,N_22129,N_22068);
nand U23133 (N_23133,N_22852,N_22763);
nor U23134 (N_23134,N_22012,N_22870);
nand U23135 (N_23135,N_22461,N_22846);
nor U23136 (N_23136,N_22529,N_22076);
nand U23137 (N_23137,N_22004,N_22509);
nor U23138 (N_23138,N_22085,N_22117);
or U23139 (N_23139,N_22911,N_22375);
and U23140 (N_23140,N_22749,N_22376);
or U23141 (N_23141,N_22396,N_22552);
and U23142 (N_23142,N_22417,N_22586);
nor U23143 (N_23143,N_22329,N_22851);
nor U23144 (N_23144,N_22135,N_22863);
xor U23145 (N_23145,N_22067,N_22017);
and U23146 (N_23146,N_22919,N_22441);
nand U23147 (N_23147,N_22235,N_22336);
and U23148 (N_23148,N_22473,N_22739);
xor U23149 (N_23149,N_22964,N_22958);
xnor U23150 (N_23150,N_22609,N_22504);
or U23151 (N_23151,N_22087,N_22016);
nor U23152 (N_23152,N_22516,N_22307);
nor U23153 (N_23153,N_22859,N_22299);
and U23154 (N_23154,N_22178,N_22700);
nor U23155 (N_23155,N_22256,N_22590);
nand U23156 (N_23156,N_22561,N_22271);
nand U23157 (N_23157,N_22039,N_22650);
and U23158 (N_23158,N_22558,N_22485);
and U23159 (N_23159,N_22345,N_22814);
nand U23160 (N_23160,N_22140,N_22547);
nand U23161 (N_23161,N_22987,N_22954);
nor U23162 (N_23162,N_22581,N_22728);
or U23163 (N_23163,N_22359,N_22643);
or U23164 (N_23164,N_22154,N_22885);
nor U23165 (N_23165,N_22092,N_22713);
and U23166 (N_23166,N_22616,N_22799);
nand U23167 (N_23167,N_22317,N_22435);
nand U23168 (N_23168,N_22978,N_22999);
and U23169 (N_23169,N_22779,N_22112);
nand U23170 (N_23170,N_22309,N_22560);
xnor U23171 (N_23171,N_22892,N_22358);
and U23172 (N_23172,N_22626,N_22284);
or U23173 (N_23173,N_22876,N_22145);
nor U23174 (N_23174,N_22670,N_22265);
xnor U23175 (N_23175,N_22631,N_22617);
xnor U23176 (N_23176,N_22137,N_22349);
or U23177 (N_23177,N_22180,N_22230);
xor U23178 (N_23178,N_22579,N_22897);
or U23179 (N_23179,N_22403,N_22095);
nand U23180 (N_23180,N_22752,N_22910);
nor U23181 (N_23181,N_22456,N_22996);
or U23182 (N_23182,N_22748,N_22288);
nand U23183 (N_23183,N_22083,N_22794);
nand U23184 (N_23184,N_22895,N_22041);
nand U23185 (N_23185,N_22891,N_22689);
xor U23186 (N_23186,N_22081,N_22893);
xor U23187 (N_23187,N_22104,N_22988);
or U23188 (N_23188,N_22111,N_22267);
nand U23189 (N_23189,N_22704,N_22599);
nor U23190 (N_23190,N_22189,N_22737);
nand U23191 (N_23191,N_22692,N_22244);
nand U23192 (N_23192,N_22900,N_22537);
nor U23193 (N_23193,N_22031,N_22680);
or U23194 (N_23194,N_22246,N_22387);
and U23195 (N_23195,N_22279,N_22384);
or U23196 (N_23196,N_22877,N_22102);
nand U23197 (N_23197,N_22418,N_22724);
nor U23198 (N_23198,N_22330,N_22727);
xor U23199 (N_23199,N_22270,N_22654);
nand U23200 (N_23200,N_22533,N_22834);
xor U23201 (N_23201,N_22777,N_22402);
xor U23202 (N_23202,N_22313,N_22405);
xor U23203 (N_23203,N_22421,N_22424);
xor U23204 (N_23204,N_22404,N_22787);
or U23205 (N_23205,N_22515,N_22212);
or U23206 (N_23206,N_22377,N_22975);
or U23207 (N_23207,N_22570,N_22002);
nand U23208 (N_23208,N_22821,N_22610);
or U23209 (N_23209,N_22046,N_22397);
or U23210 (N_23210,N_22671,N_22758);
nor U23211 (N_23211,N_22697,N_22995);
and U23212 (N_23212,N_22226,N_22114);
nor U23213 (N_23213,N_22239,N_22152);
nand U23214 (N_23214,N_22780,N_22640);
or U23215 (N_23215,N_22953,N_22013);
nor U23216 (N_23216,N_22196,N_22592);
xnor U23217 (N_23217,N_22015,N_22665);
xor U23218 (N_23218,N_22247,N_22611);
or U23219 (N_23219,N_22372,N_22472);
and U23220 (N_23220,N_22380,N_22540);
or U23221 (N_23221,N_22857,N_22746);
xnor U23222 (N_23222,N_22872,N_22287);
nand U23223 (N_23223,N_22559,N_22292);
nand U23224 (N_23224,N_22407,N_22355);
or U23225 (N_23225,N_22084,N_22091);
and U23226 (N_23226,N_22335,N_22053);
and U23227 (N_23227,N_22446,N_22211);
nand U23228 (N_23228,N_22912,N_22966);
xor U23229 (N_23229,N_22985,N_22508);
nor U23230 (N_23230,N_22229,N_22221);
xor U23231 (N_23231,N_22917,N_22243);
or U23232 (N_23232,N_22738,N_22254);
or U23233 (N_23233,N_22652,N_22078);
nand U23234 (N_23234,N_22594,N_22098);
xor U23235 (N_23235,N_22001,N_22445);
and U23236 (N_23236,N_22734,N_22628);
nand U23237 (N_23237,N_22471,N_22874);
nand U23238 (N_23238,N_22744,N_22696);
or U23239 (N_23239,N_22664,N_22320);
and U23240 (N_23240,N_22118,N_22382);
nand U23241 (N_23241,N_22416,N_22839);
xor U23242 (N_23242,N_22769,N_22119);
nor U23243 (N_23243,N_22641,N_22238);
nor U23244 (N_23244,N_22600,N_22477);
nand U23245 (N_23245,N_22542,N_22414);
and U23246 (N_23246,N_22818,N_22767);
nand U23247 (N_23247,N_22133,N_22488);
xor U23248 (N_23248,N_22865,N_22089);
and U23249 (N_23249,N_22186,N_22191);
or U23250 (N_23250,N_22730,N_22630);
xnor U23251 (N_23251,N_22969,N_22662);
nor U23252 (N_23252,N_22916,N_22981);
or U23253 (N_23253,N_22035,N_22127);
nor U23254 (N_23254,N_22056,N_22237);
nor U23255 (N_23255,N_22344,N_22967);
xor U23256 (N_23256,N_22973,N_22682);
and U23257 (N_23257,N_22331,N_22388);
and U23258 (N_23258,N_22733,N_22410);
xnor U23259 (N_23259,N_22907,N_22651);
and U23260 (N_23260,N_22462,N_22082);
nand U23261 (N_23261,N_22805,N_22116);
or U23262 (N_23262,N_22014,N_22820);
nand U23263 (N_23263,N_22902,N_22565);
xor U23264 (N_23264,N_22385,N_22666);
nand U23265 (N_23265,N_22164,N_22334);
or U23266 (N_23266,N_22593,N_22352);
xor U23267 (N_23267,N_22905,N_22580);
and U23268 (N_23268,N_22496,N_22860);
nand U23269 (N_23269,N_22873,N_22275);
or U23270 (N_23270,N_22108,N_22363);
nor U23271 (N_23271,N_22921,N_22366);
nor U23272 (N_23272,N_22183,N_22959);
or U23273 (N_23273,N_22875,N_22572);
nor U23274 (N_23274,N_22539,N_22785);
nand U23275 (N_23275,N_22064,N_22519);
nor U23276 (N_23276,N_22065,N_22368);
nand U23277 (N_23277,N_22965,N_22957);
nand U23278 (N_23278,N_22698,N_22526);
and U23279 (N_23279,N_22880,N_22510);
and U23280 (N_23280,N_22466,N_22413);
xor U23281 (N_23281,N_22107,N_22029);
xor U23282 (N_23282,N_22854,N_22686);
nor U23283 (N_23283,N_22940,N_22500);
and U23284 (N_23284,N_22094,N_22058);
or U23285 (N_23285,N_22057,N_22126);
xor U23286 (N_23286,N_22241,N_22447);
and U23287 (N_23287,N_22032,N_22216);
xnor U23288 (N_23288,N_22663,N_22918);
or U23289 (N_23289,N_22797,N_22390);
xor U23290 (N_23290,N_22920,N_22286);
or U23291 (N_23291,N_22434,N_22795);
or U23292 (N_23292,N_22026,N_22938);
or U23293 (N_23293,N_22054,N_22899);
nor U23294 (N_23294,N_22010,N_22360);
xor U23295 (N_23295,N_22451,N_22395);
nand U23296 (N_23296,N_22514,N_22888);
nand U23297 (N_23297,N_22635,N_22939);
or U23298 (N_23298,N_22438,N_22648);
and U23299 (N_23299,N_22103,N_22369);
and U23300 (N_23300,N_22507,N_22427);
nand U23301 (N_23301,N_22653,N_22148);
nand U23302 (N_23302,N_22970,N_22712);
nor U23303 (N_23303,N_22105,N_22399);
xor U23304 (N_23304,N_22639,N_22884);
and U23305 (N_23305,N_22862,N_22984);
nor U23306 (N_23306,N_22901,N_22177);
xor U23307 (N_23307,N_22312,N_22843);
nor U23308 (N_23308,N_22470,N_22400);
nand U23309 (N_23309,N_22249,N_22778);
xor U23310 (N_23310,N_22924,N_22636);
and U23311 (N_23311,N_22551,N_22142);
nand U23312 (N_23312,N_22603,N_22476);
xnor U23313 (N_23313,N_22927,N_22800);
and U23314 (N_23314,N_22555,N_22252);
or U23315 (N_23315,N_22881,N_22097);
nand U23316 (N_23316,N_22167,N_22463);
xnor U23317 (N_23317,N_22130,N_22037);
nand U23318 (N_23318,N_22695,N_22491);
or U23319 (N_23319,N_22564,N_22813);
nor U23320 (N_23320,N_22759,N_22454);
or U23321 (N_23321,N_22364,N_22645);
or U23322 (N_23322,N_22199,N_22301);
and U23323 (N_23323,N_22351,N_22448);
and U23324 (N_23324,N_22706,N_22675);
nor U23325 (N_23325,N_22303,N_22922);
nand U23326 (N_23326,N_22314,N_22179);
nor U23327 (N_23327,N_22676,N_22848);
and U23328 (N_23328,N_22589,N_22803);
and U23329 (N_23329,N_22659,N_22991);
xor U23330 (N_23330,N_22354,N_22480);
nand U23331 (N_23331,N_22864,N_22406);
xnor U23332 (N_23332,N_22931,N_22842);
nand U23333 (N_23333,N_22941,N_22687);
or U23334 (N_23334,N_22379,N_22673);
nor U23335 (N_23335,N_22512,N_22337);
xor U23336 (N_23336,N_22408,N_22725);
and U23337 (N_23337,N_22571,N_22207);
and U23338 (N_23338,N_22195,N_22949);
and U23339 (N_23339,N_22879,N_22976);
xnor U23340 (N_23340,N_22036,N_22674);
and U23341 (N_23341,N_22124,N_22228);
or U23342 (N_23342,N_22577,N_22915);
xor U23343 (N_23343,N_22158,N_22415);
and U23344 (N_23344,N_22202,N_22318);
xor U23345 (N_23345,N_22277,N_22944);
or U23346 (N_23346,N_22051,N_22047);
nor U23347 (N_23347,N_22443,N_22647);
xnor U23348 (N_23348,N_22968,N_22997);
nor U23349 (N_23349,N_22072,N_22613);
or U23350 (N_23350,N_22173,N_22113);
nor U23351 (N_23351,N_22096,N_22077);
and U23352 (N_23352,N_22232,N_22120);
nor U23353 (N_23353,N_22218,N_22619);
nor U23354 (N_23354,N_22937,N_22452);
or U23355 (N_23355,N_22071,N_22980);
xor U23356 (N_23356,N_22638,N_22726);
nand U23357 (N_23357,N_22280,N_22285);
xnor U23358 (N_23358,N_22773,N_22234);
and U23359 (N_23359,N_22030,N_22720);
and U23360 (N_23360,N_22255,N_22790);
nor U23361 (N_23361,N_22523,N_22106);
xor U23362 (N_23362,N_22736,N_22006);
nor U23363 (N_23363,N_22889,N_22310);
or U23364 (N_23364,N_22460,N_22008);
xor U23365 (N_23365,N_22622,N_22812);
xor U23366 (N_23366,N_22521,N_22849);
nand U23367 (N_23367,N_22498,N_22172);
xor U23368 (N_23368,N_22708,N_22490);
nor U23369 (N_23369,N_22990,N_22011);
nand U23370 (N_23370,N_22836,N_22690);
xnor U23371 (N_23371,N_22021,N_22101);
xor U23372 (N_23372,N_22074,N_22175);
and U23373 (N_23373,N_22867,N_22316);
or U23374 (N_23374,N_22293,N_22705);
xnor U23375 (N_23375,N_22449,N_22994);
xor U23376 (N_23376,N_22090,N_22977);
and U23377 (N_23377,N_22340,N_22745);
or U23378 (N_23378,N_22612,N_22489);
nand U23379 (N_23379,N_22826,N_22503);
nand U23380 (N_23380,N_22804,N_22266);
xor U23381 (N_23381,N_22204,N_22040);
or U23382 (N_23382,N_22717,N_22531);
or U23383 (N_23383,N_22563,N_22633);
and U23384 (N_23384,N_22022,N_22155);
or U23385 (N_23385,N_22844,N_22059);
nand U23386 (N_23386,N_22847,N_22250);
or U23387 (N_23387,N_22601,N_22624);
and U23388 (N_23388,N_22963,N_22322);
xnor U23389 (N_23389,N_22932,N_22788);
xnor U23390 (N_23390,N_22757,N_22841);
nand U23391 (N_23391,N_22464,N_22479);
nand U23392 (N_23392,N_22024,N_22573);
nor U23393 (N_23393,N_22018,N_22933);
or U23394 (N_23394,N_22604,N_22786);
nand U23395 (N_23395,N_22357,N_22546);
nand U23396 (N_23396,N_22182,N_22066);
nand U23397 (N_23397,N_22588,N_22582);
xnor U23398 (N_23398,N_22809,N_22982);
xnor U23399 (N_23399,N_22481,N_22033);
and U23400 (N_23400,N_22373,N_22986);
or U23401 (N_23401,N_22974,N_22545);
nand U23402 (N_23402,N_22783,N_22348);
or U23403 (N_23403,N_22878,N_22185);
nand U23404 (N_23404,N_22998,N_22792);
nor U23405 (N_23405,N_22850,N_22273);
and U23406 (N_23406,N_22197,N_22474);
or U23407 (N_23407,N_22522,N_22115);
nand U23408 (N_23408,N_22192,N_22153);
and U23409 (N_23409,N_22935,N_22607);
or U23410 (N_23410,N_22768,N_22832);
nor U23411 (N_23411,N_22672,N_22703);
or U23412 (N_23412,N_22315,N_22883);
and U23413 (N_23413,N_22871,N_22198);
or U23414 (N_23414,N_22934,N_22075);
nand U23415 (N_23415,N_22122,N_22045);
or U23416 (N_23416,N_22381,N_22099);
and U23417 (N_23417,N_22830,N_22667);
nor U23418 (N_23418,N_22290,N_22478);
or U23419 (N_23419,N_22791,N_22398);
and U23420 (N_23420,N_22281,N_22181);
nor U23421 (N_23421,N_22391,N_22550);
or U23422 (N_23422,N_22629,N_22781);
nand U23423 (N_23423,N_22782,N_22264);
xor U23424 (N_23424,N_22450,N_22052);
xnor U23425 (N_23425,N_22003,N_22642);
xnor U23426 (N_23426,N_22086,N_22929);
nand U23427 (N_23427,N_22819,N_22882);
xor U23428 (N_23428,N_22923,N_22428);
xnor U23429 (N_23429,N_22605,N_22827);
and U23430 (N_23430,N_22655,N_22486);
xnor U23431 (N_23431,N_22088,N_22070);
xnor U23432 (N_23432,N_22831,N_22227);
xnor U23433 (N_23433,N_22321,N_22219);
xor U23434 (N_23434,N_22263,N_22793);
and U23435 (N_23435,N_22691,N_22623);
or U23436 (N_23436,N_22411,N_22866);
xor U23437 (N_23437,N_22886,N_22983);
nor U23438 (N_23438,N_22356,N_22392);
nor U23439 (N_23439,N_22602,N_22374);
or U23440 (N_23440,N_22371,N_22825);
nor U23441 (N_23441,N_22679,N_22838);
and U23442 (N_23442,N_22444,N_22276);
nor U23443 (N_23443,N_22475,N_22157);
or U23444 (N_23444,N_22936,N_22618);
xnor U23445 (N_23445,N_22802,N_22711);
nand U23446 (N_23446,N_22716,N_22497);
xor U23447 (N_23447,N_22138,N_22188);
nor U23448 (N_23448,N_22393,N_22433);
nor U23449 (N_23449,N_22432,N_22289);
xor U23450 (N_23450,N_22493,N_22993);
or U23451 (N_23451,N_22038,N_22365);
and U23452 (N_23452,N_22278,N_22347);
or U23453 (N_23453,N_22184,N_22989);
nor U23454 (N_23454,N_22093,N_22930);
xnor U23455 (N_23455,N_22412,N_22751);
xnor U23456 (N_23456,N_22282,N_22774);
nand U23457 (N_23457,N_22494,N_22775);
or U23458 (N_23458,N_22482,N_22532);
nand U23459 (N_23459,N_22556,N_22297);
xor U23460 (N_23460,N_22943,N_22962);
xor U23461 (N_23461,N_22701,N_22326);
or U23462 (N_23462,N_22132,N_22715);
and U23463 (N_23463,N_22557,N_22735);
nand U23464 (N_23464,N_22506,N_22721);
or U23465 (N_23465,N_22627,N_22585);
nor U23466 (N_23466,N_22050,N_22614);
nor U23467 (N_23467,N_22719,N_22043);
nor U23468 (N_23468,N_22534,N_22606);
nor U23469 (N_23469,N_22342,N_22732);
xnor U23470 (N_23470,N_22165,N_22436);
and U23471 (N_23471,N_22431,N_22517);
and U23472 (N_23472,N_22430,N_22525);
and U23473 (N_23473,N_22367,N_22308);
and U23474 (N_23474,N_22952,N_22887);
xnor U23475 (N_23475,N_22898,N_22253);
or U23476 (N_23476,N_22168,N_22361);
xor U23477 (N_23477,N_22756,N_22741);
nand U23478 (N_23478,N_22743,N_22159);
and U23479 (N_23479,N_22259,N_22926);
nor U23480 (N_23480,N_22868,N_22231);
and U23481 (N_23481,N_22942,N_22378);
nand U23482 (N_23482,N_22055,N_22798);
nand U23483 (N_23483,N_22584,N_22248);
nand U23484 (N_23484,N_22750,N_22206);
xnor U23485 (N_23485,N_22268,N_22213);
xor U23486 (N_23486,N_22468,N_22677);
or U23487 (N_23487,N_22005,N_22328);
or U23488 (N_23488,N_22762,N_22258);
and U23489 (N_23489,N_22562,N_22693);
or U23490 (N_23490,N_22060,N_22383);
nor U23491 (N_23491,N_22203,N_22950);
xnor U23492 (N_23492,N_22816,N_22136);
nor U23493 (N_23493,N_22789,N_22487);
or U23494 (N_23494,N_22306,N_22492);
nor U23495 (N_23495,N_22890,N_22019);
or U23496 (N_23496,N_22298,N_22661);
xor U23497 (N_23497,N_22764,N_22061);
or U23498 (N_23498,N_22755,N_22353);
xor U23499 (N_23499,N_22553,N_22709);
or U23500 (N_23500,N_22197,N_22397);
nand U23501 (N_23501,N_22842,N_22791);
nand U23502 (N_23502,N_22309,N_22469);
nor U23503 (N_23503,N_22436,N_22212);
and U23504 (N_23504,N_22953,N_22005);
nor U23505 (N_23505,N_22055,N_22268);
nand U23506 (N_23506,N_22692,N_22024);
or U23507 (N_23507,N_22842,N_22637);
nand U23508 (N_23508,N_22082,N_22859);
xnor U23509 (N_23509,N_22554,N_22098);
and U23510 (N_23510,N_22589,N_22354);
xnor U23511 (N_23511,N_22362,N_22861);
and U23512 (N_23512,N_22193,N_22710);
nand U23513 (N_23513,N_22128,N_22962);
nand U23514 (N_23514,N_22371,N_22970);
nor U23515 (N_23515,N_22377,N_22250);
nor U23516 (N_23516,N_22923,N_22468);
and U23517 (N_23517,N_22732,N_22128);
nor U23518 (N_23518,N_22387,N_22316);
xor U23519 (N_23519,N_22158,N_22329);
nand U23520 (N_23520,N_22681,N_22734);
nor U23521 (N_23521,N_22089,N_22914);
nor U23522 (N_23522,N_22079,N_22342);
and U23523 (N_23523,N_22650,N_22654);
xnor U23524 (N_23524,N_22336,N_22490);
nand U23525 (N_23525,N_22496,N_22845);
nor U23526 (N_23526,N_22437,N_22261);
nand U23527 (N_23527,N_22738,N_22375);
and U23528 (N_23528,N_22236,N_22531);
xnor U23529 (N_23529,N_22127,N_22903);
nor U23530 (N_23530,N_22808,N_22519);
and U23531 (N_23531,N_22537,N_22543);
nand U23532 (N_23532,N_22175,N_22674);
and U23533 (N_23533,N_22682,N_22860);
xor U23534 (N_23534,N_22458,N_22523);
nand U23535 (N_23535,N_22115,N_22972);
nand U23536 (N_23536,N_22778,N_22242);
xor U23537 (N_23537,N_22671,N_22116);
or U23538 (N_23538,N_22483,N_22407);
or U23539 (N_23539,N_22659,N_22168);
nor U23540 (N_23540,N_22364,N_22651);
or U23541 (N_23541,N_22776,N_22896);
or U23542 (N_23542,N_22608,N_22264);
nor U23543 (N_23543,N_22295,N_22966);
xor U23544 (N_23544,N_22162,N_22469);
nor U23545 (N_23545,N_22603,N_22416);
xnor U23546 (N_23546,N_22256,N_22080);
nor U23547 (N_23547,N_22751,N_22638);
xor U23548 (N_23548,N_22423,N_22391);
or U23549 (N_23549,N_22282,N_22680);
nand U23550 (N_23550,N_22975,N_22039);
nor U23551 (N_23551,N_22912,N_22955);
or U23552 (N_23552,N_22863,N_22594);
nand U23553 (N_23553,N_22634,N_22742);
xnor U23554 (N_23554,N_22074,N_22550);
and U23555 (N_23555,N_22829,N_22477);
xnor U23556 (N_23556,N_22461,N_22359);
nor U23557 (N_23557,N_22195,N_22811);
nand U23558 (N_23558,N_22178,N_22980);
nand U23559 (N_23559,N_22246,N_22399);
nand U23560 (N_23560,N_22538,N_22986);
and U23561 (N_23561,N_22317,N_22187);
nor U23562 (N_23562,N_22002,N_22879);
or U23563 (N_23563,N_22609,N_22151);
xor U23564 (N_23564,N_22743,N_22427);
and U23565 (N_23565,N_22467,N_22048);
and U23566 (N_23566,N_22744,N_22721);
nor U23567 (N_23567,N_22074,N_22001);
nor U23568 (N_23568,N_22981,N_22228);
nor U23569 (N_23569,N_22864,N_22055);
nor U23570 (N_23570,N_22118,N_22529);
nor U23571 (N_23571,N_22133,N_22838);
or U23572 (N_23572,N_22155,N_22895);
xor U23573 (N_23573,N_22387,N_22207);
or U23574 (N_23574,N_22648,N_22362);
nand U23575 (N_23575,N_22123,N_22711);
nand U23576 (N_23576,N_22194,N_22253);
or U23577 (N_23577,N_22831,N_22644);
and U23578 (N_23578,N_22901,N_22470);
xor U23579 (N_23579,N_22259,N_22474);
and U23580 (N_23580,N_22140,N_22182);
nand U23581 (N_23581,N_22933,N_22207);
nor U23582 (N_23582,N_22927,N_22892);
and U23583 (N_23583,N_22558,N_22210);
xnor U23584 (N_23584,N_22342,N_22555);
and U23585 (N_23585,N_22873,N_22429);
nand U23586 (N_23586,N_22488,N_22453);
nor U23587 (N_23587,N_22719,N_22545);
nor U23588 (N_23588,N_22902,N_22919);
nand U23589 (N_23589,N_22455,N_22589);
nor U23590 (N_23590,N_22585,N_22210);
and U23591 (N_23591,N_22162,N_22700);
and U23592 (N_23592,N_22689,N_22951);
nor U23593 (N_23593,N_22615,N_22519);
nand U23594 (N_23594,N_22218,N_22846);
nor U23595 (N_23595,N_22449,N_22372);
xor U23596 (N_23596,N_22147,N_22167);
nand U23597 (N_23597,N_22036,N_22225);
xnor U23598 (N_23598,N_22834,N_22835);
nor U23599 (N_23599,N_22001,N_22680);
nor U23600 (N_23600,N_22936,N_22343);
nand U23601 (N_23601,N_22891,N_22832);
and U23602 (N_23602,N_22893,N_22788);
nand U23603 (N_23603,N_22828,N_22361);
nor U23604 (N_23604,N_22270,N_22335);
xnor U23605 (N_23605,N_22891,N_22424);
nor U23606 (N_23606,N_22498,N_22474);
and U23607 (N_23607,N_22851,N_22089);
and U23608 (N_23608,N_22451,N_22988);
nand U23609 (N_23609,N_22164,N_22767);
or U23610 (N_23610,N_22811,N_22223);
nand U23611 (N_23611,N_22390,N_22790);
nor U23612 (N_23612,N_22277,N_22919);
and U23613 (N_23613,N_22291,N_22799);
nor U23614 (N_23614,N_22346,N_22964);
or U23615 (N_23615,N_22415,N_22456);
and U23616 (N_23616,N_22142,N_22246);
or U23617 (N_23617,N_22005,N_22861);
and U23618 (N_23618,N_22136,N_22373);
nand U23619 (N_23619,N_22090,N_22614);
nand U23620 (N_23620,N_22740,N_22542);
and U23621 (N_23621,N_22115,N_22156);
nor U23622 (N_23622,N_22132,N_22946);
and U23623 (N_23623,N_22180,N_22022);
or U23624 (N_23624,N_22559,N_22542);
and U23625 (N_23625,N_22945,N_22616);
or U23626 (N_23626,N_22202,N_22304);
nor U23627 (N_23627,N_22910,N_22347);
nand U23628 (N_23628,N_22246,N_22494);
or U23629 (N_23629,N_22549,N_22699);
and U23630 (N_23630,N_22656,N_22605);
and U23631 (N_23631,N_22953,N_22382);
nand U23632 (N_23632,N_22985,N_22019);
nor U23633 (N_23633,N_22896,N_22228);
or U23634 (N_23634,N_22427,N_22900);
xor U23635 (N_23635,N_22045,N_22136);
nand U23636 (N_23636,N_22554,N_22726);
nor U23637 (N_23637,N_22111,N_22964);
xor U23638 (N_23638,N_22876,N_22304);
or U23639 (N_23639,N_22322,N_22172);
and U23640 (N_23640,N_22647,N_22195);
nand U23641 (N_23641,N_22229,N_22051);
or U23642 (N_23642,N_22415,N_22856);
xor U23643 (N_23643,N_22895,N_22172);
nor U23644 (N_23644,N_22492,N_22915);
and U23645 (N_23645,N_22590,N_22253);
xor U23646 (N_23646,N_22017,N_22590);
nand U23647 (N_23647,N_22359,N_22115);
nand U23648 (N_23648,N_22142,N_22810);
and U23649 (N_23649,N_22502,N_22996);
nand U23650 (N_23650,N_22182,N_22071);
or U23651 (N_23651,N_22816,N_22571);
or U23652 (N_23652,N_22980,N_22745);
nor U23653 (N_23653,N_22007,N_22458);
nand U23654 (N_23654,N_22146,N_22245);
or U23655 (N_23655,N_22415,N_22300);
nor U23656 (N_23656,N_22650,N_22258);
xor U23657 (N_23657,N_22615,N_22541);
or U23658 (N_23658,N_22468,N_22154);
nor U23659 (N_23659,N_22186,N_22872);
or U23660 (N_23660,N_22059,N_22175);
and U23661 (N_23661,N_22035,N_22619);
nor U23662 (N_23662,N_22293,N_22006);
xor U23663 (N_23663,N_22396,N_22650);
and U23664 (N_23664,N_22666,N_22454);
xor U23665 (N_23665,N_22933,N_22298);
nand U23666 (N_23666,N_22957,N_22749);
or U23667 (N_23667,N_22715,N_22439);
xnor U23668 (N_23668,N_22306,N_22456);
nor U23669 (N_23669,N_22254,N_22323);
xnor U23670 (N_23670,N_22277,N_22095);
and U23671 (N_23671,N_22302,N_22308);
and U23672 (N_23672,N_22298,N_22084);
or U23673 (N_23673,N_22447,N_22841);
nor U23674 (N_23674,N_22879,N_22711);
nor U23675 (N_23675,N_22552,N_22798);
and U23676 (N_23676,N_22708,N_22829);
xor U23677 (N_23677,N_22835,N_22434);
xor U23678 (N_23678,N_22026,N_22096);
and U23679 (N_23679,N_22816,N_22198);
and U23680 (N_23680,N_22228,N_22937);
or U23681 (N_23681,N_22949,N_22491);
nor U23682 (N_23682,N_22074,N_22227);
or U23683 (N_23683,N_22079,N_22351);
xor U23684 (N_23684,N_22438,N_22414);
or U23685 (N_23685,N_22593,N_22215);
nor U23686 (N_23686,N_22432,N_22575);
and U23687 (N_23687,N_22503,N_22014);
or U23688 (N_23688,N_22980,N_22827);
and U23689 (N_23689,N_22872,N_22107);
and U23690 (N_23690,N_22625,N_22732);
nor U23691 (N_23691,N_22043,N_22213);
or U23692 (N_23692,N_22358,N_22024);
and U23693 (N_23693,N_22495,N_22635);
nor U23694 (N_23694,N_22196,N_22749);
xor U23695 (N_23695,N_22559,N_22180);
and U23696 (N_23696,N_22584,N_22321);
xnor U23697 (N_23697,N_22462,N_22471);
or U23698 (N_23698,N_22908,N_22957);
nor U23699 (N_23699,N_22284,N_22744);
nand U23700 (N_23700,N_22207,N_22607);
and U23701 (N_23701,N_22197,N_22700);
and U23702 (N_23702,N_22730,N_22558);
nand U23703 (N_23703,N_22788,N_22435);
and U23704 (N_23704,N_22420,N_22363);
nor U23705 (N_23705,N_22973,N_22712);
and U23706 (N_23706,N_22913,N_22010);
or U23707 (N_23707,N_22936,N_22339);
nor U23708 (N_23708,N_22230,N_22739);
and U23709 (N_23709,N_22592,N_22146);
and U23710 (N_23710,N_22510,N_22295);
and U23711 (N_23711,N_22637,N_22874);
and U23712 (N_23712,N_22694,N_22417);
nor U23713 (N_23713,N_22657,N_22702);
and U23714 (N_23714,N_22100,N_22818);
and U23715 (N_23715,N_22324,N_22986);
nand U23716 (N_23716,N_22927,N_22443);
nand U23717 (N_23717,N_22611,N_22159);
nand U23718 (N_23718,N_22350,N_22495);
or U23719 (N_23719,N_22899,N_22332);
nand U23720 (N_23720,N_22773,N_22226);
nand U23721 (N_23721,N_22737,N_22217);
nand U23722 (N_23722,N_22698,N_22306);
xor U23723 (N_23723,N_22606,N_22365);
nor U23724 (N_23724,N_22637,N_22495);
and U23725 (N_23725,N_22805,N_22998);
and U23726 (N_23726,N_22599,N_22792);
xnor U23727 (N_23727,N_22247,N_22028);
nor U23728 (N_23728,N_22987,N_22080);
and U23729 (N_23729,N_22740,N_22061);
nor U23730 (N_23730,N_22485,N_22314);
xnor U23731 (N_23731,N_22297,N_22685);
xnor U23732 (N_23732,N_22745,N_22683);
nor U23733 (N_23733,N_22993,N_22793);
nor U23734 (N_23734,N_22219,N_22980);
nand U23735 (N_23735,N_22513,N_22417);
or U23736 (N_23736,N_22652,N_22226);
nand U23737 (N_23737,N_22508,N_22563);
nand U23738 (N_23738,N_22171,N_22642);
nor U23739 (N_23739,N_22972,N_22559);
nor U23740 (N_23740,N_22805,N_22654);
nor U23741 (N_23741,N_22574,N_22484);
xnor U23742 (N_23742,N_22653,N_22307);
xor U23743 (N_23743,N_22839,N_22079);
xor U23744 (N_23744,N_22612,N_22264);
and U23745 (N_23745,N_22123,N_22541);
nor U23746 (N_23746,N_22448,N_22980);
nand U23747 (N_23747,N_22318,N_22013);
or U23748 (N_23748,N_22595,N_22490);
nor U23749 (N_23749,N_22644,N_22270);
and U23750 (N_23750,N_22311,N_22554);
xnor U23751 (N_23751,N_22189,N_22045);
nor U23752 (N_23752,N_22239,N_22898);
nor U23753 (N_23753,N_22730,N_22100);
nand U23754 (N_23754,N_22566,N_22771);
and U23755 (N_23755,N_22504,N_22501);
nor U23756 (N_23756,N_22364,N_22376);
xnor U23757 (N_23757,N_22913,N_22997);
and U23758 (N_23758,N_22116,N_22692);
nand U23759 (N_23759,N_22566,N_22322);
nand U23760 (N_23760,N_22135,N_22837);
nor U23761 (N_23761,N_22564,N_22964);
nor U23762 (N_23762,N_22706,N_22786);
or U23763 (N_23763,N_22182,N_22209);
and U23764 (N_23764,N_22917,N_22860);
nand U23765 (N_23765,N_22328,N_22413);
xnor U23766 (N_23766,N_22113,N_22425);
nor U23767 (N_23767,N_22761,N_22679);
nor U23768 (N_23768,N_22180,N_22595);
or U23769 (N_23769,N_22696,N_22599);
or U23770 (N_23770,N_22527,N_22230);
nand U23771 (N_23771,N_22355,N_22935);
nand U23772 (N_23772,N_22360,N_22730);
and U23773 (N_23773,N_22603,N_22780);
xor U23774 (N_23774,N_22697,N_22593);
or U23775 (N_23775,N_22571,N_22329);
and U23776 (N_23776,N_22734,N_22313);
xnor U23777 (N_23777,N_22845,N_22156);
and U23778 (N_23778,N_22942,N_22112);
nor U23779 (N_23779,N_22506,N_22557);
and U23780 (N_23780,N_22048,N_22094);
and U23781 (N_23781,N_22651,N_22016);
or U23782 (N_23782,N_22017,N_22007);
xnor U23783 (N_23783,N_22888,N_22004);
nand U23784 (N_23784,N_22333,N_22081);
or U23785 (N_23785,N_22118,N_22932);
nand U23786 (N_23786,N_22984,N_22150);
xnor U23787 (N_23787,N_22027,N_22960);
or U23788 (N_23788,N_22319,N_22033);
nand U23789 (N_23789,N_22241,N_22139);
nand U23790 (N_23790,N_22108,N_22207);
xor U23791 (N_23791,N_22916,N_22608);
nand U23792 (N_23792,N_22326,N_22599);
nor U23793 (N_23793,N_22368,N_22300);
nand U23794 (N_23794,N_22625,N_22290);
or U23795 (N_23795,N_22243,N_22386);
and U23796 (N_23796,N_22761,N_22866);
xor U23797 (N_23797,N_22570,N_22997);
or U23798 (N_23798,N_22020,N_22700);
nor U23799 (N_23799,N_22540,N_22526);
xor U23800 (N_23800,N_22192,N_22032);
nand U23801 (N_23801,N_22943,N_22458);
nand U23802 (N_23802,N_22402,N_22773);
nand U23803 (N_23803,N_22007,N_22609);
xor U23804 (N_23804,N_22384,N_22635);
and U23805 (N_23805,N_22495,N_22988);
nand U23806 (N_23806,N_22950,N_22890);
nor U23807 (N_23807,N_22810,N_22261);
and U23808 (N_23808,N_22869,N_22453);
xnor U23809 (N_23809,N_22028,N_22231);
and U23810 (N_23810,N_22035,N_22480);
nand U23811 (N_23811,N_22891,N_22672);
nor U23812 (N_23812,N_22885,N_22597);
xnor U23813 (N_23813,N_22169,N_22346);
or U23814 (N_23814,N_22028,N_22380);
nand U23815 (N_23815,N_22396,N_22001);
and U23816 (N_23816,N_22960,N_22124);
and U23817 (N_23817,N_22350,N_22459);
xor U23818 (N_23818,N_22860,N_22164);
or U23819 (N_23819,N_22203,N_22434);
nor U23820 (N_23820,N_22129,N_22256);
nand U23821 (N_23821,N_22961,N_22195);
and U23822 (N_23822,N_22874,N_22033);
or U23823 (N_23823,N_22238,N_22993);
or U23824 (N_23824,N_22994,N_22025);
or U23825 (N_23825,N_22694,N_22875);
nor U23826 (N_23826,N_22203,N_22944);
xor U23827 (N_23827,N_22224,N_22392);
and U23828 (N_23828,N_22897,N_22761);
xnor U23829 (N_23829,N_22620,N_22894);
nand U23830 (N_23830,N_22625,N_22192);
nor U23831 (N_23831,N_22467,N_22495);
nand U23832 (N_23832,N_22502,N_22772);
nor U23833 (N_23833,N_22031,N_22198);
nor U23834 (N_23834,N_22820,N_22608);
xor U23835 (N_23835,N_22681,N_22411);
or U23836 (N_23836,N_22410,N_22871);
nor U23837 (N_23837,N_22425,N_22795);
xor U23838 (N_23838,N_22907,N_22418);
and U23839 (N_23839,N_22645,N_22799);
nor U23840 (N_23840,N_22392,N_22418);
nor U23841 (N_23841,N_22226,N_22116);
nor U23842 (N_23842,N_22054,N_22214);
xor U23843 (N_23843,N_22002,N_22369);
nand U23844 (N_23844,N_22891,N_22843);
xnor U23845 (N_23845,N_22721,N_22155);
and U23846 (N_23846,N_22812,N_22210);
nor U23847 (N_23847,N_22884,N_22471);
nand U23848 (N_23848,N_22498,N_22356);
nor U23849 (N_23849,N_22278,N_22981);
or U23850 (N_23850,N_22078,N_22139);
or U23851 (N_23851,N_22269,N_22072);
and U23852 (N_23852,N_22576,N_22082);
xor U23853 (N_23853,N_22148,N_22182);
nand U23854 (N_23854,N_22712,N_22093);
nand U23855 (N_23855,N_22798,N_22556);
xnor U23856 (N_23856,N_22053,N_22897);
xor U23857 (N_23857,N_22355,N_22038);
or U23858 (N_23858,N_22944,N_22708);
nand U23859 (N_23859,N_22957,N_22149);
nor U23860 (N_23860,N_22392,N_22471);
or U23861 (N_23861,N_22056,N_22359);
or U23862 (N_23862,N_22259,N_22191);
or U23863 (N_23863,N_22230,N_22426);
and U23864 (N_23864,N_22561,N_22434);
nor U23865 (N_23865,N_22889,N_22306);
and U23866 (N_23866,N_22190,N_22549);
xor U23867 (N_23867,N_22666,N_22635);
nor U23868 (N_23868,N_22021,N_22127);
nor U23869 (N_23869,N_22365,N_22757);
nand U23870 (N_23870,N_22098,N_22942);
nor U23871 (N_23871,N_22801,N_22724);
xnor U23872 (N_23872,N_22736,N_22182);
or U23873 (N_23873,N_22286,N_22676);
or U23874 (N_23874,N_22378,N_22625);
nand U23875 (N_23875,N_22595,N_22807);
nand U23876 (N_23876,N_22455,N_22280);
nand U23877 (N_23877,N_22864,N_22136);
nor U23878 (N_23878,N_22068,N_22872);
nand U23879 (N_23879,N_22427,N_22200);
nand U23880 (N_23880,N_22089,N_22394);
nor U23881 (N_23881,N_22517,N_22421);
nand U23882 (N_23882,N_22955,N_22596);
xor U23883 (N_23883,N_22208,N_22498);
xor U23884 (N_23884,N_22919,N_22759);
or U23885 (N_23885,N_22532,N_22896);
or U23886 (N_23886,N_22141,N_22016);
nand U23887 (N_23887,N_22243,N_22607);
and U23888 (N_23888,N_22094,N_22658);
nor U23889 (N_23889,N_22979,N_22389);
xnor U23890 (N_23890,N_22317,N_22190);
and U23891 (N_23891,N_22043,N_22839);
or U23892 (N_23892,N_22497,N_22112);
nor U23893 (N_23893,N_22256,N_22663);
nand U23894 (N_23894,N_22258,N_22130);
nor U23895 (N_23895,N_22335,N_22733);
or U23896 (N_23896,N_22559,N_22421);
or U23897 (N_23897,N_22177,N_22799);
nor U23898 (N_23898,N_22828,N_22398);
nor U23899 (N_23899,N_22587,N_22693);
nand U23900 (N_23900,N_22301,N_22314);
nor U23901 (N_23901,N_22567,N_22692);
xnor U23902 (N_23902,N_22186,N_22504);
and U23903 (N_23903,N_22364,N_22851);
nand U23904 (N_23904,N_22755,N_22539);
nand U23905 (N_23905,N_22643,N_22894);
and U23906 (N_23906,N_22276,N_22759);
and U23907 (N_23907,N_22674,N_22887);
nand U23908 (N_23908,N_22984,N_22200);
xor U23909 (N_23909,N_22483,N_22968);
or U23910 (N_23910,N_22044,N_22488);
nor U23911 (N_23911,N_22677,N_22275);
xnor U23912 (N_23912,N_22198,N_22885);
nor U23913 (N_23913,N_22268,N_22859);
and U23914 (N_23914,N_22382,N_22579);
and U23915 (N_23915,N_22529,N_22652);
xor U23916 (N_23916,N_22027,N_22160);
and U23917 (N_23917,N_22594,N_22872);
nand U23918 (N_23918,N_22090,N_22237);
nor U23919 (N_23919,N_22634,N_22447);
nor U23920 (N_23920,N_22867,N_22585);
and U23921 (N_23921,N_22621,N_22048);
xor U23922 (N_23922,N_22090,N_22375);
xor U23923 (N_23923,N_22508,N_22530);
or U23924 (N_23924,N_22190,N_22082);
and U23925 (N_23925,N_22971,N_22474);
xnor U23926 (N_23926,N_22102,N_22912);
and U23927 (N_23927,N_22682,N_22670);
nand U23928 (N_23928,N_22169,N_22711);
nor U23929 (N_23929,N_22422,N_22723);
and U23930 (N_23930,N_22780,N_22170);
xnor U23931 (N_23931,N_22771,N_22248);
nor U23932 (N_23932,N_22289,N_22259);
and U23933 (N_23933,N_22662,N_22758);
or U23934 (N_23934,N_22203,N_22931);
nand U23935 (N_23935,N_22755,N_22375);
nand U23936 (N_23936,N_22055,N_22793);
or U23937 (N_23937,N_22156,N_22299);
or U23938 (N_23938,N_22282,N_22301);
nor U23939 (N_23939,N_22339,N_22562);
xnor U23940 (N_23940,N_22837,N_22288);
xor U23941 (N_23941,N_22834,N_22866);
nand U23942 (N_23942,N_22994,N_22690);
xor U23943 (N_23943,N_22866,N_22414);
or U23944 (N_23944,N_22388,N_22157);
and U23945 (N_23945,N_22156,N_22001);
and U23946 (N_23946,N_22116,N_22002);
or U23947 (N_23947,N_22710,N_22325);
and U23948 (N_23948,N_22536,N_22749);
nand U23949 (N_23949,N_22004,N_22702);
or U23950 (N_23950,N_22029,N_22811);
and U23951 (N_23951,N_22077,N_22989);
nor U23952 (N_23952,N_22225,N_22158);
nand U23953 (N_23953,N_22453,N_22720);
nand U23954 (N_23954,N_22056,N_22211);
and U23955 (N_23955,N_22595,N_22368);
nand U23956 (N_23956,N_22110,N_22810);
and U23957 (N_23957,N_22329,N_22033);
nand U23958 (N_23958,N_22258,N_22973);
and U23959 (N_23959,N_22099,N_22979);
xnor U23960 (N_23960,N_22701,N_22638);
and U23961 (N_23961,N_22505,N_22859);
or U23962 (N_23962,N_22696,N_22408);
xnor U23963 (N_23963,N_22175,N_22082);
or U23964 (N_23964,N_22681,N_22613);
xor U23965 (N_23965,N_22357,N_22733);
nand U23966 (N_23966,N_22319,N_22886);
xnor U23967 (N_23967,N_22137,N_22706);
xor U23968 (N_23968,N_22315,N_22776);
xnor U23969 (N_23969,N_22611,N_22017);
or U23970 (N_23970,N_22857,N_22251);
nand U23971 (N_23971,N_22248,N_22034);
nand U23972 (N_23972,N_22148,N_22507);
or U23973 (N_23973,N_22637,N_22947);
and U23974 (N_23974,N_22584,N_22571);
xor U23975 (N_23975,N_22443,N_22412);
and U23976 (N_23976,N_22407,N_22587);
or U23977 (N_23977,N_22677,N_22953);
nand U23978 (N_23978,N_22179,N_22286);
nand U23979 (N_23979,N_22565,N_22870);
nor U23980 (N_23980,N_22499,N_22640);
and U23981 (N_23981,N_22987,N_22561);
xnor U23982 (N_23982,N_22223,N_22095);
nor U23983 (N_23983,N_22894,N_22360);
nor U23984 (N_23984,N_22321,N_22139);
nor U23985 (N_23985,N_22204,N_22368);
and U23986 (N_23986,N_22713,N_22283);
or U23987 (N_23987,N_22215,N_22456);
or U23988 (N_23988,N_22378,N_22801);
nor U23989 (N_23989,N_22680,N_22258);
and U23990 (N_23990,N_22371,N_22129);
xor U23991 (N_23991,N_22423,N_22143);
nor U23992 (N_23992,N_22112,N_22848);
xor U23993 (N_23993,N_22592,N_22113);
or U23994 (N_23994,N_22534,N_22883);
and U23995 (N_23995,N_22076,N_22730);
nand U23996 (N_23996,N_22171,N_22021);
nor U23997 (N_23997,N_22979,N_22741);
nor U23998 (N_23998,N_22816,N_22623);
nand U23999 (N_23999,N_22224,N_22935);
nor U24000 (N_24000,N_23114,N_23306);
nor U24001 (N_24001,N_23368,N_23847);
nand U24002 (N_24002,N_23593,N_23345);
or U24003 (N_24003,N_23464,N_23727);
nor U24004 (N_24004,N_23956,N_23842);
xnor U24005 (N_24005,N_23200,N_23288);
and U24006 (N_24006,N_23825,N_23874);
nor U24007 (N_24007,N_23041,N_23846);
xnor U24008 (N_24008,N_23508,N_23377);
xor U24009 (N_24009,N_23666,N_23946);
and U24010 (N_24010,N_23292,N_23927);
and U24011 (N_24011,N_23777,N_23212);
or U24012 (N_24012,N_23894,N_23559);
xor U24013 (N_24013,N_23684,N_23366);
nand U24014 (N_24014,N_23256,N_23421);
nor U24015 (N_24015,N_23098,N_23580);
or U24016 (N_24016,N_23264,N_23837);
nor U24017 (N_24017,N_23068,N_23836);
nor U24018 (N_24018,N_23605,N_23764);
nor U24019 (N_24019,N_23109,N_23036);
xnor U24020 (N_24020,N_23227,N_23574);
and U24021 (N_24021,N_23974,N_23702);
or U24022 (N_24022,N_23102,N_23970);
xnor U24023 (N_24023,N_23929,N_23881);
nor U24024 (N_24024,N_23071,N_23797);
xor U24025 (N_24025,N_23685,N_23154);
and U24026 (N_24026,N_23561,N_23058);
and U24027 (N_24027,N_23455,N_23545);
or U24028 (N_24028,N_23614,N_23745);
or U24029 (N_24029,N_23230,N_23885);
or U24030 (N_24030,N_23121,N_23748);
or U24031 (N_24031,N_23273,N_23641);
xor U24032 (N_24032,N_23689,N_23238);
nand U24033 (N_24033,N_23481,N_23059);
xnor U24034 (N_24034,N_23719,N_23184);
and U24035 (N_24035,N_23995,N_23953);
nand U24036 (N_24036,N_23002,N_23656);
nand U24037 (N_24037,N_23812,N_23699);
xor U24038 (N_24038,N_23514,N_23105);
xnor U24039 (N_24039,N_23131,N_23143);
nand U24040 (N_24040,N_23643,N_23280);
or U24041 (N_24041,N_23770,N_23549);
or U24042 (N_24042,N_23696,N_23371);
or U24043 (N_24043,N_23810,N_23274);
xor U24044 (N_24044,N_23445,N_23494);
nand U24045 (N_24045,N_23213,N_23153);
or U24046 (N_24046,N_23207,N_23983);
xnor U24047 (N_24047,N_23231,N_23729);
xor U24048 (N_24048,N_23715,N_23343);
nand U24049 (N_24049,N_23808,N_23319);
nor U24050 (N_24050,N_23909,N_23570);
nor U24051 (N_24051,N_23320,N_23356);
or U24052 (N_24052,N_23890,N_23814);
and U24053 (N_24053,N_23788,N_23316);
nand U24054 (N_24054,N_23707,N_23007);
nor U24055 (N_24055,N_23826,N_23216);
nor U24056 (N_24056,N_23205,N_23204);
nor U24057 (N_24057,N_23783,N_23222);
and U24058 (N_24058,N_23300,N_23711);
nand U24059 (N_24059,N_23916,N_23015);
nor U24060 (N_24060,N_23444,N_23518);
xor U24061 (N_24061,N_23203,N_23112);
nor U24062 (N_24062,N_23000,N_23501);
and U24063 (N_24063,N_23585,N_23528);
xor U24064 (N_24064,N_23789,N_23655);
and U24065 (N_24065,N_23296,N_23022);
nand U24066 (N_24066,N_23311,N_23811);
nor U24067 (N_24067,N_23394,N_23660);
xnor U24068 (N_24068,N_23506,N_23717);
nor U24069 (N_24069,N_23461,N_23252);
xnor U24070 (N_24070,N_23698,N_23803);
and U24071 (N_24071,N_23199,N_23893);
and U24072 (N_24072,N_23452,N_23673);
or U24073 (N_24073,N_23784,N_23647);
or U24074 (N_24074,N_23841,N_23567);
nor U24075 (N_24075,N_23492,N_23785);
xor U24076 (N_24076,N_23510,N_23820);
xnor U24077 (N_24077,N_23863,N_23755);
nor U24078 (N_24078,N_23101,N_23531);
nand U24079 (N_24079,N_23287,N_23989);
nand U24080 (N_24080,N_23569,N_23333);
nand U24081 (N_24081,N_23761,N_23185);
or U24082 (N_24082,N_23291,N_23592);
xor U24083 (N_24083,N_23683,N_23977);
nor U24084 (N_24084,N_23511,N_23395);
nand U24085 (N_24085,N_23026,N_23357);
or U24086 (N_24086,N_23600,N_23879);
nand U24087 (N_24087,N_23873,N_23503);
xor U24088 (N_24088,N_23535,N_23253);
and U24089 (N_24089,N_23383,N_23906);
and U24090 (N_24090,N_23613,N_23201);
and U24091 (N_24091,N_23821,N_23375);
nor U24092 (N_24092,N_23959,N_23313);
nand U24093 (N_24093,N_23171,N_23017);
xnor U24094 (N_24094,N_23370,N_23267);
nand U24095 (N_24095,N_23229,N_23297);
or U24096 (N_24096,N_23969,N_23393);
nor U24097 (N_24097,N_23801,N_23431);
nor U24098 (N_24098,N_23575,N_23878);
nand U24099 (N_24099,N_23215,N_23723);
nor U24100 (N_24100,N_23427,N_23588);
nand U24101 (N_24101,N_23374,N_23720);
nor U24102 (N_24102,N_23122,N_23219);
nand U24103 (N_24103,N_23178,N_23888);
or U24104 (N_24104,N_23485,N_23335);
nand U24105 (N_24105,N_23621,N_23456);
xor U24106 (N_24106,N_23539,N_23057);
nor U24107 (N_24107,N_23167,N_23609);
xnor U24108 (N_24108,N_23532,N_23314);
and U24109 (N_24109,N_23794,N_23930);
nand U24110 (N_24110,N_23671,N_23399);
xor U24111 (N_24111,N_23019,N_23623);
nor U24112 (N_24112,N_23591,N_23055);
and U24113 (N_24113,N_23355,N_23759);
nor U24114 (N_24114,N_23649,N_23008);
nor U24115 (N_24115,N_23822,N_23134);
nor U24116 (N_24116,N_23586,N_23447);
xor U24117 (N_24117,N_23118,N_23018);
nor U24118 (N_24118,N_23945,N_23413);
or U24119 (N_24119,N_23576,N_23804);
nand U24120 (N_24120,N_23617,N_23080);
nand U24121 (N_24121,N_23465,N_23910);
or U24122 (N_24122,N_23188,N_23750);
nor U24123 (N_24123,N_23376,N_23857);
nand U24124 (N_24124,N_23951,N_23861);
nor U24125 (N_24125,N_23138,N_23289);
nor U24126 (N_24126,N_23406,N_23913);
and U24127 (N_24127,N_23347,N_23218);
nand U24128 (N_24128,N_23831,N_23976);
or U24129 (N_24129,N_23217,N_23500);
nor U24130 (N_24130,N_23752,N_23560);
or U24131 (N_24131,N_23799,N_23620);
or U24132 (N_24132,N_23520,N_23780);
nand U24133 (N_24133,N_23350,N_23975);
xnor U24134 (N_24134,N_23544,N_23747);
nor U24135 (N_24135,N_23434,N_23441);
or U24136 (N_24136,N_23996,N_23607);
and U24137 (N_24137,N_23793,N_23858);
or U24138 (N_24138,N_23426,N_23984);
nand U24139 (N_24139,N_23891,N_23454);
or U24140 (N_24140,N_23190,N_23577);
xor U24141 (N_24141,N_23308,N_23092);
or U24142 (N_24142,N_23957,N_23078);
nand U24143 (N_24143,N_23373,N_23769);
and U24144 (N_24144,N_23579,N_23224);
xor U24145 (N_24145,N_23411,N_23818);
xnor U24146 (N_24146,N_23497,N_23923);
nand U24147 (N_24147,N_23733,N_23266);
or U24148 (N_24148,N_23063,N_23283);
or U24149 (N_24149,N_23795,N_23499);
xor U24150 (N_24150,N_23072,N_23304);
xor U24151 (N_24151,N_23408,N_23541);
nand U24152 (N_24152,N_23372,N_23381);
nand U24153 (N_24153,N_23833,N_23488);
and U24154 (N_24154,N_23303,N_23947);
and U24155 (N_24155,N_23941,N_23312);
or U24156 (N_24156,N_23645,N_23410);
nand U24157 (N_24157,N_23527,N_23123);
nand U24158 (N_24158,N_23270,N_23116);
xnor U24159 (N_24159,N_23151,N_23133);
nand U24160 (N_24160,N_23602,N_23104);
nand U24161 (N_24161,N_23147,N_23048);
xnor U24162 (N_24162,N_23140,N_23403);
nand U24163 (N_24163,N_23901,N_23392);
nand U24164 (N_24164,N_23150,N_23236);
and U24165 (N_24165,N_23859,N_23704);
nand U24166 (N_24166,N_23449,N_23997);
nand U24167 (N_24167,N_23220,N_23737);
or U24168 (N_24168,N_23364,N_23603);
or U24169 (N_24169,N_23043,N_23652);
or U24170 (N_24170,N_23502,N_23191);
and U24171 (N_24171,N_23039,N_23095);
xor U24172 (N_24172,N_23778,N_23630);
or U24173 (N_24173,N_23176,N_23054);
nand U24174 (N_24174,N_23337,N_23701);
or U24175 (N_24175,N_23965,N_23892);
nor U24176 (N_24176,N_23931,N_23084);
nor U24177 (N_24177,N_23644,N_23871);
and U24178 (N_24178,N_23174,N_23182);
or U24179 (N_24179,N_23265,N_23548);
and U24180 (N_24180,N_23438,N_23993);
nor U24181 (N_24181,N_23553,N_23004);
nand U24182 (N_24182,N_23523,N_23736);
or U24183 (N_24183,N_23616,N_23515);
and U24184 (N_24184,N_23936,N_23159);
nand U24185 (N_24185,N_23064,N_23360);
or U24186 (N_24186,N_23546,N_23386);
xor U24187 (N_24187,N_23233,N_23897);
nor U24188 (N_24188,N_23670,N_23418);
xnor U24189 (N_24189,N_23021,N_23954);
nor U24190 (N_24190,N_23606,N_23971);
or U24191 (N_24191,N_23024,N_23525);
xnor U24192 (N_24192,N_23415,N_23391);
or U24193 (N_24193,N_23155,N_23905);
nor U24194 (N_24194,N_23106,N_23932);
or U24195 (N_24195,N_23677,N_23866);
xor U24196 (N_24196,N_23158,N_23145);
nand U24197 (N_24197,N_23676,N_23478);
xor U24198 (N_24198,N_23091,N_23639);
xor U24199 (N_24199,N_23248,N_23246);
nor U24200 (N_24200,N_23211,N_23658);
and U24201 (N_24201,N_23542,N_23556);
nor U24202 (N_24202,N_23128,N_23470);
xor U24203 (N_24203,N_23537,N_23486);
xor U24204 (N_24204,N_23838,N_23680);
nand U24205 (N_24205,N_23782,N_23775);
nor U24206 (N_24206,N_23958,N_23848);
xnor U24207 (N_24207,N_23322,N_23615);
nor U24208 (N_24208,N_23005,N_23705);
nand U24209 (N_24209,N_23686,N_23419);
nor U24210 (N_24210,N_23436,N_23533);
xnor U24211 (N_24211,N_23309,N_23596);
xor U24212 (N_24212,N_23405,N_23519);
xor U24213 (N_24213,N_23202,N_23587);
and U24214 (N_24214,N_23193,N_23524);
nor U24215 (N_24215,N_23629,N_23754);
xnor U24216 (N_24216,N_23013,N_23214);
and U24217 (N_24217,N_23388,N_23088);
nand U24218 (N_24218,N_23380,N_23990);
nand U24219 (N_24219,N_23779,N_23853);
nand U24220 (N_24220,N_23489,N_23934);
and U24221 (N_24221,N_23498,N_23079);
or U24222 (N_24222,N_23898,N_23743);
or U24223 (N_24223,N_23664,N_23849);
xnor U24224 (N_24224,N_23166,N_23554);
nor U24225 (N_24225,N_23513,N_23295);
xnor U24226 (N_24226,N_23618,N_23242);
or U24227 (N_24227,N_23301,N_23318);
or U24228 (N_24228,N_23067,N_23282);
nand U24229 (N_24229,N_23479,N_23796);
and U24230 (N_24230,N_23966,N_23132);
and U24231 (N_24231,N_23762,N_23772);
xnor U24232 (N_24232,N_23854,N_23096);
nand U24233 (N_24233,N_23558,N_23581);
xor U24234 (N_24234,N_23305,N_23389);
nor U24235 (N_24235,N_23285,N_23526);
and U24236 (N_24236,N_23061,N_23551);
nand U24237 (N_24237,N_23344,N_23573);
nor U24238 (N_24238,N_23177,N_23255);
nand U24239 (N_24239,N_23249,N_23186);
xnor U24240 (N_24240,N_23693,N_23361);
xor U24241 (N_24241,N_23900,N_23756);
and U24242 (N_24242,N_23338,N_23033);
xor U24243 (N_24243,N_23850,N_23608);
and U24244 (N_24244,N_23964,N_23981);
nor U24245 (N_24245,N_23340,N_23099);
and U24246 (N_24246,N_23198,N_23046);
xor U24247 (N_24247,N_23272,N_23100);
nor U24248 (N_24248,N_23776,N_23991);
nand U24249 (N_24249,N_23688,N_23578);
and U24250 (N_24250,N_23823,N_23237);
and U24251 (N_24251,N_23844,N_23724);
or U24252 (N_24252,N_23787,N_23011);
or U24253 (N_24253,N_23758,N_23612);
or U24254 (N_24254,N_23922,N_23865);
or U24255 (N_24255,N_23495,N_23156);
nand U24256 (N_24256,N_23387,N_23160);
nor U24257 (N_24257,N_23307,N_23604);
or U24258 (N_24258,N_23757,N_23734);
nand U24259 (N_24259,N_23139,N_23697);
or U24260 (N_24260,N_23839,N_23740);
nor U24261 (N_24261,N_23960,N_23250);
nand U24262 (N_24262,N_23358,N_23732);
and U24263 (N_24263,N_23710,N_23721);
or U24264 (N_24264,N_23115,N_23584);
and U24265 (N_24265,N_23884,N_23328);
nor U24266 (N_24266,N_23610,N_23994);
xor U24267 (N_24267,N_23774,N_23800);
xnor U24268 (N_24268,N_23493,N_23299);
and U24269 (N_24269,N_23552,N_23654);
and U24270 (N_24270,N_23446,N_23060);
xnor U24271 (N_24271,N_23130,N_23324);
xor U24272 (N_24272,N_23195,N_23136);
nor U24273 (N_24273,N_23281,N_23753);
and U24274 (N_24274,N_23628,N_23003);
nor U24275 (N_24275,N_23944,N_23120);
nor U24276 (N_24276,N_23451,N_23565);
nor U24277 (N_24277,N_23439,N_23805);
or U24278 (N_24278,N_23365,N_23867);
or U24279 (N_24279,N_23679,N_23869);
nor U24280 (N_24280,N_23310,N_23448);
or U24281 (N_24281,N_23474,N_23051);
or U24282 (N_24282,N_23896,N_23540);
xor U24283 (N_24283,N_23261,N_23895);
xor U24284 (N_24284,N_23904,N_23962);
nor U24285 (N_24285,N_23682,N_23425);
nor U24286 (N_24286,N_23563,N_23483);
and U24287 (N_24287,N_23829,N_23924);
nor U24288 (N_24288,N_23665,N_23232);
and U24289 (N_24289,N_23903,N_23876);
and U24290 (N_24290,N_23911,N_23522);
or U24291 (N_24291,N_23512,N_23330);
or U24292 (N_24292,N_23882,N_23062);
xor U24293 (N_24293,N_23157,N_23398);
and U24294 (N_24294,N_23168,N_23937);
xor U24295 (N_24295,N_23968,N_23192);
nand U24296 (N_24296,N_23037,N_23642);
nor U24297 (N_24297,N_23332,N_23627);
nor U24298 (N_24298,N_23982,N_23572);
nand U24299 (N_24299,N_23985,N_23244);
or U24300 (N_24300,N_23416,N_23187);
and U24301 (N_24301,N_23146,N_23902);
nor U24302 (N_24302,N_23173,N_23594);
or U24303 (N_24303,N_23234,N_23065);
xnor U24304 (N_24304,N_23339,N_23735);
nor U24305 (N_24305,N_23325,N_23097);
and U24306 (N_24306,N_23183,N_23334);
nand U24307 (N_24307,N_23597,N_23920);
xor U24308 (N_24308,N_23938,N_23152);
nor U24309 (N_24309,N_23816,N_23678);
nand U24310 (N_24310,N_23504,N_23781);
nor U24311 (N_24311,N_23611,N_23362);
nor U24312 (N_24312,N_23638,N_23422);
xnor U24313 (N_24313,N_23378,N_23082);
or U24314 (N_24314,N_23496,N_23069);
or U24315 (N_24315,N_23868,N_23827);
nand U24316 (N_24316,N_23379,N_23315);
or U24317 (N_24317,N_23009,N_23221);
nand U24318 (N_24318,N_23830,N_23709);
and U24319 (N_24319,N_23137,N_23950);
nand U24320 (N_24320,N_23636,N_23353);
or U24321 (N_24321,N_23359,N_23978);
nor U24322 (N_24322,N_23988,N_23086);
or U24323 (N_24323,N_23258,N_23239);
or U24324 (N_24324,N_23010,N_23624);
xnor U24325 (N_24325,N_23703,N_23124);
nor U24326 (N_24326,N_23622,N_23491);
xnor U24327 (N_24327,N_23226,N_23731);
or U24328 (N_24328,N_23437,N_23209);
or U24329 (N_24329,N_23327,N_23087);
and U24330 (N_24330,N_23208,N_23430);
and U24331 (N_24331,N_23864,N_23329);
or U24332 (N_24332,N_23279,N_23467);
xnor U24333 (N_24333,N_23998,N_23653);
or U24334 (N_24334,N_23384,N_23807);
nor U24335 (N_24335,N_23973,N_23404);
xor U24336 (N_24336,N_23169,N_23029);
and U24337 (N_24337,N_23967,N_23103);
and U24338 (N_24338,N_23047,N_23952);
nor U24339 (N_24339,N_23521,N_23085);
or U24340 (N_24340,N_23718,N_23453);
nor U24341 (N_24341,N_23423,N_23243);
xnor U24342 (N_24342,N_23786,N_23571);
and U24343 (N_24343,N_23321,N_23766);
and U24344 (N_24344,N_23598,N_23768);
or U24345 (N_24345,N_23429,N_23883);
xnor U24346 (N_24346,N_23484,N_23284);
and U24347 (N_24347,N_23028,N_23659);
xor U24348 (N_24348,N_23443,N_23730);
and U24349 (N_24349,N_23468,N_23935);
and U24350 (N_24350,N_23241,N_23278);
nand U24351 (N_24351,N_23414,N_23030);
and U24352 (N_24352,N_23369,N_23271);
or U24353 (N_24353,N_23240,N_23228);
and U24354 (N_24354,N_23341,N_23875);
and U24355 (N_24355,N_23940,N_23856);
nand U24356 (N_24356,N_23728,N_23172);
or U24357 (N_24357,N_23401,N_23955);
or U24358 (N_24358,N_23107,N_23912);
xnor U24359 (N_24359,N_23662,N_23164);
or U24360 (N_24360,N_23110,N_23919);
or U24361 (N_24361,N_23081,N_23336);
nor U24362 (N_24362,N_23223,N_23460);
xnor U24363 (N_24363,N_23052,N_23294);
nand U24364 (N_24364,N_23075,N_23589);
nor U24365 (N_24365,N_23547,N_23536);
nand U24366 (N_24366,N_23251,N_23625);
nor U24367 (N_24367,N_23245,N_23473);
or U24368 (N_24368,N_23049,N_23089);
nand U24369 (N_24369,N_23714,N_23634);
and U24370 (N_24370,N_23619,N_23773);
nand U24371 (N_24371,N_23712,N_23765);
xor U24372 (N_24372,N_23507,N_23144);
or U24373 (N_24373,N_23949,N_23367);
xor U24374 (N_24374,N_23746,N_23396);
xnor U24375 (N_24375,N_23090,N_23135);
and U24376 (N_24376,N_23180,N_23032);
or U24377 (N_24377,N_23845,N_23025);
nor U24378 (N_24378,N_23987,N_23722);
or U24379 (N_24379,N_23262,N_23290);
or U24380 (N_24380,N_23887,N_23694);
nand U24381 (N_24381,N_23806,N_23475);
xnor U24382 (N_24382,N_23802,N_23813);
xnor U24383 (N_24383,N_23555,N_23824);
and U24384 (N_24384,N_23417,N_23351);
or U24385 (N_24385,N_23725,N_23390);
nand U24386 (N_24386,N_23832,N_23972);
nand U24387 (N_24387,N_23263,N_23477);
and U24388 (N_24388,N_23886,N_23742);
nand U24389 (N_24389,N_23538,N_23117);
or U24390 (N_24390,N_23943,N_23771);
or U24391 (N_24391,N_23420,N_23457);
nor U24392 (N_24392,N_23257,N_23534);
or U24393 (N_24393,N_23027,N_23595);
nand U24394 (N_24394,N_23323,N_23963);
xnor U24395 (N_24395,N_23469,N_23939);
or U24396 (N_24396,N_23691,N_23631);
and U24397 (N_24397,N_23031,N_23855);
or U24398 (N_24398,N_23690,N_23568);
or U24399 (N_24399,N_23342,N_23700);
and U24400 (N_24400,N_23979,N_23148);
xor U24401 (N_24401,N_23543,N_23129);
nor U24402 (N_24402,N_23001,N_23331);
nor U24403 (N_24403,N_23206,N_23409);
nor U24404 (N_24404,N_23210,N_23908);
and U24405 (N_24405,N_23668,N_23472);
nand U24406 (N_24406,N_23792,N_23663);
nor U24407 (N_24407,N_23094,N_23162);
or U24408 (N_24408,N_23165,N_23687);
nor U24409 (N_24409,N_23925,N_23111);
and U24410 (N_24410,N_23035,N_23767);
or U24411 (N_24411,N_23175,N_23834);
nand U24412 (N_24412,N_23601,N_23108);
or U24413 (N_24413,N_23661,N_23899);
and U24414 (N_24414,N_23073,N_23225);
and U24415 (N_24415,N_23860,N_23583);
nand U24416 (N_24416,N_23352,N_23161);
nor U24417 (N_24417,N_23113,N_23819);
xor U24418 (N_24418,N_23053,N_23412);
nor U24419 (N_24419,N_23760,N_23708);
nand U24420 (N_24420,N_23093,N_23509);
xor U24421 (N_24421,N_23928,N_23459);
nand U24422 (N_24422,N_23517,N_23440);
nand U24423 (N_24423,N_23326,N_23014);
or U24424 (N_24424,N_23933,N_23424);
nor U24425 (N_24425,N_23020,N_23435);
nor U24426 (N_24426,N_23741,N_23918);
nand U24427 (N_24427,N_23385,N_23458);
and U24428 (N_24428,N_23466,N_23056);
nand U24429 (N_24429,N_23828,N_23480);
and U24430 (N_24430,N_23254,N_23999);
nand U24431 (N_24431,N_23681,N_23651);
nand U24432 (N_24432,N_23400,N_23170);
xnor U24433 (N_24433,N_23482,N_23023);
and U24434 (N_24434,N_23840,N_23286);
nand U24435 (N_24435,N_23872,N_23790);
nor U24436 (N_24436,N_23040,N_23921);
or U24437 (N_24437,N_23397,N_23077);
and U24438 (N_24438,N_23042,N_23516);
and U24439 (N_24439,N_23298,N_23260);
nor U24440 (N_24440,N_23674,N_23012);
or U24441 (N_24441,N_23490,N_23083);
or U24442 (N_24442,N_23948,N_23529);
nand U24443 (N_24443,N_23126,N_23016);
xor U24444 (N_24444,N_23817,N_23635);
nand U24445 (N_24445,N_23442,N_23070);
or U24446 (N_24446,N_23276,N_23317);
or U24447 (N_24447,N_23914,N_23471);
or U24448 (N_24448,N_23889,N_23505);
nand U24449 (N_24449,N_23992,N_23259);
or U24450 (N_24450,N_23877,N_23980);
xor U24451 (N_24451,N_23348,N_23739);
xnor U24452 (N_24452,N_23942,N_23566);
xor U24453 (N_24453,N_23044,N_23582);
and U24454 (N_24454,N_23626,N_23557);
xor U24455 (N_24455,N_23706,N_23382);
xnor U24456 (N_24456,N_23293,N_23045);
nand U24457 (N_24457,N_23163,N_23749);
and U24458 (N_24458,N_23428,N_23076);
nand U24459 (N_24459,N_23763,N_23835);
and U24460 (N_24460,N_23189,N_23809);
xnor U24461 (N_24461,N_23149,N_23667);
nand U24462 (N_24462,N_23433,N_23744);
nor U24463 (N_24463,N_23179,N_23632);
or U24464 (N_24464,N_23269,N_23695);
or U24465 (N_24465,N_23181,N_23851);
nor U24466 (N_24466,N_23142,N_23066);
and U24467 (N_24467,N_23194,N_23692);
xor U24468 (N_24468,N_23986,N_23346);
nor U24469 (N_24469,N_23562,N_23349);
or U24470 (N_24470,N_23450,N_23852);
nand U24471 (N_24471,N_23648,N_23870);
xnor U24472 (N_24472,N_23034,N_23564);
xnor U24473 (N_24473,N_23268,N_23550);
nor U24474 (N_24474,N_23716,N_23127);
nand U24475 (N_24475,N_23650,N_23713);
nand U24476 (N_24476,N_23487,N_23125);
xnor U24477 (N_24477,N_23407,N_23277);
nor U24478 (N_24478,N_23926,N_23637);
nor U24479 (N_24479,N_23657,N_23751);
nand U24480 (N_24480,N_23672,N_23640);
xnor U24481 (N_24481,N_23675,N_23197);
nand U24482 (N_24482,N_23141,N_23726);
nand U24483 (N_24483,N_23599,N_23907);
nor U24484 (N_24484,N_23815,N_23354);
and U24485 (N_24485,N_23646,N_23880);
xnor U24486 (N_24486,N_23669,N_23798);
xnor U24487 (N_24487,N_23917,N_23961);
nand U24488 (N_24488,N_23275,N_23074);
nor U24489 (N_24489,N_23633,N_23196);
xnor U24490 (N_24490,N_23791,N_23363);
or U24491 (N_24491,N_23915,N_23476);
nand U24492 (N_24492,N_23119,N_23738);
or U24493 (N_24493,N_23235,N_23432);
xor U24494 (N_24494,N_23463,N_23590);
xnor U24495 (N_24495,N_23050,N_23038);
nand U24496 (N_24496,N_23402,N_23462);
and U24497 (N_24497,N_23247,N_23530);
xnor U24498 (N_24498,N_23843,N_23006);
or U24499 (N_24499,N_23302,N_23862);
xnor U24500 (N_24500,N_23921,N_23525);
or U24501 (N_24501,N_23419,N_23668);
xnor U24502 (N_24502,N_23022,N_23324);
nor U24503 (N_24503,N_23319,N_23989);
xor U24504 (N_24504,N_23902,N_23547);
nand U24505 (N_24505,N_23333,N_23046);
nand U24506 (N_24506,N_23326,N_23526);
and U24507 (N_24507,N_23761,N_23414);
or U24508 (N_24508,N_23224,N_23795);
xnor U24509 (N_24509,N_23619,N_23398);
xnor U24510 (N_24510,N_23936,N_23696);
nand U24511 (N_24511,N_23638,N_23273);
nor U24512 (N_24512,N_23161,N_23914);
or U24513 (N_24513,N_23341,N_23762);
xnor U24514 (N_24514,N_23267,N_23302);
nand U24515 (N_24515,N_23530,N_23624);
and U24516 (N_24516,N_23681,N_23011);
xnor U24517 (N_24517,N_23637,N_23053);
nand U24518 (N_24518,N_23730,N_23997);
xor U24519 (N_24519,N_23229,N_23786);
or U24520 (N_24520,N_23824,N_23641);
xnor U24521 (N_24521,N_23717,N_23930);
and U24522 (N_24522,N_23461,N_23465);
or U24523 (N_24523,N_23705,N_23090);
or U24524 (N_24524,N_23502,N_23218);
xnor U24525 (N_24525,N_23235,N_23669);
nand U24526 (N_24526,N_23869,N_23409);
xnor U24527 (N_24527,N_23615,N_23778);
or U24528 (N_24528,N_23750,N_23027);
and U24529 (N_24529,N_23206,N_23695);
nor U24530 (N_24530,N_23278,N_23648);
xor U24531 (N_24531,N_23549,N_23595);
and U24532 (N_24532,N_23682,N_23691);
xor U24533 (N_24533,N_23124,N_23677);
xor U24534 (N_24534,N_23635,N_23808);
and U24535 (N_24535,N_23049,N_23757);
nor U24536 (N_24536,N_23273,N_23836);
nor U24537 (N_24537,N_23354,N_23773);
nand U24538 (N_24538,N_23206,N_23245);
and U24539 (N_24539,N_23365,N_23425);
nor U24540 (N_24540,N_23880,N_23126);
or U24541 (N_24541,N_23810,N_23972);
or U24542 (N_24542,N_23523,N_23310);
and U24543 (N_24543,N_23982,N_23084);
xnor U24544 (N_24544,N_23015,N_23654);
nand U24545 (N_24545,N_23947,N_23968);
and U24546 (N_24546,N_23780,N_23547);
nand U24547 (N_24547,N_23573,N_23438);
xor U24548 (N_24548,N_23734,N_23182);
nand U24549 (N_24549,N_23731,N_23974);
nor U24550 (N_24550,N_23333,N_23541);
nor U24551 (N_24551,N_23293,N_23655);
xor U24552 (N_24552,N_23052,N_23152);
nor U24553 (N_24553,N_23704,N_23715);
and U24554 (N_24554,N_23496,N_23969);
nand U24555 (N_24555,N_23068,N_23012);
xor U24556 (N_24556,N_23221,N_23550);
and U24557 (N_24557,N_23912,N_23097);
or U24558 (N_24558,N_23901,N_23165);
xnor U24559 (N_24559,N_23577,N_23455);
nor U24560 (N_24560,N_23273,N_23793);
xnor U24561 (N_24561,N_23945,N_23010);
xnor U24562 (N_24562,N_23654,N_23503);
nor U24563 (N_24563,N_23651,N_23588);
and U24564 (N_24564,N_23487,N_23136);
xor U24565 (N_24565,N_23892,N_23703);
nand U24566 (N_24566,N_23110,N_23541);
and U24567 (N_24567,N_23912,N_23404);
xnor U24568 (N_24568,N_23542,N_23316);
nor U24569 (N_24569,N_23465,N_23080);
and U24570 (N_24570,N_23392,N_23174);
xor U24571 (N_24571,N_23861,N_23659);
nand U24572 (N_24572,N_23717,N_23524);
and U24573 (N_24573,N_23290,N_23654);
xnor U24574 (N_24574,N_23341,N_23114);
xnor U24575 (N_24575,N_23717,N_23161);
nand U24576 (N_24576,N_23029,N_23055);
nor U24577 (N_24577,N_23221,N_23251);
xnor U24578 (N_24578,N_23880,N_23767);
nand U24579 (N_24579,N_23194,N_23058);
and U24580 (N_24580,N_23439,N_23378);
nor U24581 (N_24581,N_23346,N_23356);
and U24582 (N_24582,N_23149,N_23698);
or U24583 (N_24583,N_23237,N_23493);
nor U24584 (N_24584,N_23506,N_23008);
and U24585 (N_24585,N_23612,N_23160);
nand U24586 (N_24586,N_23113,N_23445);
nor U24587 (N_24587,N_23162,N_23194);
nor U24588 (N_24588,N_23194,N_23464);
and U24589 (N_24589,N_23793,N_23732);
or U24590 (N_24590,N_23325,N_23618);
and U24591 (N_24591,N_23827,N_23175);
and U24592 (N_24592,N_23258,N_23036);
nand U24593 (N_24593,N_23424,N_23239);
nand U24594 (N_24594,N_23061,N_23207);
xnor U24595 (N_24595,N_23994,N_23631);
and U24596 (N_24596,N_23696,N_23023);
and U24597 (N_24597,N_23693,N_23456);
and U24598 (N_24598,N_23258,N_23545);
nand U24599 (N_24599,N_23209,N_23317);
xor U24600 (N_24600,N_23081,N_23627);
nor U24601 (N_24601,N_23575,N_23018);
and U24602 (N_24602,N_23392,N_23450);
and U24603 (N_24603,N_23986,N_23319);
nor U24604 (N_24604,N_23702,N_23029);
nor U24605 (N_24605,N_23019,N_23695);
nor U24606 (N_24606,N_23721,N_23412);
nand U24607 (N_24607,N_23237,N_23816);
and U24608 (N_24608,N_23909,N_23541);
xor U24609 (N_24609,N_23950,N_23774);
nand U24610 (N_24610,N_23569,N_23697);
and U24611 (N_24611,N_23652,N_23693);
nor U24612 (N_24612,N_23913,N_23678);
xnor U24613 (N_24613,N_23970,N_23061);
nand U24614 (N_24614,N_23747,N_23199);
nor U24615 (N_24615,N_23556,N_23890);
and U24616 (N_24616,N_23551,N_23310);
nand U24617 (N_24617,N_23186,N_23001);
xnor U24618 (N_24618,N_23659,N_23927);
nand U24619 (N_24619,N_23776,N_23597);
xnor U24620 (N_24620,N_23639,N_23900);
or U24621 (N_24621,N_23417,N_23481);
nand U24622 (N_24622,N_23946,N_23049);
and U24623 (N_24623,N_23149,N_23620);
nor U24624 (N_24624,N_23110,N_23137);
nand U24625 (N_24625,N_23243,N_23340);
nor U24626 (N_24626,N_23892,N_23896);
or U24627 (N_24627,N_23267,N_23509);
xnor U24628 (N_24628,N_23643,N_23067);
xnor U24629 (N_24629,N_23583,N_23419);
and U24630 (N_24630,N_23761,N_23643);
or U24631 (N_24631,N_23872,N_23387);
nor U24632 (N_24632,N_23369,N_23820);
nor U24633 (N_24633,N_23410,N_23008);
and U24634 (N_24634,N_23306,N_23400);
or U24635 (N_24635,N_23117,N_23865);
or U24636 (N_24636,N_23344,N_23816);
or U24637 (N_24637,N_23725,N_23976);
and U24638 (N_24638,N_23851,N_23428);
and U24639 (N_24639,N_23971,N_23881);
and U24640 (N_24640,N_23286,N_23280);
nor U24641 (N_24641,N_23120,N_23173);
and U24642 (N_24642,N_23993,N_23027);
or U24643 (N_24643,N_23452,N_23180);
and U24644 (N_24644,N_23759,N_23711);
nand U24645 (N_24645,N_23702,N_23654);
and U24646 (N_24646,N_23765,N_23340);
xnor U24647 (N_24647,N_23787,N_23888);
xor U24648 (N_24648,N_23743,N_23704);
or U24649 (N_24649,N_23750,N_23265);
nand U24650 (N_24650,N_23585,N_23771);
or U24651 (N_24651,N_23092,N_23578);
xnor U24652 (N_24652,N_23232,N_23611);
or U24653 (N_24653,N_23261,N_23736);
nand U24654 (N_24654,N_23099,N_23792);
and U24655 (N_24655,N_23044,N_23149);
nor U24656 (N_24656,N_23040,N_23114);
or U24657 (N_24657,N_23647,N_23900);
and U24658 (N_24658,N_23094,N_23972);
or U24659 (N_24659,N_23799,N_23669);
and U24660 (N_24660,N_23679,N_23580);
xor U24661 (N_24661,N_23348,N_23312);
xor U24662 (N_24662,N_23128,N_23743);
or U24663 (N_24663,N_23073,N_23320);
nand U24664 (N_24664,N_23379,N_23759);
nor U24665 (N_24665,N_23575,N_23463);
or U24666 (N_24666,N_23507,N_23929);
nand U24667 (N_24667,N_23001,N_23125);
and U24668 (N_24668,N_23870,N_23494);
or U24669 (N_24669,N_23551,N_23603);
and U24670 (N_24670,N_23551,N_23130);
and U24671 (N_24671,N_23534,N_23994);
or U24672 (N_24672,N_23912,N_23687);
and U24673 (N_24673,N_23127,N_23817);
or U24674 (N_24674,N_23663,N_23842);
xor U24675 (N_24675,N_23533,N_23347);
xnor U24676 (N_24676,N_23652,N_23093);
nor U24677 (N_24677,N_23065,N_23721);
and U24678 (N_24678,N_23445,N_23147);
nand U24679 (N_24679,N_23385,N_23443);
nor U24680 (N_24680,N_23229,N_23654);
xnor U24681 (N_24681,N_23573,N_23045);
xor U24682 (N_24682,N_23868,N_23727);
nor U24683 (N_24683,N_23209,N_23925);
and U24684 (N_24684,N_23442,N_23688);
nand U24685 (N_24685,N_23386,N_23193);
xnor U24686 (N_24686,N_23823,N_23401);
nand U24687 (N_24687,N_23114,N_23166);
and U24688 (N_24688,N_23598,N_23322);
nand U24689 (N_24689,N_23730,N_23311);
and U24690 (N_24690,N_23218,N_23353);
nand U24691 (N_24691,N_23576,N_23783);
or U24692 (N_24692,N_23645,N_23058);
nand U24693 (N_24693,N_23894,N_23878);
and U24694 (N_24694,N_23041,N_23352);
nor U24695 (N_24695,N_23750,N_23160);
and U24696 (N_24696,N_23483,N_23413);
or U24697 (N_24697,N_23738,N_23555);
or U24698 (N_24698,N_23657,N_23975);
xnor U24699 (N_24699,N_23436,N_23428);
nand U24700 (N_24700,N_23186,N_23993);
xnor U24701 (N_24701,N_23747,N_23381);
nor U24702 (N_24702,N_23520,N_23160);
and U24703 (N_24703,N_23304,N_23770);
nand U24704 (N_24704,N_23231,N_23192);
or U24705 (N_24705,N_23765,N_23660);
or U24706 (N_24706,N_23763,N_23592);
nand U24707 (N_24707,N_23187,N_23271);
xnor U24708 (N_24708,N_23052,N_23176);
or U24709 (N_24709,N_23044,N_23637);
nor U24710 (N_24710,N_23867,N_23186);
nand U24711 (N_24711,N_23918,N_23579);
xnor U24712 (N_24712,N_23847,N_23696);
and U24713 (N_24713,N_23210,N_23860);
or U24714 (N_24714,N_23748,N_23009);
or U24715 (N_24715,N_23785,N_23809);
nor U24716 (N_24716,N_23697,N_23012);
nor U24717 (N_24717,N_23612,N_23999);
or U24718 (N_24718,N_23523,N_23553);
or U24719 (N_24719,N_23502,N_23268);
nor U24720 (N_24720,N_23293,N_23813);
nor U24721 (N_24721,N_23024,N_23349);
xor U24722 (N_24722,N_23797,N_23806);
nand U24723 (N_24723,N_23070,N_23380);
or U24724 (N_24724,N_23468,N_23976);
xor U24725 (N_24725,N_23860,N_23011);
nand U24726 (N_24726,N_23500,N_23080);
or U24727 (N_24727,N_23604,N_23021);
or U24728 (N_24728,N_23208,N_23752);
nand U24729 (N_24729,N_23782,N_23556);
and U24730 (N_24730,N_23523,N_23676);
nand U24731 (N_24731,N_23694,N_23626);
or U24732 (N_24732,N_23940,N_23310);
and U24733 (N_24733,N_23722,N_23268);
nand U24734 (N_24734,N_23195,N_23263);
and U24735 (N_24735,N_23166,N_23964);
or U24736 (N_24736,N_23838,N_23336);
xnor U24737 (N_24737,N_23094,N_23283);
nand U24738 (N_24738,N_23462,N_23172);
xnor U24739 (N_24739,N_23044,N_23831);
or U24740 (N_24740,N_23229,N_23958);
nor U24741 (N_24741,N_23784,N_23614);
nor U24742 (N_24742,N_23782,N_23815);
nor U24743 (N_24743,N_23817,N_23010);
nand U24744 (N_24744,N_23550,N_23070);
xnor U24745 (N_24745,N_23111,N_23403);
and U24746 (N_24746,N_23590,N_23028);
and U24747 (N_24747,N_23387,N_23890);
nor U24748 (N_24748,N_23481,N_23397);
and U24749 (N_24749,N_23661,N_23750);
or U24750 (N_24750,N_23363,N_23090);
or U24751 (N_24751,N_23459,N_23623);
nor U24752 (N_24752,N_23299,N_23194);
xor U24753 (N_24753,N_23109,N_23081);
xnor U24754 (N_24754,N_23746,N_23740);
or U24755 (N_24755,N_23472,N_23741);
or U24756 (N_24756,N_23709,N_23399);
xnor U24757 (N_24757,N_23294,N_23274);
nand U24758 (N_24758,N_23863,N_23046);
nand U24759 (N_24759,N_23342,N_23285);
or U24760 (N_24760,N_23577,N_23161);
nor U24761 (N_24761,N_23142,N_23925);
xor U24762 (N_24762,N_23788,N_23014);
nand U24763 (N_24763,N_23928,N_23547);
xor U24764 (N_24764,N_23906,N_23354);
and U24765 (N_24765,N_23875,N_23135);
nor U24766 (N_24766,N_23209,N_23999);
nor U24767 (N_24767,N_23231,N_23801);
nor U24768 (N_24768,N_23387,N_23754);
nor U24769 (N_24769,N_23588,N_23549);
nand U24770 (N_24770,N_23819,N_23030);
nor U24771 (N_24771,N_23454,N_23934);
nor U24772 (N_24772,N_23043,N_23136);
xnor U24773 (N_24773,N_23352,N_23107);
nand U24774 (N_24774,N_23866,N_23254);
nor U24775 (N_24775,N_23095,N_23047);
or U24776 (N_24776,N_23713,N_23446);
and U24777 (N_24777,N_23209,N_23305);
nor U24778 (N_24778,N_23027,N_23021);
nor U24779 (N_24779,N_23821,N_23954);
xor U24780 (N_24780,N_23249,N_23716);
xnor U24781 (N_24781,N_23392,N_23635);
or U24782 (N_24782,N_23076,N_23484);
nor U24783 (N_24783,N_23996,N_23440);
and U24784 (N_24784,N_23928,N_23465);
nand U24785 (N_24785,N_23281,N_23136);
or U24786 (N_24786,N_23792,N_23645);
nor U24787 (N_24787,N_23996,N_23160);
or U24788 (N_24788,N_23194,N_23549);
and U24789 (N_24789,N_23498,N_23434);
nor U24790 (N_24790,N_23907,N_23942);
xnor U24791 (N_24791,N_23865,N_23631);
and U24792 (N_24792,N_23439,N_23145);
and U24793 (N_24793,N_23352,N_23047);
nor U24794 (N_24794,N_23558,N_23114);
nor U24795 (N_24795,N_23006,N_23254);
xor U24796 (N_24796,N_23068,N_23172);
or U24797 (N_24797,N_23431,N_23972);
and U24798 (N_24798,N_23367,N_23843);
and U24799 (N_24799,N_23220,N_23447);
or U24800 (N_24800,N_23168,N_23651);
xor U24801 (N_24801,N_23353,N_23015);
nor U24802 (N_24802,N_23747,N_23248);
nor U24803 (N_24803,N_23273,N_23989);
or U24804 (N_24804,N_23052,N_23053);
xnor U24805 (N_24805,N_23585,N_23412);
or U24806 (N_24806,N_23209,N_23938);
xor U24807 (N_24807,N_23696,N_23333);
or U24808 (N_24808,N_23149,N_23592);
or U24809 (N_24809,N_23209,N_23372);
or U24810 (N_24810,N_23377,N_23840);
nand U24811 (N_24811,N_23634,N_23658);
nand U24812 (N_24812,N_23858,N_23368);
xor U24813 (N_24813,N_23139,N_23531);
or U24814 (N_24814,N_23595,N_23934);
and U24815 (N_24815,N_23255,N_23020);
nand U24816 (N_24816,N_23532,N_23653);
nand U24817 (N_24817,N_23753,N_23361);
nand U24818 (N_24818,N_23486,N_23077);
xor U24819 (N_24819,N_23856,N_23131);
and U24820 (N_24820,N_23836,N_23631);
nor U24821 (N_24821,N_23242,N_23501);
nand U24822 (N_24822,N_23954,N_23410);
nand U24823 (N_24823,N_23802,N_23875);
xnor U24824 (N_24824,N_23537,N_23054);
and U24825 (N_24825,N_23786,N_23441);
and U24826 (N_24826,N_23078,N_23177);
and U24827 (N_24827,N_23814,N_23717);
nor U24828 (N_24828,N_23436,N_23890);
nand U24829 (N_24829,N_23027,N_23001);
or U24830 (N_24830,N_23120,N_23711);
and U24831 (N_24831,N_23618,N_23966);
and U24832 (N_24832,N_23070,N_23786);
nand U24833 (N_24833,N_23360,N_23508);
nand U24834 (N_24834,N_23748,N_23951);
xnor U24835 (N_24835,N_23300,N_23129);
and U24836 (N_24836,N_23348,N_23934);
or U24837 (N_24837,N_23505,N_23458);
nand U24838 (N_24838,N_23817,N_23154);
xnor U24839 (N_24839,N_23266,N_23609);
xnor U24840 (N_24840,N_23519,N_23644);
or U24841 (N_24841,N_23254,N_23000);
and U24842 (N_24842,N_23534,N_23604);
and U24843 (N_24843,N_23001,N_23179);
or U24844 (N_24844,N_23240,N_23936);
xor U24845 (N_24845,N_23643,N_23258);
xnor U24846 (N_24846,N_23345,N_23757);
or U24847 (N_24847,N_23480,N_23730);
and U24848 (N_24848,N_23519,N_23259);
nor U24849 (N_24849,N_23060,N_23567);
nor U24850 (N_24850,N_23292,N_23598);
xor U24851 (N_24851,N_23939,N_23341);
or U24852 (N_24852,N_23533,N_23032);
nor U24853 (N_24853,N_23632,N_23957);
nand U24854 (N_24854,N_23480,N_23091);
xnor U24855 (N_24855,N_23742,N_23950);
nand U24856 (N_24856,N_23986,N_23812);
nor U24857 (N_24857,N_23231,N_23302);
nor U24858 (N_24858,N_23930,N_23724);
or U24859 (N_24859,N_23178,N_23155);
or U24860 (N_24860,N_23279,N_23048);
nand U24861 (N_24861,N_23689,N_23872);
and U24862 (N_24862,N_23405,N_23502);
nor U24863 (N_24863,N_23509,N_23505);
and U24864 (N_24864,N_23095,N_23461);
or U24865 (N_24865,N_23354,N_23192);
xnor U24866 (N_24866,N_23800,N_23099);
xnor U24867 (N_24867,N_23698,N_23710);
nand U24868 (N_24868,N_23326,N_23890);
xor U24869 (N_24869,N_23929,N_23208);
xnor U24870 (N_24870,N_23059,N_23883);
and U24871 (N_24871,N_23292,N_23222);
nand U24872 (N_24872,N_23466,N_23065);
or U24873 (N_24873,N_23356,N_23285);
and U24874 (N_24874,N_23591,N_23005);
xnor U24875 (N_24875,N_23310,N_23720);
nand U24876 (N_24876,N_23731,N_23504);
or U24877 (N_24877,N_23653,N_23135);
or U24878 (N_24878,N_23169,N_23126);
xor U24879 (N_24879,N_23488,N_23329);
nor U24880 (N_24880,N_23814,N_23322);
nor U24881 (N_24881,N_23299,N_23833);
nand U24882 (N_24882,N_23119,N_23896);
or U24883 (N_24883,N_23625,N_23951);
nor U24884 (N_24884,N_23149,N_23328);
nand U24885 (N_24885,N_23514,N_23613);
xor U24886 (N_24886,N_23722,N_23327);
or U24887 (N_24887,N_23855,N_23371);
nand U24888 (N_24888,N_23485,N_23963);
xnor U24889 (N_24889,N_23337,N_23622);
nor U24890 (N_24890,N_23593,N_23967);
xor U24891 (N_24891,N_23952,N_23473);
xnor U24892 (N_24892,N_23285,N_23306);
and U24893 (N_24893,N_23236,N_23193);
xor U24894 (N_24894,N_23504,N_23544);
nor U24895 (N_24895,N_23464,N_23039);
or U24896 (N_24896,N_23232,N_23028);
and U24897 (N_24897,N_23519,N_23559);
or U24898 (N_24898,N_23120,N_23527);
or U24899 (N_24899,N_23971,N_23780);
nand U24900 (N_24900,N_23274,N_23375);
nor U24901 (N_24901,N_23807,N_23603);
nand U24902 (N_24902,N_23994,N_23603);
and U24903 (N_24903,N_23501,N_23450);
xnor U24904 (N_24904,N_23880,N_23113);
and U24905 (N_24905,N_23911,N_23386);
nand U24906 (N_24906,N_23285,N_23719);
xor U24907 (N_24907,N_23286,N_23309);
xor U24908 (N_24908,N_23822,N_23770);
and U24909 (N_24909,N_23295,N_23354);
xor U24910 (N_24910,N_23971,N_23013);
xnor U24911 (N_24911,N_23145,N_23112);
xnor U24912 (N_24912,N_23868,N_23378);
and U24913 (N_24913,N_23581,N_23006);
nor U24914 (N_24914,N_23785,N_23003);
or U24915 (N_24915,N_23253,N_23708);
nor U24916 (N_24916,N_23913,N_23860);
xor U24917 (N_24917,N_23408,N_23761);
and U24918 (N_24918,N_23972,N_23182);
xor U24919 (N_24919,N_23786,N_23277);
nand U24920 (N_24920,N_23846,N_23579);
and U24921 (N_24921,N_23648,N_23375);
nand U24922 (N_24922,N_23366,N_23885);
nor U24923 (N_24923,N_23493,N_23374);
and U24924 (N_24924,N_23033,N_23573);
or U24925 (N_24925,N_23826,N_23775);
or U24926 (N_24926,N_23273,N_23106);
nand U24927 (N_24927,N_23823,N_23229);
nand U24928 (N_24928,N_23659,N_23088);
and U24929 (N_24929,N_23486,N_23573);
or U24930 (N_24930,N_23139,N_23477);
or U24931 (N_24931,N_23933,N_23732);
and U24932 (N_24932,N_23883,N_23311);
and U24933 (N_24933,N_23883,N_23326);
nand U24934 (N_24934,N_23891,N_23000);
nand U24935 (N_24935,N_23324,N_23181);
xnor U24936 (N_24936,N_23872,N_23475);
or U24937 (N_24937,N_23245,N_23153);
nor U24938 (N_24938,N_23091,N_23712);
and U24939 (N_24939,N_23007,N_23691);
nand U24940 (N_24940,N_23667,N_23990);
nor U24941 (N_24941,N_23540,N_23703);
nand U24942 (N_24942,N_23859,N_23488);
or U24943 (N_24943,N_23283,N_23004);
nand U24944 (N_24944,N_23367,N_23519);
nor U24945 (N_24945,N_23309,N_23700);
nor U24946 (N_24946,N_23566,N_23251);
and U24947 (N_24947,N_23215,N_23996);
and U24948 (N_24948,N_23654,N_23586);
xnor U24949 (N_24949,N_23482,N_23146);
or U24950 (N_24950,N_23634,N_23833);
and U24951 (N_24951,N_23373,N_23174);
nor U24952 (N_24952,N_23964,N_23516);
nand U24953 (N_24953,N_23830,N_23656);
or U24954 (N_24954,N_23520,N_23552);
or U24955 (N_24955,N_23611,N_23344);
xor U24956 (N_24956,N_23847,N_23535);
or U24957 (N_24957,N_23686,N_23895);
nand U24958 (N_24958,N_23834,N_23079);
nand U24959 (N_24959,N_23877,N_23848);
nand U24960 (N_24960,N_23844,N_23829);
nor U24961 (N_24961,N_23847,N_23614);
and U24962 (N_24962,N_23990,N_23059);
or U24963 (N_24963,N_23270,N_23018);
nand U24964 (N_24964,N_23932,N_23808);
nand U24965 (N_24965,N_23403,N_23935);
or U24966 (N_24966,N_23019,N_23319);
and U24967 (N_24967,N_23326,N_23793);
nand U24968 (N_24968,N_23227,N_23544);
xnor U24969 (N_24969,N_23163,N_23450);
or U24970 (N_24970,N_23261,N_23795);
nand U24971 (N_24971,N_23259,N_23770);
or U24972 (N_24972,N_23479,N_23889);
or U24973 (N_24973,N_23542,N_23689);
and U24974 (N_24974,N_23605,N_23270);
or U24975 (N_24975,N_23188,N_23323);
nor U24976 (N_24976,N_23723,N_23344);
or U24977 (N_24977,N_23457,N_23640);
xnor U24978 (N_24978,N_23801,N_23305);
and U24979 (N_24979,N_23442,N_23643);
nor U24980 (N_24980,N_23060,N_23295);
and U24981 (N_24981,N_23990,N_23816);
nor U24982 (N_24982,N_23964,N_23570);
and U24983 (N_24983,N_23713,N_23919);
or U24984 (N_24984,N_23295,N_23055);
and U24985 (N_24985,N_23668,N_23200);
xor U24986 (N_24986,N_23002,N_23936);
nand U24987 (N_24987,N_23761,N_23412);
and U24988 (N_24988,N_23688,N_23855);
and U24989 (N_24989,N_23317,N_23357);
nor U24990 (N_24990,N_23951,N_23520);
nor U24991 (N_24991,N_23437,N_23460);
and U24992 (N_24992,N_23080,N_23867);
and U24993 (N_24993,N_23281,N_23175);
nand U24994 (N_24994,N_23139,N_23217);
xor U24995 (N_24995,N_23128,N_23908);
xnor U24996 (N_24996,N_23429,N_23956);
xnor U24997 (N_24997,N_23067,N_23376);
nor U24998 (N_24998,N_23359,N_23775);
xor U24999 (N_24999,N_23014,N_23328);
nand UO_0 (O_0,N_24816,N_24213);
nand UO_1 (O_1,N_24212,N_24087);
or UO_2 (O_2,N_24695,N_24219);
nor UO_3 (O_3,N_24413,N_24454);
nor UO_4 (O_4,N_24957,N_24655);
xor UO_5 (O_5,N_24833,N_24676);
nand UO_6 (O_6,N_24656,N_24943);
xor UO_7 (O_7,N_24503,N_24110);
xnor UO_8 (O_8,N_24600,N_24201);
or UO_9 (O_9,N_24462,N_24348);
nand UO_10 (O_10,N_24877,N_24936);
nand UO_11 (O_11,N_24968,N_24135);
nand UO_12 (O_12,N_24370,N_24962);
xnor UO_13 (O_13,N_24838,N_24295);
nor UO_14 (O_14,N_24054,N_24419);
and UO_15 (O_15,N_24183,N_24689);
or UO_16 (O_16,N_24312,N_24132);
or UO_17 (O_17,N_24210,N_24849);
nor UO_18 (O_18,N_24176,N_24262);
and UO_19 (O_19,N_24377,N_24100);
and UO_20 (O_20,N_24860,N_24128);
and UO_21 (O_21,N_24037,N_24512);
or UO_22 (O_22,N_24828,N_24829);
nand UO_23 (O_23,N_24387,N_24440);
xor UO_24 (O_24,N_24195,N_24354);
and UO_25 (O_25,N_24938,N_24151);
or UO_26 (O_26,N_24892,N_24079);
nor UO_27 (O_27,N_24720,N_24126);
nor UO_28 (O_28,N_24520,N_24424);
xor UO_29 (O_29,N_24493,N_24014);
and UO_30 (O_30,N_24191,N_24193);
nand UO_31 (O_31,N_24198,N_24248);
and UO_32 (O_32,N_24606,N_24867);
xnor UO_33 (O_33,N_24729,N_24551);
or UO_34 (O_34,N_24330,N_24525);
nor UO_35 (O_35,N_24663,N_24708);
xor UO_36 (O_36,N_24147,N_24499);
and UO_37 (O_37,N_24064,N_24451);
nor UO_38 (O_38,N_24339,N_24133);
nand UO_39 (O_39,N_24721,N_24716);
or UO_40 (O_40,N_24445,N_24306);
or UO_41 (O_41,N_24743,N_24659);
nor UO_42 (O_42,N_24966,N_24360);
and UO_43 (O_43,N_24935,N_24987);
and UO_44 (O_44,N_24225,N_24020);
nor UO_45 (O_45,N_24001,N_24332);
nand UO_46 (O_46,N_24947,N_24202);
and UO_47 (O_47,N_24486,N_24215);
and UO_48 (O_48,N_24915,N_24406);
nand UO_49 (O_49,N_24336,N_24157);
nand UO_50 (O_50,N_24232,N_24632);
nor UO_51 (O_51,N_24956,N_24178);
or UO_52 (O_52,N_24502,N_24245);
nor UO_53 (O_53,N_24378,N_24608);
and UO_54 (O_54,N_24182,N_24316);
nand UO_55 (O_55,N_24362,N_24224);
or UO_56 (O_56,N_24047,N_24887);
or UO_57 (O_57,N_24572,N_24866);
and UO_58 (O_58,N_24679,N_24702);
nand UO_59 (O_59,N_24117,N_24587);
nor UO_60 (O_60,N_24643,N_24408);
or UO_61 (O_61,N_24142,N_24226);
or UO_62 (O_62,N_24562,N_24620);
or UO_63 (O_63,N_24648,N_24603);
or UO_64 (O_64,N_24640,N_24837);
or UO_65 (O_65,N_24429,N_24030);
xor UO_66 (O_66,N_24988,N_24565);
xor UO_67 (O_67,N_24750,N_24083);
nor UO_68 (O_68,N_24379,N_24251);
xnor UO_69 (O_69,N_24733,N_24961);
and UO_70 (O_70,N_24143,N_24438);
nand UO_71 (O_71,N_24196,N_24651);
or UO_72 (O_72,N_24170,N_24003);
nor UO_73 (O_73,N_24229,N_24421);
xnor UO_74 (O_74,N_24150,N_24952);
or UO_75 (O_75,N_24310,N_24214);
xor UO_76 (O_76,N_24888,N_24650);
nand UO_77 (O_77,N_24570,N_24343);
or UO_78 (O_78,N_24762,N_24818);
or UO_79 (O_79,N_24169,N_24531);
and UO_80 (O_80,N_24560,N_24945);
nor UO_81 (O_81,N_24744,N_24735);
nor UO_82 (O_82,N_24345,N_24841);
or UO_83 (O_83,N_24356,N_24825);
xnor UO_84 (O_84,N_24712,N_24159);
xnor UO_85 (O_85,N_24862,N_24472);
nand UO_86 (O_86,N_24386,N_24917);
xnor UO_87 (O_87,N_24745,N_24417);
or UO_88 (O_88,N_24254,N_24645);
nand UO_89 (O_89,N_24878,N_24446);
and UO_90 (O_90,N_24719,N_24497);
nor UO_91 (O_91,N_24094,N_24216);
or UO_92 (O_92,N_24477,N_24246);
xor UO_93 (O_93,N_24209,N_24573);
xor UO_94 (O_94,N_24673,N_24097);
xnor UO_95 (O_95,N_24998,N_24685);
nor UO_96 (O_96,N_24494,N_24532);
xor UO_97 (O_97,N_24607,N_24510);
xnor UO_98 (O_98,N_24690,N_24358);
nand UO_99 (O_99,N_24767,N_24846);
xor UO_100 (O_100,N_24626,N_24882);
nor UO_101 (O_101,N_24010,N_24827);
nor UO_102 (O_102,N_24309,N_24042);
nor UO_103 (O_103,N_24918,N_24537);
and UO_104 (O_104,N_24925,N_24488);
nor UO_105 (O_105,N_24806,N_24324);
nor UO_106 (O_106,N_24292,N_24969);
nor UO_107 (O_107,N_24990,N_24124);
xor UO_108 (O_108,N_24435,N_24768);
nor UO_109 (O_109,N_24630,N_24016);
and UO_110 (O_110,N_24028,N_24759);
or UO_111 (O_111,N_24145,N_24638);
nor UO_112 (O_112,N_24253,N_24705);
or UO_113 (O_113,N_24048,N_24017);
or UO_114 (O_114,N_24807,N_24299);
and UO_115 (O_115,N_24623,N_24696);
nor UO_116 (O_116,N_24403,N_24092);
xnor UO_117 (O_117,N_24662,N_24088);
nand UO_118 (O_118,N_24830,N_24980);
nor UO_119 (O_119,N_24505,N_24973);
nand UO_120 (O_120,N_24993,N_24265);
nor UO_121 (O_121,N_24060,N_24029);
or UO_122 (O_122,N_24670,N_24948);
nand UO_123 (O_123,N_24025,N_24612);
xnor UO_124 (O_124,N_24863,N_24163);
or UO_125 (O_125,N_24236,N_24121);
and UO_126 (O_126,N_24709,N_24044);
nor UO_127 (O_127,N_24465,N_24153);
or UO_128 (O_128,N_24350,N_24749);
and UO_129 (O_129,N_24884,N_24235);
nor UO_130 (O_130,N_24864,N_24976);
xnor UO_131 (O_131,N_24255,N_24563);
nor UO_132 (O_132,N_24813,N_24741);
nand UO_133 (O_133,N_24574,N_24528);
xnor UO_134 (O_134,N_24313,N_24155);
and UO_135 (O_135,N_24858,N_24504);
or UO_136 (O_136,N_24450,N_24747);
nand UO_137 (O_137,N_24007,N_24937);
and UO_138 (O_138,N_24949,N_24898);
nor UO_139 (O_139,N_24444,N_24637);
and UO_140 (O_140,N_24461,N_24642);
or UO_141 (O_141,N_24542,N_24012);
or UO_142 (O_142,N_24548,N_24901);
xnor UO_143 (O_143,N_24649,N_24822);
or UO_144 (O_144,N_24301,N_24715);
nor UO_145 (O_145,N_24861,N_24974);
nand UO_146 (O_146,N_24188,N_24853);
xnor UO_147 (O_147,N_24355,N_24646);
xor UO_148 (O_148,N_24774,N_24801);
nor UO_149 (O_149,N_24794,N_24052);
xnor UO_150 (O_150,N_24068,N_24033);
xnor UO_151 (O_151,N_24114,N_24189);
and UO_152 (O_152,N_24983,N_24487);
nand UO_153 (O_153,N_24283,N_24041);
or UO_154 (O_154,N_24431,N_24000);
xor UO_155 (O_155,N_24826,N_24383);
nor UO_156 (O_156,N_24286,N_24290);
nor UO_157 (O_157,N_24700,N_24367);
xnor UO_158 (O_158,N_24372,N_24035);
nor UO_159 (O_159,N_24293,N_24534);
xor UO_160 (O_160,N_24591,N_24739);
and UO_161 (O_161,N_24032,N_24181);
or UO_162 (O_162,N_24628,N_24156);
nand UO_163 (O_163,N_24070,N_24970);
xor UO_164 (O_164,N_24889,N_24799);
xnor UO_165 (O_165,N_24162,N_24845);
and UO_166 (O_166,N_24361,N_24624);
nand UO_167 (O_167,N_24996,N_24699);
nand UO_168 (O_168,N_24771,N_24883);
xnor UO_169 (O_169,N_24785,N_24912);
nor UO_170 (O_170,N_24929,N_24731);
xnor UO_171 (O_171,N_24644,N_24868);
xnor UO_172 (O_172,N_24168,N_24434);
nand UO_173 (O_173,N_24404,N_24277);
nor UO_174 (O_174,N_24491,N_24895);
nand UO_175 (O_175,N_24276,N_24071);
xor UO_176 (O_176,N_24755,N_24844);
xnor UO_177 (O_177,N_24578,N_24796);
xor UO_178 (O_178,N_24713,N_24141);
or UO_179 (O_179,N_24508,N_24927);
nor UO_180 (O_180,N_24385,N_24577);
nor UO_181 (O_181,N_24390,N_24242);
xor UO_182 (O_182,N_24601,N_24122);
nand UO_183 (O_183,N_24500,N_24803);
or UO_184 (O_184,N_24284,N_24264);
or UO_185 (O_185,N_24058,N_24125);
nand UO_186 (O_186,N_24180,N_24647);
and UO_187 (O_187,N_24258,N_24657);
xnor UO_188 (O_188,N_24568,N_24507);
nor UO_189 (O_189,N_24757,N_24102);
xor UO_190 (O_190,N_24791,N_24104);
nand UO_191 (O_191,N_24772,N_24108);
nor UO_192 (O_192,N_24074,N_24409);
or UO_193 (O_193,N_24204,N_24266);
and UO_194 (O_194,N_24789,N_24013);
or UO_195 (O_195,N_24763,N_24069);
or UO_196 (O_196,N_24540,N_24631);
nor UO_197 (O_197,N_24992,N_24682);
xor UO_198 (O_198,N_24296,N_24834);
nor UO_199 (O_199,N_24959,N_24559);
or UO_200 (O_200,N_24096,N_24430);
or UO_201 (O_201,N_24683,N_24405);
nand UO_202 (O_202,N_24045,N_24769);
nor UO_203 (O_203,N_24984,N_24474);
xor UO_204 (O_204,N_24321,N_24775);
xor UO_205 (O_205,N_24717,N_24802);
or UO_206 (O_206,N_24896,N_24549);
nand UO_207 (O_207,N_24809,N_24515);
nand UO_208 (O_208,N_24804,N_24134);
and UO_209 (O_209,N_24395,N_24842);
nand UO_210 (O_210,N_24773,N_24399);
nor UO_211 (O_211,N_24365,N_24363);
nor UO_212 (O_212,N_24684,N_24514);
xor UO_213 (O_213,N_24614,N_24252);
and UO_214 (O_214,N_24031,N_24397);
nand UO_215 (O_215,N_24185,N_24975);
or UO_216 (O_216,N_24851,N_24919);
nor UO_217 (O_217,N_24872,N_24402);
or UO_218 (O_218,N_24920,N_24285);
nand UO_219 (O_219,N_24075,N_24111);
and UO_220 (O_220,N_24432,N_24589);
or UO_221 (O_221,N_24051,N_24439);
xor UO_222 (O_222,N_24605,N_24304);
nor UO_223 (O_223,N_24393,N_24173);
nor UO_224 (O_224,N_24584,N_24061);
and UO_225 (O_225,N_24536,N_24315);
or UO_226 (O_226,N_24109,N_24597);
nor UO_227 (O_227,N_24453,N_24701);
or UO_228 (O_228,N_24939,N_24473);
xnor UO_229 (O_229,N_24906,N_24672);
nor UO_230 (O_230,N_24724,N_24334);
xor UO_231 (O_231,N_24800,N_24687);
and UO_232 (O_232,N_24243,N_24057);
and UO_233 (O_233,N_24291,N_24160);
nor UO_234 (O_234,N_24999,N_24373);
and UO_235 (O_235,N_24857,N_24698);
and UO_236 (O_236,N_24981,N_24275);
nand UO_237 (O_237,N_24119,N_24184);
or UO_238 (O_238,N_24036,N_24227);
xor UO_239 (O_239,N_24836,N_24478);
xor UO_240 (O_240,N_24940,N_24049);
xor UO_241 (O_241,N_24349,N_24220);
and UO_242 (O_242,N_24617,N_24871);
or UO_243 (O_243,N_24022,N_24848);
or UO_244 (O_244,N_24524,N_24737);
xor UO_245 (O_245,N_24040,N_24269);
nor UO_246 (O_246,N_24810,N_24839);
and UO_247 (O_247,N_24783,N_24821);
nand UO_248 (O_248,N_24986,N_24034);
and UO_249 (O_249,N_24665,N_24634);
and UO_250 (O_250,N_24059,N_24703);
xor UO_251 (O_251,N_24197,N_24519);
xnor UO_252 (O_252,N_24798,N_24261);
nor UO_253 (O_253,N_24278,N_24723);
nor UO_254 (O_254,N_24411,N_24043);
or UO_255 (O_255,N_24137,N_24944);
nand UO_256 (O_256,N_24222,N_24812);
and UO_257 (O_257,N_24099,N_24758);
or UO_258 (O_258,N_24538,N_24658);
xnor UO_259 (O_259,N_24116,N_24610);
nand UO_260 (O_260,N_24543,N_24481);
and UO_261 (O_261,N_24091,N_24009);
and UO_262 (O_262,N_24641,N_24442);
and UO_263 (O_263,N_24599,N_24078);
and UO_264 (O_264,N_24625,N_24619);
nor UO_265 (O_265,N_24139,N_24470);
and UO_266 (O_266,N_24904,N_24571);
nor UO_267 (O_267,N_24566,N_24922);
or UO_268 (O_268,N_24995,N_24778);
and UO_269 (O_269,N_24675,N_24297);
nor UO_270 (O_270,N_24298,N_24722);
or UO_271 (O_271,N_24340,N_24257);
nand UO_272 (O_272,N_24250,N_24464);
or UO_273 (O_273,N_24084,N_24526);
xor UO_274 (O_274,N_24865,N_24847);
or UO_275 (O_275,N_24903,N_24376);
nor UO_276 (O_276,N_24893,N_24105);
xnor UO_277 (O_277,N_24518,N_24979);
and UO_278 (O_278,N_24437,N_24931);
nand UO_279 (O_279,N_24130,N_24909);
xor UO_280 (O_280,N_24471,N_24433);
and UO_281 (O_281,N_24530,N_24516);
or UO_282 (O_282,N_24582,N_24282);
nand UO_283 (O_283,N_24660,N_24886);
xnor UO_284 (O_284,N_24653,N_24148);
nor UO_285 (O_285,N_24192,N_24186);
nor UO_286 (O_286,N_24027,N_24460);
and UO_287 (O_287,N_24575,N_24598);
nor UO_288 (O_288,N_24905,N_24666);
nor UO_289 (O_289,N_24602,N_24899);
nand UO_290 (O_290,N_24545,N_24950);
xor UO_291 (O_291,N_24954,N_24326);
or UO_292 (O_292,N_24671,N_24635);
and UO_293 (O_293,N_24609,N_24509);
and UO_294 (O_294,N_24484,N_24955);
or UO_295 (O_295,N_24077,N_24900);
nand UO_296 (O_296,N_24555,N_24468);
nor UO_297 (O_297,N_24873,N_24629);
or UO_298 (O_298,N_24318,N_24098);
and UO_299 (O_299,N_24171,N_24407);
xor UO_300 (O_300,N_24693,N_24483);
and UO_301 (O_301,N_24311,N_24476);
and UO_302 (O_302,N_24754,N_24455);
xnor UO_303 (O_303,N_24550,N_24859);
xor UO_304 (O_304,N_24815,N_24890);
nor UO_305 (O_305,N_24113,N_24753);
nand UO_306 (O_306,N_24053,N_24305);
xnor UO_307 (O_307,N_24015,N_24174);
or UO_308 (O_308,N_24932,N_24303);
or UO_309 (O_309,N_24581,N_24725);
and UO_310 (O_310,N_24492,N_24885);
nor UO_311 (O_311,N_24357,N_24633);
or UO_312 (O_312,N_24347,N_24050);
xnor UO_313 (O_313,N_24691,N_24006);
and UO_314 (O_314,N_24780,N_24556);
xor UO_315 (O_315,N_24002,N_24466);
and UO_316 (O_316,N_24239,N_24211);
or UO_317 (O_317,N_24814,N_24485);
xor UO_318 (O_318,N_24770,N_24856);
nor UO_319 (O_319,N_24718,N_24140);
and UO_320 (O_320,N_24469,N_24971);
or UO_321 (O_321,N_24172,N_24958);
or UO_322 (O_322,N_24752,N_24942);
nand UO_323 (O_323,N_24392,N_24941);
nor UO_324 (O_324,N_24164,N_24618);
or UO_325 (O_325,N_24661,N_24797);
nand UO_326 (O_326,N_24207,N_24686);
and UO_327 (O_327,N_24322,N_24654);
or UO_328 (O_328,N_24366,N_24965);
nand UO_329 (O_329,N_24274,N_24557);
and UO_330 (O_330,N_24482,N_24681);
xor UO_331 (O_331,N_24613,N_24677);
or UO_332 (O_332,N_24089,N_24736);
and UO_333 (O_333,N_24782,N_24793);
nand UO_334 (O_334,N_24329,N_24928);
and UO_335 (O_335,N_24400,N_24320);
and UO_336 (O_336,N_24694,N_24490);
nor UO_337 (O_337,N_24820,N_24746);
nand UO_338 (O_338,N_24384,N_24832);
nor UO_339 (O_339,N_24926,N_24951);
xnor UO_340 (O_340,N_24817,N_24389);
and UO_341 (O_341,N_24217,N_24418);
and UO_342 (O_342,N_24586,N_24289);
nor UO_343 (O_343,N_24055,N_24038);
nor UO_344 (O_344,N_24790,N_24811);
xnor UO_345 (O_345,N_24452,N_24267);
and UO_346 (O_346,N_24594,N_24314);
nor UO_347 (O_347,N_24416,N_24412);
xor UO_348 (O_348,N_24154,N_24428);
or UO_349 (O_349,N_24776,N_24233);
nand UO_350 (O_350,N_24081,N_24333);
nand UO_351 (O_351,N_24697,N_24175);
nand UO_352 (O_352,N_24457,N_24344);
and UO_353 (O_353,N_24260,N_24131);
and UO_354 (O_354,N_24891,N_24127);
xnor UO_355 (O_355,N_24398,N_24352);
nor UO_356 (O_356,N_24161,N_24281);
or UO_357 (O_357,N_24910,N_24732);
and UO_358 (O_358,N_24240,N_24766);
and UO_359 (O_359,N_24394,N_24371);
and UO_360 (O_360,N_24544,N_24639);
nand UO_361 (O_361,N_24369,N_24103);
xor UO_362 (O_362,N_24115,N_24177);
nor UO_363 (O_363,N_24447,N_24669);
and UO_364 (O_364,N_24436,N_24535);
and UO_365 (O_365,N_24341,N_24692);
nand UO_366 (O_366,N_24396,N_24280);
and UO_367 (O_367,N_24095,N_24082);
or UO_368 (O_368,N_24353,N_24710);
and UO_369 (O_369,N_24787,N_24908);
and UO_370 (O_370,N_24415,N_24541);
nor UO_371 (O_371,N_24480,N_24467);
nor UO_372 (O_372,N_24085,N_24921);
and UO_373 (O_373,N_24066,N_24138);
or UO_374 (O_374,N_24228,N_24441);
and UO_375 (O_375,N_24533,N_24026);
nor UO_376 (O_376,N_24914,N_24167);
xnor UO_377 (O_377,N_24580,N_24761);
xnor UO_378 (O_378,N_24569,N_24011);
xor UO_379 (O_379,N_24337,N_24667);
nand UO_380 (O_380,N_24711,N_24596);
and UO_381 (O_381,N_24426,N_24259);
nor UO_382 (O_382,N_24706,N_24263);
xnor UO_383 (O_383,N_24786,N_24760);
xor UO_384 (O_384,N_24997,N_24223);
and UO_385 (O_385,N_24205,N_24982);
xnor UO_386 (O_386,N_24558,N_24805);
or UO_387 (O_387,N_24496,N_24852);
and UO_388 (O_388,N_24230,N_24123);
or UO_389 (O_389,N_24740,N_24985);
nand UO_390 (O_390,N_24475,N_24527);
nand UO_391 (O_391,N_24427,N_24734);
xnor UO_392 (O_392,N_24994,N_24756);
nand UO_393 (O_393,N_24552,N_24101);
and UO_394 (O_394,N_24933,N_24351);
nor UO_395 (O_395,N_24149,N_24989);
or UO_396 (O_396,N_24458,N_24194);
xor UO_397 (O_397,N_24136,N_24200);
xnor UO_398 (O_398,N_24112,N_24547);
nor UO_399 (O_399,N_24420,N_24788);
and UO_400 (O_400,N_24924,N_24005);
and UO_401 (O_401,N_24072,N_24593);
nor UO_402 (O_402,N_24425,N_24414);
nand UO_403 (O_403,N_24792,N_24585);
and UO_404 (O_404,N_24063,N_24726);
and UO_405 (O_405,N_24463,N_24271);
and UO_406 (O_406,N_24241,N_24875);
or UO_407 (O_407,N_24869,N_24328);
and UO_408 (O_408,N_24765,N_24479);
or UO_409 (O_409,N_24907,N_24308);
and UO_410 (O_410,N_24590,N_24728);
nand UO_411 (O_411,N_24894,N_24080);
and UO_412 (O_412,N_24916,N_24152);
xor UO_413 (O_413,N_24179,N_24325);
or UO_414 (O_414,N_24093,N_24678);
xor UO_415 (O_415,N_24364,N_24576);
xnor UO_416 (O_416,N_24777,N_24090);
and UO_417 (O_417,N_24972,N_24779);
xor UO_418 (O_418,N_24021,N_24268);
and UO_419 (O_419,N_24338,N_24714);
xor UO_420 (O_420,N_24317,N_24382);
xnor UO_421 (O_421,N_24323,N_24065);
and UO_422 (O_422,N_24023,N_24621);
or UO_423 (O_423,N_24840,N_24302);
nand UO_424 (O_424,N_24674,N_24237);
or UO_425 (O_425,N_24616,N_24489);
nand UO_426 (O_426,N_24203,N_24008);
xnor UO_427 (O_427,N_24118,N_24521);
or UO_428 (O_428,N_24062,N_24165);
nand UO_429 (O_429,N_24876,N_24206);
or UO_430 (O_430,N_24652,N_24234);
nand UO_431 (O_431,N_24501,N_24346);
nor UO_432 (O_432,N_24579,N_24897);
nand UO_433 (O_433,N_24748,N_24391);
nand UO_434 (O_434,N_24448,N_24707);
or UO_435 (O_435,N_24381,N_24056);
nand UO_436 (O_436,N_24960,N_24583);
xnor UO_437 (O_437,N_24300,N_24129);
or UO_438 (O_438,N_24554,N_24208);
or UO_439 (O_439,N_24553,N_24247);
nor UO_440 (O_440,N_24902,N_24604);
nand UO_441 (O_441,N_24688,N_24930);
nand UO_442 (O_442,N_24374,N_24146);
nand UO_443 (O_443,N_24668,N_24881);
xor UO_444 (O_444,N_24221,N_24561);
and UO_445 (O_445,N_24879,N_24244);
or UO_446 (O_446,N_24564,N_24368);
xnor UO_447 (O_447,N_24018,N_24158);
nand UO_448 (O_448,N_24727,N_24636);
or UO_449 (O_449,N_24459,N_24106);
nand UO_450 (O_450,N_24513,N_24611);
or UO_451 (O_451,N_24456,N_24964);
and UO_452 (O_452,N_24190,N_24319);
nor UO_453 (O_453,N_24076,N_24449);
nor UO_454 (O_454,N_24850,N_24107);
nand UO_455 (O_455,N_24831,N_24854);
nand UO_456 (O_456,N_24627,N_24279);
or UO_457 (O_457,N_24067,N_24764);
nor UO_458 (O_458,N_24231,N_24855);
nor UO_459 (O_459,N_24923,N_24978);
or UO_460 (O_460,N_24819,N_24967);
nor UO_461 (O_461,N_24946,N_24784);
and UO_462 (O_462,N_24567,N_24307);
or UO_463 (O_463,N_24511,N_24934);
nor UO_464 (O_464,N_24664,N_24911);
nor UO_465 (O_465,N_24294,N_24187);
nand UO_466 (O_466,N_24529,N_24120);
nand UO_467 (O_467,N_24288,N_24824);
nor UO_468 (O_468,N_24730,N_24073);
and UO_469 (O_469,N_24588,N_24218);
and UO_470 (O_470,N_24270,N_24823);
nand UO_471 (O_471,N_24751,N_24327);
nor UO_472 (O_472,N_24615,N_24046);
and UO_473 (O_473,N_24795,N_24517);
and UO_474 (O_474,N_24287,N_24238);
or UO_475 (O_475,N_24401,N_24019);
nand UO_476 (O_476,N_24273,N_24144);
or UO_477 (O_477,N_24506,N_24249);
xnor UO_478 (O_478,N_24522,N_24375);
nor UO_479 (O_479,N_24977,N_24704);
nor UO_480 (O_480,N_24595,N_24256);
xnor UO_481 (O_481,N_24880,N_24742);
xor UO_482 (O_482,N_24843,N_24592);
and UO_483 (O_483,N_24808,N_24953);
xor UO_484 (O_484,N_24272,N_24331);
and UO_485 (O_485,N_24039,N_24335);
and UO_486 (O_486,N_24342,N_24835);
or UO_487 (O_487,N_24546,N_24024);
and UO_488 (O_488,N_24539,N_24086);
nand UO_489 (O_489,N_24622,N_24199);
xor UO_490 (O_490,N_24004,N_24874);
xnor UO_491 (O_491,N_24680,N_24498);
and UO_492 (O_492,N_24443,N_24410);
or UO_493 (O_493,N_24991,N_24738);
nor UO_494 (O_494,N_24963,N_24870);
nand UO_495 (O_495,N_24166,N_24781);
xnor UO_496 (O_496,N_24913,N_24422);
or UO_497 (O_497,N_24388,N_24523);
or UO_498 (O_498,N_24359,N_24380);
or UO_499 (O_499,N_24423,N_24495);
or UO_500 (O_500,N_24755,N_24769);
nor UO_501 (O_501,N_24529,N_24232);
nor UO_502 (O_502,N_24377,N_24564);
nand UO_503 (O_503,N_24394,N_24750);
nand UO_504 (O_504,N_24528,N_24568);
and UO_505 (O_505,N_24023,N_24628);
or UO_506 (O_506,N_24346,N_24465);
xor UO_507 (O_507,N_24853,N_24516);
and UO_508 (O_508,N_24207,N_24053);
or UO_509 (O_509,N_24727,N_24765);
xnor UO_510 (O_510,N_24829,N_24755);
and UO_511 (O_511,N_24023,N_24844);
nor UO_512 (O_512,N_24709,N_24067);
and UO_513 (O_513,N_24527,N_24105);
or UO_514 (O_514,N_24808,N_24626);
or UO_515 (O_515,N_24559,N_24299);
nor UO_516 (O_516,N_24301,N_24353);
and UO_517 (O_517,N_24142,N_24342);
and UO_518 (O_518,N_24083,N_24801);
nand UO_519 (O_519,N_24791,N_24050);
nor UO_520 (O_520,N_24650,N_24700);
nand UO_521 (O_521,N_24286,N_24029);
or UO_522 (O_522,N_24109,N_24889);
nor UO_523 (O_523,N_24289,N_24554);
and UO_524 (O_524,N_24334,N_24917);
or UO_525 (O_525,N_24015,N_24308);
or UO_526 (O_526,N_24896,N_24265);
nand UO_527 (O_527,N_24125,N_24025);
and UO_528 (O_528,N_24222,N_24837);
xnor UO_529 (O_529,N_24487,N_24497);
xor UO_530 (O_530,N_24172,N_24237);
or UO_531 (O_531,N_24527,N_24315);
nand UO_532 (O_532,N_24362,N_24713);
nand UO_533 (O_533,N_24094,N_24633);
xnor UO_534 (O_534,N_24237,N_24181);
xor UO_535 (O_535,N_24428,N_24178);
nor UO_536 (O_536,N_24893,N_24067);
or UO_537 (O_537,N_24314,N_24615);
and UO_538 (O_538,N_24828,N_24962);
or UO_539 (O_539,N_24015,N_24037);
nor UO_540 (O_540,N_24142,N_24811);
or UO_541 (O_541,N_24026,N_24831);
or UO_542 (O_542,N_24235,N_24909);
nand UO_543 (O_543,N_24077,N_24314);
xnor UO_544 (O_544,N_24051,N_24105);
nand UO_545 (O_545,N_24416,N_24141);
nor UO_546 (O_546,N_24449,N_24430);
nand UO_547 (O_547,N_24656,N_24413);
xor UO_548 (O_548,N_24466,N_24695);
nor UO_549 (O_549,N_24511,N_24303);
and UO_550 (O_550,N_24129,N_24757);
or UO_551 (O_551,N_24935,N_24898);
nor UO_552 (O_552,N_24754,N_24766);
or UO_553 (O_553,N_24626,N_24704);
or UO_554 (O_554,N_24571,N_24084);
nor UO_555 (O_555,N_24558,N_24803);
or UO_556 (O_556,N_24122,N_24098);
and UO_557 (O_557,N_24035,N_24699);
xor UO_558 (O_558,N_24711,N_24364);
or UO_559 (O_559,N_24840,N_24609);
nand UO_560 (O_560,N_24762,N_24189);
and UO_561 (O_561,N_24041,N_24186);
xnor UO_562 (O_562,N_24070,N_24607);
nand UO_563 (O_563,N_24151,N_24708);
xor UO_564 (O_564,N_24314,N_24574);
xor UO_565 (O_565,N_24549,N_24819);
xnor UO_566 (O_566,N_24322,N_24577);
or UO_567 (O_567,N_24202,N_24055);
and UO_568 (O_568,N_24268,N_24739);
xor UO_569 (O_569,N_24928,N_24296);
nor UO_570 (O_570,N_24901,N_24776);
nand UO_571 (O_571,N_24856,N_24754);
nand UO_572 (O_572,N_24029,N_24077);
xor UO_573 (O_573,N_24165,N_24752);
or UO_574 (O_574,N_24828,N_24407);
nand UO_575 (O_575,N_24245,N_24539);
xnor UO_576 (O_576,N_24598,N_24456);
nor UO_577 (O_577,N_24318,N_24841);
xnor UO_578 (O_578,N_24061,N_24858);
or UO_579 (O_579,N_24656,N_24788);
or UO_580 (O_580,N_24480,N_24302);
nor UO_581 (O_581,N_24639,N_24365);
nor UO_582 (O_582,N_24695,N_24519);
xnor UO_583 (O_583,N_24850,N_24327);
and UO_584 (O_584,N_24844,N_24912);
nor UO_585 (O_585,N_24338,N_24495);
nor UO_586 (O_586,N_24967,N_24520);
or UO_587 (O_587,N_24975,N_24328);
xor UO_588 (O_588,N_24735,N_24474);
xor UO_589 (O_589,N_24512,N_24549);
nand UO_590 (O_590,N_24394,N_24528);
xnor UO_591 (O_591,N_24983,N_24809);
nand UO_592 (O_592,N_24920,N_24412);
nand UO_593 (O_593,N_24035,N_24278);
or UO_594 (O_594,N_24172,N_24399);
nand UO_595 (O_595,N_24578,N_24933);
or UO_596 (O_596,N_24336,N_24299);
or UO_597 (O_597,N_24680,N_24700);
nand UO_598 (O_598,N_24977,N_24626);
xnor UO_599 (O_599,N_24796,N_24494);
or UO_600 (O_600,N_24937,N_24911);
xnor UO_601 (O_601,N_24905,N_24545);
xnor UO_602 (O_602,N_24751,N_24206);
or UO_603 (O_603,N_24117,N_24803);
nor UO_604 (O_604,N_24209,N_24345);
or UO_605 (O_605,N_24405,N_24447);
nor UO_606 (O_606,N_24598,N_24373);
or UO_607 (O_607,N_24952,N_24964);
nand UO_608 (O_608,N_24645,N_24081);
and UO_609 (O_609,N_24012,N_24176);
nor UO_610 (O_610,N_24372,N_24490);
nor UO_611 (O_611,N_24936,N_24504);
and UO_612 (O_612,N_24578,N_24309);
nand UO_613 (O_613,N_24852,N_24350);
nand UO_614 (O_614,N_24494,N_24615);
nand UO_615 (O_615,N_24028,N_24957);
or UO_616 (O_616,N_24352,N_24179);
xnor UO_617 (O_617,N_24329,N_24316);
xor UO_618 (O_618,N_24108,N_24010);
xor UO_619 (O_619,N_24775,N_24670);
and UO_620 (O_620,N_24947,N_24211);
nand UO_621 (O_621,N_24189,N_24633);
xnor UO_622 (O_622,N_24445,N_24348);
or UO_623 (O_623,N_24370,N_24935);
or UO_624 (O_624,N_24191,N_24988);
xor UO_625 (O_625,N_24523,N_24889);
nand UO_626 (O_626,N_24036,N_24981);
nor UO_627 (O_627,N_24375,N_24656);
and UO_628 (O_628,N_24975,N_24731);
and UO_629 (O_629,N_24510,N_24587);
xor UO_630 (O_630,N_24576,N_24421);
and UO_631 (O_631,N_24989,N_24349);
and UO_632 (O_632,N_24727,N_24507);
xor UO_633 (O_633,N_24873,N_24834);
xor UO_634 (O_634,N_24284,N_24020);
xor UO_635 (O_635,N_24424,N_24149);
or UO_636 (O_636,N_24080,N_24435);
or UO_637 (O_637,N_24516,N_24583);
or UO_638 (O_638,N_24796,N_24277);
and UO_639 (O_639,N_24392,N_24662);
nand UO_640 (O_640,N_24503,N_24026);
and UO_641 (O_641,N_24419,N_24621);
nor UO_642 (O_642,N_24534,N_24393);
nand UO_643 (O_643,N_24788,N_24268);
nand UO_644 (O_644,N_24426,N_24816);
nor UO_645 (O_645,N_24010,N_24513);
nand UO_646 (O_646,N_24305,N_24517);
nand UO_647 (O_647,N_24107,N_24870);
or UO_648 (O_648,N_24384,N_24495);
xor UO_649 (O_649,N_24942,N_24508);
and UO_650 (O_650,N_24272,N_24150);
or UO_651 (O_651,N_24541,N_24145);
xnor UO_652 (O_652,N_24499,N_24724);
nand UO_653 (O_653,N_24478,N_24607);
and UO_654 (O_654,N_24682,N_24901);
nand UO_655 (O_655,N_24858,N_24606);
nor UO_656 (O_656,N_24328,N_24823);
or UO_657 (O_657,N_24995,N_24899);
or UO_658 (O_658,N_24023,N_24632);
nand UO_659 (O_659,N_24110,N_24468);
and UO_660 (O_660,N_24499,N_24339);
nor UO_661 (O_661,N_24642,N_24494);
nand UO_662 (O_662,N_24552,N_24176);
nand UO_663 (O_663,N_24300,N_24077);
nor UO_664 (O_664,N_24800,N_24152);
or UO_665 (O_665,N_24618,N_24593);
and UO_666 (O_666,N_24504,N_24663);
or UO_667 (O_667,N_24035,N_24204);
and UO_668 (O_668,N_24064,N_24774);
xnor UO_669 (O_669,N_24178,N_24402);
nor UO_670 (O_670,N_24601,N_24063);
nand UO_671 (O_671,N_24300,N_24731);
nor UO_672 (O_672,N_24933,N_24345);
or UO_673 (O_673,N_24442,N_24372);
or UO_674 (O_674,N_24468,N_24339);
xor UO_675 (O_675,N_24129,N_24252);
xor UO_676 (O_676,N_24288,N_24053);
nand UO_677 (O_677,N_24447,N_24283);
or UO_678 (O_678,N_24224,N_24504);
and UO_679 (O_679,N_24440,N_24819);
and UO_680 (O_680,N_24705,N_24111);
nand UO_681 (O_681,N_24431,N_24580);
nand UO_682 (O_682,N_24173,N_24611);
and UO_683 (O_683,N_24677,N_24481);
nand UO_684 (O_684,N_24063,N_24250);
nor UO_685 (O_685,N_24694,N_24398);
nor UO_686 (O_686,N_24687,N_24530);
xnor UO_687 (O_687,N_24315,N_24044);
nand UO_688 (O_688,N_24561,N_24964);
nand UO_689 (O_689,N_24136,N_24711);
nand UO_690 (O_690,N_24281,N_24810);
nor UO_691 (O_691,N_24879,N_24306);
or UO_692 (O_692,N_24525,N_24792);
xnor UO_693 (O_693,N_24913,N_24570);
and UO_694 (O_694,N_24950,N_24815);
and UO_695 (O_695,N_24397,N_24752);
nand UO_696 (O_696,N_24548,N_24831);
xor UO_697 (O_697,N_24957,N_24078);
or UO_698 (O_698,N_24357,N_24390);
or UO_699 (O_699,N_24147,N_24069);
xnor UO_700 (O_700,N_24828,N_24212);
or UO_701 (O_701,N_24835,N_24381);
nor UO_702 (O_702,N_24986,N_24239);
and UO_703 (O_703,N_24069,N_24863);
or UO_704 (O_704,N_24341,N_24610);
and UO_705 (O_705,N_24351,N_24189);
xnor UO_706 (O_706,N_24935,N_24679);
xor UO_707 (O_707,N_24762,N_24450);
nand UO_708 (O_708,N_24271,N_24483);
and UO_709 (O_709,N_24193,N_24021);
xor UO_710 (O_710,N_24247,N_24766);
and UO_711 (O_711,N_24042,N_24930);
and UO_712 (O_712,N_24631,N_24160);
and UO_713 (O_713,N_24158,N_24759);
xnor UO_714 (O_714,N_24690,N_24830);
or UO_715 (O_715,N_24574,N_24151);
nand UO_716 (O_716,N_24452,N_24175);
and UO_717 (O_717,N_24301,N_24405);
nand UO_718 (O_718,N_24916,N_24893);
or UO_719 (O_719,N_24798,N_24217);
nand UO_720 (O_720,N_24518,N_24040);
nand UO_721 (O_721,N_24605,N_24521);
nand UO_722 (O_722,N_24746,N_24791);
nand UO_723 (O_723,N_24124,N_24654);
nor UO_724 (O_724,N_24877,N_24841);
or UO_725 (O_725,N_24255,N_24558);
xor UO_726 (O_726,N_24304,N_24434);
nor UO_727 (O_727,N_24364,N_24749);
nor UO_728 (O_728,N_24784,N_24697);
and UO_729 (O_729,N_24238,N_24529);
xnor UO_730 (O_730,N_24704,N_24267);
nor UO_731 (O_731,N_24639,N_24559);
nand UO_732 (O_732,N_24960,N_24629);
and UO_733 (O_733,N_24139,N_24618);
xnor UO_734 (O_734,N_24305,N_24492);
or UO_735 (O_735,N_24668,N_24189);
and UO_736 (O_736,N_24584,N_24462);
nor UO_737 (O_737,N_24761,N_24268);
nand UO_738 (O_738,N_24163,N_24840);
xor UO_739 (O_739,N_24427,N_24742);
nand UO_740 (O_740,N_24097,N_24956);
and UO_741 (O_741,N_24774,N_24714);
and UO_742 (O_742,N_24413,N_24702);
or UO_743 (O_743,N_24225,N_24369);
nor UO_744 (O_744,N_24445,N_24387);
and UO_745 (O_745,N_24161,N_24397);
or UO_746 (O_746,N_24230,N_24969);
or UO_747 (O_747,N_24269,N_24171);
and UO_748 (O_748,N_24885,N_24645);
or UO_749 (O_749,N_24620,N_24911);
or UO_750 (O_750,N_24548,N_24083);
nor UO_751 (O_751,N_24607,N_24905);
or UO_752 (O_752,N_24611,N_24399);
nor UO_753 (O_753,N_24277,N_24611);
and UO_754 (O_754,N_24776,N_24873);
or UO_755 (O_755,N_24132,N_24015);
nor UO_756 (O_756,N_24591,N_24966);
nand UO_757 (O_757,N_24398,N_24085);
xor UO_758 (O_758,N_24282,N_24831);
and UO_759 (O_759,N_24997,N_24236);
xor UO_760 (O_760,N_24631,N_24831);
nand UO_761 (O_761,N_24177,N_24844);
nor UO_762 (O_762,N_24418,N_24577);
nand UO_763 (O_763,N_24359,N_24672);
or UO_764 (O_764,N_24633,N_24394);
nor UO_765 (O_765,N_24104,N_24529);
nand UO_766 (O_766,N_24210,N_24528);
and UO_767 (O_767,N_24425,N_24627);
nand UO_768 (O_768,N_24836,N_24687);
xor UO_769 (O_769,N_24215,N_24502);
nor UO_770 (O_770,N_24252,N_24932);
nor UO_771 (O_771,N_24537,N_24742);
nor UO_772 (O_772,N_24253,N_24163);
nor UO_773 (O_773,N_24002,N_24902);
and UO_774 (O_774,N_24496,N_24510);
nor UO_775 (O_775,N_24831,N_24851);
and UO_776 (O_776,N_24272,N_24982);
xor UO_777 (O_777,N_24914,N_24220);
and UO_778 (O_778,N_24418,N_24690);
nor UO_779 (O_779,N_24470,N_24570);
nor UO_780 (O_780,N_24749,N_24017);
and UO_781 (O_781,N_24181,N_24069);
or UO_782 (O_782,N_24296,N_24265);
or UO_783 (O_783,N_24453,N_24242);
or UO_784 (O_784,N_24643,N_24883);
nor UO_785 (O_785,N_24239,N_24528);
nor UO_786 (O_786,N_24499,N_24073);
nor UO_787 (O_787,N_24074,N_24510);
nor UO_788 (O_788,N_24633,N_24412);
nand UO_789 (O_789,N_24361,N_24439);
nand UO_790 (O_790,N_24786,N_24150);
xnor UO_791 (O_791,N_24647,N_24588);
nand UO_792 (O_792,N_24308,N_24894);
xor UO_793 (O_793,N_24033,N_24621);
nand UO_794 (O_794,N_24406,N_24823);
and UO_795 (O_795,N_24642,N_24255);
or UO_796 (O_796,N_24748,N_24790);
xnor UO_797 (O_797,N_24043,N_24395);
xnor UO_798 (O_798,N_24183,N_24550);
xnor UO_799 (O_799,N_24667,N_24929);
nor UO_800 (O_800,N_24597,N_24813);
nor UO_801 (O_801,N_24323,N_24249);
and UO_802 (O_802,N_24458,N_24147);
nand UO_803 (O_803,N_24489,N_24584);
and UO_804 (O_804,N_24473,N_24966);
or UO_805 (O_805,N_24552,N_24797);
or UO_806 (O_806,N_24022,N_24387);
and UO_807 (O_807,N_24333,N_24053);
and UO_808 (O_808,N_24541,N_24190);
nand UO_809 (O_809,N_24318,N_24230);
nand UO_810 (O_810,N_24698,N_24697);
nor UO_811 (O_811,N_24125,N_24972);
xnor UO_812 (O_812,N_24945,N_24944);
and UO_813 (O_813,N_24187,N_24356);
nand UO_814 (O_814,N_24326,N_24098);
or UO_815 (O_815,N_24927,N_24998);
nor UO_816 (O_816,N_24775,N_24965);
xnor UO_817 (O_817,N_24793,N_24285);
nor UO_818 (O_818,N_24671,N_24932);
nand UO_819 (O_819,N_24804,N_24507);
and UO_820 (O_820,N_24377,N_24480);
or UO_821 (O_821,N_24937,N_24724);
nor UO_822 (O_822,N_24612,N_24507);
nand UO_823 (O_823,N_24292,N_24591);
or UO_824 (O_824,N_24960,N_24877);
xnor UO_825 (O_825,N_24947,N_24730);
or UO_826 (O_826,N_24922,N_24145);
xor UO_827 (O_827,N_24883,N_24252);
xnor UO_828 (O_828,N_24239,N_24597);
xor UO_829 (O_829,N_24023,N_24412);
and UO_830 (O_830,N_24610,N_24105);
or UO_831 (O_831,N_24598,N_24931);
or UO_832 (O_832,N_24788,N_24293);
nand UO_833 (O_833,N_24778,N_24467);
and UO_834 (O_834,N_24091,N_24203);
or UO_835 (O_835,N_24686,N_24973);
nor UO_836 (O_836,N_24771,N_24708);
xor UO_837 (O_837,N_24171,N_24625);
nor UO_838 (O_838,N_24269,N_24716);
xor UO_839 (O_839,N_24680,N_24835);
nand UO_840 (O_840,N_24760,N_24854);
or UO_841 (O_841,N_24036,N_24650);
and UO_842 (O_842,N_24685,N_24263);
and UO_843 (O_843,N_24670,N_24517);
or UO_844 (O_844,N_24762,N_24115);
nor UO_845 (O_845,N_24393,N_24145);
nor UO_846 (O_846,N_24437,N_24729);
xor UO_847 (O_847,N_24422,N_24815);
nor UO_848 (O_848,N_24394,N_24012);
nor UO_849 (O_849,N_24817,N_24165);
or UO_850 (O_850,N_24229,N_24537);
and UO_851 (O_851,N_24848,N_24339);
and UO_852 (O_852,N_24107,N_24079);
nor UO_853 (O_853,N_24193,N_24972);
nor UO_854 (O_854,N_24800,N_24913);
and UO_855 (O_855,N_24665,N_24801);
nor UO_856 (O_856,N_24569,N_24886);
xnor UO_857 (O_857,N_24867,N_24318);
xnor UO_858 (O_858,N_24466,N_24986);
nand UO_859 (O_859,N_24769,N_24825);
or UO_860 (O_860,N_24670,N_24574);
xor UO_861 (O_861,N_24576,N_24973);
nor UO_862 (O_862,N_24699,N_24436);
and UO_863 (O_863,N_24823,N_24717);
or UO_864 (O_864,N_24411,N_24808);
xnor UO_865 (O_865,N_24604,N_24194);
xor UO_866 (O_866,N_24728,N_24610);
or UO_867 (O_867,N_24809,N_24688);
and UO_868 (O_868,N_24577,N_24918);
and UO_869 (O_869,N_24414,N_24339);
nand UO_870 (O_870,N_24985,N_24642);
xor UO_871 (O_871,N_24617,N_24038);
nand UO_872 (O_872,N_24195,N_24614);
and UO_873 (O_873,N_24700,N_24964);
xor UO_874 (O_874,N_24834,N_24376);
xor UO_875 (O_875,N_24313,N_24389);
nand UO_876 (O_876,N_24847,N_24959);
and UO_877 (O_877,N_24932,N_24098);
nand UO_878 (O_878,N_24556,N_24345);
nand UO_879 (O_879,N_24902,N_24416);
nand UO_880 (O_880,N_24432,N_24866);
nor UO_881 (O_881,N_24833,N_24825);
or UO_882 (O_882,N_24516,N_24548);
nor UO_883 (O_883,N_24076,N_24603);
nor UO_884 (O_884,N_24818,N_24565);
or UO_885 (O_885,N_24097,N_24578);
and UO_886 (O_886,N_24437,N_24276);
and UO_887 (O_887,N_24773,N_24247);
nor UO_888 (O_888,N_24972,N_24249);
or UO_889 (O_889,N_24861,N_24549);
nor UO_890 (O_890,N_24986,N_24246);
nand UO_891 (O_891,N_24638,N_24293);
or UO_892 (O_892,N_24141,N_24315);
and UO_893 (O_893,N_24272,N_24864);
xnor UO_894 (O_894,N_24496,N_24843);
nand UO_895 (O_895,N_24592,N_24105);
xnor UO_896 (O_896,N_24887,N_24226);
xnor UO_897 (O_897,N_24907,N_24337);
and UO_898 (O_898,N_24651,N_24775);
or UO_899 (O_899,N_24743,N_24800);
nand UO_900 (O_900,N_24745,N_24259);
xor UO_901 (O_901,N_24480,N_24968);
and UO_902 (O_902,N_24651,N_24866);
nor UO_903 (O_903,N_24606,N_24441);
nor UO_904 (O_904,N_24100,N_24886);
or UO_905 (O_905,N_24496,N_24700);
xnor UO_906 (O_906,N_24766,N_24710);
nor UO_907 (O_907,N_24050,N_24624);
nand UO_908 (O_908,N_24988,N_24439);
and UO_909 (O_909,N_24764,N_24568);
nand UO_910 (O_910,N_24694,N_24591);
nor UO_911 (O_911,N_24184,N_24085);
nor UO_912 (O_912,N_24821,N_24323);
nand UO_913 (O_913,N_24144,N_24984);
xnor UO_914 (O_914,N_24395,N_24502);
nand UO_915 (O_915,N_24480,N_24405);
nand UO_916 (O_916,N_24696,N_24032);
or UO_917 (O_917,N_24500,N_24508);
xnor UO_918 (O_918,N_24559,N_24773);
or UO_919 (O_919,N_24816,N_24916);
nand UO_920 (O_920,N_24257,N_24629);
or UO_921 (O_921,N_24088,N_24638);
or UO_922 (O_922,N_24274,N_24457);
and UO_923 (O_923,N_24813,N_24349);
xor UO_924 (O_924,N_24453,N_24715);
nand UO_925 (O_925,N_24288,N_24902);
nor UO_926 (O_926,N_24023,N_24689);
nor UO_927 (O_927,N_24595,N_24915);
xnor UO_928 (O_928,N_24802,N_24304);
nand UO_929 (O_929,N_24663,N_24368);
and UO_930 (O_930,N_24589,N_24152);
nand UO_931 (O_931,N_24739,N_24074);
and UO_932 (O_932,N_24478,N_24833);
nand UO_933 (O_933,N_24465,N_24630);
nor UO_934 (O_934,N_24146,N_24448);
xnor UO_935 (O_935,N_24317,N_24521);
and UO_936 (O_936,N_24991,N_24600);
xnor UO_937 (O_937,N_24846,N_24200);
xnor UO_938 (O_938,N_24366,N_24714);
nand UO_939 (O_939,N_24044,N_24310);
and UO_940 (O_940,N_24026,N_24024);
xnor UO_941 (O_941,N_24501,N_24714);
and UO_942 (O_942,N_24588,N_24936);
nor UO_943 (O_943,N_24977,N_24949);
and UO_944 (O_944,N_24757,N_24153);
nand UO_945 (O_945,N_24224,N_24921);
or UO_946 (O_946,N_24483,N_24206);
nand UO_947 (O_947,N_24975,N_24143);
xnor UO_948 (O_948,N_24446,N_24545);
and UO_949 (O_949,N_24613,N_24816);
nor UO_950 (O_950,N_24682,N_24206);
xnor UO_951 (O_951,N_24496,N_24228);
nor UO_952 (O_952,N_24022,N_24108);
nand UO_953 (O_953,N_24658,N_24192);
and UO_954 (O_954,N_24547,N_24054);
nor UO_955 (O_955,N_24745,N_24292);
xor UO_956 (O_956,N_24368,N_24196);
and UO_957 (O_957,N_24600,N_24997);
and UO_958 (O_958,N_24778,N_24587);
and UO_959 (O_959,N_24709,N_24634);
xnor UO_960 (O_960,N_24052,N_24806);
or UO_961 (O_961,N_24056,N_24011);
nor UO_962 (O_962,N_24336,N_24994);
or UO_963 (O_963,N_24418,N_24375);
nor UO_964 (O_964,N_24497,N_24604);
nor UO_965 (O_965,N_24039,N_24873);
and UO_966 (O_966,N_24529,N_24295);
or UO_967 (O_967,N_24318,N_24729);
nand UO_968 (O_968,N_24804,N_24381);
and UO_969 (O_969,N_24711,N_24991);
nand UO_970 (O_970,N_24196,N_24452);
xor UO_971 (O_971,N_24601,N_24347);
nand UO_972 (O_972,N_24839,N_24498);
nor UO_973 (O_973,N_24766,N_24592);
nor UO_974 (O_974,N_24934,N_24803);
or UO_975 (O_975,N_24001,N_24693);
nand UO_976 (O_976,N_24349,N_24192);
xor UO_977 (O_977,N_24383,N_24213);
nand UO_978 (O_978,N_24869,N_24044);
and UO_979 (O_979,N_24695,N_24427);
nor UO_980 (O_980,N_24724,N_24357);
nand UO_981 (O_981,N_24357,N_24929);
nor UO_982 (O_982,N_24805,N_24133);
xnor UO_983 (O_983,N_24242,N_24108);
nand UO_984 (O_984,N_24527,N_24926);
xnor UO_985 (O_985,N_24443,N_24905);
nand UO_986 (O_986,N_24292,N_24090);
or UO_987 (O_987,N_24644,N_24945);
nor UO_988 (O_988,N_24512,N_24644);
or UO_989 (O_989,N_24384,N_24547);
and UO_990 (O_990,N_24235,N_24039);
or UO_991 (O_991,N_24810,N_24727);
and UO_992 (O_992,N_24868,N_24875);
or UO_993 (O_993,N_24054,N_24082);
or UO_994 (O_994,N_24212,N_24044);
or UO_995 (O_995,N_24228,N_24297);
xor UO_996 (O_996,N_24899,N_24808);
nand UO_997 (O_997,N_24613,N_24237);
nand UO_998 (O_998,N_24471,N_24212);
nand UO_999 (O_999,N_24457,N_24188);
nand UO_1000 (O_1000,N_24655,N_24217);
and UO_1001 (O_1001,N_24476,N_24038);
nor UO_1002 (O_1002,N_24512,N_24868);
nand UO_1003 (O_1003,N_24516,N_24382);
xor UO_1004 (O_1004,N_24374,N_24326);
xor UO_1005 (O_1005,N_24515,N_24833);
nand UO_1006 (O_1006,N_24243,N_24044);
and UO_1007 (O_1007,N_24990,N_24776);
xnor UO_1008 (O_1008,N_24764,N_24222);
nor UO_1009 (O_1009,N_24691,N_24632);
and UO_1010 (O_1010,N_24976,N_24066);
nor UO_1011 (O_1011,N_24343,N_24358);
nand UO_1012 (O_1012,N_24803,N_24787);
nand UO_1013 (O_1013,N_24182,N_24480);
and UO_1014 (O_1014,N_24844,N_24120);
or UO_1015 (O_1015,N_24181,N_24723);
or UO_1016 (O_1016,N_24034,N_24530);
and UO_1017 (O_1017,N_24305,N_24042);
nor UO_1018 (O_1018,N_24359,N_24214);
and UO_1019 (O_1019,N_24190,N_24562);
nand UO_1020 (O_1020,N_24594,N_24466);
nor UO_1021 (O_1021,N_24655,N_24973);
xor UO_1022 (O_1022,N_24577,N_24675);
xor UO_1023 (O_1023,N_24978,N_24710);
nand UO_1024 (O_1024,N_24690,N_24663);
nand UO_1025 (O_1025,N_24692,N_24080);
xor UO_1026 (O_1026,N_24587,N_24212);
nand UO_1027 (O_1027,N_24141,N_24378);
nor UO_1028 (O_1028,N_24481,N_24547);
or UO_1029 (O_1029,N_24107,N_24698);
nand UO_1030 (O_1030,N_24253,N_24464);
xor UO_1031 (O_1031,N_24271,N_24630);
and UO_1032 (O_1032,N_24971,N_24581);
nand UO_1033 (O_1033,N_24749,N_24998);
xor UO_1034 (O_1034,N_24869,N_24480);
or UO_1035 (O_1035,N_24184,N_24622);
nor UO_1036 (O_1036,N_24194,N_24893);
xor UO_1037 (O_1037,N_24721,N_24093);
nand UO_1038 (O_1038,N_24821,N_24353);
nor UO_1039 (O_1039,N_24370,N_24764);
or UO_1040 (O_1040,N_24156,N_24027);
nand UO_1041 (O_1041,N_24723,N_24040);
xor UO_1042 (O_1042,N_24901,N_24900);
nor UO_1043 (O_1043,N_24711,N_24537);
xnor UO_1044 (O_1044,N_24885,N_24435);
and UO_1045 (O_1045,N_24068,N_24043);
or UO_1046 (O_1046,N_24279,N_24264);
and UO_1047 (O_1047,N_24966,N_24342);
nor UO_1048 (O_1048,N_24054,N_24896);
and UO_1049 (O_1049,N_24763,N_24119);
or UO_1050 (O_1050,N_24371,N_24879);
and UO_1051 (O_1051,N_24698,N_24137);
nand UO_1052 (O_1052,N_24554,N_24935);
nand UO_1053 (O_1053,N_24920,N_24145);
and UO_1054 (O_1054,N_24813,N_24389);
nor UO_1055 (O_1055,N_24772,N_24955);
nor UO_1056 (O_1056,N_24175,N_24307);
or UO_1057 (O_1057,N_24672,N_24313);
or UO_1058 (O_1058,N_24069,N_24644);
or UO_1059 (O_1059,N_24182,N_24984);
or UO_1060 (O_1060,N_24345,N_24412);
and UO_1061 (O_1061,N_24438,N_24542);
nor UO_1062 (O_1062,N_24645,N_24495);
nand UO_1063 (O_1063,N_24430,N_24059);
nor UO_1064 (O_1064,N_24169,N_24602);
and UO_1065 (O_1065,N_24095,N_24478);
and UO_1066 (O_1066,N_24173,N_24154);
nand UO_1067 (O_1067,N_24081,N_24079);
and UO_1068 (O_1068,N_24804,N_24145);
nor UO_1069 (O_1069,N_24554,N_24450);
xnor UO_1070 (O_1070,N_24985,N_24261);
nor UO_1071 (O_1071,N_24193,N_24840);
nor UO_1072 (O_1072,N_24240,N_24551);
nor UO_1073 (O_1073,N_24775,N_24188);
and UO_1074 (O_1074,N_24481,N_24912);
and UO_1075 (O_1075,N_24074,N_24398);
xnor UO_1076 (O_1076,N_24108,N_24106);
nand UO_1077 (O_1077,N_24174,N_24687);
and UO_1078 (O_1078,N_24445,N_24680);
xor UO_1079 (O_1079,N_24128,N_24926);
nor UO_1080 (O_1080,N_24027,N_24616);
nor UO_1081 (O_1081,N_24117,N_24606);
or UO_1082 (O_1082,N_24724,N_24748);
or UO_1083 (O_1083,N_24600,N_24915);
and UO_1084 (O_1084,N_24076,N_24947);
and UO_1085 (O_1085,N_24276,N_24187);
and UO_1086 (O_1086,N_24399,N_24851);
or UO_1087 (O_1087,N_24538,N_24068);
nand UO_1088 (O_1088,N_24142,N_24589);
nand UO_1089 (O_1089,N_24779,N_24451);
or UO_1090 (O_1090,N_24576,N_24297);
nor UO_1091 (O_1091,N_24464,N_24194);
xnor UO_1092 (O_1092,N_24498,N_24457);
nor UO_1093 (O_1093,N_24851,N_24766);
or UO_1094 (O_1094,N_24110,N_24032);
nor UO_1095 (O_1095,N_24836,N_24430);
and UO_1096 (O_1096,N_24698,N_24378);
nand UO_1097 (O_1097,N_24670,N_24772);
nor UO_1098 (O_1098,N_24129,N_24019);
xnor UO_1099 (O_1099,N_24716,N_24562);
and UO_1100 (O_1100,N_24720,N_24030);
and UO_1101 (O_1101,N_24530,N_24884);
and UO_1102 (O_1102,N_24722,N_24499);
or UO_1103 (O_1103,N_24855,N_24323);
or UO_1104 (O_1104,N_24589,N_24327);
and UO_1105 (O_1105,N_24429,N_24784);
and UO_1106 (O_1106,N_24419,N_24078);
nor UO_1107 (O_1107,N_24382,N_24426);
and UO_1108 (O_1108,N_24983,N_24678);
nand UO_1109 (O_1109,N_24791,N_24671);
nand UO_1110 (O_1110,N_24764,N_24913);
and UO_1111 (O_1111,N_24089,N_24480);
and UO_1112 (O_1112,N_24388,N_24565);
nor UO_1113 (O_1113,N_24739,N_24044);
xor UO_1114 (O_1114,N_24305,N_24859);
nor UO_1115 (O_1115,N_24344,N_24796);
or UO_1116 (O_1116,N_24668,N_24622);
nand UO_1117 (O_1117,N_24167,N_24800);
or UO_1118 (O_1118,N_24641,N_24325);
nand UO_1119 (O_1119,N_24445,N_24323);
or UO_1120 (O_1120,N_24826,N_24530);
or UO_1121 (O_1121,N_24430,N_24652);
nand UO_1122 (O_1122,N_24907,N_24138);
xor UO_1123 (O_1123,N_24168,N_24447);
and UO_1124 (O_1124,N_24375,N_24774);
nor UO_1125 (O_1125,N_24741,N_24331);
nor UO_1126 (O_1126,N_24749,N_24266);
nor UO_1127 (O_1127,N_24911,N_24236);
xnor UO_1128 (O_1128,N_24954,N_24957);
or UO_1129 (O_1129,N_24749,N_24826);
xor UO_1130 (O_1130,N_24683,N_24927);
or UO_1131 (O_1131,N_24179,N_24499);
or UO_1132 (O_1132,N_24521,N_24142);
xor UO_1133 (O_1133,N_24984,N_24203);
nor UO_1134 (O_1134,N_24964,N_24850);
xor UO_1135 (O_1135,N_24931,N_24648);
nor UO_1136 (O_1136,N_24542,N_24426);
and UO_1137 (O_1137,N_24258,N_24055);
xnor UO_1138 (O_1138,N_24634,N_24874);
xor UO_1139 (O_1139,N_24660,N_24991);
or UO_1140 (O_1140,N_24238,N_24258);
nand UO_1141 (O_1141,N_24012,N_24815);
xor UO_1142 (O_1142,N_24476,N_24268);
nand UO_1143 (O_1143,N_24103,N_24935);
or UO_1144 (O_1144,N_24677,N_24848);
nand UO_1145 (O_1145,N_24761,N_24903);
nand UO_1146 (O_1146,N_24682,N_24966);
nor UO_1147 (O_1147,N_24502,N_24681);
nor UO_1148 (O_1148,N_24263,N_24014);
nor UO_1149 (O_1149,N_24886,N_24483);
nand UO_1150 (O_1150,N_24183,N_24557);
nand UO_1151 (O_1151,N_24128,N_24839);
nand UO_1152 (O_1152,N_24549,N_24930);
nand UO_1153 (O_1153,N_24429,N_24531);
or UO_1154 (O_1154,N_24529,N_24950);
nand UO_1155 (O_1155,N_24271,N_24870);
nand UO_1156 (O_1156,N_24673,N_24731);
nand UO_1157 (O_1157,N_24930,N_24630);
and UO_1158 (O_1158,N_24256,N_24934);
and UO_1159 (O_1159,N_24460,N_24031);
nor UO_1160 (O_1160,N_24199,N_24098);
nand UO_1161 (O_1161,N_24657,N_24279);
and UO_1162 (O_1162,N_24754,N_24912);
nand UO_1163 (O_1163,N_24086,N_24845);
nor UO_1164 (O_1164,N_24734,N_24195);
xnor UO_1165 (O_1165,N_24630,N_24980);
nand UO_1166 (O_1166,N_24488,N_24123);
nand UO_1167 (O_1167,N_24252,N_24881);
nor UO_1168 (O_1168,N_24020,N_24251);
nor UO_1169 (O_1169,N_24515,N_24160);
or UO_1170 (O_1170,N_24213,N_24197);
nand UO_1171 (O_1171,N_24488,N_24734);
xnor UO_1172 (O_1172,N_24168,N_24585);
nor UO_1173 (O_1173,N_24098,N_24964);
or UO_1174 (O_1174,N_24084,N_24538);
nand UO_1175 (O_1175,N_24245,N_24235);
nor UO_1176 (O_1176,N_24200,N_24460);
or UO_1177 (O_1177,N_24270,N_24784);
xnor UO_1178 (O_1178,N_24500,N_24515);
xor UO_1179 (O_1179,N_24904,N_24172);
or UO_1180 (O_1180,N_24010,N_24138);
or UO_1181 (O_1181,N_24736,N_24535);
and UO_1182 (O_1182,N_24830,N_24264);
and UO_1183 (O_1183,N_24348,N_24908);
or UO_1184 (O_1184,N_24282,N_24443);
nor UO_1185 (O_1185,N_24692,N_24063);
or UO_1186 (O_1186,N_24750,N_24810);
xnor UO_1187 (O_1187,N_24034,N_24790);
xor UO_1188 (O_1188,N_24510,N_24173);
and UO_1189 (O_1189,N_24569,N_24914);
or UO_1190 (O_1190,N_24083,N_24603);
or UO_1191 (O_1191,N_24185,N_24313);
or UO_1192 (O_1192,N_24280,N_24255);
and UO_1193 (O_1193,N_24550,N_24163);
nor UO_1194 (O_1194,N_24892,N_24730);
or UO_1195 (O_1195,N_24909,N_24744);
and UO_1196 (O_1196,N_24870,N_24303);
nor UO_1197 (O_1197,N_24549,N_24257);
or UO_1198 (O_1198,N_24978,N_24616);
or UO_1199 (O_1199,N_24960,N_24402);
and UO_1200 (O_1200,N_24448,N_24515);
nand UO_1201 (O_1201,N_24474,N_24641);
xnor UO_1202 (O_1202,N_24254,N_24992);
nor UO_1203 (O_1203,N_24011,N_24919);
or UO_1204 (O_1204,N_24668,N_24066);
xnor UO_1205 (O_1205,N_24517,N_24259);
xnor UO_1206 (O_1206,N_24253,N_24324);
nand UO_1207 (O_1207,N_24254,N_24700);
xor UO_1208 (O_1208,N_24454,N_24589);
and UO_1209 (O_1209,N_24369,N_24540);
xor UO_1210 (O_1210,N_24525,N_24906);
nor UO_1211 (O_1211,N_24931,N_24132);
nand UO_1212 (O_1212,N_24961,N_24511);
and UO_1213 (O_1213,N_24926,N_24774);
xnor UO_1214 (O_1214,N_24521,N_24212);
or UO_1215 (O_1215,N_24004,N_24336);
nor UO_1216 (O_1216,N_24130,N_24278);
xor UO_1217 (O_1217,N_24244,N_24994);
nand UO_1218 (O_1218,N_24827,N_24000);
and UO_1219 (O_1219,N_24095,N_24554);
xnor UO_1220 (O_1220,N_24793,N_24897);
nor UO_1221 (O_1221,N_24384,N_24152);
or UO_1222 (O_1222,N_24686,N_24406);
xnor UO_1223 (O_1223,N_24510,N_24982);
and UO_1224 (O_1224,N_24788,N_24397);
nor UO_1225 (O_1225,N_24152,N_24180);
nor UO_1226 (O_1226,N_24235,N_24199);
and UO_1227 (O_1227,N_24971,N_24458);
nor UO_1228 (O_1228,N_24980,N_24518);
and UO_1229 (O_1229,N_24466,N_24876);
xnor UO_1230 (O_1230,N_24000,N_24143);
nand UO_1231 (O_1231,N_24006,N_24443);
or UO_1232 (O_1232,N_24916,N_24945);
nor UO_1233 (O_1233,N_24527,N_24241);
xor UO_1234 (O_1234,N_24471,N_24988);
or UO_1235 (O_1235,N_24555,N_24260);
nor UO_1236 (O_1236,N_24315,N_24719);
nand UO_1237 (O_1237,N_24635,N_24524);
nor UO_1238 (O_1238,N_24823,N_24197);
nand UO_1239 (O_1239,N_24166,N_24144);
xor UO_1240 (O_1240,N_24756,N_24876);
nor UO_1241 (O_1241,N_24578,N_24790);
nor UO_1242 (O_1242,N_24324,N_24533);
or UO_1243 (O_1243,N_24523,N_24239);
nor UO_1244 (O_1244,N_24256,N_24921);
and UO_1245 (O_1245,N_24011,N_24597);
or UO_1246 (O_1246,N_24737,N_24118);
nand UO_1247 (O_1247,N_24769,N_24956);
nand UO_1248 (O_1248,N_24516,N_24608);
and UO_1249 (O_1249,N_24375,N_24370);
or UO_1250 (O_1250,N_24306,N_24320);
xor UO_1251 (O_1251,N_24955,N_24670);
and UO_1252 (O_1252,N_24174,N_24223);
nand UO_1253 (O_1253,N_24045,N_24023);
nor UO_1254 (O_1254,N_24959,N_24200);
and UO_1255 (O_1255,N_24949,N_24930);
xor UO_1256 (O_1256,N_24754,N_24447);
or UO_1257 (O_1257,N_24430,N_24680);
nor UO_1258 (O_1258,N_24724,N_24999);
or UO_1259 (O_1259,N_24600,N_24157);
nor UO_1260 (O_1260,N_24155,N_24075);
nor UO_1261 (O_1261,N_24781,N_24329);
or UO_1262 (O_1262,N_24534,N_24633);
nand UO_1263 (O_1263,N_24656,N_24242);
or UO_1264 (O_1264,N_24888,N_24249);
and UO_1265 (O_1265,N_24256,N_24954);
and UO_1266 (O_1266,N_24831,N_24672);
and UO_1267 (O_1267,N_24064,N_24257);
nand UO_1268 (O_1268,N_24076,N_24300);
xnor UO_1269 (O_1269,N_24985,N_24250);
and UO_1270 (O_1270,N_24349,N_24812);
xor UO_1271 (O_1271,N_24674,N_24404);
or UO_1272 (O_1272,N_24724,N_24238);
and UO_1273 (O_1273,N_24787,N_24309);
and UO_1274 (O_1274,N_24656,N_24598);
nand UO_1275 (O_1275,N_24667,N_24373);
nand UO_1276 (O_1276,N_24928,N_24285);
or UO_1277 (O_1277,N_24786,N_24661);
nand UO_1278 (O_1278,N_24793,N_24915);
xor UO_1279 (O_1279,N_24895,N_24329);
or UO_1280 (O_1280,N_24721,N_24708);
and UO_1281 (O_1281,N_24336,N_24124);
xnor UO_1282 (O_1282,N_24808,N_24324);
and UO_1283 (O_1283,N_24602,N_24648);
xnor UO_1284 (O_1284,N_24424,N_24497);
and UO_1285 (O_1285,N_24659,N_24281);
nand UO_1286 (O_1286,N_24609,N_24157);
nor UO_1287 (O_1287,N_24024,N_24832);
nand UO_1288 (O_1288,N_24455,N_24327);
nor UO_1289 (O_1289,N_24071,N_24406);
or UO_1290 (O_1290,N_24537,N_24361);
or UO_1291 (O_1291,N_24876,N_24663);
nand UO_1292 (O_1292,N_24376,N_24884);
and UO_1293 (O_1293,N_24258,N_24447);
or UO_1294 (O_1294,N_24763,N_24732);
xor UO_1295 (O_1295,N_24054,N_24621);
nand UO_1296 (O_1296,N_24584,N_24234);
nor UO_1297 (O_1297,N_24176,N_24312);
or UO_1298 (O_1298,N_24074,N_24202);
nand UO_1299 (O_1299,N_24525,N_24404);
or UO_1300 (O_1300,N_24014,N_24292);
xnor UO_1301 (O_1301,N_24426,N_24082);
nand UO_1302 (O_1302,N_24062,N_24103);
or UO_1303 (O_1303,N_24734,N_24018);
nor UO_1304 (O_1304,N_24942,N_24224);
and UO_1305 (O_1305,N_24434,N_24338);
nor UO_1306 (O_1306,N_24941,N_24114);
nor UO_1307 (O_1307,N_24052,N_24969);
or UO_1308 (O_1308,N_24804,N_24072);
or UO_1309 (O_1309,N_24864,N_24771);
nor UO_1310 (O_1310,N_24810,N_24157);
or UO_1311 (O_1311,N_24204,N_24281);
xor UO_1312 (O_1312,N_24612,N_24957);
xor UO_1313 (O_1313,N_24242,N_24088);
xor UO_1314 (O_1314,N_24894,N_24462);
nand UO_1315 (O_1315,N_24619,N_24150);
nor UO_1316 (O_1316,N_24294,N_24918);
xnor UO_1317 (O_1317,N_24723,N_24909);
and UO_1318 (O_1318,N_24327,N_24098);
nand UO_1319 (O_1319,N_24842,N_24887);
xnor UO_1320 (O_1320,N_24728,N_24563);
and UO_1321 (O_1321,N_24790,N_24252);
xnor UO_1322 (O_1322,N_24560,N_24879);
xor UO_1323 (O_1323,N_24924,N_24468);
xnor UO_1324 (O_1324,N_24100,N_24646);
and UO_1325 (O_1325,N_24779,N_24530);
or UO_1326 (O_1326,N_24257,N_24005);
nor UO_1327 (O_1327,N_24399,N_24788);
xor UO_1328 (O_1328,N_24271,N_24592);
or UO_1329 (O_1329,N_24419,N_24852);
nand UO_1330 (O_1330,N_24273,N_24381);
or UO_1331 (O_1331,N_24971,N_24815);
and UO_1332 (O_1332,N_24138,N_24881);
and UO_1333 (O_1333,N_24187,N_24330);
and UO_1334 (O_1334,N_24041,N_24859);
or UO_1335 (O_1335,N_24391,N_24003);
nand UO_1336 (O_1336,N_24468,N_24375);
nand UO_1337 (O_1337,N_24801,N_24804);
and UO_1338 (O_1338,N_24487,N_24931);
or UO_1339 (O_1339,N_24337,N_24182);
xnor UO_1340 (O_1340,N_24783,N_24194);
or UO_1341 (O_1341,N_24448,N_24107);
and UO_1342 (O_1342,N_24639,N_24433);
nor UO_1343 (O_1343,N_24885,N_24767);
or UO_1344 (O_1344,N_24657,N_24027);
and UO_1345 (O_1345,N_24564,N_24720);
xnor UO_1346 (O_1346,N_24747,N_24053);
or UO_1347 (O_1347,N_24436,N_24287);
or UO_1348 (O_1348,N_24086,N_24054);
and UO_1349 (O_1349,N_24134,N_24486);
or UO_1350 (O_1350,N_24467,N_24227);
xor UO_1351 (O_1351,N_24416,N_24426);
nor UO_1352 (O_1352,N_24360,N_24389);
and UO_1353 (O_1353,N_24593,N_24507);
xnor UO_1354 (O_1354,N_24590,N_24766);
and UO_1355 (O_1355,N_24689,N_24926);
and UO_1356 (O_1356,N_24230,N_24321);
and UO_1357 (O_1357,N_24874,N_24739);
or UO_1358 (O_1358,N_24691,N_24004);
nor UO_1359 (O_1359,N_24975,N_24589);
or UO_1360 (O_1360,N_24670,N_24215);
or UO_1361 (O_1361,N_24546,N_24590);
or UO_1362 (O_1362,N_24306,N_24678);
and UO_1363 (O_1363,N_24147,N_24962);
nand UO_1364 (O_1364,N_24557,N_24085);
or UO_1365 (O_1365,N_24783,N_24118);
or UO_1366 (O_1366,N_24174,N_24968);
xnor UO_1367 (O_1367,N_24950,N_24414);
or UO_1368 (O_1368,N_24750,N_24952);
nand UO_1369 (O_1369,N_24605,N_24564);
nand UO_1370 (O_1370,N_24062,N_24501);
or UO_1371 (O_1371,N_24923,N_24835);
and UO_1372 (O_1372,N_24580,N_24870);
or UO_1373 (O_1373,N_24403,N_24496);
xor UO_1374 (O_1374,N_24408,N_24456);
and UO_1375 (O_1375,N_24894,N_24026);
or UO_1376 (O_1376,N_24902,N_24423);
or UO_1377 (O_1377,N_24031,N_24540);
nor UO_1378 (O_1378,N_24651,N_24551);
nand UO_1379 (O_1379,N_24507,N_24827);
or UO_1380 (O_1380,N_24964,N_24837);
and UO_1381 (O_1381,N_24055,N_24064);
nand UO_1382 (O_1382,N_24359,N_24424);
and UO_1383 (O_1383,N_24289,N_24669);
or UO_1384 (O_1384,N_24076,N_24154);
and UO_1385 (O_1385,N_24978,N_24005);
nor UO_1386 (O_1386,N_24613,N_24418);
or UO_1387 (O_1387,N_24814,N_24865);
and UO_1388 (O_1388,N_24171,N_24580);
and UO_1389 (O_1389,N_24213,N_24214);
xnor UO_1390 (O_1390,N_24594,N_24016);
and UO_1391 (O_1391,N_24713,N_24241);
and UO_1392 (O_1392,N_24800,N_24226);
or UO_1393 (O_1393,N_24020,N_24385);
nand UO_1394 (O_1394,N_24362,N_24151);
nor UO_1395 (O_1395,N_24884,N_24880);
or UO_1396 (O_1396,N_24375,N_24957);
xnor UO_1397 (O_1397,N_24246,N_24907);
xor UO_1398 (O_1398,N_24587,N_24485);
xor UO_1399 (O_1399,N_24731,N_24105);
xor UO_1400 (O_1400,N_24441,N_24672);
xnor UO_1401 (O_1401,N_24859,N_24717);
nand UO_1402 (O_1402,N_24779,N_24101);
nor UO_1403 (O_1403,N_24148,N_24956);
nand UO_1404 (O_1404,N_24727,N_24880);
nor UO_1405 (O_1405,N_24269,N_24874);
xor UO_1406 (O_1406,N_24715,N_24048);
xnor UO_1407 (O_1407,N_24921,N_24067);
nor UO_1408 (O_1408,N_24227,N_24976);
or UO_1409 (O_1409,N_24010,N_24722);
xnor UO_1410 (O_1410,N_24648,N_24548);
and UO_1411 (O_1411,N_24490,N_24574);
nor UO_1412 (O_1412,N_24350,N_24142);
nand UO_1413 (O_1413,N_24900,N_24317);
nor UO_1414 (O_1414,N_24557,N_24726);
and UO_1415 (O_1415,N_24917,N_24466);
or UO_1416 (O_1416,N_24281,N_24554);
xor UO_1417 (O_1417,N_24055,N_24710);
or UO_1418 (O_1418,N_24680,N_24196);
nor UO_1419 (O_1419,N_24045,N_24173);
nor UO_1420 (O_1420,N_24512,N_24073);
and UO_1421 (O_1421,N_24768,N_24623);
or UO_1422 (O_1422,N_24867,N_24167);
nor UO_1423 (O_1423,N_24068,N_24001);
nor UO_1424 (O_1424,N_24504,N_24092);
nor UO_1425 (O_1425,N_24448,N_24149);
nand UO_1426 (O_1426,N_24075,N_24456);
nand UO_1427 (O_1427,N_24337,N_24666);
nand UO_1428 (O_1428,N_24850,N_24559);
nor UO_1429 (O_1429,N_24827,N_24163);
xnor UO_1430 (O_1430,N_24228,N_24142);
nand UO_1431 (O_1431,N_24331,N_24818);
xnor UO_1432 (O_1432,N_24372,N_24493);
xnor UO_1433 (O_1433,N_24136,N_24207);
and UO_1434 (O_1434,N_24766,N_24510);
nor UO_1435 (O_1435,N_24530,N_24408);
nand UO_1436 (O_1436,N_24680,N_24149);
nand UO_1437 (O_1437,N_24697,N_24287);
and UO_1438 (O_1438,N_24408,N_24701);
nor UO_1439 (O_1439,N_24694,N_24259);
xor UO_1440 (O_1440,N_24079,N_24503);
xor UO_1441 (O_1441,N_24357,N_24040);
nor UO_1442 (O_1442,N_24692,N_24081);
and UO_1443 (O_1443,N_24468,N_24421);
xnor UO_1444 (O_1444,N_24521,N_24256);
or UO_1445 (O_1445,N_24000,N_24030);
nor UO_1446 (O_1446,N_24000,N_24757);
and UO_1447 (O_1447,N_24903,N_24999);
nor UO_1448 (O_1448,N_24762,N_24497);
nor UO_1449 (O_1449,N_24496,N_24001);
and UO_1450 (O_1450,N_24175,N_24662);
or UO_1451 (O_1451,N_24308,N_24164);
or UO_1452 (O_1452,N_24772,N_24569);
or UO_1453 (O_1453,N_24775,N_24128);
and UO_1454 (O_1454,N_24574,N_24791);
or UO_1455 (O_1455,N_24791,N_24154);
or UO_1456 (O_1456,N_24994,N_24454);
xor UO_1457 (O_1457,N_24473,N_24356);
and UO_1458 (O_1458,N_24448,N_24236);
nand UO_1459 (O_1459,N_24829,N_24287);
and UO_1460 (O_1460,N_24699,N_24886);
xnor UO_1461 (O_1461,N_24213,N_24151);
nor UO_1462 (O_1462,N_24585,N_24399);
and UO_1463 (O_1463,N_24989,N_24919);
or UO_1464 (O_1464,N_24995,N_24742);
and UO_1465 (O_1465,N_24489,N_24954);
and UO_1466 (O_1466,N_24797,N_24472);
and UO_1467 (O_1467,N_24569,N_24337);
nand UO_1468 (O_1468,N_24028,N_24543);
nor UO_1469 (O_1469,N_24605,N_24253);
xnor UO_1470 (O_1470,N_24548,N_24465);
nand UO_1471 (O_1471,N_24196,N_24266);
nand UO_1472 (O_1472,N_24098,N_24160);
or UO_1473 (O_1473,N_24975,N_24632);
or UO_1474 (O_1474,N_24864,N_24741);
xor UO_1475 (O_1475,N_24383,N_24215);
nand UO_1476 (O_1476,N_24248,N_24042);
nor UO_1477 (O_1477,N_24427,N_24049);
xor UO_1478 (O_1478,N_24993,N_24511);
nand UO_1479 (O_1479,N_24571,N_24648);
nand UO_1480 (O_1480,N_24513,N_24588);
nor UO_1481 (O_1481,N_24462,N_24796);
xor UO_1482 (O_1482,N_24584,N_24460);
xor UO_1483 (O_1483,N_24791,N_24783);
nor UO_1484 (O_1484,N_24334,N_24584);
and UO_1485 (O_1485,N_24950,N_24456);
nor UO_1486 (O_1486,N_24930,N_24775);
nand UO_1487 (O_1487,N_24127,N_24051);
or UO_1488 (O_1488,N_24951,N_24154);
xor UO_1489 (O_1489,N_24193,N_24822);
or UO_1490 (O_1490,N_24727,N_24860);
or UO_1491 (O_1491,N_24671,N_24481);
and UO_1492 (O_1492,N_24808,N_24314);
nor UO_1493 (O_1493,N_24058,N_24805);
xnor UO_1494 (O_1494,N_24743,N_24905);
nor UO_1495 (O_1495,N_24447,N_24199);
nor UO_1496 (O_1496,N_24274,N_24883);
or UO_1497 (O_1497,N_24279,N_24126);
nor UO_1498 (O_1498,N_24481,N_24085);
or UO_1499 (O_1499,N_24600,N_24813);
nand UO_1500 (O_1500,N_24118,N_24745);
and UO_1501 (O_1501,N_24394,N_24693);
or UO_1502 (O_1502,N_24353,N_24124);
nor UO_1503 (O_1503,N_24152,N_24050);
and UO_1504 (O_1504,N_24180,N_24005);
or UO_1505 (O_1505,N_24398,N_24210);
xnor UO_1506 (O_1506,N_24571,N_24070);
xor UO_1507 (O_1507,N_24935,N_24820);
xnor UO_1508 (O_1508,N_24158,N_24605);
nor UO_1509 (O_1509,N_24560,N_24266);
xor UO_1510 (O_1510,N_24128,N_24197);
and UO_1511 (O_1511,N_24005,N_24642);
and UO_1512 (O_1512,N_24359,N_24498);
and UO_1513 (O_1513,N_24805,N_24786);
or UO_1514 (O_1514,N_24859,N_24575);
nor UO_1515 (O_1515,N_24085,N_24570);
and UO_1516 (O_1516,N_24220,N_24010);
or UO_1517 (O_1517,N_24626,N_24572);
xor UO_1518 (O_1518,N_24212,N_24311);
and UO_1519 (O_1519,N_24363,N_24153);
or UO_1520 (O_1520,N_24427,N_24380);
xnor UO_1521 (O_1521,N_24538,N_24821);
or UO_1522 (O_1522,N_24271,N_24266);
nor UO_1523 (O_1523,N_24103,N_24981);
and UO_1524 (O_1524,N_24630,N_24803);
and UO_1525 (O_1525,N_24532,N_24802);
nor UO_1526 (O_1526,N_24344,N_24514);
and UO_1527 (O_1527,N_24900,N_24886);
nand UO_1528 (O_1528,N_24734,N_24257);
or UO_1529 (O_1529,N_24682,N_24170);
or UO_1530 (O_1530,N_24595,N_24035);
and UO_1531 (O_1531,N_24955,N_24349);
or UO_1532 (O_1532,N_24129,N_24886);
or UO_1533 (O_1533,N_24719,N_24865);
or UO_1534 (O_1534,N_24110,N_24686);
xor UO_1535 (O_1535,N_24740,N_24599);
or UO_1536 (O_1536,N_24240,N_24108);
xnor UO_1537 (O_1537,N_24517,N_24169);
nand UO_1538 (O_1538,N_24441,N_24479);
nand UO_1539 (O_1539,N_24402,N_24200);
xor UO_1540 (O_1540,N_24262,N_24229);
xor UO_1541 (O_1541,N_24085,N_24161);
nand UO_1542 (O_1542,N_24058,N_24214);
xor UO_1543 (O_1543,N_24338,N_24030);
nand UO_1544 (O_1544,N_24289,N_24776);
and UO_1545 (O_1545,N_24750,N_24543);
and UO_1546 (O_1546,N_24128,N_24829);
and UO_1547 (O_1547,N_24301,N_24632);
or UO_1548 (O_1548,N_24070,N_24959);
and UO_1549 (O_1549,N_24220,N_24239);
xnor UO_1550 (O_1550,N_24413,N_24806);
and UO_1551 (O_1551,N_24267,N_24753);
nand UO_1552 (O_1552,N_24833,N_24967);
nand UO_1553 (O_1553,N_24938,N_24884);
xor UO_1554 (O_1554,N_24018,N_24559);
nor UO_1555 (O_1555,N_24734,N_24303);
nor UO_1556 (O_1556,N_24488,N_24072);
or UO_1557 (O_1557,N_24669,N_24047);
xor UO_1558 (O_1558,N_24823,N_24712);
and UO_1559 (O_1559,N_24282,N_24540);
nand UO_1560 (O_1560,N_24680,N_24617);
or UO_1561 (O_1561,N_24281,N_24966);
nor UO_1562 (O_1562,N_24637,N_24230);
or UO_1563 (O_1563,N_24239,N_24970);
or UO_1564 (O_1564,N_24457,N_24696);
and UO_1565 (O_1565,N_24564,N_24072);
or UO_1566 (O_1566,N_24115,N_24941);
or UO_1567 (O_1567,N_24665,N_24788);
xnor UO_1568 (O_1568,N_24267,N_24457);
xnor UO_1569 (O_1569,N_24350,N_24412);
or UO_1570 (O_1570,N_24683,N_24071);
and UO_1571 (O_1571,N_24796,N_24989);
nor UO_1572 (O_1572,N_24520,N_24529);
nor UO_1573 (O_1573,N_24423,N_24922);
or UO_1574 (O_1574,N_24143,N_24472);
or UO_1575 (O_1575,N_24273,N_24243);
nor UO_1576 (O_1576,N_24612,N_24069);
xnor UO_1577 (O_1577,N_24317,N_24193);
nand UO_1578 (O_1578,N_24624,N_24648);
and UO_1579 (O_1579,N_24166,N_24510);
nor UO_1580 (O_1580,N_24657,N_24767);
nor UO_1581 (O_1581,N_24201,N_24886);
xnor UO_1582 (O_1582,N_24621,N_24190);
nand UO_1583 (O_1583,N_24481,N_24306);
and UO_1584 (O_1584,N_24219,N_24370);
or UO_1585 (O_1585,N_24342,N_24994);
nand UO_1586 (O_1586,N_24672,N_24187);
or UO_1587 (O_1587,N_24204,N_24291);
xnor UO_1588 (O_1588,N_24772,N_24462);
and UO_1589 (O_1589,N_24339,N_24631);
or UO_1590 (O_1590,N_24445,N_24340);
xor UO_1591 (O_1591,N_24887,N_24501);
or UO_1592 (O_1592,N_24680,N_24611);
nor UO_1593 (O_1593,N_24465,N_24763);
nand UO_1594 (O_1594,N_24760,N_24131);
and UO_1595 (O_1595,N_24409,N_24835);
nand UO_1596 (O_1596,N_24492,N_24130);
xor UO_1597 (O_1597,N_24973,N_24336);
and UO_1598 (O_1598,N_24540,N_24351);
nand UO_1599 (O_1599,N_24299,N_24492);
and UO_1600 (O_1600,N_24169,N_24430);
or UO_1601 (O_1601,N_24186,N_24188);
nand UO_1602 (O_1602,N_24703,N_24709);
xor UO_1603 (O_1603,N_24640,N_24106);
xor UO_1604 (O_1604,N_24475,N_24408);
and UO_1605 (O_1605,N_24154,N_24637);
nor UO_1606 (O_1606,N_24807,N_24020);
xor UO_1607 (O_1607,N_24029,N_24456);
xnor UO_1608 (O_1608,N_24856,N_24547);
nor UO_1609 (O_1609,N_24023,N_24948);
xnor UO_1610 (O_1610,N_24996,N_24437);
or UO_1611 (O_1611,N_24124,N_24118);
xnor UO_1612 (O_1612,N_24927,N_24156);
or UO_1613 (O_1613,N_24612,N_24706);
or UO_1614 (O_1614,N_24108,N_24556);
or UO_1615 (O_1615,N_24979,N_24382);
and UO_1616 (O_1616,N_24484,N_24566);
nor UO_1617 (O_1617,N_24261,N_24507);
nor UO_1618 (O_1618,N_24161,N_24310);
nand UO_1619 (O_1619,N_24022,N_24442);
or UO_1620 (O_1620,N_24579,N_24229);
and UO_1621 (O_1621,N_24844,N_24448);
nand UO_1622 (O_1622,N_24294,N_24579);
nor UO_1623 (O_1623,N_24182,N_24172);
xnor UO_1624 (O_1624,N_24979,N_24547);
xnor UO_1625 (O_1625,N_24755,N_24476);
xor UO_1626 (O_1626,N_24263,N_24260);
and UO_1627 (O_1627,N_24280,N_24824);
and UO_1628 (O_1628,N_24111,N_24524);
or UO_1629 (O_1629,N_24099,N_24634);
and UO_1630 (O_1630,N_24698,N_24138);
nand UO_1631 (O_1631,N_24355,N_24964);
nand UO_1632 (O_1632,N_24214,N_24412);
or UO_1633 (O_1633,N_24735,N_24628);
nor UO_1634 (O_1634,N_24682,N_24744);
and UO_1635 (O_1635,N_24666,N_24237);
xor UO_1636 (O_1636,N_24030,N_24590);
nand UO_1637 (O_1637,N_24034,N_24512);
and UO_1638 (O_1638,N_24163,N_24222);
or UO_1639 (O_1639,N_24936,N_24284);
or UO_1640 (O_1640,N_24468,N_24635);
or UO_1641 (O_1641,N_24732,N_24656);
nand UO_1642 (O_1642,N_24309,N_24445);
and UO_1643 (O_1643,N_24356,N_24267);
and UO_1644 (O_1644,N_24071,N_24638);
and UO_1645 (O_1645,N_24537,N_24768);
or UO_1646 (O_1646,N_24663,N_24868);
xnor UO_1647 (O_1647,N_24082,N_24570);
xnor UO_1648 (O_1648,N_24704,N_24407);
and UO_1649 (O_1649,N_24163,N_24739);
nor UO_1650 (O_1650,N_24571,N_24039);
nor UO_1651 (O_1651,N_24051,N_24157);
nor UO_1652 (O_1652,N_24695,N_24543);
or UO_1653 (O_1653,N_24035,N_24770);
nor UO_1654 (O_1654,N_24183,N_24287);
xnor UO_1655 (O_1655,N_24133,N_24246);
nand UO_1656 (O_1656,N_24340,N_24483);
and UO_1657 (O_1657,N_24687,N_24217);
xnor UO_1658 (O_1658,N_24732,N_24851);
or UO_1659 (O_1659,N_24363,N_24041);
nand UO_1660 (O_1660,N_24162,N_24397);
xor UO_1661 (O_1661,N_24998,N_24518);
xnor UO_1662 (O_1662,N_24034,N_24975);
xor UO_1663 (O_1663,N_24984,N_24438);
or UO_1664 (O_1664,N_24559,N_24088);
nand UO_1665 (O_1665,N_24737,N_24721);
nor UO_1666 (O_1666,N_24958,N_24818);
xor UO_1667 (O_1667,N_24032,N_24905);
xnor UO_1668 (O_1668,N_24668,N_24162);
nand UO_1669 (O_1669,N_24008,N_24620);
or UO_1670 (O_1670,N_24533,N_24583);
xor UO_1671 (O_1671,N_24347,N_24204);
xnor UO_1672 (O_1672,N_24535,N_24181);
nor UO_1673 (O_1673,N_24454,N_24133);
and UO_1674 (O_1674,N_24295,N_24662);
nor UO_1675 (O_1675,N_24133,N_24717);
and UO_1676 (O_1676,N_24974,N_24780);
or UO_1677 (O_1677,N_24252,N_24559);
or UO_1678 (O_1678,N_24651,N_24478);
nor UO_1679 (O_1679,N_24412,N_24735);
xnor UO_1680 (O_1680,N_24009,N_24995);
and UO_1681 (O_1681,N_24064,N_24047);
nand UO_1682 (O_1682,N_24598,N_24073);
xnor UO_1683 (O_1683,N_24049,N_24090);
xor UO_1684 (O_1684,N_24561,N_24279);
and UO_1685 (O_1685,N_24874,N_24864);
or UO_1686 (O_1686,N_24531,N_24087);
and UO_1687 (O_1687,N_24461,N_24179);
xnor UO_1688 (O_1688,N_24122,N_24065);
and UO_1689 (O_1689,N_24328,N_24719);
xnor UO_1690 (O_1690,N_24149,N_24167);
nand UO_1691 (O_1691,N_24185,N_24774);
nand UO_1692 (O_1692,N_24361,N_24612);
nor UO_1693 (O_1693,N_24809,N_24495);
xnor UO_1694 (O_1694,N_24695,N_24675);
nor UO_1695 (O_1695,N_24717,N_24576);
nor UO_1696 (O_1696,N_24241,N_24451);
nand UO_1697 (O_1697,N_24053,N_24038);
nor UO_1698 (O_1698,N_24073,N_24774);
and UO_1699 (O_1699,N_24267,N_24342);
nand UO_1700 (O_1700,N_24115,N_24714);
xor UO_1701 (O_1701,N_24998,N_24428);
nor UO_1702 (O_1702,N_24162,N_24471);
xnor UO_1703 (O_1703,N_24794,N_24056);
and UO_1704 (O_1704,N_24241,N_24684);
xor UO_1705 (O_1705,N_24998,N_24772);
nand UO_1706 (O_1706,N_24334,N_24983);
nand UO_1707 (O_1707,N_24261,N_24152);
and UO_1708 (O_1708,N_24925,N_24582);
xor UO_1709 (O_1709,N_24508,N_24740);
or UO_1710 (O_1710,N_24380,N_24987);
or UO_1711 (O_1711,N_24011,N_24662);
and UO_1712 (O_1712,N_24517,N_24466);
xor UO_1713 (O_1713,N_24374,N_24983);
xnor UO_1714 (O_1714,N_24460,N_24594);
nand UO_1715 (O_1715,N_24094,N_24109);
nor UO_1716 (O_1716,N_24896,N_24573);
and UO_1717 (O_1717,N_24765,N_24037);
xor UO_1718 (O_1718,N_24221,N_24523);
xnor UO_1719 (O_1719,N_24005,N_24714);
or UO_1720 (O_1720,N_24729,N_24417);
or UO_1721 (O_1721,N_24412,N_24095);
nand UO_1722 (O_1722,N_24918,N_24391);
and UO_1723 (O_1723,N_24607,N_24148);
and UO_1724 (O_1724,N_24838,N_24534);
nand UO_1725 (O_1725,N_24459,N_24988);
or UO_1726 (O_1726,N_24288,N_24116);
or UO_1727 (O_1727,N_24085,N_24309);
nand UO_1728 (O_1728,N_24696,N_24521);
xor UO_1729 (O_1729,N_24449,N_24695);
nand UO_1730 (O_1730,N_24863,N_24252);
nand UO_1731 (O_1731,N_24530,N_24572);
and UO_1732 (O_1732,N_24697,N_24897);
nand UO_1733 (O_1733,N_24133,N_24332);
or UO_1734 (O_1734,N_24962,N_24219);
or UO_1735 (O_1735,N_24835,N_24598);
xnor UO_1736 (O_1736,N_24681,N_24616);
nand UO_1737 (O_1737,N_24733,N_24547);
nand UO_1738 (O_1738,N_24427,N_24909);
and UO_1739 (O_1739,N_24975,N_24068);
or UO_1740 (O_1740,N_24636,N_24952);
or UO_1741 (O_1741,N_24086,N_24683);
xnor UO_1742 (O_1742,N_24295,N_24643);
xor UO_1743 (O_1743,N_24933,N_24222);
or UO_1744 (O_1744,N_24158,N_24284);
nand UO_1745 (O_1745,N_24190,N_24270);
nor UO_1746 (O_1746,N_24592,N_24451);
nor UO_1747 (O_1747,N_24492,N_24416);
nor UO_1748 (O_1748,N_24931,N_24074);
and UO_1749 (O_1749,N_24734,N_24494);
nor UO_1750 (O_1750,N_24822,N_24303);
or UO_1751 (O_1751,N_24764,N_24383);
xor UO_1752 (O_1752,N_24998,N_24162);
nor UO_1753 (O_1753,N_24805,N_24215);
xor UO_1754 (O_1754,N_24111,N_24081);
xor UO_1755 (O_1755,N_24802,N_24703);
xor UO_1756 (O_1756,N_24549,N_24238);
nor UO_1757 (O_1757,N_24328,N_24859);
and UO_1758 (O_1758,N_24171,N_24659);
and UO_1759 (O_1759,N_24141,N_24247);
nor UO_1760 (O_1760,N_24734,N_24562);
nand UO_1761 (O_1761,N_24468,N_24980);
xor UO_1762 (O_1762,N_24109,N_24445);
nand UO_1763 (O_1763,N_24939,N_24294);
and UO_1764 (O_1764,N_24837,N_24636);
nand UO_1765 (O_1765,N_24852,N_24954);
nand UO_1766 (O_1766,N_24140,N_24843);
nand UO_1767 (O_1767,N_24034,N_24015);
xnor UO_1768 (O_1768,N_24589,N_24126);
nor UO_1769 (O_1769,N_24151,N_24477);
nor UO_1770 (O_1770,N_24275,N_24854);
nor UO_1771 (O_1771,N_24955,N_24508);
or UO_1772 (O_1772,N_24916,N_24694);
nor UO_1773 (O_1773,N_24562,N_24816);
or UO_1774 (O_1774,N_24825,N_24053);
or UO_1775 (O_1775,N_24323,N_24146);
and UO_1776 (O_1776,N_24879,N_24921);
or UO_1777 (O_1777,N_24115,N_24416);
or UO_1778 (O_1778,N_24396,N_24071);
xor UO_1779 (O_1779,N_24992,N_24366);
xor UO_1780 (O_1780,N_24965,N_24980);
nor UO_1781 (O_1781,N_24190,N_24126);
or UO_1782 (O_1782,N_24078,N_24344);
xnor UO_1783 (O_1783,N_24101,N_24061);
nor UO_1784 (O_1784,N_24783,N_24120);
nor UO_1785 (O_1785,N_24597,N_24886);
nor UO_1786 (O_1786,N_24198,N_24386);
xnor UO_1787 (O_1787,N_24918,N_24485);
nand UO_1788 (O_1788,N_24523,N_24992);
or UO_1789 (O_1789,N_24841,N_24476);
xnor UO_1790 (O_1790,N_24515,N_24152);
nor UO_1791 (O_1791,N_24759,N_24915);
and UO_1792 (O_1792,N_24335,N_24499);
nand UO_1793 (O_1793,N_24489,N_24696);
nand UO_1794 (O_1794,N_24049,N_24980);
nor UO_1795 (O_1795,N_24022,N_24819);
nor UO_1796 (O_1796,N_24170,N_24759);
and UO_1797 (O_1797,N_24349,N_24287);
and UO_1798 (O_1798,N_24688,N_24741);
xnor UO_1799 (O_1799,N_24785,N_24284);
nand UO_1800 (O_1800,N_24351,N_24332);
nand UO_1801 (O_1801,N_24977,N_24826);
xnor UO_1802 (O_1802,N_24220,N_24850);
xor UO_1803 (O_1803,N_24779,N_24595);
and UO_1804 (O_1804,N_24986,N_24569);
and UO_1805 (O_1805,N_24142,N_24636);
nor UO_1806 (O_1806,N_24493,N_24275);
nor UO_1807 (O_1807,N_24635,N_24397);
xor UO_1808 (O_1808,N_24840,N_24028);
or UO_1809 (O_1809,N_24873,N_24372);
or UO_1810 (O_1810,N_24975,N_24646);
xor UO_1811 (O_1811,N_24977,N_24337);
nand UO_1812 (O_1812,N_24235,N_24360);
and UO_1813 (O_1813,N_24496,N_24749);
xor UO_1814 (O_1814,N_24338,N_24867);
nor UO_1815 (O_1815,N_24896,N_24695);
xor UO_1816 (O_1816,N_24430,N_24912);
and UO_1817 (O_1817,N_24211,N_24725);
xnor UO_1818 (O_1818,N_24036,N_24153);
nor UO_1819 (O_1819,N_24396,N_24422);
nor UO_1820 (O_1820,N_24899,N_24601);
nor UO_1821 (O_1821,N_24471,N_24460);
nor UO_1822 (O_1822,N_24258,N_24230);
xor UO_1823 (O_1823,N_24897,N_24245);
and UO_1824 (O_1824,N_24158,N_24627);
and UO_1825 (O_1825,N_24230,N_24342);
nor UO_1826 (O_1826,N_24475,N_24298);
and UO_1827 (O_1827,N_24865,N_24647);
nor UO_1828 (O_1828,N_24153,N_24147);
xor UO_1829 (O_1829,N_24458,N_24337);
nand UO_1830 (O_1830,N_24845,N_24569);
and UO_1831 (O_1831,N_24573,N_24420);
xnor UO_1832 (O_1832,N_24703,N_24899);
nor UO_1833 (O_1833,N_24284,N_24555);
or UO_1834 (O_1834,N_24722,N_24600);
nor UO_1835 (O_1835,N_24200,N_24958);
nand UO_1836 (O_1836,N_24241,N_24870);
nor UO_1837 (O_1837,N_24227,N_24023);
nand UO_1838 (O_1838,N_24526,N_24727);
xor UO_1839 (O_1839,N_24772,N_24303);
or UO_1840 (O_1840,N_24730,N_24967);
nor UO_1841 (O_1841,N_24579,N_24014);
and UO_1842 (O_1842,N_24638,N_24166);
or UO_1843 (O_1843,N_24696,N_24620);
or UO_1844 (O_1844,N_24324,N_24161);
nand UO_1845 (O_1845,N_24579,N_24813);
xnor UO_1846 (O_1846,N_24295,N_24439);
or UO_1847 (O_1847,N_24801,N_24143);
or UO_1848 (O_1848,N_24848,N_24930);
or UO_1849 (O_1849,N_24726,N_24268);
nor UO_1850 (O_1850,N_24776,N_24789);
or UO_1851 (O_1851,N_24052,N_24437);
and UO_1852 (O_1852,N_24351,N_24690);
nor UO_1853 (O_1853,N_24281,N_24056);
nand UO_1854 (O_1854,N_24650,N_24799);
nand UO_1855 (O_1855,N_24758,N_24708);
or UO_1856 (O_1856,N_24743,N_24897);
and UO_1857 (O_1857,N_24693,N_24124);
xor UO_1858 (O_1858,N_24821,N_24915);
xor UO_1859 (O_1859,N_24952,N_24486);
nor UO_1860 (O_1860,N_24852,N_24102);
or UO_1861 (O_1861,N_24694,N_24151);
or UO_1862 (O_1862,N_24216,N_24311);
or UO_1863 (O_1863,N_24008,N_24762);
nor UO_1864 (O_1864,N_24411,N_24748);
nor UO_1865 (O_1865,N_24729,N_24149);
or UO_1866 (O_1866,N_24382,N_24242);
and UO_1867 (O_1867,N_24732,N_24208);
or UO_1868 (O_1868,N_24594,N_24048);
nand UO_1869 (O_1869,N_24987,N_24558);
nor UO_1870 (O_1870,N_24549,N_24025);
xnor UO_1871 (O_1871,N_24599,N_24277);
xor UO_1872 (O_1872,N_24156,N_24612);
nor UO_1873 (O_1873,N_24414,N_24987);
and UO_1874 (O_1874,N_24095,N_24139);
nand UO_1875 (O_1875,N_24707,N_24096);
xor UO_1876 (O_1876,N_24600,N_24120);
xnor UO_1877 (O_1877,N_24844,N_24581);
xor UO_1878 (O_1878,N_24148,N_24582);
or UO_1879 (O_1879,N_24621,N_24545);
and UO_1880 (O_1880,N_24311,N_24871);
or UO_1881 (O_1881,N_24772,N_24892);
and UO_1882 (O_1882,N_24175,N_24000);
or UO_1883 (O_1883,N_24919,N_24627);
or UO_1884 (O_1884,N_24610,N_24436);
and UO_1885 (O_1885,N_24595,N_24290);
nor UO_1886 (O_1886,N_24149,N_24578);
xor UO_1887 (O_1887,N_24766,N_24302);
and UO_1888 (O_1888,N_24630,N_24606);
xor UO_1889 (O_1889,N_24929,N_24901);
and UO_1890 (O_1890,N_24696,N_24219);
nand UO_1891 (O_1891,N_24672,N_24394);
nand UO_1892 (O_1892,N_24405,N_24236);
nand UO_1893 (O_1893,N_24331,N_24565);
and UO_1894 (O_1894,N_24929,N_24473);
nand UO_1895 (O_1895,N_24017,N_24015);
nor UO_1896 (O_1896,N_24850,N_24272);
and UO_1897 (O_1897,N_24245,N_24338);
nand UO_1898 (O_1898,N_24081,N_24204);
nor UO_1899 (O_1899,N_24502,N_24212);
nand UO_1900 (O_1900,N_24951,N_24611);
nand UO_1901 (O_1901,N_24221,N_24395);
or UO_1902 (O_1902,N_24100,N_24761);
and UO_1903 (O_1903,N_24131,N_24243);
or UO_1904 (O_1904,N_24719,N_24062);
nor UO_1905 (O_1905,N_24967,N_24933);
or UO_1906 (O_1906,N_24056,N_24062);
nand UO_1907 (O_1907,N_24705,N_24183);
or UO_1908 (O_1908,N_24687,N_24477);
nand UO_1909 (O_1909,N_24718,N_24374);
or UO_1910 (O_1910,N_24509,N_24626);
or UO_1911 (O_1911,N_24022,N_24994);
or UO_1912 (O_1912,N_24623,N_24294);
nand UO_1913 (O_1913,N_24218,N_24844);
or UO_1914 (O_1914,N_24957,N_24813);
or UO_1915 (O_1915,N_24946,N_24169);
xnor UO_1916 (O_1916,N_24089,N_24355);
or UO_1917 (O_1917,N_24707,N_24184);
and UO_1918 (O_1918,N_24174,N_24169);
and UO_1919 (O_1919,N_24080,N_24381);
nor UO_1920 (O_1920,N_24635,N_24663);
nor UO_1921 (O_1921,N_24515,N_24086);
nand UO_1922 (O_1922,N_24061,N_24166);
and UO_1923 (O_1923,N_24289,N_24065);
and UO_1924 (O_1924,N_24397,N_24104);
nor UO_1925 (O_1925,N_24196,N_24476);
and UO_1926 (O_1926,N_24950,N_24178);
nand UO_1927 (O_1927,N_24515,N_24394);
xnor UO_1928 (O_1928,N_24336,N_24412);
or UO_1929 (O_1929,N_24171,N_24616);
or UO_1930 (O_1930,N_24718,N_24067);
and UO_1931 (O_1931,N_24012,N_24166);
nor UO_1932 (O_1932,N_24666,N_24677);
and UO_1933 (O_1933,N_24895,N_24775);
xnor UO_1934 (O_1934,N_24231,N_24723);
or UO_1935 (O_1935,N_24564,N_24642);
or UO_1936 (O_1936,N_24435,N_24943);
nand UO_1937 (O_1937,N_24988,N_24327);
and UO_1938 (O_1938,N_24956,N_24091);
and UO_1939 (O_1939,N_24793,N_24461);
nand UO_1940 (O_1940,N_24725,N_24815);
or UO_1941 (O_1941,N_24897,N_24085);
nand UO_1942 (O_1942,N_24829,N_24270);
and UO_1943 (O_1943,N_24681,N_24890);
and UO_1944 (O_1944,N_24021,N_24965);
nor UO_1945 (O_1945,N_24883,N_24656);
and UO_1946 (O_1946,N_24235,N_24363);
and UO_1947 (O_1947,N_24653,N_24652);
and UO_1948 (O_1948,N_24412,N_24949);
or UO_1949 (O_1949,N_24704,N_24194);
and UO_1950 (O_1950,N_24453,N_24455);
nand UO_1951 (O_1951,N_24606,N_24376);
xnor UO_1952 (O_1952,N_24494,N_24757);
nand UO_1953 (O_1953,N_24897,N_24194);
nand UO_1954 (O_1954,N_24953,N_24621);
nor UO_1955 (O_1955,N_24952,N_24059);
nand UO_1956 (O_1956,N_24576,N_24341);
xnor UO_1957 (O_1957,N_24605,N_24903);
and UO_1958 (O_1958,N_24998,N_24731);
nand UO_1959 (O_1959,N_24280,N_24351);
nor UO_1960 (O_1960,N_24827,N_24033);
xnor UO_1961 (O_1961,N_24987,N_24703);
and UO_1962 (O_1962,N_24777,N_24743);
nand UO_1963 (O_1963,N_24950,N_24753);
or UO_1964 (O_1964,N_24312,N_24584);
nand UO_1965 (O_1965,N_24125,N_24852);
nand UO_1966 (O_1966,N_24416,N_24200);
or UO_1967 (O_1967,N_24464,N_24782);
and UO_1968 (O_1968,N_24389,N_24945);
nand UO_1969 (O_1969,N_24991,N_24188);
and UO_1970 (O_1970,N_24689,N_24203);
nand UO_1971 (O_1971,N_24203,N_24600);
nand UO_1972 (O_1972,N_24140,N_24496);
and UO_1973 (O_1973,N_24406,N_24570);
or UO_1974 (O_1974,N_24243,N_24665);
or UO_1975 (O_1975,N_24770,N_24131);
nand UO_1976 (O_1976,N_24828,N_24741);
or UO_1977 (O_1977,N_24763,N_24106);
nor UO_1978 (O_1978,N_24823,N_24656);
xnor UO_1979 (O_1979,N_24690,N_24423);
xnor UO_1980 (O_1980,N_24476,N_24909);
nand UO_1981 (O_1981,N_24372,N_24469);
nor UO_1982 (O_1982,N_24700,N_24892);
nor UO_1983 (O_1983,N_24881,N_24865);
xnor UO_1984 (O_1984,N_24390,N_24391);
xor UO_1985 (O_1985,N_24043,N_24004);
nand UO_1986 (O_1986,N_24182,N_24726);
or UO_1987 (O_1987,N_24818,N_24864);
or UO_1988 (O_1988,N_24090,N_24124);
nand UO_1989 (O_1989,N_24007,N_24676);
nand UO_1990 (O_1990,N_24747,N_24582);
xor UO_1991 (O_1991,N_24714,N_24680);
xor UO_1992 (O_1992,N_24837,N_24146);
xnor UO_1993 (O_1993,N_24198,N_24061);
xor UO_1994 (O_1994,N_24616,N_24928);
nand UO_1995 (O_1995,N_24348,N_24020);
and UO_1996 (O_1996,N_24666,N_24373);
and UO_1997 (O_1997,N_24623,N_24820);
and UO_1998 (O_1998,N_24345,N_24928);
or UO_1999 (O_1999,N_24324,N_24232);
and UO_2000 (O_2000,N_24236,N_24094);
nand UO_2001 (O_2001,N_24326,N_24159);
nand UO_2002 (O_2002,N_24230,N_24375);
or UO_2003 (O_2003,N_24551,N_24049);
xnor UO_2004 (O_2004,N_24200,N_24140);
or UO_2005 (O_2005,N_24116,N_24330);
nor UO_2006 (O_2006,N_24750,N_24193);
or UO_2007 (O_2007,N_24138,N_24377);
nand UO_2008 (O_2008,N_24721,N_24898);
nor UO_2009 (O_2009,N_24461,N_24975);
xnor UO_2010 (O_2010,N_24024,N_24015);
xnor UO_2011 (O_2011,N_24986,N_24304);
xor UO_2012 (O_2012,N_24592,N_24712);
or UO_2013 (O_2013,N_24298,N_24601);
xor UO_2014 (O_2014,N_24323,N_24859);
nand UO_2015 (O_2015,N_24834,N_24993);
or UO_2016 (O_2016,N_24351,N_24721);
nand UO_2017 (O_2017,N_24232,N_24991);
or UO_2018 (O_2018,N_24608,N_24863);
xor UO_2019 (O_2019,N_24100,N_24348);
nand UO_2020 (O_2020,N_24234,N_24043);
nor UO_2021 (O_2021,N_24548,N_24643);
and UO_2022 (O_2022,N_24315,N_24708);
xor UO_2023 (O_2023,N_24251,N_24281);
nor UO_2024 (O_2024,N_24640,N_24060);
nand UO_2025 (O_2025,N_24437,N_24755);
nor UO_2026 (O_2026,N_24791,N_24149);
nor UO_2027 (O_2027,N_24437,N_24267);
nor UO_2028 (O_2028,N_24268,N_24225);
nand UO_2029 (O_2029,N_24909,N_24958);
or UO_2030 (O_2030,N_24579,N_24447);
or UO_2031 (O_2031,N_24347,N_24880);
and UO_2032 (O_2032,N_24069,N_24401);
nand UO_2033 (O_2033,N_24325,N_24140);
xor UO_2034 (O_2034,N_24791,N_24367);
xnor UO_2035 (O_2035,N_24895,N_24202);
and UO_2036 (O_2036,N_24735,N_24001);
and UO_2037 (O_2037,N_24171,N_24614);
xnor UO_2038 (O_2038,N_24435,N_24824);
or UO_2039 (O_2039,N_24193,N_24295);
or UO_2040 (O_2040,N_24765,N_24932);
xor UO_2041 (O_2041,N_24311,N_24095);
or UO_2042 (O_2042,N_24075,N_24471);
nor UO_2043 (O_2043,N_24261,N_24869);
or UO_2044 (O_2044,N_24679,N_24125);
or UO_2045 (O_2045,N_24973,N_24613);
xor UO_2046 (O_2046,N_24118,N_24278);
nand UO_2047 (O_2047,N_24680,N_24170);
and UO_2048 (O_2048,N_24054,N_24254);
nand UO_2049 (O_2049,N_24762,N_24760);
xnor UO_2050 (O_2050,N_24010,N_24383);
nand UO_2051 (O_2051,N_24096,N_24205);
nand UO_2052 (O_2052,N_24185,N_24731);
xor UO_2053 (O_2053,N_24047,N_24653);
nor UO_2054 (O_2054,N_24824,N_24515);
and UO_2055 (O_2055,N_24294,N_24098);
or UO_2056 (O_2056,N_24654,N_24131);
xnor UO_2057 (O_2057,N_24788,N_24277);
or UO_2058 (O_2058,N_24046,N_24073);
xnor UO_2059 (O_2059,N_24189,N_24972);
xor UO_2060 (O_2060,N_24941,N_24674);
nor UO_2061 (O_2061,N_24191,N_24495);
xnor UO_2062 (O_2062,N_24389,N_24820);
and UO_2063 (O_2063,N_24191,N_24428);
and UO_2064 (O_2064,N_24837,N_24558);
or UO_2065 (O_2065,N_24691,N_24853);
and UO_2066 (O_2066,N_24305,N_24481);
xnor UO_2067 (O_2067,N_24943,N_24896);
or UO_2068 (O_2068,N_24265,N_24579);
and UO_2069 (O_2069,N_24358,N_24407);
xnor UO_2070 (O_2070,N_24375,N_24872);
and UO_2071 (O_2071,N_24330,N_24709);
nor UO_2072 (O_2072,N_24640,N_24527);
nand UO_2073 (O_2073,N_24823,N_24639);
nor UO_2074 (O_2074,N_24370,N_24947);
nand UO_2075 (O_2075,N_24667,N_24527);
nand UO_2076 (O_2076,N_24989,N_24646);
or UO_2077 (O_2077,N_24890,N_24737);
nor UO_2078 (O_2078,N_24762,N_24712);
and UO_2079 (O_2079,N_24394,N_24319);
and UO_2080 (O_2080,N_24973,N_24866);
xor UO_2081 (O_2081,N_24740,N_24328);
xor UO_2082 (O_2082,N_24180,N_24719);
xnor UO_2083 (O_2083,N_24112,N_24106);
and UO_2084 (O_2084,N_24995,N_24560);
and UO_2085 (O_2085,N_24550,N_24420);
or UO_2086 (O_2086,N_24371,N_24796);
or UO_2087 (O_2087,N_24334,N_24668);
xor UO_2088 (O_2088,N_24329,N_24801);
xor UO_2089 (O_2089,N_24060,N_24591);
nor UO_2090 (O_2090,N_24755,N_24041);
xnor UO_2091 (O_2091,N_24699,N_24262);
or UO_2092 (O_2092,N_24494,N_24066);
or UO_2093 (O_2093,N_24965,N_24810);
or UO_2094 (O_2094,N_24788,N_24040);
nor UO_2095 (O_2095,N_24200,N_24223);
xor UO_2096 (O_2096,N_24637,N_24069);
or UO_2097 (O_2097,N_24686,N_24904);
nor UO_2098 (O_2098,N_24456,N_24609);
xor UO_2099 (O_2099,N_24923,N_24698);
or UO_2100 (O_2100,N_24909,N_24854);
nand UO_2101 (O_2101,N_24053,N_24845);
nand UO_2102 (O_2102,N_24158,N_24455);
and UO_2103 (O_2103,N_24694,N_24869);
or UO_2104 (O_2104,N_24296,N_24009);
or UO_2105 (O_2105,N_24655,N_24434);
xnor UO_2106 (O_2106,N_24528,N_24727);
nand UO_2107 (O_2107,N_24205,N_24804);
and UO_2108 (O_2108,N_24571,N_24604);
nor UO_2109 (O_2109,N_24909,N_24633);
or UO_2110 (O_2110,N_24471,N_24020);
and UO_2111 (O_2111,N_24012,N_24832);
and UO_2112 (O_2112,N_24830,N_24663);
or UO_2113 (O_2113,N_24452,N_24648);
nor UO_2114 (O_2114,N_24684,N_24412);
xnor UO_2115 (O_2115,N_24775,N_24745);
nor UO_2116 (O_2116,N_24791,N_24949);
nand UO_2117 (O_2117,N_24635,N_24074);
and UO_2118 (O_2118,N_24565,N_24427);
nor UO_2119 (O_2119,N_24007,N_24512);
or UO_2120 (O_2120,N_24727,N_24116);
xnor UO_2121 (O_2121,N_24982,N_24590);
nor UO_2122 (O_2122,N_24742,N_24704);
and UO_2123 (O_2123,N_24089,N_24527);
nand UO_2124 (O_2124,N_24188,N_24263);
and UO_2125 (O_2125,N_24431,N_24834);
nand UO_2126 (O_2126,N_24387,N_24381);
xnor UO_2127 (O_2127,N_24439,N_24580);
or UO_2128 (O_2128,N_24939,N_24069);
xor UO_2129 (O_2129,N_24966,N_24995);
xnor UO_2130 (O_2130,N_24397,N_24660);
nand UO_2131 (O_2131,N_24249,N_24054);
and UO_2132 (O_2132,N_24042,N_24704);
xor UO_2133 (O_2133,N_24315,N_24938);
nor UO_2134 (O_2134,N_24077,N_24765);
and UO_2135 (O_2135,N_24234,N_24219);
and UO_2136 (O_2136,N_24203,N_24625);
or UO_2137 (O_2137,N_24073,N_24878);
xor UO_2138 (O_2138,N_24274,N_24324);
nand UO_2139 (O_2139,N_24749,N_24215);
nand UO_2140 (O_2140,N_24183,N_24364);
and UO_2141 (O_2141,N_24030,N_24328);
nor UO_2142 (O_2142,N_24143,N_24430);
xnor UO_2143 (O_2143,N_24836,N_24709);
or UO_2144 (O_2144,N_24936,N_24472);
nor UO_2145 (O_2145,N_24336,N_24750);
or UO_2146 (O_2146,N_24707,N_24108);
nand UO_2147 (O_2147,N_24732,N_24610);
and UO_2148 (O_2148,N_24639,N_24816);
xnor UO_2149 (O_2149,N_24533,N_24878);
and UO_2150 (O_2150,N_24702,N_24305);
nor UO_2151 (O_2151,N_24104,N_24516);
or UO_2152 (O_2152,N_24522,N_24171);
or UO_2153 (O_2153,N_24460,N_24587);
nand UO_2154 (O_2154,N_24849,N_24457);
and UO_2155 (O_2155,N_24486,N_24646);
or UO_2156 (O_2156,N_24717,N_24645);
or UO_2157 (O_2157,N_24817,N_24319);
or UO_2158 (O_2158,N_24373,N_24781);
and UO_2159 (O_2159,N_24348,N_24706);
nand UO_2160 (O_2160,N_24567,N_24161);
nor UO_2161 (O_2161,N_24808,N_24298);
xor UO_2162 (O_2162,N_24667,N_24555);
nand UO_2163 (O_2163,N_24576,N_24634);
xnor UO_2164 (O_2164,N_24253,N_24453);
or UO_2165 (O_2165,N_24668,N_24723);
nor UO_2166 (O_2166,N_24540,N_24589);
and UO_2167 (O_2167,N_24253,N_24854);
xnor UO_2168 (O_2168,N_24179,N_24376);
or UO_2169 (O_2169,N_24598,N_24494);
nor UO_2170 (O_2170,N_24776,N_24978);
nor UO_2171 (O_2171,N_24217,N_24256);
nand UO_2172 (O_2172,N_24491,N_24177);
and UO_2173 (O_2173,N_24691,N_24664);
nand UO_2174 (O_2174,N_24185,N_24328);
and UO_2175 (O_2175,N_24530,N_24521);
nand UO_2176 (O_2176,N_24166,N_24356);
nor UO_2177 (O_2177,N_24090,N_24601);
nor UO_2178 (O_2178,N_24113,N_24923);
or UO_2179 (O_2179,N_24485,N_24376);
and UO_2180 (O_2180,N_24944,N_24916);
or UO_2181 (O_2181,N_24707,N_24393);
or UO_2182 (O_2182,N_24822,N_24766);
or UO_2183 (O_2183,N_24210,N_24309);
nand UO_2184 (O_2184,N_24263,N_24445);
or UO_2185 (O_2185,N_24302,N_24283);
xor UO_2186 (O_2186,N_24338,N_24206);
and UO_2187 (O_2187,N_24141,N_24095);
or UO_2188 (O_2188,N_24607,N_24612);
xor UO_2189 (O_2189,N_24669,N_24138);
nor UO_2190 (O_2190,N_24393,N_24526);
and UO_2191 (O_2191,N_24674,N_24130);
xnor UO_2192 (O_2192,N_24881,N_24564);
or UO_2193 (O_2193,N_24242,N_24259);
xnor UO_2194 (O_2194,N_24699,N_24827);
or UO_2195 (O_2195,N_24710,N_24882);
xnor UO_2196 (O_2196,N_24262,N_24438);
and UO_2197 (O_2197,N_24026,N_24042);
and UO_2198 (O_2198,N_24589,N_24739);
or UO_2199 (O_2199,N_24618,N_24736);
nor UO_2200 (O_2200,N_24171,N_24928);
nor UO_2201 (O_2201,N_24578,N_24111);
and UO_2202 (O_2202,N_24563,N_24120);
or UO_2203 (O_2203,N_24485,N_24980);
nand UO_2204 (O_2204,N_24354,N_24709);
or UO_2205 (O_2205,N_24984,N_24353);
and UO_2206 (O_2206,N_24816,N_24765);
and UO_2207 (O_2207,N_24819,N_24176);
and UO_2208 (O_2208,N_24290,N_24105);
nor UO_2209 (O_2209,N_24195,N_24394);
nand UO_2210 (O_2210,N_24456,N_24091);
or UO_2211 (O_2211,N_24055,N_24598);
nor UO_2212 (O_2212,N_24894,N_24783);
xnor UO_2213 (O_2213,N_24900,N_24834);
nor UO_2214 (O_2214,N_24099,N_24975);
and UO_2215 (O_2215,N_24746,N_24665);
nor UO_2216 (O_2216,N_24702,N_24728);
or UO_2217 (O_2217,N_24919,N_24167);
and UO_2218 (O_2218,N_24845,N_24139);
nand UO_2219 (O_2219,N_24956,N_24200);
and UO_2220 (O_2220,N_24632,N_24430);
or UO_2221 (O_2221,N_24851,N_24543);
nand UO_2222 (O_2222,N_24201,N_24071);
and UO_2223 (O_2223,N_24996,N_24180);
xor UO_2224 (O_2224,N_24652,N_24783);
and UO_2225 (O_2225,N_24197,N_24772);
nand UO_2226 (O_2226,N_24842,N_24329);
nand UO_2227 (O_2227,N_24258,N_24510);
xor UO_2228 (O_2228,N_24308,N_24967);
nor UO_2229 (O_2229,N_24378,N_24753);
nand UO_2230 (O_2230,N_24574,N_24668);
or UO_2231 (O_2231,N_24051,N_24447);
or UO_2232 (O_2232,N_24056,N_24411);
nor UO_2233 (O_2233,N_24463,N_24917);
or UO_2234 (O_2234,N_24939,N_24080);
and UO_2235 (O_2235,N_24622,N_24440);
and UO_2236 (O_2236,N_24315,N_24191);
nor UO_2237 (O_2237,N_24799,N_24741);
or UO_2238 (O_2238,N_24460,N_24935);
nand UO_2239 (O_2239,N_24762,N_24968);
and UO_2240 (O_2240,N_24401,N_24671);
and UO_2241 (O_2241,N_24456,N_24365);
or UO_2242 (O_2242,N_24388,N_24335);
nand UO_2243 (O_2243,N_24294,N_24684);
and UO_2244 (O_2244,N_24648,N_24821);
xor UO_2245 (O_2245,N_24663,N_24611);
or UO_2246 (O_2246,N_24335,N_24208);
and UO_2247 (O_2247,N_24396,N_24150);
nor UO_2248 (O_2248,N_24747,N_24407);
and UO_2249 (O_2249,N_24950,N_24241);
nor UO_2250 (O_2250,N_24779,N_24013);
nor UO_2251 (O_2251,N_24167,N_24334);
nor UO_2252 (O_2252,N_24019,N_24363);
and UO_2253 (O_2253,N_24676,N_24457);
nor UO_2254 (O_2254,N_24479,N_24679);
or UO_2255 (O_2255,N_24480,N_24824);
or UO_2256 (O_2256,N_24862,N_24135);
nand UO_2257 (O_2257,N_24149,N_24378);
nor UO_2258 (O_2258,N_24690,N_24260);
nand UO_2259 (O_2259,N_24966,N_24369);
xor UO_2260 (O_2260,N_24805,N_24891);
nand UO_2261 (O_2261,N_24420,N_24913);
or UO_2262 (O_2262,N_24260,N_24298);
nand UO_2263 (O_2263,N_24022,N_24675);
xnor UO_2264 (O_2264,N_24616,N_24267);
nand UO_2265 (O_2265,N_24079,N_24928);
xor UO_2266 (O_2266,N_24914,N_24655);
xor UO_2267 (O_2267,N_24189,N_24667);
nand UO_2268 (O_2268,N_24806,N_24396);
xor UO_2269 (O_2269,N_24013,N_24708);
xor UO_2270 (O_2270,N_24354,N_24495);
or UO_2271 (O_2271,N_24846,N_24213);
and UO_2272 (O_2272,N_24735,N_24529);
nand UO_2273 (O_2273,N_24093,N_24621);
nand UO_2274 (O_2274,N_24440,N_24317);
and UO_2275 (O_2275,N_24172,N_24298);
nand UO_2276 (O_2276,N_24259,N_24247);
xnor UO_2277 (O_2277,N_24565,N_24740);
or UO_2278 (O_2278,N_24200,N_24308);
and UO_2279 (O_2279,N_24241,N_24931);
nand UO_2280 (O_2280,N_24210,N_24085);
nand UO_2281 (O_2281,N_24284,N_24918);
nor UO_2282 (O_2282,N_24006,N_24465);
and UO_2283 (O_2283,N_24263,N_24384);
nand UO_2284 (O_2284,N_24417,N_24409);
nor UO_2285 (O_2285,N_24190,N_24255);
nand UO_2286 (O_2286,N_24884,N_24193);
nor UO_2287 (O_2287,N_24254,N_24193);
xor UO_2288 (O_2288,N_24877,N_24857);
or UO_2289 (O_2289,N_24363,N_24867);
xor UO_2290 (O_2290,N_24389,N_24913);
nand UO_2291 (O_2291,N_24056,N_24792);
nor UO_2292 (O_2292,N_24179,N_24614);
nand UO_2293 (O_2293,N_24966,N_24075);
or UO_2294 (O_2294,N_24561,N_24080);
nor UO_2295 (O_2295,N_24128,N_24715);
xnor UO_2296 (O_2296,N_24888,N_24820);
xnor UO_2297 (O_2297,N_24210,N_24859);
nand UO_2298 (O_2298,N_24400,N_24209);
nand UO_2299 (O_2299,N_24164,N_24168);
nor UO_2300 (O_2300,N_24753,N_24346);
xnor UO_2301 (O_2301,N_24572,N_24739);
nand UO_2302 (O_2302,N_24710,N_24272);
nand UO_2303 (O_2303,N_24774,N_24460);
and UO_2304 (O_2304,N_24716,N_24078);
and UO_2305 (O_2305,N_24937,N_24267);
xor UO_2306 (O_2306,N_24273,N_24861);
nor UO_2307 (O_2307,N_24590,N_24623);
xor UO_2308 (O_2308,N_24469,N_24770);
nor UO_2309 (O_2309,N_24898,N_24131);
or UO_2310 (O_2310,N_24884,N_24321);
or UO_2311 (O_2311,N_24477,N_24435);
and UO_2312 (O_2312,N_24394,N_24040);
xor UO_2313 (O_2313,N_24934,N_24958);
xor UO_2314 (O_2314,N_24130,N_24451);
and UO_2315 (O_2315,N_24034,N_24635);
xor UO_2316 (O_2316,N_24488,N_24531);
and UO_2317 (O_2317,N_24927,N_24740);
nand UO_2318 (O_2318,N_24166,N_24740);
nand UO_2319 (O_2319,N_24973,N_24238);
xnor UO_2320 (O_2320,N_24499,N_24517);
xor UO_2321 (O_2321,N_24084,N_24824);
and UO_2322 (O_2322,N_24727,N_24467);
nand UO_2323 (O_2323,N_24945,N_24150);
and UO_2324 (O_2324,N_24589,N_24366);
nand UO_2325 (O_2325,N_24316,N_24540);
nor UO_2326 (O_2326,N_24407,N_24878);
and UO_2327 (O_2327,N_24171,N_24542);
or UO_2328 (O_2328,N_24975,N_24931);
and UO_2329 (O_2329,N_24336,N_24098);
or UO_2330 (O_2330,N_24143,N_24564);
and UO_2331 (O_2331,N_24193,N_24683);
xnor UO_2332 (O_2332,N_24390,N_24970);
xor UO_2333 (O_2333,N_24311,N_24400);
xor UO_2334 (O_2334,N_24084,N_24806);
nor UO_2335 (O_2335,N_24855,N_24618);
and UO_2336 (O_2336,N_24012,N_24058);
nand UO_2337 (O_2337,N_24596,N_24438);
or UO_2338 (O_2338,N_24253,N_24041);
nand UO_2339 (O_2339,N_24165,N_24219);
or UO_2340 (O_2340,N_24328,N_24657);
nand UO_2341 (O_2341,N_24362,N_24554);
or UO_2342 (O_2342,N_24508,N_24360);
nor UO_2343 (O_2343,N_24836,N_24559);
and UO_2344 (O_2344,N_24389,N_24785);
nand UO_2345 (O_2345,N_24712,N_24217);
nor UO_2346 (O_2346,N_24699,N_24071);
and UO_2347 (O_2347,N_24153,N_24137);
nor UO_2348 (O_2348,N_24698,N_24991);
and UO_2349 (O_2349,N_24841,N_24330);
xor UO_2350 (O_2350,N_24854,N_24173);
and UO_2351 (O_2351,N_24062,N_24939);
and UO_2352 (O_2352,N_24609,N_24934);
nor UO_2353 (O_2353,N_24121,N_24235);
and UO_2354 (O_2354,N_24142,N_24809);
and UO_2355 (O_2355,N_24569,N_24553);
nand UO_2356 (O_2356,N_24647,N_24739);
nand UO_2357 (O_2357,N_24456,N_24555);
and UO_2358 (O_2358,N_24552,N_24971);
nor UO_2359 (O_2359,N_24391,N_24261);
nor UO_2360 (O_2360,N_24861,N_24350);
nor UO_2361 (O_2361,N_24131,N_24335);
and UO_2362 (O_2362,N_24383,N_24811);
and UO_2363 (O_2363,N_24326,N_24780);
nand UO_2364 (O_2364,N_24623,N_24266);
or UO_2365 (O_2365,N_24247,N_24407);
xnor UO_2366 (O_2366,N_24971,N_24129);
and UO_2367 (O_2367,N_24240,N_24870);
xor UO_2368 (O_2368,N_24277,N_24881);
nand UO_2369 (O_2369,N_24994,N_24381);
or UO_2370 (O_2370,N_24051,N_24202);
xor UO_2371 (O_2371,N_24954,N_24212);
nor UO_2372 (O_2372,N_24597,N_24683);
or UO_2373 (O_2373,N_24863,N_24707);
xnor UO_2374 (O_2374,N_24681,N_24811);
xnor UO_2375 (O_2375,N_24457,N_24851);
nand UO_2376 (O_2376,N_24709,N_24722);
and UO_2377 (O_2377,N_24414,N_24258);
nand UO_2378 (O_2378,N_24280,N_24979);
nand UO_2379 (O_2379,N_24231,N_24315);
nand UO_2380 (O_2380,N_24953,N_24632);
nor UO_2381 (O_2381,N_24788,N_24663);
xor UO_2382 (O_2382,N_24948,N_24725);
nor UO_2383 (O_2383,N_24013,N_24069);
and UO_2384 (O_2384,N_24142,N_24875);
nor UO_2385 (O_2385,N_24992,N_24196);
and UO_2386 (O_2386,N_24385,N_24789);
and UO_2387 (O_2387,N_24381,N_24044);
and UO_2388 (O_2388,N_24466,N_24069);
or UO_2389 (O_2389,N_24617,N_24573);
xor UO_2390 (O_2390,N_24010,N_24697);
nor UO_2391 (O_2391,N_24129,N_24490);
or UO_2392 (O_2392,N_24914,N_24373);
nand UO_2393 (O_2393,N_24282,N_24765);
xor UO_2394 (O_2394,N_24779,N_24572);
nor UO_2395 (O_2395,N_24515,N_24088);
xor UO_2396 (O_2396,N_24613,N_24360);
xor UO_2397 (O_2397,N_24992,N_24003);
nor UO_2398 (O_2398,N_24625,N_24240);
or UO_2399 (O_2399,N_24613,N_24039);
xor UO_2400 (O_2400,N_24592,N_24812);
nor UO_2401 (O_2401,N_24117,N_24860);
or UO_2402 (O_2402,N_24606,N_24207);
and UO_2403 (O_2403,N_24205,N_24505);
nand UO_2404 (O_2404,N_24622,N_24031);
xor UO_2405 (O_2405,N_24482,N_24587);
xor UO_2406 (O_2406,N_24733,N_24040);
or UO_2407 (O_2407,N_24922,N_24539);
nand UO_2408 (O_2408,N_24021,N_24231);
nor UO_2409 (O_2409,N_24505,N_24602);
nor UO_2410 (O_2410,N_24895,N_24327);
nand UO_2411 (O_2411,N_24450,N_24264);
nand UO_2412 (O_2412,N_24956,N_24369);
nor UO_2413 (O_2413,N_24515,N_24686);
xnor UO_2414 (O_2414,N_24116,N_24170);
nor UO_2415 (O_2415,N_24420,N_24708);
nand UO_2416 (O_2416,N_24059,N_24358);
nand UO_2417 (O_2417,N_24589,N_24331);
nor UO_2418 (O_2418,N_24722,N_24171);
and UO_2419 (O_2419,N_24625,N_24749);
nor UO_2420 (O_2420,N_24683,N_24781);
nor UO_2421 (O_2421,N_24702,N_24515);
nand UO_2422 (O_2422,N_24761,N_24436);
xnor UO_2423 (O_2423,N_24444,N_24306);
nand UO_2424 (O_2424,N_24086,N_24680);
xor UO_2425 (O_2425,N_24138,N_24586);
or UO_2426 (O_2426,N_24448,N_24324);
nand UO_2427 (O_2427,N_24190,N_24469);
or UO_2428 (O_2428,N_24939,N_24211);
and UO_2429 (O_2429,N_24578,N_24743);
xor UO_2430 (O_2430,N_24606,N_24466);
nand UO_2431 (O_2431,N_24706,N_24693);
nor UO_2432 (O_2432,N_24657,N_24082);
nand UO_2433 (O_2433,N_24175,N_24663);
or UO_2434 (O_2434,N_24555,N_24496);
or UO_2435 (O_2435,N_24486,N_24923);
and UO_2436 (O_2436,N_24800,N_24746);
or UO_2437 (O_2437,N_24227,N_24069);
xnor UO_2438 (O_2438,N_24536,N_24729);
and UO_2439 (O_2439,N_24361,N_24299);
nor UO_2440 (O_2440,N_24131,N_24436);
nand UO_2441 (O_2441,N_24181,N_24017);
nor UO_2442 (O_2442,N_24939,N_24125);
nand UO_2443 (O_2443,N_24763,N_24847);
xor UO_2444 (O_2444,N_24008,N_24964);
and UO_2445 (O_2445,N_24734,N_24984);
nor UO_2446 (O_2446,N_24166,N_24162);
nor UO_2447 (O_2447,N_24104,N_24015);
nand UO_2448 (O_2448,N_24644,N_24223);
nand UO_2449 (O_2449,N_24057,N_24665);
nor UO_2450 (O_2450,N_24766,N_24360);
xnor UO_2451 (O_2451,N_24249,N_24576);
and UO_2452 (O_2452,N_24814,N_24042);
nor UO_2453 (O_2453,N_24826,N_24392);
nor UO_2454 (O_2454,N_24160,N_24662);
xor UO_2455 (O_2455,N_24801,N_24886);
nor UO_2456 (O_2456,N_24201,N_24149);
and UO_2457 (O_2457,N_24680,N_24949);
nand UO_2458 (O_2458,N_24320,N_24225);
xnor UO_2459 (O_2459,N_24523,N_24962);
xor UO_2460 (O_2460,N_24314,N_24073);
or UO_2461 (O_2461,N_24199,N_24466);
xor UO_2462 (O_2462,N_24334,N_24973);
or UO_2463 (O_2463,N_24544,N_24270);
xnor UO_2464 (O_2464,N_24052,N_24585);
nand UO_2465 (O_2465,N_24354,N_24124);
or UO_2466 (O_2466,N_24334,N_24089);
and UO_2467 (O_2467,N_24932,N_24257);
and UO_2468 (O_2468,N_24414,N_24875);
xnor UO_2469 (O_2469,N_24318,N_24532);
nand UO_2470 (O_2470,N_24765,N_24899);
nand UO_2471 (O_2471,N_24564,N_24156);
xor UO_2472 (O_2472,N_24515,N_24687);
or UO_2473 (O_2473,N_24625,N_24926);
nand UO_2474 (O_2474,N_24320,N_24631);
nor UO_2475 (O_2475,N_24721,N_24912);
xor UO_2476 (O_2476,N_24667,N_24012);
and UO_2477 (O_2477,N_24397,N_24528);
and UO_2478 (O_2478,N_24616,N_24245);
xnor UO_2479 (O_2479,N_24711,N_24858);
nor UO_2480 (O_2480,N_24599,N_24944);
or UO_2481 (O_2481,N_24476,N_24818);
nand UO_2482 (O_2482,N_24914,N_24633);
nor UO_2483 (O_2483,N_24143,N_24922);
nand UO_2484 (O_2484,N_24095,N_24227);
nor UO_2485 (O_2485,N_24523,N_24041);
or UO_2486 (O_2486,N_24215,N_24683);
and UO_2487 (O_2487,N_24659,N_24592);
nand UO_2488 (O_2488,N_24079,N_24394);
xor UO_2489 (O_2489,N_24980,N_24525);
or UO_2490 (O_2490,N_24830,N_24231);
xnor UO_2491 (O_2491,N_24438,N_24369);
or UO_2492 (O_2492,N_24479,N_24385);
or UO_2493 (O_2493,N_24126,N_24067);
or UO_2494 (O_2494,N_24068,N_24943);
nor UO_2495 (O_2495,N_24534,N_24163);
or UO_2496 (O_2496,N_24709,N_24418);
xnor UO_2497 (O_2497,N_24773,N_24567);
or UO_2498 (O_2498,N_24680,N_24262);
nor UO_2499 (O_2499,N_24923,N_24772);
or UO_2500 (O_2500,N_24401,N_24098);
or UO_2501 (O_2501,N_24492,N_24400);
xnor UO_2502 (O_2502,N_24728,N_24073);
or UO_2503 (O_2503,N_24113,N_24333);
nand UO_2504 (O_2504,N_24951,N_24781);
xor UO_2505 (O_2505,N_24477,N_24610);
nor UO_2506 (O_2506,N_24459,N_24614);
and UO_2507 (O_2507,N_24648,N_24880);
nor UO_2508 (O_2508,N_24377,N_24447);
and UO_2509 (O_2509,N_24371,N_24375);
nor UO_2510 (O_2510,N_24352,N_24970);
xor UO_2511 (O_2511,N_24059,N_24374);
and UO_2512 (O_2512,N_24841,N_24129);
nor UO_2513 (O_2513,N_24353,N_24407);
nand UO_2514 (O_2514,N_24009,N_24073);
nand UO_2515 (O_2515,N_24273,N_24537);
nand UO_2516 (O_2516,N_24318,N_24134);
and UO_2517 (O_2517,N_24511,N_24530);
or UO_2518 (O_2518,N_24542,N_24358);
xor UO_2519 (O_2519,N_24941,N_24108);
nand UO_2520 (O_2520,N_24038,N_24595);
or UO_2521 (O_2521,N_24313,N_24128);
or UO_2522 (O_2522,N_24382,N_24435);
nand UO_2523 (O_2523,N_24196,N_24265);
and UO_2524 (O_2524,N_24743,N_24726);
or UO_2525 (O_2525,N_24660,N_24502);
or UO_2526 (O_2526,N_24379,N_24800);
xnor UO_2527 (O_2527,N_24390,N_24484);
and UO_2528 (O_2528,N_24626,N_24453);
and UO_2529 (O_2529,N_24614,N_24268);
nand UO_2530 (O_2530,N_24157,N_24197);
nor UO_2531 (O_2531,N_24476,N_24651);
or UO_2532 (O_2532,N_24130,N_24720);
and UO_2533 (O_2533,N_24889,N_24819);
nor UO_2534 (O_2534,N_24361,N_24759);
and UO_2535 (O_2535,N_24530,N_24527);
nand UO_2536 (O_2536,N_24824,N_24110);
nor UO_2537 (O_2537,N_24624,N_24366);
and UO_2538 (O_2538,N_24096,N_24232);
xor UO_2539 (O_2539,N_24033,N_24463);
or UO_2540 (O_2540,N_24318,N_24107);
nor UO_2541 (O_2541,N_24355,N_24633);
and UO_2542 (O_2542,N_24072,N_24293);
xnor UO_2543 (O_2543,N_24255,N_24483);
nand UO_2544 (O_2544,N_24020,N_24200);
xnor UO_2545 (O_2545,N_24014,N_24160);
and UO_2546 (O_2546,N_24649,N_24756);
nor UO_2547 (O_2547,N_24038,N_24155);
nand UO_2548 (O_2548,N_24569,N_24265);
nand UO_2549 (O_2549,N_24766,N_24399);
xor UO_2550 (O_2550,N_24550,N_24025);
nand UO_2551 (O_2551,N_24735,N_24766);
and UO_2552 (O_2552,N_24208,N_24812);
xnor UO_2553 (O_2553,N_24518,N_24864);
or UO_2554 (O_2554,N_24370,N_24501);
nor UO_2555 (O_2555,N_24546,N_24156);
and UO_2556 (O_2556,N_24315,N_24181);
xnor UO_2557 (O_2557,N_24964,N_24985);
nand UO_2558 (O_2558,N_24398,N_24592);
and UO_2559 (O_2559,N_24516,N_24076);
xor UO_2560 (O_2560,N_24570,N_24830);
nor UO_2561 (O_2561,N_24963,N_24627);
and UO_2562 (O_2562,N_24378,N_24784);
nand UO_2563 (O_2563,N_24416,N_24367);
and UO_2564 (O_2564,N_24046,N_24135);
and UO_2565 (O_2565,N_24063,N_24087);
xor UO_2566 (O_2566,N_24650,N_24289);
nor UO_2567 (O_2567,N_24827,N_24284);
nor UO_2568 (O_2568,N_24204,N_24355);
xnor UO_2569 (O_2569,N_24338,N_24254);
xor UO_2570 (O_2570,N_24336,N_24080);
or UO_2571 (O_2571,N_24651,N_24009);
nor UO_2572 (O_2572,N_24691,N_24545);
and UO_2573 (O_2573,N_24579,N_24008);
nor UO_2574 (O_2574,N_24509,N_24681);
nand UO_2575 (O_2575,N_24393,N_24343);
and UO_2576 (O_2576,N_24909,N_24814);
xor UO_2577 (O_2577,N_24732,N_24011);
nor UO_2578 (O_2578,N_24103,N_24227);
or UO_2579 (O_2579,N_24822,N_24540);
nand UO_2580 (O_2580,N_24321,N_24324);
or UO_2581 (O_2581,N_24440,N_24170);
nand UO_2582 (O_2582,N_24719,N_24474);
nand UO_2583 (O_2583,N_24364,N_24396);
nor UO_2584 (O_2584,N_24689,N_24858);
nor UO_2585 (O_2585,N_24729,N_24211);
or UO_2586 (O_2586,N_24433,N_24816);
xnor UO_2587 (O_2587,N_24263,N_24982);
and UO_2588 (O_2588,N_24975,N_24238);
or UO_2589 (O_2589,N_24783,N_24581);
xor UO_2590 (O_2590,N_24081,N_24677);
nand UO_2591 (O_2591,N_24972,N_24089);
nor UO_2592 (O_2592,N_24033,N_24603);
or UO_2593 (O_2593,N_24842,N_24550);
nor UO_2594 (O_2594,N_24371,N_24848);
or UO_2595 (O_2595,N_24574,N_24197);
nor UO_2596 (O_2596,N_24979,N_24441);
and UO_2597 (O_2597,N_24688,N_24162);
nand UO_2598 (O_2598,N_24276,N_24854);
nor UO_2599 (O_2599,N_24192,N_24963);
nor UO_2600 (O_2600,N_24710,N_24528);
xor UO_2601 (O_2601,N_24471,N_24344);
nor UO_2602 (O_2602,N_24474,N_24886);
or UO_2603 (O_2603,N_24844,N_24411);
or UO_2604 (O_2604,N_24929,N_24811);
xnor UO_2605 (O_2605,N_24415,N_24065);
and UO_2606 (O_2606,N_24855,N_24398);
and UO_2607 (O_2607,N_24737,N_24048);
nand UO_2608 (O_2608,N_24682,N_24876);
xor UO_2609 (O_2609,N_24845,N_24336);
or UO_2610 (O_2610,N_24825,N_24009);
nor UO_2611 (O_2611,N_24484,N_24498);
xnor UO_2612 (O_2612,N_24337,N_24695);
nand UO_2613 (O_2613,N_24237,N_24644);
or UO_2614 (O_2614,N_24961,N_24996);
nor UO_2615 (O_2615,N_24229,N_24127);
xor UO_2616 (O_2616,N_24020,N_24890);
nor UO_2617 (O_2617,N_24754,N_24138);
or UO_2618 (O_2618,N_24745,N_24070);
and UO_2619 (O_2619,N_24663,N_24878);
nor UO_2620 (O_2620,N_24264,N_24359);
or UO_2621 (O_2621,N_24688,N_24240);
and UO_2622 (O_2622,N_24260,N_24267);
and UO_2623 (O_2623,N_24089,N_24653);
nand UO_2624 (O_2624,N_24853,N_24217);
and UO_2625 (O_2625,N_24560,N_24541);
nor UO_2626 (O_2626,N_24540,N_24768);
nor UO_2627 (O_2627,N_24556,N_24038);
nand UO_2628 (O_2628,N_24625,N_24563);
and UO_2629 (O_2629,N_24667,N_24411);
xnor UO_2630 (O_2630,N_24348,N_24992);
nor UO_2631 (O_2631,N_24023,N_24935);
nor UO_2632 (O_2632,N_24168,N_24891);
and UO_2633 (O_2633,N_24169,N_24886);
and UO_2634 (O_2634,N_24628,N_24266);
or UO_2635 (O_2635,N_24597,N_24891);
or UO_2636 (O_2636,N_24950,N_24342);
nor UO_2637 (O_2637,N_24393,N_24291);
or UO_2638 (O_2638,N_24797,N_24291);
xor UO_2639 (O_2639,N_24365,N_24067);
or UO_2640 (O_2640,N_24658,N_24914);
nand UO_2641 (O_2641,N_24811,N_24471);
or UO_2642 (O_2642,N_24420,N_24797);
nor UO_2643 (O_2643,N_24118,N_24232);
nand UO_2644 (O_2644,N_24342,N_24229);
or UO_2645 (O_2645,N_24716,N_24818);
or UO_2646 (O_2646,N_24923,N_24337);
xor UO_2647 (O_2647,N_24113,N_24484);
and UO_2648 (O_2648,N_24939,N_24774);
nor UO_2649 (O_2649,N_24227,N_24948);
or UO_2650 (O_2650,N_24735,N_24758);
and UO_2651 (O_2651,N_24792,N_24176);
and UO_2652 (O_2652,N_24931,N_24929);
nand UO_2653 (O_2653,N_24674,N_24188);
nand UO_2654 (O_2654,N_24197,N_24424);
xnor UO_2655 (O_2655,N_24848,N_24882);
nor UO_2656 (O_2656,N_24802,N_24935);
and UO_2657 (O_2657,N_24671,N_24030);
or UO_2658 (O_2658,N_24040,N_24997);
nor UO_2659 (O_2659,N_24996,N_24260);
xor UO_2660 (O_2660,N_24023,N_24846);
and UO_2661 (O_2661,N_24316,N_24640);
or UO_2662 (O_2662,N_24609,N_24904);
xor UO_2663 (O_2663,N_24886,N_24604);
nor UO_2664 (O_2664,N_24540,N_24660);
and UO_2665 (O_2665,N_24970,N_24649);
xor UO_2666 (O_2666,N_24907,N_24644);
nand UO_2667 (O_2667,N_24517,N_24216);
and UO_2668 (O_2668,N_24409,N_24655);
xnor UO_2669 (O_2669,N_24475,N_24754);
and UO_2670 (O_2670,N_24419,N_24964);
or UO_2671 (O_2671,N_24881,N_24840);
or UO_2672 (O_2672,N_24316,N_24623);
or UO_2673 (O_2673,N_24373,N_24464);
nor UO_2674 (O_2674,N_24973,N_24799);
nor UO_2675 (O_2675,N_24220,N_24964);
and UO_2676 (O_2676,N_24553,N_24238);
nor UO_2677 (O_2677,N_24795,N_24339);
nand UO_2678 (O_2678,N_24945,N_24409);
nor UO_2679 (O_2679,N_24552,N_24931);
and UO_2680 (O_2680,N_24938,N_24204);
or UO_2681 (O_2681,N_24685,N_24186);
and UO_2682 (O_2682,N_24137,N_24065);
and UO_2683 (O_2683,N_24892,N_24835);
xnor UO_2684 (O_2684,N_24070,N_24458);
nand UO_2685 (O_2685,N_24819,N_24001);
xnor UO_2686 (O_2686,N_24220,N_24131);
nand UO_2687 (O_2687,N_24346,N_24093);
and UO_2688 (O_2688,N_24094,N_24058);
or UO_2689 (O_2689,N_24180,N_24568);
xnor UO_2690 (O_2690,N_24780,N_24688);
nor UO_2691 (O_2691,N_24619,N_24844);
nor UO_2692 (O_2692,N_24903,N_24552);
xnor UO_2693 (O_2693,N_24760,N_24783);
nor UO_2694 (O_2694,N_24083,N_24469);
nor UO_2695 (O_2695,N_24446,N_24117);
nand UO_2696 (O_2696,N_24153,N_24085);
or UO_2697 (O_2697,N_24116,N_24205);
or UO_2698 (O_2698,N_24911,N_24566);
xnor UO_2699 (O_2699,N_24295,N_24207);
or UO_2700 (O_2700,N_24768,N_24520);
nor UO_2701 (O_2701,N_24835,N_24723);
or UO_2702 (O_2702,N_24968,N_24908);
nor UO_2703 (O_2703,N_24630,N_24728);
nand UO_2704 (O_2704,N_24443,N_24510);
nor UO_2705 (O_2705,N_24122,N_24253);
xor UO_2706 (O_2706,N_24818,N_24685);
and UO_2707 (O_2707,N_24700,N_24996);
xnor UO_2708 (O_2708,N_24388,N_24094);
and UO_2709 (O_2709,N_24620,N_24274);
or UO_2710 (O_2710,N_24950,N_24520);
and UO_2711 (O_2711,N_24501,N_24992);
nor UO_2712 (O_2712,N_24585,N_24549);
nand UO_2713 (O_2713,N_24816,N_24167);
or UO_2714 (O_2714,N_24214,N_24823);
and UO_2715 (O_2715,N_24940,N_24462);
or UO_2716 (O_2716,N_24046,N_24306);
or UO_2717 (O_2717,N_24822,N_24523);
or UO_2718 (O_2718,N_24265,N_24330);
nor UO_2719 (O_2719,N_24197,N_24966);
xor UO_2720 (O_2720,N_24120,N_24562);
nand UO_2721 (O_2721,N_24152,N_24606);
nand UO_2722 (O_2722,N_24178,N_24954);
nand UO_2723 (O_2723,N_24567,N_24499);
nor UO_2724 (O_2724,N_24162,N_24090);
or UO_2725 (O_2725,N_24630,N_24069);
nor UO_2726 (O_2726,N_24157,N_24875);
or UO_2727 (O_2727,N_24077,N_24330);
xnor UO_2728 (O_2728,N_24856,N_24158);
and UO_2729 (O_2729,N_24384,N_24446);
nand UO_2730 (O_2730,N_24585,N_24752);
or UO_2731 (O_2731,N_24863,N_24871);
or UO_2732 (O_2732,N_24620,N_24246);
nor UO_2733 (O_2733,N_24648,N_24182);
nand UO_2734 (O_2734,N_24474,N_24394);
nand UO_2735 (O_2735,N_24990,N_24880);
and UO_2736 (O_2736,N_24147,N_24789);
nor UO_2737 (O_2737,N_24718,N_24895);
or UO_2738 (O_2738,N_24508,N_24743);
nand UO_2739 (O_2739,N_24506,N_24559);
nand UO_2740 (O_2740,N_24963,N_24116);
xor UO_2741 (O_2741,N_24731,N_24982);
and UO_2742 (O_2742,N_24211,N_24998);
nor UO_2743 (O_2743,N_24257,N_24264);
nand UO_2744 (O_2744,N_24505,N_24410);
and UO_2745 (O_2745,N_24838,N_24485);
nand UO_2746 (O_2746,N_24495,N_24073);
and UO_2747 (O_2747,N_24785,N_24635);
or UO_2748 (O_2748,N_24551,N_24100);
xor UO_2749 (O_2749,N_24004,N_24076);
and UO_2750 (O_2750,N_24460,N_24169);
or UO_2751 (O_2751,N_24202,N_24630);
and UO_2752 (O_2752,N_24601,N_24993);
nand UO_2753 (O_2753,N_24900,N_24069);
nor UO_2754 (O_2754,N_24351,N_24009);
or UO_2755 (O_2755,N_24316,N_24332);
nor UO_2756 (O_2756,N_24923,N_24351);
and UO_2757 (O_2757,N_24397,N_24327);
and UO_2758 (O_2758,N_24080,N_24721);
and UO_2759 (O_2759,N_24891,N_24181);
nand UO_2760 (O_2760,N_24003,N_24811);
xor UO_2761 (O_2761,N_24203,N_24715);
nor UO_2762 (O_2762,N_24325,N_24991);
nand UO_2763 (O_2763,N_24622,N_24669);
nand UO_2764 (O_2764,N_24617,N_24612);
or UO_2765 (O_2765,N_24153,N_24414);
or UO_2766 (O_2766,N_24003,N_24868);
nand UO_2767 (O_2767,N_24606,N_24085);
or UO_2768 (O_2768,N_24372,N_24604);
xor UO_2769 (O_2769,N_24182,N_24047);
nor UO_2770 (O_2770,N_24129,N_24427);
nand UO_2771 (O_2771,N_24685,N_24929);
nand UO_2772 (O_2772,N_24939,N_24671);
or UO_2773 (O_2773,N_24635,N_24418);
nor UO_2774 (O_2774,N_24892,N_24196);
nand UO_2775 (O_2775,N_24406,N_24673);
xnor UO_2776 (O_2776,N_24472,N_24692);
nand UO_2777 (O_2777,N_24022,N_24036);
or UO_2778 (O_2778,N_24246,N_24651);
and UO_2779 (O_2779,N_24972,N_24620);
xor UO_2780 (O_2780,N_24891,N_24812);
nor UO_2781 (O_2781,N_24395,N_24720);
nor UO_2782 (O_2782,N_24436,N_24988);
or UO_2783 (O_2783,N_24595,N_24306);
nor UO_2784 (O_2784,N_24277,N_24963);
nand UO_2785 (O_2785,N_24222,N_24760);
nor UO_2786 (O_2786,N_24744,N_24135);
or UO_2787 (O_2787,N_24590,N_24652);
nor UO_2788 (O_2788,N_24651,N_24570);
and UO_2789 (O_2789,N_24138,N_24048);
nand UO_2790 (O_2790,N_24637,N_24587);
and UO_2791 (O_2791,N_24690,N_24720);
and UO_2792 (O_2792,N_24099,N_24762);
xnor UO_2793 (O_2793,N_24015,N_24640);
xnor UO_2794 (O_2794,N_24782,N_24025);
nor UO_2795 (O_2795,N_24245,N_24863);
nand UO_2796 (O_2796,N_24960,N_24620);
nand UO_2797 (O_2797,N_24803,N_24953);
nand UO_2798 (O_2798,N_24275,N_24753);
nand UO_2799 (O_2799,N_24024,N_24894);
nand UO_2800 (O_2800,N_24864,N_24799);
nor UO_2801 (O_2801,N_24163,N_24556);
nor UO_2802 (O_2802,N_24122,N_24809);
nand UO_2803 (O_2803,N_24108,N_24988);
xnor UO_2804 (O_2804,N_24414,N_24638);
and UO_2805 (O_2805,N_24507,N_24298);
or UO_2806 (O_2806,N_24705,N_24721);
xor UO_2807 (O_2807,N_24390,N_24881);
xnor UO_2808 (O_2808,N_24767,N_24072);
nor UO_2809 (O_2809,N_24907,N_24891);
or UO_2810 (O_2810,N_24099,N_24606);
and UO_2811 (O_2811,N_24474,N_24659);
nor UO_2812 (O_2812,N_24532,N_24777);
xnor UO_2813 (O_2813,N_24674,N_24931);
nor UO_2814 (O_2814,N_24934,N_24453);
and UO_2815 (O_2815,N_24553,N_24486);
or UO_2816 (O_2816,N_24260,N_24853);
nand UO_2817 (O_2817,N_24110,N_24566);
nand UO_2818 (O_2818,N_24018,N_24637);
or UO_2819 (O_2819,N_24468,N_24773);
and UO_2820 (O_2820,N_24073,N_24775);
nand UO_2821 (O_2821,N_24770,N_24951);
nand UO_2822 (O_2822,N_24518,N_24340);
or UO_2823 (O_2823,N_24855,N_24913);
and UO_2824 (O_2824,N_24025,N_24728);
and UO_2825 (O_2825,N_24858,N_24593);
and UO_2826 (O_2826,N_24960,N_24031);
xor UO_2827 (O_2827,N_24594,N_24830);
nand UO_2828 (O_2828,N_24209,N_24488);
xnor UO_2829 (O_2829,N_24725,N_24623);
xnor UO_2830 (O_2830,N_24998,N_24155);
nor UO_2831 (O_2831,N_24562,N_24279);
nand UO_2832 (O_2832,N_24848,N_24922);
nor UO_2833 (O_2833,N_24262,N_24553);
nor UO_2834 (O_2834,N_24092,N_24813);
nand UO_2835 (O_2835,N_24481,N_24095);
xor UO_2836 (O_2836,N_24281,N_24444);
nand UO_2837 (O_2837,N_24735,N_24000);
and UO_2838 (O_2838,N_24744,N_24169);
nor UO_2839 (O_2839,N_24608,N_24079);
nand UO_2840 (O_2840,N_24821,N_24793);
and UO_2841 (O_2841,N_24737,N_24411);
and UO_2842 (O_2842,N_24313,N_24706);
and UO_2843 (O_2843,N_24818,N_24531);
nor UO_2844 (O_2844,N_24517,N_24071);
nand UO_2845 (O_2845,N_24781,N_24149);
nand UO_2846 (O_2846,N_24231,N_24298);
and UO_2847 (O_2847,N_24504,N_24314);
or UO_2848 (O_2848,N_24436,N_24981);
xor UO_2849 (O_2849,N_24062,N_24304);
nand UO_2850 (O_2850,N_24196,N_24388);
xnor UO_2851 (O_2851,N_24989,N_24080);
xor UO_2852 (O_2852,N_24535,N_24002);
nand UO_2853 (O_2853,N_24751,N_24578);
nand UO_2854 (O_2854,N_24379,N_24657);
nand UO_2855 (O_2855,N_24335,N_24916);
xor UO_2856 (O_2856,N_24544,N_24932);
nand UO_2857 (O_2857,N_24110,N_24797);
nor UO_2858 (O_2858,N_24858,N_24675);
nand UO_2859 (O_2859,N_24249,N_24587);
nand UO_2860 (O_2860,N_24203,N_24196);
and UO_2861 (O_2861,N_24761,N_24015);
and UO_2862 (O_2862,N_24783,N_24357);
and UO_2863 (O_2863,N_24707,N_24159);
or UO_2864 (O_2864,N_24511,N_24753);
nand UO_2865 (O_2865,N_24515,N_24007);
xor UO_2866 (O_2866,N_24874,N_24517);
nor UO_2867 (O_2867,N_24364,N_24532);
and UO_2868 (O_2868,N_24972,N_24727);
nand UO_2869 (O_2869,N_24016,N_24397);
nand UO_2870 (O_2870,N_24621,N_24343);
nor UO_2871 (O_2871,N_24586,N_24215);
and UO_2872 (O_2872,N_24480,N_24865);
xor UO_2873 (O_2873,N_24796,N_24177);
xnor UO_2874 (O_2874,N_24857,N_24547);
and UO_2875 (O_2875,N_24345,N_24449);
or UO_2876 (O_2876,N_24840,N_24055);
or UO_2877 (O_2877,N_24072,N_24379);
and UO_2878 (O_2878,N_24949,N_24722);
or UO_2879 (O_2879,N_24466,N_24678);
xor UO_2880 (O_2880,N_24874,N_24365);
xor UO_2881 (O_2881,N_24306,N_24724);
or UO_2882 (O_2882,N_24415,N_24162);
xor UO_2883 (O_2883,N_24572,N_24828);
nor UO_2884 (O_2884,N_24312,N_24070);
xor UO_2885 (O_2885,N_24661,N_24914);
and UO_2886 (O_2886,N_24241,N_24515);
and UO_2887 (O_2887,N_24218,N_24344);
or UO_2888 (O_2888,N_24373,N_24921);
xnor UO_2889 (O_2889,N_24040,N_24711);
and UO_2890 (O_2890,N_24294,N_24236);
xor UO_2891 (O_2891,N_24767,N_24610);
nor UO_2892 (O_2892,N_24951,N_24012);
nand UO_2893 (O_2893,N_24002,N_24232);
or UO_2894 (O_2894,N_24261,N_24558);
or UO_2895 (O_2895,N_24837,N_24265);
nand UO_2896 (O_2896,N_24630,N_24682);
and UO_2897 (O_2897,N_24295,N_24438);
nand UO_2898 (O_2898,N_24302,N_24626);
nor UO_2899 (O_2899,N_24618,N_24230);
and UO_2900 (O_2900,N_24615,N_24064);
and UO_2901 (O_2901,N_24349,N_24929);
nand UO_2902 (O_2902,N_24160,N_24570);
and UO_2903 (O_2903,N_24319,N_24056);
nor UO_2904 (O_2904,N_24027,N_24431);
nor UO_2905 (O_2905,N_24444,N_24432);
or UO_2906 (O_2906,N_24623,N_24898);
and UO_2907 (O_2907,N_24518,N_24654);
and UO_2908 (O_2908,N_24577,N_24495);
nor UO_2909 (O_2909,N_24969,N_24417);
and UO_2910 (O_2910,N_24242,N_24817);
nand UO_2911 (O_2911,N_24550,N_24088);
nand UO_2912 (O_2912,N_24212,N_24958);
xor UO_2913 (O_2913,N_24293,N_24781);
nor UO_2914 (O_2914,N_24546,N_24065);
or UO_2915 (O_2915,N_24230,N_24080);
nor UO_2916 (O_2916,N_24787,N_24321);
and UO_2917 (O_2917,N_24252,N_24036);
nor UO_2918 (O_2918,N_24023,N_24449);
nand UO_2919 (O_2919,N_24425,N_24463);
nor UO_2920 (O_2920,N_24084,N_24186);
xor UO_2921 (O_2921,N_24087,N_24191);
xnor UO_2922 (O_2922,N_24414,N_24483);
nand UO_2923 (O_2923,N_24670,N_24028);
nand UO_2924 (O_2924,N_24071,N_24131);
or UO_2925 (O_2925,N_24724,N_24979);
xor UO_2926 (O_2926,N_24458,N_24542);
nor UO_2927 (O_2927,N_24071,N_24224);
nand UO_2928 (O_2928,N_24981,N_24464);
and UO_2929 (O_2929,N_24323,N_24812);
nor UO_2930 (O_2930,N_24682,N_24925);
xor UO_2931 (O_2931,N_24189,N_24207);
and UO_2932 (O_2932,N_24617,N_24553);
and UO_2933 (O_2933,N_24726,N_24126);
nor UO_2934 (O_2934,N_24363,N_24529);
nand UO_2935 (O_2935,N_24401,N_24141);
nor UO_2936 (O_2936,N_24295,N_24198);
and UO_2937 (O_2937,N_24602,N_24912);
nor UO_2938 (O_2938,N_24581,N_24941);
xor UO_2939 (O_2939,N_24629,N_24595);
xnor UO_2940 (O_2940,N_24868,N_24104);
and UO_2941 (O_2941,N_24704,N_24947);
nor UO_2942 (O_2942,N_24449,N_24900);
xnor UO_2943 (O_2943,N_24696,N_24789);
xor UO_2944 (O_2944,N_24711,N_24962);
nand UO_2945 (O_2945,N_24977,N_24938);
nor UO_2946 (O_2946,N_24734,N_24837);
nand UO_2947 (O_2947,N_24974,N_24869);
and UO_2948 (O_2948,N_24042,N_24684);
xor UO_2949 (O_2949,N_24493,N_24833);
nand UO_2950 (O_2950,N_24087,N_24097);
nand UO_2951 (O_2951,N_24869,N_24266);
and UO_2952 (O_2952,N_24922,N_24706);
nor UO_2953 (O_2953,N_24104,N_24696);
nor UO_2954 (O_2954,N_24403,N_24130);
and UO_2955 (O_2955,N_24228,N_24838);
and UO_2956 (O_2956,N_24969,N_24810);
nor UO_2957 (O_2957,N_24302,N_24991);
or UO_2958 (O_2958,N_24234,N_24217);
nor UO_2959 (O_2959,N_24741,N_24368);
nand UO_2960 (O_2960,N_24845,N_24391);
and UO_2961 (O_2961,N_24535,N_24148);
nand UO_2962 (O_2962,N_24267,N_24071);
xnor UO_2963 (O_2963,N_24739,N_24770);
nand UO_2964 (O_2964,N_24880,N_24007);
nor UO_2965 (O_2965,N_24839,N_24471);
xnor UO_2966 (O_2966,N_24736,N_24337);
nand UO_2967 (O_2967,N_24536,N_24902);
nand UO_2968 (O_2968,N_24689,N_24447);
and UO_2969 (O_2969,N_24910,N_24870);
and UO_2970 (O_2970,N_24496,N_24779);
nor UO_2971 (O_2971,N_24309,N_24003);
and UO_2972 (O_2972,N_24742,N_24057);
xor UO_2973 (O_2973,N_24251,N_24566);
or UO_2974 (O_2974,N_24886,N_24462);
and UO_2975 (O_2975,N_24140,N_24523);
nor UO_2976 (O_2976,N_24131,N_24233);
nor UO_2977 (O_2977,N_24416,N_24738);
nor UO_2978 (O_2978,N_24671,N_24041);
nand UO_2979 (O_2979,N_24291,N_24684);
nand UO_2980 (O_2980,N_24801,N_24492);
or UO_2981 (O_2981,N_24729,N_24237);
or UO_2982 (O_2982,N_24736,N_24594);
or UO_2983 (O_2983,N_24423,N_24488);
and UO_2984 (O_2984,N_24583,N_24500);
xor UO_2985 (O_2985,N_24448,N_24465);
nand UO_2986 (O_2986,N_24562,N_24084);
nand UO_2987 (O_2987,N_24368,N_24220);
nor UO_2988 (O_2988,N_24111,N_24879);
or UO_2989 (O_2989,N_24690,N_24724);
nand UO_2990 (O_2990,N_24033,N_24128);
nor UO_2991 (O_2991,N_24105,N_24925);
xor UO_2992 (O_2992,N_24908,N_24283);
and UO_2993 (O_2993,N_24713,N_24041);
xnor UO_2994 (O_2994,N_24318,N_24168);
xor UO_2995 (O_2995,N_24862,N_24995);
xor UO_2996 (O_2996,N_24279,N_24382);
nand UO_2997 (O_2997,N_24906,N_24898);
or UO_2998 (O_2998,N_24150,N_24584);
xor UO_2999 (O_2999,N_24664,N_24109);
endmodule