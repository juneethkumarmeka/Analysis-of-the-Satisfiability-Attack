module basic_1500_15000_2000_30_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_366,In_1386);
nor U1 (N_1,In_539,In_1406);
or U2 (N_2,In_267,In_578);
nor U3 (N_3,In_873,In_1366);
and U4 (N_4,In_494,In_641);
xnor U5 (N_5,In_989,In_497);
or U6 (N_6,In_67,In_1216);
and U7 (N_7,In_848,In_14);
and U8 (N_8,In_753,In_1427);
nand U9 (N_9,In_713,In_1293);
nand U10 (N_10,In_281,In_1270);
nor U11 (N_11,In_106,In_581);
nor U12 (N_12,In_414,In_583);
or U13 (N_13,In_918,In_969);
nand U14 (N_14,In_948,In_1394);
or U15 (N_15,In_1391,In_13);
xnor U16 (N_16,In_280,In_464);
nand U17 (N_17,In_483,In_1222);
and U18 (N_18,In_1136,In_1428);
nand U19 (N_19,In_1365,In_1496);
xnor U20 (N_20,In_1200,In_1237);
nor U21 (N_21,In_580,In_1435);
and U22 (N_22,In_1350,In_812);
nor U23 (N_23,In_566,In_284);
nand U24 (N_24,In_800,In_37);
nor U25 (N_25,In_248,In_777);
nor U26 (N_26,In_41,In_1129);
and U27 (N_27,In_355,In_134);
nor U28 (N_28,In_731,In_1148);
nor U29 (N_29,In_639,In_339);
or U30 (N_30,In_43,In_1469);
or U31 (N_31,In_111,In_194);
or U32 (N_32,In_769,In_1158);
nand U33 (N_33,In_554,In_1460);
nand U34 (N_34,In_130,In_63);
nand U35 (N_35,In_18,In_147);
nand U36 (N_36,In_773,In_651);
nor U37 (N_37,In_1119,In_227);
and U38 (N_38,In_1034,In_775);
xnor U39 (N_39,In_412,In_276);
and U40 (N_40,In_335,In_1049);
or U41 (N_41,In_1240,In_20);
nand U42 (N_42,In_12,In_465);
nor U43 (N_43,In_850,In_27);
and U44 (N_44,In_653,In_505);
nor U45 (N_45,In_190,In_172);
nor U46 (N_46,In_277,In_616);
and U47 (N_47,In_923,In_1396);
nor U48 (N_48,In_84,In_1123);
and U49 (N_49,In_737,In_264);
nand U50 (N_50,In_1430,In_153);
nand U51 (N_51,In_1197,In_890);
nand U52 (N_52,In_99,In_480);
or U53 (N_53,In_1289,In_1264);
nor U54 (N_54,In_302,In_636);
and U55 (N_55,In_931,In_744);
and U56 (N_56,In_338,In_124);
nand U57 (N_57,In_760,In_1093);
nor U58 (N_58,In_495,In_1145);
or U59 (N_59,In_1392,In_169);
or U60 (N_60,In_1497,In_973);
xnor U61 (N_61,In_1111,In_656);
and U62 (N_62,In_1082,In_966);
and U63 (N_63,In_790,In_625);
or U64 (N_64,In_1384,In_678);
and U65 (N_65,In_997,In_741);
and U66 (N_66,In_897,In_1046);
and U67 (N_67,In_1141,In_121);
xnor U68 (N_68,In_60,In_1239);
xor U69 (N_69,In_21,In_176);
nor U70 (N_70,In_68,In_1190);
nand U71 (N_71,In_58,In_1055);
and U72 (N_72,In_1349,In_1387);
nor U73 (N_73,In_283,In_516);
and U74 (N_74,In_1195,In_1134);
or U75 (N_75,In_461,In_440);
or U76 (N_76,In_827,In_184);
and U77 (N_77,In_1268,In_584);
and U78 (N_78,In_1438,In_211);
xnor U79 (N_79,In_1498,In_1333);
xor U80 (N_80,In_714,In_186);
xnor U81 (N_81,In_1453,In_1328);
and U82 (N_82,In_39,In_1067);
xnor U83 (N_83,In_986,In_536);
xnor U84 (N_84,In_743,In_313);
nand U85 (N_85,In_449,In_1379);
and U86 (N_86,In_202,In_237);
and U87 (N_87,In_1159,In_23);
nor U88 (N_88,In_519,In_243);
and U89 (N_89,In_1398,In_1163);
nand U90 (N_90,In_1087,In_509);
nand U91 (N_91,In_562,In_1196);
nand U92 (N_92,In_1234,In_32);
nor U93 (N_93,In_331,In_950);
and U94 (N_94,In_633,In_1044);
and U95 (N_95,In_691,In_887);
xor U96 (N_96,In_472,In_368);
nand U97 (N_97,In_290,In_1370);
xnor U98 (N_98,In_357,In_683);
nand U99 (N_99,In_1362,In_165);
nand U100 (N_100,In_706,In_259);
and U101 (N_101,In_166,In_1079);
nand U102 (N_102,In_1088,In_537);
or U103 (N_103,In_650,In_1004);
nor U104 (N_104,In_821,In_1205);
nor U105 (N_105,In_928,In_927);
and U106 (N_106,In_780,In_847);
nand U107 (N_107,In_881,In_862);
nand U108 (N_108,In_385,In_363);
nor U109 (N_109,In_1250,In_967);
nor U110 (N_110,In_978,In_739);
or U111 (N_111,In_803,In_323);
nand U112 (N_112,In_1164,In_1201);
or U113 (N_113,In_1066,In_630);
and U114 (N_114,In_163,In_419);
nand U115 (N_115,In_1076,In_356);
and U116 (N_116,In_1098,In_858);
nand U117 (N_117,In_217,In_913);
and U118 (N_118,In_1336,In_611);
or U119 (N_119,In_7,In_299);
nand U120 (N_120,In_126,In_1363);
xor U121 (N_121,In_100,In_643);
nand U122 (N_122,In_1120,In_1375);
nor U123 (N_123,In_1285,In_1083);
nand U124 (N_124,In_224,In_136);
nor U125 (N_125,In_514,In_1221);
and U126 (N_126,In_1419,In_960);
nor U127 (N_127,In_1426,In_1227);
nor U128 (N_128,In_1086,In_535);
and U129 (N_129,In_486,In_30);
nand U130 (N_130,In_961,In_24);
and U131 (N_131,In_1053,In_1484);
nor U132 (N_132,In_628,In_1059);
nor U133 (N_133,In_994,In_1332);
nor U134 (N_134,In_957,In_1476);
nand U135 (N_135,In_369,In_1130);
and U136 (N_136,In_1133,In_332);
or U137 (N_137,In_851,In_1191);
or U138 (N_138,In_689,In_496);
xnor U139 (N_139,In_674,In_298);
nand U140 (N_140,In_151,In_146);
xor U141 (N_141,In_1425,In_820);
and U142 (N_142,In_1184,In_159);
nand U143 (N_143,In_1395,In_1211);
nor U144 (N_144,In_622,In_155);
nand U145 (N_145,In_1071,In_1016);
or U146 (N_146,In_1327,In_262);
xor U147 (N_147,In_188,In_833);
nand U148 (N_148,In_665,In_105);
and U149 (N_149,In_474,In_345);
and U150 (N_150,In_1179,In_1260);
or U151 (N_151,In_1321,In_326);
nand U152 (N_152,In_1272,In_52);
or U153 (N_153,In_836,In_1238);
and U154 (N_154,In_877,In_813);
and U155 (N_155,In_1443,In_142);
nor U156 (N_156,In_373,In_1152);
nor U157 (N_157,In_1137,In_108);
nor U158 (N_158,In_922,In_123);
nand U159 (N_159,In_1143,In_422);
and U160 (N_160,In_96,In_854);
nand U161 (N_161,In_878,In_1251);
nor U162 (N_162,In_909,In_98);
and U163 (N_163,In_1045,In_990);
or U164 (N_164,In_500,In_866);
nand U165 (N_165,In_576,In_874);
xnor U166 (N_166,In_179,In_503);
or U167 (N_167,In_160,In_132);
or U168 (N_168,In_291,In_1029);
or U169 (N_169,In_1024,In_1009);
and U170 (N_170,In_102,In_45);
and U171 (N_171,In_1275,In_863);
and U172 (N_172,In_1372,In_307);
nand U173 (N_173,In_1356,In_38);
nand U174 (N_174,In_1019,In_1403);
or U175 (N_175,In_1,In_941);
nor U176 (N_176,In_9,In_839);
xor U177 (N_177,In_1236,In_158);
nand U178 (N_178,In_387,In_430);
or U179 (N_179,In_735,In_64);
and U180 (N_180,In_508,In_1175);
and U181 (N_181,In_220,In_205);
or U182 (N_182,In_1465,In_1310);
nor U183 (N_183,In_256,In_1431);
and U184 (N_184,In_216,In_545);
nand U185 (N_185,In_46,In_1106);
or U186 (N_186,In_1373,In_548);
nor U187 (N_187,In_551,In_1005);
nand U188 (N_188,In_1172,In_6);
or U189 (N_189,In_620,In_646);
nor U190 (N_190,In_996,In_411);
and U191 (N_191,In_955,In_1099);
nor U192 (N_192,In_547,In_517);
nor U193 (N_193,In_1353,In_1292);
or U194 (N_194,In_1116,In_1153);
nand U195 (N_195,In_1262,In_1338);
xor U196 (N_196,In_62,In_502);
nor U197 (N_197,In_171,In_959);
nand U198 (N_198,In_306,In_914);
and U199 (N_199,In_384,In_565);
or U200 (N_200,In_214,In_1344);
nand U201 (N_201,In_606,In_445);
nand U202 (N_202,In_249,In_1015);
and U203 (N_203,In_784,In_415);
nand U204 (N_204,In_1080,In_33);
nor U205 (N_205,In_203,In_358);
or U206 (N_206,In_327,In_571);
nand U207 (N_207,In_676,In_705);
nand U208 (N_208,In_1173,In_1467);
nand U209 (N_209,In_1499,In_316);
and U210 (N_210,In_658,In_448);
nand U211 (N_211,In_1092,In_561);
or U212 (N_212,In_785,In_1452);
or U213 (N_213,In_175,In_1343);
nand U214 (N_214,In_399,In_530);
nand U215 (N_215,In_1400,In_1008);
xnor U216 (N_216,In_15,In_1471);
nand U217 (N_217,In_498,In_1223);
xnor U218 (N_218,In_844,In_882);
nand U219 (N_219,In_441,In_772);
xnor U220 (N_220,In_680,In_843);
or U221 (N_221,In_1101,In_1454);
xnor U222 (N_222,In_76,In_886);
and U223 (N_223,In_1423,In_869);
xnor U224 (N_224,In_44,In_193);
nor U225 (N_225,In_804,In_1481);
and U226 (N_226,In_392,In_860);
or U227 (N_227,In_1209,In_1369);
and U228 (N_228,In_1485,In_888);
and U229 (N_229,In_282,In_1410);
nand U230 (N_230,In_1028,In_402);
nand U231 (N_231,In_574,In_1269);
nand U232 (N_232,In_215,In_1219);
nor U233 (N_233,In_234,In_1048);
nand U234 (N_234,In_1036,In_670);
or U235 (N_235,In_1448,In_788);
nor U236 (N_236,In_1204,In_943);
and U237 (N_237,In_150,In_688);
nand U238 (N_238,In_25,In_437);
or U239 (N_239,In_1188,In_1255);
nor U240 (N_240,In_428,In_1376);
nand U241 (N_241,In_1382,In_22);
or U242 (N_242,In_638,In_810);
nand U243 (N_243,In_991,In_607);
or U244 (N_244,In_1266,In_479);
and U245 (N_245,In_1472,In_1060);
and U246 (N_246,In_1249,In_374);
nand U247 (N_247,In_673,In_1156);
and U248 (N_248,In_720,In_1091);
nor U249 (N_249,In_1458,In_917);
and U250 (N_250,In_138,In_92);
or U251 (N_251,In_1078,In_418);
and U252 (N_252,In_183,In_1037);
nand U253 (N_253,In_1155,In_783);
and U254 (N_254,In_522,In_1302);
nor U255 (N_255,In_72,In_912);
nor U256 (N_256,In_1303,In_329);
nand U257 (N_257,In_1324,In_431);
and U258 (N_258,In_585,In_86);
nand U259 (N_259,In_701,In_868);
xnor U260 (N_260,In_493,In_1432);
or U261 (N_261,In_453,In_1062);
or U262 (N_262,In_975,In_1478);
nor U263 (N_263,In_5,In_849);
nor U264 (N_264,In_1243,In_454);
nor U265 (N_265,In_478,In_781);
and U266 (N_266,In_352,In_1287);
nand U267 (N_267,In_1113,In_225);
nand U268 (N_268,In_178,In_786);
nor U269 (N_269,In_792,In_655);
nor U270 (N_270,In_1335,In_507);
or U271 (N_271,In_61,In_1107);
and U272 (N_272,In_322,In_1011);
xnor U273 (N_273,In_1385,In_1466);
or U274 (N_274,In_239,In_1315);
nor U275 (N_275,In_1026,In_1169);
or U276 (N_276,In_349,In_162);
and U277 (N_277,In_1215,In_1377);
nand U278 (N_278,In_1199,In_310);
nand U279 (N_279,In_900,In_702);
nand U280 (N_280,In_80,In_938);
nand U281 (N_281,In_778,In_117);
nand U282 (N_282,In_779,In_1487);
and U283 (N_283,In_1494,In_312);
nand U284 (N_284,In_654,In_1002);
nand U285 (N_285,In_1124,In_1105);
nor U286 (N_286,In_391,In_588);
or U287 (N_287,In_816,In_1288);
xnor U288 (N_288,In_956,In_0);
nand U289 (N_289,In_1323,In_1118);
nand U290 (N_290,In_409,In_755);
or U291 (N_291,In_919,In_1388);
nor U292 (N_292,In_663,In_1341);
nor U293 (N_293,In_894,In_533);
or U294 (N_294,In_181,In_1281);
nor U295 (N_295,In_808,In_1065);
nor U296 (N_296,In_254,In_1380);
or U297 (N_297,In_1461,In_1254);
nor U298 (N_298,In_1397,In_1267);
xor U299 (N_299,In_269,In_697);
nor U300 (N_300,In_748,In_838);
xor U301 (N_301,In_470,In_73);
nor U302 (N_302,In_1296,In_793);
nand U303 (N_303,In_343,In_852);
xnor U304 (N_304,In_1308,In_936);
and U305 (N_305,In_149,In_623);
or U306 (N_306,In_71,In_528);
nand U307 (N_307,In_1056,In_311);
nand U308 (N_308,In_1127,In_504);
or U309 (N_309,In_542,In_4);
nand U310 (N_310,In_634,In_1299);
or U311 (N_311,In_807,In_1300);
nor U312 (N_312,In_946,In_114);
or U313 (N_313,In_424,In_811);
and U314 (N_314,In_1473,In_1439);
nand U315 (N_315,In_1334,In_1003);
and U316 (N_316,In_795,In_93);
nand U317 (N_317,In_597,In_605);
nor U318 (N_318,In_529,In_1374);
nand U319 (N_319,In_1168,In_515);
and U320 (N_320,In_1450,In_756);
nand U321 (N_321,In_766,In_196);
or U322 (N_322,In_579,In_148);
nand U323 (N_323,In_856,In_935);
nand U324 (N_324,In_1351,In_635);
nor U325 (N_325,In_1245,In_671);
and U326 (N_326,In_1446,In_31);
nand U327 (N_327,In_139,In_1241);
or U328 (N_328,In_1486,In_118);
and U329 (N_329,In_1418,In_563);
xor U330 (N_330,In_246,In_288);
or U331 (N_331,In_1089,In_698);
nor U332 (N_332,In_1265,In_722);
xor U333 (N_333,In_586,In_905);
xor U334 (N_334,In_1140,In_416);
nand U335 (N_335,In_295,In_1283);
nand U336 (N_336,In_1279,In_704);
nor U337 (N_337,In_686,In_1000);
or U338 (N_338,In_921,In_980);
or U339 (N_339,In_1007,In_443);
and U340 (N_340,In_727,In_1198);
nand U341 (N_341,In_573,In_28);
nand U342 (N_342,In_947,In_893);
nand U343 (N_343,In_212,In_1231);
and U344 (N_344,In_932,In_1035);
or U345 (N_345,In_244,In_324);
or U346 (N_346,In_279,In_988);
xor U347 (N_347,In_1462,In_265);
nor U348 (N_348,In_53,In_724);
nor U349 (N_349,In_1025,In_487);
xor U350 (N_350,In_898,In_253);
nor U351 (N_351,In_1412,In_608);
and U352 (N_352,In_594,In_687);
and U353 (N_353,In_593,In_1447);
or U354 (N_354,In_83,In_774);
and U355 (N_355,In_377,In_910);
and U356 (N_356,In_1006,In_518);
or U357 (N_357,In_222,In_1354);
and U358 (N_358,In_589,In_26);
and U359 (N_359,In_1437,In_666);
nor U360 (N_360,In_1154,In_29);
and U361 (N_361,In_1210,In_815);
and U362 (N_362,In_119,In_1135);
or U363 (N_363,In_1167,In_541);
nor U364 (N_364,In_1075,In_524);
xor U365 (N_365,In_152,In_1381);
nor U366 (N_366,In_341,In_995);
xor U367 (N_367,In_1138,In_328);
nand U368 (N_368,In_830,In_235);
nor U369 (N_369,In_278,In_632);
and U370 (N_370,In_40,In_426);
xnor U371 (N_371,In_1208,In_1187);
and U372 (N_372,In_477,In_1110);
or U373 (N_373,In_91,In_682);
nand U374 (N_374,In_1063,In_1160);
and U375 (N_375,In_458,In_168);
or U376 (N_376,In_447,In_1407);
and U377 (N_377,In_1177,In_1401);
nand U378 (N_378,In_1217,In_285);
nand U379 (N_379,In_49,In_1073);
or U380 (N_380,In_703,In_1235);
nand U381 (N_381,In_768,In_110);
nand U382 (N_382,In_457,In_1102);
and U383 (N_383,In_765,In_915);
xnor U384 (N_384,In_1166,In_393);
nor U385 (N_385,In_195,In_317);
nand U386 (N_386,In_557,In_835);
or U387 (N_387,In_817,In_297);
nand U388 (N_388,In_1298,In_746);
or U389 (N_389,In_1339,In_81);
xnor U390 (N_390,In_116,In_1125);
and U391 (N_391,In_143,In_1314);
nand U392 (N_392,In_271,In_734);
and U393 (N_393,In_717,In_885);
nor U394 (N_394,In_1017,In_1284);
or U395 (N_395,In_174,In_823);
or U396 (N_396,In_379,In_1345);
or U397 (N_397,In_1174,In_675);
nand U398 (N_398,In_97,In_491);
nand U399 (N_399,In_1475,In_925);
nor U400 (N_400,In_526,In_1474);
or U401 (N_401,In_1393,In_274);
or U402 (N_402,In_490,In_207);
nor U403 (N_403,In_1072,In_140);
and U404 (N_404,In_340,In_875);
nand U405 (N_405,In_962,In_315);
and U406 (N_406,In_273,In_221);
or U407 (N_407,In_423,In_953);
and U408 (N_408,In_672,In_789);
xnor U409 (N_409,In_161,In_709);
xor U410 (N_410,In_857,In_135);
or U411 (N_411,In_841,In_388);
xor U412 (N_412,In_1202,In_564);
nor U413 (N_413,In_1309,In_104);
xor U414 (N_414,In_1378,In_1018);
nand U415 (N_415,In_871,In_467);
nand U416 (N_416,In_1420,In_1352);
or U417 (N_417,In_745,In_1305);
nand U418 (N_418,In_602,In_19);
nor U419 (N_419,In_79,In_964);
and U420 (N_420,In_1207,In_372);
and U421 (N_421,In_1399,In_1429);
nor U422 (N_422,In_1280,In_371);
nand U423 (N_423,In_627,In_644);
nor U424 (N_424,In_204,In_952);
or U425 (N_425,In_1258,In_657);
or U426 (N_426,In_587,In_747);
nand U427 (N_427,In_164,In_570);
or U428 (N_428,In_907,In_436);
or U429 (N_429,In_1041,In_1340);
nor U430 (N_430,In_506,In_1117);
or U431 (N_431,In_879,In_1490);
nor U432 (N_432,In_558,In_305);
and U433 (N_433,In_837,In_1242);
nor U434 (N_434,In_361,In_982);
or U435 (N_435,In_1390,In_951);
nor U436 (N_436,In_78,In_934);
nand U437 (N_437,In_365,In_407);
nor U438 (N_438,In_617,In_1347);
or U439 (N_439,In_325,In_442);
or U440 (N_440,In_476,In_1033);
and U441 (N_441,In_382,In_668);
or U442 (N_442,In_353,In_1330);
and U443 (N_443,In_473,In_799);
xnor U444 (N_444,In_95,In_1278);
and U445 (N_445,In_1449,In_754);
or U446 (N_446,In_69,In_275);
nand U447 (N_447,In_434,In_1212);
nor U448 (N_448,In_65,In_296);
or U449 (N_449,In_82,In_595);
or U450 (N_450,In_1263,In_1109);
or U451 (N_451,In_301,In_263);
nor U452 (N_452,In_1477,In_1480);
nand U453 (N_453,In_742,In_845);
or U454 (N_454,In_8,In_74);
or U455 (N_455,In_895,In_814);
and U456 (N_456,In_109,In_1442);
nor U457 (N_457,In_694,In_603);
or U458 (N_458,In_75,In_201);
nand U459 (N_459,In_1455,In_336);
or U460 (N_460,In_1357,In_872);
and U461 (N_461,In_1367,In_85);
and U462 (N_462,In_131,In_386);
nand U463 (N_463,In_420,In_719);
xnor U464 (N_464,In_621,In_930);
nor U465 (N_465,In_652,In_321);
xor U466 (N_466,In_958,In_218);
nor U467 (N_467,In_725,In_711);
nor U468 (N_468,In_1244,In_367);
and U469 (N_469,In_1220,In_805);
and U470 (N_470,In_1252,In_510);
nand U471 (N_471,In_1194,In_1189);
and U472 (N_472,In_1183,In_1050);
nor U473 (N_473,In_1013,In_197);
or U474 (N_474,In_1074,In_846);
or U475 (N_475,In_50,In_133);
and U476 (N_476,In_375,In_733);
and U477 (N_477,In_770,In_1213);
or U478 (N_478,In_729,In_47);
nand U479 (N_479,In_230,In_208);
xor U480 (N_480,In_427,In_1126);
and U481 (N_481,In_984,In_1364);
xnor U482 (N_482,In_681,In_113);
or U483 (N_483,In_405,In_1405);
nand U484 (N_484,In_42,In_1151);
nor U485 (N_485,In_1032,In_1273);
or U486 (N_486,In_1489,In_1061);
and U487 (N_487,In_1186,In_600);
xnor U488 (N_488,In_723,In_1146);
nor U489 (N_489,In_1318,In_1131);
or U490 (N_490,In_404,In_200);
nand U491 (N_491,In_289,In_1022);
and U492 (N_492,In_397,In_721);
nor U493 (N_493,In_1294,In_261);
and U494 (N_494,In_645,In_330);
xnor U495 (N_495,In_1317,In_776);
nand U496 (N_496,In_1224,In_834);
and U497 (N_497,In_591,In_693);
or U498 (N_498,In_572,In_210);
or U499 (N_499,In_185,In_699);
nand U500 (N_500,In_1361,In_1248);
xor U501 (N_501,N_173,N_401);
and U502 (N_502,N_359,In_1128);
or U503 (N_503,N_320,N_428);
nand U504 (N_504,N_160,N_431);
nand U505 (N_505,In_1147,In_255);
nor U506 (N_506,N_166,In_167);
and U507 (N_507,N_480,In_286);
nand U508 (N_508,N_456,N_149);
xnor U509 (N_509,In_1274,In_767);
nand U510 (N_510,N_462,N_177);
or U511 (N_511,In_787,N_407);
and U512 (N_512,N_333,In_173);
and U513 (N_513,N_230,N_44);
nor U514 (N_514,N_260,N_22);
or U515 (N_515,N_198,In_145);
nand U516 (N_516,In_156,In_1114);
and U517 (N_517,N_229,N_78);
nor U518 (N_518,N_50,N_358);
and U519 (N_519,N_337,N_385);
nor U520 (N_520,N_301,In_822);
nand U521 (N_521,In_400,In_180);
nor U522 (N_522,N_188,N_305);
nand U523 (N_523,In_867,N_38);
xnor U524 (N_524,N_450,In_684);
or U525 (N_525,N_352,N_444);
and U526 (N_526,In_1492,In_413);
nor U527 (N_527,In_199,In_141);
and U528 (N_528,In_107,N_317);
or U529 (N_529,N_53,N_481);
or U530 (N_530,N_473,In_48);
or U531 (N_531,In_1256,In_718);
or U532 (N_532,N_41,N_242);
and U533 (N_533,In_1306,In_451);
nand U534 (N_534,In_446,In_1014);
and U535 (N_535,N_79,N_186);
nor U536 (N_536,N_219,N_75);
and U537 (N_537,In_751,In_891);
or U538 (N_538,In_738,N_414);
or U539 (N_539,In_1290,N_483);
nand U540 (N_540,N_277,N_471);
nand U541 (N_541,N_263,In_206);
nor U542 (N_542,N_310,In_127);
or U543 (N_543,In_859,In_1132);
nor U544 (N_544,N_421,In_304);
nand U545 (N_545,In_582,In_462);
nand U546 (N_546,In_347,In_791);
nand U547 (N_547,In_937,In_806);
nor U548 (N_548,In_56,In_553);
nand U549 (N_549,In_944,N_280);
nor U550 (N_550,In_540,In_1316);
or U551 (N_551,N_101,N_218);
nor U552 (N_552,N_128,In_626);
and U553 (N_553,N_60,In_381);
and U554 (N_554,In_89,In_1371);
and U555 (N_555,In_242,N_486);
or U556 (N_556,In_115,N_9);
nand U557 (N_557,N_429,N_410);
and U558 (N_558,N_196,N_49);
xor U559 (N_559,In_899,N_304);
nand U560 (N_560,N_457,In_940);
nor U561 (N_561,In_924,In_1043);
nand U562 (N_562,In_631,N_490);
or U563 (N_563,N_90,N_353);
and U564 (N_564,N_375,In_764);
and U565 (N_565,In_1445,In_122);
and U566 (N_566,N_30,In_695);
nor U567 (N_567,N_268,In_300);
nand U568 (N_568,N_382,In_1456);
or U569 (N_569,N_356,N_228);
nand U570 (N_570,In_1482,In_1112);
nor U571 (N_571,In_942,N_118);
xor U572 (N_572,In_308,In_998);
nand U573 (N_573,N_154,In_520);
nand U574 (N_574,In_883,In_247);
nand U575 (N_575,In_1096,In_1144);
and U576 (N_576,N_485,In_459);
or U577 (N_577,In_999,N_412);
or U578 (N_578,N_281,N_430);
or U579 (N_579,N_487,In_170);
or U580 (N_580,In_1483,In_527);
nand U581 (N_581,N_283,In_534);
nand U582 (N_582,In_55,In_360);
or U583 (N_583,N_35,In_752);
or U584 (N_584,In_485,In_272);
xnor U585 (N_585,In_292,In_1348);
or U586 (N_586,N_124,N_54);
and U587 (N_587,In_1170,In_992);
nand U588 (N_588,N_138,In_842);
and U589 (N_589,In_260,In_469);
nor U590 (N_590,In_1360,N_134);
nand U591 (N_591,N_86,N_8);
nor U592 (N_592,In_389,In_1081);
or U593 (N_593,In_896,N_157);
nor U594 (N_594,N_147,In_1203);
and U595 (N_595,In_730,N_448);
or U596 (N_596,In_797,N_71);
nand U597 (N_597,In_824,In_1228);
nand U598 (N_598,In_1436,In_1261);
and U599 (N_599,In_1451,In_1054);
nand U600 (N_600,N_14,In_1085);
nand U601 (N_601,N_459,N_491);
nor U602 (N_602,In_511,In_612);
nor U603 (N_603,N_59,N_387);
xor U604 (N_604,In_710,N_18);
nor U605 (N_605,N_74,N_461);
or U606 (N_606,N_111,In_649);
or U607 (N_607,In_1185,N_241);
or U608 (N_608,N_210,N_390);
and U609 (N_609,N_66,N_318);
nor U610 (N_610,In_1493,In_1149);
or U611 (N_611,In_1021,N_326);
or U612 (N_612,In_901,In_383);
nor U613 (N_613,In_592,N_419);
nand U614 (N_614,In_1441,N_64);
xor U615 (N_615,N_298,N_307);
or U616 (N_616,In_1408,In_1181);
nand U617 (N_617,In_549,N_131);
or U618 (N_618,N_165,In_88);
or U619 (N_619,N_5,N_357);
xnor U620 (N_620,In_1039,In_1020);
and U621 (N_621,In_1417,N_181);
and U622 (N_622,In_1470,N_161);
nor U623 (N_623,N_201,N_142);
and U624 (N_624,N_164,In_1094);
or U625 (N_625,In_209,N_466);
xor U626 (N_626,N_32,In_906);
or U627 (N_627,In_1434,In_1047);
nor U628 (N_628,In_911,N_225);
nor U629 (N_629,N_266,N_293);
or U630 (N_630,In_902,N_389);
nand U631 (N_631,In_1301,N_1);
and U632 (N_632,In_359,N_87);
or U633 (N_633,N_303,In_319);
or U634 (N_634,N_411,In_855);
nand U635 (N_635,N_383,In_1307);
and U636 (N_636,In_354,N_496);
nand U637 (N_637,N_208,In_1421);
and U638 (N_638,In_1468,N_395);
and U639 (N_639,In_112,N_339);
nor U640 (N_640,N_99,N_51);
or U641 (N_641,N_309,In_559);
and U642 (N_642,N_184,In_1052);
and U643 (N_643,In_560,In_433);
nor U644 (N_644,In_240,N_61);
and U645 (N_645,In_521,In_864);
nor U646 (N_646,In_1295,In_604);
xor U647 (N_647,N_68,N_91);
or U648 (N_648,N_296,In_908);
xor U649 (N_649,In_761,N_234);
and U650 (N_650,In_685,In_456);
or U651 (N_651,N_122,In_970);
nand U652 (N_652,In_137,In_829);
nand U653 (N_653,N_438,In_1226);
or U654 (N_654,In_1023,In_236);
nor U655 (N_655,N_341,N_29);
and U656 (N_656,N_209,N_469);
nand U657 (N_657,N_213,N_312);
xor U658 (N_658,In_87,In_763);
or U659 (N_659,N_299,In_1176);
and U660 (N_660,N_396,N_235);
nand U661 (N_661,In_629,In_1389);
nor U662 (N_662,N_117,N_158);
nand U663 (N_663,In_1042,In_241);
xor U664 (N_664,In_252,In_1368);
nor U665 (N_665,In_16,In_1414);
and U666 (N_666,N_278,N_191);
and U667 (N_667,N_350,N_152);
or U668 (N_668,In_1358,In_963);
and U669 (N_669,In_501,In_1491);
and U670 (N_670,N_474,In_749);
nand U671 (N_671,N_479,N_257);
nand U672 (N_672,N_329,N_493);
and U673 (N_673,N_16,In_376);
nor U674 (N_674,In_351,N_379);
nor U675 (N_675,In_1095,In_1097);
nand U676 (N_676,N_120,In_333);
nand U677 (N_677,In_1040,N_327);
nand U678 (N_678,N_216,In_590);
and U679 (N_679,In_1150,N_367);
or U680 (N_680,In_679,In_1319);
nor U681 (N_681,In_499,N_45);
or U682 (N_682,In_659,N_418);
and U683 (N_683,N_464,N_497);
xor U684 (N_684,N_351,In_1069);
xnor U685 (N_685,N_331,N_435);
and U686 (N_686,N_433,In_187);
nor U687 (N_687,N_273,In_342);
and U688 (N_688,N_370,In_1479);
xor U689 (N_689,In_1297,N_451);
nor U690 (N_690,In_661,In_266);
nand U691 (N_691,In_1277,N_193);
or U692 (N_692,N_100,N_338);
nand U693 (N_693,In_974,N_92);
xor U694 (N_694,N_300,In_492);
xor U695 (N_695,N_254,In_154);
nand U696 (N_696,In_11,In_1171);
nor U697 (N_697,In_613,In_1077);
or U698 (N_698,In_364,N_365);
nand U699 (N_699,In_771,N_70);
and U700 (N_700,In_831,N_222);
nand U701 (N_701,N_244,In_192);
nor U702 (N_702,In_1444,N_211);
nand U703 (N_703,N_476,In_801);
nor U704 (N_704,N_37,N_40);
or U705 (N_705,In_614,N_470);
or U706 (N_706,In_257,N_460);
nand U707 (N_707,In_667,N_88);
or U708 (N_708,N_27,N_46);
nor U709 (N_709,N_465,N_467);
nor U710 (N_710,N_34,In_696);
and U711 (N_711,N_494,In_976);
and U712 (N_712,In_450,N_33);
or U713 (N_713,In_294,In_926);
nor U714 (N_714,In_1058,N_102);
nor U715 (N_715,In_543,N_499);
nand U716 (N_716,In_1084,N_449);
nand U717 (N_717,In_884,In_17);
nor U718 (N_718,N_498,N_200);
nor U719 (N_719,N_139,In_189);
and U720 (N_720,N_97,In_826);
nand U721 (N_721,In_466,N_475);
nor U722 (N_722,N_250,N_290);
nor U723 (N_723,N_321,In_624);
xnor U724 (N_724,N_488,N_195);
nand U725 (N_725,In_344,In_213);
or U726 (N_726,N_25,In_700);
or U727 (N_727,N_306,In_1233);
nor U728 (N_728,In_1383,N_443);
and U729 (N_729,In_1192,N_406);
or U730 (N_730,In_482,N_439);
and U731 (N_731,N_287,N_17);
nand U732 (N_732,In_401,N_145);
nor U733 (N_733,In_226,N_183);
nand U734 (N_734,In_1090,In_619);
nor U735 (N_735,In_320,In_968);
or U736 (N_736,N_180,In_601);
nor U737 (N_737,In_832,N_361);
xor U738 (N_738,In_94,In_965);
xnor U739 (N_739,N_223,N_214);
nor U740 (N_740,In_1214,N_212);
or U741 (N_741,In_251,N_335);
or U742 (N_742,In_432,In_728);
or U743 (N_743,N_286,N_130);
nor U744 (N_744,N_322,In_1488);
and U745 (N_745,In_987,N_452);
nor U746 (N_746,In_1416,In_396);
nand U747 (N_747,In_223,N_324);
and U748 (N_748,In_429,In_1165);
and U749 (N_749,N_119,N_384);
nand U750 (N_750,In_303,N_292);
nor U751 (N_751,In_1031,In_362);
or U752 (N_752,In_1030,N_215);
nor U753 (N_753,In_1282,N_202);
or U754 (N_754,N_69,In_334);
nand U755 (N_755,N_77,N_282);
nand U756 (N_756,N_221,N_84);
nand U757 (N_757,In_468,N_116);
nand U758 (N_758,N_187,In_318);
nand U759 (N_759,In_1320,N_434);
or U760 (N_760,N_133,In_715);
nand U761 (N_761,In_103,In_1051);
nor U762 (N_762,N_252,N_56);
and U763 (N_763,N_472,In_1057);
nor U764 (N_764,N_239,N_238);
xnor U765 (N_765,N_295,N_82);
nor U766 (N_766,In_618,In_993);
and U767 (N_767,N_362,In_876);
nor U768 (N_768,N_12,In_1291);
and U769 (N_769,N_10,In_531);
or U770 (N_770,N_343,In_929);
and U771 (N_771,In_438,N_369);
nand U772 (N_772,N_143,N_397);
nand U773 (N_773,In_615,In_794);
nand U774 (N_774,In_1193,N_94);
and U775 (N_775,In_1286,In_408);
and U776 (N_776,N_403,N_484);
nor U777 (N_777,In_1322,In_1068);
nand U778 (N_778,N_141,In_523);
xor U779 (N_779,In_798,In_532);
nand U780 (N_780,N_114,In_395);
xor U781 (N_781,In_460,N_249);
xnor U782 (N_782,N_4,In_1271);
nor U783 (N_783,N_240,N_62);
or U784 (N_784,N_489,N_227);
nand U785 (N_785,N_192,In_1313);
and U786 (N_786,In_971,In_452);
and U787 (N_787,N_48,N_400);
nand U788 (N_788,In_762,In_640);
xor U789 (N_789,In_736,In_1457);
and U790 (N_790,In_35,N_39);
and U791 (N_791,N_265,N_394);
xnor U792 (N_792,In_609,N_168);
nor U793 (N_793,In_120,In_481);
or U794 (N_794,N_95,In_677);
and U795 (N_795,N_442,In_394);
or U796 (N_796,N_73,N_163);
nand U797 (N_797,In_933,N_126);
or U798 (N_798,In_569,N_347);
xor U799 (N_799,N_262,In_157);
and U800 (N_800,In_1422,In_1404);
and U801 (N_801,In_567,In_949);
nand U802 (N_802,N_104,In_406);
xnor U803 (N_803,N_85,N_372);
nor U804 (N_804,N_224,N_468);
xor U805 (N_805,N_174,In_707);
nor U806 (N_806,In_1312,N_336);
nor U807 (N_807,In_819,In_3);
nand U808 (N_808,N_386,N_80);
nor U809 (N_809,N_482,N_334);
nand U810 (N_810,N_441,N_360);
xnor U811 (N_811,In_1424,In_314);
nor U812 (N_812,In_421,N_194);
or U813 (N_813,N_248,N_388);
or U814 (N_814,In_90,In_544);
nand U815 (N_815,N_380,N_364);
nand U816 (N_816,In_1232,N_340);
and U817 (N_817,In_233,N_264);
xor U818 (N_818,N_288,N_376);
nand U819 (N_819,N_267,N_424);
nor U820 (N_820,N_115,In_1218);
nand U821 (N_821,In_648,In_1246);
nand U822 (N_822,In_920,In_268);
nand U823 (N_823,N_15,In_1459);
nand U824 (N_824,N_175,In_1206);
nand U825 (N_825,In_238,N_405);
or U826 (N_826,N_76,In_1104);
or U827 (N_827,In_1012,N_371);
nand U828 (N_828,N_398,In_1225);
nand U829 (N_829,In_1038,N_455);
xor U830 (N_830,N_189,In_475);
nor U831 (N_831,N_7,N_121);
and U832 (N_832,In_182,N_153);
xnor U833 (N_833,N_67,N_43);
and U834 (N_834,N_251,In_101);
nor U835 (N_835,In_1108,N_463);
and U836 (N_836,In_782,In_350);
or U837 (N_837,N_427,N_89);
or U838 (N_838,N_381,N_259);
nand U839 (N_839,In_662,N_349);
or U840 (N_840,In_979,In_34);
xor U841 (N_841,N_190,N_416);
nor U842 (N_842,In_861,N_374);
nor U843 (N_843,In_939,In_398);
nor U844 (N_844,In_1304,In_403);
xor U845 (N_845,In_1359,N_113);
xnor U846 (N_846,N_217,N_125);
or U847 (N_847,In_463,N_72);
or U848 (N_848,N_346,In_370);
xor U849 (N_849,In_439,In_1142);
or U850 (N_850,N_169,N_176);
and U851 (N_851,In_985,N_311);
nand U852 (N_852,N_492,N_19);
or U853 (N_853,In_865,N_368);
nor U854 (N_854,N_106,In_758);
nand U855 (N_855,N_247,N_447);
nor U856 (N_856,In_716,N_162);
nand U857 (N_857,N_129,N_477);
or U858 (N_858,In_1103,N_137);
and U859 (N_859,N_167,N_58);
and U860 (N_860,In_796,In_853);
and U861 (N_861,N_109,N_432);
nor U862 (N_862,In_828,N_96);
xor U863 (N_863,N_151,N_323);
nor U864 (N_864,N_171,N_185);
nand U865 (N_865,In_1409,In_1326);
or U866 (N_866,N_269,N_289);
nand U867 (N_867,In_596,In_1495);
or U868 (N_868,In_1180,N_253);
nand U869 (N_869,In_538,N_205);
or U870 (N_870,N_197,N_232);
or U871 (N_871,N_302,N_319);
or U872 (N_872,In_1276,N_172);
and U873 (N_873,N_425,In_669);
nand U874 (N_874,N_436,In_1070);
and U875 (N_875,N_13,N_373);
and U876 (N_876,In_1355,N_57);
nor U877 (N_877,N_156,N_123);
nand U878 (N_878,In_425,In_1257);
and U879 (N_879,N_36,N_108);
and U880 (N_880,In_1331,N_363);
nand U881 (N_881,In_802,In_552);
nand U882 (N_882,In_647,In_390);
or U883 (N_883,N_110,In_732);
xor U884 (N_884,N_0,In_219);
or U885 (N_885,In_1402,In_1346);
nor U886 (N_886,In_1413,In_692);
nor U887 (N_887,N_105,In_916);
or U888 (N_888,N_226,N_155);
nand U889 (N_889,In_740,N_42);
and U890 (N_890,N_11,In_977);
and U891 (N_891,In_577,N_243);
xor U892 (N_892,In_555,N_261);
nor U893 (N_893,N_140,In_2);
and U894 (N_894,In_818,N_245);
and U895 (N_895,In_250,N_355);
nor U896 (N_896,In_610,N_423);
or U897 (N_897,In_229,N_231);
nand U898 (N_898,N_103,N_344);
or U899 (N_899,In_489,In_125);
nor U900 (N_900,N_233,N_21);
or U901 (N_901,In_1229,In_245);
nor U902 (N_902,N_274,In_575);
nor U903 (N_903,In_726,In_1010);
nor U904 (N_904,In_1342,In_1122);
and U905 (N_905,N_415,In_972);
nand U906 (N_906,N_204,N_52);
nor U907 (N_907,In_1433,In_380);
nor U908 (N_908,In_840,N_24);
xor U909 (N_909,In_435,In_568);
or U910 (N_910,N_332,N_203);
xor U911 (N_911,N_399,In_1139);
or U912 (N_912,In_690,N_246);
xor U913 (N_913,In_1027,N_297);
nor U914 (N_914,N_255,N_279);
nand U915 (N_915,N_392,In_455);
nand U916 (N_916,N_144,N_345);
and U917 (N_917,In_1100,N_440);
xnor U918 (N_918,N_276,In_191);
nand U919 (N_919,N_270,In_198);
nor U920 (N_920,N_426,In_128);
or U921 (N_921,N_258,In_945);
nand U922 (N_922,In_410,N_236);
or U923 (N_923,In_954,N_458);
and U924 (N_924,N_377,In_484);
or U925 (N_925,N_3,In_59);
nand U926 (N_926,In_258,In_1325);
or U927 (N_927,N_98,In_77);
or U928 (N_928,N_275,In_642);
nor U929 (N_929,In_1259,N_348);
xor U930 (N_930,In_598,In_983);
nor U931 (N_931,N_178,In_1440);
and U932 (N_932,In_809,N_272);
and U933 (N_933,N_179,In_637);
or U934 (N_934,In_1411,N_393);
or U935 (N_935,N_284,N_132);
nor U936 (N_936,N_6,In_471);
or U937 (N_937,N_81,N_445);
and U938 (N_938,N_135,In_66);
or U939 (N_939,In_57,N_314);
and U940 (N_940,N_316,In_1337);
or U941 (N_941,In_546,In_129);
or U942 (N_942,N_313,N_206);
and U943 (N_943,In_232,In_757);
nor U944 (N_944,N_159,N_199);
or U945 (N_945,In_270,In_904);
and U946 (N_946,In_889,N_330);
or U947 (N_947,N_271,N_63);
nor U948 (N_948,N_107,N_182);
nand U949 (N_949,In_550,N_291);
nor U950 (N_950,N_285,In_880);
nor U951 (N_951,N_127,In_1115);
nor U952 (N_952,In_1253,In_1001);
and U953 (N_953,In_981,In_346);
and U954 (N_954,N_2,In_1230);
nand U955 (N_955,In_750,N_112);
nor U956 (N_956,N_294,In_287);
or U957 (N_957,N_454,N_354);
or U958 (N_958,In_1415,In_870);
xor U959 (N_959,N_446,In_54);
nor U960 (N_960,In_660,In_417);
xor U961 (N_961,N_408,In_664);
nor U962 (N_962,N_378,In_1064);
or U963 (N_963,N_495,N_83);
or U964 (N_964,N_150,N_366);
xor U965 (N_965,N_28,N_342);
or U966 (N_966,In_759,N_478);
and U967 (N_967,In_599,N_93);
nor U968 (N_968,In_1182,N_20);
nor U969 (N_969,In_1162,In_1464);
nor U970 (N_970,In_1247,In_513);
xor U971 (N_971,N_420,In_1157);
nand U972 (N_972,In_70,In_825);
or U973 (N_973,In_293,In_512);
or U974 (N_974,N_65,In_51);
nand U975 (N_975,In_10,N_220);
and U976 (N_976,N_404,In_144);
or U977 (N_977,N_55,N_422);
and U978 (N_978,N_325,N_315);
nand U979 (N_979,In_712,In_309);
nor U980 (N_980,N_409,N_136);
xor U981 (N_981,In_556,In_337);
nor U982 (N_982,In_488,In_892);
nand U983 (N_983,In_1463,In_903);
nor U984 (N_984,N_437,N_170);
nand U985 (N_985,N_148,N_207);
or U986 (N_986,N_31,N_308);
nor U987 (N_987,N_417,N_146);
or U988 (N_988,In_1311,In_378);
or U989 (N_989,N_256,In_708);
xor U990 (N_990,N_453,N_413);
or U991 (N_991,In_231,In_525);
and U992 (N_992,In_1121,In_177);
nor U993 (N_993,N_47,N_23);
xnor U994 (N_994,In_36,N_328);
nor U995 (N_995,In_348,In_1178);
or U996 (N_996,In_1329,N_237);
and U997 (N_997,N_391,In_1161);
and U998 (N_998,In_444,N_26);
nand U999 (N_999,N_402,In_228);
or U1000 (N_1000,N_776,N_772);
nor U1001 (N_1001,N_720,N_986);
nand U1002 (N_1002,N_875,N_786);
or U1003 (N_1003,N_877,N_688);
or U1004 (N_1004,N_548,N_990);
and U1005 (N_1005,N_887,N_738);
nand U1006 (N_1006,N_943,N_897);
nand U1007 (N_1007,N_690,N_540);
or U1008 (N_1008,N_741,N_867);
nand U1009 (N_1009,N_658,N_632);
nor U1010 (N_1010,N_755,N_578);
and U1011 (N_1011,N_760,N_694);
nor U1012 (N_1012,N_872,N_790);
and U1013 (N_1013,N_662,N_863);
nand U1014 (N_1014,N_963,N_816);
and U1015 (N_1015,N_951,N_619);
nor U1016 (N_1016,N_998,N_671);
xnor U1017 (N_1017,N_546,N_811);
xor U1018 (N_1018,N_739,N_771);
or U1019 (N_1019,N_585,N_855);
and U1020 (N_1020,N_530,N_789);
or U1021 (N_1021,N_598,N_899);
nand U1022 (N_1022,N_653,N_997);
nand U1023 (N_1023,N_868,N_567);
and U1024 (N_1024,N_737,N_851);
xor U1025 (N_1025,N_660,N_940);
and U1026 (N_1026,N_876,N_707);
nand U1027 (N_1027,N_769,N_994);
xor U1028 (N_1028,N_807,N_929);
nand U1029 (N_1029,N_531,N_779);
or U1030 (N_1030,N_825,N_638);
or U1031 (N_1031,N_833,N_781);
and U1032 (N_1032,N_713,N_699);
and U1033 (N_1033,N_839,N_602);
or U1034 (N_1034,N_586,N_528);
and U1035 (N_1035,N_549,N_541);
xnor U1036 (N_1036,N_913,N_907);
nand U1037 (N_1037,N_703,N_879);
nor U1038 (N_1038,N_798,N_914);
and U1039 (N_1039,N_714,N_652);
and U1040 (N_1040,N_778,N_752);
or U1041 (N_1041,N_936,N_631);
and U1042 (N_1042,N_849,N_815);
and U1043 (N_1043,N_928,N_568);
nand U1044 (N_1044,N_821,N_980);
nand U1045 (N_1045,N_656,N_743);
nor U1046 (N_1046,N_972,N_523);
or U1047 (N_1047,N_818,N_952);
nand U1048 (N_1048,N_513,N_663);
nand U1049 (N_1049,N_844,N_831);
nand U1050 (N_1050,N_745,N_835);
nor U1051 (N_1051,N_604,N_923);
and U1052 (N_1052,N_941,N_608);
and U1053 (N_1053,N_926,N_733);
and U1054 (N_1054,N_894,N_950);
nor U1055 (N_1055,N_942,N_766);
and U1056 (N_1056,N_562,N_649);
nor U1057 (N_1057,N_757,N_906);
and U1058 (N_1058,N_637,N_981);
nand U1059 (N_1059,N_646,N_765);
or U1060 (N_1060,N_566,N_666);
xnor U1061 (N_1061,N_727,N_698);
nor U1062 (N_1062,N_916,N_582);
or U1063 (N_1063,N_915,N_510);
and U1064 (N_1064,N_725,N_558);
nand U1065 (N_1065,N_754,N_504);
nor U1066 (N_1066,N_642,N_596);
nor U1067 (N_1067,N_803,N_896);
and U1068 (N_1068,N_820,N_689);
or U1069 (N_1069,N_959,N_908);
nand U1070 (N_1070,N_945,N_946);
or U1071 (N_1071,N_670,N_607);
and U1072 (N_1072,N_597,N_934);
nor U1073 (N_1073,N_987,N_723);
and U1074 (N_1074,N_676,N_841);
nor U1075 (N_1075,N_756,N_960);
and U1076 (N_1076,N_937,N_822);
nand U1077 (N_1077,N_971,N_683);
xnor U1078 (N_1078,N_686,N_889);
and U1079 (N_1079,N_623,N_610);
nor U1080 (N_1080,N_931,N_561);
and U1081 (N_1081,N_672,N_594);
nor U1082 (N_1082,N_636,N_613);
nor U1083 (N_1083,N_912,N_615);
nor U1084 (N_1084,N_939,N_503);
or U1085 (N_1085,N_854,N_680);
nand U1086 (N_1086,N_810,N_518);
nand U1087 (N_1087,N_761,N_592);
or U1088 (N_1088,N_857,N_650);
nand U1089 (N_1089,N_774,N_826);
xor U1090 (N_1090,N_938,N_730);
nor U1091 (N_1091,N_520,N_587);
or U1092 (N_1092,N_988,N_728);
nor U1093 (N_1093,N_809,N_949);
nor U1094 (N_1094,N_590,N_622);
nand U1095 (N_1095,N_853,N_678);
xor U1096 (N_1096,N_957,N_932);
or U1097 (N_1097,N_977,N_555);
nor U1098 (N_1098,N_583,N_813);
nor U1099 (N_1099,N_791,N_910);
nor U1100 (N_1100,N_673,N_735);
or U1101 (N_1101,N_993,N_729);
nor U1102 (N_1102,N_991,N_535);
nor U1103 (N_1103,N_710,N_983);
nor U1104 (N_1104,N_655,N_639);
or U1105 (N_1105,N_511,N_917);
and U1106 (N_1106,N_967,N_859);
and U1107 (N_1107,N_969,N_775);
and U1108 (N_1108,N_836,N_697);
and U1109 (N_1109,N_659,N_601);
nor U1110 (N_1110,N_955,N_801);
nand U1111 (N_1111,N_711,N_804);
nor U1112 (N_1112,N_881,N_856);
nand U1113 (N_1113,N_848,N_995);
or U1114 (N_1114,N_536,N_878);
or U1115 (N_1115,N_519,N_600);
nor U1116 (N_1116,N_627,N_736);
and U1117 (N_1117,N_965,N_726);
nand U1118 (N_1118,N_814,N_514);
and U1119 (N_1119,N_973,N_534);
or U1120 (N_1120,N_614,N_862);
nor U1121 (N_1121,N_700,N_898);
xnor U1122 (N_1122,N_605,N_704);
nand U1123 (N_1123,N_800,N_606);
nor U1124 (N_1124,N_920,N_861);
or U1125 (N_1125,N_640,N_556);
nand U1126 (N_1126,N_538,N_718);
and U1127 (N_1127,N_834,N_992);
nor U1128 (N_1128,N_611,N_641);
nand U1129 (N_1129,N_964,N_956);
and U1130 (N_1130,N_968,N_695);
nand U1131 (N_1131,N_684,N_500);
nor U1132 (N_1132,N_537,N_616);
and U1133 (N_1133,N_651,N_989);
or U1134 (N_1134,N_505,N_565);
and U1135 (N_1135,N_824,N_576);
nand U1136 (N_1136,N_609,N_668);
nand U1137 (N_1137,N_524,N_681);
nand U1138 (N_1138,N_515,N_953);
nor U1139 (N_1139,N_793,N_958);
nand U1140 (N_1140,N_996,N_864);
and U1141 (N_1141,N_544,N_823);
nor U1142 (N_1142,N_591,N_512);
and U1143 (N_1143,N_630,N_827);
nand U1144 (N_1144,N_629,N_966);
nand U1145 (N_1145,N_679,N_644);
and U1146 (N_1146,N_753,N_621);
and U1147 (N_1147,N_922,N_732);
nand U1148 (N_1148,N_860,N_780);
nand U1149 (N_1149,N_719,N_665);
and U1150 (N_1150,N_724,N_522);
nor U1151 (N_1151,N_902,N_527);
and U1152 (N_1152,N_874,N_508);
and U1153 (N_1153,N_626,N_529);
and U1154 (N_1154,N_974,N_539);
and U1155 (N_1155,N_634,N_842);
xnor U1156 (N_1156,N_870,N_785);
xor U1157 (N_1157,N_802,N_970);
xnor U1158 (N_1158,N_805,N_551);
nor U1159 (N_1159,N_812,N_517);
or U1160 (N_1160,N_709,N_550);
and U1161 (N_1161,N_767,N_866);
and U1162 (N_1162,N_900,N_954);
and U1163 (N_1163,N_794,N_927);
and U1164 (N_1164,N_705,N_982);
or U1165 (N_1165,N_721,N_783);
nand U1166 (N_1166,N_748,N_506);
or U1167 (N_1167,N_888,N_930);
nor U1168 (N_1168,N_873,N_580);
xor U1169 (N_1169,N_693,N_645);
and U1170 (N_1170,N_925,N_817);
nor U1171 (N_1171,N_501,N_865);
nor U1172 (N_1172,N_533,N_643);
nand U1173 (N_1173,N_740,N_797);
xnor U1174 (N_1174,N_691,N_734);
nor U1175 (N_1175,N_708,N_846);
or U1176 (N_1176,N_784,N_883);
xor U1177 (N_1177,N_559,N_933);
and U1178 (N_1178,N_911,N_525);
and U1179 (N_1179,N_909,N_687);
or U1180 (N_1180,N_674,N_588);
or U1181 (N_1181,N_845,N_702);
xor U1182 (N_1182,N_819,N_787);
or U1183 (N_1183,N_507,N_742);
nand U1184 (N_1184,N_577,N_792);
nor U1185 (N_1185,N_978,N_944);
and U1186 (N_1186,N_543,N_984);
nor U1187 (N_1187,N_624,N_661);
or U1188 (N_1188,N_744,N_882);
xnor U1189 (N_1189,N_979,N_696);
and U1190 (N_1190,N_847,N_570);
or U1191 (N_1191,N_589,N_885);
nor U1192 (N_1192,N_837,N_575);
and U1193 (N_1193,N_795,N_840);
and U1194 (N_1194,N_773,N_962);
nor U1195 (N_1195,N_921,N_838);
or U1196 (N_1196,N_880,N_516);
nand U1197 (N_1197,N_750,N_788);
and U1198 (N_1198,N_749,N_901);
and U1199 (N_1199,N_947,N_722);
nor U1200 (N_1200,N_564,N_579);
and U1201 (N_1201,N_808,N_509);
nand U1202 (N_1202,N_892,N_692);
and U1203 (N_1203,N_985,N_843);
and U1204 (N_1204,N_560,N_904);
or U1205 (N_1205,N_669,N_764);
or U1206 (N_1206,N_893,N_948);
xor U1207 (N_1207,N_747,N_918);
nor U1208 (N_1208,N_620,N_664);
and U1209 (N_1209,N_657,N_850);
and U1210 (N_1210,N_572,N_829);
nand U1211 (N_1211,N_832,N_547);
or U1212 (N_1212,N_759,N_617);
nor U1213 (N_1213,N_770,N_799);
nand U1214 (N_1214,N_762,N_542);
or U1215 (N_1215,N_635,N_625);
or U1216 (N_1216,N_685,N_603);
or U1217 (N_1217,N_569,N_782);
or U1218 (N_1218,N_871,N_852);
and U1219 (N_1219,N_777,N_999);
or U1220 (N_1220,N_758,N_975);
xor U1221 (N_1221,N_595,N_891);
or U1222 (N_1222,N_633,N_701);
nor U1223 (N_1223,N_581,N_796);
or U1224 (N_1224,N_890,N_521);
nor U1225 (N_1225,N_716,N_706);
and U1226 (N_1226,N_571,N_667);
xor U1227 (N_1227,N_593,N_677);
nor U1228 (N_1228,N_731,N_712);
xnor U1229 (N_1229,N_905,N_903);
nor U1230 (N_1230,N_763,N_526);
nor U1231 (N_1231,N_828,N_746);
or U1232 (N_1232,N_584,N_599);
xor U1233 (N_1233,N_886,N_612);
or U1234 (N_1234,N_715,N_675);
nor U1235 (N_1235,N_919,N_717);
nor U1236 (N_1236,N_554,N_869);
nand U1237 (N_1237,N_552,N_573);
nand U1238 (N_1238,N_553,N_976);
or U1239 (N_1239,N_545,N_924);
nor U1240 (N_1240,N_654,N_563);
and U1241 (N_1241,N_618,N_858);
nor U1242 (N_1242,N_830,N_647);
and U1243 (N_1243,N_806,N_935);
and U1244 (N_1244,N_884,N_961);
nand U1245 (N_1245,N_895,N_682);
nand U1246 (N_1246,N_628,N_532);
or U1247 (N_1247,N_768,N_557);
nor U1248 (N_1248,N_648,N_574);
nor U1249 (N_1249,N_751,N_502);
nor U1250 (N_1250,N_615,N_653);
nor U1251 (N_1251,N_692,N_918);
nor U1252 (N_1252,N_757,N_977);
xnor U1253 (N_1253,N_549,N_555);
xnor U1254 (N_1254,N_591,N_887);
or U1255 (N_1255,N_851,N_965);
xor U1256 (N_1256,N_535,N_524);
or U1257 (N_1257,N_987,N_668);
or U1258 (N_1258,N_600,N_505);
and U1259 (N_1259,N_834,N_619);
xor U1260 (N_1260,N_640,N_643);
nor U1261 (N_1261,N_609,N_632);
nor U1262 (N_1262,N_551,N_835);
and U1263 (N_1263,N_974,N_858);
xor U1264 (N_1264,N_881,N_687);
xnor U1265 (N_1265,N_735,N_786);
or U1266 (N_1266,N_705,N_942);
or U1267 (N_1267,N_588,N_827);
and U1268 (N_1268,N_812,N_530);
nand U1269 (N_1269,N_505,N_720);
nor U1270 (N_1270,N_923,N_753);
or U1271 (N_1271,N_956,N_664);
and U1272 (N_1272,N_735,N_999);
and U1273 (N_1273,N_987,N_622);
nor U1274 (N_1274,N_995,N_928);
nor U1275 (N_1275,N_673,N_654);
nor U1276 (N_1276,N_893,N_929);
nand U1277 (N_1277,N_886,N_644);
nor U1278 (N_1278,N_905,N_793);
and U1279 (N_1279,N_654,N_745);
and U1280 (N_1280,N_736,N_580);
and U1281 (N_1281,N_569,N_548);
or U1282 (N_1282,N_850,N_846);
or U1283 (N_1283,N_945,N_852);
xnor U1284 (N_1284,N_761,N_954);
and U1285 (N_1285,N_630,N_815);
or U1286 (N_1286,N_648,N_651);
or U1287 (N_1287,N_605,N_781);
or U1288 (N_1288,N_585,N_823);
or U1289 (N_1289,N_978,N_749);
and U1290 (N_1290,N_705,N_686);
and U1291 (N_1291,N_714,N_725);
or U1292 (N_1292,N_684,N_555);
and U1293 (N_1293,N_583,N_798);
nand U1294 (N_1294,N_721,N_554);
or U1295 (N_1295,N_607,N_501);
or U1296 (N_1296,N_815,N_665);
and U1297 (N_1297,N_640,N_775);
nor U1298 (N_1298,N_598,N_876);
or U1299 (N_1299,N_945,N_582);
and U1300 (N_1300,N_588,N_933);
nand U1301 (N_1301,N_603,N_646);
or U1302 (N_1302,N_719,N_793);
or U1303 (N_1303,N_733,N_825);
nor U1304 (N_1304,N_562,N_530);
or U1305 (N_1305,N_669,N_507);
and U1306 (N_1306,N_923,N_762);
or U1307 (N_1307,N_994,N_946);
and U1308 (N_1308,N_813,N_875);
nor U1309 (N_1309,N_537,N_673);
nor U1310 (N_1310,N_976,N_628);
or U1311 (N_1311,N_564,N_697);
or U1312 (N_1312,N_961,N_824);
and U1313 (N_1313,N_954,N_599);
and U1314 (N_1314,N_853,N_895);
and U1315 (N_1315,N_688,N_589);
nor U1316 (N_1316,N_813,N_619);
and U1317 (N_1317,N_549,N_990);
nand U1318 (N_1318,N_800,N_622);
or U1319 (N_1319,N_998,N_894);
nand U1320 (N_1320,N_870,N_551);
or U1321 (N_1321,N_827,N_620);
or U1322 (N_1322,N_788,N_797);
or U1323 (N_1323,N_949,N_837);
nor U1324 (N_1324,N_591,N_628);
nand U1325 (N_1325,N_623,N_595);
nor U1326 (N_1326,N_911,N_795);
or U1327 (N_1327,N_794,N_740);
xnor U1328 (N_1328,N_772,N_735);
nor U1329 (N_1329,N_512,N_510);
or U1330 (N_1330,N_506,N_827);
or U1331 (N_1331,N_731,N_964);
nand U1332 (N_1332,N_927,N_536);
nor U1333 (N_1333,N_691,N_986);
or U1334 (N_1334,N_872,N_771);
nand U1335 (N_1335,N_827,N_639);
nor U1336 (N_1336,N_875,N_892);
and U1337 (N_1337,N_944,N_988);
or U1338 (N_1338,N_901,N_696);
or U1339 (N_1339,N_685,N_744);
nor U1340 (N_1340,N_837,N_958);
and U1341 (N_1341,N_831,N_561);
and U1342 (N_1342,N_894,N_637);
and U1343 (N_1343,N_819,N_662);
nand U1344 (N_1344,N_578,N_829);
and U1345 (N_1345,N_575,N_590);
or U1346 (N_1346,N_924,N_970);
nand U1347 (N_1347,N_643,N_937);
and U1348 (N_1348,N_546,N_602);
and U1349 (N_1349,N_935,N_977);
nor U1350 (N_1350,N_920,N_794);
or U1351 (N_1351,N_815,N_756);
nor U1352 (N_1352,N_812,N_983);
nand U1353 (N_1353,N_524,N_674);
and U1354 (N_1354,N_571,N_653);
and U1355 (N_1355,N_669,N_770);
xor U1356 (N_1356,N_792,N_501);
nor U1357 (N_1357,N_668,N_564);
nand U1358 (N_1358,N_978,N_780);
and U1359 (N_1359,N_766,N_652);
or U1360 (N_1360,N_936,N_510);
nor U1361 (N_1361,N_669,N_925);
and U1362 (N_1362,N_787,N_968);
or U1363 (N_1363,N_509,N_568);
or U1364 (N_1364,N_874,N_883);
xnor U1365 (N_1365,N_577,N_692);
nor U1366 (N_1366,N_835,N_810);
nor U1367 (N_1367,N_645,N_552);
xor U1368 (N_1368,N_904,N_736);
or U1369 (N_1369,N_545,N_660);
or U1370 (N_1370,N_500,N_702);
nand U1371 (N_1371,N_786,N_594);
and U1372 (N_1372,N_598,N_515);
nand U1373 (N_1373,N_846,N_578);
nor U1374 (N_1374,N_997,N_972);
or U1375 (N_1375,N_662,N_877);
and U1376 (N_1376,N_553,N_935);
nand U1377 (N_1377,N_528,N_728);
nor U1378 (N_1378,N_665,N_799);
nand U1379 (N_1379,N_566,N_665);
nand U1380 (N_1380,N_569,N_946);
nand U1381 (N_1381,N_567,N_668);
nand U1382 (N_1382,N_554,N_685);
nor U1383 (N_1383,N_903,N_545);
nor U1384 (N_1384,N_827,N_940);
and U1385 (N_1385,N_942,N_778);
xnor U1386 (N_1386,N_511,N_669);
nor U1387 (N_1387,N_769,N_520);
xor U1388 (N_1388,N_930,N_619);
or U1389 (N_1389,N_909,N_818);
nor U1390 (N_1390,N_961,N_542);
or U1391 (N_1391,N_967,N_923);
xor U1392 (N_1392,N_819,N_578);
nor U1393 (N_1393,N_795,N_969);
nor U1394 (N_1394,N_665,N_508);
xnor U1395 (N_1395,N_539,N_853);
nand U1396 (N_1396,N_714,N_780);
nand U1397 (N_1397,N_931,N_837);
or U1398 (N_1398,N_565,N_982);
and U1399 (N_1399,N_562,N_842);
or U1400 (N_1400,N_662,N_878);
nand U1401 (N_1401,N_739,N_947);
and U1402 (N_1402,N_948,N_657);
nor U1403 (N_1403,N_545,N_823);
nand U1404 (N_1404,N_770,N_949);
and U1405 (N_1405,N_739,N_628);
xnor U1406 (N_1406,N_724,N_822);
xor U1407 (N_1407,N_960,N_763);
and U1408 (N_1408,N_534,N_666);
nor U1409 (N_1409,N_947,N_964);
nand U1410 (N_1410,N_557,N_607);
nor U1411 (N_1411,N_960,N_929);
and U1412 (N_1412,N_675,N_946);
or U1413 (N_1413,N_857,N_847);
nand U1414 (N_1414,N_588,N_699);
xor U1415 (N_1415,N_541,N_753);
nor U1416 (N_1416,N_629,N_997);
nor U1417 (N_1417,N_795,N_577);
or U1418 (N_1418,N_541,N_514);
and U1419 (N_1419,N_602,N_986);
nor U1420 (N_1420,N_912,N_525);
and U1421 (N_1421,N_612,N_752);
nand U1422 (N_1422,N_814,N_706);
nor U1423 (N_1423,N_555,N_607);
nand U1424 (N_1424,N_684,N_847);
or U1425 (N_1425,N_983,N_646);
nand U1426 (N_1426,N_543,N_672);
nor U1427 (N_1427,N_907,N_516);
nand U1428 (N_1428,N_740,N_934);
and U1429 (N_1429,N_716,N_785);
and U1430 (N_1430,N_647,N_755);
xor U1431 (N_1431,N_863,N_608);
nor U1432 (N_1432,N_831,N_993);
nand U1433 (N_1433,N_802,N_688);
and U1434 (N_1434,N_561,N_593);
and U1435 (N_1435,N_654,N_990);
nor U1436 (N_1436,N_521,N_868);
nand U1437 (N_1437,N_542,N_639);
or U1438 (N_1438,N_516,N_507);
nand U1439 (N_1439,N_800,N_579);
or U1440 (N_1440,N_631,N_522);
xor U1441 (N_1441,N_960,N_545);
or U1442 (N_1442,N_758,N_779);
nor U1443 (N_1443,N_816,N_556);
xnor U1444 (N_1444,N_953,N_828);
and U1445 (N_1445,N_969,N_966);
and U1446 (N_1446,N_694,N_790);
nor U1447 (N_1447,N_954,N_671);
and U1448 (N_1448,N_664,N_541);
nor U1449 (N_1449,N_837,N_670);
and U1450 (N_1450,N_514,N_796);
nor U1451 (N_1451,N_559,N_520);
or U1452 (N_1452,N_548,N_550);
nor U1453 (N_1453,N_938,N_853);
nand U1454 (N_1454,N_894,N_901);
nor U1455 (N_1455,N_944,N_897);
or U1456 (N_1456,N_548,N_793);
xor U1457 (N_1457,N_915,N_913);
and U1458 (N_1458,N_850,N_615);
nand U1459 (N_1459,N_513,N_983);
nand U1460 (N_1460,N_951,N_992);
xor U1461 (N_1461,N_977,N_726);
xnor U1462 (N_1462,N_871,N_971);
and U1463 (N_1463,N_678,N_866);
or U1464 (N_1464,N_645,N_998);
nor U1465 (N_1465,N_748,N_827);
nor U1466 (N_1466,N_586,N_601);
nor U1467 (N_1467,N_795,N_934);
nor U1468 (N_1468,N_670,N_513);
nor U1469 (N_1469,N_583,N_716);
and U1470 (N_1470,N_835,N_809);
nand U1471 (N_1471,N_879,N_876);
and U1472 (N_1472,N_690,N_747);
nor U1473 (N_1473,N_515,N_607);
or U1474 (N_1474,N_747,N_626);
and U1475 (N_1475,N_847,N_542);
nand U1476 (N_1476,N_569,N_678);
or U1477 (N_1477,N_513,N_842);
and U1478 (N_1478,N_910,N_598);
nand U1479 (N_1479,N_691,N_861);
and U1480 (N_1480,N_510,N_506);
nand U1481 (N_1481,N_920,N_932);
and U1482 (N_1482,N_584,N_732);
or U1483 (N_1483,N_765,N_606);
and U1484 (N_1484,N_907,N_656);
nand U1485 (N_1485,N_747,N_550);
or U1486 (N_1486,N_684,N_617);
xnor U1487 (N_1487,N_698,N_692);
xnor U1488 (N_1488,N_645,N_624);
nand U1489 (N_1489,N_760,N_731);
nor U1490 (N_1490,N_759,N_593);
and U1491 (N_1491,N_954,N_630);
nor U1492 (N_1492,N_659,N_637);
xor U1493 (N_1493,N_537,N_584);
or U1494 (N_1494,N_515,N_789);
xnor U1495 (N_1495,N_613,N_694);
nor U1496 (N_1496,N_919,N_750);
nor U1497 (N_1497,N_806,N_645);
xor U1498 (N_1498,N_686,N_550);
nand U1499 (N_1499,N_762,N_931);
nand U1500 (N_1500,N_1028,N_1103);
or U1501 (N_1501,N_1313,N_1455);
nor U1502 (N_1502,N_1492,N_1369);
or U1503 (N_1503,N_1478,N_1005);
xor U1504 (N_1504,N_1305,N_1152);
and U1505 (N_1505,N_1402,N_1137);
and U1506 (N_1506,N_1422,N_1320);
nor U1507 (N_1507,N_1114,N_1116);
and U1508 (N_1508,N_1293,N_1197);
or U1509 (N_1509,N_1068,N_1363);
or U1510 (N_1510,N_1250,N_1310);
and U1511 (N_1511,N_1021,N_1392);
nand U1512 (N_1512,N_1190,N_1241);
or U1513 (N_1513,N_1272,N_1173);
nor U1514 (N_1514,N_1206,N_1202);
or U1515 (N_1515,N_1382,N_1047);
nor U1516 (N_1516,N_1358,N_1332);
nand U1517 (N_1517,N_1019,N_1093);
nand U1518 (N_1518,N_1312,N_1441);
nand U1519 (N_1519,N_1308,N_1396);
nand U1520 (N_1520,N_1487,N_1494);
nor U1521 (N_1521,N_1149,N_1483);
or U1522 (N_1522,N_1147,N_1124);
and U1523 (N_1523,N_1326,N_1423);
xnor U1524 (N_1524,N_1406,N_1348);
or U1525 (N_1525,N_1160,N_1444);
nor U1526 (N_1526,N_1006,N_1397);
nor U1527 (N_1527,N_1411,N_1234);
or U1528 (N_1528,N_1063,N_1327);
nor U1529 (N_1529,N_1178,N_1150);
xnor U1530 (N_1530,N_1323,N_1227);
nor U1531 (N_1531,N_1125,N_1373);
and U1532 (N_1532,N_1057,N_1471);
nor U1533 (N_1533,N_1346,N_1119);
nand U1534 (N_1534,N_1317,N_1242);
nand U1535 (N_1535,N_1398,N_1462);
nand U1536 (N_1536,N_1443,N_1438);
or U1537 (N_1537,N_1334,N_1284);
and U1538 (N_1538,N_1473,N_1211);
nand U1539 (N_1539,N_1044,N_1177);
or U1540 (N_1540,N_1385,N_1182);
and U1541 (N_1541,N_1266,N_1046);
nor U1542 (N_1542,N_1038,N_1184);
nand U1543 (N_1543,N_1145,N_1066);
or U1544 (N_1544,N_1430,N_1099);
nor U1545 (N_1545,N_1490,N_1153);
nor U1546 (N_1546,N_1498,N_1216);
and U1547 (N_1547,N_1257,N_1383);
nand U1548 (N_1548,N_1481,N_1096);
nor U1549 (N_1549,N_1208,N_1491);
nand U1550 (N_1550,N_1102,N_1017);
and U1551 (N_1551,N_1319,N_1192);
xor U1552 (N_1552,N_1378,N_1467);
xnor U1553 (N_1553,N_1070,N_1330);
and U1554 (N_1554,N_1280,N_1052);
nand U1555 (N_1555,N_1333,N_1246);
nand U1556 (N_1556,N_1094,N_1055);
and U1557 (N_1557,N_1078,N_1264);
xnor U1558 (N_1558,N_1338,N_1276);
or U1559 (N_1559,N_1384,N_1087);
and U1560 (N_1560,N_1418,N_1482);
nand U1561 (N_1561,N_1442,N_1133);
nor U1562 (N_1562,N_1477,N_1288);
and U1563 (N_1563,N_1059,N_1464);
nor U1564 (N_1564,N_1123,N_1067);
nand U1565 (N_1565,N_1433,N_1479);
and U1566 (N_1566,N_1045,N_1297);
nor U1567 (N_1567,N_1014,N_1292);
nor U1568 (N_1568,N_1085,N_1048);
xor U1569 (N_1569,N_1042,N_1159);
or U1570 (N_1570,N_1408,N_1156);
and U1571 (N_1571,N_1437,N_1409);
nand U1572 (N_1572,N_1457,N_1213);
nor U1573 (N_1573,N_1466,N_1340);
nor U1574 (N_1574,N_1108,N_1161);
nand U1575 (N_1575,N_1413,N_1454);
xnor U1576 (N_1576,N_1004,N_1432);
or U1577 (N_1577,N_1275,N_1254);
xnor U1578 (N_1578,N_1318,N_1082);
nand U1579 (N_1579,N_1375,N_1233);
nor U1580 (N_1580,N_1098,N_1097);
xnor U1581 (N_1581,N_1181,N_1261);
nor U1582 (N_1582,N_1435,N_1499);
nor U1583 (N_1583,N_1090,N_1458);
and U1584 (N_1584,N_1248,N_1429);
xor U1585 (N_1585,N_1031,N_1037);
nor U1586 (N_1586,N_1166,N_1355);
or U1587 (N_1587,N_1285,N_1100);
and U1588 (N_1588,N_1002,N_1106);
nand U1589 (N_1589,N_1474,N_1191);
and U1590 (N_1590,N_1361,N_1316);
nand U1591 (N_1591,N_1122,N_1476);
nand U1592 (N_1592,N_1277,N_1236);
and U1593 (N_1593,N_1407,N_1089);
and U1594 (N_1594,N_1302,N_1088);
and U1595 (N_1595,N_1165,N_1010);
and U1596 (N_1596,N_1342,N_1329);
nor U1597 (N_1597,N_1016,N_1064);
or U1598 (N_1598,N_1199,N_1401);
nand U1599 (N_1599,N_1018,N_1336);
nand U1600 (N_1600,N_1139,N_1395);
nor U1601 (N_1601,N_1239,N_1451);
or U1602 (N_1602,N_1209,N_1151);
or U1603 (N_1603,N_1309,N_1380);
nor U1604 (N_1604,N_1144,N_1475);
nor U1605 (N_1605,N_1304,N_1497);
xnor U1606 (N_1606,N_1142,N_1158);
and U1607 (N_1607,N_1130,N_1357);
nor U1608 (N_1608,N_1061,N_1172);
and U1609 (N_1609,N_1486,N_1225);
or U1610 (N_1610,N_1260,N_1495);
nand U1611 (N_1611,N_1036,N_1060);
and U1612 (N_1612,N_1343,N_1027);
and U1613 (N_1613,N_1207,N_1295);
and U1614 (N_1614,N_1115,N_1271);
and U1615 (N_1615,N_1091,N_1238);
nand U1616 (N_1616,N_1426,N_1269);
nor U1617 (N_1617,N_1472,N_1290);
xor U1618 (N_1618,N_1095,N_1170);
and U1619 (N_1619,N_1092,N_1388);
xnor U1620 (N_1620,N_1311,N_1185);
nand U1621 (N_1621,N_1243,N_1029);
nand U1622 (N_1622,N_1425,N_1394);
nor U1623 (N_1623,N_1240,N_1033);
nand U1624 (N_1624,N_1034,N_1132);
nand U1625 (N_1625,N_1452,N_1049);
nand U1626 (N_1626,N_1112,N_1352);
or U1627 (N_1627,N_1120,N_1465);
and U1628 (N_1628,N_1453,N_1350);
xnor U1629 (N_1629,N_1015,N_1403);
and U1630 (N_1630,N_1368,N_1393);
or U1631 (N_1631,N_1247,N_1134);
or U1632 (N_1632,N_1359,N_1174);
and U1633 (N_1633,N_1427,N_1104);
nand U1634 (N_1634,N_1303,N_1485);
nand U1635 (N_1635,N_1062,N_1307);
or U1636 (N_1636,N_1445,N_1187);
nand U1637 (N_1637,N_1267,N_1434);
nand U1638 (N_1638,N_1140,N_1030);
nand U1639 (N_1639,N_1344,N_1186);
or U1640 (N_1640,N_1306,N_1287);
or U1641 (N_1641,N_1154,N_1024);
nand U1642 (N_1642,N_1228,N_1224);
and U1643 (N_1643,N_1460,N_1180);
or U1644 (N_1644,N_1428,N_1025);
nor U1645 (N_1645,N_1203,N_1053);
nor U1646 (N_1646,N_1072,N_1171);
nand U1647 (N_1647,N_1218,N_1461);
nor U1648 (N_1648,N_1281,N_1440);
xor U1649 (N_1649,N_1127,N_1249);
and U1650 (N_1650,N_1283,N_1328);
or U1651 (N_1651,N_1164,N_1219);
nor U1652 (N_1652,N_1265,N_1043);
nand U1653 (N_1653,N_1337,N_1377);
nand U1654 (N_1654,N_1163,N_1289);
nor U1655 (N_1655,N_1069,N_1381);
or U1656 (N_1656,N_1222,N_1365);
and U1657 (N_1657,N_1488,N_1469);
nand U1658 (N_1658,N_1420,N_1003);
nand U1659 (N_1659,N_1489,N_1405);
and U1660 (N_1660,N_1496,N_1480);
xor U1661 (N_1661,N_1468,N_1282);
nand U1662 (N_1662,N_1107,N_1270);
and U1663 (N_1663,N_1065,N_1001);
or U1664 (N_1664,N_1000,N_1179);
nand U1665 (N_1665,N_1215,N_1077);
and U1666 (N_1666,N_1237,N_1217);
xor U1667 (N_1667,N_1195,N_1386);
nand U1668 (N_1668,N_1009,N_1155);
nand U1669 (N_1669,N_1020,N_1279);
nor U1670 (N_1670,N_1198,N_1353);
nand U1671 (N_1671,N_1362,N_1084);
nor U1672 (N_1672,N_1251,N_1109);
nand U1673 (N_1673,N_1414,N_1347);
nor U1674 (N_1674,N_1463,N_1417);
xnor U1675 (N_1675,N_1076,N_1175);
nand U1676 (N_1676,N_1446,N_1244);
nand U1677 (N_1677,N_1412,N_1349);
nand U1678 (N_1678,N_1449,N_1050);
and U1679 (N_1679,N_1448,N_1101);
nand U1680 (N_1680,N_1138,N_1071);
and U1681 (N_1681,N_1360,N_1141);
nor U1682 (N_1682,N_1117,N_1220);
nor U1683 (N_1683,N_1169,N_1210);
and U1684 (N_1684,N_1335,N_1374);
nor U1685 (N_1685,N_1274,N_1058);
or U1686 (N_1686,N_1136,N_1231);
nand U1687 (N_1687,N_1493,N_1011);
or U1688 (N_1688,N_1032,N_1314);
nor U1689 (N_1689,N_1322,N_1447);
or U1690 (N_1690,N_1135,N_1421);
nor U1691 (N_1691,N_1255,N_1339);
nor U1692 (N_1692,N_1252,N_1366);
or U1693 (N_1693,N_1229,N_1419);
or U1694 (N_1694,N_1113,N_1256);
nand U1695 (N_1695,N_1129,N_1054);
and U1696 (N_1696,N_1205,N_1410);
nor U1697 (N_1697,N_1325,N_1008);
or U1698 (N_1698,N_1111,N_1404);
and U1699 (N_1699,N_1399,N_1258);
and U1700 (N_1700,N_1204,N_1157);
nor U1701 (N_1701,N_1041,N_1364);
nand U1702 (N_1702,N_1194,N_1148);
and U1703 (N_1703,N_1431,N_1459);
xor U1704 (N_1704,N_1196,N_1273);
or U1705 (N_1705,N_1121,N_1299);
or U1706 (N_1706,N_1183,N_1226);
nor U1707 (N_1707,N_1012,N_1354);
xnor U1708 (N_1708,N_1301,N_1040);
nand U1709 (N_1709,N_1296,N_1118);
nand U1710 (N_1710,N_1086,N_1387);
xnor U1711 (N_1711,N_1212,N_1176);
nand U1712 (N_1712,N_1168,N_1026);
and U1713 (N_1713,N_1056,N_1263);
and U1714 (N_1714,N_1221,N_1013);
and U1715 (N_1715,N_1315,N_1105);
nor U1716 (N_1716,N_1143,N_1167);
or U1717 (N_1717,N_1356,N_1200);
or U1718 (N_1718,N_1223,N_1456);
nand U1719 (N_1719,N_1230,N_1075);
xnor U1720 (N_1720,N_1245,N_1367);
nand U1721 (N_1721,N_1131,N_1321);
nand U1722 (N_1722,N_1201,N_1390);
nor U1723 (N_1723,N_1193,N_1286);
nor U1724 (N_1724,N_1416,N_1341);
or U1725 (N_1725,N_1379,N_1470);
and U1726 (N_1726,N_1259,N_1389);
and U1727 (N_1727,N_1235,N_1450);
nand U1728 (N_1728,N_1415,N_1376);
xor U1729 (N_1729,N_1268,N_1146);
nand U1730 (N_1730,N_1214,N_1007);
nor U1731 (N_1731,N_1400,N_1345);
or U1732 (N_1732,N_1162,N_1035);
and U1733 (N_1733,N_1351,N_1391);
nand U1734 (N_1734,N_1324,N_1331);
nor U1735 (N_1735,N_1300,N_1436);
nand U1736 (N_1736,N_1023,N_1022);
or U1737 (N_1737,N_1126,N_1253);
and U1738 (N_1738,N_1484,N_1298);
nor U1739 (N_1739,N_1232,N_1291);
or U1740 (N_1740,N_1439,N_1262);
and U1741 (N_1741,N_1189,N_1424);
nand U1742 (N_1742,N_1278,N_1110);
or U1743 (N_1743,N_1039,N_1074);
nand U1744 (N_1744,N_1083,N_1370);
or U1745 (N_1745,N_1294,N_1081);
nor U1746 (N_1746,N_1371,N_1051);
nand U1747 (N_1747,N_1128,N_1073);
nand U1748 (N_1748,N_1188,N_1079);
nand U1749 (N_1749,N_1080,N_1372);
and U1750 (N_1750,N_1173,N_1343);
nor U1751 (N_1751,N_1082,N_1474);
and U1752 (N_1752,N_1414,N_1269);
and U1753 (N_1753,N_1393,N_1239);
or U1754 (N_1754,N_1305,N_1297);
nor U1755 (N_1755,N_1403,N_1460);
nand U1756 (N_1756,N_1469,N_1276);
or U1757 (N_1757,N_1182,N_1331);
or U1758 (N_1758,N_1472,N_1035);
and U1759 (N_1759,N_1152,N_1346);
nor U1760 (N_1760,N_1148,N_1253);
and U1761 (N_1761,N_1003,N_1058);
nand U1762 (N_1762,N_1192,N_1315);
nor U1763 (N_1763,N_1210,N_1265);
or U1764 (N_1764,N_1195,N_1353);
nor U1765 (N_1765,N_1473,N_1345);
nor U1766 (N_1766,N_1453,N_1221);
or U1767 (N_1767,N_1316,N_1092);
nor U1768 (N_1768,N_1044,N_1042);
nor U1769 (N_1769,N_1418,N_1400);
and U1770 (N_1770,N_1109,N_1478);
xnor U1771 (N_1771,N_1224,N_1494);
or U1772 (N_1772,N_1491,N_1001);
nand U1773 (N_1773,N_1358,N_1008);
or U1774 (N_1774,N_1158,N_1182);
nor U1775 (N_1775,N_1372,N_1283);
xor U1776 (N_1776,N_1170,N_1245);
nor U1777 (N_1777,N_1167,N_1236);
nand U1778 (N_1778,N_1333,N_1080);
and U1779 (N_1779,N_1078,N_1272);
nor U1780 (N_1780,N_1014,N_1030);
xnor U1781 (N_1781,N_1150,N_1443);
nor U1782 (N_1782,N_1393,N_1126);
nor U1783 (N_1783,N_1234,N_1153);
or U1784 (N_1784,N_1216,N_1462);
xnor U1785 (N_1785,N_1249,N_1106);
nor U1786 (N_1786,N_1254,N_1062);
or U1787 (N_1787,N_1251,N_1405);
nor U1788 (N_1788,N_1499,N_1144);
nand U1789 (N_1789,N_1118,N_1105);
or U1790 (N_1790,N_1479,N_1464);
or U1791 (N_1791,N_1056,N_1254);
nand U1792 (N_1792,N_1427,N_1189);
and U1793 (N_1793,N_1340,N_1211);
or U1794 (N_1794,N_1232,N_1139);
and U1795 (N_1795,N_1472,N_1036);
nor U1796 (N_1796,N_1064,N_1059);
nand U1797 (N_1797,N_1202,N_1458);
and U1798 (N_1798,N_1323,N_1195);
or U1799 (N_1799,N_1413,N_1053);
or U1800 (N_1800,N_1179,N_1445);
nand U1801 (N_1801,N_1256,N_1207);
nor U1802 (N_1802,N_1186,N_1011);
or U1803 (N_1803,N_1307,N_1337);
or U1804 (N_1804,N_1168,N_1282);
nor U1805 (N_1805,N_1438,N_1291);
nor U1806 (N_1806,N_1347,N_1366);
and U1807 (N_1807,N_1155,N_1204);
nor U1808 (N_1808,N_1013,N_1355);
and U1809 (N_1809,N_1032,N_1303);
or U1810 (N_1810,N_1401,N_1448);
nand U1811 (N_1811,N_1023,N_1448);
or U1812 (N_1812,N_1474,N_1493);
or U1813 (N_1813,N_1102,N_1057);
nand U1814 (N_1814,N_1292,N_1097);
nand U1815 (N_1815,N_1468,N_1274);
nor U1816 (N_1816,N_1444,N_1081);
xnor U1817 (N_1817,N_1124,N_1478);
nand U1818 (N_1818,N_1213,N_1196);
or U1819 (N_1819,N_1006,N_1056);
and U1820 (N_1820,N_1351,N_1081);
nor U1821 (N_1821,N_1468,N_1186);
and U1822 (N_1822,N_1063,N_1004);
or U1823 (N_1823,N_1092,N_1056);
and U1824 (N_1824,N_1353,N_1266);
nand U1825 (N_1825,N_1292,N_1040);
nand U1826 (N_1826,N_1423,N_1196);
nand U1827 (N_1827,N_1394,N_1483);
nor U1828 (N_1828,N_1370,N_1063);
and U1829 (N_1829,N_1265,N_1221);
and U1830 (N_1830,N_1294,N_1224);
or U1831 (N_1831,N_1400,N_1102);
or U1832 (N_1832,N_1469,N_1355);
or U1833 (N_1833,N_1024,N_1210);
and U1834 (N_1834,N_1433,N_1419);
or U1835 (N_1835,N_1043,N_1478);
or U1836 (N_1836,N_1085,N_1060);
xor U1837 (N_1837,N_1327,N_1040);
and U1838 (N_1838,N_1300,N_1411);
nor U1839 (N_1839,N_1333,N_1353);
and U1840 (N_1840,N_1352,N_1150);
nor U1841 (N_1841,N_1181,N_1404);
nand U1842 (N_1842,N_1028,N_1490);
and U1843 (N_1843,N_1227,N_1272);
or U1844 (N_1844,N_1256,N_1333);
nor U1845 (N_1845,N_1289,N_1395);
nand U1846 (N_1846,N_1223,N_1302);
nor U1847 (N_1847,N_1321,N_1403);
or U1848 (N_1848,N_1253,N_1247);
or U1849 (N_1849,N_1061,N_1406);
nor U1850 (N_1850,N_1410,N_1476);
nor U1851 (N_1851,N_1434,N_1038);
nor U1852 (N_1852,N_1222,N_1095);
nor U1853 (N_1853,N_1182,N_1392);
or U1854 (N_1854,N_1290,N_1408);
nor U1855 (N_1855,N_1163,N_1371);
nor U1856 (N_1856,N_1424,N_1298);
or U1857 (N_1857,N_1188,N_1487);
xnor U1858 (N_1858,N_1168,N_1060);
nand U1859 (N_1859,N_1019,N_1207);
xor U1860 (N_1860,N_1454,N_1151);
and U1861 (N_1861,N_1328,N_1479);
or U1862 (N_1862,N_1195,N_1062);
and U1863 (N_1863,N_1042,N_1438);
or U1864 (N_1864,N_1102,N_1433);
nor U1865 (N_1865,N_1387,N_1262);
nor U1866 (N_1866,N_1178,N_1490);
nor U1867 (N_1867,N_1404,N_1406);
and U1868 (N_1868,N_1254,N_1357);
or U1869 (N_1869,N_1411,N_1464);
or U1870 (N_1870,N_1311,N_1065);
and U1871 (N_1871,N_1220,N_1381);
or U1872 (N_1872,N_1272,N_1253);
nand U1873 (N_1873,N_1293,N_1373);
and U1874 (N_1874,N_1080,N_1129);
xnor U1875 (N_1875,N_1153,N_1249);
and U1876 (N_1876,N_1035,N_1071);
and U1877 (N_1877,N_1415,N_1138);
nor U1878 (N_1878,N_1012,N_1415);
and U1879 (N_1879,N_1461,N_1153);
nor U1880 (N_1880,N_1265,N_1413);
and U1881 (N_1881,N_1096,N_1330);
nor U1882 (N_1882,N_1346,N_1140);
nor U1883 (N_1883,N_1129,N_1261);
nand U1884 (N_1884,N_1255,N_1487);
nand U1885 (N_1885,N_1457,N_1186);
or U1886 (N_1886,N_1346,N_1298);
nor U1887 (N_1887,N_1470,N_1210);
nor U1888 (N_1888,N_1315,N_1491);
nand U1889 (N_1889,N_1213,N_1364);
and U1890 (N_1890,N_1079,N_1094);
or U1891 (N_1891,N_1276,N_1203);
nand U1892 (N_1892,N_1187,N_1087);
nor U1893 (N_1893,N_1445,N_1234);
nor U1894 (N_1894,N_1035,N_1216);
or U1895 (N_1895,N_1335,N_1468);
nand U1896 (N_1896,N_1167,N_1013);
nor U1897 (N_1897,N_1449,N_1297);
nor U1898 (N_1898,N_1122,N_1327);
nand U1899 (N_1899,N_1229,N_1149);
and U1900 (N_1900,N_1123,N_1483);
nor U1901 (N_1901,N_1274,N_1218);
or U1902 (N_1902,N_1119,N_1410);
nor U1903 (N_1903,N_1416,N_1028);
or U1904 (N_1904,N_1229,N_1337);
nand U1905 (N_1905,N_1080,N_1007);
or U1906 (N_1906,N_1184,N_1202);
nor U1907 (N_1907,N_1096,N_1060);
nor U1908 (N_1908,N_1483,N_1116);
nand U1909 (N_1909,N_1117,N_1382);
nand U1910 (N_1910,N_1024,N_1377);
or U1911 (N_1911,N_1316,N_1090);
and U1912 (N_1912,N_1221,N_1479);
nor U1913 (N_1913,N_1231,N_1305);
nand U1914 (N_1914,N_1310,N_1161);
nor U1915 (N_1915,N_1151,N_1137);
and U1916 (N_1916,N_1375,N_1079);
and U1917 (N_1917,N_1349,N_1079);
nand U1918 (N_1918,N_1090,N_1095);
nor U1919 (N_1919,N_1359,N_1405);
nor U1920 (N_1920,N_1316,N_1128);
xor U1921 (N_1921,N_1170,N_1111);
and U1922 (N_1922,N_1067,N_1266);
and U1923 (N_1923,N_1301,N_1420);
or U1924 (N_1924,N_1228,N_1457);
and U1925 (N_1925,N_1373,N_1127);
nor U1926 (N_1926,N_1175,N_1151);
nand U1927 (N_1927,N_1407,N_1477);
nor U1928 (N_1928,N_1143,N_1215);
nor U1929 (N_1929,N_1160,N_1043);
or U1930 (N_1930,N_1447,N_1445);
or U1931 (N_1931,N_1047,N_1035);
xnor U1932 (N_1932,N_1472,N_1211);
nand U1933 (N_1933,N_1247,N_1161);
and U1934 (N_1934,N_1304,N_1045);
or U1935 (N_1935,N_1372,N_1260);
nand U1936 (N_1936,N_1455,N_1207);
and U1937 (N_1937,N_1144,N_1408);
xnor U1938 (N_1938,N_1120,N_1037);
nor U1939 (N_1939,N_1338,N_1102);
xnor U1940 (N_1940,N_1261,N_1177);
nor U1941 (N_1941,N_1405,N_1036);
nor U1942 (N_1942,N_1217,N_1111);
nand U1943 (N_1943,N_1454,N_1183);
and U1944 (N_1944,N_1300,N_1006);
and U1945 (N_1945,N_1147,N_1414);
and U1946 (N_1946,N_1111,N_1140);
nand U1947 (N_1947,N_1075,N_1259);
nor U1948 (N_1948,N_1139,N_1267);
and U1949 (N_1949,N_1314,N_1004);
nand U1950 (N_1950,N_1353,N_1446);
nand U1951 (N_1951,N_1482,N_1413);
nor U1952 (N_1952,N_1275,N_1252);
nand U1953 (N_1953,N_1271,N_1383);
nor U1954 (N_1954,N_1443,N_1127);
nand U1955 (N_1955,N_1108,N_1286);
nand U1956 (N_1956,N_1023,N_1291);
nand U1957 (N_1957,N_1207,N_1401);
xor U1958 (N_1958,N_1235,N_1224);
and U1959 (N_1959,N_1054,N_1168);
nand U1960 (N_1960,N_1234,N_1303);
nand U1961 (N_1961,N_1499,N_1063);
nand U1962 (N_1962,N_1025,N_1220);
or U1963 (N_1963,N_1124,N_1234);
nand U1964 (N_1964,N_1335,N_1312);
nor U1965 (N_1965,N_1452,N_1078);
xnor U1966 (N_1966,N_1159,N_1151);
nor U1967 (N_1967,N_1292,N_1317);
xor U1968 (N_1968,N_1445,N_1159);
nor U1969 (N_1969,N_1093,N_1261);
nor U1970 (N_1970,N_1309,N_1472);
and U1971 (N_1971,N_1252,N_1473);
nand U1972 (N_1972,N_1208,N_1424);
nand U1973 (N_1973,N_1211,N_1205);
and U1974 (N_1974,N_1089,N_1054);
or U1975 (N_1975,N_1406,N_1294);
xor U1976 (N_1976,N_1111,N_1371);
and U1977 (N_1977,N_1333,N_1355);
nand U1978 (N_1978,N_1220,N_1082);
nor U1979 (N_1979,N_1382,N_1224);
nand U1980 (N_1980,N_1248,N_1301);
and U1981 (N_1981,N_1356,N_1365);
xor U1982 (N_1982,N_1332,N_1216);
or U1983 (N_1983,N_1178,N_1086);
nand U1984 (N_1984,N_1064,N_1396);
or U1985 (N_1985,N_1232,N_1313);
nor U1986 (N_1986,N_1213,N_1125);
and U1987 (N_1987,N_1464,N_1449);
nor U1988 (N_1988,N_1337,N_1437);
xnor U1989 (N_1989,N_1498,N_1324);
nand U1990 (N_1990,N_1351,N_1450);
and U1991 (N_1991,N_1129,N_1116);
or U1992 (N_1992,N_1001,N_1203);
nor U1993 (N_1993,N_1222,N_1126);
or U1994 (N_1994,N_1323,N_1140);
nand U1995 (N_1995,N_1438,N_1165);
or U1996 (N_1996,N_1063,N_1425);
nor U1997 (N_1997,N_1371,N_1361);
and U1998 (N_1998,N_1489,N_1161);
and U1999 (N_1999,N_1391,N_1037);
or U2000 (N_2000,N_1538,N_1814);
nand U2001 (N_2001,N_1816,N_1830);
and U2002 (N_2002,N_1823,N_1920);
nand U2003 (N_2003,N_1588,N_1973);
xnor U2004 (N_2004,N_1528,N_1811);
or U2005 (N_2005,N_1547,N_1839);
nor U2006 (N_2006,N_1789,N_1662);
or U2007 (N_2007,N_1592,N_1820);
and U2008 (N_2008,N_1618,N_1878);
xor U2009 (N_2009,N_1784,N_1772);
nand U2010 (N_2010,N_1629,N_1624);
xnor U2011 (N_2011,N_1831,N_1711);
and U2012 (N_2012,N_1518,N_1637);
nand U2013 (N_2013,N_1905,N_1634);
nand U2014 (N_2014,N_1663,N_1855);
nor U2015 (N_2015,N_1986,N_1694);
and U2016 (N_2016,N_1644,N_1529);
xor U2017 (N_2017,N_1543,N_1919);
nand U2018 (N_2018,N_1924,N_1654);
nor U2019 (N_2019,N_1950,N_1719);
nand U2020 (N_2020,N_1619,N_1642);
and U2021 (N_2021,N_1767,N_1959);
and U2022 (N_2022,N_1677,N_1628);
nor U2023 (N_2023,N_1631,N_1601);
and U2024 (N_2024,N_1550,N_1936);
nand U2025 (N_2025,N_1569,N_1896);
nor U2026 (N_2026,N_1753,N_1951);
nand U2027 (N_2027,N_1740,N_1974);
nand U2028 (N_2028,N_1791,N_1828);
nor U2029 (N_2029,N_1777,N_1698);
or U2030 (N_2030,N_1599,N_1940);
or U2031 (N_2031,N_1926,N_1724);
nor U2032 (N_2032,N_1587,N_1860);
nand U2033 (N_2033,N_1801,N_1602);
nand U2034 (N_2034,N_1612,N_1840);
nor U2035 (N_2035,N_1989,N_1848);
xnor U2036 (N_2036,N_1751,N_1763);
and U2037 (N_2037,N_1704,N_1967);
nor U2038 (N_2038,N_1870,N_1583);
and U2039 (N_2039,N_1510,N_1903);
nand U2040 (N_2040,N_1540,N_1630);
nand U2041 (N_2041,N_1858,N_1513);
or U2042 (N_2042,N_1609,N_1768);
and U2043 (N_2043,N_1982,N_1687);
nand U2044 (N_2044,N_1625,N_1682);
nor U2045 (N_2045,N_1503,N_1780);
or U2046 (N_2046,N_1552,N_1627);
nand U2047 (N_2047,N_1865,N_1721);
nand U2048 (N_2048,N_1661,N_1727);
nand U2049 (N_2049,N_1658,N_1707);
nand U2050 (N_2050,N_1509,N_1957);
and U2051 (N_2051,N_1832,N_1922);
nor U2052 (N_2052,N_1633,N_1760);
nor U2053 (N_2053,N_1668,N_1802);
nor U2054 (N_2054,N_1526,N_1966);
or U2055 (N_2055,N_1736,N_1696);
nand U2056 (N_2056,N_1758,N_1894);
and U2057 (N_2057,N_1665,N_1871);
nor U2058 (N_2058,N_1530,N_1659);
nor U2059 (N_2059,N_1866,N_1714);
and U2060 (N_2060,N_1873,N_1700);
and U2061 (N_2061,N_1891,N_1626);
or U2062 (N_2062,N_1807,N_1810);
and U2063 (N_2063,N_1614,N_1988);
or U2064 (N_2064,N_1885,N_1710);
nor U2065 (N_2065,N_1589,N_1971);
nor U2066 (N_2066,N_1799,N_1671);
nor U2067 (N_2067,N_1541,N_1676);
or U2068 (N_2068,N_1718,N_1958);
and U2069 (N_2069,N_1819,N_1506);
and U2070 (N_2070,N_1557,N_1869);
or U2071 (N_2071,N_1712,N_1693);
nand U2072 (N_2072,N_1586,N_1930);
and U2073 (N_2073,N_1527,N_1674);
and U2074 (N_2074,N_1759,N_1638);
xnor U2075 (N_2075,N_1623,N_1603);
nor U2076 (N_2076,N_1722,N_1741);
nor U2077 (N_2077,N_1742,N_1852);
nand U2078 (N_2078,N_1987,N_1549);
and U2079 (N_2079,N_1821,N_1998);
or U2080 (N_2080,N_1845,N_1516);
and U2081 (N_2081,N_1617,N_1895);
nand U2082 (N_2082,N_1666,N_1689);
and U2083 (N_2083,N_1981,N_1686);
nand U2084 (N_2084,N_1796,N_1884);
and U2085 (N_2085,N_1706,N_1641);
xnor U2086 (N_2086,N_1565,N_1771);
nand U2087 (N_2087,N_1916,N_1582);
and U2088 (N_2088,N_1846,N_1675);
nand U2089 (N_2089,N_1798,N_1766);
or U2090 (N_2090,N_1639,N_1773);
xnor U2091 (N_2091,N_1524,N_1915);
and U2092 (N_2092,N_1648,N_1572);
and U2093 (N_2093,N_1531,N_1669);
and U2094 (N_2094,N_1756,N_1782);
nand U2095 (N_2095,N_1535,N_1908);
nand U2096 (N_2096,N_1861,N_1786);
or U2097 (N_2097,N_1570,N_1836);
nor U2098 (N_2098,N_1739,N_1720);
nor U2099 (N_2099,N_1750,N_1859);
or U2100 (N_2100,N_1748,N_1523);
and U2101 (N_2101,N_1953,N_1731);
nor U2102 (N_2102,N_1948,N_1934);
nand U2103 (N_2103,N_1611,N_1684);
and U2104 (N_2104,N_1900,N_1838);
nand U2105 (N_2105,N_1598,N_1909);
nand U2106 (N_2106,N_1558,N_1923);
nor U2107 (N_2107,N_1749,N_1925);
nor U2108 (N_2108,N_1868,N_1581);
or U2109 (N_2109,N_1809,N_1702);
nor U2110 (N_2110,N_1555,N_1996);
and U2111 (N_2111,N_1508,N_1656);
and U2112 (N_2112,N_1514,N_1716);
xor U2113 (N_2113,N_1551,N_1519);
nor U2114 (N_2114,N_1833,N_1879);
nand U2115 (N_2115,N_1680,N_1822);
nand U2116 (N_2116,N_1670,N_1785);
xnor U2117 (N_2117,N_1708,N_1553);
nor U2118 (N_2118,N_1912,N_1856);
and U2119 (N_2119,N_1968,N_1571);
nor U2120 (N_2120,N_1576,N_1517);
and U2121 (N_2121,N_1781,N_1521);
nand U2122 (N_2122,N_1764,N_1537);
nand U2123 (N_2123,N_1673,N_1575);
or U2124 (N_2124,N_1824,N_1887);
and U2125 (N_2125,N_1774,N_1732);
and U2126 (N_2126,N_1790,N_1985);
nand U2127 (N_2127,N_1757,N_1688);
nor U2128 (N_2128,N_1899,N_1640);
nor U2129 (N_2129,N_1937,N_1815);
or U2130 (N_2130,N_1544,N_1844);
and U2131 (N_2131,N_1679,N_1835);
and U2132 (N_2132,N_1520,N_1596);
xor U2133 (N_2133,N_1562,N_1837);
nor U2134 (N_2134,N_1901,N_1536);
and U2135 (N_2135,N_1697,N_1882);
or U2136 (N_2136,N_1733,N_1797);
or U2137 (N_2137,N_1929,N_1853);
xor U2138 (N_2138,N_1792,N_1897);
and U2139 (N_2139,N_1761,N_1534);
and U2140 (N_2140,N_1713,N_1939);
or U2141 (N_2141,N_1862,N_1994);
or U2142 (N_2142,N_1842,N_1977);
and U2143 (N_2143,N_1995,N_1651);
nor U2144 (N_2144,N_1646,N_1608);
and U2145 (N_2145,N_1590,N_1808);
and U2146 (N_2146,N_1818,N_1867);
nand U2147 (N_2147,N_1681,N_1813);
and U2148 (N_2148,N_1843,N_1902);
nand U2149 (N_2149,N_1705,N_1613);
or U2150 (N_2150,N_1965,N_1657);
or U2151 (N_2151,N_1755,N_1573);
nand U2152 (N_2152,N_1723,N_1997);
nor U2153 (N_2153,N_1875,N_1956);
and U2154 (N_2154,N_1595,N_1672);
nor U2155 (N_2155,N_1512,N_1622);
or U2156 (N_2156,N_1765,N_1574);
nor U2157 (N_2157,N_1593,N_1970);
nand U2158 (N_2158,N_1795,N_1561);
nor U2159 (N_2159,N_1580,N_1690);
or U2160 (N_2160,N_1947,N_1804);
xor U2161 (N_2161,N_1876,N_1938);
nor U2162 (N_2162,N_1647,N_1643);
and U2163 (N_2163,N_1717,N_1505);
or U2164 (N_2164,N_1610,N_1776);
nor U2165 (N_2165,N_1730,N_1888);
nor U2166 (N_2166,N_1556,N_1964);
nor U2167 (N_2167,N_1746,N_1584);
nor U2168 (N_2168,N_1542,N_1825);
nor U2169 (N_2169,N_1931,N_1918);
xor U2170 (N_2170,N_1847,N_1744);
and U2171 (N_2171,N_1907,N_1991);
nor U2172 (N_2172,N_1525,N_1889);
nor U2173 (N_2173,N_1652,N_1921);
nand U2174 (N_2174,N_1893,N_1883);
nor U2175 (N_2175,N_1794,N_1683);
nand U2176 (N_2176,N_1747,N_1863);
nand U2177 (N_2177,N_1546,N_1726);
nor U2178 (N_2178,N_1635,N_1892);
xnor U2179 (N_2179,N_1806,N_1655);
or U2180 (N_2180,N_1660,N_1783);
xnor U2181 (N_2181,N_1649,N_1738);
nor U2182 (N_2182,N_1567,N_1913);
or U2183 (N_2183,N_1954,N_1944);
nor U2184 (N_2184,N_1984,N_1539);
nor U2185 (N_2185,N_1793,N_1961);
or U2186 (N_2186,N_1829,N_1729);
and U2187 (N_2187,N_1927,N_1645);
and U2188 (N_2188,N_1910,N_1872);
nand U2189 (N_2189,N_1577,N_1545);
and U2190 (N_2190,N_1933,N_1734);
and U2191 (N_2191,N_1701,N_1834);
or U2192 (N_2192,N_1591,N_1850);
or U2193 (N_2193,N_1743,N_1963);
nand U2194 (N_2194,N_1857,N_1864);
or U2195 (N_2195,N_1597,N_1616);
nand U2196 (N_2196,N_1501,N_1606);
nand U2197 (N_2197,N_1849,N_1880);
or U2198 (N_2198,N_1502,N_1972);
or U2199 (N_2199,N_1805,N_1621);
or U2200 (N_2200,N_1906,N_1911);
nor U2201 (N_2201,N_1980,N_1932);
xnor U2202 (N_2202,N_1678,N_1990);
nand U2203 (N_2203,N_1935,N_1955);
or U2204 (N_2204,N_1564,N_1620);
and U2205 (N_2205,N_1507,N_1600);
xor U2206 (N_2206,N_1578,N_1664);
nand U2207 (N_2207,N_1715,N_1942);
xor U2208 (N_2208,N_1969,N_1607);
nor U2209 (N_2209,N_1874,N_1917);
nand U2210 (N_2210,N_1904,N_1803);
xnor U2211 (N_2211,N_1952,N_1554);
or U2212 (N_2212,N_1500,N_1703);
xor U2213 (N_2213,N_1653,N_1841);
or U2214 (N_2214,N_1788,N_1787);
nor U2215 (N_2215,N_1594,N_1975);
or U2216 (N_2216,N_1999,N_1559);
nand U2217 (N_2217,N_1745,N_1983);
and U2218 (N_2218,N_1560,N_1737);
and U2219 (N_2219,N_1946,N_1691);
nand U2220 (N_2220,N_1886,N_1898);
nor U2221 (N_2221,N_1854,N_1754);
or U2222 (N_2222,N_1585,N_1604);
nor U2223 (N_2223,N_1881,N_1725);
and U2224 (N_2224,N_1566,N_1563);
nand U2225 (N_2225,N_1532,N_1504);
nand U2226 (N_2226,N_1812,N_1515);
and U2227 (N_2227,N_1817,N_1976);
nor U2228 (N_2228,N_1709,N_1992);
xor U2229 (N_2229,N_1778,N_1533);
and U2230 (N_2230,N_1914,N_1779);
nor U2231 (N_2231,N_1579,N_1877);
xor U2232 (N_2232,N_1941,N_1692);
or U2233 (N_2233,N_1978,N_1699);
nand U2234 (N_2234,N_1979,N_1827);
nand U2235 (N_2235,N_1615,N_1650);
or U2236 (N_2236,N_1667,N_1949);
and U2237 (N_2237,N_1775,N_1548);
nand U2238 (N_2238,N_1800,N_1685);
nand U2239 (N_2239,N_1568,N_1943);
and U2240 (N_2240,N_1960,N_1993);
and U2241 (N_2241,N_1762,N_1511);
or U2242 (N_2242,N_1695,N_1851);
nor U2243 (N_2243,N_1752,N_1769);
nand U2244 (N_2244,N_1962,N_1928);
or U2245 (N_2245,N_1728,N_1605);
nand U2246 (N_2246,N_1770,N_1890);
nor U2247 (N_2247,N_1636,N_1632);
or U2248 (N_2248,N_1945,N_1826);
and U2249 (N_2249,N_1522,N_1735);
nand U2250 (N_2250,N_1809,N_1624);
or U2251 (N_2251,N_1800,N_1975);
or U2252 (N_2252,N_1600,N_1663);
nand U2253 (N_2253,N_1618,N_1751);
or U2254 (N_2254,N_1850,N_1974);
and U2255 (N_2255,N_1835,N_1916);
nand U2256 (N_2256,N_1506,N_1781);
and U2257 (N_2257,N_1738,N_1616);
and U2258 (N_2258,N_1800,N_1615);
nand U2259 (N_2259,N_1665,N_1839);
and U2260 (N_2260,N_1824,N_1620);
or U2261 (N_2261,N_1722,N_1746);
or U2262 (N_2262,N_1577,N_1956);
nor U2263 (N_2263,N_1729,N_1749);
nand U2264 (N_2264,N_1510,N_1841);
or U2265 (N_2265,N_1690,N_1952);
and U2266 (N_2266,N_1694,N_1720);
nand U2267 (N_2267,N_1564,N_1956);
or U2268 (N_2268,N_1797,N_1625);
or U2269 (N_2269,N_1658,N_1796);
xnor U2270 (N_2270,N_1786,N_1918);
and U2271 (N_2271,N_1951,N_1676);
or U2272 (N_2272,N_1790,N_1812);
and U2273 (N_2273,N_1922,N_1731);
or U2274 (N_2274,N_1591,N_1612);
xor U2275 (N_2275,N_1939,N_1625);
and U2276 (N_2276,N_1968,N_1709);
nand U2277 (N_2277,N_1949,N_1611);
nand U2278 (N_2278,N_1627,N_1761);
and U2279 (N_2279,N_1880,N_1886);
and U2280 (N_2280,N_1698,N_1903);
and U2281 (N_2281,N_1791,N_1920);
and U2282 (N_2282,N_1516,N_1829);
or U2283 (N_2283,N_1726,N_1559);
or U2284 (N_2284,N_1760,N_1623);
nor U2285 (N_2285,N_1537,N_1853);
nand U2286 (N_2286,N_1763,N_1990);
nor U2287 (N_2287,N_1622,N_1846);
xor U2288 (N_2288,N_1574,N_1666);
xnor U2289 (N_2289,N_1849,N_1845);
nand U2290 (N_2290,N_1766,N_1924);
xnor U2291 (N_2291,N_1797,N_1964);
nor U2292 (N_2292,N_1932,N_1600);
nor U2293 (N_2293,N_1811,N_1533);
nand U2294 (N_2294,N_1866,N_1701);
or U2295 (N_2295,N_1611,N_1516);
nor U2296 (N_2296,N_1527,N_1517);
nand U2297 (N_2297,N_1842,N_1810);
nand U2298 (N_2298,N_1678,N_1950);
nand U2299 (N_2299,N_1703,N_1862);
nor U2300 (N_2300,N_1729,N_1974);
or U2301 (N_2301,N_1925,N_1637);
and U2302 (N_2302,N_1582,N_1885);
or U2303 (N_2303,N_1518,N_1770);
nand U2304 (N_2304,N_1739,N_1856);
nand U2305 (N_2305,N_1536,N_1533);
nor U2306 (N_2306,N_1605,N_1747);
nand U2307 (N_2307,N_1827,N_1637);
nand U2308 (N_2308,N_1531,N_1874);
or U2309 (N_2309,N_1534,N_1592);
xor U2310 (N_2310,N_1502,N_1722);
and U2311 (N_2311,N_1867,N_1975);
or U2312 (N_2312,N_1751,N_1721);
nor U2313 (N_2313,N_1996,N_1823);
nor U2314 (N_2314,N_1864,N_1871);
xnor U2315 (N_2315,N_1910,N_1582);
or U2316 (N_2316,N_1785,N_1520);
and U2317 (N_2317,N_1544,N_1792);
nor U2318 (N_2318,N_1589,N_1945);
nand U2319 (N_2319,N_1906,N_1659);
nand U2320 (N_2320,N_1937,N_1645);
or U2321 (N_2321,N_1998,N_1693);
nand U2322 (N_2322,N_1747,N_1716);
nand U2323 (N_2323,N_1870,N_1859);
or U2324 (N_2324,N_1669,N_1602);
or U2325 (N_2325,N_1828,N_1741);
or U2326 (N_2326,N_1833,N_1515);
nand U2327 (N_2327,N_1897,N_1621);
and U2328 (N_2328,N_1550,N_1735);
nor U2329 (N_2329,N_1570,N_1782);
and U2330 (N_2330,N_1900,N_1603);
nand U2331 (N_2331,N_1797,N_1992);
and U2332 (N_2332,N_1813,N_1761);
nand U2333 (N_2333,N_1585,N_1870);
and U2334 (N_2334,N_1838,N_1779);
and U2335 (N_2335,N_1982,N_1915);
nor U2336 (N_2336,N_1751,N_1689);
or U2337 (N_2337,N_1872,N_1717);
or U2338 (N_2338,N_1594,N_1579);
and U2339 (N_2339,N_1517,N_1971);
and U2340 (N_2340,N_1522,N_1555);
and U2341 (N_2341,N_1827,N_1729);
nor U2342 (N_2342,N_1900,N_1942);
nand U2343 (N_2343,N_1841,N_1561);
nand U2344 (N_2344,N_1824,N_1692);
and U2345 (N_2345,N_1556,N_1821);
nor U2346 (N_2346,N_1796,N_1922);
nor U2347 (N_2347,N_1582,N_1743);
and U2348 (N_2348,N_1905,N_1955);
or U2349 (N_2349,N_1525,N_1513);
and U2350 (N_2350,N_1590,N_1579);
and U2351 (N_2351,N_1612,N_1912);
and U2352 (N_2352,N_1763,N_1650);
nand U2353 (N_2353,N_1979,N_1633);
nor U2354 (N_2354,N_1665,N_1951);
and U2355 (N_2355,N_1567,N_1743);
and U2356 (N_2356,N_1570,N_1881);
xnor U2357 (N_2357,N_1828,N_1576);
and U2358 (N_2358,N_1907,N_1732);
or U2359 (N_2359,N_1647,N_1895);
and U2360 (N_2360,N_1811,N_1894);
and U2361 (N_2361,N_1651,N_1638);
nand U2362 (N_2362,N_1547,N_1729);
or U2363 (N_2363,N_1562,N_1689);
or U2364 (N_2364,N_1827,N_1529);
xnor U2365 (N_2365,N_1563,N_1876);
nand U2366 (N_2366,N_1818,N_1570);
or U2367 (N_2367,N_1519,N_1716);
nand U2368 (N_2368,N_1609,N_1742);
and U2369 (N_2369,N_1817,N_1642);
xnor U2370 (N_2370,N_1593,N_1544);
or U2371 (N_2371,N_1654,N_1669);
nand U2372 (N_2372,N_1556,N_1790);
nor U2373 (N_2373,N_1657,N_1865);
or U2374 (N_2374,N_1668,N_1938);
nand U2375 (N_2375,N_1952,N_1754);
or U2376 (N_2376,N_1530,N_1845);
nand U2377 (N_2377,N_1725,N_1873);
nand U2378 (N_2378,N_1581,N_1890);
and U2379 (N_2379,N_1747,N_1535);
nor U2380 (N_2380,N_1601,N_1821);
nor U2381 (N_2381,N_1721,N_1850);
and U2382 (N_2382,N_1963,N_1668);
nor U2383 (N_2383,N_1635,N_1605);
and U2384 (N_2384,N_1617,N_1832);
nor U2385 (N_2385,N_1914,N_1638);
or U2386 (N_2386,N_1742,N_1970);
xor U2387 (N_2387,N_1948,N_1885);
nand U2388 (N_2388,N_1533,N_1672);
nand U2389 (N_2389,N_1891,N_1836);
and U2390 (N_2390,N_1884,N_1582);
or U2391 (N_2391,N_1847,N_1721);
and U2392 (N_2392,N_1861,N_1950);
nor U2393 (N_2393,N_1507,N_1627);
nor U2394 (N_2394,N_1620,N_1924);
or U2395 (N_2395,N_1551,N_1910);
xor U2396 (N_2396,N_1811,N_1561);
nor U2397 (N_2397,N_1652,N_1873);
and U2398 (N_2398,N_1803,N_1711);
and U2399 (N_2399,N_1949,N_1591);
and U2400 (N_2400,N_1911,N_1687);
nor U2401 (N_2401,N_1967,N_1521);
and U2402 (N_2402,N_1665,N_1791);
xor U2403 (N_2403,N_1992,N_1991);
nand U2404 (N_2404,N_1753,N_1599);
nand U2405 (N_2405,N_1663,N_1515);
or U2406 (N_2406,N_1766,N_1920);
or U2407 (N_2407,N_1835,N_1704);
nor U2408 (N_2408,N_1627,N_1585);
nand U2409 (N_2409,N_1625,N_1662);
nand U2410 (N_2410,N_1740,N_1563);
nand U2411 (N_2411,N_1882,N_1902);
nand U2412 (N_2412,N_1793,N_1604);
nand U2413 (N_2413,N_1699,N_1657);
or U2414 (N_2414,N_1540,N_1957);
or U2415 (N_2415,N_1805,N_1597);
nand U2416 (N_2416,N_1728,N_1851);
nand U2417 (N_2417,N_1905,N_1694);
xor U2418 (N_2418,N_1514,N_1726);
and U2419 (N_2419,N_1891,N_1844);
or U2420 (N_2420,N_1804,N_1628);
or U2421 (N_2421,N_1980,N_1773);
nand U2422 (N_2422,N_1994,N_1626);
or U2423 (N_2423,N_1616,N_1774);
and U2424 (N_2424,N_1785,N_1534);
nand U2425 (N_2425,N_1882,N_1813);
or U2426 (N_2426,N_1988,N_1901);
nand U2427 (N_2427,N_1616,N_1747);
and U2428 (N_2428,N_1581,N_1615);
and U2429 (N_2429,N_1652,N_1747);
nand U2430 (N_2430,N_1956,N_1537);
or U2431 (N_2431,N_1729,N_1807);
nor U2432 (N_2432,N_1980,N_1984);
or U2433 (N_2433,N_1600,N_1763);
nor U2434 (N_2434,N_1699,N_1901);
nand U2435 (N_2435,N_1586,N_1547);
nor U2436 (N_2436,N_1725,N_1616);
and U2437 (N_2437,N_1920,N_1767);
and U2438 (N_2438,N_1625,N_1572);
or U2439 (N_2439,N_1980,N_1615);
and U2440 (N_2440,N_1684,N_1649);
xor U2441 (N_2441,N_1721,N_1733);
and U2442 (N_2442,N_1918,N_1658);
nand U2443 (N_2443,N_1950,N_1740);
and U2444 (N_2444,N_1802,N_1551);
nand U2445 (N_2445,N_1822,N_1560);
or U2446 (N_2446,N_1890,N_1523);
nand U2447 (N_2447,N_1953,N_1786);
nor U2448 (N_2448,N_1740,N_1907);
or U2449 (N_2449,N_1837,N_1880);
nor U2450 (N_2450,N_1652,N_1646);
and U2451 (N_2451,N_1877,N_1550);
and U2452 (N_2452,N_1570,N_1662);
nand U2453 (N_2453,N_1788,N_1688);
or U2454 (N_2454,N_1750,N_1668);
and U2455 (N_2455,N_1966,N_1698);
and U2456 (N_2456,N_1690,N_1931);
and U2457 (N_2457,N_1993,N_1715);
or U2458 (N_2458,N_1815,N_1510);
nand U2459 (N_2459,N_1795,N_1881);
nand U2460 (N_2460,N_1959,N_1664);
or U2461 (N_2461,N_1890,N_1595);
nor U2462 (N_2462,N_1727,N_1838);
nor U2463 (N_2463,N_1661,N_1655);
or U2464 (N_2464,N_1661,N_1981);
nand U2465 (N_2465,N_1980,N_1538);
nor U2466 (N_2466,N_1873,N_1734);
nor U2467 (N_2467,N_1865,N_1562);
and U2468 (N_2468,N_1733,N_1918);
or U2469 (N_2469,N_1709,N_1759);
nand U2470 (N_2470,N_1757,N_1594);
or U2471 (N_2471,N_1565,N_1956);
nor U2472 (N_2472,N_1556,N_1574);
and U2473 (N_2473,N_1944,N_1889);
nand U2474 (N_2474,N_1594,N_1881);
or U2475 (N_2475,N_1646,N_1515);
and U2476 (N_2476,N_1888,N_1986);
nor U2477 (N_2477,N_1598,N_1606);
xnor U2478 (N_2478,N_1901,N_1714);
xnor U2479 (N_2479,N_1541,N_1960);
nor U2480 (N_2480,N_1820,N_1541);
nand U2481 (N_2481,N_1773,N_1889);
nand U2482 (N_2482,N_1857,N_1684);
nand U2483 (N_2483,N_1797,N_1840);
nor U2484 (N_2484,N_1544,N_1526);
nand U2485 (N_2485,N_1827,N_1907);
nand U2486 (N_2486,N_1528,N_1974);
nand U2487 (N_2487,N_1506,N_1948);
and U2488 (N_2488,N_1618,N_1757);
xor U2489 (N_2489,N_1775,N_1818);
nor U2490 (N_2490,N_1753,N_1879);
xnor U2491 (N_2491,N_1871,N_1666);
nor U2492 (N_2492,N_1646,N_1916);
and U2493 (N_2493,N_1823,N_1952);
and U2494 (N_2494,N_1623,N_1994);
or U2495 (N_2495,N_1603,N_1531);
nor U2496 (N_2496,N_1881,N_1809);
and U2497 (N_2497,N_1822,N_1793);
nor U2498 (N_2498,N_1762,N_1964);
nor U2499 (N_2499,N_1725,N_1713);
nand U2500 (N_2500,N_2460,N_2041);
or U2501 (N_2501,N_2065,N_2341);
nand U2502 (N_2502,N_2149,N_2194);
or U2503 (N_2503,N_2406,N_2461);
and U2504 (N_2504,N_2304,N_2383);
and U2505 (N_2505,N_2411,N_2221);
nor U2506 (N_2506,N_2392,N_2052);
nand U2507 (N_2507,N_2332,N_2315);
xnor U2508 (N_2508,N_2213,N_2000);
and U2509 (N_2509,N_2334,N_2366);
xnor U2510 (N_2510,N_2220,N_2265);
and U2511 (N_2511,N_2437,N_2188);
nor U2512 (N_2512,N_2124,N_2358);
and U2513 (N_2513,N_2039,N_2011);
nand U2514 (N_2514,N_2360,N_2009);
or U2515 (N_2515,N_2307,N_2320);
nand U2516 (N_2516,N_2174,N_2339);
nand U2517 (N_2517,N_2270,N_2291);
xnor U2518 (N_2518,N_2131,N_2138);
nor U2519 (N_2519,N_2072,N_2473);
nor U2520 (N_2520,N_2378,N_2365);
nand U2521 (N_2521,N_2495,N_2431);
nand U2522 (N_2522,N_2099,N_2491);
or U2523 (N_2523,N_2081,N_2187);
nand U2524 (N_2524,N_2349,N_2104);
nor U2525 (N_2525,N_2295,N_2191);
nor U2526 (N_2526,N_2274,N_2425);
or U2527 (N_2527,N_2494,N_2238);
or U2528 (N_2528,N_2248,N_2449);
or U2529 (N_2529,N_2147,N_2323);
nand U2530 (N_2530,N_2035,N_2372);
nand U2531 (N_2531,N_2397,N_2088);
nor U2532 (N_2532,N_2227,N_2250);
or U2533 (N_2533,N_2199,N_2350);
or U2534 (N_2534,N_2002,N_2245);
or U2535 (N_2535,N_2169,N_2239);
and U2536 (N_2536,N_2448,N_2243);
or U2537 (N_2537,N_2217,N_2017);
and U2538 (N_2538,N_2288,N_2290);
and U2539 (N_2539,N_2389,N_2167);
nor U2540 (N_2540,N_2413,N_2278);
nand U2541 (N_2541,N_2393,N_2443);
nor U2542 (N_2542,N_2381,N_2314);
or U2543 (N_2543,N_2159,N_2402);
and U2544 (N_2544,N_2456,N_2216);
xnor U2545 (N_2545,N_2478,N_2135);
or U2546 (N_2546,N_2019,N_2020);
and U2547 (N_2547,N_2340,N_2190);
nor U2548 (N_2548,N_2309,N_2060);
nand U2549 (N_2549,N_2403,N_2094);
nand U2550 (N_2550,N_2369,N_2244);
nand U2551 (N_2551,N_2271,N_2166);
or U2552 (N_2552,N_2076,N_2022);
and U2553 (N_2553,N_2045,N_2370);
or U2554 (N_2554,N_2260,N_2102);
and U2555 (N_2555,N_2367,N_2162);
nand U2556 (N_2556,N_2419,N_2241);
nor U2557 (N_2557,N_2001,N_2294);
or U2558 (N_2558,N_2204,N_2405);
nand U2559 (N_2559,N_2132,N_2298);
nand U2560 (N_2560,N_2115,N_2096);
nor U2561 (N_2561,N_2127,N_2352);
or U2562 (N_2562,N_2480,N_2106);
or U2563 (N_2563,N_2119,N_2417);
nand U2564 (N_2564,N_2142,N_2273);
nor U2565 (N_2565,N_2027,N_2496);
nor U2566 (N_2566,N_2141,N_2123);
nor U2567 (N_2567,N_2388,N_2459);
and U2568 (N_2568,N_2353,N_2414);
nor U2569 (N_2569,N_2212,N_2242);
nand U2570 (N_2570,N_2037,N_2329);
nand U2571 (N_2571,N_2322,N_2319);
xnor U2572 (N_2572,N_2256,N_2058);
nor U2573 (N_2573,N_2268,N_2318);
nand U2574 (N_2574,N_2005,N_2021);
and U2575 (N_2575,N_2264,N_2292);
and U2576 (N_2576,N_2454,N_2423);
nor U2577 (N_2577,N_2283,N_2084);
or U2578 (N_2578,N_2053,N_2144);
or U2579 (N_2579,N_2497,N_2492);
and U2580 (N_2580,N_2198,N_2408);
nand U2581 (N_2581,N_2089,N_2136);
nand U2582 (N_2582,N_2368,N_2062);
nand U2583 (N_2583,N_2409,N_2145);
or U2584 (N_2584,N_2028,N_2252);
or U2585 (N_2585,N_2087,N_2276);
nor U2586 (N_2586,N_2003,N_2433);
nand U2587 (N_2587,N_2156,N_2071);
and U2588 (N_2588,N_2297,N_2015);
nor U2589 (N_2589,N_2176,N_2181);
nor U2590 (N_2590,N_2371,N_2308);
xnor U2591 (N_2591,N_2462,N_2237);
xor U2592 (N_2592,N_2385,N_2412);
nand U2593 (N_2593,N_2168,N_2476);
or U2594 (N_2594,N_2063,N_2157);
and U2595 (N_2595,N_2343,N_2185);
or U2596 (N_2596,N_2184,N_2356);
nor U2597 (N_2597,N_2057,N_2434);
nand U2598 (N_2598,N_2200,N_2224);
nand U2599 (N_2599,N_2186,N_2023);
or U2600 (N_2600,N_2122,N_2208);
nor U2601 (N_2601,N_2316,N_2386);
or U2602 (N_2602,N_2326,N_2090);
nand U2603 (N_2603,N_2183,N_2078);
and U2604 (N_2604,N_2346,N_2007);
nor U2605 (N_2605,N_2344,N_2055);
or U2606 (N_2606,N_2296,N_2266);
or U2607 (N_2607,N_2435,N_2333);
xnor U2608 (N_2608,N_2391,N_2446);
nand U2609 (N_2609,N_2463,N_2455);
or U2610 (N_2610,N_2285,N_2038);
and U2611 (N_2611,N_2482,N_2233);
and U2612 (N_2612,N_2355,N_2487);
or U2613 (N_2613,N_2148,N_2440);
nand U2614 (N_2614,N_2107,N_2254);
and U2615 (N_2615,N_2086,N_2032);
nor U2616 (N_2616,N_2228,N_2486);
and U2617 (N_2617,N_2010,N_2428);
nor U2618 (N_2618,N_2301,N_2125);
nand U2619 (N_2619,N_2044,N_2080);
nor U2620 (N_2620,N_2240,N_2493);
nor U2621 (N_2621,N_2429,N_2430);
or U2622 (N_2622,N_2061,N_2120);
and U2623 (N_2623,N_2114,N_2117);
nand U2624 (N_2624,N_2049,N_2261);
nand U2625 (N_2625,N_2215,N_2281);
and U2626 (N_2626,N_2453,N_2130);
or U2627 (N_2627,N_2426,N_2277);
nor U2628 (N_2628,N_2209,N_2279);
nand U2629 (N_2629,N_2040,N_2140);
nand U2630 (N_2630,N_2253,N_2267);
or U2631 (N_2631,N_2470,N_2085);
and U2632 (N_2632,N_2490,N_2012);
nor U2633 (N_2633,N_2236,N_2287);
or U2634 (N_2634,N_2471,N_2154);
and U2635 (N_2635,N_2342,N_2093);
nor U2636 (N_2636,N_2070,N_2300);
nand U2637 (N_2637,N_2442,N_2311);
and U2638 (N_2638,N_2146,N_2247);
nor U2639 (N_2639,N_2205,N_2054);
xnor U2640 (N_2640,N_2262,N_2079);
nor U2641 (N_2641,N_2373,N_2394);
nand U2642 (N_2642,N_2110,N_2137);
nor U2643 (N_2643,N_2016,N_2445);
nand U2644 (N_2644,N_2293,N_2231);
nor U2645 (N_2645,N_2375,N_2230);
nor U2646 (N_2646,N_2282,N_2284);
or U2647 (N_2647,N_2014,N_2427);
nor U2648 (N_2648,N_2150,N_2303);
nand U2649 (N_2649,N_2472,N_2073);
and U2650 (N_2650,N_2031,N_2347);
nand U2651 (N_2651,N_2152,N_2330);
nand U2652 (N_2652,N_2483,N_2421);
nand U2653 (N_2653,N_2474,N_2203);
or U2654 (N_2654,N_2064,N_2111);
and U2655 (N_2655,N_2398,N_2348);
or U2656 (N_2656,N_2499,N_2118);
or U2657 (N_2657,N_2207,N_2218);
or U2658 (N_2658,N_2112,N_2100);
and U2659 (N_2659,N_2202,N_2180);
nor U2660 (N_2660,N_2128,N_2451);
and U2661 (N_2661,N_2321,N_2404);
nand U2662 (N_2662,N_2206,N_2259);
nor U2663 (N_2663,N_2336,N_2195);
xnor U2664 (N_2664,N_2489,N_2488);
and U2665 (N_2665,N_2139,N_2395);
nor U2666 (N_2666,N_2382,N_2179);
nor U2667 (N_2667,N_2477,N_2197);
nand U2668 (N_2668,N_2351,N_2165);
nor U2669 (N_2669,N_2407,N_2075);
and U2670 (N_2670,N_2438,N_2312);
and U2671 (N_2671,N_2313,N_2173);
and U2672 (N_2672,N_2095,N_2143);
and U2673 (N_2673,N_2286,N_2498);
or U2674 (N_2674,N_2177,N_2068);
or U2675 (N_2675,N_2067,N_2222);
nor U2676 (N_2676,N_2467,N_2105);
and U2677 (N_2677,N_2251,N_2401);
and U2678 (N_2678,N_2004,N_2468);
and U2679 (N_2679,N_2246,N_2317);
xor U2680 (N_2680,N_2066,N_2121);
nand U2681 (N_2681,N_2331,N_2214);
nor U2682 (N_2682,N_2447,N_2289);
and U2683 (N_2683,N_2424,N_2439);
nor U2684 (N_2684,N_2361,N_2432);
and U2685 (N_2685,N_2335,N_2153);
nand U2686 (N_2686,N_2160,N_2229);
xnor U2687 (N_2687,N_2310,N_2376);
nor U2688 (N_2688,N_2384,N_2097);
nor U2689 (N_2689,N_2327,N_2013);
or U2690 (N_2690,N_2475,N_2164);
nand U2691 (N_2691,N_2219,N_2420);
nand U2692 (N_2692,N_2302,N_2299);
nor U2693 (N_2693,N_2324,N_2379);
nand U2694 (N_2694,N_2034,N_2481);
or U2695 (N_2695,N_2363,N_2091);
and U2696 (N_2696,N_2196,N_2235);
or U2697 (N_2697,N_2056,N_2042);
or U2698 (N_2698,N_2026,N_2211);
nand U2699 (N_2699,N_2484,N_2345);
or U2700 (N_2700,N_2018,N_2029);
and U2701 (N_2701,N_2083,N_2024);
or U2702 (N_2702,N_2410,N_2452);
or U2703 (N_2703,N_2255,N_2006);
or U2704 (N_2704,N_2101,N_2306);
xor U2705 (N_2705,N_2399,N_2458);
nand U2706 (N_2706,N_2390,N_2047);
or U2707 (N_2707,N_2077,N_2082);
or U2708 (N_2708,N_2325,N_2436);
or U2709 (N_2709,N_2465,N_2129);
nor U2710 (N_2710,N_2036,N_2133);
nor U2711 (N_2711,N_2280,N_2364);
nor U2712 (N_2712,N_2134,N_2171);
xnor U2713 (N_2713,N_2485,N_2172);
and U2714 (N_2714,N_2048,N_2441);
xnor U2715 (N_2715,N_2362,N_2464);
nand U2716 (N_2716,N_2210,N_2069);
and U2717 (N_2717,N_2354,N_2151);
and U2718 (N_2718,N_2444,N_2377);
nand U2719 (N_2719,N_2074,N_2103);
xor U2720 (N_2720,N_2051,N_2008);
or U2721 (N_2721,N_2466,N_2415);
or U2722 (N_2722,N_2257,N_2025);
and U2723 (N_2723,N_2226,N_2046);
xnor U2724 (N_2724,N_2108,N_2182);
xnor U2725 (N_2725,N_2050,N_2201);
or U2726 (N_2726,N_2113,N_2030);
nand U2727 (N_2727,N_2234,N_2396);
and U2728 (N_2728,N_2457,N_2374);
xnor U2729 (N_2729,N_2043,N_2450);
nor U2730 (N_2730,N_2357,N_2223);
nand U2731 (N_2731,N_2338,N_2175);
and U2732 (N_2732,N_2269,N_2249);
and U2733 (N_2733,N_2098,N_2418);
nor U2734 (N_2734,N_2422,N_2192);
or U2735 (N_2735,N_2126,N_2469);
nor U2736 (N_2736,N_2170,N_2387);
and U2737 (N_2737,N_2232,N_2033);
nand U2738 (N_2738,N_2328,N_2272);
and U2739 (N_2739,N_2305,N_2059);
or U2740 (N_2740,N_2158,N_2225);
nor U2741 (N_2741,N_2359,N_2400);
and U2742 (N_2742,N_2109,N_2275);
or U2743 (N_2743,N_2263,N_2189);
nor U2744 (N_2744,N_2479,N_2092);
xor U2745 (N_2745,N_2116,N_2380);
nor U2746 (N_2746,N_2163,N_2161);
or U2747 (N_2747,N_2193,N_2258);
nand U2748 (N_2748,N_2155,N_2337);
and U2749 (N_2749,N_2416,N_2178);
nand U2750 (N_2750,N_2253,N_2038);
xor U2751 (N_2751,N_2390,N_2054);
or U2752 (N_2752,N_2372,N_2437);
or U2753 (N_2753,N_2290,N_2306);
or U2754 (N_2754,N_2269,N_2222);
xor U2755 (N_2755,N_2422,N_2098);
or U2756 (N_2756,N_2408,N_2175);
and U2757 (N_2757,N_2195,N_2210);
or U2758 (N_2758,N_2454,N_2269);
nand U2759 (N_2759,N_2033,N_2011);
and U2760 (N_2760,N_2176,N_2191);
and U2761 (N_2761,N_2043,N_2088);
and U2762 (N_2762,N_2267,N_2410);
nor U2763 (N_2763,N_2294,N_2363);
or U2764 (N_2764,N_2170,N_2084);
and U2765 (N_2765,N_2459,N_2314);
nand U2766 (N_2766,N_2296,N_2374);
and U2767 (N_2767,N_2336,N_2012);
or U2768 (N_2768,N_2424,N_2071);
and U2769 (N_2769,N_2375,N_2179);
and U2770 (N_2770,N_2103,N_2326);
or U2771 (N_2771,N_2476,N_2159);
and U2772 (N_2772,N_2300,N_2117);
or U2773 (N_2773,N_2302,N_2124);
or U2774 (N_2774,N_2289,N_2089);
and U2775 (N_2775,N_2457,N_2085);
nor U2776 (N_2776,N_2492,N_2379);
xor U2777 (N_2777,N_2284,N_2421);
nand U2778 (N_2778,N_2388,N_2291);
and U2779 (N_2779,N_2135,N_2239);
or U2780 (N_2780,N_2296,N_2001);
nor U2781 (N_2781,N_2064,N_2280);
nand U2782 (N_2782,N_2142,N_2090);
nor U2783 (N_2783,N_2092,N_2270);
xor U2784 (N_2784,N_2070,N_2469);
nor U2785 (N_2785,N_2113,N_2174);
nand U2786 (N_2786,N_2262,N_2385);
or U2787 (N_2787,N_2103,N_2075);
nor U2788 (N_2788,N_2072,N_2073);
and U2789 (N_2789,N_2264,N_2282);
and U2790 (N_2790,N_2198,N_2030);
and U2791 (N_2791,N_2202,N_2472);
xor U2792 (N_2792,N_2028,N_2031);
and U2793 (N_2793,N_2214,N_2279);
xnor U2794 (N_2794,N_2172,N_2135);
and U2795 (N_2795,N_2462,N_2324);
nand U2796 (N_2796,N_2070,N_2056);
nor U2797 (N_2797,N_2316,N_2326);
or U2798 (N_2798,N_2036,N_2106);
nand U2799 (N_2799,N_2489,N_2106);
or U2800 (N_2800,N_2307,N_2285);
nor U2801 (N_2801,N_2432,N_2446);
nor U2802 (N_2802,N_2413,N_2362);
nand U2803 (N_2803,N_2062,N_2195);
nand U2804 (N_2804,N_2258,N_2237);
or U2805 (N_2805,N_2191,N_2151);
and U2806 (N_2806,N_2103,N_2220);
nand U2807 (N_2807,N_2321,N_2415);
nor U2808 (N_2808,N_2291,N_2159);
nand U2809 (N_2809,N_2140,N_2387);
xnor U2810 (N_2810,N_2344,N_2486);
nor U2811 (N_2811,N_2492,N_2420);
xnor U2812 (N_2812,N_2414,N_2379);
nor U2813 (N_2813,N_2130,N_2399);
xor U2814 (N_2814,N_2128,N_2358);
and U2815 (N_2815,N_2053,N_2119);
or U2816 (N_2816,N_2055,N_2334);
nor U2817 (N_2817,N_2389,N_2229);
and U2818 (N_2818,N_2110,N_2431);
and U2819 (N_2819,N_2370,N_2357);
nor U2820 (N_2820,N_2052,N_2179);
xnor U2821 (N_2821,N_2430,N_2155);
xnor U2822 (N_2822,N_2300,N_2036);
or U2823 (N_2823,N_2075,N_2285);
nand U2824 (N_2824,N_2377,N_2422);
nand U2825 (N_2825,N_2444,N_2003);
and U2826 (N_2826,N_2462,N_2381);
and U2827 (N_2827,N_2039,N_2456);
or U2828 (N_2828,N_2366,N_2438);
nand U2829 (N_2829,N_2173,N_2126);
nand U2830 (N_2830,N_2276,N_2027);
or U2831 (N_2831,N_2199,N_2204);
and U2832 (N_2832,N_2181,N_2360);
nor U2833 (N_2833,N_2174,N_2178);
or U2834 (N_2834,N_2036,N_2143);
and U2835 (N_2835,N_2389,N_2005);
or U2836 (N_2836,N_2073,N_2453);
and U2837 (N_2837,N_2437,N_2363);
and U2838 (N_2838,N_2319,N_2367);
nand U2839 (N_2839,N_2270,N_2192);
and U2840 (N_2840,N_2155,N_2260);
nor U2841 (N_2841,N_2315,N_2297);
and U2842 (N_2842,N_2261,N_2246);
xnor U2843 (N_2843,N_2014,N_2439);
nand U2844 (N_2844,N_2085,N_2423);
nand U2845 (N_2845,N_2447,N_2151);
or U2846 (N_2846,N_2227,N_2440);
nor U2847 (N_2847,N_2402,N_2069);
or U2848 (N_2848,N_2424,N_2022);
and U2849 (N_2849,N_2249,N_2148);
nor U2850 (N_2850,N_2484,N_2057);
nand U2851 (N_2851,N_2131,N_2183);
nand U2852 (N_2852,N_2455,N_2434);
nor U2853 (N_2853,N_2309,N_2016);
xor U2854 (N_2854,N_2375,N_2110);
nor U2855 (N_2855,N_2278,N_2425);
nand U2856 (N_2856,N_2421,N_2013);
or U2857 (N_2857,N_2068,N_2018);
nand U2858 (N_2858,N_2239,N_2261);
or U2859 (N_2859,N_2450,N_2282);
nand U2860 (N_2860,N_2314,N_2062);
nand U2861 (N_2861,N_2493,N_2400);
nor U2862 (N_2862,N_2151,N_2277);
and U2863 (N_2863,N_2305,N_2110);
xor U2864 (N_2864,N_2452,N_2073);
or U2865 (N_2865,N_2017,N_2386);
xor U2866 (N_2866,N_2025,N_2473);
and U2867 (N_2867,N_2029,N_2165);
or U2868 (N_2868,N_2163,N_2282);
nor U2869 (N_2869,N_2240,N_2102);
and U2870 (N_2870,N_2471,N_2135);
xor U2871 (N_2871,N_2086,N_2216);
nand U2872 (N_2872,N_2206,N_2141);
or U2873 (N_2873,N_2443,N_2448);
or U2874 (N_2874,N_2299,N_2384);
nor U2875 (N_2875,N_2211,N_2448);
and U2876 (N_2876,N_2000,N_2390);
and U2877 (N_2877,N_2280,N_2367);
and U2878 (N_2878,N_2370,N_2437);
nand U2879 (N_2879,N_2220,N_2179);
nor U2880 (N_2880,N_2288,N_2260);
or U2881 (N_2881,N_2143,N_2196);
or U2882 (N_2882,N_2059,N_2482);
nor U2883 (N_2883,N_2499,N_2317);
or U2884 (N_2884,N_2404,N_2114);
xor U2885 (N_2885,N_2253,N_2206);
nor U2886 (N_2886,N_2498,N_2205);
and U2887 (N_2887,N_2160,N_2047);
or U2888 (N_2888,N_2204,N_2192);
or U2889 (N_2889,N_2389,N_2141);
and U2890 (N_2890,N_2356,N_2324);
and U2891 (N_2891,N_2038,N_2225);
or U2892 (N_2892,N_2139,N_2274);
or U2893 (N_2893,N_2353,N_2407);
nand U2894 (N_2894,N_2111,N_2304);
nor U2895 (N_2895,N_2409,N_2294);
nor U2896 (N_2896,N_2124,N_2381);
and U2897 (N_2897,N_2362,N_2393);
and U2898 (N_2898,N_2412,N_2160);
xor U2899 (N_2899,N_2046,N_2079);
or U2900 (N_2900,N_2497,N_2131);
nor U2901 (N_2901,N_2295,N_2404);
and U2902 (N_2902,N_2196,N_2247);
and U2903 (N_2903,N_2417,N_2025);
nand U2904 (N_2904,N_2329,N_2046);
and U2905 (N_2905,N_2447,N_2465);
and U2906 (N_2906,N_2370,N_2212);
nand U2907 (N_2907,N_2017,N_2008);
and U2908 (N_2908,N_2084,N_2092);
and U2909 (N_2909,N_2067,N_2367);
xnor U2910 (N_2910,N_2176,N_2475);
nor U2911 (N_2911,N_2021,N_2244);
and U2912 (N_2912,N_2484,N_2235);
or U2913 (N_2913,N_2092,N_2123);
and U2914 (N_2914,N_2322,N_2473);
and U2915 (N_2915,N_2469,N_2268);
nand U2916 (N_2916,N_2462,N_2150);
nor U2917 (N_2917,N_2361,N_2287);
and U2918 (N_2918,N_2005,N_2168);
xnor U2919 (N_2919,N_2042,N_2195);
nor U2920 (N_2920,N_2311,N_2409);
xnor U2921 (N_2921,N_2172,N_2053);
nor U2922 (N_2922,N_2256,N_2293);
nand U2923 (N_2923,N_2142,N_2454);
nand U2924 (N_2924,N_2122,N_2203);
and U2925 (N_2925,N_2401,N_2297);
nor U2926 (N_2926,N_2096,N_2324);
and U2927 (N_2927,N_2366,N_2091);
or U2928 (N_2928,N_2310,N_2168);
nand U2929 (N_2929,N_2273,N_2370);
and U2930 (N_2930,N_2295,N_2248);
xor U2931 (N_2931,N_2271,N_2344);
or U2932 (N_2932,N_2106,N_2422);
nor U2933 (N_2933,N_2322,N_2175);
nor U2934 (N_2934,N_2264,N_2459);
nor U2935 (N_2935,N_2476,N_2006);
and U2936 (N_2936,N_2196,N_2110);
and U2937 (N_2937,N_2236,N_2433);
and U2938 (N_2938,N_2085,N_2109);
nand U2939 (N_2939,N_2355,N_2444);
and U2940 (N_2940,N_2303,N_2492);
nand U2941 (N_2941,N_2382,N_2196);
nand U2942 (N_2942,N_2209,N_2021);
and U2943 (N_2943,N_2147,N_2273);
or U2944 (N_2944,N_2470,N_2302);
nor U2945 (N_2945,N_2453,N_2266);
xor U2946 (N_2946,N_2159,N_2171);
xor U2947 (N_2947,N_2001,N_2064);
nand U2948 (N_2948,N_2420,N_2097);
or U2949 (N_2949,N_2363,N_2280);
or U2950 (N_2950,N_2416,N_2131);
nand U2951 (N_2951,N_2378,N_2338);
nor U2952 (N_2952,N_2482,N_2080);
or U2953 (N_2953,N_2251,N_2222);
nand U2954 (N_2954,N_2282,N_2196);
nand U2955 (N_2955,N_2408,N_2360);
and U2956 (N_2956,N_2293,N_2198);
or U2957 (N_2957,N_2185,N_2149);
and U2958 (N_2958,N_2041,N_2245);
or U2959 (N_2959,N_2451,N_2249);
nor U2960 (N_2960,N_2398,N_2155);
nor U2961 (N_2961,N_2385,N_2311);
or U2962 (N_2962,N_2128,N_2064);
nor U2963 (N_2963,N_2199,N_2464);
and U2964 (N_2964,N_2235,N_2138);
or U2965 (N_2965,N_2151,N_2027);
nor U2966 (N_2966,N_2377,N_2011);
xnor U2967 (N_2967,N_2311,N_2148);
nor U2968 (N_2968,N_2252,N_2231);
xor U2969 (N_2969,N_2445,N_2181);
or U2970 (N_2970,N_2484,N_2245);
nor U2971 (N_2971,N_2338,N_2235);
nor U2972 (N_2972,N_2267,N_2467);
or U2973 (N_2973,N_2303,N_2350);
xnor U2974 (N_2974,N_2427,N_2340);
and U2975 (N_2975,N_2011,N_2458);
nor U2976 (N_2976,N_2272,N_2408);
nand U2977 (N_2977,N_2044,N_2473);
or U2978 (N_2978,N_2153,N_2267);
nand U2979 (N_2979,N_2267,N_2462);
or U2980 (N_2980,N_2437,N_2305);
or U2981 (N_2981,N_2300,N_2146);
nand U2982 (N_2982,N_2197,N_2261);
nand U2983 (N_2983,N_2498,N_2010);
and U2984 (N_2984,N_2078,N_2115);
nor U2985 (N_2985,N_2394,N_2066);
and U2986 (N_2986,N_2399,N_2179);
nand U2987 (N_2987,N_2055,N_2261);
and U2988 (N_2988,N_2393,N_2016);
nand U2989 (N_2989,N_2108,N_2125);
or U2990 (N_2990,N_2045,N_2330);
nand U2991 (N_2991,N_2097,N_2418);
nand U2992 (N_2992,N_2476,N_2066);
nor U2993 (N_2993,N_2117,N_2205);
or U2994 (N_2994,N_2291,N_2481);
and U2995 (N_2995,N_2184,N_2261);
or U2996 (N_2996,N_2095,N_2478);
and U2997 (N_2997,N_2060,N_2233);
and U2998 (N_2998,N_2000,N_2009);
xnor U2999 (N_2999,N_2290,N_2197);
xnor U3000 (N_3000,N_2659,N_2861);
nand U3001 (N_3001,N_2556,N_2757);
xnor U3002 (N_3002,N_2763,N_2751);
and U3003 (N_3003,N_2571,N_2777);
nor U3004 (N_3004,N_2838,N_2525);
xnor U3005 (N_3005,N_2543,N_2917);
or U3006 (N_3006,N_2611,N_2669);
or U3007 (N_3007,N_2947,N_2626);
nand U3008 (N_3008,N_2889,N_2969);
or U3009 (N_3009,N_2656,N_2736);
nor U3010 (N_3010,N_2743,N_2651);
and U3011 (N_3011,N_2649,N_2899);
and U3012 (N_3012,N_2738,N_2828);
and U3013 (N_3013,N_2805,N_2692);
nand U3014 (N_3014,N_2912,N_2622);
nor U3015 (N_3015,N_2689,N_2982);
and U3016 (N_3016,N_2764,N_2939);
nor U3017 (N_3017,N_2923,N_2699);
nor U3018 (N_3018,N_2740,N_2636);
nor U3019 (N_3019,N_2986,N_2895);
xor U3020 (N_3020,N_2867,N_2635);
xor U3021 (N_3021,N_2882,N_2795);
and U3022 (N_3022,N_2517,N_2682);
and U3023 (N_3023,N_2501,N_2521);
nand U3024 (N_3024,N_2594,N_2700);
nor U3025 (N_3025,N_2715,N_2579);
and U3026 (N_3026,N_2625,N_2948);
nand U3027 (N_3027,N_2825,N_2730);
nor U3028 (N_3028,N_2788,N_2811);
and U3029 (N_3029,N_2835,N_2584);
and U3030 (N_3030,N_2978,N_2914);
nor U3031 (N_3031,N_2507,N_2879);
or U3032 (N_3032,N_2735,N_2902);
nand U3033 (N_3033,N_2870,N_2657);
nor U3034 (N_3034,N_2619,N_2799);
xor U3035 (N_3035,N_2675,N_2865);
xnor U3036 (N_3036,N_2845,N_2863);
xor U3037 (N_3037,N_2816,N_2710);
xnor U3038 (N_3038,N_2990,N_2557);
nand U3039 (N_3039,N_2970,N_2809);
nor U3040 (N_3040,N_2620,N_2893);
nor U3041 (N_3041,N_2972,N_2908);
nor U3042 (N_3042,N_2952,N_2536);
nand U3043 (N_3043,N_2667,N_2672);
or U3044 (N_3044,N_2734,N_2903);
xnor U3045 (N_3045,N_2820,N_2938);
and U3046 (N_3046,N_2529,N_2823);
nand U3047 (N_3047,N_2508,N_2964);
or U3048 (N_3048,N_2563,N_2989);
and U3049 (N_3049,N_2997,N_2968);
nor U3050 (N_3050,N_2916,N_2790);
nor U3051 (N_3051,N_2802,N_2909);
nand U3052 (N_3052,N_2642,N_2897);
xnor U3053 (N_3053,N_2604,N_2535);
or U3054 (N_3054,N_2711,N_2609);
nor U3055 (N_3055,N_2505,N_2780);
or U3056 (N_3056,N_2506,N_2639);
nand U3057 (N_3057,N_2509,N_2515);
nand U3058 (N_3058,N_2630,N_2588);
or U3059 (N_3059,N_2684,N_2567);
and U3060 (N_3060,N_2974,N_2851);
nand U3061 (N_3061,N_2878,N_2927);
and U3062 (N_3062,N_2668,N_2576);
nand U3063 (N_3063,N_2663,N_2920);
or U3064 (N_3064,N_2518,N_2648);
or U3065 (N_3065,N_2856,N_2800);
nor U3066 (N_3066,N_2600,N_2558);
nor U3067 (N_3067,N_2717,N_2991);
nor U3068 (N_3068,N_2652,N_2599);
or U3069 (N_3069,N_2634,N_2841);
nand U3070 (N_3070,N_2842,N_2704);
and U3071 (N_3071,N_2775,N_2686);
and U3072 (N_3072,N_2713,N_2707);
and U3073 (N_3073,N_2754,N_2866);
and U3074 (N_3074,N_2729,N_2971);
nor U3075 (N_3075,N_2615,N_2725);
or U3076 (N_3076,N_2608,N_2546);
nor U3077 (N_3077,N_2712,N_2834);
and U3078 (N_3078,N_2674,N_2796);
or U3079 (N_3079,N_2943,N_2647);
or U3080 (N_3080,N_2539,N_2907);
nand U3081 (N_3081,N_2748,N_2690);
xor U3082 (N_3082,N_2637,N_2847);
nor U3083 (N_3083,N_2698,N_2540);
or U3084 (N_3084,N_2922,N_2808);
or U3085 (N_3085,N_2880,N_2658);
or U3086 (N_3086,N_2665,N_2771);
nand U3087 (N_3087,N_2602,N_2785);
and U3088 (N_3088,N_2919,N_2618);
nor U3089 (N_3089,N_2791,N_2854);
nand U3090 (N_3090,N_2770,N_2614);
nand U3091 (N_3091,N_2901,N_2522);
nand U3092 (N_3092,N_2766,N_2623);
and U3093 (N_3093,N_2818,N_2601);
nand U3094 (N_3094,N_2941,N_2554);
nand U3095 (N_3095,N_2678,N_2890);
nor U3096 (N_3096,N_2987,N_2593);
nor U3097 (N_3097,N_2701,N_2877);
or U3098 (N_3098,N_2531,N_2732);
nor U3099 (N_3099,N_2679,N_2580);
and U3100 (N_3100,N_2650,N_2504);
and U3101 (N_3101,N_2998,N_2570);
or U3102 (N_3102,N_2703,N_2512);
nand U3103 (N_3103,N_2774,N_2560);
or U3104 (N_3104,N_2849,N_2883);
xnor U3105 (N_3105,N_2822,N_2526);
or U3106 (N_3106,N_2610,N_2681);
nor U3107 (N_3107,N_2896,N_2961);
nor U3108 (N_3108,N_2804,N_2850);
nor U3109 (N_3109,N_2644,N_2924);
and U3110 (N_3110,N_2653,N_2886);
or U3111 (N_3111,N_2815,N_2769);
nand U3112 (N_3112,N_2597,N_2731);
or U3113 (N_3113,N_2733,N_2551);
nor U3114 (N_3114,N_2801,N_2846);
and U3115 (N_3115,N_2613,N_2930);
or U3116 (N_3116,N_2942,N_2607);
nor U3117 (N_3117,N_2817,N_2953);
and U3118 (N_3118,N_2836,N_2513);
xor U3119 (N_3119,N_2705,N_2843);
xor U3120 (N_3120,N_2829,N_2857);
or U3121 (N_3121,N_2789,N_2862);
and U3122 (N_3122,N_2624,N_2528);
nor U3123 (N_3123,N_2918,N_2562);
nand U3124 (N_3124,N_2661,N_2821);
or U3125 (N_3125,N_2633,N_2537);
nor U3126 (N_3126,N_2547,N_2932);
nor U3127 (N_3127,N_2812,N_2956);
nor U3128 (N_3128,N_2577,N_2632);
nor U3129 (N_3129,N_2612,N_2868);
nand U3130 (N_3130,N_2758,N_2853);
or U3131 (N_3131,N_2848,N_2519);
nor U3132 (N_3132,N_2510,N_2544);
nand U3133 (N_3133,N_2944,N_2793);
or U3134 (N_3134,N_2747,N_2995);
nand U3135 (N_3135,N_2871,N_2545);
and U3136 (N_3136,N_2589,N_2827);
xor U3137 (N_3137,N_2858,N_2831);
nor U3138 (N_3138,N_2586,N_2581);
nor U3139 (N_3139,N_2977,N_2727);
xnor U3140 (N_3140,N_2931,N_2530);
nor U3141 (N_3141,N_2864,N_2915);
or U3142 (N_3142,N_2646,N_2814);
nand U3143 (N_3143,N_2739,N_2685);
and U3144 (N_3144,N_2561,N_2984);
nand U3145 (N_3145,N_2884,N_2532);
or U3146 (N_3146,N_2975,N_2959);
or U3147 (N_3147,N_2683,N_2603);
nor U3148 (N_3148,N_2994,N_2832);
or U3149 (N_3149,N_2660,N_2755);
nor U3150 (N_3150,N_2677,N_2583);
xnor U3151 (N_3151,N_2552,N_2750);
and U3152 (N_3152,N_2533,N_2824);
xnor U3153 (N_3153,N_2979,N_2794);
nor U3154 (N_3154,N_2721,N_2541);
or U3155 (N_3155,N_2759,N_2980);
xor U3156 (N_3156,N_2773,N_2892);
nor U3157 (N_3157,N_2728,N_2502);
xnor U3158 (N_3158,N_2524,N_2957);
nand U3159 (N_3159,N_2662,N_2925);
or U3160 (N_3160,N_2905,N_2792);
nor U3161 (N_3161,N_2582,N_2673);
or U3162 (N_3162,N_2676,N_2641);
xor U3163 (N_3163,N_2745,N_2714);
nor U3164 (N_3164,N_2573,N_2640);
or U3165 (N_3165,N_2840,N_2960);
nor U3166 (N_3166,N_2873,N_2963);
nor U3167 (N_3167,N_2687,N_2949);
nand U3168 (N_3168,N_2926,N_2569);
or U3169 (N_3169,N_2876,N_2904);
nand U3170 (N_3170,N_2523,N_2578);
nor U3171 (N_3171,N_2783,N_2753);
or U3172 (N_3172,N_2940,N_2776);
nor U3173 (N_3173,N_2538,N_2720);
nand U3174 (N_3174,N_2726,N_2937);
and U3175 (N_3175,N_2559,N_2999);
and U3176 (N_3176,N_2629,N_2950);
or U3177 (N_3177,N_2967,N_2706);
and U3178 (N_3178,N_2810,N_2621);
nor U3179 (N_3179,N_2976,N_2973);
nand U3180 (N_3180,N_2722,N_2671);
or U3181 (N_3181,N_2833,N_2761);
or U3182 (N_3182,N_2590,N_2881);
nor U3183 (N_3183,N_2844,N_2936);
nor U3184 (N_3184,N_2894,N_2591);
or U3185 (N_3185,N_2830,N_2962);
or U3186 (N_3186,N_2520,N_2500);
or U3187 (N_3187,N_2913,N_2911);
or U3188 (N_3188,N_2781,N_2988);
nand U3189 (N_3189,N_2826,N_2813);
or U3190 (N_3190,N_2741,N_2724);
and U3191 (N_3191,N_2768,N_2598);
nand U3192 (N_3192,N_2954,N_2587);
and U3193 (N_3193,N_2951,N_2568);
or U3194 (N_3194,N_2885,N_2534);
nor U3195 (N_3195,N_2906,N_2859);
nand U3196 (N_3196,N_2549,N_2806);
nand U3197 (N_3197,N_2869,N_2566);
and U3198 (N_3198,N_2888,N_2746);
and U3199 (N_3199,N_2803,N_2616);
or U3200 (N_3200,N_2898,N_2933);
and U3201 (N_3201,N_2742,N_2565);
nor U3202 (N_3202,N_2955,N_2585);
or U3203 (N_3203,N_2553,N_2935);
or U3204 (N_3204,N_2575,N_2511);
xnor U3205 (N_3205,N_2807,N_2670);
nor U3206 (N_3206,N_2574,N_2654);
xor U3207 (N_3207,N_2680,N_2592);
nand U3208 (N_3208,N_2737,N_2837);
nand U3209 (N_3209,N_2860,N_2928);
nor U3210 (N_3210,N_2550,N_2718);
nand U3211 (N_3211,N_2772,N_2645);
or U3212 (N_3212,N_2782,N_2762);
nor U3213 (N_3213,N_2983,N_2910);
or U3214 (N_3214,N_2631,N_2760);
or U3215 (N_3215,N_2697,N_2852);
and U3216 (N_3216,N_2744,N_2752);
nand U3217 (N_3217,N_2688,N_2992);
xor U3218 (N_3218,N_2542,N_2784);
nor U3219 (N_3219,N_2617,N_2946);
or U3220 (N_3220,N_2875,N_2719);
or U3221 (N_3221,N_2708,N_2765);
nor U3222 (N_3222,N_2985,N_2514);
or U3223 (N_3223,N_2767,N_2945);
nor U3224 (N_3224,N_2628,N_2605);
nand U3225 (N_3225,N_2934,N_2516);
and U3226 (N_3226,N_2643,N_2694);
nor U3227 (N_3227,N_2716,N_2655);
and U3228 (N_3228,N_2756,N_2993);
nand U3229 (N_3229,N_2749,N_2779);
or U3230 (N_3230,N_2797,N_2702);
nor U3231 (N_3231,N_2891,N_2723);
nor U3232 (N_3232,N_2595,N_2596);
and U3233 (N_3233,N_2958,N_2564);
and U3234 (N_3234,N_2929,N_2798);
nor U3235 (N_3235,N_2696,N_2503);
xnor U3236 (N_3236,N_2709,N_2887);
and U3237 (N_3237,N_2555,N_2787);
or U3238 (N_3238,N_2981,N_2572);
nand U3239 (N_3239,N_2921,N_2606);
or U3240 (N_3240,N_2872,N_2627);
xor U3241 (N_3241,N_2839,N_2855);
or U3242 (N_3242,N_2664,N_2638);
nor U3243 (N_3243,N_2786,N_2527);
or U3244 (N_3244,N_2666,N_2996);
and U3245 (N_3245,N_2900,N_2691);
or U3246 (N_3246,N_2778,N_2548);
nor U3247 (N_3247,N_2966,N_2695);
xor U3248 (N_3248,N_2819,N_2693);
or U3249 (N_3249,N_2965,N_2874);
or U3250 (N_3250,N_2862,N_2513);
and U3251 (N_3251,N_2864,N_2824);
or U3252 (N_3252,N_2717,N_2941);
and U3253 (N_3253,N_2893,N_2859);
and U3254 (N_3254,N_2608,N_2797);
nor U3255 (N_3255,N_2798,N_2590);
and U3256 (N_3256,N_2929,N_2519);
xor U3257 (N_3257,N_2562,N_2961);
nand U3258 (N_3258,N_2737,N_2945);
or U3259 (N_3259,N_2573,N_2662);
nand U3260 (N_3260,N_2584,N_2781);
and U3261 (N_3261,N_2873,N_2623);
xnor U3262 (N_3262,N_2594,N_2986);
nand U3263 (N_3263,N_2651,N_2630);
nand U3264 (N_3264,N_2892,N_2605);
and U3265 (N_3265,N_2854,N_2843);
xnor U3266 (N_3266,N_2778,N_2796);
and U3267 (N_3267,N_2572,N_2738);
nand U3268 (N_3268,N_2912,N_2852);
nor U3269 (N_3269,N_2590,N_2936);
and U3270 (N_3270,N_2847,N_2778);
nor U3271 (N_3271,N_2505,N_2852);
and U3272 (N_3272,N_2971,N_2711);
xnor U3273 (N_3273,N_2542,N_2523);
nand U3274 (N_3274,N_2726,N_2864);
or U3275 (N_3275,N_2849,N_2517);
nor U3276 (N_3276,N_2876,N_2788);
nor U3277 (N_3277,N_2970,N_2897);
or U3278 (N_3278,N_2780,N_2536);
nor U3279 (N_3279,N_2633,N_2812);
nor U3280 (N_3280,N_2686,N_2951);
nand U3281 (N_3281,N_2810,N_2594);
or U3282 (N_3282,N_2665,N_2749);
or U3283 (N_3283,N_2855,N_2860);
nor U3284 (N_3284,N_2831,N_2721);
or U3285 (N_3285,N_2777,N_2977);
and U3286 (N_3286,N_2627,N_2512);
or U3287 (N_3287,N_2918,N_2785);
and U3288 (N_3288,N_2856,N_2561);
nand U3289 (N_3289,N_2759,N_2993);
and U3290 (N_3290,N_2879,N_2623);
xnor U3291 (N_3291,N_2883,N_2991);
nor U3292 (N_3292,N_2548,N_2611);
and U3293 (N_3293,N_2845,N_2718);
xnor U3294 (N_3294,N_2706,N_2674);
nand U3295 (N_3295,N_2641,N_2662);
and U3296 (N_3296,N_2921,N_2894);
nand U3297 (N_3297,N_2729,N_2676);
xor U3298 (N_3298,N_2811,N_2596);
or U3299 (N_3299,N_2953,N_2668);
nor U3300 (N_3300,N_2572,N_2728);
or U3301 (N_3301,N_2884,N_2523);
nor U3302 (N_3302,N_2784,N_2851);
nand U3303 (N_3303,N_2743,N_2553);
and U3304 (N_3304,N_2861,N_2657);
xnor U3305 (N_3305,N_2603,N_2696);
and U3306 (N_3306,N_2946,N_2692);
nor U3307 (N_3307,N_2993,N_2691);
and U3308 (N_3308,N_2846,N_2998);
and U3309 (N_3309,N_2809,N_2938);
and U3310 (N_3310,N_2554,N_2753);
nand U3311 (N_3311,N_2640,N_2622);
xor U3312 (N_3312,N_2670,N_2748);
nand U3313 (N_3313,N_2798,N_2703);
nand U3314 (N_3314,N_2990,N_2985);
or U3315 (N_3315,N_2894,N_2926);
and U3316 (N_3316,N_2666,N_2815);
nor U3317 (N_3317,N_2674,N_2552);
or U3318 (N_3318,N_2676,N_2835);
or U3319 (N_3319,N_2594,N_2510);
and U3320 (N_3320,N_2849,N_2699);
and U3321 (N_3321,N_2614,N_2714);
nand U3322 (N_3322,N_2945,N_2629);
nor U3323 (N_3323,N_2754,N_2750);
and U3324 (N_3324,N_2798,N_2705);
nor U3325 (N_3325,N_2914,N_2878);
and U3326 (N_3326,N_2720,N_2914);
or U3327 (N_3327,N_2916,N_2639);
and U3328 (N_3328,N_2885,N_2590);
and U3329 (N_3329,N_2502,N_2632);
and U3330 (N_3330,N_2526,N_2776);
xnor U3331 (N_3331,N_2967,N_2758);
or U3332 (N_3332,N_2632,N_2836);
xor U3333 (N_3333,N_2670,N_2769);
xnor U3334 (N_3334,N_2573,N_2591);
nand U3335 (N_3335,N_2927,N_2597);
and U3336 (N_3336,N_2838,N_2827);
or U3337 (N_3337,N_2728,N_2966);
nand U3338 (N_3338,N_2813,N_2708);
and U3339 (N_3339,N_2875,N_2540);
nand U3340 (N_3340,N_2533,N_2733);
nand U3341 (N_3341,N_2745,N_2710);
or U3342 (N_3342,N_2831,N_2963);
and U3343 (N_3343,N_2852,N_2751);
nand U3344 (N_3344,N_2869,N_2812);
or U3345 (N_3345,N_2617,N_2696);
or U3346 (N_3346,N_2562,N_2884);
or U3347 (N_3347,N_2940,N_2579);
or U3348 (N_3348,N_2947,N_2567);
or U3349 (N_3349,N_2874,N_2560);
nor U3350 (N_3350,N_2969,N_2886);
nor U3351 (N_3351,N_2865,N_2526);
xnor U3352 (N_3352,N_2696,N_2802);
and U3353 (N_3353,N_2875,N_2974);
or U3354 (N_3354,N_2910,N_2761);
and U3355 (N_3355,N_2600,N_2934);
or U3356 (N_3356,N_2756,N_2504);
or U3357 (N_3357,N_2909,N_2812);
nand U3358 (N_3358,N_2812,N_2985);
or U3359 (N_3359,N_2738,N_2714);
nor U3360 (N_3360,N_2632,N_2916);
nor U3361 (N_3361,N_2626,N_2925);
xor U3362 (N_3362,N_2730,N_2582);
nand U3363 (N_3363,N_2942,N_2787);
xnor U3364 (N_3364,N_2762,N_2539);
or U3365 (N_3365,N_2642,N_2816);
and U3366 (N_3366,N_2763,N_2765);
or U3367 (N_3367,N_2714,N_2791);
and U3368 (N_3368,N_2803,N_2812);
or U3369 (N_3369,N_2546,N_2693);
or U3370 (N_3370,N_2639,N_2761);
and U3371 (N_3371,N_2840,N_2650);
nand U3372 (N_3372,N_2764,N_2591);
or U3373 (N_3373,N_2795,N_2967);
nor U3374 (N_3374,N_2589,N_2553);
nand U3375 (N_3375,N_2508,N_2800);
nand U3376 (N_3376,N_2625,N_2759);
nand U3377 (N_3377,N_2804,N_2665);
nor U3378 (N_3378,N_2977,N_2643);
and U3379 (N_3379,N_2972,N_2854);
nor U3380 (N_3380,N_2793,N_2779);
nand U3381 (N_3381,N_2786,N_2738);
or U3382 (N_3382,N_2616,N_2859);
nor U3383 (N_3383,N_2663,N_2632);
or U3384 (N_3384,N_2635,N_2745);
or U3385 (N_3385,N_2668,N_2692);
xnor U3386 (N_3386,N_2827,N_2950);
nor U3387 (N_3387,N_2741,N_2946);
nor U3388 (N_3388,N_2699,N_2677);
and U3389 (N_3389,N_2573,N_2902);
nor U3390 (N_3390,N_2555,N_2926);
or U3391 (N_3391,N_2675,N_2561);
or U3392 (N_3392,N_2870,N_2963);
nor U3393 (N_3393,N_2669,N_2904);
nor U3394 (N_3394,N_2807,N_2786);
or U3395 (N_3395,N_2742,N_2508);
nor U3396 (N_3396,N_2744,N_2810);
or U3397 (N_3397,N_2976,N_2809);
or U3398 (N_3398,N_2968,N_2783);
nand U3399 (N_3399,N_2891,N_2875);
nor U3400 (N_3400,N_2871,N_2714);
or U3401 (N_3401,N_2830,N_2510);
or U3402 (N_3402,N_2691,N_2685);
nand U3403 (N_3403,N_2754,N_2986);
and U3404 (N_3404,N_2910,N_2566);
or U3405 (N_3405,N_2736,N_2703);
nor U3406 (N_3406,N_2531,N_2884);
or U3407 (N_3407,N_2831,N_2979);
nand U3408 (N_3408,N_2968,N_2875);
or U3409 (N_3409,N_2865,N_2510);
or U3410 (N_3410,N_2943,N_2738);
or U3411 (N_3411,N_2828,N_2878);
and U3412 (N_3412,N_2546,N_2900);
and U3413 (N_3413,N_2596,N_2769);
nor U3414 (N_3414,N_2969,N_2891);
nor U3415 (N_3415,N_2575,N_2726);
and U3416 (N_3416,N_2576,N_2699);
nor U3417 (N_3417,N_2958,N_2554);
and U3418 (N_3418,N_2892,N_2913);
and U3419 (N_3419,N_2853,N_2838);
and U3420 (N_3420,N_2781,N_2835);
or U3421 (N_3421,N_2766,N_2950);
nand U3422 (N_3422,N_2672,N_2916);
xnor U3423 (N_3423,N_2713,N_2658);
and U3424 (N_3424,N_2647,N_2659);
xor U3425 (N_3425,N_2779,N_2635);
nand U3426 (N_3426,N_2927,N_2537);
and U3427 (N_3427,N_2856,N_2533);
nor U3428 (N_3428,N_2823,N_2514);
nand U3429 (N_3429,N_2993,N_2549);
nor U3430 (N_3430,N_2575,N_2557);
nor U3431 (N_3431,N_2700,N_2914);
or U3432 (N_3432,N_2979,N_2512);
nand U3433 (N_3433,N_2715,N_2901);
nand U3434 (N_3434,N_2659,N_2641);
and U3435 (N_3435,N_2709,N_2774);
nand U3436 (N_3436,N_2961,N_2519);
nor U3437 (N_3437,N_2654,N_2550);
nand U3438 (N_3438,N_2858,N_2855);
and U3439 (N_3439,N_2971,N_2832);
nand U3440 (N_3440,N_2860,N_2753);
and U3441 (N_3441,N_2717,N_2635);
nor U3442 (N_3442,N_2829,N_2555);
nor U3443 (N_3443,N_2768,N_2717);
and U3444 (N_3444,N_2809,N_2721);
xor U3445 (N_3445,N_2870,N_2668);
or U3446 (N_3446,N_2653,N_2735);
nor U3447 (N_3447,N_2705,N_2942);
nand U3448 (N_3448,N_2805,N_2627);
and U3449 (N_3449,N_2761,N_2646);
xor U3450 (N_3450,N_2537,N_2721);
nor U3451 (N_3451,N_2872,N_2835);
nor U3452 (N_3452,N_2604,N_2599);
and U3453 (N_3453,N_2517,N_2661);
nor U3454 (N_3454,N_2504,N_2909);
nor U3455 (N_3455,N_2805,N_2558);
nor U3456 (N_3456,N_2563,N_2650);
nand U3457 (N_3457,N_2783,N_2539);
and U3458 (N_3458,N_2543,N_2951);
nand U3459 (N_3459,N_2725,N_2525);
nor U3460 (N_3460,N_2524,N_2522);
or U3461 (N_3461,N_2819,N_2802);
and U3462 (N_3462,N_2963,N_2800);
nor U3463 (N_3463,N_2858,N_2540);
and U3464 (N_3464,N_2939,N_2844);
or U3465 (N_3465,N_2785,N_2798);
or U3466 (N_3466,N_2784,N_2811);
nand U3467 (N_3467,N_2524,N_2846);
or U3468 (N_3468,N_2845,N_2594);
or U3469 (N_3469,N_2956,N_2607);
or U3470 (N_3470,N_2820,N_2606);
nand U3471 (N_3471,N_2864,N_2641);
or U3472 (N_3472,N_2789,N_2787);
nor U3473 (N_3473,N_2779,N_2557);
nor U3474 (N_3474,N_2713,N_2870);
nor U3475 (N_3475,N_2699,N_2611);
xor U3476 (N_3476,N_2886,N_2864);
nand U3477 (N_3477,N_2672,N_2626);
and U3478 (N_3478,N_2833,N_2952);
or U3479 (N_3479,N_2629,N_2588);
xor U3480 (N_3480,N_2836,N_2817);
xor U3481 (N_3481,N_2866,N_2935);
and U3482 (N_3482,N_2861,N_2811);
and U3483 (N_3483,N_2945,N_2873);
and U3484 (N_3484,N_2820,N_2908);
nand U3485 (N_3485,N_2682,N_2725);
or U3486 (N_3486,N_2961,N_2661);
and U3487 (N_3487,N_2711,N_2892);
nand U3488 (N_3488,N_2959,N_2656);
or U3489 (N_3489,N_2535,N_2881);
or U3490 (N_3490,N_2564,N_2771);
and U3491 (N_3491,N_2511,N_2507);
or U3492 (N_3492,N_2677,N_2560);
nor U3493 (N_3493,N_2641,N_2809);
or U3494 (N_3494,N_2855,N_2800);
nor U3495 (N_3495,N_2840,N_2699);
nor U3496 (N_3496,N_2683,N_2925);
nor U3497 (N_3497,N_2900,N_2713);
and U3498 (N_3498,N_2932,N_2601);
xor U3499 (N_3499,N_2991,N_2534);
and U3500 (N_3500,N_3223,N_3481);
nand U3501 (N_3501,N_3188,N_3114);
nor U3502 (N_3502,N_3135,N_3306);
or U3503 (N_3503,N_3294,N_3151);
nand U3504 (N_3504,N_3133,N_3457);
nor U3505 (N_3505,N_3022,N_3439);
or U3506 (N_3506,N_3371,N_3462);
or U3507 (N_3507,N_3435,N_3218);
nand U3508 (N_3508,N_3139,N_3428);
or U3509 (N_3509,N_3450,N_3455);
xor U3510 (N_3510,N_3061,N_3083);
and U3511 (N_3511,N_3473,N_3434);
nand U3512 (N_3512,N_3251,N_3249);
or U3513 (N_3513,N_3447,N_3275);
xnor U3514 (N_3514,N_3357,N_3209);
nor U3515 (N_3515,N_3366,N_3208);
nand U3516 (N_3516,N_3383,N_3395);
and U3517 (N_3517,N_3464,N_3363);
or U3518 (N_3518,N_3090,N_3191);
or U3519 (N_3519,N_3169,N_3325);
nand U3520 (N_3520,N_3041,N_3417);
and U3521 (N_3521,N_3107,N_3027);
and U3522 (N_3522,N_3475,N_3305);
nand U3523 (N_3523,N_3403,N_3192);
nand U3524 (N_3524,N_3477,N_3486);
or U3525 (N_3525,N_3045,N_3051);
and U3526 (N_3526,N_3350,N_3073);
or U3527 (N_3527,N_3173,N_3063);
nor U3528 (N_3528,N_3004,N_3418);
and U3529 (N_3529,N_3245,N_3315);
and U3530 (N_3530,N_3202,N_3131);
xnor U3531 (N_3531,N_3399,N_3287);
or U3532 (N_3532,N_3240,N_3229);
xor U3533 (N_3533,N_3016,N_3256);
nand U3534 (N_3534,N_3343,N_3308);
nor U3535 (N_3535,N_3364,N_3310);
nor U3536 (N_3536,N_3204,N_3289);
or U3537 (N_3537,N_3127,N_3242);
or U3538 (N_3538,N_3085,N_3230);
or U3539 (N_3539,N_3424,N_3433);
and U3540 (N_3540,N_3125,N_3214);
nand U3541 (N_3541,N_3471,N_3194);
nor U3542 (N_3542,N_3316,N_3049);
or U3543 (N_3543,N_3117,N_3300);
nand U3544 (N_3544,N_3332,N_3410);
and U3545 (N_3545,N_3312,N_3373);
nor U3546 (N_3546,N_3291,N_3241);
nor U3547 (N_3547,N_3277,N_3437);
nor U3548 (N_3548,N_3033,N_3148);
or U3549 (N_3549,N_3220,N_3165);
or U3550 (N_3550,N_3124,N_3335);
and U3551 (N_3551,N_3452,N_3468);
xor U3552 (N_3552,N_3014,N_3311);
or U3553 (N_3553,N_3039,N_3062);
nor U3554 (N_3554,N_3258,N_3448);
nand U3555 (N_3555,N_3374,N_3094);
nor U3556 (N_3556,N_3175,N_3196);
and U3557 (N_3557,N_3381,N_3222);
nand U3558 (N_3558,N_3327,N_3384);
nand U3559 (N_3559,N_3239,N_3146);
nand U3560 (N_3560,N_3338,N_3358);
nand U3561 (N_3561,N_3326,N_3487);
or U3562 (N_3562,N_3040,N_3162);
and U3563 (N_3563,N_3279,N_3183);
nor U3564 (N_3564,N_3420,N_3172);
nor U3565 (N_3565,N_3147,N_3382);
or U3566 (N_3566,N_3212,N_3260);
nor U3567 (N_3567,N_3262,N_3496);
and U3568 (N_3568,N_3012,N_3421);
nand U3569 (N_3569,N_3054,N_3353);
nor U3570 (N_3570,N_3484,N_3330);
xor U3571 (N_3571,N_3203,N_3155);
xor U3572 (N_3572,N_3415,N_3419);
nand U3573 (N_3573,N_3375,N_3231);
nor U3574 (N_3574,N_3334,N_3390);
or U3575 (N_3575,N_3170,N_3317);
nand U3576 (N_3576,N_3344,N_3370);
and U3577 (N_3577,N_3337,N_3152);
or U3578 (N_3578,N_3154,N_3436);
or U3579 (N_3579,N_3044,N_3086);
xor U3580 (N_3580,N_3138,N_3093);
nand U3581 (N_3581,N_3368,N_3206);
and U3582 (N_3582,N_3032,N_3128);
xor U3583 (N_3583,N_3098,N_3122);
xor U3584 (N_3584,N_3372,N_3431);
nand U3585 (N_3585,N_3442,N_3469);
or U3586 (N_3586,N_3187,N_3323);
or U3587 (N_3587,N_3143,N_3215);
nor U3588 (N_3588,N_3309,N_3362);
and U3589 (N_3589,N_3365,N_3461);
nand U3590 (N_3590,N_3048,N_3485);
or U3591 (N_3591,N_3081,N_3059);
nand U3592 (N_3592,N_3095,N_3414);
and U3593 (N_3593,N_3159,N_3346);
or U3594 (N_3594,N_3112,N_3401);
nor U3595 (N_3595,N_3376,N_3444);
nor U3596 (N_3596,N_3084,N_3109);
nand U3597 (N_3597,N_3184,N_3149);
nor U3598 (N_3598,N_3068,N_3168);
xnor U3599 (N_3599,N_3460,N_3440);
or U3600 (N_3600,N_3288,N_3299);
or U3601 (N_3601,N_3087,N_3181);
and U3602 (N_3602,N_3341,N_3029);
and U3603 (N_3603,N_3195,N_3019);
xor U3604 (N_3604,N_3120,N_3478);
or U3605 (N_3605,N_3186,N_3285);
nor U3606 (N_3606,N_3367,N_3225);
nor U3607 (N_3607,N_3438,N_3250);
nor U3608 (N_3608,N_3035,N_3066);
nor U3609 (N_3609,N_3456,N_3198);
xnor U3610 (N_3610,N_3210,N_3342);
nor U3611 (N_3611,N_3157,N_3071);
or U3612 (N_3612,N_3103,N_3318);
and U3613 (N_3613,N_3331,N_3489);
or U3614 (N_3614,N_3216,N_3314);
nor U3615 (N_3615,N_3409,N_3321);
nor U3616 (N_3616,N_3479,N_3179);
nor U3617 (N_3617,N_3483,N_3282);
nor U3618 (N_3618,N_3011,N_3339);
nor U3619 (N_3619,N_3036,N_3388);
or U3620 (N_3620,N_3057,N_3190);
nand U3621 (N_3621,N_3176,N_3246);
xnor U3622 (N_3622,N_3089,N_3056);
or U3623 (N_3623,N_3096,N_3322);
nor U3624 (N_3624,N_3392,N_3271);
xor U3625 (N_3625,N_3150,N_3009);
and U3626 (N_3626,N_3118,N_3058);
nor U3627 (N_3627,N_3145,N_3272);
nand U3628 (N_3628,N_3088,N_3425);
nor U3629 (N_3629,N_3293,N_3072);
or U3630 (N_3630,N_3377,N_3007);
nand U3631 (N_3631,N_3261,N_3319);
nand U3632 (N_3632,N_3449,N_3351);
or U3633 (N_3633,N_3497,N_3008);
and U3634 (N_3634,N_3278,N_3298);
xor U3635 (N_3635,N_3174,N_3281);
nand U3636 (N_3636,N_3394,N_3263);
nand U3637 (N_3637,N_3284,N_3295);
and U3638 (N_3638,N_3432,N_3013);
and U3639 (N_3639,N_3047,N_3043);
xor U3640 (N_3640,N_3270,N_3416);
nand U3641 (N_3641,N_3182,N_3385);
and U3642 (N_3642,N_3389,N_3329);
nand U3643 (N_3643,N_3467,N_3158);
nand U3644 (N_3644,N_3034,N_3052);
nand U3645 (N_3645,N_3453,N_3177);
nor U3646 (N_3646,N_3255,N_3280);
and U3647 (N_3647,N_3313,N_3021);
or U3648 (N_3648,N_3104,N_3472);
nor U3649 (N_3649,N_3380,N_3193);
nand U3650 (N_3650,N_3200,N_3402);
nor U3651 (N_3651,N_3099,N_3064);
or U3652 (N_3652,N_3266,N_3247);
or U3653 (N_3653,N_3053,N_3378);
nand U3654 (N_3654,N_3030,N_3235);
xnor U3655 (N_3655,N_3077,N_3466);
nand U3656 (N_3656,N_3470,N_3274);
nor U3657 (N_3657,N_3110,N_3207);
nor U3658 (N_3658,N_3493,N_3498);
nor U3659 (N_3659,N_3387,N_3221);
nand U3660 (N_3660,N_3273,N_3050);
and U3661 (N_3661,N_3345,N_3166);
xnor U3662 (N_3662,N_3348,N_3324);
or U3663 (N_3663,N_3199,N_3038);
or U3664 (N_3664,N_3031,N_3082);
or U3665 (N_3665,N_3140,N_3115);
and U3666 (N_3666,N_3163,N_3328);
and U3667 (N_3667,N_3228,N_3265);
nor U3668 (N_3668,N_3101,N_3304);
and U3669 (N_3669,N_3001,N_3010);
nor U3670 (N_3670,N_3296,N_3205);
nor U3671 (N_3671,N_3026,N_3015);
and U3672 (N_3672,N_3025,N_3423);
or U3673 (N_3673,N_3491,N_3268);
or U3674 (N_3674,N_3142,N_3290);
nand U3675 (N_3675,N_3474,N_3233);
nand U3676 (N_3676,N_3189,N_3136);
or U3677 (N_3677,N_3046,N_3356);
nand U3678 (N_3678,N_3259,N_3232);
or U3679 (N_3679,N_3113,N_3495);
nand U3680 (N_3680,N_3404,N_3267);
xor U3681 (N_3681,N_3126,N_3426);
nand U3682 (N_3682,N_3217,N_3134);
nor U3683 (N_3683,N_3091,N_3352);
nand U3684 (N_3684,N_3121,N_3340);
nor U3685 (N_3685,N_3076,N_3005);
or U3686 (N_3686,N_3024,N_3119);
nor U3687 (N_3687,N_3445,N_3028);
or U3688 (N_3688,N_3349,N_3441);
or U3689 (N_3689,N_3406,N_3161);
nor U3690 (N_3690,N_3347,N_3069);
nor U3691 (N_3691,N_3248,N_3396);
nor U3692 (N_3692,N_3405,N_3123);
xor U3693 (N_3693,N_3292,N_3160);
or U3694 (N_3694,N_3037,N_3197);
nor U3695 (N_3695,N_3301,N_3302);
and U3696 (N_3696,N_3320,N_3137);
nand U3697 (N_3697,N_3018,N_3129);
and U3698 (N_3698,N_3499,N_3067);
nor U3699 (N_3699,N_3430,N_3237);
xnor U3700 (N_3700,N_3454,N_3476);
xor U3701 (N_3701,N_3333,N_3156);
nor U3702 (N_3702,N_3354,N_3264);
nand U3703 (N_3703,N_3482,N_3042);
or U3704 (N_3704,N_3480,N_3391);
and U3705 (N_3705,N_3269,N_3070);
nand U3706 (N_3706,N_3398,N_3201);
and U3707 (N_3707,N_3253,N_3065);
nand U3708 (N_3708,N_3429,N_3243);
and U3709 (N_3709,N_3244,N_3141);
nor U3710 (N_3710,N_3060,N_3361);
nor U3711 (N_3711,N_3413,N_3020);
nor U3712 (N_3712,N_3283,N_3458);
and U3713 (N_3713,N_3451,N_3297);
xor U3714 (N_3714,N_3336,N_3097);
nor U3715 (N_3715,N_3130,N_3074);
or U3716 (N_3716,N_3360,N_3185);
nand U3717 (N_3717,N_3397,N_3488);
nor U3718 (N_3718,N_3369,N_3355);
nand U3719 (N_3719,N_3227,N_3080);
nor U3720 (N_3720,N_3407,N_3055);
and U3721 (N_3721,N_3379,N_3422);
or U3722 (N_3722,N_3393,N_3144);
nand U3723 (N_3723,N_3075,N_3153);
nand U3724 (N_3724,N_3252,N_3002);
and U3725 (N_3725,N_3006,N_3234);
and U3726 (N_3726,N_3459,N_3000);
nor U3727 (N_3727,N_3400,N_3236);
nor U3728 (N_3728,N_3446,N_3359);
nand U3729 (N_3729,N_3219,N_3132);
and U3730 (N_3730,N_3111,N_3427);
xnor U3731 (N_3731,N_3463,N_3286);
nand U3732 (N_3732,N_3254,N_3492);
nand U3733 (N_3733,N_3303,N_3017);
nor U3734 (N_3734,N_3003,N_3092);
and U3735 (N_3735,N_3226,N_3167);
and U3736 (N_3736,N_3465,N_3023);
and U3737 (N_3737,N_3224,N_3116);
or U3738 (N_3738,N_3238,N_3102);
xnor U3739 (N_3739,N_3494,N_3180);
or U3740 (N_3740,N_3100,N_3412);
nand U3741 (N_3741,N_3307,N_3490);
nor U3742 (N_3742,N_3171,N_3257);
nand U3743 (N_3743,N_3211,N_3443);
and U3744 (N_3744,N_3105,N_3276);
or U3745 (N_3745,N_3164,N_3078);
nand U3746 (N_3746,N_3213,N_3079);
nor U3747 (N_3747,N_3108,N_3106);
and U3748 (N_3748,N_3411,N_3386);
or U3749 (N_3749,N_3178,N_3408);
xor U3750 (N_3750,N_3241,N_3418);
nor U3751 (N_3751,N_3249,N_3377);
nand U3752 (N_3752,N_3185,N_3213);
nor U3753 (N_3753,N_3118,N_3130);
nor U3754 (N_3754,N_3440,N_3149);
nor U3755 (N_3755,N_3440,N_3010);
or U3756 (N_3756,N_3157,N_3460);
or U3757 (N_3757,N_3324,N_3095);
xor U3758 (N_3758,N_3385,N_3436);
nor U3759 (N_3759,N_3022,N_3446);
nand U3760 (N_3760,N_3002,N_3437);
nand U3761 (N_3761,N_3295,N_3219);
nand U3762 (N_3762,N_3253,N_3362);
or U3763 (N_3763,N_3188,N_3028);
nand U3764 (N_3764,N_3230,N_3402);
xnor U3765 (N_3765,N_3012,N_3357);
nand U3766 (N_3766,N_3406,N_3341);
or U3767 (N_3767,N_3293,N_3408);
and U3768 (N_3768,N_3144,N_3497);
and U3769 (N_3769,N_3072,N_3174);
or U3770 (N_3770,N_3322,N_3109);
and U3771 (N_3771,N_3434,N_3132);
or U3772 (N_3772,N_3273,N_3332);
or U3773 (N_3773,N_3429,N_3116);
or U3774 (N_3774,N_3317,N_3448);
nor U3775 (N_3775,N_3088,N_3321);
or U3776 (N_3776,N_3287,N_3338);
or U3777 (N_3777,N_3458,N_3285);
nor U3778 (N_3778,N_3146,N_3057);
and U3779 (N_3779,N_3252,N_3125);
nand U3780 (N_3780,N_3134,N_3471);
and U3781 (N_3781,N_3267,N_3476);
and U3782 (N_3782,N_3210,N_3000);
nand U3783 (N_3783,N_3229,N_3046);
nor U3784 (N_3784,N_3070,N_3191);
nor U3785 (N_3785,N_3440,N_3445);
or U3786 (N_3786,N_3108,N_3495);
or U3787 (N_3787,N_3345,N_3175);
nand U3788 (N_3788,N_3191,N_3302);
or U3789 (N_3789,N_3174,N_3399);
nand U3790 (N_3790,N_3465,N_3256);
nand U3791 (N_3791,N_3298,N_3287);
and U3792 (N_3792,N_3061,N_3213);
and U3793 (N_3793,N_3185,N_3423);
and U3794 (N_3794,N_3199,N_3051);
nand U3795 (N_3795,N_3108,N_3068);
or U3796 (N_3796,N_3082,N_3316);
nand U3797 (N_3797,N_3496,N_3253);
nor U3798 (N_3798,N_3053,N_3135);
nor U3799 (N_3799,N_3018,N_3252);
nand U3800 (N_3800,N_3178,N_3052);
nor U3801 (N_3801,N_3234,N_3235);
nand U3802 (N_3802,N_3020,N_3343);
nor U3803 (N_3803,N_3335,N_3091);
and U3804 (N_3804,N_3441,N_3080);
nand U3805 (N_3805,N_3232,N_3099);
or U3806 (N_3806,N_3370,N_3012);
nor U3807 (N_3807,N_3271,N_3168);
nand U3808 (N_3808,N_3415,N_3405);
or U3809 (N_3809,N_3139,N_3145);
or U3810 (N_3810,N_3075,N_3178);
and U3811 (N_3811,N_3043,N_3474);
xor U3812 (N_3812,N_3405,N_3446);
nor U3813 (N_3813,N_3411,N_3309);
nor U3814 (N_3814,N_3128,N_3286);
nand U3815 (N_3815,N_3283,N_3046);
nor U3816 (N_3816,N_3056,N_3182);
or U3817 (N_3817,N_3243,N_3294);
or U3818 (N_3818,N_3197,N_3214);
nand U3819 (N_3819,N_3036,N_3283);
and U3820 (N_3820,N_3099,N_3479);
nor U3821 (N_3821,N_3406,N_3347);
or U3822 (N_3822,N_3465,N_3461);
and U3823 (N_3823,N_3119,N_3314);
nor U3824 (N_3824,N_3115,N_3060);
nor U3825 (N_3825,N_3431,N_3376);
nor U3826 (N_3826,N_3485,N_3068);
nor U3827 (N_3827,N_3102,N_3051);
nor U3828 (N_3828,N_3108,N_3485);
or U3829 (N_3829,N_3467,N_3161);
and U3830 (N_3830,N_3431,N_3476);
or U3831 (N_3831,N_3020,N_3004);
nand U3832 (N_3832,N_3119,N_3011);
or U3833 (N_3833,N_3027,N_3012);
and U3834 (N_3834,N_3179,N_3260);
nor U3835 (N_3835,N_3450,N_3018);
and U3836 (N_3836,N_3191,N_3271);
xor U3837 (N_3837,N_3231,N_3139);
and U3838 (N_3838,N_3046,N_3350);
or U3839 (N_3839,N_3041,N_3093);
and U3840 (N_3840,N_3184,N_3159);
and U3841 (N_3841,N_3308,N_3360);
and U3842 (N_3842,N_3077,N_3259);
nor U3843 (N_3843,N_3433,N_3271);
or U3844 (N_3844,N_3001,N_3335);
nand U3845 (N_3845,N_3016,N_3389);
or U3846 (N_3846,N_3315,N_3146);
nor U3847 (N_3847,N_3175,N_3279);
and U3848 (N_3848,N_3293,N_3228);
nand U3849 (N_3849,N_3221,N_3423);
or U3850 (N_3850,N_3281,N_3032);
nand U3851 (N_3851,N_3328,N_3314);
nand U3852 (N_3852,N_3405,N_3112);
nor U3853 (N_3853,N_3037,N_3484);
nor U3854 (N_3854,N_3222,N_3114);
nand U3855 (N_3855,N_3150,N_3065);
or U3856 (N_3856,N_3372,N_3222);
and U3857 (N_3857,N_3039,N_3483);
nand U3858 (N_3858,N_3311,N_3463);
nor U3859 (N_3859,N_3055,N_3188);
nor U3860 (N_3860,N_3046,N_3355);
nor U3861 (N_3861,N_3210,N_3464);
and U3862 (N_3862,N_3264,N_3101);
or U3863 (N_3863,N_3416,N_3282);
nand U3864 (N_3864,N_3121,N_3225);
or U3865 (N_3865,N_3268,N_3015);
nand U3866 (N_3866,N_3456,N_3122);
nand U3867 (N_3867,N_3185,N_3236);
nor U3868 (N_3868,N_3237,N_3250);
or U3869 (N_3869,N_3455,N_3492);
nand U3870 (N_3870,N_3023,N_3098);
nor U3871 (N_3871,N_3458,N_3434);
and U3872 (N_3872,N_3041,N_3472);
and U3873 (N_3873,N_3333,N_3063);
and U3874 (N_3874,N_3372,N_3184);
or U3875 (N_3875,N_3153,N_3089);
nor U3876 (N_3876,N_3238,N_3088);
nor U3877 (N_3877,N_3130,N_3127);
nor U3878 (N_3878,N_3256,N_3144);
nand U3879 (N_3879,N_3105,N_3462);
or U3880 (N_3880,N_3364,N_3360);
and U3881 (N_3881,N_3136,N_3054);
nor U3882 (N_3882,N_3200,N_3125);
or U3883 (N_3883,N_3427,N_3106);
xnor U3884 (N_3884,N_3425,N_3008);
or U3885 (N_3885,N_3067,N_3401);
nor U3886 (N_3886,N_3323,N_3309);
or U3887 (N_3887,N_3018,N_3167);
and U3888 (N_3888,N_3178,N_3110);
and U3889 (N_3889,N_3403,N_3032);
nand U3890 (N_3890,N_3040,N_3240);
and U3891 (N_3891,N_3210,N_3388);
xnor U3892 (N_3892,N_3129,N_3116);
nand U3893 (N_3893,N_3092,N_3006);
or U3894 (N_3894,N_3085,N_3364);
and U3895 (N_3895,N_3049,N_3051);
nand U3896 (N_3896,N_3326,N_3372);
and U3897 (N_3897,N_3321,N_3286);
xnor U3898 (N_3898,N_3387,N_3054);
and U3899 (N_3899,N_3115,N_3498);
and U3900 (N_3900,N_3147,N_3200);
nand U3901 (N_3901,N_3386,N_3261);
and U3902 (N_3902,N_3276,N_3112);
nand U3903 (N_3903,N_3330,N_3342);
or U3904 (N_3904,N_3409,N_3167);
nand U3905 (N_3905,N_3057,N_3105);
nand U3906 (N_3906,N_3346,N_3037);
and U3907 (N_3907,N_3176,N_3479);
nand U3908 (N_3908,N_3352,N_3201);
or U3909 (N_3909,N_3454,N_3338);
nand U3910 (N_3910,N_3465,N_3018);
xnor U3911 (N_3911,N_3228,N_3184);
nor U3912 (N_3912,N_3310,N_3478);
nor U3913 (N_3913,N_3129,N_3034);
nor U3914 (N_3914,N_3457,N_3041);
and U3915 (N_3915,N_3298,N_3036);
nand U3916 (N_3916,N_3228,N_3180);
nor U3917 (N_3917,N_3312,N_3073);
or U3918 (N_3918,N_3467,N_3274);
or U3919 (N_3919,N_3405,N_3122);
and U3920 (N_3920,N_3086,N_3373);
and U3921 (N_3921,N_3341,N_3049);
or U3922 (N_3922,N_3443,N_3474);
or U3923 (N_3923,N_3010,N_3452);
or U3924 (N_3924,N_3347,N_3430);
and U3925 (N_3925,N_3039,N_3337);
nand U3926 (N_3926,N_3468,N_3007);
or U3927 (N_3927,N_3471,N_3083);
and U3928 (N_3928,N_3396,N_3334);
and U3929 (N_3929,N_3189,N_3114);
nor U3930 (N_3930,N_3041,N_3480);
and U3931 (N_3931,N_3227,N_3367);
and U3932 (N_3932,N_3328,N_3445);
xnor U3933 (N_3933,N_3314,N_3075);
and U3934 (N_3934,N_3025,N_3184);
nor U3935 (N_3935,N_3247,N_3391);
and U3936 (N_3936,N_3301,N_3403);
nand U3937 (N_3937,N_3052,N_3176);
or U3938 (N_3938,N_3296,N_3213);
and U3939 (N_3939,N_3082,N_3070);
nor U3940 (N_3940,N_3404,N_3219);
nor U3941 (N_3941,N_3180,N_3036);
or U3942 (N_3942,N_3281,N_3442);
nand U3943 (N_3943,N_3055,N_3356);
nor U3944 (N_3944,N_3352,N_3096);
nor U3945 (N_3945,N_3421,N_3094);
nor U3946 (N_3946,N_3196,N_3005);
or U3947 (N_3947,N_3193,N_3084);
nand U3948 (N_3948,N_3349,N_3192);
and U3949 (N_3949,N_3032,N_3235);
or U3950 (N_3950,N_3076,N_3371);
nand U3951 (N_3951,N_3164,N_3366);
nand U3952 (N_3952,N_3021,N_3360);
and U3953 (N_3953,N_3387,N_3488);
or U3954 (N_3954,N_3076,N_3288);
and U3955 (N_3955,N_3344,N_3153);
and U3956 (N_3956,N_3248,N_3496);
or U3957 (N_3957,N_3017,N_3124);
or U3958 (N_3958,N_3361,N_3413);
xnor U3959 (N_3959,N_3391,N_3436);
or U3960 (N_3960,N_3145,N_3210);
nor U3961 (N_3961,N_3363,N_3276);
nor U3962 (N_3962,N_3051,N_3088);
nor U3963 (N_3963,N_3243,N_3453);
or U3964 (N_3964,N_3417,N_3486);
nand U3965 (N_3965,N_3045,N_3093);
nor U3966 (N_3966,N_3425,N_3055);
or U3967 (N_3967,N_3494,N_3002);
nand U3968 (N_3968,N_3323,N_3197);
nor U3969 (N_3969,N_3355,N_3152);
and U3970 (N_3970,N_3057,N_3212);
nand U3971 (N_3971,N_3439,N_3118);
and U3972 (N_3972,N_3158,N_3078);
nor U3973 (N_3973,N_3045,N_3317);
or U3974 (N_3974,N_3207,N_3164);
nor U3975 (N_3975,N_3483,N_3304);
or U3976 (N_3976,N_3392,N_3425);
and U3977 (N_3977,N_3480,N_3118);
or U3978 (N_3978,N_3296,N_3166);
and U3979 (N_3979,N_3426,N_3226);
nand U3980 (N_3980,N_3393,N_3244);
and U3981 (N_3981,N_3152,N_3295);
and U3982 (N_3982,N_3125,N_3051);
or U3983 (N_3983,N_3161,N_3219);
nor U3984 (N_3984,N_3013,N_3296);
xnor U3985 (N_3985,N_3354,N_3477);
nor U3986 (N_3986,N_3345,N_3348);
and U3987 (N_3987,N_3023,N_3377);
xnor U3988 (N_3988,N_3190,N_3406);
xnor U3989 (N_3989,N_3114,N_3268);
and U3990 (N_3990,N_3492,N_3225);
or U3991 (N_3991,N_3322,N_3490);
nor U3992 (N_3992,N_3163,N_3157);
nor U3993 (N_3993,N_3207,N_3307);
xnor U3994 (N_3994,N_3122,N_3050);
and U3995 (N_3995,N_3487,N_3029);
nand U3996 (N_3996,N_3135,N_3062);
nor U3997 (N_3997,N_3347,N_3084);
and U3998 (N_3998,N_3221,N_3404);
nand U3999 (N_3999,N_3292,N_3331);
nand U4000 (N_4000,N_3561,N_3716);
nand U4001 (N_4001,N_3682,N_3557);
or U4002 (N_4002,N_3672,N_3519);
nand U4003 (N_4003,N_3888,N_3920);
or U4004 (N_4004,N_3507,N_3902);
nor U4005 (N_4005,N_3663,N_3714);
or U4006 (N_4006,N_3758,N_3547);
nand U4007 (N_4007,N_3743,N_3580);
nand U4008 (N_4008,N_3844,N_3983);
and U4009 (N_4009,N_3807,N_3855);
nor U4010 (N_4010,N_3554,N_3717);
xnor U4011 (N_4011,N_3850,N_3726);
or U4012 (N_4012,N_3738,N_3598);
nand U4013 (N_4013,N_3503,N_3962);
and U4014 (N_4014,N_3674,N_3898);
nand U4015 (N_4015,N_3552,N_3804);
or U4016 (N_4016,N_3708,N_3529);
and U4017 (N_4017,N_3742,N_3915);
xor U4018 (N_4018,N_3560,N_3876);
or U4019 (N_4019,N_3836,N_3764);
xnor U4020 (N_4020,N_3950,N_3949);
nand U4021 (N_4021,N_3628,N_3927);
xnor U4022 (N_4022,N_3740,N_3750);
nand U4023 (N_4023,N_3860,N_3651);
or U4024 (N_4024,N_3562,N_3734);
xor U4025 (N_4025,N_3930,N_3774);
nand U4026 (N_4026,N_3765,N_3683);
or U4027 (N_4027,N_3614,N_3918);
nand U4028 (N_4028,N_3586,N_3730);
xor U4029 (N_4029,N_3642,N_3718);
nor U4030 (N_4030,N_3572,N_3892);
and U4031 (N_4031,N_3869,N_3942);
nand U4032 (N_4032,N_3737,N_3986);
nor U4033 (N_4033,N_3558,N_3867);
nand U4034 (N_4034,N_3537,N_3591);
nor U4035 (N_4035,N_3822,N_3788);
nand U4036 (N_4036,N_3505,N_3813);
nor U4037 (N_4037,N_3875,N_3512);
and U4038 (N_4038,N_3864,N_3951);
and U4039 (N_4039,N_3555,N_3859);
xnor U4040 (N_4040,N_3973,N_3854);
nor U4041 (N_4041,N_3751,N_3964);
or U4042 (N_4042,N_3511,N_3709);
nor U4043 (N_4043,N_3666,N_3881);
or U4044 (N_4044,N_3904,N_3522);
nor U4045 (N_4045,N_3833,N_3939);
and U4046 (N_4046,N_3946,N_3545);
and U4047 (N_4047,N_3821,N_3638);
nor U4048 (N_4048,N_3749,N_3935);
nand U4049 (N_4049,N_3612,N_3992);
and U4050 (N_4050,N_3744,N_3584);
nor U4051 (N_4051,N_3798,N_3914);
or U4052 (N_4052,N_3923,N_3766);
nand U4053 (N_4053,N_3961,N_3903);
and U4054 (N_4054,N_3908,N_3994);
or U4055 (N_4055,N_3632,N_3910);
or U4056 (N_4056,N_3606,N_3999);
nand U4057 (N_4057,N_3840,N_3582);
and U4058 (N_4058,N_3891,N_3513);
nor U4059 (N_4059,N_3814,N_3803);
or U4060 (N_4060,N_3775,N_3787);
nor U4061 (N_4061,N_3616,N_3877);
nor U4062 (N_4062,N_3795,N_3544);
or U4063 (N_4063,N_3963,N_3812);
nor U4064 (N_4064,N_3553,N_3634);
or U4065 (N_4065,N_3509,N_3593);
nand U4066 (N_4066,N_3954,N_3669);
xnor U4067 (N_4067,N_3622,N_3633);
xor U4068 (N_4068,N_3667,N_3694);
and U4069 (N_4069,N_3835,N_3549);
xor U4070 (N_4070,N_3928,N_3834);
nand U4071 (N_4071,N_3601,N_3525);
and U4072 (N_4072,N_3665,N_3783);
and U4073 (N_4073,N_3801,N_3579);
nand U4074 (N_4074,N_3689,N_3662);
and U4075 (N_4075,N_3504,N_3782);
nand U4076 (N_4076,N_3701,N_3873);
or U4077 (N_4077,N_3648,N_3976);
nand U4078 (N_4078,N_3851,N_3500);
or U4079 (N_4079,N_3531,N_3621);
nor U4080 (N_4080,N_3733,N_3583);
xor U4081 (N_4081,N_3828,N_3546);
and U4082 (N_4082,N_3917,N_3780);
nor U4083 (N_4083,N_3594,N_3720);
or U4084 (N_4084,N_3874,N_3664);
nand U4085 (N_4085,N_3684,N_3965);
xnor U4086 (N_4086,N_3559,N_3631);
and U4087 (N_4087,N_3995,N_3657);
nand U4088 (N_4088,N_3956,N_3985);
or U4089 (N_4089,N_3732,N_3517);
or U4090 (N_4090,N_3686,N_3792);
nor U4091 (N_4091,N_3880,N_3602);
and U4092 (N_4092,N_3970,N_3652);
nand U4093 (N_4093,N_3568,N_3567);
nand U4094 (N_4094,N_3696,N_3654);
or U4095 (N_4095,N_3748,N_3817);
nand U4096 (N_4096,N_3745,N_3838);
nor U4097 (N_4097,N_3725,N_3897);
xnor U4098 (N_4098,N_3808,N_3896);
nor U4099 (N_4099,N_3526,N_3925);
or U4100 (N_4100,N_3929,N_3574);
nor U4101 (N_4101,N_3636,N_3747);
nand U4102 (N_4102,N_3911,N_3894);
or U4103 (N_4103,N_3722,N_3856);
or U4104 (N_4104,N_3786,N_3916);
and U4105 (N_4105,N_3789,N_3988);
nand U4106 (N_4106,N_3996,N_3573);
or U4107 (N_4107,N_3752,N_3791);
nor U4108 (N_4108,N_3972,N_3827);
and U4109 (N_4109,N_3960,N_3906);
nand U4110 (N_4110,N_3589,N_3809);
xor U4111 (N_4111,N_3527,N_3763);
nand U4112 (N_4112,N_3797,N_3576);
nor U4113 (N_4113,N_3596,N_3937);
nor U4114 (N_4114,N_3532,N_3624);
nor U4115 (N_4115,N_3980,N_3820);
xnor U4116 (N_4116,N_3846,N_3770);
and U4117 (N_4117,N_3618,N_3967);
xnor U4118 (N_4118,N_3842,N_3687);
nand U4119 (N_4119,N_3691,N_3623);
or U4120 (N_4120,N_3771,N_3518);
and U4121 (N_4121,N_3768,N_3806);
and U4122 (N_4122,N_3974,N_3700);
nand U4123 (N_4123,N_3776,N_3830);
xnor U4124 (N_4124,N_3890,N_3843);
or U4125 (N_4125,N_3556,N_3551);
xor U4126 (N_4126,N_3831,N_3760);
nand U4127 (N_4127,N_3533,N_3577);
and U4128 (N_4128,N_3826,N_3767);
nand U4129 (N_4129,N_3948,N_3704);
nand U4130 (N_4130,N_3521,N_3530);
nor U4131 (N_4131,N_3565,N_3943);
and U4132 (N_4132,N_3799,N_3993);
and U4133 (N_4133,N_3516,N_3805);
nor U4134 (N_4134,N_3922,N_3587);
nand U4135 (N_4135,N_3907,N_3697);
xor U4136 (N_4136,N_3884,N_3947);
nand U4137 (N_4137,N_3761,N_3878);
nor U4138 (N_4138,N_3868,N_3938);
xor U4139 (N_4139,N_3865,N_3909);
nand U4140 (N_4140,N_3944,N_3588);
nand U4141 (N_4141,N_3832,N_3955);
and U4142 (N_4142,N_3581,N_3773);
and U4143 (N_4143,N_3713,N_3816);
nand U4144 (N_4144,N_3595,N_3848);
nand U4145 (N_4145,N_3536,N_3541);
or U4146 (N_4146,N_3655,N_3613);
and U4147 (N_4147,N_3645,N_3515);
and U4148 (N_4148,N_3534,N_3887);
or U4149 (N_4149,N_3857,N_3818);
nor U4150 (N_4150,N_3695,N_3932);
xor U4151 (N_4151,N_3940,N_3668);
nand U4152 (N_4152,N_3627,N_3506);
nor U4153 (N_4153,N_3570,N_3755);
or U4154 (N_4154,N_3688,N_3921);
or U4155 (N_4155,N_3735,N_3736);
and U4156 (N_4156,N_3597,N_3550);
and U4157 (N_4157,N_3762,N_3790);
and U4158 (N_4158,N_3607,N_3862);
and U4159 (N_4159,N_3571,N_3629);
or U4160 (N_4160,N_3997,N_3705);
nand U4161 (N_4161,N_3680,N_3698);
nand U4162 (N_4162,N_3702,N_3987);
nor U4163 (N_4163,N_3895,N_3777);
and U4164 (N_4164,N_3893,N_3501);
nor U4165 (N_4165,N_3968,N_3913);
or U4166 (N_4166,N_3870,N_3958);
nand U4167 (N_4167,N_3977,N_3510);
nor U4168 (N_4168,N_3919,N_3741);
nor U4169 (N_4169,N_3824,N_3615);
nand U4170 (N_4170,N_3866,N_3883);
nor U4171 (N_4171,N_3975,N_3899);
or U4172 (N_4172,N_3900,N_3600);
nor U4173 (N_4173,N_3670,N_3528);
and U4174 (N_4174,N_3540,N_3811);
nor U4175 (N_4175,N_3847,N_3685);
nand U4176 (N_4176,N_3535,N_3957);
nor U4177 (N_4177,N_3991,N_3539);
and U4178 (N_4178,N_3711,N_3653);
or U4179 (N_4179,N_3990,N_3508);
nand U4180 (N_4180,N_3658,N_3966);
or U4181 (N_4181,N_3759,N_3781);
or U4182 (N_4182,N_3679,N_3605);
nand U4183 (N_4183,N_3608,N_3656);
and U4184 (N_4184,N_3724,N_3959);
nand U4185 (N_4185,N_3619,N_3710);
xnor U4186 (N_4186,N_3969,N_3578);
nand U4187 (N_4187,N_3644,N_3675);
nor U4188 (N_4188,N_3739,N_3603);
or U4189 (N_4189,N_3659,N_3754);
nand U4190 (N_4190,N_3924,N_3845);
nor U4191 (N_4191,N_3729,N_3637);
nor U4192 (N_4192,N_3849,N_3671);
or U4193 (N_4193,N_3978,N_3590);
or U4194 (N_4194,N_3643,N_3989);
nand U4195 (N_4195,N_3731,N_3649);
or U4196 (N_4196,N_3693,N_3564);
and U4197 (N_4197,N_3640,N_3837);
nand U4198 (N_4198,N_3728,N_3889);
and U4199 (N_4199,N_3723,N_3769);
xnor U4200 (N_4200,N_3626,N_3617);
nand U4201 (N_4201,N_3520,N_3661);
and U4202 (N_4202,N_3901,N_3639);
and U4203 (N_4203,N_3707,N_3746);
nor U4204 (N_4204,N_3998,N_3926);
or U4205 (N_4205,N_3514,N_3794);
or U4206 (N_4206,N_3953,N_3931);
nand U4207 (N_4207,N_3563,N_3523);
xor U4208 (N_4208,N_3871,N_3971);
or U4209 (N_4209,N_3952,N_3819);
or U4210 (N_4210,N_3610,N_3861);
nor U4211 (N_4211,N_3647,N_3678);
or U4212 (N_4212,N_3542,N_3650);
and U4213 (N_4213,N_3945,N_3858);
and U4214 (N_4214,N_3800,N_3785);
and U4215 (N_4215,N_3620,N_3784);
xor U4216 (N_4216,N_3885,N_3625);
xnor U4217 (N_4217,N_3706,N_3715);
or U4218 (N_4218,N_3681,N_3793);
or U4219 (N_4219,N_3852,N_3604);
xnor U4220 (N_4220,N_3756,N_3839);
nor U4221 (N_4221,N_3524,N_3905);
nor U4222 (N_4222,N_3779,N_3585);
nor U4223 (N_4223,N_3592,N_3712);
nand U4224 (N_4224,N_3676,N_3863);
or U4225 (N_4225,N_3841,N_3981);
xnor U4226 (N_4226,N_3502,N_3611);
or U4227 (N_4227,N_3810,N_3727);
or U4228 (N_4228,N_3941,N_3543);
or U4229 (N_4229,N_3802,N_3660);
nand U4230 (N_4230,N_3548,N_3699);
nand U4231 (N_4231,N_3721,N_3872);
nand U4232 (N_4232,N_3719,N_3912);
or U4233 (N_4233,N_3677,N_3646);
nor U4234 (N_4234,N_3575,N_3753);
nand U4235 (N_4235,N_3979,N_3569);
xnor U4236 (N_4236,N_3882,N_3641);
and U4237 (N_4237,N_3566,N_3984);
nor U4238 (N_4238,N_3886,N_3673);
nand U4239 (N_4239,N_3825,N_3982);
nor U4240 (N_4240,N_3796,N_3692);
and U4241 (N_4241,N_3879,N_3772);
or U4242 (N_4242,N_3853,N_3936);
or U4243 (N_4243,N_3829,N_3933);
xnor U4244 (N_4244,N_3630,N_3609);
and U4245 (N_4245,N_3599,N_3757);
and U4246 (N_4246,N_3815,N_3778);
nor U4247 (N_4247,N_3934,N_3703);
and U4248 (N_4248,N_3823,N_3538);
nand U4249 (N_4249,N_3635,N_3690);
nand U4250 (N_4250,N_3791,N_3767);
or U4251 (N_4251,N_3998,N_3753);
and U4252 (N_4252,N_3762,N_3812);
or U4253 (N_4253,N_3884,N_3614);
nand U4254 (N_4254,N_3753,N_3600);
nor U4255 (N_4255,N_3759,N_3895);
xnor U4256 (N_4256,N_3933,N_3567);
nand U4257 (N_4257,N_3683,N_3508);
nand U4258 (N_4258,N_3717,N_3577);
nor U4259 (N_4259,N_3624,N_3824);
nand U4260 (N_4260,N_3967,N_3643);
and U4261 (N_4261,N_3961,N_3756);
nor U4262 (N_4262,N_3995,N_3891);
or U4263 (N_4263,N_3796,N_3682);
xnor U4264 (N_4264,N_3712,N_3908);
xor U4265 (N_4265,N_3593,N_3942);
and U4266 (N_4266,N_3811,N_3670);
xor U4267 (N_4267,N_3784,N_3906);
and U4268 (N_4268,N_3759,N_3692);
or U4269 (N_4269,N_3977,N_3743);
or U4270 (N_4270,N_3807,N_3729);
or U4271 (N_4271,N_3927,N_3737);
and U4272 (N_4272,N_3507,N_3868);
nor U4273 (N_4273,N_3995,N_3635);
or U4274 (N_4274,N_3758,N_3718);
or U4275 (N_4275,N_3712,N_3533);
nor U4276 (N_4276,N_3848,N_3978);
or U4277 (N_4277,N_3699,N_3655);
or U4278 (N_4278,N_3585,N_3580);
nand U4279 (N_4279,N_3613,N_3771);
xnor U4280 (N_4280,N_3789,N_3621);
or U4281 (N_4281,N_3777,N_3862);
nand U4282 (N_4282,N_3658,N_3963);
and U4283 (N_4283,N_3621,N_3974);
or U4284 (N_4284,N_3702,N_3819);
nor U4285 (N_4285,N_3815,N_3565);
and U4286 (N_4286,N_3786,N_3852);
nor U4287 (N_4287,N_3777,N_3893);
or U4288 (N_4288,N_3896,N_3859);
nand U4289 (N_4289,N_3546,N_3571);
and U4290 (N_4290,N_3887,N_3717);
nor U4291 (N_4291,N_3711,N_3789);
nand U4292 (N_4292,N_3980,N_3795);
nand U4293 (N_4293,N_3536,N_3854);
or U4294 (N_4294,N_3736,N_3561);
xnor U4295 (N_4295,N_3743,N_3586);
or U4296 (N_4296,N_3614,N_3993);
nand U4297 (N_4297,N_3622,N_3584);
nor U4298 (N_4298,N_3506,N_3921);
or U4299 (N_4299,N_3798,N_3857);
xor U4300 (N_4300,N_3709,N_3666);
nor U4301 (N_4301,N_3721,N_3949);
and U4302 (N_4302,N_3625,N_3758);
nand U4303 (N_4303,N_3623,N_3961);
xor U4304 (N_4304,N_3672,N_3682);
nor U4305 (N_4305,N_3752,N_3641);
xnor U4306 (N_4306,N_3757,N_3805);
or U4307 (N_4307,N_3795,N_3838);
nor U4308 (N_4308,N_3976,N_3592);
and U4309 (N_4309,N_3955,N_3614);
nand U4310 (N_4310,N_3682,N_3913);
nand U4311 (N_4311,N_3671,N_3969);
nor U4312 (N_4312,N_3563,N_3833);
nor U4313 (N_4313,N_3587,N_3556);
and U4314 (N_4314,N_3505,N_3628);
or U4315 (N_4315,N_3595,N_3686);
nor U4316 (N_4316,N_3778,N_3709);
nor U4317 (N_4317,N_3695,N_3675);
and U4318 (N_4318,N_3505,N_3731);
nor U4319 (N_4319,N_3545,N_3543);
and U4320 (N_4320,N_3607,N_3684);
nand U4321 (N_4321,N_3703,N_3621);
and U4322 (N_4322,N_3703,N_3557);
and U4323 (N_4323,N_3964,N_3727);
and U4324 (N_4324,N_3783,N_3929);
and U4325 (N_4325,N_3870,N_3975);
and U4326 (N_4326,N_3728,N_3960);
nand U4327 (N_4327,N_3814,N_3980);
and U4328 (N_4328,N_3966,N_3839);
and U4329 (N_4329,N_3802,N_3911);
and U4330 (N_4330,N_3688,N_3611);
nand U4331 (N_4331,N_3767,N_3922);
and U4332 (N_4332,N_3994,N_3981);
or U4333 (N_4333,N_3620,N_3785);
nor U4334 (N_4334,N_3536,N_3570);
and U4335 (N_4335,N_3644,N_3566);
or U4336 (N_4336,N_3786,N_3674);
and U4337 (N_4337,N_3786,N_3991);
or U4338 (N_4338,N_3589,N_3673);
nand U4339 (N_4339,N_3654,N_3589);
nor U4340 (N_4340,N_3881,N_3986);
and U4341 (N_4341,N_3608,N_3699);
nor U4342 (N_4342,N_3684,N_3892);
and U4343 (N_4343,N_3502,N_3535);
nand U4344 (N_4344,N_3632,N_3550);
and U4345 (N_4345,N_3872,N_3826);
nand U4346 (N_4346,N_3843,N_3546);
nand U4347 (N_4347,N_3551,N_3550);
nand U4348 (N_4348,N_3851,N_3949);
nand U4349 (N_4349,N_3993,N_3535);
nor U4350 (N_4350,N_3984,N_3669);
or U4351 (N_4351,N_3921,N_3650);
nor U4352 (N_4352,N_3687,N_3805);
and U4353 (N_4353,N_3819,N_3997);
xor U4354 (N_4354,N_3802,N_3782);
nor U4355 (N_4355,N_3714,N_3821);
or U4356 (N_4356,N_3984,N_3707);
and U4357 (N_4357,N_3752,N_3533);
or U4358 (N_4358,N_3971,N_3885);
nor U4359 (N_4359,N_3578,N_3755);
xor U4360 (N_4360,N_3830,N_3908);
and U4361 (N_4361,N_3575,N_3783);
and U4362 (N_4362,N_3583,N_3655);
or U4363 (N_4363,N_3868,N_3677);
or U4364 (N_4364,N_3513,N_3744);
or U4365 (N_4365,N_3654,N_3802);
or U4366 (N_4366,N_3835,N_3677);
nand U4367 (N_4367,N_3647,N_3853);
and U4368 (N_4368,N_3776,N_3940);
and U4369 (N_4369,N_3713,N_3763);
nand U4370 (N_4370,N_3662,N_3763);
and U4371 (N_4371,N_3929,N_3983);
and U4372 (N_4372,N_3590,N_3764);
and U4373 (N_4373,N_3710,N_3500);
or U4374 (N_4374,N_3566,N_3561);
nand U4375 (N_4375,N_3804,N_3859);
xor U4376 (N_4376,N_3840,N_3694);
xnor U4377 (N_4377,N_3841,N_3577);
and U4378 (N_4378,N_3808,N_3824);
and U4379 (N_4379,N_3737,N_3526);
xnor U4380 (N_4380,N_3822,N_3875);
xnor U4381 (N_4381,N_3592,N_3564);
or U4382 (N_4382,N_3681,N_3850);
nor U4383 (N_4383,N_3714,N_3869);
nand U4384 (N_4384,N_3628,N_3583);
or U4385 (N_4385,N_3801,N_3714);
or U4386 (N_4386,N_3794,N_3768);
nor U4387 (N_4387,N_3506,N_3734);
and U4388 (N_4388,N_3886,N_3706);
xor U4389 (N_4389,N_3577,N_3883);
or U4390 (N_4390,N_3835,N_3753);
xor U4391 (N_4391,N_3935,N_3622);
nand U4392 (N_4392,N_3875,N_3613);
or U4393 (N_4393,N_3709,N_3573);
and U4394 (N_4394,N_3913,N_3847);
nor U4395 (N_4395,N_3942,N_3940);
and U4396 (N_4396,N_3558,N_3739);
nand U4397 (N_4397,N_3882,N_3739);
or U4398 (N_4398,N_3809,N_3609);
and U4399 (N_4399,N_3785,N_3810);
nor U4400 (N_4400,N_3608,N_3504);
nor U4401 (N_4401,N_3650,N_3884);
xnor U4402 (N_4402,N_3988,N_3839);
and U4403 (N_4403,N_3640,N_3767);
and U4404 (N_4404,N_3699,N_3816);
xnor U4405 (N_4405,N_3510,N_3833);
nand U4406 (N_4406,N_3894,N_3788);
and U4407 (N_4407,N_3511,N_3799);
nand U4408 (N_4408,N_3822,N_3974);
nor U4409 (N_4409,N_3854,N_3648);
or U4410 (N_4410,N_3962,N_3796);
xor U4411 (N_4411,N_3861,N_3752);
xor U4412 (N_4412,N_3989,N_3716);
xnor U4413 (N_4413,N_3634,N_3958);
or U4414 (N_4414,N_3606,N_3596);
nand U4415 (N_4415,N_3547,N_3925);
nor U4416 (N_4416,N_3906,N_3980);
or U4417 (N_4417,N_3836,N_3703);
nand U4418 (N_4418,N_3529,N_3998);
and U4419 (N_4419,N_3763,N_3992);
or U4420 (N_4420,N_3895,N_3782);
and U4421 (N_4421,N_3605,N_3683);
xnor U4422 (N_4422,N_3602,N_3630);
xnor U4423 (N_4423,N_3717,N_3595);
or U4424 (N_4424,N_3879,N_3543);
nand U4425 (N_4425,N_3785,N_3963);
and U4426 (N_4426,N_3755,N_3579);
and U4427 (N_4427,N_3781,N_3679);
xnor U4428 (N_4428,N_3524,N_3645);
nor U4429 (N_4429,N_3821,N_3910);
or U4430 (N_4430,N_3941,N_3644);
and U4431 (N_4431,N_3683,N_3951);
nand U4432 (N_4432,N_3711,N_3889);
and U4433 (N_4433,N_3638,N_3630);
or U4434 (N_4434,N_3757,N_3723);
nand U4435 (N_4435,N_3862,N_3576);
nand U4436 (N_4436,N_3623,N_3519);
or U4437 (N_4437,N_3818,N_3883);
or U4438 (N_4438,N_3929,N_3533);
xnor U4439 (N_4439,N_3743,N_3838);
nor U4440 (N_4440,N_3512,N_3764);
nand U4441 (N_4441,N_3903,N_3867);
or U4442 (N_4442,N_3757,N_3873);
or U4443 (N_4443,N_3664,N_3791);
and U4444 (N_4444,N_3524,N_3640);
nor U4445 (N_4445,N_3954,N_3992);
and U4446 (N_4446,N_3607,N_3963);
xor U4447 (N_4447,N_3910,N_3662);
nor U4448 (N_4448,N_3976,N_3944);
nand U4449 (N_4449,N_3749,N_3914);
nand U4450 (N_4450,N_3833,N_3660);
xor U4451 (N_4451,N_3630,N_3681);
and U4452 (N_4452,N_3711,N_3684);
xor U4453 (N_4453,N_3820,N_3743);
nor U4454 (N_4454,N_3917,N_3714);
and U4455 (N_4455,N_3954,N_3659);
and U4456 (N_4456,N_3676,N_3926);
nand U4457 (N_4457,N_3567,N_3930);
nand U4458 (N_4458,N_3823,N_3580);
nand U4459 (N_4459,N_3906,N_3870);
or U4460 (N_4460,N_3777,N_3759);
nor U4461 (N_4461,N_3815,N_3648);
and U4462 (N_4462,N_3676,N_3690);
xor U4463 (N_4463,N_3831,N_3505);
nand U4464 (N_4464,N_3792,N_3673);
and U4465 (N_4465,N_3512,N_3573);
xnor U4466 (N_4466,N_3992,N_3648);
nand U4467 (N_4467,N_3662,N_3634);
or U4468 (N_4468,N_3925,N_3604);
and U4469 (N_4469,N_3871,N_3864);
nand U4470 (N_4470,N_3983,N_3836);
or U4471 (N_4471,N_3500,N_3575);
and U4472 (N_4472,N_3573,N_3730);
or U4473 (N_4473,N_3842,N_3666);
nor U4474 (N_4474,N_3830,N_3724);
nand U4475 (N_4475,N_3961,N_3768);
nand U4476 (N_4476,N_3876,N_3995);
nand U4477 (N_4477,N_3532,N_3653);
or U4478 (N_4478,N_3500,N_3763);
or U4479 (N_4479,N_3839,N_3582);
and U4480 (N_4480,N_3828,N_3946);
and U4481 (N_4481,N_3663,N_3585);
nand U4482 (N_4482,N_3746,N_3786);
xnor U4483 (N_4483,N_3766,N_3571);
nor U4484 (N_4484,N_3722,N_3756);
and U4485 (N_4485,N_3551,N_3623);
or U4486 (N_4486,N_3956,N_3977);
and U4487 (N_4487,N_3718,N_3589);
xor U4488 (N_4488,N_3639,N_3719);
xor U4489 (N_4489,N_3932,N_3975);
or U4490 (N_4490,N_3868,N_3983);
or U4491 (N_4491,N_3501,N_3517);
nand U4492 (N_4492,N_3841,N_3976);
and U4493 (N_4493,N_3549,N_3909);
xnor U4494 (N_4494,N_3954,N_3857);
nor U4495 (N_4495,N_3620,N_3721);
or U4496 (N_4496,N_3953,N_3629);
or U4497 (N_4497,N_3627,N_3521);
nand U4498 (N_4498,N_3875,N_3719);
nor U4499 (N_4499,N_3859,N_3772);
nand U4500 (N_4500,N_4218,N_4487);
xor U4501 (N_4501,N_4355,N_4426);
nand U4502 (N_4502,N_4269,N_4351);
nand U4503 (N_4503,N_4094,N_4195);
or U4504 (N_4504,N_4140,N_4170);
or U4505 (N_4505,N_4276,N_4247);
or U4506 (N_4506,N_4145,N_4138);
and U4507 (N_4507,N_4229,N_4273);
xor U4508 (N_4508,N_4440,N_4163);
and U4509 (N_4509,N_4471,N_4271);
and U4510 (N_4510,N_4021,N_4046);
xor U4511 (N_4511,N_4244,N_4014);
and U4512 (N_4512,N_4016,N_4148);
or U4513 (N_4513,N_4442,N_4408);
nor U4514 (N_4514,N_4372,N_4431);
xor U4515 (N_4515,N_4373,N_4449);
or U4516 (N_4516,N_4039,N_4209);
nor U4517 (N_4517,N_4083,N_4305);
nor U4518 (N_4518,N_4360,N_4074);
nor U4519 (N_4519,N_4466,N_4425);
nor U4520 (N_4520,N_4378,N_4320);
or U4521 (N_4521,N_4042,N_4026);
or U4522 (N_4522,N_4230,N_4226);
nand U4523 (N_4523,N_4497,N_4142);
and U4524 (N_4524,N_4203,N_4322);
nand U4525 (N_4525,N_4369,N_4422);
nor U4526 (N_4526,N_4296,N_4479);
or U4527 (N_4527,N_4265,N_4285);
and U4528 (N_4528,N_4240,N_4396);
or U4529 (N_4529,N_4414,N_4109);
or U4530 (N_4530,N_4091,N_4491);
nor U4531 (N_4531,N_4312,N_4224);
xnor U4532 (N_4532,N_4190,N_4119);
xor U4533 (N_4533,N_4153,N_4188);
nand U4534 (N_4534,N_4353,N_4071);
and U4535 (N_4535,N_4358,N_4111);
nor U4536 (N_4536,N_4388,N_4079);
nand U4537 (N_4537,N_4473,N_4059);
and U4538 (N_4538,N_4291,N_4318);
nor U4539 (N_4539,N_4215,N_4084);
xnor U4540 (N_4540,N_4401,N_4420);
nor U4541 (N_4541,N_4376,N_4185);
nor U4542 (N_4542,N_4100,N_4087);
and U4543 (N_4543,N_4453,N_4356);
nor U4544 (N_4544,N_4311,N_4278);
and U4545 (N_4545,N_4104,N_4354);
nor U4546 (N_4546,N_4078,N_4151);
or U4547 (N_4547,N_4448,N_4347);
nand U4548 (N_4548,N_4191,N_4266);
nand U4549 (N_4549,N_4259,N_4030);
and U4550 (N_4550,N_4202,N_4267);
or U4551 (N_4551,N_4122,N_4001);
nand U4552 (N_4552,N_4346,N_4136);
nor U4553 (N_4553,N_4162,N_4103);
nor U4554 (N_4554,N_4044,N_4261);
or U4555 (N_4555,N_4382,N_4018);
nor U4556 (N_4556,N_4054,N_4464);
nand U4557 (N_4557,N_4306,N_4057);
nor U4558 (N_4558,N_4424,N_4033);
nand U4559 (N_4559,N_4069,N_4410);
xnor U4560 (N_4560,N_4475,N_4330);
or U4561 (N_4561,N_4251,N_4255);
and U4562 (N_4562,N_4027,N_4254);
nand U4563 (N_4563,N_4379,N_4152);
or U4564 (N_4564,N_4395,N_4117);
and U4565 (N_4565,N_4297,N_4436);
nor U4566 (N_4566,N_4061,N_4234);
xnor U4567 (N_4567,N_4416,N_4433);
nor U4568 (N_4568,N_4031,N_4008);
nand U4569 (N_4569,N_4300,N_4304);
and U4570 (N_4570,N_4315,N_4004);
nor U4571 (N_4571,N_4493,N_4349);
nor U4572 (N_4572,N_4238,N_4051);
nand U4573 (N_4573,N_4309,N_4052);
nand U4574 (N_4574,N_4387,N_4478);
or U4575 (N_4575,N_4200,N_4490);
nand U4576 (N_4576,N_4256,N_4066);
or U4577 (N_4577,N_4280,N_4384);
nor U4578 (N_4578,N_4193,N_4221);
nor U4579 (N_4579,N_4263,N_4481);
and U4580 (N_4580,N_4187,N_4303);
or U4581 (N_4581,N_4123,N_4390);
nor U4582 (N_4582,N_4035,N_4105);
and U4583 (N_4583,N_4386,N_4038);
or U4584 (N_4584,N_4468,N_4321);
xnor U4585 (N_4585,N_4367,N_4099);
nand U4586 (N_4586,N_4411,N_4380);
nor U4587 (N_4587,N_4129,N_4277);
or U4588 (N_4588,N_4456,N_4338);
nand U4589 (N_4589,N_4150,N_4437);
and U4590 (N_4590,N_4486,N_4025);
or U4591 (N_4591,N_4498,N_4371);
nor U4592 (N_4592,N_4462,N_4310);
or U4593 (N_4593,N_4370,N_4428);
nand U4594 (N_4594,N_4043,N_4060);
xor U4595 (N_4595,N_4146,N_4272);
and U4596 (N_4596,N_4154,N_4217);
and U4597 (N_4597,N_4093,N_4270);
xor U4598 (N_4598,N_4461,N_4308);
or U4599 (N_4599,N_4144,N_4298);
nor U4600 (N_4600,N_4392,N_4460);
nor U4601 (N_4601,N_4295,N_4333);
nor U4602 (N_4602,N_4458,N_4045);
or U4603 (N_4603,N_4164,N_4365);
or U4604 (N_4604,N_4492,N_4115);
or U4605 (N_4605,N_4274,N_4106);
and U4606 (N_4606,N_4173,N_4455);
nor U4607 (N_4607,N_4081,N_4036);
nand U4608 (N_4608,N_4000,N_4143);
nand U4609 (N_4609,N_4214,N_4092);
nand U4610 (N_4610,N_4124,N_4292);
xor U4611 (N_4611,N_4324,N_4350);
xor U4612 (N_4612,N_4332,N_4257);
or U4613 (N_4613,N_4107,N_4239);
or U4614 (N_4614,N_4198,N_4262);
and U4615 (N_4615,N_4137,N_4417);
nand U4616 (N_4616,N_4007,N_4463);
nand U4617 (N_4617,N_4053,N_4469);
or U4618 (N_4618,N_4113,N_4070);
nand U4619 (N_4619,N_4037,N_4086);
or U4620 (N_4620,N_4389,N_4180);
or U4621 (N_4621,N_4488,N_4245);
and U4622 (N_4622,N_4192,N_4169);
nor U4623 (N_4623,N_4160,N_4445);
nor U4624 (N_4624,N_4116,N_4364);
nor U4625 (N_4625,N_4208,N_4009);
and U4626 (N_4626,N_4253,N_4077);
or U4627 (N_4627,N_4062,N_4006);
or U4628 (N_4628,N_4194,N_4327);
nor U4629 (N_4629,N_4340,N_4141);
nand U4630 (N_4630,N_4275,N_4168);
or U4631 (N_4631,N_4206,N_4236);
and U4632 (N_4632,N_4454,N_4155);
or U4633 (N_4633,N_4423,N_4182);
nor U4634 (N_4634,N_4472,N_4334);
or U4635 (N_4635,N_4049,N_4176);
nand U4636 (N_4636,N_4178,N_4175);
nand U4637 (N_4637,N_4363,N_4485);
nor U4638 (N_4638,N_4406,N_4028);
nand U4639 (N_4639,N_4325,N_4063);
nand U4640 (N_4640,N_4480,N_4073);
nor U4641 (N_4641,N_4199,N_4402);
and U4642 (N_4642,N_4301,N_4098);
xor U4643 (N_4643,N_4494,N_4213);
xor U4644 (N_4644,N_4316,N_4344);
or U4645 (N_4645,N_4211,N_4210);
nor U4646 (N_4646,N_4432,N_4288);
and U4647 (N_4647,N_4065,N_4101);
nor U4648 (N_4648,N_4149,N_4317);
nand U4649 (N_4649,N_4232,N_4383);
xnor U4650 (N_4650,N_4375,N_4393);
or U4651 (N_4651,N_4147,N_4055);
and U4652 (N_4652,N_4096,N_4366);
nor U4653 (N_4653,N_4158,N_4450);
and U4654 (N_4654,N_4452,N_4017);
or U4655 (N_4655,N_4075,N_4336);
nand U4656 (N_4656,N_4499,N_4430);
nand U4657 (N_4657,N_4249,N_4237);
or U4658 (N_4658,N_4201,N_4076);
nor U4659 (N_4659,N_4407,N_4241);
and U4660 (N_4660,N_4451,N_4120);
and U4661 (N_4661,N_4032,N_4484);
nand U4662 (N_4662,N_4398,N_4342);
xnor U4663 (N_4663,N_4228,N_4112);
and U4664 (N_4664,N_4345,N_4167);
nor U4665 (N_4665,N_4482,N_4319);
nor U4666 (N_4666,N_4391,N_4118);
nor U4667 (N_4667,N_4013,N_4446);
and U4668 (N_4668,N_4283,N_4010);
nand U4669 (N_4669,N_4467,N_4293);
nor U4670 (N_4670,N_4132,N_4290);
nor U4671 (N_4671,N_4231,N_4177);
nor U4672 (N_4672,N_4284,N_4068);
nand U4673 (N_4673,N_4405,N_4216);
and U4674 (N_4674,N_4415,N_4050);
or U4675 (N_4675,N_4156,N_4429);
nand U4676 (N_4676,N_4385,N_4323);
nand U4677 (N_4677,N_4368,N_4281);
or U4678 (N_4678,N_4447,N_4307);
nand U4679 (N_4679,N_4020,N_4166);
xor U4680 (N_4680,N_4268,N_4012);
nand U4681 (N_4681,N_4029,N_4339);
nand U4682 (N_4682,N_4067,N_4225);
nor U4683 (N_4683,N_4443,N_4034);
and U4684 (N_4684,N_4047,N_4089);
or U4685 (N_4685,N_4496,N_4418);
or U4686 (N_4686,N_4212,N_4130);
nor U4687 (N_4687,N_4181,N_4427);
nor U4688 (N_4688,N_4419,N_4197);
nand U4689 (N_4689,N_4331,N_4082);
or U4690 (N_4690,N_4474,N_4127);
and U4691 (N_4691,N_4003,N_4489);
nor U4692 (N_4692,N_4361,N_4457);
nor U4693 (N_4693,N_4223,N_4222);
nor U4694 (N_4694,N_4134,N_4056);
nor U4695 (N_4695,N_4343,N_4439);
xor U4696 (N_4696,N_4441,N_4023);
nand U4697 (N_4697,N_4205,N_4337);
nand U4698 (N_4698,N_4131,N_4133);
and U4699 (N_4699,N_4097,N_4302);
nor U4700 (N_4700,N_4243,N_4348);
and U4701 (N_4701,N_4495,N_4359);
or U4702 (N_4702,N_4048,N_4041);
nor U4703 (N_4703,N_4444,N_4326);
nor U4704 (N_4704,N_4220,N_4328);
and U4705 (N_4705,N_4121,N_4183);
nand U4706 (N_4706,N_4090,N_4072);
or U4707 (N_4707,N_4362,N_4135);
nor U4708 (N_4708,N_4011,N_4381);
nor U4709 (N_4709,N_4477,N_4250);
nand U4710 (N_4710,N_4314,N_4329);
nand U4711 (N_4711,N_4219,N_4260);
nand U4712 (N_4712,N_4352,N_4126);
or U4713 (N_4713,N_4299,N_4024);
and U4714 (N_4714,N_4171,N_4357);
or U4715 (N_4715,N_4080,N_4470);
nor U4716 (N_4716,N_4196,N_4264);
nor U4717 (N_4717,N_4374,N_4279);
and U4718 (N_4718,N_4412,N_4227);
and U4719 (N_4719,N_4108,N_4161);
nand U4720 (N_4720,N_4242,N_4159);
xnor U4721 (N_4721,N_4413,N_4040);
nand U4722 (N_4722,N_4128,N_4400);
and U4723 (N_4723,N_4022,N_4174);
and U4724 (N_4724,N_4172,N_4102);
or U4725 (N_4725,N_4005,N_4397);
and U4726 (N_4726,N_4287,N_4313);
and U4727 (N_4727,N_4438,N_4258);
xnor U4728 (N_4728,N_4335,N_4204);
or U4729 (N_4729,N_4286,N_4341);
nand U4730 (N_4730,N_4483,N_4282);
and U4731 (N_4731,N_4125,N_4465);
or U4732 (N_4732,N_4246,N_4435);
nor U4733 (N_4733,N_4088,N_4235);
and U4734 (N_4734,N_4409,N_4186);
nor U4735 (N_4735,N_4095,N_4404);
nor U4736 (N_4736,N_4085,N_4233);
xor U4737 (N_4737,N_4403,N_4189);
or U4738 (N_4738,N_4064,N_4015);
nand U4739 (N_4739,N_4252,N_4184);
nor U4740 (N_4740,N_4248,N_4165);
nand U4741 (N_4741,N_4421,N_4114);
nand U4742 (N_4742,N_4459,N_4394);
and U4743 (N_4743,N_4179,N_4399);
or U4744 (N_4744,N_4002,N_4157);
or U4745 (N_4745,N_4476,N_4058);
nand U4746 (N_4746,N_4110,N_4019);
nor U4747 (N_4747,N_4207,N_4289);
xor U4748 (N_4748,N_4377,N_4139);
and U4749 (N_4749,N_4434,N_4294);
xnor U4750 (N_4750,N_4448,N_4131);
xor U4751 (N_4751,N_4187,N_4240);
nand U4752 (N_4752,N_4130,N_4385);
nand U4753 (N_4753,N_4013,N_4457);
or U4754 (N_4754,N_4237,N_4153);
nor U4755 (N_4755,N_4057,N_4033);
nor U4756 (N_4756,N_4344,N_4427);
nand U4757 (N_4757,N_4293,N_4056);
and U4758 (N_4758,N_4223,N_4228);
xor U4759 (N_4759,N_4240,N_4099);
nand U4760 (N_4760,N_4415,N_4151);
or U4761 (N_4761,N_4033,N_4279);
nor U4762 (N_4762,N_4004,N_4485);
and U4763 (N_4763,N_4263,N_4264);
nor U4764 (N_4764,N_4385,N_4111);
and U4765 (N_4765,N_4332,N_4054);
nand U4766 (N_4766,N_4401,N_4448);
xnor U4767 (N_4767,N_4435,N_4168);
or U4768 (N_4768,N_4343,N_4204);
and U4769 (N_4769,N_4049,N_4253);
and U4770 (N_4770,N_4236,N_4190);
and U4771 (N_4771,N_4263,N_4031);
nand U4772 (N_4772,N_4295,N_4445);
or U4773 (N_4773,N_4333,N_4216);
nand U4774 (N_4774,N_4291,N_4207);
nor U4775 (N_4775,N_4228,N_4044);
xnor U4776 (N_4776,N_4325,N_4275);
nand U4777 (N_4777,N_4265,N_4166);
or U4778 (N_4778,N_4273,N_4050);
nor U4779 (N_4779,N_4318,N_4086);
or U4780 (N_4780,N_4374,N_4498);
and U4781 (N_4781,N_4212,N_4105);
nor U4782 (N_4782,N_4292,N_4485);
and U4783 (N_4783,N_4340,N_4476);
nand U4784 (N_4784,N_4461,N_4236);
nand U4785 (N_4785,N_4312,N_4385);
nand U4786 (N_4786,N_4260,N_4203);
xnor U4787 (N_4787,N_4222,N_4169);
xor U4788 (N_4788,N_4018,N_4276);
nand U4789 (N_4789,N_4003,N_4416);
nand U4790 (N_4790,N_4332,N_4032);
and U4791 (N_4791,N_4372,N_4226);
or U4792 (N_4792,N_4268,N_4277);
and U4793 (N_4793,N_4197,N_4251);
or U4794 (N_4794,N_4274,N_4332);
nand U4795 (N_4795,N_4213,N_4409);
or U4796 (N_4796,N_4080,N_4214);
nand U4797 (N_4797,N_4430,N_4216);
and U4798 (N_4798,N_4378,N_4309);
or U4799 (N_4799,N_4260,N_4160);
or U4800 (N_4800,N_4298,N_4171);
nand U4801 (N_4801,N_4288,N_4418);
and U4802 (N_4802,N_4454,N_4494);
nand U4803 (N_4803,N_4348,N_4334);
and U4804 (N_4804,N_4240,N_4468);
or U4805 (N_4805,N_4298,N_4351);
and U4806 (N_4806,N_4306,N_4366);
nor U4807 (N_4807,N_4458,N_4049);
or U4808 (N_4808,N_4185,N_4062);
or U4809 (N_4809,N_4055,N_4424);
nand U4810 (N_4810,N_4011,N_4356);
nor U4811 (N_4811,N_4311,N_4222);
nor U4812 (N_4812,N_4373,N_4367);
nor U4813 (N_4813,N_4326,N_4202);
or U4814 (N_4814,N_4206,N_4104);
or U4815 (N_4815,N_4254,N_4021);
xor U4816 (N_4816,N_4094,N_4333);
nor U4817 (N_4817,N_4492,N_4047);
xnor U4818 (N_4818,N_4364,N_4428);
and U4819 (N_4819,N_4459,N_4341);
and U4820 (N_4820,N_4293,N_4129);
or U4821 (N_4821,N_4312,N_4044);
and U4822 (N_4822,N_4353,N_4219);
nand U4823 (N_4823,N_4136,N_4258);
nand U4824 (N_4824,N_4402,N_4048);
nand U4825 (N_4825,N_4186,N_4404);
nor U4826 (N_4826,N_4155,N_4058);
nor U4827 (N_4827,N_4098,N_4381);
xor U4828 (N_4828,N_4050,N_4211);
and U4829 (N_4829,N_4282,N_4386);
nor U4830 (N_4830,N_4289,N_4341);
xnor U4831 (N_4831,N_4165,N_4094);
xnor U4832 (N_4832,N_4208,N_4178);
nand U4833 (N_4833,N_4438,N_4068);
and U4834 (N_4834,N_4216,N_4047);
or U4835 (N_4835,N_4281,N_4342);
xnor U4836 (N_4836,N_4111,N_4036);
xor U4837 (N_4837,N_4493,N_4412);
or U4838 (N_4838,N_4161,N_4051);
and U4839 (N_4839,N_4492,N_4176);
or U4840 (N_4840,N_4128,N_4343);
nor U4841 (N_4841,N_4346,N_4229);
or U4842 (N_4842,N_4097,N_4371);
and U4843 (N_4843,N_4483,N_4013);
or U4844 (N_4844,N_4164,N_4097);
nand U4845 (N_4845,N_4233,N_4246);
or U4846 (N_4846,N_4237,N_4187);
nand U4847 (N_4847,N_4256,N_4451);
nor U4848 (N_4848,N_4170,N_4430);
and U4849 (N_4849,N_4121,N_4377);
or U4850 (N_4850,N_4173,N_4318);
nor U4851 (N_4851,N_4292,N_4144);
nand U4852 (N_4852,N_4290,N_4498);
nand U4853 (N_4853,N_4182,N_4060);
and U4854 (N_4854,N_4192,N_4396);
or U4855 (N_4855,N_4463,N_4293);
and U4856 (N_4856,N_4054,N_4447);
nor U4857 (N_4857,N_4140,N_4220);
xor U4858 (N_4858,N_4208,N_4469);
nor U4859 (N_4859,N_4337,N_4393);
xor U4860 (N_4860,N_4139,N_4060);
nand U4861 (N_4861,N_4223,N_4149);
xor U4862 (N_4862,N_4333,N_4035);
nor U4863 (N_4863,N_4285,N_4456);
nand U4864 (N_4864,N_4335,N_4323);
xor U4865 (N_4865,N_4049,N_4111);
or U4866 (N_4866,N_4052,N_4400);
nor U4867 (N_4867,N_4265,N_4498);
nor U4868 (N_4868,N_4492,N_4437);
nor U4869 (N_4869,N_4350,N_4414);
nand U4870 (N_4870,N_4370,N_4028);
and U4871 (N_4871,N_4054,N_4213);
nor U4872 (N_4872,N_4290,N_4186);
and U4873 (N_4873,N_4070,N_4307);
and U4874 (N_4874,N_4052,N_4356);
xnor U4875 (N_4875,N_4207,N_4281);
or U4876 (N_4876,N_4351,N_4445);
nand U4877 (N_4877,N_4497,N_4293);
and U4878 (N_4878,N_4127,N_4133);
and U4879 (N_4879,N_4308,N_4194);
or U4880 (N_4880,N_4239,N_4143);
nand U4881 (N_4881,N_4445,N_4190);
nand U4882 (N_4882,N_4065,N_4405);
or U4883 (N_4883,N_4344,N_4477);
and U4884 (N_4884,N_4466,N_4327);
and U4885 (N_4885,N_4163,N_4067);
or U4886 (N_4886,N_4160,N_4271);
or U4887 (N_4887,N_4166,N_4248);
nand U4888 (N_4888,N_4492,N_4023);
nor U4889 (N_4889,N_4180,N_4343);
and U4890 (N_4890,N_4098,N_4297);
nand U4891 (N_4891,N_4222,N_4112);
and U4892 (N_4892,N_4017,N_4435);
nor U4893 (N_4893,N_4068,N_4339);
nor U4894 (N_4894,N_4192,N_4343);
nand U4895 (N_4895,N_4125,N_4048);
or U4896 (N_4896,N_4049,N_4387);
nand U4897 (N_4897,N_4093,N_4042);
and U4898 (N_4898,N_4325,N_4309);
nor U4899 (N_4899,N_4471,N_4202);
nor U4900 (N_4900,N_4354,N_4077);
and U4901 (N_4901,N_4264,N_4064);
or U4902 (N_4902,N_4422,N_4330);
and U4903 (N_4903,N_4347,N_4394);
or U4904 (N_4904,N_4339,N_4101);
nand U4905 (N_4905,N_4424,N_4075);
nor U4906 (N_4906,N_4355,N_4386);
nand U4907 (N_4907,N_4452,N_4377);
and U4908 (N_4908,N_4157,N_4332);
nand U4909 (N_4909,N_4414,N_4235);
or U4910 (N_4910,N_4315,N_4248);
or U4911 (N_4911,N_4333,N_4210);
nor U4912 (N_4912,N_4201,N_4040);
and U4913 (N_4913,N_4075,N_4240);
nor U4914 (N_4914,N_4294,N_4428);
and U4915 (N_4915,N_4350,N_4365);
or U4916 (N_4916,N_4299,N_4413);
nand U4917 (N_4917,N_4373,N_4191);
xnor U4918 (N_4918,N_4037,N_4124);
and U4919 (N_4919,N_4301,N_4144);
xnor U4920 (N_4920,N_4221,N_4487);
nor U4921 (N_4921,N_4429,N_4495);
nand U4922 (N_4922,N_4021,N_4419);
nor U4923 (N_4923,N_4049,N_4209);
nor U4924 (N_4924,N_4317,N_4326);
or U4925 (N_4925,N_4175,N_4463);
or U4926 (N_4926,N_4011,N_4478);
and U4927 (N_4927,N_4377,N_4346);
and U4928 (N_4928,N_4152,N_4378);
nand U4929 (N_4929,N_4144,N_4484);
or U4930 (N_4930,N_4447,N_4188);
or U4931 (N_4931,N_4260,N_4236);
and U4932 (N_4932,N_4393,N_4171);
nand U4933 (N_4933,N_4436,N_4412);
nand U4934 (N_4934,N_4018,N_4119);
or U4935 (N_4935,N_4400,N_4495);
xor U4936 (N_4936,N_4151,N_4030);
nand U4937 (N_4937,N_4195,N_4325);
nor U4938 (N_4938,N_4043,N_4356);
or U4939 (N_4939,N_4046,N_4414);
and U4940 (N_4940,N_4427,N_4304);
nor U4941 (N_4941,N_4354,N_4347);
xor U4942 (N_4942,N_4283,N_4482);
nand U4943 (N_4943,N_4223,N_4271);
or U4944 (N_4944,N_4490,N_4286);
xor U4945 (N_4945,N_4117,N_4339);
and U4946 (N_4946,N_4318,N_4141);
or U4947 (N_4947,N_4338,N_4199);
nand U4948 (N_4948,N_4111,N_4033);
nand U4949 (N_4949,N_4369,N_4127);
or U4950 (N_4950,N_4257,N_4105);
and U4951 (N_4951,N_4119,N_4221);
and U4952 (N_4952,N_4354,N_4152);
nor U4953 (N_4953,N_4425,N_4187);
and U4954 (N_4954,N_4197,N_4425);
and U4955 (N_4955,N_4446,N_4385);
nor U4956 (N_4956,N_4085,N_4027);
nand U4957 (N_4957,N_4148,N_4283);
and U4958 (N_4958,N_4092,N_4487);
and U4959 (N_4959,N_4418,N_4106);
nand U4960 (N_4960,N_4389,N_4219);
or U4961 (N_4961,N_4037,N_4406);
nand U4962 (N_4962,N_4118,N_4263);
or U4963 (N_4963,N_4444,N_4405);
or U4964 (N_4964,N_4089,N_4294);
nand U4965 (N_4965,N_4361,N_4077);
and U4966 (N_4966,N_4153,N_4407);
nor U4967 (N_4967,N_4192,N_4305);
or U4968 (N_4968,N_4015,N_4038);
or U4969 (N_4969,N_4480,N_4363);
and U4970 (N_4970,N_4191,N_4144);
or U4971 (N_4971,N_4088,N_4184);
or U4972 (N_4972,N_4048,N_4158);
nor U4973 (N_4973,N_4488,N_4300);
or U4974 (N_4974,N_4161,N_4315);
or U4975 (N_4975,N_4298,N_4383);
or U4976 (N_4976,N_4404,N_4485);
nor U4977 (N_4977,N_4300,N_4060);
nand U4978 (N_4978,N_4048,N_4114);
nand U4979 (N_4979,N_4036,N_4417);
xor U4980 (N_4980,N_4401,N_4007);
nor U4981 (N_4981,N_4269,N_4000);
or U4982 (N_4982,N_4271,N_4437);
and U4983 (N_4983,N_4039,N_4093);
nand U4984 (N_4984,N_4390,N_4026);
nand U4985 (N_4985,N_4466,N_4161);
xnor U4986 (N_4986,N_4212,N_4082);
xor U4987 (N_4987,N_4075,N_4495);
nand U4988 (N_4988,N_4239,N_4497);
or U4989 (N_4989,N_4290,N_4458);
or U4990 (N_4990,N_4219,N_4174);
nand U4991 (N_4991,N_4399,N_4177);
and U4992 (N_4992,N_4263,N_4407);
and U4993 (N_4993,N_4404,N_4397);
or U4994 (N_4994,N_4246,N_4448);
nor U4995 (N_4995,N_4415,N_4448);
or U4996 (N_4996,N_4168,N_4346);
or U4997 (N_4997,N_4312,N_4396);
or U4998 (N_4998,N_4395,N_4064);
or U4999 (N_4999,N_4286,N_4178);
or U5000 (N_5000,N_4898,N_4849);
and U5001 (N_5001,N_4527,N_4672);
and U5002 (N_5002,N_4891,N_4526);
nor U5003 (N_5003,N_4860,N_4575);
nor U5004 (N_5004,N_4576,N_4836);
or U5005 (N_5005,N_4681,N_4518);
xnor U5006 (N_5006,N_4921,N_4905);
nor U5007 (N_5007,N_4769,N_4904);
nor U5008 (N_5008,N_4911,N_4539);
nand U5009 (N_5009,N_4550,N_4816);
and U5010 (N_5010,N_4739,N_4880);
nand U5011 (N_5011,N_4743,N_4704);
nand U5012 (N_5012,N_4830,N_4917);
nor U5013 (N_5013,N_4730,N_4593);
nand U5014 (N_5014,N_4581,N_4888);
and U5015 (N_5015,N_4953,N_4815);
nand U5016 (N_5016,N_4781,N_4696);
and U5017 (N_5017,N_4948,N_4626);
or U5018 (N_5018,N_4560,N_4750);
or U5019 (N_5019,N_4877,N_4597);
nor U5020 (N_5020,N_4813,N_4933);
nor U5021 (N_5021,N_4929,N_4635);
or U5022 (N_5022,N_4683,N_4827);
nor U5023 (N_5023,N_4798,N_4610);
or U5024 (N_5024,N_4852,N_4817);
nor U5025 (N_5025,N_4747,N_4745);
nor U5026 (N_5026,N_4862,N_4649);
and U5027 (N_5027,N_4624,N_4936);
nor U5028 (N_5028,N_4677,N_4780);
and U5029 (N_5029,N_4603,N_4991);
xor U5030 (N_5030,N_4790,N_4759);
nand U5031 (N_5031,N_4967,N_4820);
xnor U5032 (N_5032,N_4809,N_4796);
nor U5033 (N_5033,N_4744,N_4612);
nand U5034 (N_5034,N_4731,N_4679);
nand U5035 (N_5035,N_4647,N_4927);
nand U5036 (N_5036,N_4515,N_4655);
nor U5037 (N_5037,N_4963,N_4653);
xor U5038 (N_5038,N_4695,N_4505);
nor U5039 (N_5039,N_4667,N_4713);
xor U5040 (N_5040,N_4767,N_4588);
or U5041 (N_5041,N_4686,N_4900);
nor U5042 (N_5042,N_4940,N_4664);
and U5043 (N_5043,N_4674,N_4724);
or U5044 (N_5044,N_4645,N_4971);
and U5045 (N_5045,N_4595,N_4574);
nor U5046 (N_5046,N_4670,N_4512);
nor U5047 (N_5047,N_4707,N_4886);
nor U5048 (N_5048,N_4785,N_4972);
nand U5049 (N_5049,N_4719,N_4738);
nand U5050 (N_5050,N_4910,N_4969);
xnor U5051 (N_5051,N_4625,N_4666);
nor U5052 (N_5052,N_4544,N_4985);
nor U5053 (N_5053,N_4962,N_4826);
and U5054 (N_5054,N_4628,N_4659);
or U5055 (N_5055,N_4629,N_4831);
and U5056 (N_5056,N_4878,N_4640);
nor U5057 (N_5057,N_4631,N_4714);
nor U5058 (N_5058,N_4858,N_4841);
nand U5059 (N_5059,N_4792,N_4685);
xor U5060 (N_5060,N_4541,N_4632);
and U5061 (N_5061,N_4840,N_4863);
or U5062 (N_5062,N_4992,N_4954);
or U5063 (N_5063,N_4935,N_4913);
nor U5064 (N_5064,N_4673,N_4501);
and U5065 (N_5065,N_4513,N_4591);
or U5066 (N_5066,N_4979,N_4600);
and U5067 (N_5067,N_4671,N_4521);
and U5068 (N_5068,N_4651,N_4876);
nor U5069 (N_5069,N_4930,N_4545);
or U5070 (N_5070,N_4688,N_4643);
and U5071 (N_5071,N_4509,N_4723);
or U5072 (N_5072,N_4722,N_4834);
or U5073 (N_5073,N_4956,N_4765);
xor U5074 (N_5074,N_4937,N_4735);
nor U5075 (N_5075,N_4500,N_4549);
and U5076 (N_5076,N_4536,N_4627);
nand U5077 (N_5077,N_4596,N_4543);
or U5078 (N_5078,N_4973,N_4517);
or U5079 (N_5079,N_4583,N_4838);
xor U5080 (N_5080,N_4734,N_4968);
xnor U5081 (N_5081,N_4872,N_4994);
nand U5082 (N_5082,N_4571,N_4528);
xnor U5083 (N_5083,N_4693,N_4703);
and U5084 (N_5084,N_4990,N_4751);
or U5085 (N_5085,N_4939,N_4906);
nand U5086 (N_5086,N_4652,N_4959);
nor U5087 (N_5087,N_4709,N_4656);
or U5088 (N_5088,N_4949,N_4561);
and U5089 (N_5089,N_4895,N_4770);
nand U5090 (N_5090,N_4957,N_4533);
nand U5091 (N_5091,N_4601,N_4650);
xor U5092 (N_5092,N_4800,N_4899);
or U5093 (N_5093,N_4995,N_4503);
nand U5094 (N_5094,N_4964,N_4639);
and U5095 (N_5095,N_4675,N_4566);
nand U5096 (N_5096,N_4534,N_4996);
nor U5097 (N_5097,N_4828,N_4502);
or U5098 (N_5098,N_4740,N_4851);
nand U5099 (N_5099,N_4660,N_4865);
and U5100 (N_5100,N_4507,N_4814);
nand U5101 (N_5101,N_4897,N_4975);
nor U5102 (N_5102,N_4636,N_4808);
nand U5103 (N_5103,N_4733,N_4774);
or U5104 (N_5104,N_4641,N_4570);
xor U5105 (N_5105,N_4947,N_4567);
nand U5106 (N_5106,N_4586,N_4926);
and U5107 (N_5107,N_4787,N_4902);
nor U5108 (N_5108,N_4915,N_4942);
and U5109 (N_5109,N_4853,N_4987);
xnor U5110 (N_5110,N_4960,N_4997);
nand U5111 (N_5111,N_4847,N_4710);
and U5112 (N_5112,N_4892,N_4859);
nand U5113 (N_5113,N_4662,N_4896);
nor U5114 (N_5114,N_4978,N_4608);
xor U5115 (N_5115,N_4871,N_4909);
nor U5116 (N_5116,N_4619,N_4606);
nor U5117 (N_5117,N_4661,N_4778);
nor U5118 (N_5118,N_4755,N_4621);
or U5119 (N_5119,N_4557,N_4654);
or U5120 (N_5120,N_4572,N_4614);
xnor U5121 (N_5121,N_4562,N_4889);
nor U5122 (N_5122,N_4870,N_4864);
and U5123 (N_5123,N_4883,N_4764);
or U5124 (N_5124,N_4623,N_4506);
and U5125 (N_5125,N_4775,N_4793);
nor U5126 (N_5126,N_4955,N_4950);
xor U5127 (N_5127,N_4881,N_4689);
xnor U5128 (N_5128,N_4845,N_4810);
and U5129 (N_5129,N_4986,N_4565);
or U5130 (N_5130,N_4715,N_4868);
nand U5131 (N_5131,N_4749,N_4611);
or U5132 (N_5132,N_4680,N_4773);
or U5133 (N_5133,N_4622,N_4832);
and U5134 (N_5134,N_4690,N_4779);
and U5135 (N_5135,N_4806,N_4568);
nand U5136 (N_5136,N_4546,N_4691);
nor U5137 (N_5137,N_4989,N_4726);
nand U5138 (N_5138,N_4676,N_4776);
nor U5139 (N_5139,N_4842,N_4946);
nor U5140 (N_5140,N_4737,N_4717);
or U5141 (N_5141,N_4579,N_4999);
nor U5142 (N_5142,N_4616,N_4928);
nor U5143 (N_5143,N_4604,N_4618);
nand U5144 (N_5144,N_4558,N_4522);
or U5145 (N_5145,N_4736,N_4559);
or U5146 (N_5146,N_4777,N_4794);
nand U5147 (N_5147,N_4584,N_4916);
nor U5148 (N_5148,N_4577,N_4523);
nor U5149 (N_5149,N_4524,N_4762);
xnor U5150 (N_5150,N_4801,N_4598);
nor U5151 (N_5151,N_4843,N_4811);
and U5152 (N_5152,N_4894,N_4564);
nand U5153 (N_5153,N_4923,N_4637);
and U5154 (N_5154,N_4537,N_4783);
or U5155 (N_5155,N_4580,N_4720);
or U5156 (N_5156,N_4525,N_4587);
or U5157 (N_5157,N_4742,N_4799);
xnor U5158 (N_5158,N_4694,N_4547);
or U5159 (N_5159,N_4516,N_4705);
nor U5160 (N_5160,N_4725,N_4687);
and U5161 (N_5161,N_4786,N_4869);
xor U5162 (N_5162,N_4844,N_4941);
or U5163 (N_5163,N_4702,N_4757);
nor U5164 (N_5164,N_4981,N_4839);
nor U5165 (N_5165,N_4829,N_4520);
xnor U5166 (N_5166,N_4998,N_4753);
or U5167 (N_5167,N_4768,N_4741);
nor U5168 (N_5168,N_4804,N_4556);
and U5169 (N_5169,N_4914,N_4663);
nor U5170 (N_5170,N_4805,N_4569);
nand U5171 (N_5171,N_4976,N_4812);
nand U5172 (N_5172,N_4578,N_4712);
or U5173 (N_5173,N_4548,N_4607);
or U5174 (N_5174,N_4553,N_4856);
nand U5175 (N_5175,N_4825,N_4630);
and U5176 (N_5176,N_4620,N_4903);
nor U5177 (N_5177,N_4706,N_4692);
nand U5178 (N_5178,N_4965,N_4818);
or U5179 (N_5179,N_4819,N_4970);
and U5180 (N_5180,N_4701,N_4846);
or U5181 (N_5181,N_4760,N_4634);
nor U5182 (N_5182,N_4728,N_4938);
nor U5183 (N_5183,N_4925,N_4802);
or U5184 (N_5184,N_4824,N_4761);
and U5185 (N_5185,N_4638,N_4882);
or U5186 (N_5186,N_4504,N_4835);
xnor U5187 (N_5187,N_4884,N_4958);
and U5188 (N_5188,N_4589,N_4885);
and U5189 (N_5189,N_4982,N_4658);
and U5190 (N_5190,N_4823,N_4901);
xnor U5191 (N_5191,N_4582,N_4554);
nand U5192 (N_5192,N_4912,N_4922);
xor U5193 (N_5193,N_4711,N_4716);
nand U5194 (N_5194,N_4605,N_4594);
nand U5195 (N_5195,N_4529,N_4531);
xnor U5196 (N_5196,N_4684,N_4754);
nand U5197 (N_5197,N_4931,N_4519);
xor U5198 (N_5198,N_4943,N_4585);
or U5199 (N_5199,N_4893,N_4752);
or U5200 (N_5200,N_4850,N_4945);
nor U5201 (N_5201,N_4668,N_4974);
or U5202 (N_5202,N_4613,N_4807);
or U5203 (N_5203,N_4797,N_4669);
nor U5204 (N_5204,N_4908,N_4857);
and U5205 (N_5205,N_4718,N_4822);
nor U5206 (N_5206,N_4821,N_4646);
nand U5207 (N_5207,N_4538,N_4599);
or U5208 (N_5208,N_4833,N_4602);
xor U5209 (N_5209,N_4866,N_4727);
and U5210 (N_5210,N_4682,N_4551);
xnor U5211 (N_5211,N_4920,N_4803);
or U5212 (N_5212,N_4771,N_4784);
or U5213 (N_5213,N_4848,N_4721);
nor U5214 (N_5214,N_4944,N_4708);
or U5215 (N_5215,N_4746,N_4890);
and U5216 (N_5216,N_4657,N_4988);
nand U5217 (N_5217,N_4615,N_4795);
nor U5218 (N_5218,N_4609,N_4932);
and U5219 (N_5219,N_4980,N_4508);
nor U5220 (N_5220,N_4873,N_4875);
nor U5221 (N_5221,N_4861,N_4563);
nand U5222 (N_5222,N_4642,N_4918);
nand U5223 (N_5223,N_4984,N_4697);
or U5224 (N_5224,N_4919,N_4510);
or U5225 (N_5225,N_4952,N_4552);
xnor U5226 (N_5226,N_4766,N_4837);
nand U5227 (N_5227,N_4732,N_4678);
nor U5228 (N_5228,N_4951,N_4633);
nor U5229 (N_5229,N_4758,N_4874);
or U5230 (N_5230,N_4966,N_4514);
or U5231 (N_5231,N_4700,N_4748);
or U5232 (N_5232,N_4530,N_4772);
or U5233 (N_5233,N_4617,N_4782);
and U5234 (N_5234,N_4854,N_4590);
nand U5235 (N_5235,N_4592,N_4540);
xnor U5236 (N_5236,N_4532,N_4879);
nor U5237 (N_5237,N_4977,N_4644);
and U5238 (N_5238,N_4648,N_4555);
nor U5239 (N_5239,N_4855,N_4573);
or U5240 (N_5240,N_4934,N_4542);
or U5241 (N_5241,N_4788,N_4699);
xor U5242 (N_5242,N_4763,N_4983);
nor U5243 (N_5243,N_4993,N_4907);
nor U5244 (N_5244,N_4924,N_4535);
xnor U5245 (N_5245,N_4756,N_4665);
or U5246 (N_5246,N_4887,N_4867);
and U5247 (N_5247,N_4961,N_4791);
or U5248 (N_5248,N_4511,N_4698);
nand U5249 (N_5249,N_4729,N_4789);
nand U5250 (N_5250,N_4807,N_4811);
and U5251 (N_5251,N_4995,N_4960);
and U5252 (N_5252,N_4653,N_4918);
and U5253 (N_5253,N_4798,N_4700);
or U5254 (N_5254,N_4998,N_4560);
nor U5255 (N_5255,N_4847,N_4697);
nand U5256 (N_5256,N_4946,N_4617);
or U5257 (N_5257,N_4674,N_4939);
nand U5258 (N_5258,N_4748,N_4875);
nand U5259 (N_5259,N_4878,N_4509);
nor U5260 (N_5260,N_4664,N_4703);
and U5261 (N_5261,N_4668,N_4671);
nor U5262 (N_5262,N_4630,N_4856);
nand U5263 (N_5263,N_4749,N_4811);
nor U5264 (N_5264,N_4663,N_4972);
or U5265 (N_5265,N_4816,N_4654);
and U5266 (N_5266,N_4573,N_4500);
or U5267 (N_5267,N_4636,N_4819);
and U5268 (N_5268,N_4983,N_4960);
or U5269 (N_5269,N_4617,N_4979);
or U5270 (N_5270,N_4505,N_4725);
or U5271 (N_5271,N_4749,N_4734);
nand U5272 (N_5272,N_4571,N_4736);
and U5273 (N_5273,N_4679,N_4891);
nor U5274 (N_5274,N_4572,N_4909);
and U5275 (N_5275,N_4593,N_4824);
or U5276 (N_5276,N_4662,N_4874);
or U5277 (N_5277,N_4931,N_4903);
and U5278 (N_5278,N_4943,N_4975);
and U5279 (N_5279,N_4795,N_4882);
xor U5280 (N_5280,N_4937,N_4850);
nand U5281 (N_5281,N_4914,N_4529);
nor U5282 (N_5282,N_4507,N_4892);
and U5283 (N_5283,N_4709,N_4636);
xnor U5284 (N_5284,N_4568,N_4787);
xnor U5285 (N_5285,N_4629,N_4643);
and U5286 (N_5286,N_4773,N_4655);
nand U5287 (N_5287,N_4537,N_4893);
or U5288 (N_5288,N_4744,N_4508);
nand U5289 (N_5289,N_4617,N_4913);
or U5290 (N_5290,N_4616,N_4840);
nand U5291 (N_5291,N_4857,N_4801);
nand U5292 (N_5292,N_4805,N_4593);
nor U5293 (N_5293,N_4690,N_4678);
xnor U5294 (N_5294,N_4642,N_4638);
nand U5295 (N_5295,N_4853,N_4514);
nand U5296 (N_5296,N_4643,N_4832);
and U5297 (N_5297,N_4962,N_4681);
or U5298 (N_5298,N_4520,N_4697);
or U5299 (N_5299,N_4558,N_4981);
nand U5300 (N_5300,N_4692,N_4678);
nor U5301 (N_5301,N_4523,N_4607);
and U5302 (N_5302,N_4656,N_4897);
nand U5303 (N_5303,N_4572,N_4871);
or U5304 (N_5304,N_4896,N_4833);
nand U5305 (N_5305,N_4561,N_4841);
xnor U5306 (N_5306,N_4769,N_4700);
and U5307 (N_5307,N_4901,N_4942);
nand U5308 (N_5308,N_4757,N_4742);
nor U5309 (N_5309,N_4926,N_4538);
nand U5310 (N_5310,N_4769,N_4555);
nand U5311 (N_5311,N_4935,N_4542);
or U5312 (N_5312,N_4550,N_4531);
nand U5313 (N_5313,N_4696,N_4655);
or U5314 (N_5314,N_4542,N_4521);
and U5315 (N_5315,N_4719,N_4635);
nor U5316 (N_5316,N_4935,N_4523);
nand U5317 (N_5317,N_4818,N_4653);
nor U5318 (N_5318,N_4736,N_4743);
nor U5319 (N_5319,N_4938,N_4710);
and U5320 (N_5320,N_4728,N_4780);
nor U5321 (N_5321,N_4542,N_4641);
nand U5322 (N_5322,N_4640,N_4976);
nand U5323 (N_5323,N_4812,N_4629);
xor U5324 (N_5324,N_4876,N_4867);
xnor U5325 (N_5325,N_4606,N_4834);
or U5326 (N_5326,N_4853,N_4540);
xnor U5327 (N_5327,N_4550,N_4640);
xnor U5328 (N_5328,N_4684,N_4828);
nor U5329 (N_5329,N_4604,N_4807);
nand U5330 (N_5330,N_4695,N_4891);
or U5331 (N_5331,N_4920,N_4812);
or U5332 (N_5332,N_4665,N_4975);
or U5333 (N_5333,N_4994,N_4733);
or U5334 (N_5334,N_4664,N_4952);
or U5335 (N_5335,N_4642,N_4954);
xnor U5336 (N_5336,N_4711,N_4954);
and U5337 (N_5337,N_4550,N_4725);
and U5338 (N_5338,N_4638,N_4990);
nor U5339 (N_5339,N_4518,N_4917);
or U5340 (N_5340,N_4550,N_4691);
or U5341 (N_5341,N_4968,N_4632);
nor U5342 (N_5342,N_4711,N_4712);
or U5343 (N_5343,N_4618,N_4749);
and U5344 (N_5344,N_4991,N_4632);
nand U5345 (N_5345,N_4701,N_4836);
nand U5346 (N_5346,N_4696,N_4684);
or U5347 (N_5347,N_4922,N_4744);
nand U5348 (N_5348,N_4999,N_4501);
or U5349 (N_5349,N_4942,N_4515);
and U5350 (N_5350,N_4675,N_4839);
xor U5351 (N_5351,N_4571,N_4962);
or U5352 (N_5352,N_4882,N_4796);
nand U5353 (N_5353,N_4950,N_4824);
or U5354 (N_5354,N_4918,N_4606);
and U5355 (N_5355,N_4692,N_4804);
xnor U5356 (N_5356,N_4964,N_4741);
nor U5357 (N_5357,N_4666,N_4617);
and U5358 (N_5358,N_4865,N_4641);
nor U5359 (N_5359,N_4619,N_4591);
and U5360 (N_5360,N_4722,N_4997);
nor U5361 (N_5361,N_4619,N_4600);
and U5362 (N_5362,N_4521,N_4770);
nand U5363 (N_5363,N_4539,N_4721);
nand U5364 (N_5364,N_4552,N_4629);
and U5365 (N_5365,N_4913,N_4609);
or U5366 (N_5366,N_4927,N_4771);
nand U5367 (N_5367,N_4738,N_4811);
and U5368 (N_5368,N_4673,N_4530);
and U5369 (N_5369,N_4928,N_4791);
and U5370 (N_5370,N_4972,N_4550);
nor U5371 (N_5371,N_4637,N_4953);
nor U5372 (N_5372,N_4915,N_4658);
xnor U5373 (N_5373,N_4957,N_4902);
nor U5374 (N_5374,N_4893,N_4567);
nor U5375 (N_5375,N_4764,N_4817);
nor U5376 (N_5376,N_4829,N_4638);
or U5377 (N_5377,N_4505,N_4796);
nand U5378 (N_5378,N_4916,N_4884);
xnor U5379 (N_5379,N_4613,N_4926);
nor U5380 (N_5380,N_4662,N_4974);
and U5381 (N_5381,N_4875,N_4932);
nor U5382 (N_5382,N_4823,N_4681);
and U5383 (N_5383,N_4758,N_4757);
and U5384 (N_5384,N_4626,N_4731);
nor U5385 (N_5385,N_4585,N_4891);
and U5386 (N_5386,N_4888,N_4574);
or U5387 (N_5387,N_4609,N_4740);
nor U5388 (N_5388,N_4965,N_4540);
or U5389 (N_5389,N_4590,N_4939);
nor U5390 (N_5390,N_4996,N_4845);
or U5391 (N_5391,N_4860,N_4681);
and U5392 (N_5392,N_4601,N_4966);
or U5393 (N_5393,N_4836,N_4624);
nand U5394 (N_5394,N_4565,N_4932);
nor U5395 (N_5395,N_4896,N_4801);
or U5396 (N_5396,N_4790,N_4928);
nor U5397 (N_5397,N_4720,N_4666);
nor U5398 (N_5398,N_4559,N_4552);
and U5399 (N_5399,N_4508,N_4915);
and U5400 (N_5400,N_4905,N_4785);
and U5401 (N_5401,N_4965,N_4648);
nor U5402 (N_5402,N_4883,N_4970);
and U5403 (N_5403,N_4606,N_4536);
and U5404 (N_5404,N_4655,N_4793);
nand U5405 (N_5405,N_4960,N_4700);
nor U5406 (N_5406,N_4900,N_4802);
and U5407 (N_5407,N_4708,N_4554);
nand U5408 (N_5408,N_4526,N_4787);
and U5409 (N_5409,N_4573,N_4632);
or U5410 (N_5410,N_4842,N_4710);
nand U5411 (N_5411,N_4654,N_4838);
nor U5412 (N_5412,N_4800,N_4657);
xnor U5413 (N_5413,N_4905,N_4798);
and U5414 (N_5414,N_4543,N_4848);
or U5415 (N_5415,N_4878,N_4821);
nand U5416 (N_5416,N_4766,N_4993);
or U5417 (N_5417,N_4845,N_4643);
nor U5418 (N_5418,N_4841,N_4892);
and U5419 (N_5419,N_4961,N_4640);
nand U5420 (N_5420,N_4681,N_4840);
and U5421 (N_5421,N_4908,N_4592);
and U5422 (N_5422,N_4935,N_4920);
xnor U5423 (N_5423,N_4912,N_4848);
and U5424 (N_5424,N_4820,N_4790);
xnor U5425 (N_5425,N_4654,N_4675);
and U5426 (N_5426,N_4506,N_4680);
nand U5427 (N_5427,N_4940,N_4953);
xor U5428 (N_5428,N_4828,N_4914);
and U5429 (N_5429,N_4755,N_4503);
nor U5430 (N_5430,N_4917,N_4802);
nand U5431 (N_5431,N_4861,N_4994);
nand U5432 (N_5432,N_4776,N_4522);
nand U5433 (N_5433,N_4982,N_4864);
nand U5434 (N_5434,N_4590,N_4852);
nor U5435 (N_5435,N_4601,N_4979);
nand U5436 (N_5436,N_4973,N_4558);
and U5437 (N_5437,N_4518,N_4679);
and U5438 (N_5438,N_4908,N_4812);
nand U5439 (N_5439,N_4614,N_4656);
nand U5440 (N_5440,N_4887,N_4577);
nand U5441 (N_5441,N_4826,N_4786);
nand U5442 (N_5442,N_4836,N_4644);
xnor U5443 (N_5443,N_4548,N_4870);
nand U5444 (N_5444,N_4794,N_4503);
nor U5445 (N_5445,N_4768,N_4552);
and U5446 (N_5446,N_4929,N_4707);
and U5447 (N_5447,N_4993,N_4876);
and U5448 (N_5448,N_4911,N_4858);
nand U5449 (N_5449,N_4747,N_4893);
xnor U5450 (N_5450,N_4837,N_4650);
and U5451 (N_5451,N_4727,N_4587);
and U5452 (N_5452,N_4691,N_4670);
and U5453 (N_5453,N_4531,N_4673);
or U5454 (N_5454,N_4766,N_4964);
and U5455 (N_5455,N_4952,N_4657);
or U5456 (N_5456,N_4832,N_4770);
and U5457 (N_5457,N_4707,N_4505);
and U5458 (N_5458,N_4514,N_4900);
xnor U5459 (N_5459,N_4968,N_4892);
or U5460 (N_5460,N_4766,N_4882);
nand U5461 (N_5461,N_4849,N_4665);
nand U5462 (N_5462,N_4634,N_4997);
and U5463 (N_5463,N_4569,N_4767);
or U5464 (N_5464,N_4825,N_4579);
nand U5465 (N_5465,N_4541,N_4519);
or U5466 (N_5466,N_4515,N_4907);
nor U5467 (N_5467,N_4736,N_4818);
nand U5468 (N_5468,N_4950,N_4680);
nand U5469 (N_5469,N_4701,N_4505);
or U5470 (N_5470,N_4967,N_4666);
and U5471 (N_5471,N_4967,N_4768);
and U5472 (N_5472,N_4601,N_4852);
nand U5473 (N_5473,N_4811,N_4681);
nor U5474 (N_5474,N_4880,N_4847);
or U5475 (N_5475,N_4687,N_4796);
nor U5476 (N_5476,N_4729,N_4529);
or U5477 (N_5477,N_4922,N_4927);
nor U5478 (N_5478,N_4832,N_4892);
nor U5479 (N_5479,N_4664,N_4620);
nor U5480 (N_5480,N_4570,N_4527);
nor U5481 (N_5481,N_4907,N_4874);
xnor U5482 (N_5482,N_4985,N_4831);
and U5483 (N_5483,N_4611,N_4774);
and U5484 (N_5484,N_4995,N_4679);
nand U5485 (N_5485,N_4540,N_4773);
nor U5486 (N_5486,N_4808,N_4547);
xor U5487 (N_5487,N_4611,N_4526);
nand U5488 (N_5488,N_4808,N_4510);
and U5489 (N_5489,N_4523,N_4691);
and U5490 (N_5490,N_4547,N_4675);
nor U5491 (N_5491,N_4867,N_4850);
or U5492 (N_5492,N_4773,N_4915);
or U5493 (N_5493,N_4837,N_4708);
nor U5494 (N_5494,N_4584,N_4520);
and U5495 (N_5495,N_4754,N_4866);
nor U5496 (N_5496,N_4502,N_4567);
and U5497 (N_5497,N_4601,N_4582);
nor U5498 (N_5498,N_4553,N_4857);
xnor U5499 (N_5499,N_4964,N_4561);
and U5500 (N_5500,N_5449,N_5327);
nor U5501 (N_5501,N_5288,N_5253);
nor U5502 (N_5502,N_5082,N_5363);
nand U5503 (N_5503,N_5463,N_5427);
nand U5504 (N_5504,N_5368,N_5283);
nand U5505 (N_5505,N_5409,N_5186);
or U5506 (N_5506,N_5256,N_5115);
xor U5507 (N_5507,N_5488,N_5418);
nand U5508 (N_5508,N_5485,N_5043);
or U5509 (N_5509,N_5041,N_5497);
xnor U5510 (N_5510,N_5262,N_5429);
nand U5511 (N_5511,N_5328,N_5339);
nor U5512 (N_5512,N_5338,N_5047);
nor U5513 (N_5513,N_5029,N_5104);
nand U5514 (N_5514,N_5393,N_5162);
nand U5515 (N_5515,N_5150,N_5317);
nand U5516 (N_5516,N_5441,N_5438);
nand U5517 (N_5517,N_5039,N_5038);
xor U5518 (N_5518,N_5059,N_5026);
nor U5519 (N_5519,N_5298,N_5171);
and U5520 (N_5520,N_5087,N_5491);
xnor U5521 (N_5521,N_5017,N_5079);
nor U5522 (N_5522,N_5408,N_5224);
or U5523 (N_5523,N_5010,N_5354);
and U5524 (N_5524,N_5030,N_5221);
nand U5525 (N_5525,N_5278,N_5349);
xor U5526 (N_5526,N_5143,N_5398);
nor U5527 (N_5527,N_5451,N_5410);
or U5528 (N_5528,N_5154,N_5309);
nor U5529 (N_5529,N_5064,N_5137);
or U5530 (N_5530,N_5119,N_5467);
xnor U5531 (N_5531,N_5261,N_5267);
or U5532 (N_5532,N_5051,N_5434);
and U5533 (N_5533,N_5108,N_5345);
and U5534 (N_5534,N_5306,N_5003);
nand U5535 (N_5535,N_5037,N_5226);
xor U5536 (N_5536,N_5413,N_5056);
nor U5537 (N_5537,N_5084,N_5357);
nand U5538 (N_5538,N_5300,N_5236);
nand U5539 (N_5539,N_5383,N_5123);
and U5540 (N_5540,N_5350,N_5227);
nor U5541 (N_5541,N_5053,N_5023);
nor U5542 (N_5542,N_5378,N_5360);
nand U5543 (N_5543,N_5273,N_5117);
or U5544 (N_5544,N_5331,N_5476);
and U5545 (N_5545,N_5099,N_5479);
nor U5546 (N_5546,N_5042,N_5089);
and U5547 (N_5547,N_5091,N_5424);
nor U5548 (N_5548,N_5321,N_5381);
and U5549 (N_5549,N_5179,N_5276);
or U5550 (N_5550,N_5055,N_5344);
or U5551 (N_5551,N_5191,N_5075);
nor U5552 (N_5552,N_5456,N_5260);
and U5553 (N_5553,N_5114,N_5021);
nand U5554 (N_5554,N_5196,N_5389);
or U5555 (N_5555,N_5454,N_5135);
or U5556 (N_5556,N_5462,N_5012);
or U5557 (N_5557,N_5478,N_5238);
nor U5558 (N_5558,N_5131,N_5397);
nor U5559 (N_5559,N_5007,N_5359);
nand U5560 (N_5560,N_5483,N_5230);
nor U5561 (N_5561,N_5248,N_5151);
and U5562 (N_5562,N_5365,N_5444);
nand U5563 (N_5563,N_5414,N_5466);
nand U5564 (N_5564,N_5129,N_5384);
nand U5565 (N_5565,N_5379,N_5149);
xor U5566 (N_5566,N_5181,N_5197);
or U5567 (N_5567,N_5493,N_5474);
nand U5568 (N_5568,N_5094,N_5235);
or U5569 (N_5569,N_5140,N_5455);
or U5570 (N_5570,N_5223,N_5044);
nor U5571 (N_5571,N_5161,N_5097);
nor U5572 (N_5572,N_5165,N_5178);
nand U5573 (N_5573,N_5277,N_5022);
nand U5574 (N_5574,N_5296,N_5341);
or U5575 (N_5575,N_5347,N_5486);
or U5576 (N_5576,N_5167,N_5318);
nor U5577 (N_5577,N_5013,N_5305);
xnor U5578 (N_5578,N_5289,N_5286);
or U5579 (N_5579,N_5078,N_5387);
or U5580 (N_5580,N_5473,N_5401);
nor U5581 (N_5581,N_5279,N_5127);
and U5582 (N_5582,N_5433,N_5330);
nor U5583 (N_5583,N_5049,N_5126);
or U5584 (N_5584,N_5291,N_5172);
nand U5585 (N_5585,N_5133,N_5430);
and U5586 (N_5586,N_5332,N_5085);
nand U5587 (N_5587,N_5005,N_5470);
nor U5588 (N_5588,N_5122,N_5292);
and U5589 (N_5589,N_5081,N_5271);
nand U5590 (N_5590,N_5313,N_5245);
nand U5591 (N_5591,N_5353,N_5180);
nor U5592 (N_5592,N_5006,N_5396);
or U5593 (N_5593,N_5045,N_5018);
xnor U5594 (N_5594,N_5281,N_5024);
and U5595 (N_5595,N_5185,N_5184);
nand U5596 (N_5596,N_5304,N_5217);
nor U5597 (N_5597,N_5355,N_5069);
and U5598 (N_5598,N_5132,N_5020);
nand U5599 (N_5599,N_5495,N_5343);
nor U5600 (N_5600,N_5333,N_5169);
and U5601 (N_5601,N_5297,N_5405);
and U5602 (N_5602,N_5210,N_5426);
nor U5603 (N_5603,N_5372,N_5105);
nand U5604 (N_5604,N_5314,N_5376);
and U5605 (N_5605,N_5086,N_5416);
nor U5606 (N_5606,N_5361,N_5116);
nand U5607 (N_5607,N_5062,N_5035);
nor U5608 (N_5608,N_5390,N_5229);
xnor U5609 (N_5609,N_5120,N_5257);
nand U5610 (N_5610,N_5176,N_5275);
nand U5611 (N_5611,N_5205,N_5465);
nor U5612 (N_5612,N_5490,N_5412);
and U5613 (N_5613,N_5420,N_5498);
or U5614 (N_5614,N_5329,N_5046);
nand U5615 (N_5615,N_5083,N_5282);
nor U5616 (N_5616,N_5395,N_5322);
or U5617 (N_5617,N_5336,N_5400);
nor U5618 (N_5618,N_5472,N_5061);
xnor U5619 (N_5619,N_5048,N_5301);
nor U5620 (N_5620,N_5323,N_5373);
nand U5621 (N_5621,N_5188,N_5284);
nand U5622 (N_5622,N_5160,N_5431);
and U5623 (N_5623,N_5411,N_5002);
nand U5624 (N_5624,N_5028,N_5302);
and U5625 (N_5625,N_5362,N_5234);
and U5626 (N_5626,N_5442,N_5219);
and U5627 (N_5627,N_5446,N_5057);
nand U5628 (N_5628,N_5204,N_5246);
nor U5629 (N_5629,N_5208,N_5175);
and U5630 (N_5630,N_5432,N_5098);
or U5631 (N_5631,N_5011,N_5337);
nand U5632 (N_5632,N_5158,N_5088);
or U5633 (N_5633,N_5074,N_5369);
nand U5634 (N_5634,N_5212,N_5453);
and U5635 (N_5635,N_5419,N_5268);
or U5636 (N_5636,N_5443,N_5215);
nand U5637 (N_5637,N_5112,N_5093);
and U5638 (N_5638,N_5287,N_5136);
and U5639 (N_5639,N_5040,N_5452);
xnor U5640 (N_5640,N_5063,N_5377);
xnor U5641 (N_5641,N_5170,N_5388);
and U5642 (N_5642,N_5280,N_5095);
nor U5643 (N_5643,N_5436,N_5475);
and U5644 (N_5644,N_5319,N_5241);
or U5645 (N_5645,N_5071,N_5148);
nand U5646 (N_5646,N_5494,N_5183);
nand U5647 (N_5647,N_5209,N_5073);
or U5648 (N_5648,N_5233,N_5407);
and U5649 (N_5649,N_5134,N_5144);
or U5650 (N_5650,N_5375,N_5076);
or U5651 (N_5651,N_5058,N_5067);
or U5652 (N_5652,N_5484,N_5458);
nor U5653 (N_5653,N_5145,N_5207);
nand U5654 (N_5654,N_5285,N_5404);
and U5655 (N_5655,N_5421,N_5386);
and U5656 (N_5656,N_5100,N_5250);
nand U5657 (N_5657,N_5066,N_5316);
nand U5658 (N_5658,N_5159,N_5324);
and U5659 (N_5659,N_5311,N_5168);
and U5660 (N_5660,N_5008,N_5367);
nand U5661 (N_5661,N_5118,N_5310);
or U5662 (N_5662,N_5106,N_5263);
nand U5663 (N_5663,N_5096,N_5101);
nand U5664 (N_5664,N_5193,N_5054);
nand U5665 (N_5665,N_5403,N_5001);
nor U5666 (N_5666,N_5468,N_5258);
and U5667 (N_5667,N_5239,N_5060);
nor U5668 (N_5668,N_5199,N_5231);
nor U5669 (N_5669,N_5270,N_5157);
xor U5670 (N_5670,N_5004,N_5489);
xor U5671 (N_5671,N_5206,N_5200);
or U5672 (N_5672,N_5218,N_5356);
nand U5673 (N_5673,N_5153,N_5340);
xnor U5674 (N_5674,N_5195,N_5255);
nor U5675 (N_5675,N_5128,N_5351);
nor U5676 (N_5676,N_5482,N_5146);
and U5677 (N_5677,N_5294,N_5342);
or U5678 (N_5678,N_5190,N_5480);
nand U5679 (N_5679,N_5244,N_5050);
and U5680 (N_5680,N_5382,N_5358);
nand U5681 (N_5681,N_5192,N_5033);
and U5682 (N_5682,N_5392,N_5177);
and U5683 (N_5683,N_5174,N_5251);
nand U5684 (N_5684,N_5371,N_5166);
xnor U5685 (N_5685,N_5293,N_5110);
nor U5686 (N_5686,N_5138,N_5471);
or U5687 (N_5687,N_5399,N_5448);
nor U5688 (N_5688,N_5499,N_5141);
xnor U5689 (N_5689,N_5366,N_5307);
or U5690 (N_5690,N_5068,N_5187);
nor U5691 (N_5691,N_5189,N_5266);
and U5692 (N_5692,N_5163,N_5461);
and U5693 (N_5693,N_5065,N_5080);
or U5694 (N_5694,N_5334,N_5460);
nand U5695 (N_5695,N_5222,N_5070);
nand U5696 (N_5696,N_5259,N_5173);
and U5697 (N_5697,N_5036,N_5225);
or U5698 (N_5698,N_5102,N_5370);
xnor U5699 (N_5699,N_5481,N_5147);
nor U5700 (N_5700,N_5031,N_5155);
nor U5701 (N_5701,N_5220,N_5121);
nand U5702 (N_5702,N_5457,N_5380);
nand U5703 (N_5703,N_5016,N_5103);
or U5704 (N_5704,N_5417,N_5269);
nand U5705 (N_5705,N_5213,N_5014);
and U5706 (N_5706,N_5090,N_5464);
and U5707 (N_5707,N_5113,N_5364);
xnor U5708 (N_5708,N_5124,N_5437);
nand U5709 (N_5709,N_5303,N_5032);
xor U5710 (N_5710,N_5402,N_5142);
xnor U5711 (N_5711,N_5320,N_5445);
and U5712 (N_5712,N_5406,N_5077);
and U5713 (N_5713,N_5496,N_5156);
or U5714 (N_5714,N_5312,N_5348);
or U5715 (N_5715,N_5492,N_5295);
or U5716 (N_5716,N_5182,N_5202);
and U5717 (N_5717,N_5092,N_5425);
and U5718 (N_5718,N_5019,N_5237);
or U5719 (N_5719,N_5109,N_5216);
nand U5720 (N_5720,N_5240,N_5346);
and U5721 (N_5721,N_5325,N_5264);
or U5722 (N_5722,N_5247,N_5194);
nor U5723 (N_5723,N_5125,N_5391);
nand U5724 (N_5724,N_5265,N_5447);
nand U5725 (N_5725,N_5450,N_5290);
or U5726 (N_5726,N_5477,N_5394);
nand U5727 (N_5727,N_5428,N_5228);
nor U5728 (N_5728,N_5211,N_5232);
nor U5729 (N_5729,N_5487,N_5459);
and U5730 (N_5730,N_5214,N_5152);
nand U5731 (N_5731,N_5052,N_5326);
and U5732 (N_5732,N_5439,N_5015);
nand U5733 (N_5733,N_5107,N_5072);
nand U5734 (N_5734,N_5164,N_5027);
nor U5735 (N_5735,N_5335,N_5025);
nor U5736 (N_5736,N_5034,N_5440);
or U5737 (N_5737,N_5139,N_5274);
nand U5738 (N_5738,N_5000,N_5203);
or U5739 (N_5739,N_5435,N_5315);
and U5740 (N_5740,N_5469,N_5308);
xor U5741 (N_5741,N_5130,N_5415);
nand U5742 (N_5742,N_5352,N_5254);
nand U5743 (N_5743,N_5423,N_5201);
nand U5744 (N_5744,N_5249,N_5272);
nand U5745 (N_5745,N_5385,N_5009);
or U5746 (N_5746,N_5198,N_5299);
xnor U5747 (N_5747,N_5252,N_5243);
or U5748 (N_5748,N_5242,N_5374);
nor U5749 (N_5749,N_5422,N_5111);
or U5750 (N_5750,N_5048,N_5229);
nor U5751 (N_5751,N_5074,N_5482);
nand U5752 (N_5752,N_5411,N_5093);
nand U5753 (N_5753,N_5025,N_5328);
nand U5754 (N_5754,N_5161,N_5110);
or U5755 (N_5755,N_5139,N_5428);
and U5756 (N_5756,N_5033,N_5315);
and U5757 (N_5757,N_5098,N_5469);
and U5758 (N_5758,N_5390,N_5366);
and U5759 (N_5759,N_5201,N_5238);
or U5760 (N_5760,N_5477,N_5324);
or U5761 (N_5761,N_5180,N_5129);
or U5762 (N_5762,N_5112,N_5206);
and U5763 (N_5763,N_5153,N_5460);
and U5764 (N_5764,N_5434,N_5406);
or U5765 (N_5765,N_5266,N_5190);
and U5766 (N_5766,N_5326,N_5059);
nor U5767 (N_5767,N_5234,N_5286);
or U5768 (N_5768,N_5104,N_5341);
nand U5769 (N_5769,N_5491,N_5281);
and U5770 (N_5770,N_5490,N_5353);
or U5771 (N_5771,N_5222,N_5181);
nor U5772 (N_5772,N_5094,N_5166);
xor U5773 (N_5773,N_5016,N_5477);
nand U5774 (N_5774,N_5275,N_5255);
nand U5775 (N_5775,N_5432,N_5317);
or U5776 (N_5776,N_5218,N_5347);
nor U5777 (N_5777,N_5227,N_5093);
or U5778 (N_5778,N_5001,N_5493);
and U5779 (N_5779,N_5108,N_5416);
xnor U5780 (N_5780,N_5007,N_5246);
nand U5781 (N_5781,N_5360,N_5293);
nor U5782 (N_5782,N_5225,N_5367);
nand U5783 (N_5783,N_5184,N_5013);
nor U5784 (N_5784,N_5140,N_5262);
nand U5785 (N_5785,N_5489,N_5076);
nand U5786 (N_5786,N_5089,N_5088);
nor U5787 (N_5787,N_5093,N_5436);
nand U5788 (N_5788,N_5399,N_5026);
or U5789 (N_5789,N_5225,N_5012);
nand U5790 (N_5790,N_5229,N_5345);
nand U5791 (N_5791,N_5342,N_5242);
xnor U5792 (N_5792,N_5130,N_5406);
or U5793 (N_5793,N_5406,N_5186);
or U5794 (N_5794,N_5483,N_5446);
nor U5795 (N_5795,N_5139,N_5410);
nand U5796 (N_5796,N_5273,N_5245);
nand U5797 (N_5797,N_5274,N_5122);
nand U5798 (N_5798,N_5309,N_5057);
or U5799 (N_5799,N_5196,N_5028);
nand U5800 (N_5800,N_5361,N_5422);
nand U5801 (N_5801,N_5451,N_5136);
xor U5802 (N_5802,N_5437,N_5481);
nand U5803 (N_5803,N_5395,N_5161);
or U5804 (N_5804,N_5246,N_5471);
nand U5805 (N_5805,N_5026,N_5467);
nand U5806 (N_5806,N_5304,N_5459);
and U5807 (N_5807,N_5086,N_5169);
nand U5808 (N_5808,N_5423,N_5118);
nand U5809 (N_5809,N_5251,N_5113);
or U5810 (N_5810,N_5123,N_5405);
nand U5811 (N_5811,N_5101,N_5172);
and U5812 (N_5812,N_5244,N_5152);
or U5813 (N_5813,N_5491,N_5137);
or U5814 (N_5814,N_5253,N_5431);
nand U5815 (N_5815,N_5351,N_5089);
nor U5816 (N_5816,N_5211,N_5389);
nand U5817 (N_5817,N_5389,N_5131);
nand U5818 (N_5818,N_5179,N_5447);
nand U5819 (N_5819,N_5333,N_5241);
or U5820 (N_5820,N_5215,N_5437);
nand U5821 (N_5821,N_5323,N_5437);
nand U5822 (N_5822,N_5221,N_5380);
nor U5823 (N_5823,N_5261,N_5288);
or U5824 (N_5824,N_5336,N_5124);
or U5825 (N_5825,N_5245,N_5401);
nor U5826 (N_5826,N_5163,N_5148);
nor U5827 (N_5827,N_5497,N_5300);
nor U5828 (N_5828,N_5260,N_5420);
and U5829 (N_5829,N_5136,N_5184);
or U5830 (N_5830,N_5024,N_5431);
and U5831 (N_5831,N_5370,N_5318);
nor U5832 (N_5832,N_5176,N_5399);
and U5833 (N_5833,N_5498,N_5283);
nor U5834 (N_5834,N_5362,N_5386);
nor U5835 (N_5835,N_5206,N_5082);
nor U5836 (N_5836,N_5485,N_5025);
nor U5837 (N_5837,N_5029,N_5360);
and U5838 (N_5838,N_5212,N_5330);
or U5839 (N_5839,N_5298,N_5388);
or U5840 (N_5840,N_5466,N_5139);
nor U5841 (N_5841,N_5180,N_5363);
nor U5842 (N_5842,N_5111,N_5371);
xor U5843 (N_5843,N_5043,N_5144);
nand U5844 (N_5844,N_5418,N_5046);
and U5845 (N_5845,N_5265,N_5219);
nor U5846 (N_5846,N_5256,N_5095);
nand U5847 (N_5847,N_5295,N_5096);
or U5848 (N_5848,N_5222,N_5355);
nor U5849 (N_5849,N_5185,N_5189);
or U5850 (N_5850,N_5201,N_5040);
nor U5851 (N_5851,N_5023,N_5443);
nand U5852 (N_5852,N_5179,N_5065);
xnor U5853 (N_5853,N_5371,N_5483);
and U5854 (N_5854,N_5215,N_5147);
xnor U5855 (N_5855,N_5175,N_5484);
and U5856 (N_5856,N_5254,N_5248);
or U5857 (N_5857,N_5248,N_5204);
xor U5858 (N_5858,N_5230,N_5485);
or U5859 (N_5859,N_5189,N_5073);
nor U5860 (N_5860,N_5118,N_5035);
nor U5861 (N_5861,N_5285,N_5321);
nor U5862 (N_5862,N_5181,N_5398);
and U5863 (N_5863,N_5043,N_5385);
and U5864 (N_5864,N_5370,N_5122);
xnor U5865 (N_5865,N_5281,N_5015);
nand U5866 (N_5866,N_5356,N_5363);
and U5867 (N_5867,N_5062,N_5086);
nor U5868 (N_5868,N_5391,N_5201);
xnor U5869 (N_5869,N_5342,N_5020);
and U5870 (N_5870,N_5139,N_5413);
and U5871 (N_5871,N_5300,N_5443);
or U5872 (N_5872,N_5286,N_5365);
or U5873 (N_5873,N_5443,N_5310);
nor U5874 (N_5874,N_5219,N_5385);
nand U5875 (N_5875,N_5421,N_5246);
or U5876 (N_5876,N_5253,N_5352);
nand U5877 (N_5877,N_5257,N_5219);
nor U5878 (N_5878,N_5488,N_5415);
and U5879 (N_5879,N_5056,N_5175);
or U5880 (N_5880,N_5292,N_5417);
xnor U5881 (N_5881,N_5439,N_5294);
or U5882 (N_5882,N_5444,N_5413);
and U5883 (N_5883,N_5157,N_5215);
or U5884 (N_5884,N_5372,N_5119);
nor U5885 (N_5885,N_5254,N_5133);
or U5886 (N_5886,N_5345,N_5334);
or U5887 (N_5887,N_5329,N_5008);
nor U5888 (N_5888,N_5096,N_5432);
nor U5889 (N_5889,N_5248,N_5108);
or U5890 (N_5890,N_5166,N_5255);
nand U5891 (N_5891,N_5177,N_5445);
xor U5892 (N_5892,N_5092,N_5144);
nand U5893 (N_5893,N_5022,N_5286);
nor U5894 (N_5894,N_5433,N_5238);
or U5895 (N_5895,N_5007,N_5358);
nand U5896 (N_5896,N_5438,N_5217);
nand U5897 (N_5897,N_5109,N_5336);
and U5898 (N_5898,N_5304,N_5257);
nor U5899 (N_5899,N_5212,N_5304);
or U5900 (N_5900,N_5164,N_5403);
or U5901 (N_5901,N_5037,N_5164);
and U5902 (N_5902,N_5099,N_5297);
or U5903 (N_5903,N_5458,N_5364);
nor U5904 (N_5904,N_5050,N_5331);
nand U5905 (N_5905,N_5173,N_5071);
nand U5906 (N_5906,N_5274,N_5223);
xor U5907 (N_5907,N_5025,N_5286);
nand U5908 (N_5908,N_5246,N_5263);
and U5909 (N_5909,N_5338,N_5363);
or U5910 (N_5910,N_5290,N_5124);
or U5911 (N_5911,N_5470,N_5132);
and U5912 (N_5912,N_5445,N_5395);
nand U5913 (N_5913,N_5304,N_5282);
and U5914 (N_5914,N_5386,N_5013);
nand U5915 (N_5915,N_5420,N_5208);
and U5916 (N_5916,N_5082,N_5306);
or U5917 (N_5917,N_5079,N_5409);
or U5918 (N_5918,N_5388,N_5261);
nand U5919 (N_5919,N_5288,N_5221);
nor U5920 (N_5920,N_5002,N_5455);
or U5921 (N_5921,N_5108,N_5278);
and U5922 (N_5922,N_5023,N_5333);
or U5923 (N_5923,N_5288,N_5473);
or U5924 (N_5924,N_5406,N_5322);
nand U5925 (N_5925,N_5340,N_5008);
and U5926 (N_5926,N_5274,N_5421);
and U5927 (N_5927,N_5345,N_5386);
nand U5928 (N_5928,N_5140,N_5399);
or U5929 (N_5929,N_5486,N_5450);
and U5930 (N_5930,N_5329,N_5015);
nand U5931 (N_5931,N_5422,N_5032);
nand U5932 (N_5932,N_5330,N_5488);
and U5933 (N_5933,N_5010,N_5168);
or U5934 (N_5934,N_5175,N_5476);
and U5935 (N_5935,N_5138,N_5163);
and U5936 (N_5936,N_5022,N_5118);
nor U5937 (N_5937,N_5336,N_5063);
and U5938 (N_5938,N_5320,N_5178);
or U5939 (N_5939,N_5209,N_5329);
and U5940 (N_5940,N_5434,N_5380);
and U5941 (N_5941,N_5434,N_5011);
or U5942 (N_5942,N_5399,N_5030);
xor U5943 (N_5943,N_5182,N_5048);
nor U5944 (N_5944,N_5239,N_5481);
nor U5945 (N_5945,N_5042,N_5436);
and U5946 (N_5946,N_5032,N_5132);
xnor U5947 (N_5947,N_5295,N_5123);
or U5948 (N_5948,N_5132,N_5130);
xnor U5949 (N_5949,N_5378,N_5457);
nor U5950 (N_5950,N_5154,N_5306);
nand U5951 (N_5951,N_5104,N_5146);
xnor U5952 (N_5952,N_5468,N_5026);
nand U5953 (N_5953,N_5043,N_5241);
nor U5954 (N_5954,N_5424,N_5178);
or U5955 (N_5955,N_5232,N_5052);
nor U5956 (N_5956,N_5024,N_5360);
nor U5957 (N_5957,N_5130,N_5382);
nand U5958 (N_5958,N_5078,N_5259);
nor U5959 (N_5959,N_5116,N_5426);
or U5960 (N_5960,N_5159,N_5078);
and U5961 (N_5961,N_5414,N_5491);
nand U5962 (N_5962,N_5350,N_5224);
or U5963 (N_5963,N_5012,N_5002);
and U5964 (N_5964,N_5234,N_5233);
nand U5965 (N_5965,N_5004,N_5324);
xnor U5966 (N_5966,N_5315,N_5386);
nor U5967 (N_5967,N_5221,N_5066);
and U5968 (N_5968,N_5412,N_5024);
and U5969 (N_5969,N_5394,N_5183);
and U5970 (N_5970,N_5363,N_5207);
or U5971 (N_5971,N_5062,N_5453);
nor U5972 (N_5972,N_5470,N_5301);
and U5973 (N_5973,N_5145,N_5178);
nand U5974 (N_5974,N_5229,N_5211);
nor U5975 (N_5975,N_5165,N_5075);
or U5976 (N_5976,N_5019,N_5010);
nand U5977 (N_5977,N_5122,N_5491);
nand U5978 (N_5978,N_5261,N_5322);
nor U5979 (N_5979,N_5219,N_5238);
nand U5980 (N_5980,N_5267,N_5372);
and U5981 (N_5981,N_5056,N_5346);
and U5982 (N_5982,N_5295,N_5109);
nor U5983 (N_5983,N_5385,N_5348);
and U5984 (N_5984,N_5403,N_5224);
nor U5985 (N_5985,N_5038,N_5268);
and U5986 (N_5986,N_5355,N_5231);
nand U5987 (N_5987,N_5461,N_5030);
nor U5988 (N_5988,N_5333,N_5173);
or U5989 (N_5989,N_5493,N_5448);
and U5990 (N_5990,N_5190,N_5364);
or U5991 (N_5991,N_5132,N_5363);
and U5992 (N_5992,N_5087,N_5128);
or U5993 (N_5993,N_5033,N_5313);
or U5994 (N_5994,N_5416,N_5018);
xnor U5995 (N_5995,N_5068,N_5017);
xnor U5996 (N_5996,N_5191,N_5026);
nand U5997 (N_5997,N_5331,N_5313);
or U5998 (N_5998,N_5480,N_5123);
xnor U5999 (N_5999,N_5364,N_5283);
and U6000 (N_6000,N_5766,N_5657);
nand U6001 (N_6001,N_5851,N_5823);
nor U6002 (N_6002,N_5763,N_5857);
nand U6003 (N_6003,N_5606,N_5953);
and U6004 (N_6004,N_5966,N_5647);
or U6005 (N_6005,N_5644,N_5888);
nand U6006 (N_6006,N_5554,N_5856);
xor U6007 (N_6007,N_5912,N_5829);
or U6008 (N_6008,N_5863,N_5787);
and U6009 (N_6009,N_5867,N_5854);
xnor U6010 (N_6010,N_5963,N_5738);
xor U6011 (N_6011,N_5747,N_5646);
or U6012 (N_6012,N_5926,N_5513);
nand U6013 (N_6013,N_5550,N_5741);
or U6014 (N_6014,N_5777,N_5874);
or U6015 (N_6015,N_5698,N_5725);
or U6016 (N_6016,N_5835,N_5693);
nand U6017 (N_6017,N_5502,N_5555);
nor U6018 (N_6018,N_5560,N_5806);
nor U6019 (N_6019,N_5969,N_5997);
nand U6020 (N_6020,N_5993,N_5954);
nand U6021 (N_6021,N_5733,N_5946);
nand U6022 (N_6022,N_5506,N_5553);
or U6023 (N_6023,N_5855,N_5539);
and U6024 (N_6024,N_5753,N_5962);
or U6025 (N_6025,N_5967,N_5790);
xnor U6026 (N_6026,N_5751,N_5933);
xor U6027 (N_6027,N_5818,N_5822);
nand U6028 (N_6028,N_5648,N_5841);
nor U6029 (N_6029,N_5930,N_5533);
nor U6030 (N_6030,N_5569,N_5571);
and U6031 (N_6031,N_5624,N_5690);
nand U6032 (N_6032,N_5729,N_5797);
and U6033 (N_6033,N_5783,N_5759);
nand U6034 (N_6034,N_5634,N_5552);
xnor U6035 (N_6035,N_5592,N_5789);
nand U6036 (N_6036,N_5580,N_5680);
nor U6037 (N_6037,N_5718,N_5542);
nor U6038 (N_6038,N_5671,N_5934);
or U6039 (N_6039,N_5547,N_5973);
or U6040 (N_6040,N_5957,N_5629);
and U6041 (N_6041,N_5814,N_5697);
or U6042 (N_6042,N_5859,N_5556);
nand U6043 (N_6043,N_5519,N_5794);
or U6044 (N_6044,N_5663,N_5911);
nand U6045 (N_6045,N_5607,N_5650);
and U6046 (N_6046,N_5535,N_5804);
xor U6047 (N_6047,N_5769,N_5514);
xnor U6048 (N_6048,N_5727,N_5767);
nand U6049 (N_6049,N_5645,N_5723);
and U6050 (N_6050,N_5736,N_5931);
and U6051 (N_6051,N_5743,N_5775);
and U6052 (N_6052,N_5627,N_5847);
or U6053 (N_6053,N_5520,N_5941);
nand U6054 (N_6054,N_5879,N_5617);
or U6055 (N_6055,N_5609,N_5722);
and U6056 (N_6056,N_5708,N_5834);
or U6057 (N_6057,N_5896,N_5992);
and U6058 (N_6058,N_5892,N_5816);
or U6059 (N_6059,N_5684,N_5705);
and U6060 (N_6060,N_5530,N_5576);
nand U6061 (N_6061,N_5828,N_5976);
nand U6062 (N_6062,N_5567,N_5824);
and U6063 (N_6063,N_5669,N_5864);
nor U6064 (N_6064,N_5802,N_5516);
and U6065 (N_6065,N_5574,N_5665);
or U6066 (N_6066,N_5603,N_5631);
nand U6067 (N_6067,N_5701,N_5632);
and U6068 (N_6068,N_5950,N_5532);
nor U6069 (N_6069,N_5876,N_5838);
and U6070 (N_6070,N_5799,N_5939);
and U6071 (N_6071,N_5651,N_5803);
nor U6072 (N_6072,N_5654,N_5961);
or U6073 (N_6073,N_5642,N_5712);
nor U6074 (N_6074,N_5836,N_5735);
nor U6075 (N_6075,N_5903,N_5959);
and U6076 (N_6076,N_5662,N_5521);
and U6077 (N_6077,N_5922,N_5906);
and U6078 (N_6078,N_5996,N_5915);
and U6079 (N_6079,N_5508,N_5541);
nand U6080 (N_6080,N_5702,N_5932);
nand U6081 (N_6081,N_5754,N_5745);
and U6082 (N_6082,N_5817,N_5998);
and U6083 (N_6083,N_5726,N_5827);
and U6084 (N_6084,N_5820,N_5910);
and U6085 (N_6085,N_5589,N_5882);
nor U6086 (N_6086,N_5782,N_5604);
nand U6087 (N_6087,N_5614,N_5572);
or U6088 (N_6088,N_5652,N_5507);
or U6089 (N_6089,N_5659,N_5951);
and U6090 (N_6090,N_5699,N_5655);
nand U6091 (N_6091,N_5522,N_5948);
nor U6092 (N_6092,N_5781,N_5732);
xor U6093 (N_6093,N_5594,N_5566);
xor U6094 (N_6094,N_5762,N_5975);
and U6095 (N_6095,N_5917,N_5749);
and U6096 (N_6096,N_5980,N_5528);
and U6097 (N_6097,N_5942,N_5921);
or U6098 (N_6098,N_5501,N_5890);
and U6099 (N_6099,N_5675,N_5633);
nor U6100 (N_6100,N_5798,N_5593);
nor U6101 (N_6101,N_5784,N_5598);
and U6102 (N_6102,N_5866,N_5653);
nand U6103 (N_6103,N_5565,N_5986);
nor U6104 (N_6104,N_5810,N_5907);
xor U6105 (N_6105,N_5955,N_5868);
and U6106 (N_6106,N_5600,N_5979);
and U6107 (N_6107,N_5793,N_5870);
xnor U6108 (N_6108,N_5731,N_5785);
nand U6109 (N_6109,N_5830,N_5720);
and U6110 (N_6110,N_5918,N_5815);
or U6111 (N_6111,N_5691,N_5916);
and U6112 (N_6112,N_5686,N_5536);
nand U6113 (N_6113,N_5586,N_5608);
or U6114 (N_6114,N_5706,N_5551);
xnor U6115 (N_6115,N_5964,N_5666);
nor U6116 (N_6116,N_5658,N_5861);
or U6117 (N_6117,N_5584,N_5801);
or U6118 (N_6118,N_5805,N_5778);
and U6119 (N_6119,N_5623,N_5613);
or U6120 (N_6120,N_5661,N_5581);
nand U6121 (N_6121,N_5618,N_5509);
nand U6122 (N_6122,N_5656,N_5744);
nand U6123 (N_6123,N_5672,N_5602);
and U6124 (N_6124,N_5852,N_5889);
or U6125 (N_6125,N_5517,N_5760);
and U6126 (N_6126,N_5813,N_5515);
and U6127 (N_6127,N_5999,N_5737);
or U6128 (N_6128,N_5643,N_5902);
and U6129 (N_6129,N_5544,N_5640);
or U6130 (N_6130,N_5905,N_5780);
or U6131 (N_6131,N_5591,N_5928);
nand U6132 (N_6132,N_5557,N_5562);
or U6133 (N_6133,N_5582,N_5842);
nand U6134 (N_6134,N_5779,N_5538);
and U6135 (N_6135,N_5843,N_5761);
nand U6136 (N_6136,N_5994,N_5641);
nor U6137 (N_6137,N_5674,N_5636);
and U6138 (N_6138,N_5683,N_5628);
nor U6139 (N_6139,N_5770,N_5893);
nor U6140 (N_6140,N_5837,N_5548);
and U6141 (N_6141,N_5850,N_5710);
nand U6142 (N_6142,N_5925,N_5711);
and U6143 (N_6143,N_5714,N_5730);
and U6144 (N_6144,N_5518,N_5881);
or U6145 (N_6145,N_5908,N_5877);
or U6146 (N_6146,N_5685,N_5742);
nand U6147 (N_6147,N_5715,N_5746);
nand U6148 (N_6148,N_5792,N_5619);
or U6149 (N_6149,N_5833,N_5549);
nand U6150 (N_6150,N_5597,N_5512);
nand U6151 (N_6151,N_5692,N_5800);
nand U6152 (N_6152,N_5831,N_5839);
xnor U6153 (N_6153,N_5970,N_5898);
and U6154 (N_6154,N_5990,N_5897);
nor U6155 (N_6155,N_5811,N_5694);
nor U6156 (N_6156,N_5679,N_5947);
or U6157 (N_6157,N_5878,N_5758);
nand U6158 (N_6158,N_5807,N_5626);
nor U6159 (N_6159,N_5853,N_5958);
and U6160 (N_6160,N_5599,N_5630);
xor U6161 (N_6161,N_5860,N_5531);
and U6162 (N_6162,N_5840,N_5523);
and U6163 (N_6163,N_5622,N_5740);
nor U6164 (N_6164,N_5844,N_5772);
xnor U6165 (N_6165,N_5610,N_5949);
and U6166 (N_6166,N_5717,N_5575);
nor U6167 (N_6167,N_5920,N_5543);
and U6168 (N_6168,N_5500,N_5616);
nand U6169 (N_6169,N_5704,N_5559);
nor U6170 (N_6170,N_5660,N_5995);
nor U6171 (N_6171,N_5703,N_5707);
xnor U6172 (N_6172,N_5936,N_5875);
or U6173 (N_6173,N_5670,N_5972);
or U6174 (N_6174,N_5849,N_5564);
or U6175 (N_6175,N_5873,N_5750);
nor U6176 (N_6176,N_5590,N_5757);
and U6177 (N_6177,N_5637,N_5526);
nor U6178 (N_6178,N_5568,N_5667);
nand U6179 (N_6179,N_5865,N_5681);
and U6180 (N_6180,N_5529,N_5913);
and U6181 (N_6181,N_5595,N_5924);
or U6182 (N_6182,N_5695,N_5688);
xor U6183 (N_6183,N_5558,N_5919);
nand U6184 (N_6184,N_5676,N_5601);
xnor U6185 (N_6185,N_5677,N_5649);
or U6186 (N_6186,N_5596,N_5724);
and U6187 (N_6187,N_5887,N_5687);
or U6188 (N_6188,N_5612,N_5635);
xnor U6189 (N_6189,N_5621,N_5982);
nor U6190 (N_6190,N_5796,N_5579);
nor U6191 (N_6191,N_5987,N_5899);
nor U6192 (N_6192,N_5588,N_5923);
or U6193 (N_6193,N_5668,N_5944);
nand U6194 (N_6194,N_5937,N_5977);
and U6195 (N_6195,N_5578,N_5615);
xnor U6196 (N_6196,N_5795,N_5786);
nand U6197 (N_6197,N_5776,N_5895);
nor U6198 (N_6198,N_5605,N_5678);
nand U6199 (N_6199,N_5886,N_5938);
and U6200 (N_6200,N_5884,N_5524);
xnor U6201 (N_6201,N_5952,N_5985);
nand U6202 (N_6202,N_5620,N_5540);
and U6203 (N_6203,N_5885,N_5577);
or U6204 (N_6204,N_5587,N_5625);
and U6205 (N_6205,N_5988,N_5788);
nor U6206 (N_6206,N_5713,N_5689);
or U6207 (N_6207,N_5974,N_5901);
nand U6208 (N_6208,N_5504,N_5546);
nand U6209 (N_6209,N_5862,N_5956);
or U6210 (N_6210,N_5771,N_5611);
or U6211 (N_6211,N_5819,N_5943);
or U6212 (N_6212,N_5821,N_5752);
and U6213 (N_6213,N_5709,N_5929);
and U6214 (N_6214,N_5585,N_5832);
or U6215 (N_6215,N_5894,N_5505);
or U6216 (N_6216,N_5664,N_5791);
and U6217 (N_6217,N_5700,N_5755);
and U6218 (N_6218,N_5983,N_5638);
xnor U6219 (N_6219,N_5812,N_5858);
and U6220 (N_6220,N_5968,N_5991);
xnor U6221 (N_6221,N_5845,N_5940);
or U6222 (N_6222,N_5965,N_5981);
xnor U6223 (N_6223,N_5503,N_5719);
nand U6224 (N_6224,N_5808,N_5534);
and U6225 (N_6225,N_5971,N_5773);
nand U6226 (N_6226,N_5721,N_5945);
nor U6227 (N_6227,N_5891,N_5511);
or U6228 (N_6228,N_5561,N_5682);
nand U6229 (N_6229,N_5872,N_5871);
or U6230 (N_6230,N_5825,N_5935);
nand U6231 (N_6231,N_5756,N_5728);
nand U6232 (N_6232,N_5563,N_5696);
nor U6233 (N_6233,N_5639,N_5739);
nand U6234 (N_6234,N_5570,N_5989);
nand U6235 (N_6235,N_5583,N_5909);
nor U6236 (N_6236,N_5927,N_5527);
nand U6237 (N_6237,N_5960,N_5525);
or U6238 (N_6238,N_5984,N_5748);
nor U6239 (N_6239,N_5914,N_5848);
and U6240 (N_6240,N_5809,N_5673);
nand U6241 (N_6241,N_5537,N_5768);
nor U6242 (N_6242,N_5869,N_5734);
and U6243 (N_6243,N_5510,N_5900);
nor U6244 (N_6244,N_5774,N_5545);
and U6245 (N_6245,N_5765,N_5573);
nand U6246 (N_6246,N_5883,N_5978);
or U6247 (N_6247,N_5826,N_5764);
and U6248 (N_6248,N_5846,N_5880);
and U6249 (N_6249,N_5716,N_5904);
or U6250 (N_6250,N_5806,N_5815);
nor U6251 (N_6251,N_5959,N_5580);
nor U6252 (N_6252,N_5892,N_5817);
and U6253 (N_6253,N_5668,N_5577);
nand U6254 (N_6254,N_5712,N_5730);
and U6255 (N_6255,N_5652,N_5682);
nand U6256 (N_6256,N_5850,N_5982);
xnor U6257 (N_6257,N_5575,N_5657);
nor U6258 (N_6258,N_5506,N_5850);
or U6259 (N_6259,N_5783,N_5721);
and U6260 (N_6260,N_5881,N_5980);
or U6261 (N_6261,N_5626,N_5507);
nor U6262 (N_6262,N_5615,N_5995);
nand U6263 (N_6263,N_5593,N_5674);
or U6264 (N_6264,N_5688,N_5896);
nor U6265 (N_6265,N_5882,N_5559);
or U6266 (N_6266,N_5583,N_5653);
or U6267 (N_6267,N_5866,N_5710);
nor U6268 (N_6268,N_5582,N_5623);
nand U6269 (N_6269,N_5866,N_5506);
or U6270 (N_6270,N_5610,N_5805);
or U6271 (N_6271,N_5597,N_5867);
nor U6272 (N_6272,N_5603,N_5658);
nor U6273 (N_6273,N_5517,N_5574);
or U6274 (N_6274,N_5631,N_5597);
and U6275 (N_6275,N_5770,N_5737);
and U6276 (N_6276,N_5521,N_5916);
or U6277 (N_6277,N_5835,N_5584);
xnor U6278 (N_6278,N_5793,N_5983);
or U6279 (N_6279,N_5687,N_5637);
nand U6280 (N_6280,N_5888,N_5944);
nor U6281 (N_6281,N_5997,N_5777);
and U6282 (N_6282,N_5581,N_5798);
or U6283 (N_6283,N_5629,N_5756);
nor U6284 (N_6284,N_5736,N_5883);
nand U6285 (N_6285,N_5925,N_5772);
xnor U6286 (N_6286,N_5998,N_5620);
or U6287 (N_6287,N_5807,N_5740);
nor U6288 (N_6288,N_5811,N_5685);
or U6289 (N_6289,N_5621,N_5719);
or U6290 (N_6290,N_5981,N_5601);
or U6291 (N_6291,N_5701,N_5764);
or U6292 (N_6292,N_5914,N_5820);
nand U6293 (N_6293,N_5623,N_5575);
or U6294 (N_6294,N_5775,N_5753);
or U6295 (N_6295,N_5985,N_5596);
nor U6296 (N_6296,N_5849,N_5676);
nor U6297 (N_6297,N_5650,N_5785);
or U6298 (N_6298,N_5574,N_5507);
or U6299 (N_6299,N_5856,N_5839);
nand U6300 (N_6300,N_5991,N_5654);
or U6301 (N_6301,N_5872,N_5624);
and U6302 (N_6302,N_5952,N_5877);
or U6303 (N_6303,N_5807,N_5605);
xor U6304 (N_6304,N_5570,N_5975);
nand U6305 (N_6305,N_5801,N_5971);
nor U6306 (N_6306,N_5876,N_5766);
and U6307 (N_6307,N_5724,N_5675);
nor U6308 (N_6308,N_5684,N_5987);
nand U6309 (N_6309,N_5639,N_5533);
and U6310 (N_6310,N_5654,N_5635);
nor U6311 (N_6311,N_5636,N_5793);
and U6312 (N_6312,N_5656,N_5562);
xor U6313 (N_6313,N_5825,N_5950);
nor U6314 (N_6314,N_5724,N_5593);
nor U6315 (N_6315,N_5778,N_5772);
nor U6316 (N_6316,N_5588,N_5627);
and U6317 (N_6317,N_5690,N_5938);
or U6318 (N_6318,N_5578,N_5754);
or U6319 (N_6319,N_5590,N_5993);
xor U6320 (N_6320,N_5565,N_5836);
and U6321 (N_6321,N_5916,N_5588);
nand U6322 (N_6322,N_5870,N_5611);
nor U6323 (N_6323,N_5649,N_5773);
nand U6324 (N_6324,N_5568,N_5910);
nand U6325 (N_6325,N_5501,N_5656);
or U6326 (N_6326,N_5548,N_5902);
or U6327 (N_6327,N_5508,N_5902);
xnor U6328 (N_6328,N_5526,N_5779);
nand U6329 (N_6329,N_5943,N_5664);
nand U6330 (N_6330,N_5607,N_5633);
and U6331 (N_6331,N_5521,N_5668);
nand U6332 (N_6332,N_5815,N_5764);
or U6333 (N_6333,N_5553,N_5891);
nand U6334 (N_6334,N_5605,N_5660);
xor U6335 (N_6335,N_5664,N_5828);
or U6336 (N_6336,N_5872,N_5614);
and U6337 (N_6337,N_5663,N_5894);
and U6338 (N_6338,N_5731,N_5585);
and U6339 (N_6339,N_5976,N_5662);
xnor U6340 (N_6340,N_5853,N_5987);
and U6341 (N_6341,N_5641,N_5839);
or U6342 (N_6342,N_5598,N_5654);
or U6343 (N_6343,N_5679,N_5827);
or U6344 (N_6344,N_5601,N_5633);
nand U6345 (N_6345,N_5639,N_5717);
xnor U6346 (N_6346,N_5912,N_5782);
or U6347 (N_6347,N_5749,N_5885);
or U6348 (N_6348,N_5704,N_5797);
nor U6349 (N_6349,N_5964,N_5877);
nand U6350 (N_6350,N_5731,N_5988);
xnor U6351 (N_6351,N_5845,N_5604);
nand U6352 (N_6352,N_5935,N_5942);
or U6353 (N_6353,N_5805,N_5620);
nor U6354 (N_6354,N_5677,N_5785);
and U6355 (N_6355,N_5527,N_5696);
or U6356 (N_6356,N_5777,N_5761);
nor U6357 (N_6357,N_5547,N_5582);
nand U6358 (N_6358,N_5755,N_5921);
nor U6359 (N_6359,N_5959,N_5904);
nor U6360 (N_6360,N_5842,N_5919);
and U6361 (N_6361,N_5928,N_5891);
nor U6362 (N_6362,N_5932,N_5535);
nand U6363 (N_6363,N_5765,N_5612);
nor U6364 (N_6364,N_5882,N_5609);
nand U6365 (N_6365,N_5796,N_5972);
nand U6366 (N_6366,N_5880,N_5666);
nand U6367 (N_6367,N_5700,N_5932);
or U6368 (N_6368,N_5727,N_5681);
and U6369 (N_6369,N_5662,N_5938);
nor U6370 (N_6370,N_5939,N_5609);
or U6371 (N_6371,N_5785,N_5937);
xor U6372 (N_6372,N_5750,N_5529);
or U6373 (N_6373,N_5960,N_5722);
or U6374 (N_6374,N_5836,N_5736);
xor U6375 (N_6375,N_5517,N_5912);
xnor U6376 (N_6376,N_5747,N_5517);
xnor U6377 (N_6377,N_5783,N_5972);
xnor U6378 (N_6378,N_5815,N_5645);
nor U6379 (N_6379,N_5682,N_5700);
nand U6380 (N_6380,N_5604,N_5833);
or U6381 (N_6381,N_5794,N_5762);
nand U6382 (N_6382,N_5547,N_5744);
nor U6383 (N_6383,N_5585,N_5729);
nand U6384 (N_6384,N_5690,N_5578);
and U6385 (N_6385,N_5616,N_5944);
and U6386 (N_6386,N_5863,N_5636);
or U6387 (N_6387,N_5716,N_5944);
nand U6388 (N_6388,N_5858,N_5694);
xnor U6389 (N_6389,N_5577,N_5945);
xor U6390 (N_6390,N_5806,N_5573);
xor U6391 (N_6391,N_5561,N_5730);
nor U6392 (N_6392,N_5556,N_5936);
nor U6393 (N_6393,N_5796,N_5886);
and U6394 (N_6394,N_5743,N_5849);
xor U6395 (N_6395,N_5898,N_5508);
or U6396 (N_6396,N_5647,N_5704);
nor U6397 (N_6397,N_5641,N_5579);
nor U6398 (N_6398,N_5971,N_5912);
or U6399 (N_6399,N_5657,N_5530);
nand U6400 (N_6400,N_5730,N_5705);
and U6401 (N_6401,N_5900,N_5583);
nor U6402 (N_6402,N_5823,N_5927);
nand U6403 (N_6403,N_5620,N_5510);
nor U6404 (N_6404,N_5807,N_5738);
nor U6405 (N_6405,N_5536,N_5966);
xnor U6406 (N_6406,N_5568,N_5549);
or U6407 (N_6407,N_5871,N_5570);
nand U6408 (N_6408,N_5780,N_5544);
and U6409 (N_6409,N_5805,N_5842);
xor U6410 (N_6410,N_5718,N_5678);
nor U6411 (N_6411,N_5548,N_5703);
and U6412 (N_6412,N_5519,N_5613);
xor U6413 (N_6413,N_5706,N_5790);
nand U6414 (N_6414,N_5529,N_5916);
nor U6415 (N_6415,N_5840,N_5756);
xnor U6416 (N_6416,N_5631,N_5550);
and U6417 (N_6417,N_5740,N_5726);
nor U6418 (N_6418,N_5706,N_5832);
nor U6419 (N_6419,N_5972,N_5964);
or U6420 (N_6420,N_5690,N_5925);
nand U6421 (N_6421,N_5916,N_5836);
nor U6422 (N_6422,N_5966,N_5824);
nor U6423 (N_6423,N_5935,N_5652);
or U6424 (N_6424,N_5859,N_5689);
and U6425 (N_6425,N_5598,N_5646);
nand U6426 (N_6426,N_5738,N_5626);
or U6427 (N_6427,N_5861,N_5678);
nor U6428 (N_6428,N_5944,N_5853);
nand U6429 (N_6429,N_5759,N_5544);
and U6430 (N_6430,N_5608,N_5966);
or U6431 (N_6431,N_5870,N_5997);
xor U6432 (N_6432,N_5966,N_5642);
nor U6433 (N_6433,N_5820,N_5631);
xor U6434 (N_6434,N_5723,N_5867);
nor U6435 (N_6435,N_5585,N_5713);
nor U6436 (N_6436,N_5688,N_5962);
xnor U6437 (N_6437,N_5544,N_5971);
nor U6438 (N_6438,N_5545,N_5876);
and U6439 (N_6439,N_5884,N_5862);
and U6440 (N_6440,N_5545,N_5760);
xor U6441 (N_6441,N_5501,N_5594);
and U6442 (N_6442,N_5853,N_5833);
nand U6443 (N_6443,N_5887,N_5753);
xor U6444 (N_6444,N_5608,N_5954);
or U6445 (N_6445,N_5664,N_5593);
nand U6446 (N_6446,N_5537,N_5559);
nor U6447 (N_6447,N_5953,N_5864);
nand U6448 (N_6448,N_5582,N_5560);
nand U6449 (N_6449,N_5768,N_5877);
and U6450 (N_6450,N_5653,N_5680);
nand U6451 (N_6451,N_5827,N_5811);
nor U6452 (N_6452,N_5685,N_5763);
and U6453 (N_6453,N_5576,N_5724);
nand U6454 (N_6454,N_5881,N_5825);
nor U6455 (N_6455,N_5766,N_5658);
nand U6456 (N_6456,N_5722,N_5562);
nor U6457 (N_6457,N_5608,N_5884);
nand U6458 (N_6458,N_5615,N_5742);
and U6459 (N_6459,N_5704,N_5593);
and U6460 (N_6460,N_5970,N_5622);
or U6461 (N_6461,N_5569,N_5711);
or U6462 (N_6462,N_5914,N_5936);
and U6463 (N_6463,N_5897,N_5890);
or U6464 (N_6464,N_5511,N_5690);
nand U6465 (N_6465,N_5960,N_5917);
xor U6466 (N_6466,N_5906,N_5828);
nor U6467 (N_6467,N_5648,N_5544);
xor U6468 (N_6468,N_5917,N_5975);
nor U6469 (N_6469,N_5924,N_5538);
nand U6470 (N_6470,N_5859,N_5830);
nand U6471 (N_6471,N_5640,N_5964);
xor U6472 (N_6472,N_5671,N_5854);
and U6473 (N_6473,N_5746,N_5770);
nor U6474 (N_6474,N_5819,N_5931);
nand U6475 (N_6475,N_5906,N_5917);
nor U6476 (N_6476,N_5713,N_5704);
or U6477 (N_6477,N_5856,N_5678);
or U6478 (N_6478,N_5940,N_5945);
or U6479 (N_6479,N_5772,N_5608);
and U6480 (N_6480,N_5981,N_5744);
nand U6481 (N_6481,N_5858,N_5536);
nor U6482 (N_6482,N_5805,N_5907);
and U6483 (N_6483,N_5896,N_5765);
and U6484 (N_6484,N_5632,N_5830);
nand U6485 (N_6485,N_5884,N_5602);
nand U6486 (N_6486,N_5821,N_5601);
or U6487 (N_6487,N_5626,N_5837);
nor U6488 (N_6488,N_5888,N_5735);
nor U6489 (N_6489,N_5948,N_5734);
and U6490 (N_6490,N_5984,N_5568);
or U6491 (N_6491,N_5864,N_5781);
nand U6492 (N_6492,N_5635,N_5681);
or U6493 (N_6493,N_5973,N_5594);
nor U6494 (N_6494,N_5503,N_5634);
and U6495 (N_6495,N_5838,N_5956);
or U6496 (N_6496,N_5605,N_5983);
or U6497 (N_6497,N_5868,N_5909);
nor U6498 (N_6498,N_5653,N_5968);
nor U6499 (N_6499,N_5698,N_5754);
and U6500 (N_6500,N_6248,N_6331);
and U6501 (N_6501,N_6262,N_6082);
or U6502 (N_6502,N_6119,N_6183);
or U6503 (N_6503,N_6268,N_6241);
nand U6504 (N_6504,N_6252,N_6024);
and U6505 (N_6505,N_6058,N_6462);
nor U6506 (N_6506,N_6013,N_6429);
and U6507 (N_6507,N_6489,N_6473);
xnor U6508 (N_6508,N_6387,N_6243);
or U6509 (N_6509,N_6079,N_6449);
nand U6510 (N_6510,N_6091,N_6299);
or U6511 (N_6511,N_6470,N_6061);
nand U6512 (N_6512,N_6386,N_6276);
and U6513 (N_6513,N_6414,N_6355);
nor U6514 (N_6514,N_6270,N_6143);
or U6515 (N_6515,N_6128,N_6096);
and U6516 (N_6516,N_6413,N_6316);
nand U6517 (N_6517,N_6069,N_6221);
or U6518 (N_6518,N_6344,N_6365);
xor U6519 (N_6519,N_6232,N_6236);
nor U6520 (N_6520,N_6379,N_6178);
or U6521 (N_6521,N_6360,N_6432);
nand U6522 (N_6522,N_6324,N_6488);
nand U6523 (N_6523,N_6201,N_6154);
nor U6524 (N_6524,N_6147,N_6076);
nor U6525 (N_6525,N_6300,N_6021);
nor U6526 (N_6526,N_6494,N_6396);
nor U6527 (N_6527,N_6491,N_6454);
and U6528 (N_6528,N_6030,N_6066);
nand U6529 (N_6529,N_6005,N_6308);
or U6530 (N_6530,N_6274,N_6216);
or U6531 (N_6531,N_6409,N_6310);
and U6532 (N_6532,N_6080,N_6466);
nand U6533 (N_6533,N_6017,N_6105);
nor U6534 (N_6534,N_6417,N_6335);
nor U6535 (N_6535,N_6203,N_6407);
nand U6536 (N_6536,N_6109,N_6338);
and U6537 (N_6537,N_6351,N_6347);
or U6538 (N_6538,N_6271,N_6135);
nand U6539 (N_6539,N_6468,N_6229);
nor U6540 (N_6540,N_6411,N_6204);
nand U6541 (N_6541,N_6141,N_6370);
xnor U6542 (N_6542,N_6403,N_6312);
or U6543 (N_6543,N_6043,N_6492);
nand U6544 (N_6544,N_6341,N_6261);
or U6545 (N_6545,N_6198,N_6189);
or U6546 (N_6546,N_6438,N_6071);
and U6547 (N_6547,N_6170,N_6125);
or U6548 (N_6548,N_6213,N_6228);
xor U6549 (N_6549,N_6004,N_6340);
nor U6550 (N_6550,N_6377,N_6426);
or U6551 (N_6551,N_6002,N_6155);
or U6552 (N_6552,N_6456,N_6254);
nand U6553 (N_6553,N_6251,N_6223);
nand U6554 (N_6554,N_6484,N_6244);
nor U6555 (N_6555,N_6081,N_6307);
nor U6556 (N_6556,N_6177,N_6023);
and U6557 (N_6557,N_6418,N_6332);
nor U6558 (N_6558,N_6019,N_6016);
and U6559 (N_6559,N_6317,N_6477);
xnor U6560 (N_6560,N_6471,N_6394);
nor U6561 (N_6561,N_6326,N_6156);
and U6562 (N_6562,N_6346,N_6441);
xnor U6563 (N_6563,N_6085,N_6388);
nand U6564 (N_6564,N_6286,N_6137);
nor U6565 (N_6565,N_6455,N_6068);
or U6566 (N_6566,N_6117,N_6301);
nor U6567 (N_6567,N_6288,N_6138);
and U6568 (N_6568,N_6263,N_6020);
and U6569 (N_6569,N_6089,N_6195);
and U6570 (N_6570,N_6490,N_6062);
and U6571 (N_6571,N_6405,N_6196);
nor U6572 (N_6572,N_6364,N_6412);
or U6573 (N_6573,N_6498,N_6160);
or U6574 (N_6574,N_6187,N_6088);
or U6575 (N_6575,N_6097,N_6011);
nand U6576 (N_6576,N_6210,N_6130);
or U6577 (N_6577,N_6115,N_6336);
nand U6578 (N_6578,N_6486,N_6159);
or U6579 (N_6579,N_6110,N_6293);
xor U6580 (N_6580,N_6014,N_6199);
or U6581 (N_6581,N_6361,N_6450);
xnor U6582 (N_6582,N_6028,N_6285);
or U6583 (N_6583,N_6362,N_6112);
and U6584 (N_6584,N_6144,N_6295);
xor U6585 (N_6585,N_6146,N_6242);
or U6586 (N_6586,N_6026,N_6313);
nor U6587 (N_6587,N_6381,N_6496);
nor U6588 (N_6588,N_6101,N_6006);
nor U6589 (N_6589,N_6174,N_6493);
nand U6590 (N_6590,N_6345,N_6162);
nand U6591 (N_6591,N_6132,N_6458);
nor U6592 (N_6592,N_6027,N_6292);
nor U6593 (N_6593,N_6395,N_6401);
nand U6594 (N_6594,N_6305,N_6298);
and U6595 (N_6595,N_6445,N_6264);
nor U6596 (N_6596,N_6476,N_6083);
xnor U6597 (N_6597,N_6102,N_6060);
nand U6598 (N_6598,N_6397,N_6250);
xor U6599 (N_6599,N_6190,N_6054);
xor U6600 (N_6600,N_6038,N_6368);
or U6601 (N_6601,N_6186,N_6461);
nand U6602 (N_6602,N_6098,N_6367);
xor U6603 (N_6603,N_6009,N_6289);
and U6604 (N_6604,N_6444,N_6194);
nor U6605 (N_6605,N_6419,N_6291);
or U6606 (N_6606,N_6151,N_6166);
and U6607 (N_6607,N_6051,N_6129);
and U6608 (N_6608,N_6318,N_6463);
nand U6609 (N_6609,N_6042,N_6099);
and U6610 (N_6610,N_6281,N_6095);
and U6611 (N_6611,N_6328,N_6440);
nor U6612 (N_6612,N_6480,N_6049);
nor U6613 (N_6613,N_6003,N_6337);
nand U6614 (N_6614,N_6349,N_6245);
nand U6615 (N_6615,N_6055,N_6257);
and U6616 (N_6616,N_6033,N_6075);
and U6617 (N_6617,N_6380,N_6384);
nand U6618 (N_6618,N_6230,N_6279);
and U6619 (N_6619,N_6267,N_6453);
nand U6620 (N_6620,N_6339,N_6392);
nor U6621 (N_6621,N_6459,N_6474);
nand U6622 (N_6622,N_6447,N_6176);
nor U6623 (N_6623,N_6200,N_6217);
nor U6624 (N_6624,N_6278,N_6202);
nand U6625 (N_6625,N_6385,N_6070);
xnor U6626 (N_6626,N_6406,N_6108);
nand U6627 (N_6627,N_6382,N_6207);
and U6628 (N_6628,N_6094,N_6435);
nor U6629 (N_6629,N_6065,N_6327);
nand U6630 (N_6630,N_6104,N_6427);
nor U6631 (N_6631,N_6424,N_6415);
and U6632 (N_6632,N_6495,N_6443);
nor U6633 (N_6633,N_6269,N_6398);
and U6634 (N_6634,N_6272,N_6040);
nor U6635 (N_6635,N_6452,N_6436);
nor U6636 (N_6636,N_6126,N_6249);
or U6637 (N_6637,N_6175,N_6481);
and U6638 (N_6638,N_6334,N_6359);
nand U6639 (N_6639,N_6294,N_6022);
nor U6640 (N_6640,N_6133,N_6180);
or U6641 (N_6641,N_6029,N_6164);
or U6642 (N_6642,N_6234,N_6311);
nand U6643 (N_6643,N_6067,N_6182);
nand U6644 (N_6644,N_6479,N_6322);
or U6645 (N_6645,N_6410,N_6304);
nand U6646 (N_6646,N_6446,N_6191);
nand U6647 (N_6647,N_6265,N_6168);
and U6648 (N_6648,N_6472,N_6373);
nand U6649 (N_6649,N_6158,N_6220);
and U6650 (N_6650,N_6400,N_6193);
or U6651 (N_6651,N_6163,N_6148);
nand U6652 (N_6652,N_6136,N_6059);
nand U6653 (N_6653,N_6072,N_6087);
and U6654 (N_6654,N_6134,N_6399);
or U6655 (N_6655,N_6007,N_6127);
nand U6656 (N_6656,N_6323,N_6325);
or U6657 (N_6657,N_6342,N_6343);
xnor U6658 (N_6658,N_6330,N_6448);
nand U6659 (N_6659,N_6483,N_6314);
nand U6660 (N_6660,N_6048,N_6391);
nor U6661 (N_6661,N_6010,N_6092);
or U6662 (N_6662,N_6114,N_6000);
and U6663 (N_6663,N_6100,N_6366);
nor U6664 (N_6664,N_6356,N_6214);
nand U6665 (N_6665,N_6064,N_6173);
or U6666 (N_6666,N_6255,N_6416);
nor U6667 (N_6667,N_6260,N_6063);
nor U6668 (N_6668,N_6482,N_6046);
or U6669 (N_6669,N_6499,N_6320);
nand U6670 (N_6670,N_6259,N_6103);
nor U6671 (N_6671,N_6056,N_6422);
nor U6672 (N_6672,N_6372,N_6425);
and U6673 (N_6673,N_6212,N_6297);
and U6674 (N_6674,N_6116,N_6035);
and U6675 (N_6675,N_6485,N_6077);
nand U6676 (N_6676,N_6451,N_6460);
and U6677 (N_6677,N_6266,N_6122);
xnor U6678 (N_6678,N_6179,N_6393);
xnor U6679 (N_6679,N_6389,N_6222);
and U6680 (N_6680,N_6209,N_6015);
or U6681 (N_6681,N_6284,N_6197);
xnor U6682 (N_6682,N_6124,N_6233);
nor U6683 (N_6683,N_6231,N_6073);
nor U6684 (N_6684,N_6431,N_6041);
xnor U6685 (N_6685,N_6239,N_6090);
nand U6686 (N_6686,N_6383,N_6034);
nand U6687 (N_6687,N_6036,N_6031);
and U6688 (N_6688,N_6277,N_6378);
or U6689 (N_6689,N_6258,N_6434);
nand U6690 (N_6690,N_6302,N_6211);
nand U6691 (N_6691,N_6282,N_6423);
nor U6692 (N_6692,N_6167,N_6206);
or U6693 (N_6693,N_6172,N_6145);
or U6694 (N_6694,N_6188,N_6497);
nand U6695 (N_6695,N_6321,N_6374);
or U6696 (N_6696,N_6001,N_6185);
or U6697 (N_6697,N_6296,N_6247);
and U6698 (N_6698,N_6044,N_6333);
or U6699 (N_6699,N_6475,N_6237);
and U6700 (N_6700,N_6350,N_6037);
xor U6701 (N_6701,N_6139,N_6430);
or U6702 (N_6702,N_6235,N_6121);
nor U6703 (N_6703,N_6487,N_6348);
or U6704 (N_6704,N_6084,N_6181);
nand U6705 (N_6705,N_6329,N_6169);
nand U6706 (N_6706,N_6192,N_6052);
nor U6707 (N_6707,N_6306,N_6142);
nand U6708 (N_6708,N_6153,N_6246);
and U6709 (N_6709,N_6240,N_6149);
or U6710 (N_6710,N_6113,N_6354);
nor U6711 (N_6711,N_6226,N_6157);
nor U6712 (N_6712,N_6273,N_6358);
and U6713 (N_6713,N_6256,N_6224);
nor U6714 (N_6714,N_6283,N_6227);
and U6715 (N_6715,N_6478,N_6106);
nand U6716 (N_6716,N_6253,N_6018);
nor U6717 (N_6717,N_6439,N_6467);
and U6718 (N_6718,N_6012,N_6215);
or U6719 (N_6719,N_6111,N_6408);
or U6720 (N_6720,N_6165,N_6402);
nand U6721 (N_6721,N_6218,N_6421);
nand U6722 (N_6722,N_6238,N_6219);
xnor U6723 (N_6723,N_6376,N_6074);
or U6724 (N_6724,N_6131,N_6371);
nand U6725 (N_6725,N_6008,N_6047);
nand U6726 (N_6726,N_6039,N_6363);
nor U6727 (N_6727,N_6465,N_6053);
xnor U6728 (N_6728,N_6032,N_6225);
nand U6729 (N_6729,N_6280,N_6442);
nor U6730 (N_6730,N_6152,N_6078);
nand U6731 (N_6731,N_6287,N_6057);
xnor U6732 (N_6732,N_6093,N_6390);
nor U6733 (N_6733,N_6433,N_6025);
nand U6734 (N_6734,N_6290,N_6161);
nor U6735 (N_6735,N_6428,N_6357);
nor U6736 (N_6736,N_6086,N_6469);
or U6737 (N_6737,N_6420,N_6319);
and U6738 (N_6738,N_6150,N_6184);
or U6739 (N_6739,N_6107,N_6315);
xor U6740 (N_6740,N_6140,N_6123);
nor U6741 (N_6741,N_6208,N_6404);
nor U6742 (N_6742,N_6437,N_6352);
or U6743 (N_6743,N_6050,N_6171);
nor U6744 (N_6744,N_6375,N_6275);
or U6745 (N_6745,N_6457,N_6464);
nor U6746 (N_6746,N_6205,N_6303);
nor U6747 (N_6747,N_6045,N_6369);
nand U6748 (N_6748,N_6353,N_6120);
xnor U6749 (N_6749,N_6309,N_6118);
nand U6750 (N_6750,N_6290,N_6005);
and U6751 (N_6751,N_6461,N_6381);
nor U6752 (N_6752,N_6121,N_6103);
xnor U6753 (N_6753,N_6272,N_6473);
and U6754 (N_6754,N_6226,N_6463);
nand U6755 (N_6755,N_6476,N_6312);
nand U6756 (N_6756,N_6417,N_6082);
nand U6757 (N_6757,N_6380,N_6326);
and U6758 (N_6758,N_6421,N_6364);
xnor U6759 (N_6759,N_6495,N_6217);
nor U6760 (N_6760,N_6296,N_6415);
nor U6761 (N_6761,N_6048,N_6012);
nor U6762 (N_6762,N_6454,N_6282);
nand U6763 (N_6763,N_6475,N_6176);
and U6764 (N_6764,N_6488,N_6298);
nor U6765 (N_6765,N_6186,N_6304);
or U6766 (N_6766,N_6485,N_6011);
nor U6767 (N_6767,N_6215,N_6015);
and U6768 (N_6768,N_6492,N_6112);
and U6769 (N_6769,N_6435,N_6019);
nand U6770 (N_6770,N_6144,N_6401);
nand U6771 (N_6771,N_6047,N_6312);
and U6772 (N_6772,N_6482,N_6122);
or U6773 (N_6773,N_6052,N_6200);
or U6774 (N_6774,N_6388,N_6358);
nor U6775 (N_6775,N_6310,N_6014);
or U6776 (N_6776,N_6140,N_6188);
and U6777 (N_6777,N_6339,N_6428);
or U6778 (N_6778,N_6354,N_6282);
nand U6779 (N_6779,N_6030,N_6395);
or U6780 (N_6780,N_6144,N_6179);
nor U6781 (N_6781,N_6180,N_6277);
nor U6782 (N_6782,N_6365,N_6394);
xor U6783 (N_6783,N_6417,N_6371);
or U6784 (N_6784,N_6419,N_6131);
or U6785 (N_6785,N_6365,N_6156);
nand U6786 (N_6786,N_6094,N_6160);
or U6787 (N_6787,N_6166,N_6318);
or U6788 (N_6788,N_6033,N_6176);
and U6789 (N_6789,N_6279,N_6123);
nand U6790 (N_6790,N_6390,N_6488);
nor U6791 (N_6791,N_6483,N_6060);
nand U6792 (N_6792,N_6161,N_6035);
or U6793 (N_6793,N_6047,N_6076);
or U6794 (N_6794,N_6186,N_6092);
nor U6795 (N_6795,N_6135,N_6221);
xnor U6796 (N_6796,N_6282,N_6205);
xor U6797 (N_6797,N_6293,N_6216);
and U6798 (N_6798,N_6456,N_6377);
and U6799 (N_6799,N_6482,N_6338);
and U6800 (N_6800,N_6052,N_6252);
nor U6801 (N_6801,N_6490,N_6068);
or U6802 (N_6802,N_6379,N_6047);
or U6803 (N_6803,N_6137,N_6242);
nor U6804 (N_6804,N_6439,N_6360);
and U6805 (N_6805,N_6155,N_6218);
xnor U6806 (N_6806,N_6143,N_6273);
nand U6807 (N_6807,N_6246,N_6395);
nand U6808 (N_6808,N_6399,N_6033);
and U6809 (N_6809,N_6272,N_6400);
or U6810 (N_6810,N_6462,N_6033);
or U6811 (N_6811,N_6326,N_6158);
or U6812 (N_6812,N_6150,N_6380);
xor U6813 (N_6813,N_6039,N_6083);
or U6814 (N_6814,N_6499,N_6259);
and U6815 (N_6815,N_6136,N_6074);
or U6816 (N_6816,N_6216,N_6206);
nor U6817 (N_6817,N_6291,N_6047);
and U6818 (N_6818,N_6062,N_6273);
and U6819 (N_6819,N_6185,N_6081);
nand U6820 (N_6820,N_6229,N_6255);
or U6821 (N_6821,N_6239,N_6081);
and U6822 (N_6822,N_6140,N_6127);
nor U6823 (N_6823,N_6458,N_6225);
xor U6824 (N_6824,N_6113,N_6484);
nor U6825 (N_6825,N_6071,N_6120);
or U6826 (N_6826,N_6424,N_6108);
or U6827 (N_6827,N_6375,N_6192);
or U6828 (N_6828,N_6362,N_6325);
nor U6829 (N_6829,N_6481,N_6224);
xnor U6830 (N_6830,N_6091,N_6172);
or U6831 (N_6831,N_6103,N_6190);
and U6832 (N_6832,N_6282,N_6371);
nor U6833 (N_6833,N_6146,N_6286);
nand U6834 (N_6834,N_6398,N_6217);
xnor U6835 (N_6835,N_6335,N_6073);
and U6836 (N_6836,N_6033,N_6104);
nand U6837 (N_6837,N_6022,N_6031);
nor U6838 (N_6838,N_6239,N_6499);
xnor U6839 (N_6839,N_6352,N_6043);
and U6840 (N_6840,N_6168,N_6129);
nor U6841 (N_6841,N_6205,N_6174);
or U6842 (N_6842,N_6124,N_6033);
nor U6843 (N_6843,N_6401,N_6397);
nor U6844 (N_6844,N_6392,N_6084);
nor U6845 (N_6845,N_6344,N_6381);
nand U6846 (N_6846,N_6354,N_6328);
nor U6847 (N_6847,N_6045,N_6020);
nand U6848 (N_6848,N_6373,N_6120);
and U6849 (N_6849,N_6429,N_6196);
nor U6850 (N_6850,N_6364,N_6136);
or U6851 (N_6851,N_6120,N_6445);
nor U6852 (N_6852,N_6424,N_6408);
xor U6853 (N_6853,N_6147,N_6213);
and U6854 (N_6854,N_6046,N_6437);
and U6855 (N_6855,N_6212,N_6466);
nand U6856 (N_6856,N_6431,N_6358);
nor U6857 (N_6857,N_6377,N_6102);
nand U6858 (N_6858,N_6029,N_6329);
nand U6859 (N_6859,N_6168,N_6195);
nor U6860 (N_6860,N_6385,N_6332);
and U6861 (N_6861,N_6418,N_6411);
and U6862 (N_6862,N_6193,N_6342);
or U6863 (N_6863,N_6124,N_6290);
nand U6864 (N_6864,N_6217,N_6223);
xor U6865 (N_6865,N_6202,N_6440);
or U6866 (N_6866,N_6060,N_6410);
nor U6867 (N_6867,N_6348,N_6458);
nor U6868 (N_6868,N_6248,N_6339);
and U6869 (N_6869,N_6201,N_6196);
nor U6870 (N_6870,N_6167,N_6011);
or U6871 (N_6871,N_6063,N_6193);
nand U6872 (N_6872,N_6092,N_6323);
nor U6873 (N_6873,N_6347,N_6383);
nor U6874 (N_6874,N_6375,N_6065);
or U6875 (N_6875,N_6337,N_6429);
nand U6876 (N_6876,N_6365,N_6309);
xnor U6877 (N_6877,N_6081,N_6335);
nand U6878 (N_6878,N_6263,N_6252);
nor U6879 (N_6879,N_6316,N_6160);
and U6880 (N_6880,N_6466,N_6202);
nand U6881 (N_6881,N_6258,N_6053);
and U6882 (N_6882,N_6014,N_6204);
nand U6883 (N_6883,N_6269,N_6362);
and U6884 (N_6884,N_6390,N_6033);
and U6885 (N_6885,N_6405,N_6488);
nor U6886 (N_6886,N_6491,N_6308);
and U6887 (N_6887,N_6123,N_6097);
and U6888 (N_6888,N_6117,N_6362);
or U6889 (N_6889,N_6165,N_6083);
nand U6890 (N_6890,N_6210,N_6477);
nand U6891 (N_6891,N_6397,N_6039);
or U6892 (N_6892,N_6100,N_6194);
and U6893 (N_6893,N_6294,N_6160);
and U6894 (N_6894,N_6479,N_6474);
or U6895 (N_6895,N_6206,N_6296);
nand U6896 (N_6896,N_6063,N_6120);
nand U6897 (N_6897,N_6028,N_6076);
or U6898 (N_6898,N_6052,N_6166);
nand U6899 (N_6899,N_6032,N_6260);
nand U6900 (N_6900,N_6251,N_6118);
or U6901 (N_6901,N_6287,N_6461);
nor U6902 (N_6902,N_6421,N_6412);
nand U6903 (N_6903,N_6424,N_6062);
and U6904 (N_6904,N_6141,N_6001);
and U6905 (N_6905,N_6474,N_6112);
nor U6906 (N_6906,N_6401,N_6350);
xor U6907 (N_6907,N_6168,N_6114);
nand U6908 (N_6908,N_6284,N_6006);
nand U6909 (N_6909,N_6036,N_6407);
or U6910 (N_6910,N_6230,N_6043);
nor U6911 (N_6911,N_6044,N_6010);
nand U6912 (N_6912,N_6082,N_6317);
and U6913 (N_6913,N_6378,N_6242);
or U6914 (N_6914,N_6174,N_6090);
or U6915 (N_6915,N_6275,N_6111);
and U6916 (N_6916,N_6207,N_6295);
xnor U6917 (N_6917,N_6384,N_6263);
and U6918 (N_6918,N_6389,N_6407);
nor U6919 (N_6919,N_6355,N_6117);
and U6920 (N_6920,N_6098,N_6137);
and U6921 (N_6921,N_6484,N_6499);
xor U6922 (N_6922,N_6184,N_6208);
nand U6923 (N_6923,N_6363,N_6284);
nor U6924 (N_6924,N_6344,N_6364);
nand U6925 (N_6925,N_6462,N_6183);
xnor U6926 (N_6926,N_6464,N_6254);
nand U6927 (N_6927,N_6276,N_6009);
nor U6928 (N_6928,N_6380,N_6453);
or U6929 (N_6929,N_6429,N_6179);
nand U6930 (N_6930,N_6025,N_6386);
nand U6931 (N_6931,N_6341,N_6453);
nor U6932 (N_6932,N_6237,N_6060);
nor U6933 (N_6933,N_6078,N_6438);
nor U6934 (N_6934,N_6079,N_6256);
nand U6935 (N_6935,N_6083,N_6188);
nor U6936 (N_6936,N_6178,N_6123);
or U6937 (N_6937,N_6429,N_6188);
nor U6938 (N_6938,N_6167,N_6178);
xnor U6939 (N_6939,N_6380,N_6120);
nor U6940 (N_6940,N_6222,N_6499);
and U6941 (N_6941,N_6275,N_6402);
and U6942 (N_6942,N_6490,N_6240);
nand U6943 (N_6943,N_6244,N_6047);
and U6944 (N_6944,N_6176,N_6206);
nand U6945 (N_6945,N_6186,N_6278);
xor U6946 (N_6946,N_6032,N_6360);
xnor U6947 (N_6947,N_6182,N_6144);
nand U6948 (N_6948,N_6342,N_6496);
and U6949 (N_6949,N_6418,N_6190);
and U6950 (N_6950,N_6268,N_6482);
and U6951 (N_6951,N_6167,N_6448);
nand U6952 (N_6952,N_6333,N_6118);
xnor U6953 (N_6953,N_6172,N_6382);
or U6954 (N_6954,N_6158,N_6190);
nor U6955 (N_6955,N_6162,N_6442);
nand U6956 (N_6956,N_6261,N_6030);
nand U6957 (N_6957,N_6199,N_6422);
or U6958 (N_6958,N_6273,N_6364);
and U6959 (N_6959,N_6368,N_6095);
or U6960 (N_6960,N_6031,N_6135);
and U6961 (N_6961,N_6440,N_6334);
nor U6962 (N_6962,N_6359,N_6466);
and U6963 (N_6963,N_6042,N_6121);
nor U6964 (N_6964,N_6074,N_6054);
nor U6965 (N_6965,N_6098,N_6149);
nand U6966 (N_6966,N_6216,N_6166);
or U6967 (N_6967,N_6324,N_6297);
nor U6968 (N_6968,N_6427,N_6193);
or U6969 (N_6969,N_6230,N_6440);
nand U6970 (N_6970,N_6479,N_6432);
nor U6971 (N_6971,N_6293,N_6158);
nor U6972 (N_6972,N_6234,N_6395);
or U6973 (N_6973,N_6469,N_6379);
or U6974 (N_6974,N_6322,N_6284);
nand U6975 (N_6975,N_6362,N_6206);
xnor U6976 (N_6976,N_6041,N_6420);
xor U6977 (N_6977,N_6039,N_6213);
nand U6978 (N_6978,N_6355,N_6281);
or U6979 (N_6979,N_6395,N_6259);
or U6980 (N_6980,N_6479,N_6102);
or U6981 (N_6981,N_6236,N_6247);
or U6982 (N_6982,N_6188,N_6410);
nand U6983 (N_6983,N_6031,N_6495);
nand U6984 (N_6984,N_6030,N_6262);
nand U6985 (N_6985,N_6337,N_6108);
nand U6986 (N_6986,N_6037,N_6015);
nor U6987 (N_6987,N_6276,N_6297);
or U6988 (N_6988,N_6260,N_6449);
nor U6989 (N_6989,N_6206,N_6018);
nor U6990 (N_6990,N_6004,N_6371);
nor U6991 (N_6991,N_6385,N_6271);
nor U6992 (N_6992,N_6267,N_6065);
xnor U6993 (N_6993,N_6312,N_6235);
and U6994 (N_6994,N_6260,N_6322);
nand U6995 (N_6995,N_6014,N_6052);
and U6996 (N_6996,N_6062,N_6045);
xnor U6997 (N_6997,N_6094,N_6455);
nor U6998 (N_6998,N_6062,N_6257);
nand U6999 (N_6999,N_6042,N_6419);
and U7000 (N_7000,N_6775,N_6741);
nor U7001 (N_7001,N_6765,N_6630);
nor U7002 (N_7002,N_6557,N_6795);
xor U7003 (N_7003,N_6653,N_6929);
nor U7004 (N_7004,N_6908,N_6678);
nor U7005 (N_7005,N_6705,N_6767);
or U7006 (N_7006,N_6545,N_6882);
nor U7007 (N_7007,N_6528,N_6598);
nand U7008 (N_7008,N_6671,N_6638);
nand U7009 (N_7009,N_6854,N_6805);
and U7010 (N_7010,N_6619,N_6660);
and U7011 (N_7011,N_6592,N_6806);
nand U7012 (N_7012,N_6532,N_6951);
or U7013 (N_7013,N_6622,N_6914);
xor U7014 (N_7014,N_6569,N_6746);
nor U7015 (N_7015,N_6916,N_6611);
or U7016 (N_7016,N_6708,N_6563);
nand U7017 (N_7017,N_6949,N_6605);
or U7018 (N_7018,N_6631,N_6885);
or U7019 (N_7019,N_6587,N_6596);
or U7020 (N_7020,N_6924,N_6947);
or U7021 (N_7021,N_6868,N_6506);
and U7022 (N_7022,N_6716,N_6675);
nand U7023 (N_7023,N_6603,N_6910);
nor U7024 (N_7024,N_6559,N_6859);
nor U7025 (N_7025,N_6753,N_6721);
nand U7026 (N_7026,N_6970,N_6504);
xor U7027 (N_7027,N_6588,N_6778);
nor U7028 (N_7028,N_6773,N_6965);
or U7029 (N_7029,N_6831,N_6920);
or U7030 (N_7030,N_6998,N_6870);
and U7031 (N_7031,N_6547,N_6833);
nand U7032 (N_7032,N_6742,N_6688);
nor U7033 (N_7033,N_6768,N_6537);
or U7034 (N_7034,N_6521,N_6689);
or U7035 (N_7035,N_6756,N_6883);
and U7036 (N_7036,N_6729,N_6793);
and U7037 (N_7037,N_6702,N_6894);
nand U7038 (N_7038,N_6683,N_6810);
nand U7039 (N_7039,N_6955,N_6770);
nor U7040 (N_7040,N_6527,N_6735);
xor U7041 (N_7041,N_6944,N_6983);
nand U7042 (N_7042,N_6749,N_6591);
and U7043 (N_7043,N_6509,N_6643);
nor U7044 (N_7044,N_6941,N_6938);
nand U7045 (N_7045,N_6820,N_6516);
nor U7046 (N_7046,N_6813,N_6518);
nor U7047 (N_7047,N_6693,N_6962);
nor U7048 (N_7048,N_6604,N_6792);
and U7049 (N_7049,N_6620,N_6972);
and U7050 (N_7050,N_6862,N_6730);
and U7051 (N_7051,N_6906,N_6990);
xnor U7052 (N_7052,N_6761,N_6915);
or U7053 (N_7053,N_6714,N_6762);
nor U7054 (N_7054,N_6709,N_6732);
and U7055 (N_7055,N_6782,N_6835);
nor U7056 (N_7056,N_6738,N_6572);
or U7057 (N_7057,N_6836,N_6907);
nor U7058 (N_7058,N_6979,N_6994);
or U7059 (N_7059,N_6551,N_6945);
or U7060 (N_7060,N_6874,N_6780);
xnor U7061 (N_7061,N_6856,N_6988);
nor U7062 (N_7062,N_6912,N_6999);
nor U7063 (N_7063,N_6621,N_6565);
xor U7064 (N_7064,N_6535,N_6758);
or U7065 (N_7065,N_6802,N_6961);
nand U7066 (N_7066,N_6623,N_6826);
xnor U7067 (N_7067,N_6501,N_6614);
and U7068 (N_7068,N_6838,N_6566);
and U7069 (N_7069,N_6873,N_6879);
or U7070 (N_7070,N_6893,N_6948);
nor U7071 (N_7071,N_6866,N_6713);
and U7072 (N_7072,N_6562,N_6887);
and U7073 (N_7073,N_6971,N_6851);
or U7074 (N_7074,N_6834,N_6748);
and U7075 (N_7075,N_6724,N_6692);
or U7076 (N_7076,N_6917,N_6684);
and U7077 (N_7077,N_6739,N_6832);
xnor U7078 (N_7078,N_6734,N_6803);
or U7079 (N_7079,N_6892,N_6553);
or U7080 (N_7080,N_6601,N_6695);
nor U7081 (N_7081,N_6909,N_6744);
nand U7082 (N_7082,N_6989,N_6645);
xor U7083 (N_7083,N_6896,N_6554);
or U7084 (N_7084,N_6898,N_6530);
or U7085 (N_7085,N_6777,N_6799);
or U7086 (N_7086,N_6957,N_6552);
and U7087 (N_7087,N_6818,N_6752);
nor U7088 (N_7088,N_6980,N_6590);
xor U7089 (N_7089,N_6911,N_6847);
and U7090 (N_7090,N_6581,N_6943);
xor U7091 (N_7091,N_6626,N_6788);
nor U7092 (N_7092,N_6798,N_6939);
or U7093 (N_7093,N_6697,N_6698);
or U7094 (N_7094,N_6586,N_6804);
nor U7095 (N_7095,N_6934,N_6617);
nor U7096 (N_7096,N_6928,N_6636);
nor U7097 (N_7097,N_6568,N_6993);
xor U7098 (N_7098,N_6825,N_6878);
or U7099 (N_7099,N_6737,N_6772);
nand U7100 (N_7100,N_6567,N_6687);
and U7101 (N_7101,N_6731,N_6754);
nor U7102 (N_7102,N_6649,N_6844);
nor U7103 (N_7103,N_6710,N_6507);
or U7104 (N_7104,N_6968,N_6700);
or U7105 (N_7105,N_6776,N_6919);
or U7106 (N_7106,N_6637,N_6644);
nand U7107 (N_7107,N_6578,N_6529);
nor U7108 (N_7108,N_6715,N_6861);
nand U7109 (N_7109,N_6502,N_6658);
nor U7110 (N_7110,N_6650,N_6582);
nand U7111 (N_7111,N_6659,N_6515);
and U7112 (N_7112,N_6670,N_6869);
or U7113 (N_7113,N_6736,N_6876);
or U7114 (N_7114,N_6639,N_6935);
nand U7115 (N_7115,N_6546,N_6648);
nor U7116 (N_7116,N_6613,N_6727);
nor U7117 (N_7117,N_6807,N_6743);
or U7118 (N_7118,N_6867,N_6995);
or U7119 (N_7119,N_6886,N_6992);
or U7120 (N_7120,N_6664,N_6575);
and U7121 (N_7121,N_6872,N_6550);
or U7122 (N_7122,N_6642,N_6607);
xnor U7123 (N_7123,N_6977,N_6556);
and U7124 (N_7124,N_6895,N_6723);
nand U7125 (N_7125,N_6889,N_6794);
nand U7126 (N_7126,N_6984,N_6774);
nor U7127 (N_7127,N_6791,N_6871);
or U7128 (N_7128,N_6815,N_6503);
or U7129 (N_7129,N_6913,N_6950);
xnor U7130 (N_7130,N_6789,N_6875);
nand U7131 (N_7131,N_6514,N_6769);
and U7132 (N_7132,N_6850,N_6819);
xnor U7133 (N_7133,N_6900,N_6956);
nor U7134 (N_7134,N_6864,N_6986);
and U7135 (N_7135,N_6830,N_6661);
or U7136 (N_7136,N_6858,N_6760);
and U7137 (N_7137,N_6967,N_6654);
xor U7138 (N_7138,N_6814,N_6570);
nor U7139 (N_7139,N_6843,N_6933);
nand U7140 (N_7140,N_6808,N_6848);
or U7141 (N_7141,N_6618,N_6641);
nand U7142 (N_7142,N_6975,N_6978);
xnor U7143 (N_7143,N_6652,N_6722);
nor U7144 (N_7144,N_6707,N_6897);
nor U7145 (N_7145,N_6863,N_6615);
or U7146 (N_7146,N_6931,N_6517);
nand U7147 (N_7147,N_6669,N_6573);
nand U7148 (N_7148,N_6719,N_6599);
and U7149 (N_7149,N_6921,N_6534);
nor U7150 (N_7150,N_6881,N_6936);
nor U7151 (N_7151,N_6519,N_6583);
nor U7152 (N_7152,N_6901,N_6728);
nor U7153 (N_7153,N_6536,N_6712);
nand U7154 (N_7154,N_6531,N_6817);
nor U7155 (N_7155,N_6655,N_6682);
or U7156 (N_7156,N_6662,N_6829);
or U7157 (N_7157,N_6558,N_6960);
or U7158 (N_7158,N_6828,N_6969);
or U7159 (N_7159,N_6884,N_6634);
nand U7160 (N_7160,N_6905,N_6512);
or U7161 (N_7161,N_6747,N_6564);
and U7162 (N_7162,N_6681,N_6902);
nand U7163 (N_7163,N_6677,N_6673);
or U7164 (N_7164,N_6667,N_6629);
nor U7165 (N_7165,N_6942,N_6610);
nor U7166 (N_7166,N_6690,N_6811);
nor U7167 (N_7167,N_6890,N_6781);
nand U7168 (N_7168,N_6840,N_6628);
nand U7169 (N_7169,N_6540,N_6680);
nor U7170 (N_7170,N_6755,N_6751);
and U7171 (N_7171,N_6927,N_6633);
or U7172 (N_7172,N_6510,N_6593);
or U7173 (N_7173,N_6757,N_6842);
nor U7174 (N_7174,N_6699,N_6904);
or U7175 (N_7175,N_6865,N_6696);
xnor U7176 (N_7176,N_6685,N_6926);
or U7177 (N_7177,N_6560,N_6891);
and U7178 (N_7178,N_6668,N_6606);
and U7179 (N_7179,N_6663,N_6824);
nor U7180 (N_7180,N_6500,N_6538);
or U7181 (N_7181,N_6796,N_6525);
nor U7182 (N_7182,N_6541,N_6783);
or U7183 (N_7183,N_6571,N_6849);
nor U7184 (N_7184,N_6585,N_6539);
nand U7185 (N_7185,N_6852,N_6561);
and U7186 (N_7186,N_6646,N_6816);
or U7187 (N_7187,N_6549,N_6635);
xor U7188 (N_7188,N_6766,N_6932);
nand U7189 (N_7189,N_6717,N_6976);
and U7190 (N_7190,N_6676,N_6701);
nand U7191 (N_7191,N_6846,N_6800);
nand U7192 (N_7192,N_6997,N_6764);
or U7193 (N_7193,N_6787,N_6740);
nor U7194 (N_7194,N_6505,N_6959);
xor U7195 (N_7195,N_6544,N_6837);
xnor U7196 (N_7196,N_6612,N_6925);
and U7197 (N_7197,N_6632,N_6520);
and U7198 (N_7198,N_6982,N_6853);
and U7199 (N_7199,N_6855,N_6839);
nor U7200 (N_7200,N_6577,N_6627);
nor U7201 (N_7201,N_6857,N_6579);
or U7202 (N_7202,N_6899,N_6651);
nand U7203 (N_7203,N_6542,N_6877);
nor U7204 (N_7204,N_6745,N_6786);
nor U7205 (N_7205,N_6797,N_6589);
and U7206 (N_7206,N_6822,N_6903);
nand U7207 (N_7207,N_6952,N_6996);
nand U7208 (N_7208,N_6625,N_6548);
and U7209 (N_7209,N_6711,N_6974);
and U7210 (N_7210,N_6657,N_6602);
nand U7211 (N_7211,N_6779,N_6691);
nand U7212 (N_7212,N_6964,N_6523);
nand U7213 (N_7213,N_6946,N_6543);
and U7214 (N_7214,N_6513,N_6597);
nand U7215 (N_7215,N_6812,N_6580);
or U7216 (N_7216,N_6930,N_6785);
nand U7217 (N_7217,N_6860,N_6790);
or U7218 (N_7218,N_6616,N_6726);
and U7219 (N_7219,N_6987,N_6533);
or U7220 (N_7220,N_6720,N_6555);
or U7221 (N_7221,N_6845,N_6595);
and U7222 (N_7222,N_6940,N_6524);
and U7223 (N_7223,N_6574,N_6963);
nand U7224 (N_7224,N_6600,N_6686);
nor U7225 (N_7225,N_6704,N_6718);
and U7226 (N_7226,N_6647,N_6763);
nor U7227 (N_7227,N_6576,N_6594);
or U7228 (N_7228,N_6666,N_6880);
and U7229 (N_7229,N_6665,N_6674);
nand U7230 (N_7230,N_6888,N_6694);
nand U7231 (N_7231,N_6985,N_6733);
or U7232 (N_7232,N_6584,N_6809);
nand U7233 (N_7233,N_6609,N_6522);
nor U7234 (N_7234,N_6953,N_6759);
nor U7235 (N_7235,N_6973,N_6750);
and U7236 (N_7236,N_6966,N_6725);
and U7237 (N_7237,N_6991,N_6624);
nand U7238 (N_7238,N_6937,N_6706);
nand U7239 (N_7239,N_6954,N_6981);
nor U7240 (N_7240,N_6608,N_6511);
nand U7241 (N_7241,N_6703,N_6672);
or U7242 (N_7242,N_6526,N_6656);
and U7243 (N_7243,N_6801,N_6841);
or U7244 (N_7244,N_6918,N_6823);
or U7245 (N_7245,N_6827,N_6821);
nand U7246 (N_7246,N_6771,N_6922);
nor U7247 (N_7247,N_6958,N_6923);
and U7248 (N_7248,N_6640,N_6508);
and U7249 (N_7249,N_6784,N_6679);
nor U7250 (N_7250,N_6831,N_6652);
nor U7251 (N_7251,N_6854,N_6507);
nand U7252 (N_7252,N_6927,N_6596);
nand U7253 (N_7253,N_6980,N_6735);
or U7254 (N_7254,N_6959,N_6643);
nand U7255 (N_7255,N_6818,N_6809);
nand U7256 (N_7256,N_6834,N_6553);
nor U7257 (N_7257,N_6788,N_6840);
and U7258 (N_7258,N_6888,N_6689);
nor U7259 (N_7259,N_6732,N_6506);
or U7260 (N_7260,N_6567,N_6872);
nand U7261 (N_7261,N_6834,N_6937);
and U7262 (N_7262,N_6817,N_6589);
or U7263 (N_7263,N_6943,N_6913);
nor U7264 (N_7264,N_6804,N_6828);
xnor U7265 (N_7265,N_6906,N_6518);
nand U7266 (N_7266,N_6510,N_6830);
nor U7267 (N_7267,N_6705,N_6759);
or U7268 (N_7268,N_6840,N_6645);
nand U7269 (N_7269,N_6746,N_6686);
nor U7270 (N_7270,N_6760,N_6754);
nand U7271 (N_7271,N_6743,N_6869);
nand U7272 (N_7272,N_6943,N_6632);
or U7273 (N_7273,N_6848,N_6707);
nor U7274 (N_7274,N_6710,N_6817);
nand U7275 (N_7275,N_6654,N_6913);
nand U7276 (N_7276,N_6737,N_6633);
or U7277 (N_7277,N_6702,N_6892);
nor U7278 (N_7278,N_6742,N_6713);
nand U7279 (N_7279,N_6896,N_6632);
nand U7280 (N_7280,N_6613,N_6720);
nor U7281 (N_7281,N_6944,N_6609);
or U7282 (N_7282,N_6514,N_6657);
nand U7283 (N_7283,N_6766,N_6658);
or U7284 (N_7284,N_6712,N_6903);
xnor U7285 (N_7285,N_6559,N_6936);
xnor U7286 (N_7286,N_6814,N_6962);
or U7287 (N_7287,N_6603,N_6783);
or U7288 (N_7288,N_6670,N_6777);
or U7289 (N_7289,N_6533,N_6513);
and U7290 (N_7290,N_6621,N_6868);
and U7291 (N_7291,N_6747,N_6825);
and U7292 (N_7292,N_6733,N_6565);
xor U7293 (N_7293,N_6563,N_6970);
or U7294 (N_7294,N_6845,N_6935);
nor U7295 (N_7295,N_6763,N_6820);
and U7296 (N_7296,N_6617,N_6556);
nor U7297 (N_7297,N_6771,N_6935);
and U7298 (N_7298,N_6974,N_6818);
or U7299 (N_7299,N_6865,N_6729);
and U7300 (N_7300,N_6619,N_6760);
nor U7301 (N_7301,N_6681,N_6687);
nand U7302 (N_7302,N_6548,N_6825);
nor U7303 (N_7303,N_6660,N_6969);
or U7304 (N_7304,N_6858,N_6835);
and U7305 (N_7305,N_6544,N_6901);
and U7306 (N_7306,N_6889,N_6901);
nor U7307 (N_7307,N_6799,N_6940);
or U7308 (N_7308,N_6637,N_6760);
nor U7309 (N_7309,N_6963,N_6666);
or U7310 (N_7310,N_6635,N_6619);
nand U7311 (N_7311,N_6728,N_6663);
and U7312 (N_7312,N_6763,N_6719);
and U7313 (N_7313,N_6528,N_6792);
and U7314 (N_7314,N_6586,N_6939);
nand U7315 (N_7315,N_6889,N_6768);
nor U7316 (N_7316,N_6515,N_6865);
nor U7317 (N_7317,N_6744,N_6999);
nand U7318 (N_7318,N_6853,N_6624);
or U7319 (N_7319,N_6677,N_6808);
xnor U7320 (N_7320,N_6979,N_6928);
nor U7321 (N_7321,N_6757,N_6830);
xor U7322 (N_7322,N_6564,N_6808);
and U7323 (N_7323,N_6630,N_6663);
nand U7324 (N_7324,N_6503,N_6552);
and U7325 (N_7325,N_6590,N_6934);
nor U7326 (N_7326,N_6680,N_6649);
nand U7327 (N_7327,N_6560,N_6761);
and U7328 (N_7328,N_6695,N_6524);
and U7329 (N_7329,N_6885,N_6769);
or U7330 (N_7330,N_6990,N_6998);
nand U7331 (N_7331,N_6750,N_6856);
and U7332 (N_7332,N_6508,N_6833);
and U7333 (N_7333,N_6565,N_6682);
nor U7334 (N_7334,N_6707,N_6997);
nor U7335 (N_7335,N_6831,N_6547);
nand U7336 (N_7336,N_6766,N_6812);
nor U7337 (N_7337,N_6839,N_6534);
nand U7338 (N_7338,N_6825,N_6955);
nor U7339 (N_7339,N_6595,N_6919);
or U7340 (N_7340,N_6769,N_6905);
nand U7341 (N_7341,N_6581,N_6802);
xnor U7342 (N_7342,N_6588,N_6911);
and U7343 (N_7343,N_6856,N_6903);
and U7344 (N_7344,N_6757,N_6918);
nand U7345 (N_7345,N_6959,N_6888);
nand U7346 (N_7346,N_6945,N_6626);
and U7347 (N_7347,N_6936,N_6715);
or U7348 (N_7348,N_6754,N_6612);
nand U7349 (N_7349,N_6667,N_6604);
and U7350 (N_7350,N_6776,N_6869);
and U7351 (N_7351,N_6735,N_6516);
nand U7352 (N_7352,N_6688,N_6862);
or U7353 (N_7353,N_6709,N_6591);
nor U7354 (N_7354,N_6574,N_6700);
nor U7355 (N_7355,N_6558,N_6907);
nand U7356 (N_7356,N_6815,N_6683);
nor U7357 (N_7357,N_6916,N_6689);
xor U7358 (N_7358,N_6923,N_6890);
or U7359 (N_7359,N_6528,N_6670);
or U7360 (N_7360,N_6896,N_6598);
nand U7361 (N_7361,N_6651,N_6891);
nand U7362 (N_7362,N_6583,N_6715);
and U7363 (N_7363,N_6935,N_6605);
nand U7364 (N_7364,N_6921,N_6576);
or U7365 (N_7365,N_6704,N_6649);
or U7366 (N_7366,N_6679,N_6692);
and U7367 (N_7367,N_6686,N_6768);
xor U7368 (N_7368,N_6967,N_6690);
nand U7369 (N_7369,N_6577,N_6793);
nand U7370 (N_7370,N_6852,N_6851);
or U7371 (N_7371,N_6572,N_6791);
nand U7372 (N_7372,N_6938,N_6633);
and U7373 (N_7373,N_6962,N_6972);
or U7374 (N_7374,N_6556,N_6638);
or U7375 (N_7375,N_6837,N_6755);
nor U7376 (N_7376,N_6806,N_6631);
nand U7377 (N_7377,N_6745,N_6599);
nor U7378 (N_7378,N_6599,N_6912);
and U7379 (N_7379,N_6779,N_6951);
nand U7380 (N_7380,N_6956,N_6735);
or U7381 (N_7381,N_6994,N_6845);
nand U7382 (N_7382,N_6511,N_6683);
or U7383 (N_7383,N_6602,N_6603);
and U7384 (N_7384,N_6964,N_6979);
nand U7385 (N_7385,N_6728,N_6702);
xnor U7386 (N_7386,N_6761,N_6508);
nor U7387 (N_7387,N_6796,N_6888);
and U7388 (N_7388,N_6539,N_6860);
nor U7389 (N_7389,N_6559,N_6840);
and U7390 (N_7390,N_6827,N_6759);
or U7391 (N_7391,N_6835,N_6678);
nand U7392 (N_7392,N_6825,N_6930);
and U7393 (N_7393,N_6805,N_6552);
nor U7394 (N_7394,N_6633,N_6798);
nand U7395 (N_7395,N_6657,N_6647);
or U7396 (N_7396,N_6676,N_6784);
xnor U7397 (N_7397,N_6953,N_6719);
and U7398 (N_7398,N_6917,N_6560);
nand U7399 (N_7399,N_6824,N_6543);
nor U7400 (N_7400,N_6726,N_6876);
or U7401 (N_7401,N_6510,N_6905);
or U7402 (N_7402,N_6765,N_6885);
or U7403 (N_7403,N_6670,N_6820);
or U7404 (N_7404,N_6858,N_6514);
and U7405 (N_7405,N_6834,N_6730);
nand U7406 (N_7406,N_6639,N_6766);
xor U7407 (N_7407,N_6512,N_6933);
nor U7408 (N_7408,N_6684,N_6979);
or U7409 (N_7409,N_6952,N_6747);
xor U7410 (N_7410,N_6580,N_6839);
xnor U7411 (N_7411,N_6997,N_6795);
and U7412 (N_7412,N_6782,N_6786);
and U7413 (N_7413,N_6833,N_6778);
and U7414 (N_7414,N_6807,N_6672);
nor U7415 (N_7415,N_6854,N_6597);
and U7416 (N_7416,N_6967,N_6733);
and U7417 (N_7417,N_6814,N_6766);
nand U7418 (N_7418,N_6720,N_6911);
and U7419 (N_7419,N_6653,N_6930);
xnor U7420 (N_7420,N_6580,N_6953);
or U7421 (N_7421,N_6868,N_6553);
or U7422 (N_7422,N_6580,N_6594);
or U7423 (N_7423,N_6771,N_6808);
and U7424 (N_7424,N_6901,N_6906);
nand U7425 (N_7425,N_6943,N_6769);
xor U7426 (N_7426,N_6907,N_6505);
and U7427 (N_7427,N_6865,N_6782);
nor U7428 (N_7428,N_6729,N_6838);
nor U7429 (N_7429,N_6951,N_6751);
nand U7430 (N_7430,N_6733,N_6971);
nand U7431 (N_7431,N_6883,N_6801);
or U7432 (N_7432,N_6775,N_6914);
nor U7433 (N_7433,N_6685,N_6623);
nand U7434 (N_7434,N_6785,N_6965);
or U7435 (N_7435,N_6560,N_6768);
or U7436 (N_7436,N_6705,N_6520);
or U7437 (N_7437,N_6504,N_6997);
nor U7438 (N_7438,N_6761,N_6716);
nand U7439 (N_7439,N_6824,N_6596);
nor U7440 (N_7440,N_6623,N_6894);
and U7441 (N_7441,N_6821,N_6662);
or U7442 (N_7442,N_6783,N_6974);
nor U7443 (N_7443,N_6995,N_6523);
or U7444 (N_7444,N_6548,N_6931);
nor U7445 (N_7445,N_6594,N_6613);
nor U7446 (N_7446,N_6592,N_6651);
and U7447 (N_7447,N_6784,N_6666);
or U7448 (N_7448,N_6581,N_6632);
nand U7449 (N_7449,N_6570,N_6600);
nand U7450 (N_7450,N_6653,N_6604);
and U7451 (N_7451,N_6973,N_6556);
nand U7452 (N_7452,N_6906,N_6779);
nor U7453 (N_7453,N_6771,N_6765);
nor U7454 (N_7454,N_6641,N_6610);
and U7455 (N_7455,N_6818,N_6755);
xnor U7456 (N_7456,N_6973,N_6864);
and U7457 (N_7457,N_6955,N_6812);
or U7458 (N_7458,N_6732,N_6653);
or U7459 (N_7459,N_6784,N_6881);
or U7460 (N_7460,N_6536,N_6835);
nand U7461 (N_7461,N_6939,N_6529);
xor U7462 (N_7462,N_6950,N_6918);
nor U7463 (N_7463,N_6980,N_6920);
nand U7464 (N_7464,N_6985,N_6901);
xnor U7465 (N_7465,N_6862,N_6548);
nor U7466 (N_7466,N_6682,N_6553);
nand U7467 (N_7467,N_6809,N_6525);
nand U7468 (N_7468,N_6931,N_6668);
or U7469 (N_7469,N_6945,N_6777);
nor U7470 (N_7470,N_6805,N_6731);
or U7471 (N_7471,N_6982,N_6746);
xor U7472 (N_7472,N_6536,N_6842);
and U7473 (N_7473,N_6604,N_6618);
and U7474 (N_7474,N_6742,N_6962);
nand U7475 (N_7475,N_6675,N_6753);
and U7476 (N_7476,N_6549,N_6615);
nand U7477 (N_7477,N_6748,N_6656);
or U7478 (N_7478,N_6816,N_6897);
nor U7479 (N_7479,N_6528,N_6770);
and U7480 (N_7480,N_6994,N_6824);
or U7481 (N_7481,N_6985,N_6896);
nor U7482 (N_7482,N_6701,N_6757);
xor U7483 (N_7483,N_6630,N_6829);
nand U7484 (N_7484,N_6538,N_6804);
nand U7485 (N_7485,N_6596,N_6509);
and U7486 (N_7486,N_6700,N_6746);
nand U7487 (N_7487,N_6902,N_6791);
and U7488 (N_7488,N_6874,N_6518);
nand U7489 (N_7489,N_6593,N_6687);
xor U7490 (N_7490,N_6609,N_6874);
and U7491 (N_7491,N_6818,N_6647);
nand U7492 (N_7492,N_6733,N_6579);
and U7493 (N_7493,N_6804,N_6925);
nand U7494 (N_7494,N_6654,N_6644);
xor U7495 (N_7495,N_6861,N_6590);
or U7496 (N_7496,N_6541,N_6737);
nor U7497 (N_7497,N_6563,N_6725);
nor U7498 (N_7498,N_6518,N_6731);
nor U7499 (N_7499,N_6742,N_6858);
or U7500 (N_7500,N_7377,N_7423);
and U7501 (N_7501,N_7331,N_7396);
nand U7502 (N_7502,N_7038,N_7058);
nand U7503 (N_7503,N_7360,N_7273);
and U7504 (N_7504,N_7264,N_7265);
or U7505 (N_7505,N_7088,N_7049);
or U7506 (N_7506,N_7458,N_7294);
nor U7507 (N_7507,N_7041,N_7017);
nor U7508 (N_7508,N_7206,N_7400);
nand U7509 (N_7509,N_7418,N_7225);
or U7510 (N_7510,N_7305,N_7483);
and U7511 (N_7511,N_7327,N_7196);
and U7512 (N_7512,N_7412,N_7208);
nand U7513 (N_7513,N_7008,N_7101);
nand U7514 (N_7514,N_7303,N_7301);
xor U7515 (N_7515,N_7089,N_7119);
nor U7516 (N_7516,N_7220,N_7202);
xor U7517 (N_7517,N_7257,N_7253);
or U7518 (N_7518,N_7075,N_7329);
nand U7519 (N_7519,N_7092,N_7241);
and U7520 (N_7520,N_7201,N_7459);
or U7521 (N_7521,N_7326,N_7321);
xnor U7522 (N_7522,N_7441,N_7036);
and U7523 (N_7523,N_7037,N_7317);
xnor U7524 (N_7524,N_7368,N_7192);
xnor U7525 (N_7525,N_7133,N_7182);
nor U7526 (N_7526,N_7123,N_7230);
and U7527 (N_7527,N_7187,N_7299);
or U7528 (N_7528,N_7367,N_7014);
nand U7529 (N_7529,N_7043,N_7354);
xnor U7530 (N_7530,N_7068,N_7486);
nand U7531 (N_7531,N_7315,N_7071);
nor U7532 (N_7532,N_7138,N_7312);
and U7533 (N_7533,N_7078,N_7232);
and U7534 (N_7534,N_7086,N_7353);
or U7535 (N_7535,N_7336,N_7385);
nor U7536 (N_7536,N_7141,N_7332);
nor U7537 (N_7537,N_7032,N_7019);
xnor U7538 (N_7538,N_7384,N_7286);
xor U7539 (N_7539,N_7494,N_7283);
nor U7540 (N_7540,N_7455,N_7203);
and U7541 (N_7541,N_7454,N_7076);
nor U7542 (N_7542,N_7247,N_7373);
or U7543 (N_7543,N_7406,N_7463);
and U7544 (N_7544,N_7467,N_7000);
nand U7545 (N_7545,N_7204,N_7226);
nor U7546 (N_7546,N_7309,N_7491);
or U7547 (N_7547,N_7419,N_7444);
or U7548 (N_7548,N_7006,N_7124);
nor U7549 (N_7549,N_7340,N_7474);
nand U7550 (N_7550,N_7300,N_7167);
nand U7551 (N_7551,N_7288,N_7083);
xnor U7552 (N_7552,N_7482,N_7456);
nor U7553 (N_7553,N_7460,N_7324);
nand U7554 (N_7554,N_7057,N_7344);
or U7555 (N_7555,N_7306,N_7371);
or U7556 (N_7556,N_7284,N_7310);
and U7557 (N_7557,N_7224,N_7087);
nor U7558 (N_7558,N_7343,N_7484);
and U7559 (N_7559,N_7015,N_7157);
nand U7560 (N_7560,N_7448,N_7297);
xnor U7561 (N_7561,N_7012,N_7277);
and U7562 (N_7562,N_7422,N_7304);
or U7563 (N_7563,N_7302,N_7117);
or U7564 (N_7564,N_7378,N_7465);
nand U7565 (N_7565,N_7154,N_7366);
nor U7566 (N_7566,N_7433,N_7073);
and U7567 (N_7567,N_7079,N_7211);
or U7568 (N_7568,N_7109,N_7148);
nand U7569 (N_7569,N_7357,N_7060);
nor U7570 (N_7570,N_7488,N_7369);
nand U7571 (N_7571,N_7260,N_7404);
nor U7572 (N_7572,N_7447,N_7213);
nand U7573 (N_7573,N_7296,N_7023);
or U7574 (N_7574,N_7108,N_7389);
or U7575 (N_7575,N_7116,N_7162);
nor U7576 (N_7576,N_7240,N_7199);
nand U7577 (N_7577,N_7269,N_7335);
and U7578 (N_7578,N_7183,N_7308);
nand U7579 (N_7579,N_7420,N_7325);
and U7580 (N_7580,N_7047,N_7009);
or U7581 (N_7581,N_7387,N_7097);
nand U7582 (N_7582,N_7349,N_7276);
nor U7583 (N_7583,N_7114,N_7067);
nand U7584 (N_7584,N_7016,N_7129);
nor U7585 (N_7585,N_7328,N_7070);
nor U7586 (N_7586,N_7118,N_7480);
and U7587 (N_7587,N_7055,N_7405);
nor U7588 (N_7588,N_7184,N_7190);
nand U7589 (N_7589,N_7359,N_7151);
nand U7590 (N_7590,N_7053,N_7236);
and U7591 (N_7591,N_7051,N_7319);
and U7592 (N_7592,N_7263,N_7440);
nand U7593 (N_7593,N_7379,N_7239);
nor U7594 (N_7594,N_7275,N_7207);
and U7595 (N_7595,N_7391,N_7497);
and U7596 (N_7596,N_7293,N_7125);
xnor U7597 (N_7597,N_7111,N_7080);
and U7598 (N_7598,N_7272,N_7210);
or U7599 (N_7599,N_7330,N_7180);
nor U7600 (N_7600,N_7429,N_7443);
nor U7601 (N_7601,N_7394,N_7155);
or U7602 (N_7602,N_7018,N_7383);
nand U7603 (N_7603,N_7228,N_7091);
and U7604 (N_7604,N_7198,N_7168);
and U7605 (N_7605,N_7289,N_7365);
or U7606 (N_7606,N_7449,N_7066);
nor U7607 (N_7607,N_7375,N_7156);
or U7608 (N_7608,N_7082,N_7231);
or U7609 (N_7609,N_7243,N_7475);
or U7610 (N_7610,N_7255,N_7256);
or U7611 (N_7611,N_7476,N_7414);
and U7612 (N_7612,N_7139,N_7234);
nor U7613 (N_7613,N_7323,N_7030);
nand U7614 (N_7614,N_7040,N_7372);
or U7615 (N_7615,N_7471,N_7258);
nor U7616 (N_7616,N_7376,N_7022);
and U7617 (N_7617,N_7218,N_7472);
nor U7618 (N_7618,N_7110,N_7136);
and U7619 (N_7619,N_7285,N_7397);
nand U7620 (N_7620,N_7492,N_7178);
nor U7621 (N_7621,N_7158,N_7222);
xor U7622 (N_7622,N_7442,N_7451);
nand U7623 (N_7623,N_7238,N_7435);
nor U7624 (N_7624,N_7386,N_7363);
nor U7625 (N_7625,N_7216,N_7341);
nand U7626 (N_7626,N_7411,N_7364);
nand U7627 (N_7627,N_7496,N_7350);
nand U7628 (N_7628,N_7176,N_7085);
and U7629 (N_7629,N_7246,N_7096);
nand U7630 (N_7630,N_7056,N_7398);
nand U7631 (N_7631,N_7069,N_7399);
xnor U7632 (N_7632,N_7267,N_7165);
nor U7633 (N_7633,N_7237,N_7095);
or U7634 (N_7634,N_7464,N_7031);
xor U7635 (N_7635,N_7142,N_7077);
and U7636 (N_7636,N_7307,N_7254);
or U7637 (N_7637,N_7351,N_7197);
nor U7638 (N_7638,N_7421,N_7462);
or U7639 (N_7639,N_7487,N_7259);
nor U7640 (N_7640,N_7113,N_7024);
nor U7641 (N_7641,N_7150,N_7450);
nor U7642 (N_7642,N_7099,N_7282);
nand U7643 (N_7643,N_7356,N_7126);
xor U7644 (N_7644,N_7334,N_7153);
xor U7645 (N_7645,N_7424,N_7159);
or U7646 (N_7646,N_7278,N_7145);
and U7647 (N_7647,N_7170,N_7426);
and U7648 (N_7648,N_7021,N_7205);
or U7649 (N_7649,N_7002,N_7445);
and U7650 (N_7650,N_7065,N_7064);
nor U7651 (N_7651,N_7172,N_7195);
or U7652 (N_7652,N_7026,N_7251);
nor U7653 (N_7653,N_7045,N_7274);
or U7654 (N_7654,N_7481,N_7410);
nand U7655 (N_7655,N_7403,N_7061);
xnor U7656 (N_7656,N_7181,N_7245);
or U7657 (N_7657,N_7427,N_7059);
nand U7658 (N_7658,N_7010,N_7416);
or U7659 (N_7659,N_7291,N_7347);
and U7660 (N_7660,N_7011,N_7250);
nor U7661 (N_7661,N_7219,N_7169);
nand U7662 (N_7662,N_7215,N_7163);
or U7663 (N_7663,N_7362,N_7042);
or U7664 (N_7664,N_7313,N_7348);
or U7665 (N_7665,N_7229,N_7127);
or U7666 (N_7666,N_7437,N_7122);
nor U7667 (N_7667,N_7295,N_7052);
nand U7668 (N_7668,N_7166,N_7374);
and U7669 (N_7669,N_7160,N_7479);
nand U7670 (N_7670,N_7425,N_7177);
or U7671 (N_7671,N_7143,N_7290);
nor U7672 (N_7672,N_7025,N_7007);
xor U7673 (N_7673,N_7185,N_7098);
nand U7674 (N_7674,N_7131,N_7407);
or U7675 (N_7675,N_7271,N_7320);
or U7676 (N_7676,N_7287,N_7013);
or U7677 (N_7677,N_7094,N_7311);
and U7678 (N_7678,N_7495,N_7001);
and U7679 (N_7679,N_7100,N_7415);
nor U7680 (N_7680,N_7469,N_7227);
or U7681 (N_7681,N_7452,N_7355);
nand U7682 (N_7682,N_7402,N_7316);
xor U7683 (N_7683,N_7081,N_7346);
or U7684 (N_7684,N_7453,N_7054);
nor U7685 (N_7685,N_7242,N_7214);
nand U7686 (N_7686,N_7034,N_7408);
or U7687 (N_7687,N_7191,N_7050);
nor U7688 (N_7688,N_7135,N_7490);
and U7689 (N_7689,N_7048,N_7493);
nor U7690 (N_7690,N_7244,N_7161);
and U7691 (N_7691,N_7409,N_7164);
or U7692 (N_7692,N_7438,N_7147);
and U7693 (N_7693,N_7105,N_7028);
nand U7694 (N_7694,N_7189,N_7186);
and U7695 (N_7695,N_7132,N_7345);
nand U7696 (N_7696,N_7428,N_7361);
nand U7697 (N_7697,N_7046,N_7370);
and U7698 (N_7698,N_7430,N_7498);
or U7699 (N_7699,N_7063,N_7130);
nand U7700 (N_7700,N_7298,N_7128);
and U7701 (N_7701,N_7112,N_7221);
nand U7702 (N_7702,N_7318,N_7292);
nor U7703 (N_7703,N_7217,N_7107);
nand U7704 (N_7704,N_7261,N_7106);
nor U7705 (N_7705,N_7212,N_7431);
and U7706 (N_7706,N_7279,N_7235);
or U7707 (N_7707,N_7439,N_7020);
and U7708 (N_7708,N_7248,N_7392);
and U7709 (N_7709,N_7174,N_7200);
nor U7710 (N_7710,N_7266,N_7004);
nor U7711 (N_7711,N_7268,N_7035);
nor U7712 (N_7712,N_7314,N_7352);
nor U7713 (N_7713,N_7104,N_7342);
nand U7714 (N_7714,N_7477,N_7390);
nand U7715 (N_7715,N_7461,N_7417);
nor U7716 (N_7716,N_7074,N_7149);
and U7717 (N_7717,N_7223,N_7194);
or U7718 (N_7718,N_7358,N_7033);
and U7719 (N_7719,N_7380,N_7144);
nor U7720 (N_7720,N_7262,N_7134);
or U7721 (N_7721,N_7473,N_7270);
or U7722 (N_7722,N_7281,N_7121);
and U7723 (N_7723,N_7003,N_7436);
nor U7724 (N_7724,N_7382,N_7209);
xor U7725 (N_7725,N_7062,N_7044);
nor U7726 (N_7726,N_7485,N_7084);
nand U7727 (N_7727,N_7103,N_7188);
or U7728 (N_7728,N_7120,N_7478);
or U7729 (N_7729,N_7090,N_7499);
xor U7730 (N_7730,N_7280,N_7388);
or U7731 (N_7731,N_7027,N_7146);
or U7732 (N_7732,N_7401,N_7193);
nand U7733 (N_7733,N_7179,N_7233);
xnor U7734 (N_7734,N_7072,N_7337);
nand U7735 (N_7735,N_7381,N_7137);
xor U7736 (N_7736,N_7093,N_7489);
and U7737 (N_7737,N_7468,N_7333);
nand U7738 (N_7738,N_7470,N_7338);
nor U7739 (N_7739,N_7152,N_7249);
or U7740 (N_7740,N_7039,N_7140);
xor U7741 (N_7741,N_7115,N_7322);
and U7742 (N_7742,N_7029,N_7171);
nand U7743 (N_7743,N_7434,N_7339);
xnor U7744 (N_7744,N_7413,N_7393);
nor U7745 (N_7745,N_7432,N_7446);
or U7746 (N_7746,N_7252,N_7395);
and U7747 (N_7747,N_7175,N_7005);
and U7748 (N_7748,N_7466,N_7102);
or U7749 (N_7749,N_7173,N_7457);
nand U7750 (N_7750,N_7300,N_7133);
or U7751 (N_7751,N_7115,N_7360);
or U7752 (N_7752,N_7178,N_7272);
and U7753 (N_7753,N_7087,N_7371);
nand U7754 (N_7754,N_7068,N_7130);
nand U7755 (N_7755,N_7406,N_7218);
or U7756 (N_7756,N_7258,N_7307);
and U7757 (N_7757,N_7360,N_7173);
nand U7758 (N_7758,N_7448,N_7385);
and U7759 (N_7759,N_7483,N_7206);
or U7760 (N_7760,N_7355,N_7125);
nand U7761 (N_7761,N_7071,N_7209);
nand U7762 (N_7762,N_7296,N_7457);
nand U7763 (N_7763,N_7159,N_7034);
xnor U7764 (N_7764,N_7491,N_7323);
and U7765 (N_7765,N_7432,N_7198);
or U7766 (N_7766,N_7419,N_7344);
nand U7767 (N_7767,N_7345,N_7180);
nor U7768 (N_7768,N_7134,N_7053);
or U7769 (N_7769,N_7084,N_7017);
or U7770 (N_7770,N_7187,N_7315);
nor U7771 (N_7771,N_7494,N_7298);
nor U7772 (N_7772,N_7023,N_7321);
nor U7773 (N_7773,N_7253,N_7246);
and U7774 (N_7774,N_7393,N_7248);
or U7775 (N_7775,N_7389,N_7474);
nor U7776 (N_7776,N_7341,N_7387);
or U7777 (N_7777,N_7362,N_7399);
and U7778 (N_7778,N_7302,N_7179);
nor U7779 (N_7779,N_7131,N_7324);
and U7780 (N_7780,N_7144,N_7286);
and U7781 (N_7781,N_7432,N_7060);
nand U7782 (N_7782,N_7064,N_7430);
nand U7783 (N_7783,N_7411,N_7166);
nor U7784 (N_7784,N_7466,N_7428);
nor U7785 (N_7785,N_7209,N_7226);
nor U7786 (N_7786,N_7209,N_7493);
nand U7787 (N_7787,N_7225,N_7064);
or U7788 (N_7788,N_7040,N_7126);
xor U7789 (N_7789,N_7356,N_7253);
and U7790 (N_7790,N_7081,N_7178);
and U7791 (N_7791,N_7467,N_7027);
and U7792 (N_7792,N_7347,N_7178);
nand U7793 (N_7793,N_7139,N_7119);
xor U7794 (N_7794,N_7154,N_7111);
nand U7795 (N_7795,N_7234,N_7254);
nor U7796 (N_7796,N_7014,N_7407);
nor U7797 (N_7797,N_7399,N_7460);
xor U7798 (N_7798,N_7150,N_7478);
and U7799 (N_7799,N_7415,N_7284);
or U7800 (N_7800,N_7044,N_7289);
and U7801 (N_7801,N_7318,N_7361);
nor U7802 (N_7802,N_7496,N_7192);
nor U7803 (N_7803,N_7441,N_7424);
or U7804 (N_7804,N_7409,N_7093);
nand U7805 (N_7805,N_7353,N_7175);
and U7806 (N_7806,N_7094,N_7236);
nor U7807 (N_7807,N_7026,N_7488);
xor U7808 (N_7808,N_7197,N_7344);
nor U7809 (N_7809,N_7040,N_7150);
nor U7810 (N_7810,N_7072,N_7271);
or U7811 (N_7811,N_7373,N_7276);
nand U7812 (N_7812,N_7433,N_7002);
or U7813 (N_7813,N_7192,N_7085);
nand U7814 (N_7814,N_7090,N_7101);
or U7815 (N_7815,N_7483,N_7169);
nand U7816 (N_7816,N_7153,N_7080);
and U7817 (N_7817,N_7365,N_7152);
xor U7818 (N_7818,N_7101,N_7050);
or U7819 (N_7819,N_7005,N_7339);
nand U7820 (N_7820,N_7293,N_7285);
or U7821 (N_7821,N_7428,N_7045);
or U7822 (N_7822,N_7454,N_7470);
and U7823 (N_7823,N_7071,N_7004);
nor U7824 (N_7824,N_7352,N_7487);
xnor U7825 (N_7825,N_7186,N_7184);
and U7826 (N_7826,N_7469,N_7401);
and U7827 (N_7827,N_7416,N_7226);
and U7828 (N_7828,N_7098,N_7265);
xor U7829 (N_7829,N_7209,N_7395);
nor U7830 (N_7830,N_7085,N_7197);
nand U7831 (N_7831,N_7067,N_7342);
nand U7832 (N_7832,N_7015,N_7380);
or U7833 (N_7833,N_7108,N_7047);
xor U7834 (N_7834,N_7013,N_7300);
xor U7835 (N_7835,N_7098,N_7079);
and U7836 (N_7836,N_7262,N_7150);
nand U7837 (N_7837,N_7219,N_7231);
nand U7838 (N_7838,N_7100,N_7484);
or U7839 (N_7839,N_7257,N_7082);
nor U7840 (N_7840,N_7011,N_7028);
nand U7841 (N_7841,N_7372,N_7409);
and U7842 (N_7842,N_7105,N_7491);
nor U7843 (N_7843,N_7301,N_7289);
nor U7844 (N_7844,N_7123,N_7438);
and U7845 (N_7845,N_7145,N_7153);
nand U7846 (N_7846,N_7339,N_7277);
nor U7847 (N_7847,N_7114,N_7021);
nor U7848 (N_7848,N_7090,N_7383);
or U7849 (N_7849,N_7031,N_7111);
or U7850 (N_7850,N_7319,N_7355);
and U7851 (N_7851,N_7304,N_7416);
nand U7852 (N_7852,N_7433,N_7213);
and U7853 (N_7853,N_7158,N_7084);
or U7854 (N_7854,N_7319,N_7446);
or U7855 (N_7855,N_7373,N_7053);
and U7856 (N_7856,N_7412,N_7153);
or U7857 (N_7857,N_7469,N_7292);
and U7858 (N_7858,N_7323,N_7386);
nand U7859 (N_7859,N_7493,N_7352);
nor U7860 (N_7860,N_7095,N_7272);
nor U7861 (N_7861,N_7221,N_7164);
and U7862 (N_7862,N_7048,N_7492);
and U7863 (N_7863,N_7067,N_7364);
nor U7864 (N_7864,N_7236,N_7128);
nand U7865 (N_7865,N_7063,N_7374);
or U7866 (N_7866,N_7444,N_7304);
or U7867 (N_7867,N_7229,N_7272);
nand U7868 (N_7868,N_7204,N_7174);
and U7869 (N_7869,N_7185,N_7406);
nand U7870 (N_7870,N_7030,N_7217);
or U7871 (N_7871,N_7375,N_7291);
or U7872 (N_7872,N_7380,N_7080);
and U7873 (N_7873,N_7297,N_7265);
or U7874 (N_7874,N_7499,N_7311);
or U7875 (N_7875,N_7040,N_7355);
nor U7876 (N_7876,N_7338,N_7070);
and U7877 (N_7877,N_7187,N_7312);
and U7878 (N_7878,N_7388,N_7364);
nand U7879 (N_7879,N_7052,N_7298);
nand U7880 (N_7880,N_7022,N_7006);
or U7881 (N_7881,N_7460,N_7475);
nand U7882 (N_7882,N_7240,N_7443);
nand U7883 (N_7883,N_7348,N_7076);
nand U7884 (N_7884,N_7375,N_7483);
nand U7885 (N_7885,N_7318,N_7287);
nand U7886 (N_7886,N_7133,N_7276);
or U7887 (N_7887,N_7345,N_7121);
nor U7888 (N_7888,N_7095,N_7492);
and U7889 (N_7889,N_7172,N_7150);
nand U7890 (N_7890,N_7415,N_7177);
and U7891 (N_7891,N_7030,N_7393);
or U7892 (N_7892,N_7100,N_7336);
or U7893 (N_7893,N_7421,N_7245);
and U7894 (N_7894,N_7101,N_7234);
or U7895 (N_7895,N_7258,N_7070);
nand U7896 (N_7896,N_7060,N_7118);
nand U7897 (N_7897,N_7018,N_7377);
nand U7898 (N_7898,N_7088,N_7204);
or U7899 (N_7899,N_7370,N_7375);
nand U7900 (N_7900,N_7096,N_7188);
nand U7901 (N_7901,N_7092,N_7316);
xnor U7902 (N_7902,N_7154,N_7070);
nand U7903 (N_7903,N_7204,N_7443);
nand U7904 (N_7904,N_7230,N_7205);
and U7905 (N_7905,N_7352,N_7325);
and U7906 (N_7906,N_7363,N_7028);
and U7907 (N_7907,N_7087,N_7482);
nor U7908 (N_7908,N_7243,N_7269);
or U7909 (N_7909,N_7349,N_7153);
nand U7910 (N_7910,N_7108,N_7234);
nand U7911 (N_7911,N_7485,N_7346);
nand U7912 (N_7912,N_7243,N_7102);
and U7913 (N_7913,N_7104,N_7131);
nand U7914 (N_7914,N_7499,N_7011);
nor U7915 (N_7915,N_7485,N_7497);
nor U7916 (N_7916,N_7210,N_7212);
or U7917 (N_7917,N_7454,N_7021);
nand U7918 (N_7918,N_7113,N_7448);
nand U7919 (N_7919,N_7001,N_7000);
and U7920 (N_7920,N_7237,N_7084);
or U7921 (N_7921,N_7309,N_7276);
nor U7922 (N_7922,N_7097,N_7002);
or U7923 (N_7923,N_7309,N_7095);
nor U7924 (N_7924,N_7402,N_7006);
xnor U7925 (N_7925,N_7240,N_7385);
nand U7926 (N_7926,N_7490,N_7007);
nand U7927 (N_7927,N_7098,N_7135);
nor U7928 (N_7928,N_7036,N_7053);
nand U7929 (N_7929,N_7147,N_7172);
nand U7930 (N_7930,N_7003,N_7174);
nand U7931 (N_7931,N_7186,N_7209);
and U7932 (N_7932,N_7184,N_7183);
xnor U7933 (N_7933,N_7017,N_7184);
nor U7934 (N_7934,N_7427,N_7185);
xor U7935 (N_7935,N_7231,N_7410);
and U7936 (N_7936,N_7168,N_7242);
or U7937 (N_7937,N_7210,N_7229);
and U7938 (N_7938,N_7253,N_7035);
and U7939 (N_7939,N_7106,N_7266);
and U7940 (N_7940,N_7376,N_7151);
or U7941 (N_7941,N_7252,N_7262);
or U7942 (N_7942,N_7097,N_7353);
and U7943 (N_7943,N_7227,N_7401);
nor U7944 (N_7944,N_7040,N_7207);
nor U7945 (N_7945,N_7349,N_7159);
or U7946 (N_7946,N_7024,N_7235);
nand U7947 (N_7947,N_7118,N_7363);
nand U7948 (N_7948,N_7384,N_7395);
or U7949 (N_7949,N_7216,N_7094);
and U7950 (N_7950,N_7395,N_7101);
nor U7951 (N_7951,N_7020,N_7328);
nand U7952 (N_7952,N_7288,N_7466);
or U7953 (N_7953,N_7372,N_7338);
or U7954 (N_7954,N_7226,N_7398);
or U7955 (N_7955,N_7250,N_7106);
and U7956 (N_7956,N_7415,N_7495);
or U7957 (N_7957,N_7076,N_7135);
nor U7958 (N_7958,N_7287,N_7241);
and U7959 (N_7959,N_7441,N_7127);
and U7960 (N_7960,N_7249,N_7188);
xnor U7961 (N_7961,N_7042,N_7195);
nor U7962 (N_7962,N_7070,N_7209);
or U7963 (N_7963,N_7197,N_7465);
and U7964 (N_7964,N_7270,N_7145);
and U7965 (N_7965,N_7496,N_7424);
or U7966 (N_7966,N_7067,N_7390);
nand U7967 (N_7967,N_7146,N_7314);
and U7968 (N_7968,N_7307,N_7134);
or U7969 (N_7969,N_7346,N_7311);
xor U7970 (N_7970,N_7425,N_7206);
nor U7971 (N_7971,N_7474,N_7052);
and U7972 (N_7972,N_7099,N_7268);
and U7973 (N_7973,N_7211,N_7261);
and U7974 (N_7974,N_7328,N_7055);
and U7975 (N_7975,N_7152,N_7197);
or U7976 (N_7976,N_7142,N_7113);
nor U7977 (N_7977,N_7088,N_7031);
or U7978 (N_7978,N_7198,N_7071);
and U7979 (N_7979,N_7398,N_7107);
or U7980 (N_7980,N_7478,N_7029);
nand U7981 (N_7981,N_7167,N_7032);
nor U7982 (N_7982,N_7014,N_7294);
or U7983 (N_7983,N_7218,N_7114);
or U7984 (N_7984,N_7039,N_7346);
and U7985 (N_7985,N_7317,N_7344);
xnor U7986 (N_7986,N_7061,N_7007);
or U7987 (N_7987,N_7123,N_7019);
or U7988 (N_7988,N_7471,N_7357);
nand U7989 (N_7989,N_7104,N_7434);
and U7990 (N_7990,N_7337,N_7211);
or U7991 (N_7991,N_7010,N_7126);
and U7992 (N_7992,N_7442,N_7410);
or U7993 (N_7993,N_7102,N_7346);
and U7994 (N_7994,N_7169,N_7467);
nor U7995 (N_7995,N_7429,N_7014);
nor U7996 (N_7996,N_7309,N_7347);
and U7997 (N_7997,N_7193,N_7283);
nor U7998 (N_7998,N_7321,N_7184);
nor U7999 (N_7999,N_7322,N_7055);
or U8000 (N_8000,N_7716,N_7556);
nor U8001 (N_8001,N_7818,N_7824);
and U8002 (N_8002,N_7681,N_7904);
nand U8003 (N_8003,N_7910,N_7685);
or U8004 (N_8004,N_7687,N_7867);
or U8005 (N_8005,N_7709,N_7680);
or U8006 (N_8006,N_7649,N_7714);
or U8007 (N_8007,N_7984,N_7719);
nor U8008 (N_8008,N_7917,N_7964);
nand U8009 (N_8009,N_7752,N_7540);
nand U8010 (N_8010,N_7953,N_7675);
and U8011 (N_8011,N_7574,N_7857);
and U8012 (N_8012,N_7784,N_7554);
xnor U8013 (N_8013,N_7549,N_7771);
nor U8014 (N_8014,N_7885,N_7564);
xor U8015 (N_8015,N_7624,N_7977);
and U8016 (N_8016,N_7897,N_7656);
nand U8017 (N_8017,N_7503,N_7748);
or U8018 (N_8018,N_7844,N_7889);
nand U8019 (N_8019,N_7912,N_7536);
nor U8020 (N_8020,N_7699,N_7636);
nor U8021 (N_8021,N_7873,N_7901);
or U8022 (N_8022,N_7941,N_7756);
nor U8023 (N_8023,N_7583,N_7836);
and U8024 (N_8024,N_7573,N_7981);
xnor U8025 (N_8025,N_7864,N_7866);
and U8026 (N_8026,N_7999,N_7787);
xnor U8027 (N_8027,N_7957,N_7563);
nor U8028 (N_8028,N_7750,N_7820);
or U8029 (N_8029,N_7821,N_7913);
xnor U8030 (N_8030,N_7923,N_7764);
nand U8031 (N_8031,N_7770,N_7749);
or U8032 (N_8032,N_7918,N_7751);
and U8033 (N_8033,N_7880,N_7978);
nor U8034 (N_8034,N_7516,N_7755);
nand U8035 (N_8035,N_7620,N_7562);
xnor U8036 (N_8036,N_7733,N_7965);
nand U8037 (N_8037,N_7854,N_7850);
xor U8038 (N_8038,N_7872,N_7853);
nor U8039 (N_8039,N_7782,N_7829);
nand U8040 (N_8040,N_7647,N_7689);
nand U8041 (N_8041,N_7623,N_7790);
xor U8042 (N_8042,N_7543,N_7676);
and U8043 (N_8043,N_7891,N_7786);
nand U8044 (N_8044,N_7712,N_7892);
xor U8045 (N_8045,N_7519,N_7505);
nor U8046 (N_8046,N_7518,N_7870);
nor U8047 (N_8047,N_7906,N_7930);
nand U8048 (N_8048,N_7601,N_7724);
nor U8049 (N_8049,N_7753,N_7665);
nor U8050 (N_8050,N_7718,N_7527);
nand U8051 (N_8051,N_7808,N_7572);
and U8052 (N_8052,N_7560,N_7881);
nand U8053 (N_8053,N_7736,N_7937);
nor U8054 (N_8054,N_7781,N_7926);
nand U8055 (N_8055,N_7759,N_7640);
nand U8056 (N_8056,N_7666,N_7667);
xor U8057 (N_8057,N_7807,N_7785);
or U8058 (N_8058,N_7883,N_7994);
nor U8059 (N_8059,N_7534,N_7946);
nand U8060 (N_8060,N_7542,N_7991);
or U8061 (N_8061,N_7731,N_7529);
and U8062 (N_8062,N_7566,N_7802);
or U8063 (N_8063,N_7662,N_7945);
nand U8064 (N_8064,N_7960,N_7581);
nor U8065 (N_8065,N_7805,N_7793);
xnor U8066 (N_8066,N_7874,N_7695);
or U8067 (N_8067,N_7800,N_7696);
nor U8068 (N_8068,N_7679,N_7828);
nor U8069 (N_8069,N_7561,N_7803);
nor U8070 (N_8070,N_7940,N_7924);
or U8071 (N_8071,N_7952,N_7726);
or U8072 (N_8072,N_7638,N_7763);
and U8073 (N_8073,N_7688,N_7510);
xnor U8074 (N_8074,N_7641,N_7979);
nand U8075 (N_8075,N_7730,N_7773);
nand U8076 (N_8076,N_7980,N_7630);
nor U8077 (N_8077,N_7590,N_7502);
and U8078 (N_8078,N_7603,N_7970);
nor U8079 (N_8079,N_7959,N_7929);
nand U8080 (N_8080,N_7740,N_7531);
and U8081 (N_8081,N_7919,N_7791);
and U8082 (N_8082,N_7944,N_7758);
or U8083 (N_8083,N_7890,N_7963);
nor U8084 (N_8084,N_7839,N_7512);
and U8085 (N_8085,N_7810,N_7899);
nand U8086 (N_8086,N_7742,N_7522);
or U8087 (N_8087,N_7673,N_7815);
xnor U8088 (N_8088,N_7738,N_7727);
nand U8089 (N_8089,N_7767,N_7723);
nand U8090 (N_8090,N_7911,N_7938);
or U8091 (N_8091,N_7691,N_7859);
nor U8092 (N_8092,N_7831,N_7863);
and U8093 (N_8093,N_7615,N_7703);
nor U8094 (N_8094,N_7878,N_7697);
and U8095 (N_8095,N_7648,N_7580);
nor U8096 (N_8096,N_7823,N_7757);
or U8097 (N_8097,N_7969,N_7795);
xnor U8098 (N_8098,N_7548,N_7611);
nor U8099 (N_8099,N_7928,N_7506);
or U8100 (N_8100,N_7642,N_7639);
or U8101 (N_8101,N_7879,N_7565);
and U8102 (N_8102,N_7520,N_7700);
or U8103 (N_8103,N_7760,N_7794);
and U8104 (N_8104,N_7728,N_7812);
nand U8105 (N_8105,N_7706,N_7674);
or U8106 (N_8106,N_7544,N_7582);
and U8107 (N_8107,N_7567,N_7684);
nor U8108 (N_8108,N_7663,N_7898);
or U8109 (N_8109,N_7729,N_7942);
nand U8110 (N_8110,N_7600,N_7933);
xnor U8111 (N_8111,N_7998,N_7985);
and U8112 (N_8112,N_7597,N_7916);
and U8113 (N_8113,N_7683,N_7775);
and U8114 (N_8114,N_7816,N_7806);
xnor U8115 (N_8115,N_7652,N_7523);
or U8116 (N_8116,N_7988,N_7651);
nor U8117 (N_8117,N_7949,N_7954);
or U8118 (N_8118,N_7989,N_7504);
nand U8119 (N_8119,N_7833,N_7846);
or U8120 (N_8120,N_7826,N_7672);
or U8121 (N_8121,N_7605,N_7845);
nor U8122 (N_8122,N_7875,N_7990);
nand U8123 (N_8123,N_7576,N_7704);
nor U8124 (N_8124,N_7765,N_7653);
nand U8125 (N_8125,N_7609,N_7788);
and U8126 (N_8126,N_7645,N_7617);
nand U8127 (N_8127,N_7628,N_7589);
nor U8128 (N_8128,N_7678,N_7779);
nor U8129 (N_8129,N_7511,N_7555);
and U8130 (N_8130,N_7721,N_7622);
or U8131 (N_8131,N_7995,N_7902);
or U8132 (N_8132,N_7961,N_7837);
and U8133 (N_8133,N_7903,N_7849);
nor U8134 (N_8134,N_7587,N_7643);
nand U8135 (N_8135,N_7635,N_7947);
xnor U8136 (N_8136,N_7974,N_7508);
and U8137 (N_8137,N_7705,N_7896);
nand U8138 (N_8138,N_7644,N_7943);
or U8139 (N_8139,N_7914,N_7935);
nand U8140 (N_8140,N_7967,N_7876);
nor U8141 (N_8141,N_7661,N_7655);
nor U8142 (N_8142,N_7993,N_7578);
and U8143 (N_8143,N_7625,N_7690);
nor U8144 (N_8144,N_7936,N_7834);
or U8145 (N_8145,N_7804,N_7595);
nor U8146 (N_8146,N_7732,N_7575);
nor U8147 (N_8147,N_7746,N_7925);
and U8148 (N_8148,N_7801,N_7702);
nor U8149 (N_8149,N_7677,N_7830);
or U8150 (N_8150,N_7517,N_7530);
nand U8151 (N_8151,N_7604,N_7692);
or U8152 (N_8152,N_7737,N_7743);
and U8153 (N_8153,N_7822,N_7934);
nor U8154 (N_8154,N_7832,N_7840);
nand U8155 (N_8155,N_7907,N_7921);
or U8156 (N_8156,N_7533,N_7707);
or U8157 (N_8157,N_7766,N_7900);
or U8158 (N_8158,N_7621,N_7966);
nand U8159 (N_8159,N_7618,N_7931);
and U8160 (N_8160,N_7825,N_7847);
or U8161 (N_8161,N_7976,N_7722);
nand U8162 (N_8162,N_7525,N_7660);
nand U8163 (N_8163,N_7552,N_7658);
nand U8164 (N_8164,N_7893,N_7762);
nand U8165 (N_8165,N_7813,N_7586);
or U8166 (N_8166,N_7860,N_7524);
and U8167 (N_8167,N_7588,N_7777);
or U8168 (N_8168,N_7594,N_7986);
nand U8169 (N_8169,N_7962,N_7789);
xor U8170 (N_8170,N_7670,N_7838);
or U8171 (N_8171,N_7550,N_7532);
xnor U8172 (N_8172,N_7598,N_7778);
and U8173 (N_8173,N_7920,N_7637);
and U8174 (N_8174,N_7915,N_7591);
nor U8175 (N_8175,N_7553,N_7894);
and U8176 (N_8176,N_7886,N_7772);
xnor U8177 (N_8177,N_7796,N_7535);
or U8178 (N_8178,N_7541,N_7577);
nor U8179 (N_8179,N_7814,N_7877);
nor U8180 (N_8180,N_7711,N_7708);
nand U8181 (N_8181,N_7551,N_7629);
nor U8182 (N_8182,N_7528,N_7570);
nor U8183 (N_8183,N_7848,N_7776);
or U8184 (N_8184,N_7811,N_7659);
nor U8185 (N_8185,N_7817,N_7694);
and U8186 (N_8186,N_7614,N_7932);
or U8187 (N_8187,N_7507,N_7725);
or U8188 (N_8188,N_7513,N_7698);
or U8189 (N_8189,N_7858,N_7654);
nor U8190 (N_8190,N_7558,N_7693);
nand U8191 (N_8191,N_7851,N_7871);
nand U8192 (N_8192,N_7927,N_7747);
and U8193 (N_8193,N_7869,N_7633);
or U8194 (N_8194,N_7909,N_7882);
nand U8195 (N_8195,N_7809,N_7599);
or U8196 (N_8196,N_7739,N_7593);
nor U8197 (N_8197,N_7741,N_7717);
nor U8198 (N_8198,N_7735,N_7884);
nand U8199 (N_8199,N_7514,N_7987);
nand U8200 (N_8200,N_7922,N_7650);
and U8201 (N_8201,N_7610,N_7626);
and U8202 (N_8202,N_7657,N_7632);
or U8203 (N_8203,N_7571,N_7557);
nand U8204 (N_8204,N_7537,N_7612);
and U8205 (N_8205,N_7955,N_7865);
or U8206 (N_8206,N_7956,N_7569);
nand U8207 (N_8207,N_7862,N_7861);
and U8208 (N_8208,N_7819,N_7501);
nor U8209 (N_8209,N_7843,N_7579);
and U8210 (N_8210,N_7592,N_7547);
or U8211 (N_8211,N_7608,N_7734);
or U8212 (N_8212,N_7888,N_7546);
or U8213 (N_8213,N_7968,N_7631);
nor U8214 (N_8214,N_7958,N_7526);
and U8215 (N_8215,N_7613,N_7539);
or U8216 (N_8216,N_7842,N_7792);
and U8217 (N_8217,N_7701,N_7798);
xnor U8218 (N_8218,N_7634,N_7686);
or U8219 (N_8219,N_7559,N_7973);
or U8220 (N_8220,N_7852,N_7538);
or U8221 (N_8221,N_7521,N_7768);
xnor U8222 (N_8222,N_7500,N_7908);
or U8223 (N_8223,N_7744,N_7887);
or U8224 (N_8224,N_7568,N_7948);
nand U8225 (N_8225,N_7783,N_7545);
nor U8226 (N_8226,N_7671,N_7754);
and U8227 (N_8227,N_7509,N_7616);
nor U8228 (N_8228,N_7585,N_7596);
and U8229 (N_8229,N_7905,N_7682);
and U8230 (N_8230,N_7627,N_7607);
nor U8231 (N_8231,N_7950,N_7895);
or U8232 (N_8232,N_7799,N_7606);
nand U8233 (N_8233,N_7983,N_7515);
nand U8234 (N_8234,N_7835,N_7996);
nand U8235 (N_8235,N_7797,N_7856);
or U8236 (N_8236,N_7713,N_7715);
nand U8237 (N_8237,N_7975,N_7939);
xnor U8238 (N_8238,N_7720,N_7972);
or U8239 (N_8239,N_7710,N_7669);
xnor U8240 (N_8240,N_7780,N_7868);
nor U8241 (N_8241,N_7584,N_7992);
xor U8242 (N_8242,N_7971,N_7769);
or U8243 (N_8243,N_7664,N_7668);
nor U8244 (N_8244,N_7602,N_7841);
or U8245 (N_8245,N_7827,N_7982);
or U8246 (N_8246,N_7774,N_7997);
or U8247 (N_8247,N_7619,N_7951);
nand U8248 (N_8248,N_7855,N_7745);
nand U8249 (N_8249,N_7646,N_7761);
nor U8250 (N_8250,N_7645,N_7751);
nor U8251 (N_8251,N_7754,N_7998);
and U8252 (N_8252,N_7740,N_7921);
nand U8253 (N_8253,N_7609,N_7501);
nand U8254 (N_8254,N_7863,N_7989);
xnor U8255 (N_8255,N_7964,N_7642);
or U8256 (N_8256,N_7807,N_7929);
nor U8257 (N_8257,N_7706,N_7610);
and U8258 (N_8258,N_7790,N_7684);
xnor U8259 (N_8259,N_7979,N_7953);
nor U8260 (N_8260,N_7589,N_7630);
or U8261 (N_8261,N_7967,N_7904);
xnor U8262 (N_8262,N_7599,N_7795);
and U8263 (N_8263,N_7941,N_7819);
nor U8264 (N_8264,N_7938,N_7853);
xnor U8265 (N_8265,N_7902,N_7765);
or U8266 (N_8266,N_7953,N_7869);
or U8267 (N_8267,N_7758,N_7936);
nand U8268 (N_8268,N_7948,N_7710);
nor U8269 (N_8269,N_7935,N_7793);
nand U8270 (N_8270,N_7755,N_7807);
nand U8271 (N_8271,N_7637,N_7554);
nor U8272 (N_8272,N_7869,N_7559);
nand U8273 (N_8273,N_7674,N_7812);
nor U8274 (N_8274,N_7791,N_7993);
and U8275 (N_8275,N_7665,N_7594);
and U8276 (N_8276,N_7729,N_7566);
or U8277 (N_8277,N_7730,N_7822);
and U8278 (N_8278,N_7757,N_7648);
nand U8279 (N_8279,N_7615,N_7595);
xnor U8280 (N_8280,N_7989,N_7677);
or U8281 (N_8281,N_7902,N_7920);
or U8282 (N_8282,N_7579,N_7858);
nor U8283 (N_8283,N_7706,N_7752);
or U8284 (N_8284,N_7766,N_7853);
nand U8285 (N_8285,N_7734,N_7710);
nand U8286 (N_8286,N_7603,N_7581);
nand U8287 (N_8287,N_7780,N_7840);
nor U8288 (N_8288,N_7795,N_7886);
nand U8289 (N_8289,N_7904,N_7976);
nor U8290 (N_8290,N_7512,N_7914);
or U8291 (N_8291,N_7670,N_7830);
nor U8292 (N_8292,N_7582,N_7785);
nor U8293 (N_8293,N_7967,N_7510);
nand U8294 (N_8294,N_7890,N_7766);
nand U8295 (N_8295,N_7545,N_7784);
nand U8296 (N_8296,N_7560,N_7750);
nor U8297 (N_8297,N_7713,N_7975);
or U8298 (N_8298,N_7950,N_7746);
and U8299 (N_8299,N_7885,N_7722);
and U8300 (N_8300,N_7619,N_7999);
nor U8301 (N_8301,N_7838,N_7532);
nor U8302 (N_8302,N_7549,N_7564);
or U8303 (N_8303,N_7746,N_7751);
nand U8304 (N_8304,N_7907,N_7737);
nor U8305 (N_8305,N_7575,N_7876);
nand U8306 (N_8306,N_7606,N_7749);
nand U8307 (N_8307,N_7786,N_7772);
nand U8308 (N_8308,N_7582,N_7808);
nor U8309 (N_8309,N_7606,N_7876);
nor U8310 (N_8310,N_7692,N_7854);
nor U8311 (N_8311,N_7584,N_7632);
nand U8312 (N_8312,N_7742,N_7663);
xnor U8313 (N_8313,N_7914,N_7936);
or U8314 (N_8314,N_7611,N_7659);
or U8315 (N_8315,N_7636,N_7768);
nor U8316 (N_8316,N_7654,N_7795);
and U8317 (N_8317,N_7565,N_7514);
and U8318 (N_8318,N_7990,N_7548);
or U8319 (N_8319,N_7806,N_7900);
nand U8320 (N_8320,N_7802,N_7578);
and U8321 (N_8321,N_7981,N_7990);
or U8322 (N_8322,N_7787,N_7627);
nand U8323 (N_8323,N_7579,N_7519);
nand U8324 (N_8324,N_7519,N_7555);
or U8325 (N_8325,N_7575,N_7627);
nor U8326 (N_8326,N_7747,N_7698);
and U8327 (N_8327,N_7566,N_7633);
nand U8328 (N_8328,N_7731,N_7634);
xnor U8329 (N_8329,N_7731,N_7796);
nor U8330 (N_8330,N_7977,N_7981);
or U8331 (N_8331,N_7553,N_7664);
and U8332 (N_8332,N_7884,N_7826);
nand U8333 (N_8333,N_7945,N_7674);
nand U8334 (N_8334,N_7735,N_7526);
or U8335 (N_8335,N_7905,N_7945);
or U8336 (N_8336,N_7778,N_7938);
nor U8337 (N_8337,N_7602,N_7811);
or U8338 (N_8338,N_7989,N_7755);
and U8339 (N_8339,N_7534,N_7914);
and U8340 (N_8340,N_7645,N_7582);
xor U8341 (N_8341,N_7582,N_7973);
and U8342 (N_8342,N_7953,N_7815);
nand U8343 (N_8343,N_7757,N_7733);
nor U8344 (N_8344,N_7830,N_7601);
nand U8345 (N_8345,N_7794,N_7645);
nand U8346 (N_8346,N_7856,N_7813);
or U8347 (N_8347,N_7544,N_7877);
nand U8348 (N_8348,N_7648,N_7898);
or U8349 (N_8349,N_7511,N_7507);
nand U8350 (N_8350,N_7746,N_7693);
or U8351 (N_8351,N_7801,N_7579);
or U8352 (N_8352,N_7702,N_7617);
nor U8353 (N_8353,N_7779,N_7840);
xnor U8354 (N_8354,N_7621,N_7528);
nor U8355 (N_8355,N_7746,N_7601);
and U8356 (N_8356,N_7777,N_7972);
nor U8357 (N_8357,N_7813,N_7845);
and U8358 (N_8358,N_7767,N_7914);
and U8359 (N_8359,N_7848,N_7727);
nand U8360 (N_8360,N_7944,N_7710);
xnor U8361 (N_8361,N_7883,N_7548);
and U8362 (N_8362,N_7650,N_7966);
nor U8363 (N_8363,N_7599,N_7856);
or U8364 (N_8364,N_7811,N_7993);
or U8365 (N_8365,N_7836,N_7892);
nor U8366 (N_8366,N_7570,N_7898);
nor U8367 (N_8367,N_7541,N_7622);
nand U8368 (N_8368,N_7542,N_7978);
and U8369 (N_8369,N_7578,N_7607);
or U8370 (N_8370,N_7855,N_7634);
xor U8371 (N_8371,N_7898,N_7527);
nand U8372 (N_8372,N_7601,N_7815);
nor U8373 (N_8373,N_7594,N_7638);
and U8374 (N_8374,N_7926,N_7829);
or U8375 (N_8375,N_7903,N_7751);
nor U8376 (N_8376,N_7936,N_7871);
nand U8377 (N_8377,N_7963,N_7742);
or U8378 (N_8378,N_7965,N_7639);
or U8379 (N_8379,N_7663,N_7609);
nand U8380 (N_8380,N_7528,N_7926);
nor U8381 (N_8381,N_7780,N_7591);
and U8382 (N_8382,N_7804,N_7874);
nand U8383 (N_8383,N_7506,N_7594);
xnor U8384 (N_8384,N_7540,N_7655);
and U8385 (N_8385,N_7511,N_7691);
xnor U8386 (N_8386,N_7822,N_7965);
xor U8387 (N_8387,N_7990,N_7529);
or U8388 (N_8388,N_7978,N_7955);
nor U8389 (N_8389,N_7782,N_7837);
nor U8390 (N_8390,N_7602,N_7994);
and U8391 (N_8391,N_7639,N_7898);
or U8392 (N_8392,N_7707,N_7518);
and U8393 (N_8393,N_7928,N_7622);
nor U8394 (N_8394,N_7926,N_7658);
nand U8395 (N_8395,N_7518,N_7716);
nand U8396 (N_8396,N_7807,N_7616);
nand U8397 (N_8397,N_7604,N_7919);
nor U8398 (N_8398,N_7519,N_7806);
nand U8399 (N_8399,N_7958,N_7601);
nor U8400 (N_8400,N_7918,N_7645);
nand U8401 (N_8401,N_7667,N_7719);
nand U8402 (N_8402,N_7641,N_7523);
or U8403 (N_8403,N_7671,N_7594);
nand U8404 (N_8404,N_7899,N_7974);
xnor U8405 (N_8405,N_7899,N_7504);
nor U8406 (N_8406,N_7973,N_7736);
xor U8407 (N_8407,N_7804,N_7562);
nand U8408 (N_8408,N_7944,N_7504);
nand U8409 (N_8409,N_7803,N_7751);
or U8410 (N_8410,N_7550,N_7862);
nand U8411 (N_8411,N_7843,N_7598);
nor U8412 (N_8412,N_7529,N_7605);
and U8413 (N_8413,N_7838,N_7649);
nor U8414 (N_8414,N_7599,N_7995);
or U8415 (N_8415,N_7984,N_7674);
and U8416 (N_8416,N_7779,N_7882);
nor U8417 (N_8417,N_7635,N_7934);
xnor U8418 (N_8418,N_7863,N_7591);
and U8419 (N_8419,N_7517,N_7983);
nand U8420 (N_8420,N_7788,N_7653);
nand U8421 (N_8421,N_7772,N_7979);
nand U8422 (N_8422,N_7595,N_7581);
and U8423 (N_8423,N_7677,N_7905);
nand U8424 (N_8424,N_7861,N_7883);
or U8425 (N_8425,N_7879,N_7651);
nand U8426 (N_8426,N_7677,N_7894);
nor U8427 (N_8427,N_7809,N_7954);
nor U8428 (N_8428,N_7861,N_7511);
nor U8429 (N_8429,N_7587,N_7729);
nor U8430 (N_8430,N_7519,N_7523);
nor U8431 (N_8431,N_7674,N_7808);
and U8432 (N_8432,N_7596,N_7720);
or U8433 (N_8433,N_7697,N_7957);
and U8434 (N_8434,N_7632,N_7638);
or U8435 (N_8435,N_7961,N_7736);
and U8436 (N_8436,N_7744,N_7503);
xnor U8437 (N_8437,N_7661,N_7958);
nand U8438 (N_8438,N_7562,N_7506);
nand U8439 (N_8439,N_7710,N_7712);
nor U8440 (N_8440,N_7504,N_7545);
or U8441 (N_8441,N_7966,N_7849);
nand U8442 (N_8442,N_7770,N_7898);
nand U8443 (N_8443,N_7977,N_7993);
and U8444 (N_8444,N_7740,N_7557);
nand U8445 (N_8445,N_7604,N_7950);
nor U8446 (N_8446,N_7639,N_7760);
or U8447 (N_8447,N_7599,N_7593);
nand U8448 (N_8448,N_7703,N_7707);
nor U8449 (N_8449,N_7898,N_7932);
or U8450 (N_8450,N_7835,N_7792);
nand U8451 (N_8451,N_7752,N_7597);
and U8452 (N_8452,N_7828,N_7723);
and U8453 (N_8453,N_7619,N_7981);
nor U8454 (N_8454,N_7823,N_7959);
or U8455 (N_8455,N_7733,N_7682);
nor U8456 (N_8456,N_7651,N_7994);
xor U8457 (N_8457,N_7670,N_7978);
nor U8458 (N_8458,N_7598,N_7518);
and U8459 (N_8459,N_7638,N_7926);
nor U8460 (N_8460,N_7941,N_7948);
nand U8461 (N_8461,N_7768,N_7619);
xor U8462 (N_8462,N_7501,N_7733);
xnor U8463 (N_8463,N_7618,N_7815);
nor U8464 (N_8464,N_7809,N_7535);
or U8465 (N_8465,N_7988,N_7635);
nor U8466 (N_8466,N_7785,N_7932);
nand U8467 (N_8467,N_7693,N_7776);
and U8468 (N_8468,N_7693,N_7902);
and U8469 (N_8469,N_7702,N_7594);
xnor U8470 (N_8470,N_7837,N_7768);
xor U8471 (N_8471,N_7748,N_7679);
or U8472 (N_8472,N_7510,N_7859);
nor U8473 (N_8473,N_7928,N_7864);
or U8474 (N_8474,N_7553,N_7592);
nor U8475 (N_8475,N_7910,N_7694);
nor U8476 (N_8476,N_7864,N_7548);
or U8477 (N_8477,N_7631,N_7703);
nor U8478 (N_8478,N_7879,N_7710);
nand U8479 (N_8479,N_7697,N_7765);
nand U8480 (N_8480,N_7956,N_7592);
and U8481 (N_8481,N_7508,N_7729);
or U8482 (N_8482,N_7681,N_7616);
nand U8483 (N_8483,N_7993,N_7581);
and U8484 (N_8484,N_7542,N_7820);
or U8485 (N_8485,N_7646,N_7901);
nand U8486 (N_8486,N_7662,N_7678);
or U8487 (N_8487,N_7994,N_7946);
or U8488 (N_8488,N_7955,N_7983);
and U8489 (N_8489,N_7773,N_7883);
nor U8490 (N_8490,N_7898,N_7718);
nor U8491 (N_8491,N_7584,N_7681);
nand U8492 (N_8492,N_7882,N_7535);
and U8493 (N_8493,N_7770,N_7792);
or U8494 (N_8494,N_7878,N_7557);
or U8495 (N_8495,N_7929,N_7919);
and U8496 (N_8496,N_7829,N_7572);
nand U8497 (N_8497,N_7986,N_7640);
and U8498 (N_8498,N_7557,N_7849);
or U8499 (N_8499,N_7764,N_7927);
or U8500 (N_8500,N_8396,N_8031);
or U8501 (N_8501,N_8280,N_8029);
and U8502 (N_8502,N_8171,N_8145);
nand U8503 (N_8503,N_8248,N_8271);
and U8504 (N_8504,N_8320,N_8426);
nand U8505 (N_8505,N_8012,N_8188);
nand U8506 (N_8506,N_8090,N_8002);
nor U8507 (N_8507,N_8139,N_8018);
nand U8508 (N_8508,N_8008,N_8128);
nand U8509 (N_8509,N_8075,N_8352);
xor U8510 (N_8510,N_8085,N_8350);
nand U8511 (N_8511,N_8419,N_8296);
or U8512 (N_8512,N_8198,N_8456);
nand U8513 (N_8513,N_8308,N_8366);
nor U8514 (N_8514,N_8066,N_8205);
nor U8515 (N_8515,N_8411,N_8123);
nand U8516 (N_8516,N_8047,N_8038);
nor U8517 (N_8517,N_8292,N_8192);
or U8518 (N_8518,N_8381,N_8473);
or U8519 (N_8519,N_8255,N_8273);
nor U8520 (N_8520,N_8096,N_8362);
and U8521 (N_8521,N_8001,N_8113);
nor U8522 (N_8522,N_8226,N_8187);
nor U8523 (N_8523,N_8441,N_8234);
nand U8524 (N_8524,N_8247,N_8448);
and U8525 (N_8525,N_8332,N_8121);
or U8526 (N_8526,N_8376,N_8369);
nand U8527 (N_8527,N_8081,N_8256);
and U8528 (N_8528,N_8203,N_8404);
xor U8529 (N_8529,N_8379,N_8326);
nor U8530 (N_8530,N_8418,N_8499);
nand U8531 (N_8531,N_8231,N_8457);
and U8532 (N_8532,N_8216,N_8471);
nor U8533 (N_8533,N_8071,N_8353);
nor U8534 (N_8534,N_8070,N_8080);
and U8535 (N_8535,N_8475,N_8218);
nand U8536 (N_8536,N_8427,N_8005);
and U8537 (N_8537,N_8264,N_8275);
and U8538 (N_8538,N_8485,N_8133);
or U8539 (N_8539,N_8345,N_8351);
xor U8540 (N_8540,N_8490,N_8309);
and U8541 (N_8541,N_8470,N_8385);
nand U8542 (N_8542,N_8030,N_8207);
nand U8543 (N_8543,N_8194,N_8233);
nor U8544 (N_8544,N_8295,N_8115);
nand U8545 (N_8545,N_8152,N_8259);
nand U8546 (N_8546,N_8151,N_8342);
nand U8547 (N_8547,N_8331,N_8043);
and U8548 (N_8548,N_8314,N_8103);
xor U8549 (N_8549,N_8484,N_8267);
and U8550 (N_8550,N_8368,N_8229);
or U8551 (N_8551,N_8202,N_8444);
nor U8552 (N_8552,N_8023,N_8169);
xor U8553 (N_8553,N_8108,N_8057);
and U8554 (N_8554,N_8114,N_8390);
and U8555 (N_8555,N_8330,N_8349);
nand U8556 (N_8556,N_8091,N_8336);
nor U8557 (N_8557,N_8403,N_8304);
and U8558 (N_8558,N_8482,N_8027);
or U8559 (N_8559,N_8084,N_8069);
nor U8560 (N_8560,N_8011,N_8321);
and U8561 (N_8561,N_8469,N_8293);
nand U8562 (N_8562,N_8380,N_8065);
nand U8563 (N_8563,N_8285,N_8077);
and U8564 (N_8564,N_8373,N_8180);
or U8565 (N_8565,N_8028,N_8250);
nand U8566 (N_8566,N_8260,N_8239);
or U8567 (N_8567,N_8118,N_8127);
nand U8568 (N_8568,N_8061,N_8409);
xnor U8569 (N_8569,N_8261,N_8182);
or U8570 (N_8570,N_8044,N_8442);
and U8571 (N_8571,N_8476,N_8064);
nand U8572 (N_8572,N_8284,N_8372);
nand U8573 (N_8573,N_8214,N_8463);
nor U8574 (N_8574,N_8060,N_8094);
and U8575 (N_8575,N_8324,N_8245);
and U8576 (N_8576,N_8298,N_8278);
nand U8577 (N_8577,N_8241,N_8343);
or U8578 (N_8578,N_8240,N_8365);
and U8579 (N_8579,N_8399,N_8126);
nand U8580 (N_8580,N_8270,N_8022);
nor U8581 (N_8581,N_8257,N_8406);
and U8582 (N_8582,N_8004,N_8143);
xor U8583 (N_8583,N_8333,N_8106);
nor U8584 (N_8584,N_8179,N_8007);
nor U8585 (N_8585,N_8410,N_8196);
nand U8586 (N_8586,N_8281,N_8166);
xor U8587 (N_8587,N_8052,N_8048);
nand U8588 (N_8588,N_8093,N_8167);
nor U8589 (N_8589,N_8003,N_8291);
nand U8590 (N_8590,N_8498,N_8032);
or U8591 (N_8591,N_8383,N_8104);
nand U8592 (N_8592,N_8224,N_8204);
and U8593 (N_8593,N_8420,N_8491);
or U8594 (N_8594,N_8402,N_8397);
or U8595 (N_8595,N_8083,N_8120);
or U8596 (N_8596,N_8217,N_8367);
xor U8597 (N_8597,N_8184,N_8000);
and U8598 (N_8598,N_8450,N_8340);
xor U8599 (N_8599,N_8100,N_8432);
nor U8600 (N_8600,N_8480,N_8357);
nor U8601 (N_8601,N_8394,N_8462);
xor U8602 (N_8602,N_8088,N_8172);
xor U8603 (N_8603,N_8181,N_8253);
nand U8604 (N_8604,N_8299,N_8493);
or U8605 (N_8605,N_8276,N_8235);
nand U8606 (N_8606,N_8178,N_8098);
nand U8607 (N_8607,N_8429,N_8497);
nor U8608 (N_8608,N_8370,N_8460);
nor U8609 (N_8609,N_8040,N_8486);
nand U8610 (N_8610,N_8288,N_8254);
and U8611 (N_8611,N_8466,N_8223);
and U8612 (N_8612,N_8417,N_8119);
nand U8613 (N_8613,N_8160,N_8142);
nand U8614 (N_8614,N_8162,N_8252);
nand U8615 (N_8615,N_8072,N_8488);
and U8616 (N_8616,N_8458,N_8496);
nor U8617 (N_8617,N_8209,N_8236);
nor U8618 (N_8618,N_8101,N_8360);
and U8619 (N_8619,N_8305,N_8148);
nand U8620 (N_8620,N_8438,N_8301);
or U8621 (N_8621,N_8361,N_8033);
nor U8622 (N_8622,N_8307,N_8176);
or U8623 (N_8623,N_8416,N_8358);
and U8624 (N_8624,N_8492,N_8318);
nor U8625 (N_8625,N_8439,N_8338);
nor U8626 (N_8626,N_8147,N_8435);
nor U8627 (N_8627,N_8423,N_8054);
xnor U8628 (N_8628,N_8258,N_8265);
nand U8629 (N_8629,N_8489,N_8487);
nor U8630 (N_8630,N_8325,N_8455);
and U8631 (N_8631,N_8316,N_8452);
nand U8632 (N_8632,N_8042,N_8335);
or U8633 (N_8633,N_8251,N_8386);
nor U8634 (N_8634,N_8019,N_8282);
nand U8635 (N_8635,N_8479,N_8051);
nand U8636 (N_8636,N_8274,N_8206);
or U8637 (N_8637,N_8377,N_8097);
nor U8638 (N_8638,N_8193,N_8400);
or U8639 (N_8639,N_8222,N_8237);
nand U8640 (N_8640,N_8451,N_8220);
and U8641 (N_8641,N_8315,N_8459);
or U8642 (N_8642,N_8374,N_8401);
or U8643 (N_8643,N_8443,N_8262);
xor U8644 (N_8644,N_8313,N_8164);
nor U8645 (N_8645,N_8186,N_8347);
and U8646 (N_8646,N_8129,N_8110);
and U8647 (N_8647,N_8323,N_8190);
nor U8648 (N_8648,N_8134,N_8195);
and U8649 (N_8649,N_8159,N_8344);
and U8650 (N_8650,N_8478,N_8039);
nand U8651 (N_8651,N_8337,N_8269);
nand U8652 (N_8652,N_8062,N_8464);
nand U8653 (N_8653,N_8339,N_8076);
or U8654 (N_8654,N_8465,N_8481);
nand U8655 (N_8655,N_8297,N_8405);
and U8656 (N_8656,N_8170,N_8107);
and U8657 (N_8657,N_8290,N_8006);
nand U8658 (N_8658,N_8440,N_8073);
nor U8659 (N_8659,N_8068,N_8494);
nor U8660 (N_8660,N_8215,N_8355);
and U8661 (N_8661,N_8132,N_8163);
nor U8662 (N_8662,N_8025,N_8446);
xnor U8663 (N_8663,N_8428,N_8310);
and U8664 (N_8664,N_8395,N_8045);
xor U8665 (N_8665,N_8136,N_8173);
nor U8666 (N_8666,N_8294,N_8391);
and U8667 (N_8667,N_8067,N_8221);
nor U8668 (N_8668,N_8130,N_8208);
nand U8669 (N_8669,N_8017,N_8200);
nor U8670 (N_8670,N_8249,N_8328);
or U8671 (N_8671,N_8375,N_8363);
or U8672 (N_8672,N_8300,N_8049);
nor U8673 (N_8673,N_8449,N_8212);
or U8674 (N_8674,N_8302,N_8289);
xor U8675 (N_8675,N_8201,N_8015);
and U8676 (N_8676,N_8138,N_8431);
and U8677 (N_8677,N_8079,N_8327);
or U8678 (N_8678,N_8131,N_8306);
nor U8679 (N_8679,N_8021,N_8227);
nor U8680 (N_8680,N_8228,N_8424);
and U8681 (N_8681,N_8063,N_8116);
nor U8682 (N_8682,N_8161,N_8112);
and U8683 (N_8683,N_8445,N_8225);
nand U8684 (N_8684,N_8453,N_8263);
nor U8685 (N_8685,N_8177,N_8407);
or U8686 (N_8686,N_8074,N_8388);
nand U8687 (N_8687,N_8158,N_8086);
nand U8688 (N_8688,N_8140,N_8219);
nand U8689 (N_8689,N_8354,N_8117);
and U8690 (N_8690,N_8243,N_8009);
or U8691 (N_8691,N_8050,N_8144);
xor U8692 (N_8692,N_8189,N_8412);
xnor U8693 (N_8693,N_8322,N_8111);
nor U8694 (N_8694,N_8211,N_8232);
and U8695 (N_8695,N_8135,N_8387);
or U8696 (N_8696,N_8371,N_8286);
and U8697 (N_8697,N_8059,N_8382);
nor U8698 (N_8698,N_8092,N_8437);
or U8699 (N_8699,N_8413,N_8026);
xnor U8700 (N_8700,N_8037,N_8454);
xor U8701 (N_8701,N_8191,N_8334);
or U8702 (N_8702,N_8056,N_8156);
or U8703 (N_8703,N_8041,N_8312);
nand U8704 (N_8704,N_8185,N_8474);
nor U8705 (N_8705,N_8238,N_8346);
nor U8706 (N_8706,N_8472,N_8146);
xor U8707 (N_8707,N_8421,N_8279);
nand U8708 (N_8708,N_8356,N_8199);
nor U8709 (N_8709,N_8175,N_8430);
and U8710 (N_8710,N_8389,N_8213);
or U8711 (N_8711,N_8125,N_8272);
or U8712 (N_8712,N_8311,N_8434);
and U8713 (N_8713,N_8053,N_8122);
or U8714 (N_8714,N_8102,N_8183);
and U8715 (N_8715,N_8244,N_8414);
and U8716 (N_8716,N_8364,N_8014);
and U8717 (N_8717,N_8468,N_8174);
nor U8718 (N_8718,N_8013,N_8137);
and U8719 (N_8719,N_8154,N_8150);
xnor U8720 (N_8720,N_8141,N_8020);
nor U8721 (N_8721,N_8392,N_8082);
nor U8722 (N_8722,N_8283,N_8436);
or U8723 (N_8723,N_8277,N_8035);
nand U8724 (N_8724,N_8398,N_8197);
nand U8725 (N_8725,N_8495,N_8089);
xor U8726 (N_8726,N_8319,N_8268);
or U8727 (N_8727,N_8483,N_8210);
and U8728 (N_8728,N_8055,N_8242);
and U8729 (N_8729,N_8168,N_8078);
or U8730 (N_8730,N_8359,N_8095);
and U8731 (N_8731,N_8153,N_8317);
or U8732 (N_8732,N_8266,N_8433);
xor U8733 (N_8733,N_8393,N_8467);
xor U8734 (N_8734,N_8099,N_8461);
and U8735 (N_8735,N_8378,N_8303);
and U8736 (N_8736,N_8124,N_8155);
or U8737 (N_8737,N_8046,N_8149);
xnor U8738 (N_8738,N_8105,N_8425);
xnor U8739 (N_8739,N_8016,N_8246);
nor U8740 (N_8740,N_8447,N_8024);
or U8741 (N_8741,N_8034,N_8010);
nor U8742 (N_8742,N_8157,N_8036);
nand U8743 (N_8743,N_8058,N_8477);
xor U8744 (N_8744,N_8087,N_8341);
and U8745 (N_8745,N_8287,N_8408);
and U8746 (N_8746,N_8329,N_8422);
xor U8747 (N_8747,N_8415,N_8109);
or U8748 (N_8748,N_8348,N_8165);
xnor U8749 (N_8749,N_8384,N_8230);
nand U8750 (N_8750,N_8149,N_8174);
nand U8751 (N_8751,N_8341,N_8145);
or U8752 (N_8752,N_8168,N_8448);
nand U8753 (N_8753,N_8202,N_8254);
or U8754 (N_8754,N_8359,N_8423);
and U8755 (N_8755,N_8077,N_8339);
and U8756 (N_8756,N_8197,N_8434);
xor U8757 (N_8757,N_8184,N_8449);
xnor U8758 (N_8758,N_8117,N_8218);
and U8759 (N_8759,N_8424,N_8387);
nand U8760 (N_8760,N_8092,N_8035);
and U8761 (N_8761,N_8021,N_8160);
nor U8762 (N_8762,N_8289,N_8249);
and U8763 (N_8763,N_8205,N_8273);
nand U8764 (N_8764,N_8013,N_8206);
nor U8765 (N_8765,N_8424,N_8479);
and U8766 (N_8766,N_8404,N_8122);
xnor U8767 (N_8767,N_8377,N_8444);
nand U8768 (N_8768,N_8209,N_8344);
or U8769 (N_8769,N_8404,N_8251);
and U8770 (N_8770,N_8388,N_8465);
nor U8771 (N_8771,N_8053,N_8328);
or U8772 (N_8772,N_8193,N_8124);
nand U8773 (N_8773,N_8463,N_8376);
and U8774 (N_8774,N_8399,N_8213);
xor U8775 (N_8775,N_8152,N_8343);
xnor U8776 (N_8776,N_8387,N_8189);
nor U8777 (N_8777,N_8281,N_8484);
nor U8778 (N_8778,N_8342,N_8303);
or U8779 (N_8779,N_8365,N_8219);
nor U8780 (N_8780,N_8386,N_8162);
and U8781 (N_8781,N_8150,N_8297);
nand U8782 (N_8782,N_8013,N_8058);
nand U8783 (N_8783,N_8043,N_8078);
or U8784 (N_8784,N_8000,N_8214);
nor U8785 (N_8785,N_8120,N_8455);
xor U8786 (N_8786,N_8211,N_8395);
xor U8787 (N_8787,N_8158,N_8117);
and U8788 (N_8788,N_8126,N_8197);
nor U8789 (N_8789,N_8477,N_8049);
nor U8790 (N_8790,N_8367,N_8269);
nor U8791 (N_8791,N_8272,N_8208);
nand U8792 (N_8792,N_8491,N_8387);
nor U8793 (N_8793,N_8170,N_8440);
and U8794 (N_8794,N_8450,N_8310);
nor U8795 (N_8795,N_8096,N_8262);
or U8796 (N_8796,N_8316,N_8165);
nand U8797 (N_8797,N_8480,N_8143);
or U8798 (N_8798,N_8219,N_8047);
nand U8799 (N_8799,N_8320,N_8236);
nor U8800 (N_8800,N_8201,N_8184);
nor U8801 (N_8801,N_8094,N_8011);
or U8802 (N_8802,N_8102,N_8346);
or U8803 (N_8803,N_8050,N_8247);
nor U8804 (N_8804,N_8065,N_8389);
xor U8805 (N_8805,N_8272,N_8050);
and U8806 (N_8806,N_8041,N_8275);
or U8807 (N_8807,N_8047,N_8362);
nand U8808 (N_8808,N_8329,N_8350);
nor U8809 (N_8809,N_8307,N_8136);
xor U8810 (N_8810,N_8410,N_8297);
nor U8811 (N_8811,N_8265,N_8427);
and U8812 (N_8812,N_8241,N_8353);
nand U8813 (N_8813,N_8018,N_8180);
and U8814 (N_8814,N_8312,N_8050);
nor U8815 (N_8815,N_8000,N_8331);
nor U8816 (N_8816,N_8300,N_8444);
or U8817 (N_8817,N_8163,N_8109);
and U8818 (N_8818,N_8327,N_8217);
and U8819 (N_8819,N_8032,N_8256);
and U8820 (N_8820,N_8233,N_8429);
nand U8821 (N_8821,N_8369,N_8497);
or U8822 (N_8822,N_8238,N_8047);
nand U8823 (N_8823,N_8431,N_8418);
nand U8824 (N_8824,N_8475,N_8383);
nor U8825 (N_8825,N_8045,N_8006);
nor U8826 (N_8826,N_8279,N_8114);
and U8827 (N_8827,N_8015,N_8279);
or U8828 (N_8828,N_8353,N_8406);
nor U8829 (N_8829,N_8316,N_8423);
nand U8830 (N_8830,N_8495,N_8257);
and U8831 (N_8831,N_8092,N_8169);
nand U8832 (N_8832,N_8044,N_8189);
nor U8833 (N_8833,N_8157,N_8436);
nor U8834 (N_8834,N_8018,N_8487);
xnor U8835 (N_8835,N_8234,N_8058);
xor U8836 (N_8836,N_8305,N_8427);
or U8837 (N_8837,N_8182,N_8133);
xnor U8838 (N_8838,N_8138,N_8234);
nand U8839 (N_8839,N_8297,N_8035);
nor U8840 (N_8840,N_8327,N_8277);
nand U8841 (N_8841,N_8479,N_8328);
nor U8842 (N_8842,N_8028,N_8155);
nand U8843 (N_8843,N_8386,N_8468);
nand U8844 (N_8844,N_8223,N_8097);
or U8845 (N_8845,N_8402,N_8427);
nand U8846 (N_8846,N_8002,N_8105);
nor U8847 (N_8847,N_8076,N_8230);
nand U8848 (N_8848,N_8498,N_8195);
xnor U8849 (N_8849,N_8153,N_8325);
nand U8850 (N_8850,N_8135,N_8101);
or U8851 (N_8851,N_8189,N_8209);
nor U8852 (N_8852,N_8150,N_8450);
or U8853 (N_8853,N_8337,N_8338);
or U8854 (N_8854,N_8169,N_8393);
nand U8855 (N_8855,N_8145,N_8192);
or U8856 (N_8856,N_8069,N_8011);
xor U8857 (N_8857,N_8008,N_8270);
and U8858 (N_8858,N_8320,N_8186);
and U8859 (N_8859,N_8482,N_8042);
and U8860 (N_8860,N_8421,N_8348);
nor U8861 (N_8861,N_8346,N_8148);
and U8862 (N_8862,N_8110,N_8304);
nand U8863 (N_8863,N_8173,N_8299);
nor U8864 (N_8864,N_8039,N_8197);
or U8865 (N_8865,N_8323,N_8067);
or U8866 (N_8866,N_8264,N_8192);
nand U8867 (N_8867,N_8148,N_8048);
nor U8868 (N_8868,N_8059,N_8498);
nand U8869 (N_8869,N_8066,N_8336);
nand U8870 (N_8870,N_8216,N_8052);
nand U8871 (N_8871,N_8383,N_8201);
nor U8872 (N_8872,N_8293,N_8161);
or U8873 (N_8873,N_8396,N_8460);
nor U8874 (N_8874,N_8448,N_8411);
nor U8875 (N_8875,N_8352,N_8378);
nor U8876 (N_8876,N_8314,N_8368);
or U8877 (N_8877,N_8127,N_8428);
and U8878 (N_8878,N_8313,N_8017);
nand U8879 (N_8879,N_8084,N_8094);
and U8880 (N_8880,N_8488,N_8380);
nor U8881 (N_8881,N_8197,N_8229);
and U8882 (N_8882,N_8339,N_8215);
or U8883 (N_8883,N_8115,N_8078);
or U8884 (N_8884,N_8223,N_8155);
and U8885 (N_8885,N_8135,N_8281);
nor U8886 (N_8886,N_8480,N_8251);
nor U8887 (N_8887,N_8287,N_8032);
or U8888 (N_8888,N_8460,N_8339);
nor U8889 (N_8889,N_8213,N_8124);
or U8890 (N_8890,N_8340,N_8005);
or U8891 (N_8891,N_8101,N_8197);
xnor U8892 (N_8892,N_8377,N_8084);
and U8893 (N_8893,N_8184,N_8439);
nand U8894 (N_8894,N_8442,N_8339);
or U8895 (N_8895,N_8372,N_8158);
xnor U8896 (N_8896,N_8398,N_8163);
and U8897 (N_8897,N_8344,N_8335);
nor U8898 (N_8898,N_8332,N_8300);
xor U8899 (N_8899,N_8234,N_8463);
nor U8900 (N_8900,N_8269,N_8033);
nand U8901 (N_8901,N_8461,N_8003);
xor U8902 (N_8902,N_8121,N_8090);
nor U8903 (N_8903,N_8202,N_8111);
nand U8904 (N_8904,N_8499,N_8025);
nand U8905 (N_8905,N_8342,N_8388);
and U8906 (N_8906,N_8092,N_8281);
or U8907 (N_8907,N_8163,N_8221);
nor U8908 (N_8908,N_8322,N_8271);
and U8909 (N_8909,N_8308,N_8394);
nand U8910 (N_8910,N_8205,N_8487);
nor U8911 (N_8911,N_8423,N_8336);
nand U8912 (N_8912,N_8430,N_8333);
nand U8913 (N_8913,N_8102,N_8187);
nand U8914 (N_8914,N_8390,N_8396);
or U8915 (N_8915,N_8317,N_8089);
xnor U8916 (N_8916,N_8253,N_8238);
nand U8917 (N_8917,N_8117,N_8269);
nor U8918 (N_8918,N_8151,N_8011);
nand U8919 (N_8919,N_8269,N_8111);
nand U8920 (N_8920,N_8344,N_8454);
and U8921 (N_8921,N_8015,N_8273);
nand U8922 (N_8922,N_8404,N_8105);
nor U8923 (N_8923,N_8270,N_8049);
xnor U8924 (N_8924,N_8419,N_8152);
or U8925 (N_8925,N_8475,N_8374);
nand U8926 (N_8926,N_8064,N_8024);
or U8927 (N_8927,N_8490,N_8041);
or U8928 (N_8928,N_8357,N_8053);
nor U8929 (N_8929,N_8359,N_8077);
or U8930 (N_8930,N_8331,N_8066);
and U8931 (N_8931,N_8073,N_8150);
xor U8932 (N_8932,N_8009,N_8029);
and U8933 (N_8933,N_8386,N_8069);
nand U8934 (N_8934,N_8053,N_8214);
nor U8935 (N_8935,N_8146,N_8130);
nand U8936 (N_8936,N_8258,N_8233);
or U8937 (N_8937,N_8467,N_8291);
nand U8938 (N_8938,N_8267,N_8108);
and U8939 (N_8939,N_8348,N_8061);
nor U8940 (N_8940,N_8257,N_8185);
nand U8941 (N_8941,N_8218,N_8173);
and U8942 (N_8942,N_8070,N_8245);
or U8943 (N_8943,N_8119,N_8396);
nor U8944 (N_8944,N_8235,N_8298);
nor U8945 (N_8945,N_8259,N_8080);
xor U8946 (N_8946,N_8382,N_8390);
nor U8947 (N_8947,N_8353,N_8332);
nand U8948 (N_8948,N_8075,N_8402);
nand U8949 (N_8949,N_8007,N_8334);
xnor U8950 (N_8950,N_8366,N_8321);
and U8951 (N_8951,N_8473,N_8153);
nand U8952 (N_8952,N_8024,N_8236);
or U8953 (N_8953,N_8008,N_8498);
nand U8954 (N_8954,N_8104,N_8041);
nor U8955 (N_8955,N_8426,N_8423);
and U8956 (N_8956,N_8492,N_8388);
or U8957 (N_8957,N_8245,N_8000);
and U8958 (N_8958,N_8455,N_8398);
or U8959 (N_8959,N_8380,N_8334);
or U8960 (N_8960,N_8305,N_8131);
nor U8961 (N_8961,N_8378,N_8463);
and U8962 (N_8962,N_8431,N_8043);
and U8963 (N_8963,N_8226,N_8222);
and U8964 (N_8964,N_8070,N_8454);
nand U8965 (N_8965,N_8342,N_8164);
and U8966 (N_8966,N_8175,N_8239);
and U8967 (N_8967,N_8154,N_8290);
nand U8968 (N_8968,N_8166,N_8303);
or U8969 (N_8969,N_8024,N_8105);
and U8970 (N_8970,N_8323,N_8141);
or U8971 (N_8971,N_8396,N_8079);
or U8972 (N_8972,N_8376,N_8159);
and U8973 (N_8973,N_8228,N_8426);
and U8974 (N_8974,N_8330,N_8324);
and U8975 (N_8975,N_8152,N_8115);
nor U8976 (N_8976,N_8110,N_8090);
nand U8977 (N_8977,N_8404,N_8061);
nand U8978 (N_8978,N_8306,N_8168);
or U8979 (N_8979,N_8471,N_8309);
nor U8980 (N_8980,N_8086,N_8383);
xnor U8981 (N_8981,N_8229,N_8321);
or U8982 (N_8982,N_8209,N_8375);
and U8983 (N_8983,N_8464,N_8180);
nand U8984 (N_8984,N_8361,N_8345);
or U8985 (N_8985,N_8188,N_8132);
and U8986 (N_8986,N_8429,N_8074);
or U8987 (N_8987,N_8268,N_8025);
and U8988 (N_8988,N_8419,N_8155);
nor U8989 (N_8989,N_8473,N_8057);
and U8990 (N_8990,N_8436,N_8166);
or U8991 (N_8991,N_8045,N_8397);
nor U8992 (N_8992,N_8046,N_8034);
and U8993 (N_8993,N_8331,N_8424);
or U8994 (N_8994,N_8116,N_8317);
nor U8995 (N_8995,N_8382,N_8070);
and U8996 (N_8996,N_8009,N_8458);
nor U8997 (N_8997,N_8242,N_8115);
nand U8998 (N_8998,N_8405,N_8323);
nand U8999 (N_8999,N_8024,N_8323);
nor U9000 (N_9000,N_8657,N_8864);
and U9001 (N_9001,N_8652,N_8882);
and U9002 (N_9002,N_8526,N_8975);
nand U9003 (N_9003,N_8567,N_8531);
nor U9004 (N_9004,N_8602,N_8649);
or U9005 (N_9005,N_8768,N_8901);
or U9006 (N_9006,N_8769,N_8852);
nor U9007 (N_9007,N_8801,N_8983);
nor U9008 (N_9008,N_8871,N_8723);
and U9009 (N_9009,N_8844,N_8785);
or U9010 (N_9010,N_8937,N_8540);
nand U9011 (N_9011,N_8626,N_8784);
and U9012 (N_9012,N_8790,N_8638);
nand U9013 (N_9013,N_8955,N_8842);
nor U9014 (N_9014,N_8958,N_8881);
or U9015 (N_9015,N_8666,N_8672);
and U9016 (N_9016,N_8906,N_8524);
nand U9017 (N_9017,N_8775,N_8800);
and U9018 (N_9018,N_8551,N_8596);
nand U9019 (N_9019,N_8564,N_8814);
and U9020 (N_9020,N_8591,N_8663);
or U9021 (N_9021,N_8875,N_8577);
or U9022 (N_9022,N_8789,N_8942);
nand U9023 (N_9023,N_8987,N_8770);
nand U9024 (N_9024,N_8588,N_8939);
nand U9025 (N_9025,N_8808,N_8758);
and U9026 (N_9026,N_8890,N_8530);
or U9027 (N_9027,N_8573,N_8945);
nor U9028 (N_9028,N_8587,N_8760);
or U9029 (N_9029,N_8632,N_8609);
xor U9030 (N_9030,N_8959,N_8919);
nand U9031 (N_9031,N_8741,N_8914);
or U9032 (N_9032,N_8651,N_8989);
or U9033 (N_9033,N_8931,N_8645);
xor U9034 (N_9034,N_8988,N_8671);
and U9035 (N_9035,N_8913,N_8675);
or U9036 (N_9036,N_8927,N_8934);
nand U9037 (N_9037,N_8619,N_8970);
nand U9038 (N_9038,N_8971,N_8765);
and U9039 (N_9039,N_8574,N_8678);
nor U9040 (N_9040,N_8992,N_8838);
and U9041 (N_9041,N_8685,N_8973);
xnor U9042 (N_9042,N_8656,N_8745);
or U9043 (N_9043,N_8984,N_8755);
nand U9044 (N_9044,N_8565,N_8583);
or U9045 (N_9045,N_8997,N_8816);
and U9046 (N_9046,N_8905,N_8584);
and U9047 (N_9047,N_8550,N_8534);
and U9048 (N_9048,N_8862,N_8623);
or U9049 (N_9049,N_8729,N_8529);
nor U9050 (N_9050,N_8659,N_8917);
nand U9051 (N_9051,N_8807,N_8582);
nor U9052 (N_9052,N_8654,N_8527);
or U9053 (N_9053,N_8980,N_8507);
or U9054 (N_9054,N_8786,N_8508);
xnor U9055 (N_9055,N_8899,N_8925);
nand U9056 (N_9056,N_8912,N_8521);
or U9057 (N_9057,N_8506,N_8581);
nand U9058 (N_9058,N_8904,N_8689);
xnor U9059 (N_9059,N_8616,N_8764);
nor U9060 (N_9060,N_8606,N_8796);
or U9061 (N_9061,N_8707,N_8859);
and U9062 (N_9062,N_8629,N_8598);
and U9063 (N_9063,N_8819,N_8798);
and U9064 (N_9064,N_8879,N_8885);
nand U9065 (N_9065,N_8886,N_8776);
or U9066 (N_9066,N_8512,N_8818);
or U9067 (N_9067,N_8525,N_8777);
or U9068 (N_9068,N_8727,N_8560);
and U9069 (N_9069,N_8898,N_8722);
or U9070 (N_9070,N_8835,N_8676);
or U9071 (N_9071,N_8738,N_8752);
and U9072 (N_9072,N_8979,N_8806);
and U9073 (N_9073,N_8982,N_8940);
nand U9074 (N_9074,N_8554,N_8909);
xnor U9075 (N_9075,N_8799,N_8668);
and U9076 (N_9076,N_8721,N_8648);
or U9077 (N_9077,N_8921,N_8795);
and U9078 (N_9078,N_8747,N_8993);
nand U9079 (N_9079,N_8624,N_8762);
nand U9080 (N_9080,N_8922,N_8981);
nand U9081 (N_9081,N_8712,N_8545);
or U9082 (N_9082,N_8590,N_8612);
and U9083 (N_9083,N_8968,N_8972);
or U9084 (N_9084,N_8597,N_8604);
nand U9085 (N_9085,N_8586,N_8815);
and U9086 (N_9086,N_8936,N_8757);
nand U9087 (N_9087,N_8620,N_8744);
or U9088 (N_9088,N_8827,N_8846);
nand U9089 (N_9089,N_8687,N_8599);
nor U9090 (N_9090,N_8701,N_8944);
nand U9091 (N_9091,N_8603,N_8860);
nand U9092 (N_9092,N_8613,N_8843);
nor U9093 (N_9093,N_8966,N_8932);
or U9094 (N_9094,N_8566,N_8926);
xor U9095 (N_9095,N_8630,N_8903);
nor U9096 (N_9096,N_8523,N_8547);
nor U9097 (N_9097,N_8878,N_8887);
xnor U9098 (N_9098,N_8924,N_8779);
nor U9099 (N_9099,N_8617,N_8908);
nor U9100 (N_9100,N_8829,N_8684);
xnor U9101 (N_9101,N_8548,N_8642);
and U9102 (N_9102,N_8910,N_8810);
and U9103 (N_9103,N_8643,N_8963);
or U9104 (N_9104,N_8856,N_8888);
and U9105 (N_9105,N_8639,N_8719);
or U9106 (N_9106,N_8711,N_8869);
nand U9107 (N_9107,N_8781,N_8828);
or U9108 (N_9108,N_8873,N_8704);
nor U9109 (N_9109,N_8830,N_8950);
or U9110 (N_9110,N_8509,N_8694);
nand U9111 (N_9111,N_8683,N_8670);
and U9112 (N_9112,N_8715,N_8717);
or U9113 (N_9113,N_8947,N_8953);
xor U9114 (N_9114,N_8977,N_8539);
or U9115 (N_9115,N_8610,N_8870);
and U9116 (N_9116,N_8965,N_8836);
and U9117 (N_9117,N_8802,N_8708);
nand U9118 (N_9118,N_8511,N_8631);
and U9119 (N_9119,N_8528,N_8960);
nand U9120 (N_9120,N_8964,N_8695);
and U9121 (N_9121,N_8740,N_8673);
and U9122 (N_9122,N_8804,N_8991);
or U9123 (N_9123,N_8920,N_8553);
and U9124 (N_9124,N_8823,N_8969);
nor U9125 (N_9125,N_8641,N_8692);
nor U9126 (N_9126,N_8933,N_8505);
and U9127 (N_9127,N_8611,N_8572);
or U9128 (N_9128,N_8621,N_8967);
and U9129 (N_9129,N_8634,N_8763);
nor U9130 (N_9130,N_8995,N_8957);
xnor U9131 (N_9131,N_8848,N_8915);
or U9132 (N_9132,N_8661,N_8883);
or U9133 (N_9133,N_8834,N_8569);
or U9134 (N_9134,N_8739,N_8923);
nand U9135 (N_9135,N_8990,N_8748);
nand U9136 (N_9136,N_8614,N_8794);
or U9137 (N_9137,N_8513,N_8737);
and U9138 (N_9138,N_8767,N_8900);
nor U9139 (N_9139,N_8891,N_8681);
nand U9140 (N_9140,N_8578,N_8674);
nor U9141 (N_9141,N_8976,N_8698);
xnor U9142 (N_9142,N_8749,N_8601);
or U9143 (N_9143,N_8669,N_8532);
or U9144 (N_9144,N_8622,N_8831);
nand U9145 (N_9145,N_8866,N_8691);
or U9146 (N_9146,N_8854,N_8850);
nor U9147 (N_9147,N_8724,N_8974);
and U9148 (N_9148,N_8595,N_8627);
and U9149 (N_9149,N_8771,N_8996);
nand U9150 (N_9150,N_8865,N_8849);
nand U9151 (N_9151,N_8894,N_8742);
nor U9152 (N_9152,N_8504,N_8677);
or U9153 (N_9153,N_8826,N_8877);
or U9154 (N_9154,N_8702,N_8880);
or U9155 (N_9155,N_8787,N_8697);
or U9156 (N_9156,N_8640,N_8935);
nor U9157 (N_9157,N_8985,N_8761);
nor U9158 (N_9158,N_8593,N_8520);
nand U9159 (N_9159,N_8793,N_8733);
and U9160 (N_9160,N_8705,N_8607);
nand U9161 (N_9161,N_8662,N_8930);
nor U9162 (N_9162,N_8517,N_8778);
or U9163 (N_9163,N_8680,N_8699);
xor U9164 (N_9164,N_8952,N_8688);
nor U9165 (N_9165,N_8570,N_8700);
xor U9166 (N_9166,N_8928,N_8946);
nand U9167 (N_9167,N_8501,N_8999);
and U9168 (N_9168,N_8543,N_8876);
nand U9169 (N_9169,N_8813,N_8907);
nand U9170 (N_9170,N_8559,N_8664);
nor U9171 (N_9171,N_8575,N_8867);
or U9172 (N_9172,N_8986,N_8803);
or U9173 (N_9173,N_8825,N_8710);
and U9174 (N_9174,N_8774,N_8874);
or U9175 (N_9175,N_8576,N_8858);
or U9176 (N_9176,N_8897,N_8589);
or U9177 (N_9177,N_8655,N_8792);
and U9178 (N_9178,N_8902,N_8746);
xnor U9179 (N_9179,N_8518,N_8929);
and U9180 (N_9180,N_8556,N_8766);
xnor U9181 (N_9181,N_8962,N_8552);
or U9182 (N_9182,N_8667,N_8500);
and U9183 (N_9183,N_8571,N_8896);
nor U9184 (N_9184,N_8514,N_8658);
nor U9185 (N_9185,N_8994,N_8845);
nand U9186 (N_9186,N_8788,N_8646);
or U9187 (N_9187,N_8743,N_8726);
or U9188 (N_9188,N_8686,N_8943);
nor U9189 (N_9189,N_8868,N_8720);
and U9190 (N_9190,N_8892,N_8718);
or U9191 (N_9191,N_8839,N_8637);
or U9192 (N_9192,N_8773,N_8889);
nor U9193 (N_9193,N_8759,N_8579);
and U9194 (N_9194,N_8951,N_8522);
nand U9195 (N_9195,N_8555,N_8750);
xnor U9196 (N_9196,N_8714,N_8660);
and U9197 (N_9197,N_8633,N_8893);
or U9198 (N_9198,N_8805,N_8948);
and U9199 (N_9199,N_8824,N_8515);
nor U9200 (N_9200,N_8730,N_8644);
xor U9201 (N_9201,N_8561,N_8709);
or U9202 (N_9202,N_8938,N_8585);
nor U9203 (N_9203,N_8562,N_8535);
nand U9204 (N_9204,N_8546,N_8544);
nor U9205 (N_9205,N_8847,N_8812);
and U9206 (N_9206,N_8536,N_8756);
nor U9207 (N_9207,N_8821,N_8533);
nor U9208 (N_9208,N_8822,N_8557);
nor U9209 (N_9209,N_8840,N_8797);
and U9210 (N_9210,N_8780,N_8736);
nor U9211 (N_9211,N_8956,N_8772);
and U9212 (N_9212,N_8911,N_8857);
and U9213 (N_9213,N_8696,N_8665);
nand U9214 (N_9214,N_8592,N_8863);
or U9215 (N_9215,N_8782,N_8538);
nand U9216 (N_9216,N_8884,N_8713);
or U9217 (N_9217,N_8841,N_8600);
nand U9218 (N_9218,N_8519,N_8594);
nand U9219 (N_9219,N_8731,N_8542);
nor U9220 (N_9220,N_8861,N_8791);
nor U9221 (N_9221,N_8941,N_8502);
and U9222 (N_9222,N_8851,N_8820);
and U9223 (N_9223,N_8961,N_8837);
and U9224 (N_9224,N_8809,N_8833);
and U9225 (N_9225,N_8541,N_8735);
and U9226 (N_9226,N_8682,N_8647);
nor U9227 (N_9227,N_8563,N_8537);
nor U9228 (N_9228,N_8725,N_8817);
or U9229 (N_9229,N_8716,N_8706);
nand U9230 (N_9230,N_8605,N_8568);
xor U9231 (N_9231,N_8998,N_8949);
and U9232 (N_9232,N_8728,N_8703);
nand U9233 (N_9233,N_8895,N_8853);
and U9234 (N_9234,N_8732,N_8650);
and U9235 (N_9235,N_8558,N_8549);
xor U9236 (N_9236,N_8811,N_8618);
and U9237 (N_9237,N_8832,N_8734);
nor U9238 (N_9238,N_8918,N_8636);
nand U9239 (N_9239,N_8503,N_8753);
nand U9240 (N_9240,N_8751,N_8625);
xor U9241 (N_9241,N_8608,N_8783);
nor U9242 (N_9242,N_8580,N_8628);
nor U9243 (N_9243,N_8510,N_8679);
nand U9244 (N_9244,N_8754,N_8954);
nand U9245 (N_9245,N_8855,N_8653);
or U9246 (N_9246,N_8916,N_8635);
nand U9247 (N_9247,N_8693,N_8690);
nor U9248 (N_9248,N_8872,N_8615);
nand U9249 (N_9249,N_8978,N_8516);
and U9250 (N_9250,N_8503,N_8646);
nor U9251 (N_9251,N_8724,N_8832);
nor U9252 (N_9252,N_8986,N_8898);
and U9253 (N_9253,N_8505,N_8672);
xor U9254 (N_9254,N_8970,N_8845);
and U9255 (N_9255,N_8761,N_8911);
nor U9256 (N_9256,N_8648,N_8802);
or U9257 (N_9257,N_8504,N_8775);
nor U9258 (N_9258,N_8810,N_8628);
and U9259 (N_9259,N_8882,N_8825);
or U9260 (N_9260,N_8657,N_8814);
or U9261 (N_9261,N_8555,N_8567);
xor U9262 (N_9262,N_8542,N_8951);
or U9263 (N_9263,N_8994,N_8865);
nor U9264 (N_9264,N_8743,N_8783);
or U9265 (N_9265,N_8530,N_8643);
and U9266 (N_9266,N_8821,N_8982);
xnor U9267 (N_9267,N_8531,N_8987);
nor U9268 (N_9268,N_8525,N_8770);
and U9269 (N_9269,N_8921,N_8543);
or U9270 (N_9270,N_8775,N_8729);
or U9271 (N_9271,N_8692,N_8996);
nand U9272 (N_9272,N_8965,N_8650);
or U9273 (N_9273,N_8857,N_8504);
nand U9274 (N_9274,N_8611,N_8646);
nor U9275 (N_9275,N_8789,N_8669);
and U9276 (N_9276,N_8684,N_8513);
nand U9277 (N_9277,N_8521,N_8505);
or U9278 (N_9278,N_8781,N_8821);
xor U9279 (N_9279,N_8736,N_8505);
and U9280 (N_9280,N_8831,N_8503);
and U9281 (N_9281,N_8779,N_8909);
nor U9282 (N_9282,N_8823,N_8624);
nand U9283 (N_9283,N_8896,N_8770);
or U9284 (N_9284,N_8959,N_8748);
and U9285 (N_9285,N_8733,N_8786);
and U9286 (N_9286,N_8937,N_8862);
xor U9287 (N_9287,N_8862,N_8857);
or U9288 (N_9288,N_8532,N_8772);
or U9289 (N_9289,N_8519,N_8792);
or U9290 (N_9290,N_8727,N_8612);
xnor U9291 (N_9291,N_8543,N_8908);
xor U9292 (N_9292,N_8987,N_8941);
nor U9293 (N_9293,N_8649,N_8982);
nand U9294 (N_9294,N_8612,N_8572);
and U9295 (N_9295,N_8659,N_8924);
nand U9296 (N_9296,N_8665,N_8807);
nor U9297 (N_9297,N_8988,N_8849);
xnor U9298 (N_9298,N_8962,N_8988);
nand U9299 (N_9299,N_8540,N_8963);
xor U9300 (N_9300,N_8963,N_8859);
and U9301 (N_9301,N_8671,N_8903);
nor U9302 (N_9302,N_8981,N_8505);
and U9303 (N_9303,N_8645,N_8530);
or U9304 (N_9304,N_8683,N_8585);
nor U9305 (N_9305,N_8737,N_8764);
nand U9306 (N_9306,N_8750,N_8646);
nand U9307 (N_9307,N_8866,N_8845);
nand U9308 (N_9308,N_8704,N_8695);
nand U9309 (N_9309,N_8664,N_8526);
nand U9310 (N_9310,N_8816,N_8744);
and U9311 (N_9311,N_8594,N_8880);
and U9312 (N_9312,N_8673,N_8942);
or U9313 (N_9313,N_8522,N_8996);
and U9314 (N_9314,N_8891,N_8528);
nand U9315 (N_9315,N_8945,N_8926);
or U9316 (N_9316,N_8619,N_8575);
and U9317 (N_9317,N_8758,N_8930);
nand U9318 (N_9318,N_8757,N_8699);
or U9319 (N_9319,N_8754,N_8798);
nor U9320 (N_9320,N_8774,N_8629);
nor U9321 (N_9321,N_8792,N_8654);
and U9322 (N_9322,N_8746,N_8909);
xnor U9323 (N_9323,N_8704,N_8519);
or U9324 (N_9324,N_8782,N_8838);
nor U9325 (N_9325,N_8705,N_8687);
nand U9326 (N_9326,N_8573,N_8533);
and U9327 (N_9327,N_8885,N_8998);
nand U9328 (N_9328,N_8582,N_8640);
and U9329 (N_9329,N_8621,N_8810);
nor U9330 (N_9330,N_8667,N_8955);
or U9331 (N_9331,N_8898,N_8748);
nor U9332 (N_9332,N_8829,N_8552);
or U9333 (N_9333,N_8915,N_8788);
nor U9334 (N_9334,N_8931,N_8697);
nand U9335 (N_9335,N_8650,N_8894);
nand U9336 (N_9336,N_8529,N_8859);
nor U9337 (N_9337,N_8509,N_8727);
nand U9338 (N_9338,N_8697,N_8921);
and U9339 (N_9339,N_8711,N_8633);
nor U9340 (N_9340,N_8884,N_8847);
nand U9341 (N_9341,N_8631,N_8584);
xor U9342 (N_9342,N_8868,N_8546);
xnor U9343 (N_9343,N_8502,N_8983);
and U9344 (N_9344,N_8949,N_8569);
xnor U9345 (N_9345,N_8689,N_8912);
xor U9346 (N_9346,N_8889,N_8684);
nand U9347 (N_9347,N_8985,N_8774);
xnor U9348 (N_9348,N_8792,N_8586);
and U9349 (N_9349,N_8704,N_8894);
or U9350 (N_9350,N_8827,N_8502);
nand U9351 (N_9351,N_8913,N_8845);
and U9352 (N_9352,N_8728,N_8697);
or U9353 (N_9353,N_8604,N_8510);
or U9354 (N_9354,N_8622,N_8522);
xnor U9355 (N_9355,N_8941,N_8692);
nand U9356 (N_9356,N_8508,N_8886);
nand U9357 (N_9357,N_8651,N_8862);
nand U9358 (N_9358,N_8848,N_8666);
and U9359 (N_9359,N_8711,N_8570);
or U9360 (N_9360,N_8845,N_8719);
nor U9361 (N_9361,N_8514,N_8673);
or U9362 (N_9362,N_8987,N_8669);
nand U9363 (N_9363,N_8541,N_8974);
nand U9364 (N_9364,N_8891,N_8762);
nor U9365 (N_9365,N_8871,N_8517);
xor U9366 (N_9366,N_8885,N_8843);
or U9367 (N_9367,N_8724,N_8532);
nor U9368 (N_9368,N_8546,N_8980);
and U9369 (N_9369,N_8679,N_8507);
nor U9370 (N_9370,N_8965,N_8562);
and U9371 (N_9371,N_8922,N_8858);
nand U9372 (N_9372,N_8980,N_8611);
xnor U9373 (N_9373,N_8643,N_8793);
nor U9374 (N_9374,N_8888,N_8523);
and U9375 (N_9375,N_8706,N_8932);
nand U9376 (N_9376,N_8764,N_8595);
and U9377 (N_9377,N_8704,N_8988);
nor U9378 (N_9378,N_8600,N_8650);
nor U9379 (N_9379,N_8876,N_8853);
nand U9380 (N_9380,N_8715,N_8961);
and U9381 (N_9381,N_8984,N_8962);
nor U9382 (N_9382,N_8863,N_8848);
nand U9383 (N_9383,N_8705,N_8690);
nor U9384 (N_9384,N_8517,N_8866);
nor U9385 (N_9385,N_8874,N_8960);
nand U9386 (N_9386,N_8563,N_8875);
nor U9387 (N_9387,N_8923,N_8858);
nor U9388 (N_9388,N_8580,N_8733);
or U9389 (N_9389,N_8564,N_8692);
and U9390 (N_9390,N_8823,N_8934);
nor U9391 (N_9391,N_8542,N_8632);
nand U9392 (N_9392,N_8713,N_8628);
or U9393 (N_9393,N_8833,N_8722);
and U9394 (N_9394,N_8694,N_8766);
nor U9395 (N_9395,N_8671,N_8719);
nand U9396 (N_9396,N_8561,N_8864);
nor U9397 (N_9397,N_8558,N_8625);
or U9398 (N_9398,N_8615,N_8739);
and U9399 (N_9399,N_8916,N_8642);
nand U9400 (N_9400,N_8984,N_8774);
nand U9401 (N_9401,N_8639,N_8527);
nand U9402 (N_9402,N_8675,N_8537);
nor U9403 (N_9403,N_8993,N_8521);
and U9404 (N_9404,N_8900,N_8844);
or U9405 (N_9405,N_8793,N_8591);
nor U9406 (N_9406,N_8994,N_8656);
and U9407 (N_9407,N_8674,N_8677);
and U9408 (N_9408,N_8987,N_8837);
nand U9409 (N_9409,N_8685,N_8825);
or U9410 (N_9410,N_8502,N_8930);
nand U9411 (N_9411,N_8739,N_8526);
nor U9412 (N_9412,N_8508,N_8632);
xor U9413 (N_9413,N_8985,N_8757);
xnor U9414 (N_9414,N_8655,N_8878);
nor U9415 (N_9415,N_8516,N_8592);
and U9416 (N_9416,N_8871,N_8778);
and U9417 (N_9417,N_8585,N_8803);
and U9418 (N_9418,N_8623,N_8739);
and U9419 (N_9419,N_8554,N_8810);
xnor U9420 (N_9420,N_8952,N_8687);
nor U9421 (N_9421,N_8754,N_8625);
xor U9422 (N_9422,N_8656,N_8603);
or U9423 (N_9423,N_8874,N_8615);
or U9424 (N_9424,N_8742,N_8820);
nand U9425 (N_9425,N_8893,N_8533);
nor U9426 (N_9426,N_8728,N_8972);
nand U9427 (N_9427,N_8802,N_8899);
or U9428 (N_9428,N_8729,N_8870);
nand U9429 (N_9429,N_8683,N_8693);
or U9430 (N_9430,N_8990,N_8649);
nand U9431 (N_9431,N_8726,N_8731);
or U9432 (N_9432,N_8625,N_8680);
nand U9433 (N_9433,N_8746,N_8784);
or U9434 (N_9434,N_8818,N_8622);
and U9435 (N_9435,N_8635,N_8922);
or U9436 (N_9436,N_8683,N_8956);
nand U9437 (N_9437,N_8785,N_8845);
nor U9438 (N_9438,N_8643,N_8555);
nor U9439 (N_9439,N_8791,N_8545);
xor U9440 (N_9440,N_8608,N_8771);
or U9441 (N_9441,N_8928,N_8613);
or U9442 (N_9442,N_8920,N_8883);
or U9443 (N_9443,N_8911,N_8803);
nor U9444 (N_9444,N_8590,N_8755);
nand U9445 (N_9445,N_8746,N_8911);
or U9446 (N_9446,N_8771,N_8509);
nor U9447 (N_9447,N_8845,N_8805);
and U9448 (N_9448,N_8821,N_8532);
nand U9449 (N_9449,N_8754,N_8731);
and U9450 (N_9450,N_8674,N_8834);
nor U9451 (N_9451,N_8521,N_8634);
nand U9452 (N_9452,N_8623,N_8958);
or U9453 (N_9453,N_8504,N_8608);
nand U9454 (N_9454,N_8629,N_8554);
xnor U9455 (N_9455,N_8869,N_8596);
nor U9456 (N_9456,N_8653,N_8720);
xor U9457 (N_9457,N_8600,N_8511);
and U9458 (N_9458,N_8961,N_8943);
or U9459 (N_9459,N_8908,N_8804);
nand U9460 (N_9460,N_8533,N_8840);
nand U9461 (N_9461,N_8671,N_8579);
xnor U9462 (N_9462,N_8591,N_8945);
and U9463 (N_9463,N_8829,N_8702);
nor U9464 (N_9464,N_8733,N_8716);
nor U9465 (N_9465,N_8922,N_8703);
and U9466 (N_9466,N_8788,N_8536);
nor U9467 (N_9467,N_8619,N_8516);
or U9468 (N_9468,N_8758,N_8826);
or U9469 (N_9469,N_8885,N_8897);
nand U9470 (N_9470,N_8621,N_8539);
nand U9471 (N_9471,N_8939,N_8786);
or U9472 (N_9472,N_8747,N_8590);
and U9473 (N_9473,N_8847,N_8795);
and U9474 (N_9474,N_8710,N_8560);
nor U9475 (N_9475,N_8578,N_8782);
nand U9476 (N_9476,N_8966,N_8541);
nor U9477 (N_9477,N_8607,N_8553);
nor U9478 (N_9478,N_8783,N_8850);
or U9479 (N_9479,N_8588,N_8915);
xnor U9480 (N_9480,N_8865,N_8841);
nand U9481 (N_9481,N_8816,N_8711);
and U9482 (N_9482,N_8953,N_8750);
nand U9483 (N_9483,N_8687,N_8690);
or U9484 (N_9484,N_8982,N_8535);
nand U9485 (N_9485,N_8701,N_8677);
xor U9486 (N_9486,N_8736,N_8806);
nand U9487 (N_9487,N_8738,N_8937);
and U9488 (N_9488,N_8633,N_8797);
and U9489 (N_9489,N_8843,N_8593);
xnor U9490 (N_9490,N_8570,N_8854);
nor U9491 (N_9491,N_8600,N_8918);
nor U9492 (N_9492,N_8813,N_8625);
nand U9493 (N_9493,N_8989,N_8672);
or U9494 (N_9494,N_8918,N_8797);
and U9495 (N_9495,N_8838,N_8798);
nand U9496 (N_9496,N_8822,N_8842);
or U9497 (N_9497,N_8651,N_8767);
or U9498 (N_9498,N_8852,N_8951);
and U9499 (N_9499,N_8965,N_8934);
xor U9500 (N_9500,N_9039,N_9332);
or U9501 (N_9501,N_9494,N_9230);
nand U9502 (N_9502,N_9471,N_9477);
nand U9503 (N_9503,N_9236,N_9265);
nor U9504 (N_9504,N_9475,N_9330);
nand U9505 (N_9505,N_9358,N_9211);
or U9506 (N_9506,N_9322,N_9003);
xor U9507 (N_9507,N_9185,N_9337);
and U9508 (N_9508,N_9262,N_9142);
or U9509 (N_9509,N_9239,N_9267);
nor U9510 (N_9510,N_9270,N_9361);
or U9511 (N_9511,N_9086,N_9227);
nand U9512 (N_9512,N_9394,N_9010);
and U9513 (N_9513,N_9282,N_9049);
and U9514 (N_9514,N_9410,N_9149);
xor U9515 (N_9515,N_9338,N_9373);
nor U9516 (N_9516,N_9176,N_9177);
and U9517 (N_9517,N_9382,N_9045);
nand U9518 (N_9518,N_9229,N_9492);
and U9519 (N_9519,N_9150,N_9452);
or U9520 (N_9520,N_9459,N_9392);
or U9521 (N_9521,N_9388,N_9480);
and U9522 (N_9522,N_9159,N_9179);
xnor U9523 (N_9523,N_9481,N_9071);
nand U9524 (N_9524,N_9024,N_9387);
xnor U9525 (N_9525,N_9339,N_9449);
xor U9526 (N_9526,N_9155,N_9428);
nor U9527 (N_9527,N_9138,N_9034);
and U9528 (N_9528,N_9276,N_9136);
xor U9529 (N_9529,N_9425,N_9336);
and U9530 (N_9530,N_9146,N_9303);
and U9531 (N_9531,N_9088,N_9264);
nor U9532 (N_9532,N_9334,N_9020);
nand U9533 (N_9533,N_9117,N_9404);
nand U9534 (N_9534,N_9467,N_9061);
nor U9535 (N_9535,N_9367,N_9040);
or U9536 (N_9536,N_9285,N_9160);
and U9537 (N_9537,N_9363,N_9172);
nor U9538 (N_9538,N_9105,N_9310);
and U9539 (N_9539,N_9209,N_9257);
xor U9540 (N_9540,N_9067,N_9495);
or U9541 (N_9541,N_9309,N_9151);
or U9542 (N_9542,N_9198,N_9068);
or U9543 (N_9543,N_9346,N_9043);
and U9544 (N_9544,N_9140,N_9390);
xnor U9545 (N_9545,N_9318,N_9087);
and U9546 (N_9546,N_9197,N_9401);
nor U9547 (N_9547,N_9201,N_9167);
and U9548 (N_9548,N_9275,N_9121);
or U9549 (N_9549,N_9395,N_9203);
nor U9550 (N_9550,N_9094,N_9238);
nor U9551 (N_9551,N_9462,N_9396);
nor U9552 (N_9552,N_9059,N_9228);
or U9553 (N_9553,N_9375,N_9080);
nand U9554 (N_9554,N_9496,N_9165);
or U9555 (N_9555,N_9497,N_9370);
xnor U9556 (N_9556,N_9108,N_9162);
and U9557 (N_9557,N_9362,N_9103);
or U9558 (N_9558,N_9443,N_9408);
xnor U9559 (N_9559,N_9397,N_9488);
or U9560 (N_9560,N_9182,N_9189);
nor U9561 (N_9561,N_9109,N_9082);
nand U9562 (N_9562,N_9391,N_9299);
or U9563 (N_9563,N_9154,N_9125);
and U9564 (N_9564,N_9127,N_9400);
and U9565 (N_9565,N_9261,N_9000);
or U9566 (N_9566,N_9491,N_9307);
or U9567 (N_9567,N_9356,N_9118);
nor U9568 (N_9568,N_9412,N_9453);
or U9569 (N_9569,N_9269,N_9335);
and U9570 (N_9570,N_9419,N_9123);
nand U9571 (N_9571,N_9450,N_9217);
xor U9572 (N_9572,N_9207,N_9403);
nor U9573 (N_9573,N_9323,N_9406);
or U9574 (N_9574,N_9178,N_9381);
nand U9575 (N_9575,N_9472,N_9208);
nand U9576 (N_9576,N_9025,N_9240);
or U9577 (N_9577,N_9035,N_9430);
xnor U9578 (N_9578,N_9432,N_9305);
or U9579 (N_9579,N_9026,N_9004);
xnor U9580 (N_9580,N_9325,N_9484);
nand U9581 (N_9581,N_9101,N_9316);
nor U9582 (N_9582,N_9251,N_9078);
nor U9583 (N_9583,N_9458,N_9005);
or U9584 (N_9584,N_9090,N_9083);
or U9585 (N_9585,N_9456,N_9050);
nand U9586 (N_9586,N_9427,N_9487);
and U9587 (N_9587,N_9205,N_9313);
and U9588 (N_9588,N_9327,N_9292);
nand U9589 (N_9589,N_9306,N_9181);
and U9590 (N_9590,N_9417,N_9107);
or U9591 (N_9591,N_9393,N_9196);
or U9592 (N_9592,N_9097,N_9170);
or U9593 (N_9593,N_9037,N_9455);
or U9594 (N_9594,N_9290,N_9293);
or U9595 (N_9595,N_9161,N_9187);
xor U9596 (N_9596,N_9438,N_9032);
nand U9597 (N_9597,N_9143,N_9435);
or U9598 (N_9598,N_9231,N_9468);
nor U9599 (N_9599,N_9463,N_9277);
nand U9600 (N_9600,N_9242,N_9175);
and U9601 (N_9601,N_9399,N_9225);
nor U9602 (N_9602,N_9402,N_9280);
nand U9603 (N_9603,N_9232,N_9469);
nor U9604 (N_9604,N_9499,N_9365);
xnor U9605 (N_9605,N_9411,N_9111);
and U9606 (N_9606,N_9352,N_9145);
nand U9607 (N_9607,N_9465,N_9156);
nor U9608 (N_9608,N_9204,N_9206);
nor U9609 (N_9609,N_9131,N_9429);
or U9610 (N_9610,N_9355,N_9116);
nor U9611 (N_9611,N_9442,N_9298);
and U9612 (N_9612,N_9055,N_9038);
nor U9613 (N_9613,N_9321,N_9194);
nand U9614 (N_9614,N_9283,N_9173);
and U9615 (N_9615,N_9398,N_9058);
xnor U9616 (N_9616,N_9011,N_9461);
nor U9617 (N_9617,N_9202,N_9188);
xnor U9618 (N_9618,N_9268,N_9376);
or U9619 (N_9619,N_9247,N_9389);
nand U9620 (N_9620,N_9106,N_9021);
and U9621 (N_9621,N_9072,N_9098);
or U9622 (N_9622,N_9183,N_9315);
xor U9623 (N_9623,N_9027,N_9493);
nor U9624 (N_9624,N_9056,N_9057);
or U9625 (N_9625,N_9420,N_9424);
nor U9626 (N_9626,N_9383,N_9371);
and U9627 (N_9627,N_9148,N_9431);
nand U9628 (N_9628,N_9126,N_9139);
and U9629 (N_9629,N_9129,N_9446);
and U9630 (N_9630,N_9384,N_9485);
nand U9631 (N_9631,N_9368,N_9498);
xor U9632 (N_9632,N_9284,N_9213);
nand U9633 (N_9633,N_9234,N_9448);
nor U9634 (N_9634,N_9447,N_9163);
nand U9635 (N_9635,N_9437,N_9253);
or U9636 (N_9636,N_9222,N_9066);
and U9637 (N_9637,N_9184,N_9200);
or U9638 (N_9638,N_9483,N_9444);
and U9639 (N_9639,N_9278,N_9304);
nor U9640 (N_9640,N_9019,N_9244);
nor U9641 (N_9641,N_9351,N_9343);
nand U9642 (N_9642,N_9291,N_9281);
nor U9643 (N_9643,N_9100,N_9302);
and U9644 (N_9644,N_9379,N_9342);
nand U9645 (N_9645,N_9147,N_9122);
or U9646 (N_9646,N_9296,N_9054);
nand U9647 (N_9647,N_9135,N_9099);
and U9648 (N_9648,N_9348,N_9454);
xnor U9649 (N_9649,N_9297,N_9473);
and U9650 (N_9650,N_9013,N_9490);
or U9651 (N_9651,N_9445,N_9044);
nand U9652 (N_9652,N_9295,N_9120);
nand U9653 (N_9653,N_9423,N_9434);
or U9654 (N_9654,N_9091,N_9354);
xnor U9655 (N_9655,N_9360,N_9065);
and U9656 (N_9656,N_9036,N_9333);
and U9657 (N_9657,N_9474,N_9312);
xnor U9658 (N_9658,N_9357,N_9029);
nor U9659 (N_9659,N_9093,N_9418);
and U9660 (N_9660,N_9349,N_9215);
and U9661 (N_9661,N_9137,N_9069);
and U9662 (N_9662,N_9457,N_9124);
nor U9663 (N_9663,N_9079,N_9128);
nor U9664 (N_9664,N_9254,N_9060);
and U9665 (N_9665,N_9002,N_9110);
xnor U9666 (N_9666,N_9252,N_9369);
and U9667 (N_9667,N_9018,N_9074);
or U9668 (N_9668,N_9152,N_9378);
and U9669 (N_9669,N_9405,N_9214);
nor U9670 (N_9670,N_9219,N_9130);
xnor U9671 (N_9671,N_9216,N_9256);
nor U9672 (N_9672,N_9301,N_9479);
or U9673 (N_9673,N_9451,N_9171);
nor U9674 (N_9674,N_9246,N_9377);
nor U9675 (N_9675,N_9077,N_9350);
and U9676 (N_9676,N_9364,N_9063);
xnor U9677 (N_9677,N_9241,N_9133);
nor U9678 (N_9678,N_9324,N_9075);
nor U9679 (N_9679,N_9180,N_9046);
nand U9680 (N_9680,N_9199,N_9289);
nand U9681 (N_9681,N_9112,N_9266);
nor U9682 (N_9682,N_9115,N_9274);
or U9683 (N_9683,N_9248,N_9144);
and U9684 (N_9684,N_9329,N_9288);
or U9685 (N_9685,N_9192,N_9092);
nor U9686 (N_9686,N_9314,N_9191);
nor U9687 (N_9687,N_9053,N_9051);
and U9688 (N_9688,N_9070,N_9157);
nor U9689 (N_9689,N_9073,N_9001);
and U9690 (N_9690,N_9353,N_9081);
and U9691 (N_9691,N_9102,N_9320);
and U9692 (N_9692,N_9153,N_9460);
nand U9693 (N_9693,N_9440,N_9028);
nor U9694 (N_9694,N_9042,N_9441);
nor U9695 (N_9695,N_9015,N_9195);
xnor U9696 (N_9696,N_9317,N_9439);
nand U9697 (N_9697,N_9014,N_9486);
nor U9698 (N_9698,N_9260,N_9210);
or U9699 (N_9699,N_9052,N_9319);
or U9700 (N_9700,N_9344,N_9223);
nand U9701 (N_9701,N_9212,N_9466);
or U9702 (N_9702,N_9012,N_9031);
nor U9703 (N_9703,N_9249,N_9258);
xor U9704 (N_9704,N_9478,N_9235);
or U9705 (N_9705,N_9385,N_9273);
xnor U9706 (N_9706,N_9114,N_9030);
and U9707 (N_9707,N_9017,N_9263);
nand U9708 (N_9708,N_9008,N_9006);
or U9709 (N_9709,N_9407,N_9164);
nor U9710 (N_9710,N_9422,N_9169);
nor U9711 (N_9711,N_9007,N_9476);
and U9712 (N_9712,N_9464,N_9416);
nand U9713 (N_9713,N_9374,N_9237);
and U9714 (N_9714,N_9096,N_9166);
nand U9715 (N_9715,N_9433,N_9250);
nand U9716 (N_9716,N_9345,N_9326);
xor U9717 (N_9717,N_9016,N_9119);
nor U9718 (N_9718,N_9064,N_9347);
or U9719 (N_9719,N_9372,N_9186);
or U9720 (N_9720,N_9141,N_9409);
or U9721 (N_9721,N_9272,N_9294);
nor U9722 (N_9722,N_9041,N_9023);
nor U9723 (N_9723,N_9009,N_9413);
nand U9724 (N_9724,N_9089,N_9287);
nor U9725 (N_9725,N_9168,N_9255);
nor U9726 (N_9726,N_9436,N_9193);
or U9727 (N_9727,N_9113,N_9489);
or U9728 (N_9728,N_9233,N_9414);
and U9729 (N_9729,N_9328,N_9259);
and U9730 (N_9730,N_9386,N_9243);
or U9731 (N_9731,N_9085,N_9415);
nor U9732 (N_9732,N_9095,N_9104);
xor U9733 (N_9733,N_9340,N_9359);
or U9734 (N_9734,N_9341,N_9311);
or U9735 (N_9735,N_9470,N_9271);
nor U9736 (N_9736,N_9190,N_9380);
and U9737 (N_9737,N_9286,N_9048);
nand U9738 (N_9738,N_9076,N_9221);
nand U9739 (N_9739,N_9421,N_9174);
and U9740 (N_9740,N_9482,N_9218);
nor U9741 (N_9741,N_9224,N_9220);
and U9742 (N_9742,N_9426,N_9062);
and U9743 (N_9743,N_9308,N_9226);
nand U9744 (N_9744,N_9279,N_9132);
nand U9745 (N_9745,N_9033,N_9331);
or U9746 (N_9746,N_9022,N_9245);
nand U9747 (N_9747,N_9158,N_9084);
nand U9748 (N_9748,N_9366,N_9134);
nor U9749 (N_9749,N_9047,N_9300);
and U9750 (N_9750,N_9066,N_9478);
or U9751 (N_9751,N_9284,N_9110);
nand U9752 (N_9752,N_9132,N_9037);
xor U9753 (N_9753,N_9254,N_9117);
and U9754 (N_9754,N_9404,N_9308);
and U9755 (N_9755,N_9131,N_9172);
xor U9756 (N_9756,N_9015,N_9275);
nand U9757 (N_9757,N_9361,N_9183);
nor U9758 (N_9758,N_9280,N_9102);
nor U9759 (N_9759,N_9099,N_9351);
or U9760 (N_9760,N_9210,N_9202);
nand U9761 (N_9761,N_9148,N_9001);
nand U9762 (N_9762,N_9247,N_9430);
nand U9763 (N_9763,N_9017,N_9387);
or U9764 (N_9764,N_9067,N_9003);
or U9765 (N_9765,N_9116,N_9138);
nor U9766 (N_9766,N_9282,N_9135);
or U9767 (N_9767,N_9498,N_9274);
and U9768 (N_9768,N_9045,N_9374);
nand U9769 (N_9769,N_9002,N_9204);
or U9770 (N_9770,N_9274,N_9411);
or U9771 (N_9771,N_9271,N_9299);
nor U9772 (N_9772,N_9403,N_9321);
nand U9773 (N_9773,N_9032,N_9419);
nand U9774 (N_9774,N_9322,N_9012);
and U9775 (N_9775,N_9489,N_9187);
or U9776 (N_9776,N_9281,N_9243);
or U9777 (N_9777,N_9362,N_9093);
xor U9778 (N_9778,N_9411,N_9150);
xor U9779 (N_9779,N_9488,N_9440);
nor U9780 (N_9780,N_9209,N_9491);
xnor U9781 (N_9781,N_9275,N_9429);
or U9782 (N_9782,N_9487,N_9401);
xnor U9783 (N_9783,N_9409,N_9183);
or U9784 (N_9784,N_9117,N_9024);
nor U9785 (N_9785,N_9479,N_9404);
and U9786 (N_9786,N_9111,N_9142);
nor U9787 (N_9787,N_9257,N_9035);
xnor U9788 (N_9788,N_9361,N_9201);
nor U9789 (N_9789,N_9290,N_9033);
or U9790 (N_9790,N_9042,N_9185);
and U9791 (N_9791,N_9459,N_9298);
xor U9792 (N_9792,N_9403,N_9220);
nand U9793 (N_9793,N_9385,N_9051);
nor U9794 (N_9794,N_9307,N_9488);
nand U9795 (N_9795,N_9093,N_9060);
and U9796 (N_9796,N_9381,N_9188);
nand U9797 (N_9797,N_9249,N_9184);
nand U9798 (N_9798,N_9057,N_9261);
nor U9799 (N_9799,N_9453,N_9296);
and U9800 (N_9800,N_9275,N_9101);
or U9801 (N_9801,N_9358,N_9128);
or U9802 (N_9802,N_9129,N_9005);
nor U9803 (N_9803,N_9462,N_9291);
or U9804 (N_9804,N_9282,N_9294);
nor U9805 (N_9805,N_9283,N_9353);
and U9806 (N_9806,N_9076,N_9265);
or U9807 (N_9807,N_9136,N_9271);
or U9808 (N_9808,N_9323,N_9207);
and U9809 (N_9809,N_9183,N_9241);
nand U9810 (N_9810,N_9471,N_9299);
nand U9811 (N_9811,N_9394,N_9108);
or U9812 (N_9812,N_9340,N_9442);
nor U9813 (N_9813,N_9138,N_9486);
or U9814 (N_9814,N_9152,N_9086);
nor U9815 (N_9815,N_9432,N_9402);
or U9816 (N_9816,N_9282,N_9315);
nor U9817 (N_9817,N_9207,N_9099);
nand U9818 (N_9818,N_9364,N_9469);
nand U9819 (N_9819,N_9425,N_9337);
and U9820 (N_9820,N_9324,N_9416);
nand U9821 (N_9821,N_9069,N_9314);
xor U9822 (N_9822,N_9176,N_9350);
and U9823 (N_9823,N_9056,N_9304);
xnor U9824 (N_9824,N_9380,N_9489);
xor U9825 (N_9825,N_9162,N_9085);
xor U9826 (N_9826,N_9060,N_9353);
xor U9827 (N_9827,N_9461,N_9163);
nand U9828 (N_9828,N_9387,N_9088);
or U9829 (N_9829,N_9331,N_9112);
and U9830 (N_9830,N_9210,N_9137);
or U9831 (N_9831,N_9274,N_9192);
nor U9832 (N_9832,N_9177,N_9494);
nor U9833 (N_9833,N_9414,N_9023);
or U9834 (N_9834,N_9228,N_9208);
nor U9835 (N_9835,N_9312,N_9135);
or U9836 (N_9836,N_9214,N_9406);
nand U9837 (N_9837,N_9460,N_9304);
or U9838 (N_9838,N_9047,N_9493);
and U9839 (N_9839,N_9373,N_9352);
or U9840 (N_9840,N_9218,N_9380);
nor U9841 (N_9841,N_9417,N_9284);
or U9842 (N_9842,N_9447,N_9219);
nand U9843 (N_9843,N_9006,N_9499);
and U9844 (N_9844,N_9136,N_9132);
nand U9845 (N_9845,N_9339,N_9448);
and U9846 (N_9846,N_9083,N_9324);
and U9847 (N_9847,N_9461,N_9167);
or U9848 (N_9848,N_9413,N_9481);
and U9849 (N_9849,N_9153,N_9047);
nor U9850 (N_9850,N_9389,N_9126);
nand U9851 (N_9851,N_9192,N_9199);
and U9852 (N_9852,N_9268,N_9454);
nand U9853 (N_9853,N_9079,N_9199);
or U9854 (N_9854,N_9161,N_9168);
or U9855 (N_9855,N_9411,N_9139);
nor U9856 (N_9856,N_9388,N_9497);
xnor U9857 (N_9857,N_9403,N_9423);
and U9858 (N_9858,N_9123,N_9273);
nor U9859 (N_9859,N_9417,N_9027);
or U9860 (N_9860,N_9176,N_9340);
and U9861 (N_9861,N_9152,N_9104);
or U9862 (N_9862,N_9440,N_9206);
or U9863 (N_9863,N_9065,N_9084);
nand U9864 (N_9864,N_9413,N_9181);
and U9865 (N_9865,N_9144,N_9391);
nor U9866 (N_9866,N_9418,N_9174);
nand U9867 (N_9867,N_9328,N_9332);
or U9868 (N_9868,N_9232,N_9348);
xor U9869 (N_9869,N_9465,N_9280);
nor U9870 (N_9870,N_9063,N_9144);
nor U9871 (N_9871,N_9172,N_9352);
xor U9872 (N_9872,N_9137,N_9163);
nor U9873 (N_9873,N_9217,N_9002);
nand U9874 (N_9874,N_9194,N_9170);
nor U9875 (N_9875,N_9266,N_9486);
or U9876 (N_9876,N_9101,N_9453);
nor U9877 (N_9877,N_9408,N_9469);
or U9878 (N_9878,N_9149,N_9283);
nand U9879 (N_9879,N_9115,N_9406);
and U9880 (N_9880,N_9458,N_9070);
nor U9881 (N_9881,N_9427,N_9328);
nor U9882 (N_9882,N_9210,N_9204);
nand U9883 (N_9883,N_9004,N_9481);
and U9884 (N_9884,N_9265,N_9029);
and U9885 (N_9885,N_9012,N_9356);
or U9886 (N_9886,N_9287,N_9327);
or U9887 (N_9887,N_9247,N_9444);
nor U9888 (N_9888,N_9048,N_9155);
nand U9889 (N_9889,N_9086,N_9455);
and U9890 (N_9890,N_9450,N_9386);
nand U9891 (N_9891,N_9411,N_9043);
nor U9892 (N_9892,N_9097,N_9328);
or U9893 (N_9893,N_9264,N_9114);
xnor U9894 (N_9894,N_9033,N_9286);
or U9895 (N_9895,N_9461,N_9050);
xnor U9896 (N_9896,N_9265,N_9077);
nor U9897 (N_9897,N_9236,N_9302);
nor U9898 (N_9898,N_9404,N_9030);
and U9899 (N_9899,N_9405,N_9437);
xnor U9900 (N_9900,N_9460,N_9284);
nand U9901 (N_9901,N_9228,N_9118);
nand U9902 (N_9902,N_9010,N_9183);
and U9903 (N_9903,N_9179,N_9113);
or U9904 (N_9904,N_9031,N_9120);
nand U9905 (N_9905,N_9445,N_9286);
xor U9906 (N_9906,N_9194,N_9153);
xor U9907 (N_9907,N_9484,N_9167);
and U9908 (N_9908,N_9244,N_9210);
nand U9909 (N_9909,N_9380,N_9142);
xnor U9910 (N_9910,N_9392,N_9174);
or U9911 (N_9911,N_9395,N_9001);
nand U9912 (N_9912,N_9058,N_9393);
nor U9913 (N_9913,N_9302,N_9438);
or U9914 (N_9914,N_9349,N_9310);
or U9915 (N_9915,N_9424,N_9301);
nor U9916 (N_9916,N_9207,N_9186);
nand U9917 (N_9917,N_9095,N_9371);
or U9918 (N_9918,N_9071,N_9284);
and U9919 (N_9919,N_9010,N_9005);
nor U9920 (N_9920,N_9492,N_9485);
or U9921 (N_9921,N_9466,N_9493);
or U9922 (N_9922,N_9457,N_9213);
xnor U9923 (N_9923,N_9017,N_9170);
nand U9924 (N_9924,N_9228,N_9241);
nand U9925 (N_9925,N_9142,N_9088);
nand U9926 (N_9926,N_9008,N_9120);
nor U9927 (N_9927,N_9129,N_9488);
and U9928 (N_9928,N_9476,N_9159);
xor U9929 (N_9929,N_9008,N_9150);
nor U9930 (N_9930,N_9194,N_9179);
or U9931 (N_9931,N_9172,N_9480);
nand U9932 (N_9932,N_9002,N_9361);
or U9933 (N_9933,N_9175,N_9271);
xor U9934 (N_9934,N_9119,N_9267);
and U9935 (N_9935,N_9232,N_9202);
nand U9936 (N_9936,N_9019,N_9148);
nor U9937 (N_9937,N_9346,N_9428);
nand U9938 (N_9938,N_9287,N_9102);
nand U9939 (N_9939,N_9456,N_9093);
and U9940 (N_9940,N_9027,N_9380);
or U9941 (N_9941,N_9065,N_9223);
xnor U9942 (N_9942,N_9362,N_9455);
nand U9943 (N_9943,N_9039,N_9003);
nor U9944 (N_9944,N_9114,N_9454);
or U9945 (N_9945,N_9225,N_9344);
nand U9946 (N_9946,N_9295,N_9417);
nor U9947 (N_9947,N_9232,N_9425);
nand U9948 (N_9948,N_9006,N_9019);
nor U9949 (N_9949,N_9127,N_9024);
and U9950 (N_9950,N_9372,N_9404);
and U9951 (N_9951,N_9043,N_9272);
and U9952 (N_9952,N_9172,N_9338);
or U9953 (N_9953,N_9345,N_9124);
xnor U9954 (N_9954,N_9143,N_9341);
or U9955 (N_9955,N_9408,N_9412);
nor U9956 (N_9956,N_9108,N_9110);
nor U9957 (N_9957,N_9433,N_9176);
nand U9958 (N_9958,N_9454,N_9438);
and U9959 (N_9959,N_9121,N_9017);
nor U9960 (N_9960,N_9185,N_9081);
or U9961 (N_9961,N_9473,N_9484);
nor U9962 (N_9962,N_9100,N_9341);
or U9963 (N_9963,N_9441,N_9112);
or U9964 (N_9964,N_9323,N_9444);
and U9965 (N_9965,N_9200,N_9020);
nor U9966 (N_9966,N_9360,N_9039);
nand U9967 (N_9967,N_9002,N_9436);
or U9968 (N_9968,N_9497,N_9416);
and U9969 (N_9969,N_9438,N_9278);
or U9970 (N_9970,N_9417,N_9021);
or U9971 (N_9971,N_9456,N_9266);
nand U9972 (N_9972,N_9057,N_9065);
nor U9973 (N_9973,N_9021,N_9327);
nand U9974 (N_9974,N_9103,N_9022);
and U9975 (N_9975,N_9011,N_9073);
nand U9976 (N_9976,N_9089,N_9203);
nand U9977 (N_9977,N_9174,N_9324);
xnor U9978 (N_9978,N_9224,N_9084);
and U9979 (N_9979,N_9403,N_9084);
nor U9980 (N_9980,N_9069,N_9032);
xnor U9981 (N_9981,N_9089,N_9371);
nor U9982 (N_9982,N_9045,N_9049);
or U9983 (N_9983,N_9148,N_9460);
nand U9984 (N_9984,N_9024,N_9003);
or U9985 (N_9985,N_9294,N_9318);
nand U9986 (N_9986,N_9480,N_9025);
and U9987 (N_9987,N_9386,N_9091);
and U9988 (N_9988,N_9376,N_9220);
and U9989 (N_9989,N_9294,N_9214);
or U9990 (N_9990,N_9148,N_9027);
or U9991 (N_9991,N_9380,N_9420);
or U9992 (N_9992,N_9383,N_9450);
nand U9993 (N_9993,N_9173,N_9121);
nor U9994 (N_9994,N_9159,N_9049);
nor U9995 (N_9995,N_9091,N_9352);
and U9996 (N_9996,N_9180,N_9261);
nor U9997 (N_9997,N_9116,N_9072);
nor U9998 (N_9998,N_9148,N_9327);
and U9999 (N_9999,N_9112,N_9293);
nand U10000 (N_10000,N_9637,N_9956);
or U10001 (N_10001,N_9911,N_9536);
and U10002 (N_10002,N_9561,N_9793);
and U10003 (N_10003,N_9665,N_9722);
nor U10004 (N_10004,N_9878,N_9917);
or U10005 (N_10005,N_9539,N_9875);
or U10006 (N_10006,N_9629,N_9585);
nand U10007 (N_10007,N_9945,N_9803);
nor U10008 (N_10008,N_9814,N_9997);
nor U10009 (N_10009,N_9867,N_9932);
and U10010 (N_10010,N_9720,N_9656);
nor U10011 (N_10011,N_9916,N_9923);
nor U10012 (N_10012,N_9526,N_9896);
nor U10013 (N_10013,N_9568,N_9571);
or U10014 (N_10014,N_9602,N_9952);
nand U10015 (N_10015,N_9920,N_9745);
or U10016 (N_10016,N_9654,N_9548);
or U10017 (N_10017,N_9596,N_9749);
nor U10018 (N_10018,N_9870,N_9826);
nor U10019 (N_10019,N_9809,N_9759);
or U10020 (N_10020,N_9634,N_9753);
xor U10021 (N_10021,N_9884,N_9863);
and U10022 (N_10022,N_9808,N_9984);
and U10023 (N_10023,N_9892,N_9635);
or U10024 (N_10024,N_9847,N_9992);
and U10025 (N_10025,N_9591,N_9671);
xor U10026 (N_10026,N_9550,N_9915);
and U10027 (N_10027,N_9855,N_9523);
nor U10028 (N_10028,N_9924,N_9633);
nand U10029 (N_10029,N_9704,N_9948);
or U10030 (N_10030,N_9609,N_9850);
nand U10031 (N_10031,N_9686,N_9670);
nand U10032 (N_10032,N_9623,N_9786);
and U10033 (N_10033,N_9765,N_9569);
and U10034 (N_10034,N_9725,N_9528);
nor U10035 (N_10035,N_9873,N_9811);
nor U10036 (N_10036,N_9921,N_9513);
and U10037 (N_10037,N_9594,N_9740);
or U10038 (N_10038,N_9677,N_9607);
and U10039 (N_10039,N_9859,N_9869);
or U10040 (N_10040,N_9780,N_9868);
and U10041 (N_10041,N_9913,N_9564);
nand U10042 (N_10042,N_9897,N_9937);
and U10043 (N_10043,N_9746,N_9584);
or U10044 (N_10044,N_9903,N_9515);
nand U10045 (N_10045,N_9895,N_9621);
or U10046 (N_10046,N_9519,N_9522);
or U10047 (N_10047,N_9620,N_9919);
nor U10048 (N_10048,N_9643,N_9936);
or U10049 (N_10049,N_9974,N_9821);
nor U10050 (N_10050,N_9905,N_9706);
or U10051 (N_10051,N_9805,N_9611);
nand U10052 (N_10052,N_9701,N_9632);
nand U10053 (N_10053,N_9510,N_9800);
xor U10054 (N_10054,N_9710,N_9781);
and U10055 (N_10055,N_9727,N_9879);
nor U10056 (N_10056,N_9739,N_9991);
and U10057 (N_10057,N_9852,N_9846);
or U10058 (N_10058,N_9723,N_9978);
or U10059 (N_10059,N_9653,N_9731);
and U10060 (N_10060,N_9856,N_9538);
and U10061 (N_10061,N_9963,N_9711);
or U10062 (N_10062,N_9823,N_9505);
nand U10063 (N_10063,N_9807,N_9982);
or U10064 (N_10064,N_9999,N_9719);
and U10065 (N_10065,N_9950,N_9586);
and U10066 (N_10066,N_9552,N_9625);
and U10067 (N_10067,N_9973,N_9819);
nor U10068 (N_10068,N_9693,N_9681);
nor U10069 (N_10069,N_9648,N_9549);
or U10070 (N_10070,N_9883,N_9672);
nand U10071 (N_10071,N_9601,N_9931);
or U10072 (N_10072,N_9766,N_9810);
nor U10073 (N_10073,N_9597,N_9589);
xor U10074 (N_10074,N_9957,N_9553);
xor U10075 (N_10075,N_9871,N_9705);
or U10076 (N_10076,N_9646,N_9631);
and U10077 (N_10077,N_9688,N_9860);
nor U10078 (N_10078,N_9960,N_9815);
and U10079 (N_10079,N_9764,N_9575);
xnor U10080 (N_10080,N_9730,N_9881);
nand U10081 (N_10081,N_9941,N_9799);
nand U10082 (N_10082,N_9858,N_9985);
or U10083 (N_10083,N_9679,N_9747);
nand U10084 (N_10084,N_9876,N_9975);
or U10085 (N_10085,N_9946,N_9694);
nand U10086 (N_10086,N_9912,N_9885);
nor U10087 (N_10087,N_9544,N_9582);
nand U10088 (N_10088,N_9980,N_9794);
nand U10089 (N_10089,N_9728,N_9587);
nor U10090 (N_10090,N_9790,N_9954);
or U10091 (N_10091,N_9752,N_9914);
or U10092 (N_10092,N_9851,N_9817);
nand U10093 (N_10093,N_9741,N_9567);
and U10094 (N_10094,N_9675,N_9669);
and U10095 (N_10095,N_9576,N_9877);
or U10096 (N_10096,N_9806,N_9667);
and U10097 (N_10097,N_9848,N_9525);
nand U10098 (N_10098,N_9690,N_9755);
nor U10099 (N_10099,N_9713,N_9909);
nand U10100 (N_10100,N_9599,N_9530);
and U10101 (N_10101,N_9760,N_9717);
nand U10102 (N_10102,N_9647,N_9762);
nor U10103 (N_10103,N_9773,N_9829);
nand U10104 (N_10104,N_9529,N_9804);
and U10105 (N_10105,N_9674,N_9733);
or U10106 (N_10106,N_9813,N_9619);
nor U10107 (N_10107,N_9506,N_9904);
and U10108 (N_10108,N_9559,N_9865);
nand U10109 (N_10109,N_9666,N_9951);
nand U10110 (N_10110,N_9732,N_9907);
or U10111 (N_10111,N_9577,N_9610);
nor U10112 (N_10112,N_9827,N_9535);
nand U10113 (N_10113,N_9579,N_9930);
or U10114 (N_10114,N_9664,N_9708);
nand U10115 (N_10115,N_9612,N_9540);
or U10116 (N_10116,N_9614,N_9928);
and U10117 (N_10117,N_9668,N_9685);
nand U10118 (N_10118,N_9798,N_9583);
nand U10119 (N_10119,N_9650,N_9716);
nand U10120 (N_10120,N_9862,N_9703);
or U10121 (N_10121,N_9958,N_9812);
nand U10122 (N_10122,N_9545,N_9508);
nor U10123 (N_10123,N_9709,N_9906);
xor U10124 (N_10124,N_9959,N_9645);
nand U10125 (N_10125,N_9615,N_9593);
or U10126 (N_10126,N_9788,N_9758);
and U10127 (N_10127,N_9825,N_9830);
xnor U10128 (N_10128,N_9588,N_9757);
nor U10129 (N_10129,N_9659,N_9735);
or U10130 (N_10130,N_9696,N_9961);
nor U10131 (N_10131,N_9533,N_9543);
or U10132 (N_10132,N_9922,N_9843);
nor U10133 (N_10133,N_9501,N_9699);
or U10134 (N_10134,N_9581,N_9898);
and U10135 (N_10135,N_9616,N_9617);
or U10136 (N_10136,N_9763,N_9784);
nand U10137 (N_10137,N_9831,N_9866);
or U10138 (N_10138,N_9792,N_9700);
xnor U10139 (N_10139,N_9775,N_9857);
and U10140 (N_10140,N_9642,N_9853);
nor U10141 (N_10141,N_9874,N_9592);
or U10142 (N_10142,N_9649,N_9558);
nand U10143 (N_10143,N_9887,N_9729);
or U10144 (N_10144,N_9880,N_9743);
nor U10145 (N_10145,N_9531,N_9901);
xnor U10146 (N_10146,N_9692,N_9964);
xor U10147 (N_10147,N_9943,N_9570);
and U10148 (N_10148,N_9556,N_9899);
nor U10149 (N_10149,N_9840,N_9524);
and U10150 (N_10150,N_9834,N_9551);
or U10151 (N_10151,N_9971,N_9657);
nand U10152 (N_10152,N_9787,N_9748);
and U10153 (N_10153,N_9547,N_9605);
nand U10154 (N_10154,N_9768,N_9707);
or U10155 (N_10155,N_9844,N_9507);
and U10156 (N_10156,N_9562,N_9691);
nand U10157 (N_10157,N_9718,N_9998);
nand U10158 (N_10158,N_9761,N_9689);
xor U10159 (N_10159,N_9640,N_9702);
and U10160 (N_10160,N_9949,N_9795);
and U10161 (N_10161,N_9514,N_9776);
and U10162 (N_10162,N_9512,N_9734);
and U10163 (N_10163,N_9680,N_9608);
nor U10164 (N_10164,N_9947,N_9563);
nor U10165 (N_10165,N_9972,N_9796);
xor U10166 (N_10166,N_9600,N_9944);
or U10167 (N_10167,N_9996,N_9777);
nor U10168 (N_10168,N_9993,N_9663);
nor U10169 (N_10169,N_9767,N_9890);
xnor U10170 (N_10170,N_9966,N_9824);
xnor U10171 (N_10171,N_9983,N_9864);
nand U10172 (N_10172,N_9933,N_9782);
nor U10173 (N_10173,N_9791,N_9894);
nand U10174 (N_10174,N_9908,N_9662);
xnor U10175 (N_10175,N_9990,N_9988);
nand U10176 (N_10176,N_9683,N_9517);
or U10177 (N_10177,N_9839,N_9835);
nor U10178 (N_10178,N_9560,N_9977);
or U10179 (N_10179,N_9886,N_9698);
or U10180 (N_10180,N_9801,N_9836);
xnor U10181 (N_10181,N_9816,N_9989);
or U10182 (N_10182,N_9500,N_9968);
and U10183 (N_10183,N_9622,N_9687);
nand U10184 (N_10184,N_9516,N_9965);
and U10185 (N_10185,N_9606,N_9527);
nand U10186 (N_10186,N_9572,N_9818);
and U10187 (N_10187,N_9891,N_9918);
xor U10188 (N_10188,N_9861,N_9627);
xor U10189 (N_10189,N_9833,N_9888);
or U10190 (N_10190,N_9603,N_9882);
and U10191 (N_10191,N_9967,N_9715);
or U10192 (N_10192,N_9981,N_9573);
or U10193 (N_10193,N_9638,N_9938);
and U10194 (N_10194,N_9541,N_9987);
nor U10195 (N_10195,N_9976,N_9969);
or U10196 (N_10196,N_9845,N_9756);
and U10197 (N_10197,N_9737,N_9953);
or U10198 (N_10198,N_9789,N_9721);
or U10199 (N_10199,N_9511,N_9682);
nand U10200 (N_10200,N_9520,N_9566);
and U10201 (N_10201,N_9636,N_9962);
nand U10202 (N_10202,N_9652,N_9769);
xor U10203 (N_10203,N_9695,N_9546);
and U10204 (N_10204,N_9772,N_9678);
or U10205 (N_10205,N_9574,N_9750);
and U10206 (N_10206,N_9641,N_9939);
or U10207 (N_10207,N_9509,N_9841);
xnor U10208 (N_10208,N_9578,N_9580);
nand U10209 (N_10209,N_9712,N_9837);
xnor U10210 (N_10210,N_9661,N_9714);
and U10211 (N_10211,N_9935,N_9742);
and U10212 (N_10212,N_9828,N_9502);
nand U10213 (N_10213,N_9854,N_9630);
nor U10214 (N_10214,N_9521,N_9557);
nand U10215 (N_10215,N_9751,N_9555);
and U10216 (N_10216,N_9849,N_9503);
nor U10217 (N_10217,N_9684,N_9639);
nand U10218 (N_10218,N_9926,N_9925);
xor U10219 (N_10219,N_9942,N_9628);
and U10220 (N_10220,N_9779,N_9774);
and U10221 (N_10221,N_9726,N_9658);
and U10222 (N_10222,N_9820,N_9783);
and U10223 (N_10223,N_9532,N_9832);
nand U10224 (N_10224,N_9979,N_9534);
nand U10225 (N_10225,N_9934,N_9771);
xor U10226 (N_10226,N_9644,N_9595);
or U10227 (N_10227,N_9673,N_9955);
and U10228 (N_10228,N_9565,N_9900);
and U10229 (N_10229,N_9598,N_9724);
and U10230 (N_10230,N_9744,N_9626);
nor U10231 (N_10231,N_9590,N_9994);
nand U10232 (N_10232,N_9655,N_9929);
nor U10233 (N_10233,N_9537,N_9778);
nor U10234 (N_10234,N_9651,N_9660);
or U10235 (N_10235,N_9613,N_9554);
xnor U10236 (N_10236,N_9872,N_9940);
nor U10237 (N_10237,N_9754,N_9738);
nand U10238 (N_10238,N_9986,N_9838);
nand U10239 (N_10239,N_9736,N_9802);
and U10240 (N_10240,N_9893,N_9902);
or U10241 (N_10241,N_9504,N_9785);
nand U10242 (N_10242,N_9676,N_9770);
nand U10243 (N_10243,N_9604,N_9542);
or U10244 (N_10244,N_9624,N_9618);
xor U10245 (N_10245,N_9797,N_9518);
nor U10246 (N_10246,N_9889,N_9970);
or U10247 (N_10247,N_9995,N_9842);
nor U10248 (N_10248,N_9697,N_9910);
and U10249 (N_10249,N_9822,N_9927);
and U10250 (N_10250,N_9986,N_9991);
or U10251 (N_10251,N_9578,N_9943);
nor U10252 (N_10252,N_9643,N_9816);
and U10253 (N_10253,N_9785,N_9512);
nand U10254 (N_10254,N_9755,N_9875);
nor U10255 (N_10255,N_9542,N_9975);
nand U10256 (N_10256,N_9882,N_9573);
nor U10257 (N_10257,N_9894,N_9551);
nor U10258 (N_10258,N_9851,N_9870);
or U10259 (N_10259,N_9541,N_9595);
and U10260 (N_10260,N_9567,N_9917);
or U10261 (N_10261,N_9608,N_9627);
and U10262 (N_10262,N_9941,N_9847);
nand U10263 (N_10263,N_9646,N_9784);
nor U10264 (N_10264,N_9560,N_9673);
nor U10265 (N_10265,N_9616,N_9729);
or U10266 (N_10266,N_9973,N_9523);
or U10267 (N_10267,N_9958,N_9989);
xnor U10268 (N_10268,N_9751,N_9673);
or U10269 (N_10269,N_9791,N_9710);
or U10270 (N_10270,N_9516,N_9921);
nor U10271 (N_10271,N_9724,N_9723);
or U10272 (N_10272,N_9528,N_9775);
nand U10273 (N_10273,N_9518,N_9695);
nor U10274 (N_10274,N_9605,N_9970);
nor U10275 (N_10275,N_9710,N_9648);
or U10276 (N_10276,N_9557,N_9931);
or U10277 (N_10277,N_9618,N_9803);
nor U10278 (N_10278,N_9979,N_9600);
or U10279 (N_10279,N_9839,N_9713);
or U10280 (N_10280,N_9685,N_9616);
or U10281 (N_10281,N_9950,N_9632);
nand U10282 (N_10282,N_9649,N_9958);
xnor U10283 (N_10283,N_9932,N_9648);
or U10284 (N_10284,N_9979,N_9674);
and U10285 (N_10285,N_9743,N_9989);
nor U10286 (N_10286,N_9790,N_9908);
nor U10287 (N_10287,N_9675,N_9963);
nand U10288 (N_10288,N_9993,N_9706);
and U10289 (N_10289,N_9526,N_9596);
xor U10290 (N_10290,N_9789,N_9904);
nor U10291 (N_10291,N_9659,N_9884);
and U10292 (N_10292,N_9527,N_9743);
or U10293 (N_10293,N_9730,N_9622);
and U10294 (N_10294,N_9850,N_9879);
and U10295 (N_10295,N_9949,N_9730);
and U10296 (N_10296,N_9706,N_9918);
or U10297 (N_10297,N_9681,N_9618);
or U10298 (N_10298,N_9993,N_9821);
nor U10299 (N_10299,N_9671,N_9805);
xor U10300 (N_10300,N_9550,N_9874);
nor U10301 (N_10301,N_9963,N_9611);
and U10302 (N_10302,N_9996,N_9727);
or U10303 (N_10303,N_9947,N_9953);
and U10304 (N_10304,N_9715,N_9547);
and U10305 (N_10305,N_9577,N_9776);
nor U10306 (N_10306,N_9731,N_9566);
xor U10307 (N_10307,N_9847,N_9886);
nand U10308 (N_10308,N_9804,N_9997);
nand U10309 (N_10309,N_9853,N_9611);
nand U10310 (N_10310,N_9905,N_9611);
and U10311 (N_10311,N_9659,N_9681);
nand U10312 (N_10312,N_9846,N_9969);
or U10313 (N_10313,N_9829,N_9908);
nor U10314 (N_10314,N_9751,N_9500);
or U10315 (N_10315,N_9569,N_9745);
and U10316 (N_10316,N_9531,N_9838);
or U10317 (N_10317,N_9756,N_9568);
and U10318 (N_10318,N_9830,N_9611);
or U10319 (N_10319,N_9860,N_9966);
and U10320 (N_10320,N_9798,N_9606);
xor U10321 (N_10321,N_9884,N_9707);
xor U10322 (N_10322,N_9837,N_9789);
xnor U10323 (N_10323,N_9777,N_9686);
or U10324 (N_10324,N_9869,N_9560);
nand U10325 (N_10325,N_9556,N_9949);
and U10326 (N_10326,N_9862,N_9898);
nor U10327 (N_10327,N_9943,N_9533);
or U10328 (N_10328,N_9662,N_9817);
nor U10329 (N_10329,N_9998,N_9649);
and U10330 (N_10330,N_9685,N_9660);
xnor U10331 (N_10331,N_9741,N_9780);
nand U10332 (N_10332,N_9563,N_9517);
nand U10333 (N_10333,N_9650,N_9800);
and U10334 (N_10334,N_9817,N_9501);
nand U10335 (N_10335,N_9744,N_9618);
nand U10336 (N_10336,N_9552,N_9995);
and U10337 (N_10337,N_9950,N_9674);
or U10338 (N_10338,N_9613,N_9551);
and U10339 (N_10339,N_9617,N_9729);
nand U10340 (N_10340,N_9782,N_9775);
and U10341 (N_10341,N_9863,N_9504);
and U10342 (N_10342,N_9746,N_9690);
nor U10343 (N_10343,N_9956,N_9841);
nor U10344 (N_10344,N_9899,N_9747);
or U10345 (N_10345,N_9655,N_9841);
nand U10346 (N_10346,N_9572,N_9641);
or U10347 (N_10347,N_9855,N_9843);
or U10348 (N_10348,N_9560,N_9597);
or U10349 (N_10349,N_9842,N_9732);
and U10350 (N_10350,N_9549,N_9847);
and U10351 (N_10351,N_9771,N_9656);
xnor U10352 (N_10352,N_9806,N_9885);
nand U10353 (N_10353,N_9507,N_9850);
nand U10354 (N_10354,N_9609,N_9801);
nor U10355 (N_10355,N_9547,N_9972);
or U10356 (N_10356,N_9927,N_9940);
nand U10357 (N_10357,N_9933,N_9913);
and U10358 (N_10358,N_9923,N_9954);
nor U10359 (N_10359,N_9743,N_9641);
nand U10360 (N_10360,N_9900,N_9579);
nor U10361 (N_10361,N_9769,N_9913);
nor U10362 (N_10362,N_9971,N_9946);
nand U10363 (N_10363,N_9856,N_9696);
nor U10364 (N_10364,N_9748,N_9678);
or U10365 (N_10365,N_9713,N_9932);
nand U10366 (N_10366,N_9699,N_9878);
nor U10367 (N_10367,N_9660,N_9850);
nand U10368 (N_10368,N_9825,N_9572);
nand U10369 (N_10369,N_9942,N_9696);
and U10370 (N_10370,N_9828,N_9721);
and U10371 (N_10371,N_9612,N_9697);
and U10372 (N_10372,N_9554,N_9555);
nor U10373 (N_10373,N_9513,N_9593);
nor U10374 (N_10374,N_9751,N_9545);
and U10375 (N_10375,N_9787,N_9871);
or U10376 (N_10376,N_9761,N_9580);
nand U10377 (N_10377,N_9682,N_9846);
nand U10378 (N_10378,N_9999,N_9665);
nand U10379 (N_10379,N_9841,N_9597);
xnor U10380 (N_10380,N_9703,N_9971);
and U10381 (N_10381,N_9565,N_9989);
xnor U10382 (N_10382,N_9727,N_9708);
nand U10383 (N_10383,N_9966,N_9952);
and U10384 (N_10384,N_9519,N_9794);
or U10385 (N_10385,N_9553,N_9846);
and U10386 (N_10386,N_9743,N_9728);
or U10387 (N_10387,N_9588,N_9897);
and U10388 (N_10388,N_9922,N_9504);
or U10389 (N_10389,N_9601,N_9884);
nand U10390 (N_10390,N_9518,N_9948);
and U10391 (N_10391,N_9697,N_9547);
and U10392 (N_10392,N_9721,N_9983);
nor U10393 (N_10393,N_9977,N_9637);
nand U10394 (N_10394,N_9824,N_9961);
or U10395 (N_10395,N_9774,N_9787);
and U10396 (N_10396,N_9869,N_9523);
and U10397 (N_10397,N_9894,N_9521);
and U10398 (N_10398,N_9663,N_9784);
or U10399 (N_10399,N_9636,N_9575);
nand U10400 (N_10400,N_9774,N_9595);
nand U10401 (N_10401,N_9765,N_9845);
nand U10402 (N_10402,N_9748,N_9708);
or U10403 (N_10403,N_9911,N_9938);
or U10404 (N_10404,N_9973,N_9633);
nor U10405 (N_10405,N_9631,N_9812);
and U10406 (N_10406,N_9783,N_9941);
or U10407 (N_10407,N_9818,N_9695);
nor U10408 (N_10408,N_9736,N_9746);
or U10409 (N_10409,N_9910,N_9851);
nor U10410 (N_10410,N_9808,N_9548);
nand U10411 (N_10411,N_9709,N_9729);
and U10412 (N_10412,N_9775,N_9566);
or U10413 (N_10413,N_9703,N_9681);
nand U10414 (N_10414,N_9777,N_9569);
nand U10415 (N_10415,N_9781,N_9973);
or U10416 (N_10416,N_9755,N_9594);
or U10417 (N_10417,N_9743,N_9622);
nand U10418 (N_10418,N_9783,N_9588);
or U10419 (N_10419,N_9901,N_9555);
nor U10420 (N_10420,N_9560,N_9611);
or U10421 (N_10421,N_9941,N_9717);
nor U10422 (N_10422,N_9954,N_9744);
nor U10423 (N_10423,N_9842,N_9834);
nor U10424 (N_10424,N_9565,N_9729);
or U10425 (N_10425,N_9768,N_9765);
or U10426 (N_10426,N_9668,N_9884);
and U10427 (N_10427,N_9870,N_9694);
xor U10428 (N_10428,N_9943,N_9689);
nor U10429 (N_10429,N_9626,N_9519);
and U10430 (N_10430,N_9895,N_9500);
or U10431 (N_10431,N_9903,N_9773);
and U10432 (N_10432,N_9743,N_9978);
nand U10433 (N_10433,N_9596,N_9620);
xnor U10434 (N_10434,N_9741,N_9668);
and U10435 (N_10435,N_9956,N_9546);
and U10436 (N_10436,N_9724,N_9505);
and U10437 (N_10437,N_9800,N_9913);
nor U10438 (N_10438,N_9569,N_9717);
or U10439 (N_10439,N_9717,N_9944);
or U10440 (N_10440,N_9935,N_9900);
or U10441 (N_10441,N_9536,N_9769);
or U10442 (N_10442,N_9780,N_9730);
or U10443 (N_10443,N_9529,N_9563);
nor U10444 (N_10444,N_9835,N_9578);
nor U10445 (N_10445,N_9917,N_9828);
and U10446 (N_10446,N_9778,N_9878);
or U10447 (N_10447,N_9815,N_9592);
nand U10448 (N_10448,N_9702,N_9676);
or U10449 (N_10449,N_9846,N_9959);
nor U10450 (N_10450,N_9861,N_9712);
and U10451 (N_10451,N_9670,N_9812);
nand U10452 (N_10452,N_9905,N_9980);
nand U10453 (N_10453,N_9992,N_9951);
nand U10454 (N_10454,N_9563,N_9672);
and U10455 (N_10455,N_9873,N_9613);
or U10456 (N_10456,N_9829,N_9778);
or U10457 (N_10457,N_9681,N_9780);
nor U10458 (N_10458,N_9832,N_9609);
or U10459 (N_10459,N_9928,N_9883);
nand U10460 (N_10460,N_9577,N_9903);
nor U10461 (N_10461,N_9931,N_9776);
nand U10462 (N_10462,N_9731,N_9504);
xnor U10463 (N_10463,N_9805,N_9724);
or U10464 (N_10464,N_9797,N_9864);
nand U10465 (N_10465,N_9947,N_9940);
nor U10466 (N_10466,N_9943,N_9860);
and U10467 (N_10467,N_9572,N_9551);
and U10468 (N_10468,N_9810,N_9788);
and U10469 (N_10469,N_9838,N_9512);
or U10470 (N_10470,N_9682,N_9501);
or U10471 (N_10471,N_9726,N_9690);
and U10472 (N_10472,N_9947,N_9510);
xor U10473 (N_10473,N_9658,N_9715);
nand U10474 (N_10474,N_9678,N_9809);
xnor U10475 (N_10475,N_9663,N_9909);
nor U10476 (N_10476,N_9869,N_9617);
or U10477 (N_10477,N_9734,N_9997);
and U10478 (N_10478,N_9673,N_9562);
or U10479 (N_10479,N_9853,N_9995);
nor U10480 (N_10480,N_9522,N_9999);
or U10481 (N_10481,N_9606,N_9739);
xnor U10482 (N_10482,N_9514,N_9725);
and U10483 (N_10483,N_9635,N_9902);
nand U10484 (N_10484,N_9676,N_9647);
or U10485 (N_10485,N_9823,N_9500);
and U10486 (N_10486,N_9938,N_9769);
and U10487 (N_10487,N_9730,N_9993);
or U10488 (N_10488,N_9650,N_9525);
or U10489 (N_10489,N_9552,N_9814);
or U10490 (N_10490,N_9552,N_9697);
xnor U10491 (N_10491,N_9602,N_9877);
and U10492 (N_10492,N_9922,N_9661);
or U10493 (N_10493,N_9666,N_9628);
and U10494 (N_10494,N_9582,N_9975);
or U10495 (N_10495,N_9950,N_9845);
or U10496 (N_10496,N_9811,N_9609);
nor U10497 (N_10497,N_9732,N_9658);
nor U10498 (N_10498,N_9610,N_9863);
nor U10499 (N_10499,N_9648,N_9604);
xor U10500 (N_10500,N_10214,N_10189);
or U10501 (N_10501,N_10253,N_10219);
nand U10502 (N_10502,N_10074,N_10043);
nand U10503 (N_10503,N_10309,N_10421);
or U10504 (N_10504,N_10291,N_10297);
nand U10505 (N_10505,N_10484,N_10248);
or U10506 (N_10506,N_10403,N_10141);
and U10507 (N_10507,N_10488,N_10075);
nand U10508 (N_10508,N_10149,N_10486);
and U10509 (N_10509,N_10479,N_10265);
nor U10510 (N_10510,N_10213,N_10031);
nor U10511 (N_10511,N_10122,N_10208);
nand U10512 (N_10512,N_10015,N_10279);
xnor U10513 (N_10513,N_10295,N_10281);
nor U10514 (N_10514,N_10400,N_10084);
and U10515 (N_10515,N_10076,N_10044);
nand U10516 (N_10516,N_10337,N_10409);
or U10517 (N_10517,N_10086,N_10264);
nor U10518 (N_10518,N_10046,N_10103);
or U10519 (N_10519,N_10331,N_10407);
nor U10520 (N_10520,N_10161,N_10092);
or U10521 (N_10521,N_10380,N_10470);
or U10522 (N_10522,N_10474,N_10019);
xnor U10523 (N_10523,N_10244,N_10093);
and U10524 (N_10524,N_10229,N_10465);
and U10525 (N_10525,N_10481,N_10146);
nor U10526 (N_10526,N_10017,N_10196);
nand U10527 (N_10527,N_10289,N_10237);
nand U10528 (N_10528,N_10322,N_10143);
and U10529 (N_10529,N_10471,N_10088);
and U10530 (N_10530,N_10449,N_10406);
xor U10531 (N_10531,N_10356,N_10355);
nor U10532 (N_10532,N_10414,N_10447);
and U10533 (N_10533,N_10452,N_10095);
or U10534 (N_10534,N_10311,N_10178);
or U10535 (N_10535,N_10433,N_10105);
and U10536 (N_10536,N_10317,N_10169);
nand U10537 (N_10537,N_10390,N_10206);
and U10538 (N_10538,N_10170,N_10341);
nand U10539 (N_10539,N_10137,N_10024);
and U10540 (N_10540,N_10358,N_10333);
nand U10541 (N_10541,N_10345,N_10454);
or U10542 (N_10542,N_10118,N_10321);
nand U10543 (N_10543,N_10401,N_10393);
or U10544 (N_10544,N_10307,N_10426);
or U10545 (N_10545,N_10000,N_10293);
xor U10546 (N_10546,N_10082,N_10312);
and U10547 (N_10547,N_10362,N_10197);
or U10548 (N_10548,N_10363,N_10437);
nand U10549 (N_10549,N_10218,N_10418);
nand U10550 (N_10550,N_10368,N_10370);
and U10551 (N_10551,N_10202,N_10032);
and U10552 (N_10552,N_10156,N_10282);
and U10553 (N_10553,N_10379,N_10480);
and U10554 (N_10554,N_10301,N_10065);
or U10555 (N_10555,N_10090,N_10242);
and U10556 (N_10556,N_10062,N_10008);
nor U10557 (N_10557,N_10323,N_10305);
or U10558 (N_10558,N_10115,N_10059);
nand U10559 (N_10559,N_10306,N_10273);
xor U10560 (N_10560,N_10274,N_10376);
and U10561 (N_10561,N_10124,N_10190);
and U10562 (N_10562,N_10014,N_10034);
and U10563 (N_10563,N_10210,N_10316);
nor U10564 (N_10564,N_10155,N_10159);
nand U10565 (N_10565,N_10334,N_10441);
nor U10566 (N_10566,N_10292,N_10233);
and U10567 (N_10567,N_10226,N_10119);
nor U10568 (N_10568,N_10182,N_10395);
nor U10569 (N_10569,N_10250,N_10187);
nand U10570 (N_10570,N_10058,N_10440);
or U10571 (N_10571,N_10123,N_10108);
or U10572 (N_10572,N_10147,N_10113);
or U10573 (N_10573,N_10102,N_10021);
xor U10574 (N_10574,N_10361,N_10016);
nand U10575 (N_10575,N_10462,N_10377);
nor U10576 (N_10576,N_10194,N_10201);
nand U10577 (N_10577,N_10410,N_10192);
and U10578 (N_10578,N_10114,N_10129);
and U10579 (N_10579,N_10396,N_10445);
or U10580 (N_10580,N_10041,N_10221);
nor U10581 (N_10581,N_10397,N_10402);
nor U10582 (N_10582,N_10227,N_10033);
nand U10583 (N_10583,N_10405,N_10284);
nand U10584 (N_10584,N_10029,N_10097);
nand U10585 (N_10585,N_10139,N_10286);
and U10586 (N_10586,N_10104,N_10223);
and U10587 (N_10587,N_10061,N_10298);
nand U10588 (N_10588,N_10175,N_10472);
nand U10589 (N_10589,N_10039,N_10080);
and U10590 (N_10590,N_10257,N_10158);
nand U10591 (N_10591,N_10482,N_10398);
nor U10592 (N_10592,N_10374,N_10007);
and U10593 (N_10593,N_10300,N_10430);
or U10594 (N_10594,N_10364,N_10205);
nand U10595 (N_10595,N_10375,N_10270);
or U10596 (N_10596,N_10348,N_10340);
or U10597 (N_10597,N_10243,N_10168);
xnor U10598 (N_10598,N_10290,N_10199);
and U10599 (N_10599,N_10180,N_10249);
or U10600 (N_10600,N_10408,N_10325);
or U10601 (N_10601,N_10132,N_10451);
or U10602 (N_10602,N_10278,N_10195);
nand U10603 (N_10603,N_10391,N_10036);
nor U10604 (N_10604,N_10394,N_10424);
nor U10605 (N_10605,N_10277,N_10164);
and U10606 (N_10606,N_10037,N_10354);
xor U10607 (N_10607,N_10177,N_10204);
xor U10608 (N_10608,N_10176,N_10018);
or U10609 (N_10609,N_10171,N_10269);
nand U10610 (N_10610,N_10130,N_10497);
nand U10611 (N_10611,N_10438,N_10285);
nor U10612 (N_10612,N_10150,N_10186);
nand U10613 (N_10613,N_10381,N_10372);
and U10614 (N_10614,N_10385,N_10200);
nand U10615 (N_10615,N_10496,N_10136);
nor U10616 (N_10616,N_10078,N_10121);
or U10617 (N_10617,N_10045,N_10296);
and U10618 (N_10618,N_10425,N_10431);
nand U10619 (N_10619,N_10299,N_10271);
nor U10620 (N_10620,N_10079,N_10209);
nor U10621 (N_10621,N_10070,N_10366);
nor U10622 (N_10622,N_10392,N_10020);
nor U10623 (N_10623,N_10461,N_10220);
or U10624 (N_10624,N_10254,N_10140);
or U10625 (N_10625,N_10085,N_10399);
or U10626 (N_10626,N_10083,N_10326);
nand U10627 (N_10627,N_10157,N_10047);
nand U10628 (N_10628,N_10099,N_10423);
nor U10629 (N_10629,N_10126,N_10288);
nand U10630 (N_10630,N_10303,N_10359);
nand U10631 (N_10631,N_10003,N_10420);
and U10632 (N_10632,N_10067,N_10049);
or U10633 (N_10633,N_10138,N_10444);
and U10634 (N_10634,N_10324,N_10346);
and U10635 (N_10635,N_10276,N_10238);
or U10636 (N_10636,N_10001,N_10128);
and U10637 (N_10637,N_10263,N_10258);
or U10638 (N_10638,N_10225,N_10330);
and U10639 (N_10639,N_10495,N_10283);
and U10640 (N_10640,N_10153,N_10308);
and U10641 (N_10641,N_10055,N_10371);
xor U10642 (N_10642,N_10148,N_10328);
nor U10643 (N_10643,N_10310,N_10228);
nand U10644 (N_10644,N_10280,N_10339);
or U10645 (N_10645,N_10173,N_10203);
xnor U10646 (N_10646,N_10260,N_10096);
or U10647 (N_10647,N_10357,N_10107);
and U10648 (N_10648,N_10456,N_10051);
nand U10649 (N_10649,N_10490,N_10477);
or U10650 (N_10650,N_10439,N_10131);
nor U10651 (N_10651,N_10347,N_10302);
or U10652 (N_10652,N_10351,N_10411);
and U10653 (N_10653,N_10338,N_10378);
nand U10654 (N_10654,N_10382,N_10010);
and U10655 (N_10655,N_10224,N_10460);
and U10656 (N_10656,N_10335,N_10446);
or U10657 (N_10657,N_10434,N_10476);
nor U10658 (N_10658,N_10314,N_10185);
xnor U10659 (N_10659,N_10360,N_10125);
and U10660 (N_10660,N_10499,N_10184);
nand U10661 (N_10661,N_10081,N_10116);
nand U10662 (N_10662,N_10054,N_10230);
and U10663 (N_10663,N_10268,N_10012);
nor U10664 (N_10664,N_10135,N_10193);
and U10665 (N_10665,N_10167,N_10313);
nor U10666 (N_10666,N_10384,N_10367);
or U10667 (N_10667,N_10256,N_10098);
nand U10668 (N_10668,N_10231,N_10198);
nand U10669 (N_10669,N_10013,N_10365);
or U10670 (N_10670,N_10207,N_10174);
nand U10671 (N_10671,N_10110,N_10318);
nand U10672 (N_10672,N_10412,N_10152);
or U10673 (N_10673,N_10216,N_10235);
nor U10674 (N_10674,N_10315,N_10154);
nand U10675 (N_10675,N_10166,N_10240);
nor U10676 (N_10676,N_10071,N_10053);
nand U10677 (N_10677,N_10272,N_10142);
xor U10678 (N_10678,N_10191,N_10320);
xnor U10679 (N_10679,N_10179,N_10188);
and U10680 (N_10680,N_10383,N_10060);
and U10681 (N_10681,N_10011,N_10232);
nor U10682 (N_10682,N_10101,N_10415);
xnor U10683 (N_10683,N_10443,N_10127);
nor U10684 (N_10684,N_10035,N_10498);
or U10685 (N_10685,N_10112,N_10493);
or U10686 (N_10686,N_10120,N_10222);
nand U10687 (N_10687,N_10064,N_10491);
nand U10688 (N_10688,N_10261,N_10181);
xor U10689 (N_10689,N_10464,N_10485);
and U10690 (N_10690,N_10422,N_10077);
and U10691 (N_10691,N_10106,N_10294);
or U10692 (N_10692,N_10234,N_10212);
nor U10693 (N_10693,N_10009,N_10109);
nor U10694 (N_10694,N_10004,N_10432);
or U10695 (N_10695,N_10267,N_10483);
and U10696 (N_10696,N_10040,N_10068);
and U10697 (N_10697,N_10151,N_10404);
nor U10698 (N_10698,N_10344,N_10163);
nand U10699 (N_10699,N_10442,N_10030);
and U10700 (N_10700,N_10448,N_10255);
and U10701 (N_10701,N_10162,N_10072);
nand U10702 (N_10702,N_10183,N_10466);
or U10703 (N_10703,N_10387,N_10038);
nor U10704 (N_10704,N_10275,N_10353);
xnor U10705 (N_10705,N_10467,N_10429);
nand U10706 (N_10706,N_10006,N_10027);
and U10707 (N_10707,N_10057,N_10336);
or U10708 (N_10708,N_10246,N_10050);
nand U10709 (N_10709,N_10487,N_10259);
and U10710 (N_10710,N_10100,N_10022);
or U10711 (N_10711,N_10089,N_10469);
nor U10712 (N_10712,N_10427,N_10245);
or U10713 (N_10713,N_10066,N_10492);
nor U10714 (N_10714,N_10239,N_10450);
nand U10715 (N_10715,N_10428,N_10236);
and U10716 (N_10716,N_10073,N_10416);
nand U10717 (N_10717,N_10247,N_10494);
nor U10718 (N_10718,N_10063,N_10069);
or U10719 (N_10719,N_10087,N_10145);
nand U10720 (N_10720,N_10266,N_10342);
or U10721 (N_10721,N_10459,N_10028);
nand U10722 (N_10722,N_10094,N_10251);
nand U10723 (N_10723,N_10436,N_10160);
or U10724 (N_10724,N_10025,N_10026);
nor U10725 (N_10725,N_10475,N_10457);
and U10726 (N_10726,N_10134,N_10489);
nand U10727 (N_10727,N_10473,N_10349);
and U10728 (N_10728,N_10388,N_10369);
and U10729 (N_10729,N_10350,N_10252);
nand U10730 (N_10730,N_10048,N_10343);
or U10731 (N_10731,N_10165,N_10042);
or U10732 (N_10732,N_10417,N_10455);
and U10733 (N_10733,N_10217,N_10111);
nand U10734 (N_10734,N_10413,N_10386);
or U10735 (N_10735,N_10052,N_10091);
and U10736 (N_10736,N_10329,N_10389);
or U10737 (N_10737,N_10211,N_10133);
nand U10738 (N_10738,N_10419,N_10287);
xnor U10739 (N_10739,N_10373,N_10304);
nor U10740 (N_10740,N_10172,N_10478);
nand U10741 (N_10741,N_10241,N_10327);
nor U10742 (N_10742,N_10023,N_10262);
or U10743 (N_10743,N_10352,N_10144);
or U10744 (N_10744,N_10117,N_10435);
nor U10745 (N_10745,N_10005,N_10215);
nand U10746 (N_10746,N_10463,N_10458);
or U10747 (N_10747,N_10056,N_10332);
or U10748 (N_10748,N_10319,N_10453);
nand U10749 (N_10749,N_10002,N_10468);
or U10750 (N_10750,N_10039,N_10025);
xor U10751 (N_10751,N_10243,N_10412);
and U10752 (N_10752,N_10301,N_10019);
nand U10753 (N_10753,N_10068,N_10413);
and U10754 (N_10754,N_10312,N_10471);
nand U10755 (N_10755,N_10200,N_10441);
nor U10756 (N_10756,N_10422,N_10234);
or U10757 (N_10757,N_10027,N_10026);
nor U10758 (N_10758,N_10257,N_10478);
or U10759 (N_10759,N_10126,N_10147);
and U10760 (N_10760,N_10394,N_10326);
or U10761 (N_10761,N_10023,N_10149);
nand U10762 (N_10762,N_10304,N_10106);
and U10763 (N_10763,N_10138,N_10080);
and U10764 (N_10764,N_10010,N_10321);
nor U10765 (N_10765,N_10099,N_10120);
nand U10766 (N_10766,N_10490,N_10133);
nor U10767 (N_10767,N_10158,N_10159);
and U10768 (N_10768,N_10420,N_10135);
nor U10769 (N_10769,N_10256,N_10335);
nor U10770 (N_10770,N_10342,N_10026);
nor U10771 (N_10771,N_10017,N_10002);
or U10772 (N_10772,N_10061,N_10453);
nor U10773 (N_10773,N_10492,N_10082);
nand U10774 (N_10774,N_10127,N_10165);
or U10775 (N_10775,N_10290,N_10132);
nand U10776 (N_10776,N_10474,N_10166);
nor U10777 (N_10777,N_10377,N_10025);
and U10778 (N_10778,N_10402,N_10026);
nand U10779 (N_10779,N_10206,N_10159);
nand U10780 (N_10780,N_10312,N_10271);
nor U10781 (N_10781,N_10049,N_10429);
or U10782 (N_10782,N_10045,N_10499);
nor U10783 (N_10783,N_10412,N_10459);
and U10784 (N_10784,N_10466,N_10469);
and U10785 (N_10785,N_10472,N_10174);
or U10786 (N_10786,N_10052,N_10441);
nand U10787 (N_10787,N_10256,N_10328);
nor U10788 (N_10788,N_10027,N_10401);
nor U10789 (N_10789,N_10016,N_10014);
nor U10790 (N_10790,N_10232,N_10336);
and U10791 (N_10791,N_10064,N_10468);
nand U10792 (N_10792,N_10003,N_10110);
or U10793 (N_10793,N_10238,N_10189);
nand U10794 (N_10794,N_10409,N_10099);
or U10795 (N_10795,N_10332,N_10250);
nand U10796 (N_10796,N_10462,N_10248);
and U10797 (N_10797,N_10041,N_10298);
nand U10798 (N_10798,N_10101,N_10000);
nand U10799 (N_10799,N_10078,N_10290);
or U10800 (N_10800,N_10028,N_10200);
nor U10801 (N_10801,N_10123,N_10098);
nand U10802 (N_10802,N_10387,N_10215);
xor U10803 (N_10803,N_10016,N_10167);
or U10804 (N_10804,N_10118,N_10057);
nor U10805 (N_10805,N_10224,N_10123);
nor U10806 (N_10806,N_10049,N_10428);
and U10807 (N_10807,N_10463,N_10077);
nor U10808 (N_10808,N_10490,N_10393);
or U10809 (N_10809,N_10096,N_10061);
nor U10810 (N_10810,N_10389,N_10450);
nand U10811 (N_10811,N_10325,N_10002);
and U10812 (N_10812,N_10071,N_10263);
nand U10813 (N_10813,N_10130,N_10312);
nand U10814 (N_10814,N_10176,N_10012);
and U10815 (N_10815,N_10134,N_10060);
or U10816 (N_10816,N_10230,N_10274);
and U10817 (N_10817,N_10220,N_10419);
or U10818 (N_10818,N_10242,N_10285);
nor U10819 (N_10819,N_10087,N_10170);
or U10820 (N_10820,N_10485,N_10295);
nand U10821 (N_10821,N_10113,N_10365);
or U10822 (N_10822,N_10375,N_10422);
nor U10823 (N_10823,N_10167,N_10326);
nor U10824 (N_10824,N_10199,N_10286);
nor U10825 (N_10825,N_10348,N_10109);
xnor U10826 (N_10826,N_10039,N_10351);
nand U10827 (N_10827,N_10469,N_10474);
nor U10828 (N_10828,N_10043,N_10060);
and U10829 (N_10829,N_10323,N_10441);
nand U10830 (N_10830,N_10315,N_10406);
nand U10831 (N_10831,N_10345,N_10048);
and U10832 (N_10832,N_10122,N_10362);
nand U10833 (N_10833,N_10274,N_10232);
and U10834 (N_10834,N_10185,N_10385);
nor U10835 (N_10835,N_10011,N_10352);
or U10836 (N_10836,N_10259,N_10112);
or U10837 (N_10837,N_10063,N_10169);
nand U10838 (N_10838,N_10310,N_10009);
or U10839 (N_10839,N_10445,N_10099);
or U10840 (N_10840,N_10409,N_10195);
and U10841 (N_10841,N_10198,N_10171);
and U10842 (N_10842,N_10027,N_10111);
or U10843 (N_10843,N_10088,N_10283);
nand U10844 (N_10844,N_10374,N_10406);
and U10845 (N_10845,N_10138,N_10242);
nor U10846 (N_10846,N_10449,N_10408);
and U10847 (N_10847,N_10081,N_10196);
nand U10848 (N_10848,N_10186,N_10035);
nor U10849 (N_10849,N_10254,N_10451);
and U10850 (N_10850,N_10476,N_10004);
nand U10851 (N_10851,N_10095,N_10242);
and U10852 (N_10852,N_10477,N_10107);
and U10853 (N_10853,N_10060,N_10059);
or U10854 (N_10854,N_10295,N_10337);
nor U10855 (N_10855,N_10113,N_10227);
xor U10856 (N_10856,N_10492,N_10485);
nand U10857 (N_10857,N_10017,N_10147);
and U10858 (N_10858,N_10129,N_10205);
xnor U10859 (N_10859,N_10268,N_10043);
nor U10860 (N_10860,N_10075,N_10454);
nor U10861 (N_10861,N_10364,N_10344);
or U10862 (N_10862,N_10182,N_10224);
nand U10863 (N_10863,N_10448,N_10246);
nand U10864 (N_10864,N_10224,N_10485);
nand U10865 (N_10865,N_10067,N_10080);
nor U10866 (N_10866,N_10319,N_10309);
or U10867 (N_10867,N_10078,N_10416);
nor U10868 (N_10868,N_10235,N_10101);
xor U10869 (N_10869,N_10132,N_10322);
and U10870 (N_10870,N_10206,N_10210);
nor U10871 (N_10871,N_10010,N_10049);
nand U10872 (N_10872,N_10398,N_10354);
xor U10873 (N_10873,N_10295,N_10369);
or U10874 (N_10874,N_10029,N_10074);
or U10875 (N_10875,N_10108,N_10350);
or U10876 (N_10876,N_10254,N_10319);
nor U10877 (N_10877,N_10373,N_10394);
and U10878 (N_10878,N_10317,N_10106);
or U10879 (N_10879,N_10319,N_10292);
or U10880 (N_10880,N_10298,N_10246);
and U10881 (N_10881,N_10116,N_10104);
or U10882 (N_10882,N_10371,N_10307);
xor U10883 (N_10883,N_10180,N_10401);
nor U10884 (N_10884,N_10205,N_10437);
or U10885 (N_10885,N_10423,N_10221);
or U10886 (N_10886,N_10001,N_10486);
or U10887 (N_10887,N_10143,N_10496);
and U10888 (N_10888,N_10444,N_10005);
and U10889 (N_10889,N_10115,N_10343);
or U10890 (N_10890,N_10043,N_10492);
nand U10891 (N_10891,N_10385,N_10153);
and U10892 (N_10892,N_10152,N_10470);
nor U10893 (N_10893,N_10409,N_10214);
nor U10894 (N_10894,N_10309,N_10392);
or U10895 (N_10895,N_10361,N_10351);
nand U10896 (N_10896,N_10400,N_10184);
nand U10897 (N_10897,N_10367,N_10209);
nand U10898 (N_10898,N_10097,N_10075);
and U10899 (N_10899,N_10411,N_10144);
nand U10900 (N_10900,N_10371,N_10106);
or U10901 (N_10901,N_10210,N_10399);
and U10902 (N_10902,N_10447,N_10165);
nor U10903 (N_10903,N_10227,N_10335);
xnor U10904 (N_10904,N_10229,N_10388);
nor U10905 (N_10905,N_10012,N_10188);
nand U10906 (N_10906,N_10286,N_10257);
xor U10907 (N_10907,N_10375,N_10496);
and U10908 (N_10908,N_10270,N_10428);
and U10909 (N_10909,N_10493,N_10005);
and U10910 (N_10910,N_10421,N_10487);
and U10911 (N_10911,N_10217,N_10340);
nand U10912 (N_10912,N_10491,N_10134);
nor U10913 (N_10913,N_10231,N_10273);
and U10914 (N_10914,N_10486,N_10415);
nor U10915 (N_10915,N_10205,N_10229);
nor U10916 (N_10916,N_10466,N_10461);
nand U10917 (N_10917,N_10056,N_10219);
nor U10918 (N_10918,N_10194,N_10002);
or U10919 (N_10919,N_10353,N_10419);
xor U10920 (N_10920,N_10110,N_10257);
and U10921 (N_10921,N_10073,N_10261);
or U10922 (N_10922,N_10311,N_10452);
xnor U10923 (N_10923,N_10164,N_10324);
nor U10924 (N_10924,N_10109,N_10084);
and U10925 (N_10925,N_10298,N_10227);
xnor U10926 (N_10926,N_10013,N_10150);
or U10927 (N_10927,N_10456,N_10492);
or U10928 (N_10928,N_10142,N_10230);
xor U10929 (N_10929,N_10034,N_10224);
and U10930 (N_10930,N_10397,N_10165);
nor U10931 (N_10931,N_10166,N_10395);
xnor U10932 (N_10932,N_10150,N_10092);
nand U10933 (N_10933,N_10239,N_10095);
nand U10934 (N_10934,N_10127,N_10153);
xnor U10935 (N_10935,N_10079,N_10308);
nand U10936 (N_10936,N_10165,N_10100);
or U10937 (N_10937,N_10388,N_10233);
and U10938 (N_10938,N_10219,N_10365);
and U10939 (N_10939,N_10106,N_10366);
or U10940 (N_10940,N_10276,N_10232);
nand U10941 (N_10941,N_10202,N_10035);
nor U10942 (N_10942,N_10430,N_10255);
nor U10943 (N_10943,N_10235,N_10124);
nor U10944 (N_10944,N_10354,N_10468);
and U10945 (N_10945,N_10028,N_10328);
and U10946 (N_10946,N_10079,N_10210);
and U10947 (N_10947,N_10313,N_10050);
or U10948 (N_10948,N_10041,N_10424);
nor U10949 (N_10949,N_10055,N_10283);
nand U10950 (N_10950,N_10457,N_10498);
or U10951 (N_10951,N_10023,N_10371);
nand U10952 (N_10952,N_10316,N_10257);
xnor U10953 (N_10953,N_10372,N_10403);
nand U10954 (N_10954,N_10448,N_10180);
xnor U10955 (N_10955,N_10487,N_10350);
or U10956 (N_10956,N_10490,N_10173);
and U10957 (N_10957,N_10274,N_10119);
nor U10958 (N_10958,N_10034,N_10254);
or U10959 (N_10959,N_10280,N_10459);
nor U10960 (N_10960,N_10434,N_10170);
nor U10961 (N_10961,N_10379,N_10408);
and U10962 (N_10962,N_10169,N_10355);
and U10963 (N_10963,N_10036,N_10085);
and U10964 (N_10964,N_10226,N_10479);
and U10965 (N_10965,N_10474,N_10287);
nor U10966 (N_10966,N_10027,N_10476);
nor U10967 (N_10967,N_10007,N_10298);
nand U10968 (N_10968,N_10260,N_10296);
or U10969 (N_10969,N_10087,N_10213);
nor U10970 (N_10970,N_10131,N_10471);
or U10971 (N_10971,N_10168,N_10327);
nand U10972 (N_10972,N_10089,N_10201);
nand U10973 (N_10973,N_10150,N_10180);
nand U10974 (N_10974,N_10116,N_10271);
nand U10975 (N_10975,N_10156,N_10207);
or U10976 (N_10976,N_10286,N_10366);
nor U10977 (N_10977,N_10429,N_10350);
nand U10978 (N_10978,N_10285,N_10026);
xnor U10979 (N_10979,N_10443,N_10424);
nand U10980 (N_10980,N_10395,N_10468);
and U10981 (N_10981,N_10498,N_10390);
nand U10982 (N_10982,N_10292,N_10256);
xnor U10983 (N_10983,N_10390,N_10115);
xnor U10984 (N_10984,N_10427,N_10334);
or U10985 (N_10985,N_10104,N_10236);
or U10986 (N_10986,N_10249,N_10348);
and U10987 (N_10987,N_10294,N_10126);
and U10988 (N_10988,N_10086,N_10355);
nand U10989 (N_10989,N_10033,N_10428);
nand U10990 (N_10990,N_10205,N_10482);
xor U10991 (N_10991,N_10217,N_10411);
and U10992 (N_10992,N_10185,N_10120);
xnor U10993 (N_10993,N_10255,N_10461);
nand U10994 (N_10994,N_10091,N_10365);
and U10995 (N_10995,N_10284,N_10091);
nand U10996 (N_10996,N_10450,N_10347);
nand U10997 (N_10997,N_10077,N_10259);
or U10998 (N_10998,N_10023,N_10465);
nand U10999 (N_10999,N_10469,N_10017);
nor U11000 (N_11000,N_10722,N_10716);
or U11001 (N_11001,N_10618,N_10892);
and U11002 (N_11002,N_10608,N_10523);
xnor U11003 (N_11003,N_10568,N_10954);
or U11004 (N_11004,N_10729,N_10742);
and U11005 (N_11005,N_10919,N_10735);
nand U11006 (N_11006,N_10793,N_10524);
or U11007 (N_11007,N_10534,N_10656);
and U11008 (N_11008,N_10841,N_10518);
or U11009 (N_11009,N_10593,N_10748);
nor U11010 (N_11010,N_10786,N_10563);
and U11011 (N_11011,N_10631,N_10611);
and U11012 (N_11012,N_10548,N_10941);
nand U11013 (N_11013,N_10779,N_10581);
nor U11014 (N_11014,N_10997,N_10702);
and U11015 (N_11015,N_10605,N_10638);
nand U11016 (N_11016,N_10528,N_10531);
or U11017 (N_11017,N_10945,N_10637);
and U11018 (N_11018,N_10507,N_10942);
nand U11019 (N_11019,N_10699,N_10595);
and U11020 (N_11020,N_10944,N_10519);
nor U11021 (N_11021,N_10923,N_10741);
and U11022 (N_11022,N_10759,N_10824);
nor U11023 (N_11023,N_10577,N_10926);
and U11024 (N_11024,N_10774,N_10603);
xnor U11025 (N_11025,N_10682,N_10701);
and U11026 (N_11026,N_10922,N_10693);
or U11027 (N_11027,N_10683,N_10935);
xor U11028 (N_11028,N_10773,N_10738);
nand U11029 (N_11029,N_10842,N_10908);
nor U11030 (N_11030,N_10753,N_10799);
nand U11031 (N_11031,N_10585,N_10902);
xor U11032 (N_11032,N_10540,N_10517);
nor U11033 (N_11033,N_10878,N_10732);
nand U11034 (N_11034,N_10614,N_10879);
nor U11035 (N_11035,N_10943,N_10950);
nor U11036 (N_11036,N_10996,N_10870);
or U11037 (N_11037,N_10622,N_10809);
nand U11038 (N_11038,N_10733,N_10711);
or U11039 (N_11039,N_10916,N_10578);
or U11040 (N_11040,N_10526,N_10994);
or U11041 (N_11041,N_10600,N_10851);
and U11042 (N_11042,N_10802,N_10616);
xor U11043 (N_11043,N_10867,N_10790);
nand U11044 (N_11044,N_10658,N_10887);
and U11045 (N_11045,N_10521,N_10921);
nand U11046 (N_11046,N_10731,N_10740);
or U11047 (N_11047,N_10647,N_10552);
or U11048 (N_11048,N_10549,N_10963);
or U11049 (N_11049,N_10789,N_10760);
nand U11050 (N_11050,N_10932,N_10826);
and U11051 (N_11051,N_10896,N_10956);
and U11052 (N_11052,N_10884,N_10686);
xnor U11053 (N_11053,N_10990,N_10610);
or U11054 (N_11054,N_10697,N_10857);
nor U11055 (N_11055,N_10906,N_10854);
nor U11056 (N_11056,N_10527,N_10642);
nor U11057 (N_11057,N_10972,N_10558);
nand U11058 (N_11058,N_10883,N_10734);
and U11059 (N_11059,N_10776,N_10727);
and U11060 (N_11060,N_10565,N_10508);
and U11061 (N_11061,N_10560,N_10666);
or U11062 (N_11062,N_10951,N_10708);
nor U11063 (N_11063,N_10920,N_10624);
or U11064 (N_11064,N_10959,N_10743);
nand U11065 (N_11065,N_10901,N_10690);
nor U11066 (N_11066,N_10859,N_10978);
nor U11067 (N_11067,N_10844,N_10678);
and U11068 (N_11068,N_10939,N_10555);
nand U11069 (N_11069,N_10787,N_10962);
nor U11070 (N_11070,N_10849,N_10582);
nor U11071 (N_11071,N_10709,N_10537);
xnor U11072 (N_11072,N_10977,N_10781);
or U11073 (N_11073,N_10783,N_10900);
or U11074 (N_11074,N_10737,N_10609);
or U11075 (N_11075,N_10506,N_10876);
and U11076 (N_11076,N_10866,N_10655);
or U11077 (N_11077,N_10937,N_10672);
nand U11078 (N_11078,N_10691,N_10795);
nor U11079 (N_11079,N_10712,N_10777);
nor U11080 (N_11080,N_10931,N_10522);
nor U11081 (N_11081,N_10520,N_10668);
or U11082 (N_11082,N_10752,N_10834);
nand U11083 (N_11083,N_10848,N_10723);
nor U11084 (N_11084,N_10910,N_10986);
nand U11085 (N_11085,N_10669,N_10514);
or U11086 (N_11086,N_10830,N_10971);
nor U11087 (N_11087,N_10653,N_10645);
or U11088 (N_11088,N_10904,N_10553);
nor U11089 (N_11089,N_10832,N_10586);
nor U11090 (N_11090,N_10794,N_10685);
and U11091 (N_11091,N_10805,N_10596);
or U11092 (N_11092,N_10505,N_10704);
or U11093 (N_11093,N_10829,N_10784);
nand U11094 (N_11094,N_10980,N_10957);
nor U11095 (N_11095,N_10765,N_10684);
or U11096 (N_11096,N_10648,N_10652);
and U11097 (N_11097,N_10969,N_10736);
nand U11098 (N_11098,N_10858,N_10989);
nor U11099 (N_11099,N_10911,N_10688);
and U11100 (N_11100,N_10974,N_10594);
or U11101 (N_11101,N_10579,N_10775);
nand U11102 (N_11102,N_10659,N_10635);
or U11103 (N_11103,N_10967,N_10681);
and U11104 (N_11104,N_10649,N_10903);
and U11105 (N_11105,N_10907,N_10509);
nor U11106 (N_11106,N_10675,N_10880);
xnor U11107 (N_11107,N_10564,N_10751);
and U11108 (N_11108,N_10890,N_10885);
xnor U11109 (N_11109,N_10550,N_10807);
nand U11110 (N_11110,N_10864,N_10717);
xor U11111 (N_11111,N_10575,N_10891);
or U11112 (N_11112,N_10623,N_10918);
nor U11113 (N_11113,N_10503,N_10513);
nor U11114 (N_11114,N_10592,N_10515);
or U11115 (N_11115,N_10964,N_10730);
xnor U11116 (N_11116,N_10501,N_10557);
or U11117 (N_11117,N_10650,N_10914);
and U11118 (N_11118,N_10539,N_10567);
or U11119 (N_11119,N_10821,N_10689);
or U11120 (N_11120,N_10543,N_10991);
nand U11121 (N_11121,N_10847,N_10780);
nand U11122 (N_11122,N_10671,N_10569);
and U11123 (N_11123,N_10670,N_10580);
nand U11124 (N_11124,N_10825,N_10516);
and U11125 (N_11125,N_10952,N_10687);
or U11126 (N_11126,N_10813,N_10823);
or U11127 (N_11127,N_10798,N_10835);
nand U11128 (N_11128,N_10541,N_10895);
and U11129 (N_11129,N_10547,N_10551);
nand U11130 (N_11130,N_10763,N_10772);
or U11131 (N_11131,N_10767,N_10597);
xnor U11132 (N_11132,N_10993,N_10960);
and U11133 (N_11133,N_10888,N_10633);
xnor U11134 (N_11134,N_10694,N_10984);
nand U11135 (N_11135,N_10801,N_10961);
nor U11136 (N_11136,N_10874,N_10816);
nand U11137 (N_11137,N_10927,N_10634);
nor U11138 (N_11138,N_10948,N_10654);
or U11139 (N_11139,N_10756,N_10791);
nor U11140 (N_11140,N_10946,N_10629);
and U11141 (N_11141,N_10981,N_10706);
or U11142 (N_11142,N_10815,N_10949);
and U11143 (N_11143,N_10856,N_10894);
xor U11144 (N_11144,N_10651,N_10640);
nor U11145 (N_11145,N_10863,N_10797);
or U11146 (N_11146,N_10535,N_10725);
nand U11147 (N_11147,N_10833,N_10837);
nor U11148 (N_11148,N_10881,N_10889);
or U11149 (N_11149,N_10800,N_10584);
nand U11150 (N_11150,N_10840,N_10719);
nand U11151 (N_11151,N_10607,N_10983);
xor U11152 (N_11152,N_10680,N_10529);
and U11153 (N_11153,N_10992,N_10976);
and U11154 (N_11154,N_10912,N_10836);
nand U11155 (N_11155,N_10757,N_10715);
or U11156 (N_11156,N_10796,N_10755);
or U11157 (N_11157,N_10749,N_10764);
nand U11158 (N_11158,N_10808,N_10999);
or U11159 (N_11159,N_10570,N_10818);
nor U11160 (N_11160,N_10975,N_10530);
nand U11161 (N_11161,N_10615,N_10566);
nor U11162 (N_11162,N_10855,N_10546);
and U11163 (N_11163,N_10696,N_10814);
and U11164 (N_11164,N_10728,N_10532);
nor U11165 (N_11165,N_10822,N_10679);
nor U11166 (N_11166,N_10810,N_10724);
nand U11167 (N_11167,N_10613,N_10533);
and U11168 (N_11168,N_10591,N_10925);
nor U11169 (N_11169,N_10574,N_10771);
nand U11170 (N_11170,N_10940,N_10747);
nor U11171 (N_11171,N_10871,N_10620);
nand U11172 (N_11172,N_10739,N_10502);
nand U11173 (N_11173,N_10663,N_10559);
nand U11174 (N_11174,N_10510,N_10571);
and U11175 (N_11175,N_10998,N_10869);
and U11176 (N_11176,N_10745,N_10831);
or U11177 (N_11177,N_10692,N_10525);
and U11178 (N_11178,N_10965,N_10710);
nand U11179 (N_11179,N_10758,N_10588);
or U11180 (N_11180,N_10636,N_10665);
and U11181 (N_11181,N_10713,N_10554);
nand U11182 (N_11182,N_10601,N_10556);
or U11183 (N_11183,N_10820,N_10700);
nor U11184 (N_11184,N_10958,N_10707);
and U11185 (N_11185,N_10598,N_10966);
nor U11186 (N_11186,N_10660,N_10632);
and U11187 (N_11187,N_10627,N_10504);
and U11188 (N_11188,N_10933,N_10644);
xor U11189 (N_11189,N_10676,N_10843);
or U11190 (N_11190,N_10806,N_10968);
nor U11191 (N_11191,N_10590,N_10803);
nor U11192 (N_11192,N_10512,N_10817);
and U11193 (N_11193,N_10893,N_10664);
nor U11194 (N_11194,N_10750,N_10587);
or U11195 (N_11195,N_10852,N_10985);
xor U11196 (N_11196,N_10953,N_10938);
nand U11197 (N_11197,N_10630,N_10917);
and U11198 (N_11198,N_10838,N_10877);
or U11199 (N_11199,N_10617,N_10726);
and U11200 (N_11200,N_10827,N_10905);
nor U11201 (N_11201,N_10639,N_10705);
nand U11202 (N_11202,N_10754,N_10761);
or U11203 (N_11203,N_10899,N_10673);
or U11204 (N_11204,N_10657,N_10536);
and U11205 (N_11205,N_10970,N_10850);
nand U11206 (N_11206,N_10511,N_10861);
or U11207 (N_11207,N_10770,N_10778);
or U11208 (N_11208,N_10846,N_10619);
nand U11209 (N_11209,N_10674,N_10839);
and U11210 (N_11210,N_10929,N_10930);
or U11211 (N_11211,N_10788,N_10572);
or U11212 (N_11212,N_10987,N_10979);
or U11213 (N_11213,N_10819,N_10898);
and U11214 (N_11214,N_10545,N_10576);
nand U11215 (N_11215,N_10544,N_10853);
or U11216 (N_11216,N_10661,N_10860);
and U11217 (N_11217,N_10982,N_10875);
and U11218 (N_11218,N_10886,N_10625);
nand U11219 (N_11219,N_10955,N_10538);
xor U11220 (N_11220,N_10621,N_10868);
and U11221 (N_11221,N_10718,N_10720);
or U11222 (N_11222,N_10612,N_10909);
and U11223 (N_11223,N_10862,N_10882);
nor U11224 (N_11224,N_10845,N_10573);
or U11225 (N_11225,N_10928,N_10604);
nor U11226 (N_11226,N_10973,N_10606);
or U11227 (N_11227,N_10913,N_10599);
nand U11228 (N_11228,N_10602,N_10561);
nand U11229 (N_11229,N_10628,N_10915);
nand U11230 (N_11230,N_10643,N_10721);
xor U11231 (N_11231,N_10936,N_10626);
and U11232 (N_11232,N_10714,N_10703);
nand U11233 (N_11233,N_10924,N_10589);
or U11234 (N_11234,N_10947,N_10873);
nor U11235 (N_11235,N_10746,N_10500);
or U11236 (N_11236,N_10695,N_10804);
nand U11237 (N_11237,N_10812,N_10811);
nor U11238 (N_11238,N_10542,N_10785);
and U11239 (N_11239,N_10762,N_10934);
xor U11240 (N_11240,N_10768,N_10865);
nor U11241 (N_11241,N_10698,N_10677);
or U11242 (N_11242,N_10792,N_10995);
or U11243 (N_11243,N_10782,N_10744);
and U11244 (N_11244,N_10872,N_10897);
nand U11245 (N_11245,N_10828,N_10988);
nor U11246 (N_11246,N_10766,N_10562);
nand U11247 (N_11247,N_10583,N_10769);
nor U11248 (N_11248,N_10641,N_10662);
nand U11249 (N_11249,N_10667,N_10646);
nor U11250 (N_11250,N_10878,N_10945);
or U11251 (N_11251,N_10821,N_10611);
and U11252 (N_11252,N_10787,N_10791);
and U11253 (N_11253,N_10677,N_10522);
or U11254 (N_11254,N_10835,N_10986);
nand U11255 (N_11255,N_10715,N_10703);
and U11256 (N_11256,N_10687,N_10516);
and U11257 (N_11257,N_10666,N_10522);
nand U11258 (N_11258,N_10856,N_10959);
nor U11259 (N_11259,N_10766,N_10763);
nor U11260 (N_11260,N_10929,N_10823);
xnor U11261 (N_11261,N_10829,N_10965);
nand U11262 (N_11262,N_10533,N_10549);
or U11263 (N_11263,N_10716,N_10862);
and U11264 (N_11264,N_10860,N_10574);
nand U11265 (N_11265,N_10529,N_10933);
xnor U11266 (N_11266,N_10884,N_10814);
nor U11267 (N_11267,N_10687,N_10984);
and U11268 (N_11268,N_10957,N_10772);
nor U11269 (N_11269,N_10691,N_10686);
nand U11270 (N_11270,N_10726,N_10914);
xor U11271 (N_11271,N_10578,N_10655);
nand U11272 (N_11272,N_10682,N_10611);
nand U11273 (N_11273,N_10958,N_10786);
nand U11274 (N_11274,N_10734,N_10716);
and U11275 (N_11275,N_10671,N_10682);
nor U11276 (N_11276,N_10674,N_10969);
and U11277 (N_11277,N_10824,N_10867);
xnor U11278 (N_11278,N_10524,N_10676);
nor U11279 (N_11279,N_10868,N_10528);
nand U11280 (N_11280,N_10885,N_10748);
xnor U11281 (N_11281,N_10770,N_10913);
nor U11282 (N_11282,N_10572,N_10674);
xor U11283 (N_11283,N_10515,N_10537);
nor U11284 (N_11284,N_10935,N_10829);
or U11285 (N_11285,N_10500,N_10734);
nand U11286 (N_11286,N_10870,N_10871);
nand U11287 (N_11287,N_10538,N_10926);
nand U11288 (N_11288,N_10988,N_10555);
or U11289 (N_11289,N_10684,N_10902);
or U11290 (N_11290,N_10586,N_10507);
xnor U11291 (N_11291,N_10936,N_10852);
or U11292 (N_11292,N_10641,N_10917);
and U11293 (N_11293,N_10636,N_10544);
and U11294 (N_11294,N_10526,N_10955);
nand U11295 (N_11295,N_10593,N_10940);
or U11296 (N_11296,N_10867,N_10579);
nand U11297 (N_11297,N_10813,N_10546);
xnor U11298 (N_11298,N_10585,N_10500);
or U11299 (N_11299,N_10872,N_10762);
nand U11300 (N_11300,N_10691,N_10713);
nor U11301 (N_11301,N_10646,N_10575);
nand U11302 (N_11302,N_10831,N_10931);
nor U11303 (N_11303,N_10615,N_10921);
and U11304 (N_11304,N_10963,N_10831);
nor U11305 (N_11305,N_10825,N_10733);
nor U11306 (N_11306,N_10686,N_10748);
nor U11307 (N_11307,N_10979,N_10598);
and U11308 (N_11308,N_10997,N_10976);
or U11309 (N_11309,N_10692,N_10993);
nor U11310 (N_11310,N_10562,N_10713);
nand U11311 (N_11311,N_10959,N_10732);
xnor U11312 (N_11312,N_10986,N_10837);
nand U11313 (N_11313,N_10997,N_10915);
nand U11314 (N_11314,N_10903,N_10909);
nand U11315 (N_11315,N_10881,N_10560);
and U11316 (N_11316,N_10691,N_10886);
or U11317 (N_11317,N_10690,N_10931);
nand U11318 (N_11318,N_10595,N_10508);
or U11319 (N_11319,N_10562,N_10676);
xnor U11320 (N_11320,N_10633,N_10536);
nand U11321 (N_11321,N_10513,N_10816);
nor U11322 (N_11322,N_10784,N_10912);
and U11323 (N_11323,N_10658,N_10800);
and U11324 (N_11324,N_10521,N_10774);
nand U11325 (N_11325,N_10692,N_10877);
or U11326 (N_11326,N_10828,N_10709);
or U11327 (N_11327,N_10996,N_10558);
xor U11328 (N_11328,N_10649,N_10913);
nand U11329 (N_11329,N_10692,N_10509);
nor U11330 (N_11330,N_10830,N_10562);
nor U11331 (N_11331,N_10912,N_10685);
xnor U11332 (N_11332,N_10902,N_10732);
nand U11333 (N_11333,N_10820,N_10728);
nand U11334 (N_11334,N_10526,N_10976);
xor U11335 (N_11335,N_10547,N_10569);
and U11336 (N_11336,N_10509,N_10950);
or U11337 (N_11337,N_10737,N_10602);
nand U11338 (N_11338,N_10567,N_10611);
or U11339 (N_11339,N_10911,N_10589);
nor U11340 (N_11340,N_10986,N_10850);
or U11341 (N_11341,N_10780,N_10946);
and U11342 (N_11342,N_10680,N_10894);
nor U11343 (N_11343,N_10718,N_10645);
or U11344 (N_11344,N_10643,N_10884);
or U11345 (N_11345,N_10935,N_10645);
or U11346 (N_11346,N_10617,N_10636);
or U11347 (N_11347,N_10849,N_10673);
or U11348 (N_11348,N_10598,N_10852);
and U11349 (N_11349,N_10765,N_10970);
and U11350 (N_11350,N_10787,N_10597);
and U11351 (N_11351,N_10973,N_10626);
or U11352 (N_11352,N_10564,N_10849);
and U11353 (N_11353,N_10520,N_10604);
nor U11354 (N_11354,N_10568,N_10891);
xor U11355 (N_11355,N_10809,N_10981);
xnor U11356 (N_11356,N_10571,N_10748);
or U11357 (N_11357,N_10536,N_10629);
nand U11358 (N_11358,N_10536,N_10731);
or U11359 (N_11359,N_10654,N_10698);
nor U11360 (N_11360,N_10736,N_10597);
nor U11361 (N_11361,N_10673,N_10871);
and U11362 (N_11362,N_10616,N_10950);
xnor U11363 (N_11363,N_10619,N_10765);
nor U11364 (N_11364,N_10766,N_10857);
nor U11365 (N_11365,N_10983,N_10553);
nand U11366 (N_11366,N_10612,N_10633);
nand U11367 (N_11367,N_10605,N_10701);
or U11368 (N_11368,N_10608,N_10646);
or U11369 (N_11369,N_10709,N_10793);
xor U11370 (N_11370,N_10554,N_10823);
xnor U11371 (N_11371,N_10519,N_10629);
nor U11372 (N_11372,N_10648,N_10931);
nand U11373 (N_11373,N_10933,N_10707);
and U11374 (N_11374,N_10610,N_10675);
or U11375 (N_11375,N_10983,N_10771);
and U11376 (N_11376,N_10718,N_10979);
nor U11377 (N_11377,N_10692,N_10893);
nand U11378 (N_11378,N_10505,N_10730);
nor U11379 (N_11379,N_10545,N_10569);
or U11380 (N_11380,N_10763,N_10827);
nor U11381 (N_11381,N_10700,N_10534);
or U11382 (N_11382,N_10526,N_10715);
nand U11383 (N_11383,N_10541,N_10990);
or U11384 (N_11384,N_10997,N_10758);
or U11385 (N_11385,N_10796,N_10586);
nand U11386 (N_11386,N_10913,N_10800);
xnor U11387 (N_11387,N_10735,N_10905);
and U11388 (N_11388,N_10911,N_10794);
or U11389 (N_11389,N_10871,N_10817);
or U11390 (N_11390,N_10881,N_10719);
nor U11391 (N_11391,N_10747,N_10779);
and U11392 (N_11392,N_10833,N_10517);
nand U11393 (N_11393,N_10780,N_10901);
nor U11394 (N_11394,N_10633,N_10501);
or U11395 (N_11395,N_10905,N_10618);
xor U11396 (N_11396,N_10665,N_10608);
and U11397 (N_11397,N_10777,N_10811);
or U11398 (N_11398,N_10827,N_10745);
nor U11399 (N_11399,N_10516,N_10588);
nor U11400 (N_11400,N_10682,N_10704);
nor U11401 (N_11401,N_10995,N_10968);
and U11402 (N_11402,N_10793,N_10521);
nor U11403 (N_11403,N_10875,N_10915);
and U11404 (N_11404,N_10687,N_10639);
xnor U11405 (N_11405,N_10549,N_10986);
nand U11406 (N_11406,N_10969,N_10700);
nor U11407 (N_11407,N_10664,N_10723);
nor U11408 (N_11408,N_10925,N_10755);
and U11409 (N_11409,N_10743,N_10776);
nor U11410 (N_11410,N_10573,N_10905);
and U11411 (N_11411,N_10583,N_10831);
and U11412 (N_11412,N_10708,N_10776);
nor U11413 (N_11413,N_10678,N_10917);
or U11414 (N_11414,N_10727,N_10561);
and U11415 (N_11415,N_10775,N_10610);
nand U11416 (N_11416,N_10978,N_10710);
nand U11417 (N_11417,N_10535,N_10758);
nand U11418 (N_11418,N_10937,N_10882);
and U11419 (N_11419,N_10565,N_10852);
nor U11420 (N_11420,N_10661,N_10761);
or U11421 (N_11421,N_10877,N_10991);
and U11422 (N_11422,N_10590,N_10860);
nand U11423 (N_11423,N_10804,N_10541);
or U11424 (N_11424,N_10833,N_10721);
or U11425 (N_11425,N_10847,N_10757);
and U11426 (N_11426,N_10620,N_10880);
and U11427 (N_11427,N_10810,N_10830);
nor U11428 (N_11428,N_10621,N_10569);
and U11429 (N_11429,N_10702,N_10663);
xnor U11430 (N_11430,N_10647,N_10778);
or U11431 (N_11431,N_10700,N_10927);
and U11432 (N_11432,N_10936,N_10742);
or U11433 (N_11433,N_10721,N_10611);
or U11434 (N_11434,N_10853,N_10904);
or U11435 (N_11435,N_10834,N_10646);
nand U11436 (N_11436,N_10773,N_10701);
and U11437 (N_11437,N_10800,N_10662);
nand U11438 (N_11438,N_10896,N_10874);
or U11439 (N_11439,N_10770,N_10572);
nor U11440 (N_11440,N_10825,N_10590);
nor U11441 (N_11441,N_10591,N_10687);
and U11442 (N_11442,N_10725,N_10510);
and U11443 (N_11443,N_10720,N_10997);
or U11444 (N_11444,N_10509,N_10873);
nand U11445 (N_11445,N_10639,N_10901);
nor U11446 (N_11446,N_10592,N_10783);
or U11447 (N_11447,N_10868,N_10893);
and U11448 (N_11448,N_10615,N_10798);
nand U11449 (N_11449,N_10895,N_10842);
nand U11450 (N_11450,N_10837,N_10850);
nor U11451 (N_11451,N_10999,N_10987);
or U11452 (N_11452,N_10576,N_10804);
or U11453 (N_11453,N_10536,N_10701);
nand U11454 (N_11454,N_10636,N_10997);
nor U11455 (N_11455,N_10603,N_10990);
or U11456 (N_11456,N_10751,N_10827);
nand U11457 (N_11457,N_10503,N_10879);
or U11458 (N_11458,N_10500,N_10655);
or U11459 (N_11459,N_10973,N_10635);
nand U11460 (N_11460,N_10750,N_10973);
and U11461 (N_11461,N_10778,N_10757);
nand U11462 (N_11462,N_10826,N_10891);
xnor U11463 (N_11463,N_10638,N_10899);
nor U11464 (N_11464,N_10550,N_10636);
or U11465 (N_11465,N_10568,N_10913);
or U11466 (N_11466,N_10665,N_10959);
or U11467 (N_11467,N_10776,N_10967);
and U11468 (N_11468,N_10573,N_10947);
and U11469 (N_11469,N_10934,N_10564);
xor U11470 (N_11470,N_10535,N_10501);
nor U11471 (N_11471,N_10938,N_10734);
or U11472 (N_11472,N_10526,N_10759);
and U11473 (N_11473,N_10726,N_10608);
or U11474 (N_11474,N_10839,N_10508);
nand U11475 (N_11475,N_10627,N_10560);
xor U11476 (N_11476,N_10803,N_10881);
nor U11477 (N_11477,N_10610,N_10934);
and U11478 (N_11478,N_10771,N_10510);
and U11479 (N_11479,N_10774,N_10963);
or U11480 (N_11480,N_10963,N_10501);
nor U11481 (N_11481,N_10962,N_10632);
nor U11482 (N_11482,N_10706,N_10516);
and U11483 (N_11483,N_10727,N_10684);
and U11484 (N_11484,N_10973,N_10703);
or U11485 (N_11485,N_10949,N_10688);
nand U11486 (N_11486,N_10893,N_10682);
xnor U11487 (N_11487,N_10576,N_10933);
or U11488 (N_11488,N_10601,N_10937);
and U11489 (N_11489,N_10979,N_10933);
and U11490 (N_11490,N_10948,N_10616);
nor U11491 (N_11491,N_10827,N_10585);
nand U11492 (N_11492,N_10832,N_10880);
and U11493 (N_11493,N_10921,N_10531);
and U11494 (N_11494,N_10743,N_10920);
nand U11495 (N_11495,N_10791,N_10979);
and U11496 (N_11496,N_10587,N_10922);
and U11497 (N_11497,N_10666,N_10918);
nand U11498 (N_11498,N_10832,N_10947);
or U11499 (N_11499,N_10846,N_10951);
or U11500 (N_11500,N_11219,N_11379);
and U11501 (N_11501,N_11481,N_11146);
and U11502 (N_11502,N_11380,N_11210);
or U11503 (N_11503,N_11207,N_11047);
nand U11504 (N_11504,N_11319,N_11054);
nand U11505 (N_11505,N_11203,N_11104);
nand U11506 (N_11506,N_11034,N_11198);
nand U11507 (N_11507,N_11342,N_11193);
nand U11508 (N_11508,N_11249,N_11488);
xor U11509 (N_11509,N_11429,N_11329);
nor U11510 (N_11510,N_11307,N_11313);
or U11511 (N_11511,N_11406,N_11163);
and U11512 (N_11512,N_11366,N_11273);
or U11513 (N_11513,N_11402,N_11142);
nor U11514 (N_11514,N_11020,N_11356);
or U11515 (N_11515,N_11037,N_11318);
and U11516 (N_11516,N_11343,N_11216);
or U11517 (N_11517,N_11295,N_11227);
xor U11518 (N_11518,N_11173,N_11261);
nor U11519 (N_11519,N_11033,N_11444);
xor U11520 (N_11520,N_11188,N_11135);
xor U11521 (N_11521,N_11076,N_11004);
nand U11522 (N_11522,N_11215,N_11016);
and U11523 (N_11523,N_11200,N_11109);
or U11524 (N_11524,N_11434,N_11057);
xor U11525 (N_11525,N_11115,N_11330);
xnor U11526 (N_11526,N_11206,N_11498);
and U11527 (N_11527,N_11151,N_11013);
nand U11528 (N_11528,N_11349,N_11238);
nor U11529 (N_11529,N_11376,N_11068);
and U11530 (N_11530,N_11248,N_11241);
nor U11531 (N_11531,N_11214,N_11259);
or U11532 (N_11532,N_11257,N_11422);
nor U11533 (N_11533,N_11412,N_11137);
nand U11534 (N_11534,N_11149,N_11111);
and U11535 (N_11535,N_11050,N_11258);
nand U11536 (N_11536,N_11096,N_11029);
or U11537 (N_11537,N_11445,N_11280);
and U11538 (N_11538,N_11125,N_11457);
nor U11539 (N_11539,N_11092,N_11036);
nand U11540 (N_11540,N_11094,N_11126);
and U11541 (N_11541,N_11011,N_11140);
nor U11542 (N_11542,N_11156,N_11053);
nand U11543 (N_11543,N_11382,N_11452);
or U11544 (N_11544,N_11089,N_11217);
and U11545 (N_11545,N_11022,N_11174);
nor U11546 (N_11546,N_11080,N_11351);
nor U11547 (N_11547,N_11254,N_11473);
or U11548 (N_11548,N_11401,N_11107);
nand U11549 (N_11549,N_11453,N_11097);
nand U11550 (N_11550,N_11272,N_11066);
and U11551 (N_11551,N_11180,N_11463);
xnor U11552 (N_11552,N_11244,N_11339);
nor U11553 (N_11553,N_11440,N_11236);
nor U11554 (N_11554,N_11121,N_11212);
nor U11555 (N_11555,N_11170,N_11314);
nor U11556 (N_11556,N_11370,N_11364);
xor U11557 (N_11557,N_11178,N_11350);
nor U11558 (N_11558,N_11186,N_11347);
nand U11559 (N_11559,N_11276,N_11478);
nor U11560 (N_11560,N_11308,N_11363);
or U11561 (N_11561,N_11185,N_11369);
and U11562 (N_11562,N_11194,N_11493);
xor U11563 (N_11563,N_11411,N_11040);
or U11564 (N_11564,N_11014,N_11102);
nand U11565 (N_11565,N_11472,N_11002);
and U11566 (N_11566,N_11041,N_11116);
or U11567 (N_11567,N_11264,N_11341);
nor U11568 (N_11568,N_11362,N_11449);
nand U11569 (N_11569,N_11322,N_11413);
xor U11570 (N_11570,N_11389,N_11153);
nor U11571 (N_11571,N_11228,N_11270);
and U11572 (N_11572,N_11242,N_11304);
nand U11573 (N_11573,N_11316,N_11381);
and U11574 (N_11574,N_11042,N_11487);
nand U11575 (N_11575,N_11384,N_11371);
nor U11576 (N_11576,N_11101,N_11046);
or U11577 (N_11577,N_11442,N_11133);
or U11578 (N_11578,N_11325,N_11263);
or U11579 (N_11579,N_11265,N_11480);
or U11580 (N_11580,N_11483,N_11485);
xnor U11581 (N_11581,N_11327,N_11438);
nor U11582 (N_11582,N_11315,N_11328);
nand U11583 (N_11583,N_11456,N_11451);
xnor U11584 (N_11584,N_11299,N_11072);
and U11585 (N_11585,N_11117,N_11255);
or U11586 (N_11586,N_11129,N_11179);
or U11587 (N_11587,N_11250,N_11398);
and U11588 (N_11588,N_11394,N_11496);
or U11589 (N_11589,N_11099,N_11465);
or U11590 (N_11590,N_11320,N_11204);
or U11591 (N_11591,N_11021,N_11288);
or U11592 (N_11592,N_11144,N_11035);
nor U11593 (N_11593,N_11197,N_11045);
and U11594 (N_11594,N_11470,N_11058);
nand U11595 (N_11595,N_11158,N_11240);
and U11596 (N_11596,N_11134,N_11428);
nor U11597 (N_11597,N_11348,N_11399);
nor U11598 (N_11598,N_11297,N_11205);
and U11599 (N_11599,N_11132,N_11281);
nand U11600 (N_11600,N_11139,N_11383);
nand U11601 (N_11601,N_11298,N_11077);
nor U11602 (N_11602,N_11291,N_11468);
or U11603 (N_11603,N_11410,N_11252);
nor U11604 (N_11604,N_11495,N_11172);
nor U11605 (N_11605,N_11436,N_11494);
and U11606 (N_11606,N_11462,N_11286);
and U11607 (N_11607,N_11344,N_11497);
or U11608 (N_11608,N_11078,N_11489);
nand U11609 (N_11609,N_11420,N_11333);
or U11610 (N_11610,N_11385,N_11368);
and U11611 (N_11611,N_11332,N_11237);
or U11612 (N_11612,N_11337,N_11051);
nor U11613 (N_11613,N_11340,N_11491);
nor U11614 (N_11614,N_11311,N_11317);
or U11615 (N_11615,N_11195,N_11044);
and U11616 (N_11616,N_11310,N_11375);
or U11617 (N_11617,N_11052,N_11063);
nand U11618 (N_11618,N_11419,N_11028);
or U11619 (N_11619,N_11269,N_11475);
xnor U11620 (N_11620,N_11367,N_11071);
and U11621 (N_11621,N_11305,N_11448);
nor U11622 (N_11622,N_11418,N_11171);
or U11623 (N_11623,N_11079,N_11282);
and U11624 (N_11624,N_11414,N_11147);
and U11625 (N_11625,N_11098,N_11397);
or U11626 (N_11626,N_11431,N_11335);
and U11627 (N_11627,N_11416,N_11441);
nand U11628 (N_11628,N_11395,N_11354);
nand U11629 (N_11629,N_11136,N_11018);
and U11630 (N_11630,N_11155,N_11199);
and U11631 (N_11631,N_11233,N_11458);
nand U11632 (N_11632,N_11081,N_11017);
xor U11633 (N_11633,N_11027,N_11201);
nand U11634 (N_11634,N_11223,N_11471);
xnor U11635 (N_11635,N_11148,N_11119);
or U11636 (N_11636,N_11157,N_11302);
and U11637 (N_11637,N_11226,N_11113);
and U11638 (N_11638,N_11191,N_11001);
or U11639 (N_11639,N_11176,N_11128);
nor U11640 (N_11640,N_11143,N_11105);
nand U11641 (N_11641,N_11127,N_11359);
and U11642 (N_11642,N_11256,N_11060);
nor U11643 (N_11643,N_11222,N_11459);
and U11644 (N_11644,N_11377,N_11166);
and U11645 (N_11645,N_11443,N_11211);
nor U11646 (N_11646,N_11486,N_11426);
or U11647 (N_11647,N_11218,N_11415);
nand U11648 (N_11648,N_11091,N_11246);
or U11649 (N_11649,N_11387,N_11296);
and U11650 (N_11650,N_11067,N_11423);
nor U11651 (N_11651,N_11043,N_11360);
and U11652 (N_11652,N_11235,N_11124);
nor U11653 (N_11653,N_11492,N_11479);
nand U11654 (N_11654,N_11232,N_11239);
nand U11655 (N_11655,N_11221,N_11141);
or U11656 (N_11656,N_11287,N_11294);
or U11657 (N_11657,N_11482,N_11455);
nand U11658 (N_11658,N_11277,N_11353);
or U11659 (N_11659,N_11039,N_11289);
and U11660 (N_11660,N_11225,N_11477);
or U11661 (N_11661,N_11461,N_11408);
and U11662 (N_11662,N_11167,N_11467);
and U11663 (N_11663,N_11184,N_11301);
or U11664 (N_11664,N_11358,N_11106);
nor U11665 (N_11665,N_11292,N_11208);
nor U11666 (N_11666,N_11450,N_11283);
nor U11667 (N_11667,N_11086,N_11293);
or U11668 (N_11668,N_11083,N_11012);
nand U11669 (N_11669,N_11260,N_11231);
or U11670 (N_11670,N_11464,N_11396);
nor U11671 (N_11671,N_11245,N_11271);
nor U11672 (N_11672,N_11405,N_11010);
and U11673 (N_11673,N_11378,N_11407);
nand U11674 (N_11674,N_11251,N_11112);
and U11675 (N_11675,N_11152,N_11075);
nor U11676 (N_11676,N_11323,N_11009);
nand U11677 (N_11677,N_11230,N_11192);
nor U11678 (N_11678,N_11372,N_11490);
xor U11679 (N_11679,N_11164,N_11321);
nand U11680 (N_11680,N_11073,N_11196);
nand U11681 (N_11681,N_11159,N_11131);
nor U11682 (N_11682,N_11070,N_11409);
nand U11683 (N_11683,N_11209,N_11000);
nor U11684 (N_11684,N_11082,N_11160);
xnor U11685 (N_11685,N_11474,N_11345);
or U11686 (N_11686,N_11460,N_11386);
or U11687 (N_11687,N_11229,N_11447);
nor U11688 (N_11688,N_11326,N_11123);
or U11689 (N_11689,N_11120,N_11103);
and U11690 (N_11690,N_11336,N_11061);
nand U11691 (N_11691,N_11114,N_11023);
nor U11692 (N_11692,N_11088,N_11253);
nand U11693 (N_11693,N_11190,N_11433);
nand U11694 (N_11694,N_11476,N_11003);
xnor U11695 (N_11695,N_11267,N_11031);
and U11696 (N_11696,N_11024,N_11404);
nand U11697 (N_11697,N_11285,N_11324);
and U11698 (N_11698,N_11108,N_11048);
or U11699 (N_11699,N_11085,N_11312);
xnor U11700 (N_11700,N_11038,N_11365);
nor U11701 (N_11701,N_11446,N_11005);
nand U11702 (N_11702,N_11187,N_11065);
nor U11703 (N_11703,N_11268,N_11425);
or U11704 (N_11704,N_11224,N_11430);
nand U11705 (N_11705,N_11019,N_11435);
or U11706 (N_11706,N_11403,N_11262);
nor U11707 (N_11707,N_11374,N_11346);
nand U11708 (N_11708,N_11421,N_11373);
nor U11709 (N_11709,N_11355,N_11390);
or U11710 (N_11710,N_11306,N_11026);
nand U11711 (N_11711,N_11122,N_11338);
nand U11712 (N_11712,N_11100,N_11279);
nand U11713 (N_11713,N_11331,N_11484);
or U11714 (N_11714,N_11182,N_11162);
and U11715 (N_11715,N_11145,N_11499);
nand U11716 (N_11716,N_11469,N_11432);
nor U11717 (N_11717,N_11030,N_11303);
or U11718 (N_11718,N_11161,N_11357);
nor U11719 (N_11719,N_11284,N_11243);
and U11720 (N_11720,N_11059,N_11352);
nor U11721 (N_11721,N_11118,N_11247);
nor U11722 (N_11722,N_11424,N_11175);
or U11723 (N_11723,N_11008,N_11213);
nand U11724 (N_11724,N_11025,N_11202);
nor U11725 (N_11725,N_11278,N_11234);
and U11726 (N_11726,N_11056,N_11417);
nand U11727 (N_11727,N_11015,N_11393);
or U11728 (N_11728,N_11049,N_11062);
nand U11729 (N_11729,N_11169,N_11400);
nor U11730 (N_11730,N_11181,N_11220);
nand U11731 (N_11731,N_11064,N_11183);
nand U11732 (N_11732,N_11274,N_11290);
and U11733 (N_11733,N_11138,N_11007);
and U11734 (N_11734,N_11361,N_11150);
and U11735 (N_11735,N_11309,N_11074);
nor U11736 (N_11736,N_11093,N_11069);
and U11737 (N_11737,N_11168,N_11266);
nand U11738 (N_11738,N_11095,N_11466);
and U11739 (N_11739,N_11087,N_11439);
and U11740 (N_11740,N_11275,N_11154);
and U11741 (N_11741,N_11388,N_11391);
nand U11742 (N_11742,N_11090,N_11084);
and U11743 (N_11743,N_11006,N_11130);
and U11744 (N_11744,N_11300,N_11177);
and U11745 (N_11745,N_11110,N_11427);
nor U11746 (N_11746,N_11189,N_11055);
nor U11747 (N_11747,N_11454,N_11392);
nand U11748 (N_11748,N_11032,N_11334);
nor U11749 (N_11749,N_11165,N_11437);
and U11750 (N_11750,N_11385,N_11418);
and U11751 (N_11751,N_11064,N_11014);
nand U11752 (N_11752,N_11163,N_11033);
nor U11753 (N_11753,N_11417,N_11243);
nand U11754 (N_11754,N_11084,N_11028);
nor U11755 (N_11755,N_11265,N_11367);
nand U11756 (N_11756,N_11368,N_11242);
xnor U11757 (N_11757,N_11033,N_11312);
nand U11758 (N_11758,N_11483,N_11106);
and U11759 (N_11759,N_11345,N_11057);
or U11760 (N_11760,N_11454,N_11236);
nand U11761 (N_11761,N_11352,N_11336);
nor U11762 (N_11762,N_11255,N_11397);
and U11763 (N_11763,N_11041,N_11147);
nand U11764 (N_11764,N_11354,N_11494);
and U11765 (N_11765,N_11070,N_11185);
nor U11766 (N_11766,N_11221,N_11218);
nor U11767 (N_11767,N_11163,N_11172);
nor U11768 (N_11768,N_11375,N_11094);
nand U11769 (N_11769,N_11251,N_11093);
and U11770 (N_11770,N_11025,N_11328);
xor U11771 (N_11771,N_11087,N_11479);
or U11772 (N_11772,N_11293,N_11077);
nand U11773 (N_11773,N_11338,N_11205);
or U11774 (N_11774,N_11249,N_11435);
nand U11775 (N_11775,N_11440,N_11446);
or U11776 (N_11776,N_11392,N_11253);
or U11777 (N_11777,N_11072,N_11268);
or U11778 (N_11778,N_11255,N_11455);
nor U11779 (N_11779,N_11163,N_11045);
and U11780 (N_11780,N_11154,N_11091);
or U11781 (N_11781,N_11078,N_11372);
nand U11782 (N_11782,N_11082,N_11449);
xor U11783 (N_11783,N_11194,N_11213);
xor U11784 (N_11784,N_11491,N_11262);
and U11785 (N_11785,N_11156,N_11414);
or U11786 (N_11786,N_11191,N_11030);
or U11787 (N_11787,N_11362,N_11008);
and U11788 (N_11788,N_11121,N_11301);
xor U11789 (N_11789,N_11205,N_11477);
nor U11790 (N_11790,N_11239,N_11112);
or U11791 (N_11791,N_11060,N_11007);
or U11792 (N_11792,N_11164,N_11315);
nand U11793 (N_11793,N_11477,N_11184);
and U11794 (N_11794,N_11468,N_11262);
xor U11795 (N_11795,N_11427,N_11393);
nand U11796 (N_11796,N_11163,N_11345);
nand U11797 (N_11797,N_11043,N_11349);
nor U11798 (N_11798,N_11095,N_11269);
or U11799 (N_11799,N_11219,N_11320);
and U11800 (N_11800,N_11188,N_11042);
and U11801 (N_11801,N_11137,N_11292);
and U11802 (N_11802,N_11014,N_11495);
and U11803 (N_11803,N_11015,N_11146);
xnor U11804 (N_11804,N_11440,N_11148);
xor U11805 (N_11805,N_11257,N_11251);
nand U11806 (N_11806,N_11033,N_11162);
nand U11807 (N_11807,N_11183,N_11469);
and U11808 (N_11808,N_11113,N_11374);
or U11809 (N_11809,N_11043,N_11173);
nor U11810 (N_11810,N_11142,N_11093);
xnor U11811 (N_11811,N_11132,N_11404);
nand U11812 (N_11812,N_11320,N_11207);
and U11813 (N_11813,N_11017,N_11197);
nor U11814 (N_11814,N_11429,N_11145);
or U11815 (N_11815,N_11337,N_11072);
or U11816 (N_11816,N_11332,N_11353);
nand U11817 (N_11817,N_11086,N_11014);
nor U11818 (N_11818,N_11422,N_11121);
xnor U11819 (N_11819,N_11435,N_11467);
or U11820 (N_11820,N_11414,N_11323);
nor U11821 (N_11821,N_11121,N_11178);
or U11822 (N_11822,N_11068,N_11084);
and U11823 (N_11823,N_11250,N_11136);
nand U11824 (N_11824,N_11211,N_11142);
or U11825 (N_11825,N_11447,N_11496);
nor U11826 (N_11826,N_11230,N_11377);
or U11827 (N_11827,N_11161,N_11378);
and U11828 (N_11828,N_11037,N_11255);
xor U11829 (N_11829,N_11427,N_11013);
and U11830 (N_11830,N_11493,N_11480);
or U11831 (N_11831,N_11375,N_11268);
nand U11832 (N_11832,N_11120,N_11264);
xnor U11833 (N_11833,N_11173,N_11101);
xor U11834 (N_11834,N_11267,N_11193);
and U11835 (N_11835,N_11142,N_11377);
and U11836 (N_11836,N_11172,N_11186);
nor U11837 (N_11837,N_11297,N_11017);
or U11838 (N_11838,N_11022,N_11309);
nand U11839 (N_11839,N_11345,N_11048);
nand U11840 (N_11840,N_11028,N_11117);
and U11841 (N_11841,N_11203,N_11489);
and U11842 (N_11842,N_11006,N_11392);
nand U11843 (N_11843,N_11169,N_11323);
nor U11844 (N_11844,N_11076,N_11115);
or U11845 (N_11845,N_11274,N_11027);
nand U11846 (N_11846,N_11497,N_11451);
or U11847 (N_11847,N_11407,N_11260);
and U11848 (N_11848,N_11443,N_11164);
nand U11849 (N_11849,N_11273,N_11471);
xnor U11850 (N_11850,N_11375,N_11355);
nor U11851 (N_11851,N_11131,N_11330);
nor U11852 (N_11852,N_11126,N_11135);
and U11853 (N_11853,N_11258,N_11172);
nor U11854 (N_11854,N_11012,N_11372);
or U11855 (N_11855,N_11423,N_11321);
xor U11856 (N_11856,N_11333,N_11242);
or U11857 (N_11857,N_11417,N_11430);
nand U11858 (N_11858,N_11451,N_11185);
and U11859 (N_11859,N_11429,N_11160);
nand U11860 (N_11860,N_11126,N_11427);
xnor U11861 (N_11861,N_11372,N_11050);
and U11862 (N_11862,N_11057,N_11062);
and U11863 (N_11863,N_11170,N_11078);
or U11864 (N_11864,N_11167,N_11440);
or U11865 (N_11865,N_11458,N_11351);
and U11866 (N_11866,N_11022,N_11423);
nor U11867 (N_11867,N_11019,N_11346);
and U11868 (N_11868,N_11409,N_11435);
and U11869 (N_11869,N_11011,N_11190);
nand U11870 (N_11870,N_11246,N_11252);
or U11871 (N_11871,N_11328,N_11261);
and U11872 (N_11872,N_11060,N_11267);
or U11873 (N_11873,N_11146,N_11123);
xnor U11874 (N_11874,N_11415,N_11290);
xor U11875 (N_11875,N_11134,N_11446);
nor U11876 (N_11876,N_11327,N_11487);
nor U11877 (N_11877,N_11155,N_11324);
nand U11878 (N_11878,N_11449,N_11261);
nor U11879 (N_11879,N_11183,N_11169);
or U11880 (N_11880,N_11095,N_11182);
and U11881 (N_11881,N_11340,N_11277);
nand U11882 (N_11882,N_11459,N_11178);
and U11883 (N_11883,N_11183,N_11108);
nor U11884 (N_11884,N_11202,N_11252);
nand U11885 (N_11885,N_11191,N_11434);
nand U11886 (N_11886,N_11061,N_11202);
nand U11887 (N_11887,N_11155,N_11183);
nor U11888 (N_11888,N_11218,N_11056);
and U11889 (N_11889,N_11055,N_11363);
nand U11890 (N_11890,N_11493,N_11261);
and U11891 (N_11891,N_11195,N_11372);
nand U11892 (N_11892,N_11423,N_11083);
nand U11893 (N_11893,N_11116,N_11259);
nand U11894 (N_11894,N_11255,N_11267);
nor U11895 (N_11895,N_11128,N_11079);
and U11896 (N_11896,N_11274,N_11329);
nor U11897 (N_11897,N_11044,N_11043);
nor U11898 (N_11898,N_11246,N_11016);
or U11899 (N_11899,N_11368,N_11006);
nand U11900 (N_11900,N_11321,N_11298);
nor U11901 (N_11901,N_11270,N_11280);
or U11902 (N_11902,N_11378,N_11408);
and U11903 (N_11903,N_11406,N_11295);
nand U11904 (N_11904,N_11340,N_11090);
nand U11905 (N_11905,N_11427,N_11296);
and U11906 (N_11906,N_11027,N_11364);
or U11907 (N_11907,N_11144,N_11097);
nand U11908 (N_11908,N_11234,N_11126);
nor U11909 (N_11909,N_11110,N_11066);
nand U11910 (N_11910,N_11373,N_11417);
or U11911 (N_11911,N_11437,N_11269);
and U11912 (N_11912,N_11426,N_11411);
and U11913 (N_11913,N_11180,N_11197);
and U11914 (N_11914,N_11474,N_11105);
and U11915 (N_11915,N_11445,N_11295);
and U11916 (N_11916,N_11430,N_11404);
or U11917 (N_11917,N_11418,N_11179);
and U11918 (N_11918,N_11116,N_11039);
xnor U11919 (N_11919,N_11058,N_11122);
nand U11920 (N_11920,N_11291,N_11344);
nor U11921 (N_11921,N_11260,N_11492);
and U11922 (N_11922,N_11475,N_11136);
or U11923 (N_11923,N_11345,N_11338);
or U11924 (N_11924,N_11268,N_11423);
xnor U11925 (N_11925,N_11428,N_11171);
or U11926 (N_11926,N_11245,N_11440);
nor U11927 (N_11927,N_11400,N_11403);
and U11928 (N_11928,N_11260,N_11130);
or U11929 (N_11929,N_11083,N_11264);
nand U11930 (N_11930,N_11429,N_11187);
nand U11931 (N_11931,N_11210,N_11075);
or U11932 (N_11932,N_11479,N_11324);
nand U11933 (N_11933,N_11173,N_11019);
xor U11934 (N_11934,N_11399,N_11494);
nand U11935 (N_11935,N_11497,N_11117);
or U11936 (N_11936,N_11230,N_11145);
or U11937 (N_11937,N_11422,N_11499);
nor U11938 (N_11938,N_11291,N_11494);
nand U11939 (N_11939,N_11008,N_11066);
and U11940 (N_11940,N_11375,N_11198);
or U11941 (N_11941,N_11400,N_11343);
or U11942 (N_11942,N_11214,N_11092);
and U11943 (N_11943,N_11306,N_11015);
nor U11944 (N_11944,N_11423,N_11184);
or U11945 (N_11945,N_11031,N_11081);
or U11946 (N_11946,N_11020,N_11413);
and U11947 (N_11947,N_11254,N_11138);
or U11948 (N_11948,N_11104,N_11253);
xor U11949 (N_11949,N_11449,N_11216);
nand U11950 (N_11950,N_11126,N_11262);
nor U11951 (N_11951,N_11367,N_11207);
nor U11952 (N_11952,N_11112,N_11363);
xor U11953 (N_11953,N_11287,N_11074);
nor U11954 (N_11954,N_11299,N_11311);
nor U11955 (N_11955,N_11096,N_11268);
nand U11956 (N_11956,N_11343,N_11431);
or U11957 (N_11957,N_11365,N_11237);
xnor U11958 (N_11958,N_11297,N_11453);
nand U11959 (N_11959,N_11199,N_11462);
xor U11960 (N_11960,N_11032,N_11055);
or U11961 (N_11961,N_11245,N_11205);
and U11962 (N_11962,N_11269,N_11406);
xor U11963 (N_11963,N_11316,N_11277);
and U11964 (N_11964,N_11364,N_11353);
and U11965 (N_11965,N_11445,N_11019);
nand U11966 (N_11966,N_11457,N_11088);
or U11967 (N_11967,N_11120,N_11316);
nand U11968 (N_11968,N_11150,N_11024);
nand U11969 (N_11969,N_11060,N_11454);
or U11970 (N_11970,N_11039,N_11272);
nand U11971 (N_11971,N_11227,N_11427);
or U11972 (N_11972,N_11062,N_11343);
nor U11973 (N_11973,N_11441,N_11031);
nand U11974 (N_11974,N_11480,N_11473);
nor U11975 (N_11975,N_11397,N_11341);
xor U11976 (N_11976,N_11111,N_11306);
nor U11977 (N_11977,N_11471,N_11332);
and U11978 (N_11978,N_11044,N_11295);
and U11979 (N_11979,N_11298,N_11103);
nor U11980 (N_11980,N_11461,N_11041);
and U11981 (N_11981,N_11197,N_11081);
or U11982 (N_11982,N_11042,N_11044);
nor U11983 (N_11983,N_11493,N_11272);
or U11984 (N_11984,N_11353,N_11211);
or U11985 (N_11985,N_11230,N_11321);
or U11986 (N_11986,N_11302,N_11090);
and U11987 (N_11987,N_11464,N_11364);
nor U11988 (N_11988,N_11463,N_11426);
nor U11989 (N_11989,N_11496,N_11018);
nand U11990 (N_11990,N_11453,N_11325);
or U11991 (N_11991,N_11044,N_11422);
or U11992 (N_11992,N_11226,N_11109);
and U11993 (N_11993,N_11413,N_11179);
or U11994 (N_11994,N_11361,N_11435);
nand U11995 (N_11995,N_11271,N_11394);
nand U11996 (N_11996,N_11377,N_11318);
nor U11997 (N_11997,N_11487,N_11074);
or U11998 (N_11998,N_11285,N_11160);
nand U11999 (N_11999,N_11492,N_11295);
nand U12000 (N_12000,N_11801,N_11539);
or U12001 (N_12001,N_11748,N_11635);
nor U12002 (N_12002,N_11812,N_11746);
or U12003 (N_12003,N_11650,N_11515);
and U12004 (N_12004,N_11928,N_11626);
or U12005 (N_12005,N_11716,N_11825);
nor U12006 (N_12006,N_11987,N_11548);
and U12007 (N_12007,N_11949,N_11624);
nand U12008 (N_12008,N_11594,N_11938);
and U12009 (N_12009,N_11772,N_11702);
nand U12010 (N_12010,N_11981,N_11512);
nor U12011 (N_12011,N_11931,N_11851);
nor U12012 (N_12012,N_11781,N_11526);
and U12013 (N_12013,N_11875,N_11671);
nand U12014 (N_12014,N_11845,N_11970);
and U12015 (N_12015,N_11842,N_11856);
nor U12016 (N_12016,N_11819,N_11621);
or U12017 (N_12017,N_11735,N_11955);
or U12018 (N_12018,N_11606,N_11742);
or U12019 (N_12019,N_11571,N_11761);
nor U12020 (N_12020,N_11925,N_11718);
or U12021 (N_12021,N_11881,N_11706);
nand U12022 (N_12022,N_11904,N_11976);
nor U12023 (N_12023,N_11800,N_11648);
nand U12024 (N_12024,N_11561,N_11877);
or U12025 (N_12025,N_11942,N_11973);
nand U12026 (N_12026,N_11791,N_11803);
nor U12027 (N_12027,N_11897,N_11866);
and U12028 (N_12028,N_11972,N_11874);
nor U12029 (N_12029,N_11661,N_11672);
nor U12030 (N_12030,N_11757,N_11598);
nor U12031 (N_12031,N_11787,N_11550);
and U12032 (N_12032,N_11788,N_11708);
nor U12033 (N_12033,N_11604,N_11783);
and U12034 (N_12034,N_11560,N_11950);
or U12035 (N_12035,N_11755,N_11717);
nand U12036 (N_12036,N_11597,N_11815);
nand U12037 (N_12037,N_11760,N_11599);
nor U12038 (N_12038,N_11872,N_11634);
or U12039 (N_12039,N_11617,N_11922);
nand U12040 (N_12040,N_11618,N_11502);
or U12041 (N_12041,N_11688,N_11847);
and U12042 (N_12042,N_11699,N_11587);
nand U12043 (N_12043,N_11971,N_11577);
xnor U12044 (N_12044,N_11697,N_11632);
nand U12045 (N_12045,N_11883,N_11643);
and U12046 (N_12046,N_11703,N_11542);
and U12047 (N_12047,N_11558,N_11764);
nand U12048 (N_12048,N_11848,N_11712);
nor U12049 (N_12049,N_11951,N_11727);
xnor U12050 (N_12050,N_11930,N_11743);
nor U12051 (N_12051,N_11568,N_11553);
nand U12052 (N_12052,N_11696,N_11513);
or U12053 (N_12053,N_11879,N_11850);
nor U12054 (N_12054,N_11592,N_11892);
nand U12055 (N_12055,N_11580,N_11582);
or U12056 (N_12056,N_11555,N_11779);
nor U12057 (N_12057,N_11777,N_11609);
nand U12058 (N_12058,N_11878,N_11759);
nand U12059 (N_12059,N_11989,N_11816);
nand U12060 (N_12060,N_11682,N_11530);
or U12061 (N_12061,N_11694,N_11662);
and U12062 (N_12062,N_11993,N_11956);
xor U12063 (N_12063,N_11821,N_11957);
and U12064 (N_12064,N_11893,N_11572);
and U12065 (N_12065,N_11503,N_11614);
or U12066 (N_12066,N_11836,N_11969);
nor U12067 (N_12067,N_11645,N_11522);
or U12068 (N_12068,N_11932,N_11722);
nand U12069 (N_12069,N_11982,N_11730);
nand U12070 (N_12070,N_11911,N_11670);
nand U12071 (N_12071,N_11880,N_11983);
and U12072 (N_12072,N_11998,N_11758);
nor U12073 (N_12073,N_11538,N_11543);
and U12074 (N_12074,N_11826,N_11595);
nor U12075 (N_12075,N_11858,N_11683);
and U12076 (N_12076,N_11705,N_11979);
xnor U12077 (N_12077,N_11666,N_11610);
nand U12078 (N_12078,N_11792,N_11546);
and U12079 (N_12079,N_11860,N_11615);
nor U12080 (N_12080,N_11778,N_11590);
nand U12081 (N_12081,N_11707,N_11579);
nor U12082 (N_12082,N_11769,N_11766);
xor U12083 (N_12083,N_11934,N_11745);
and U12084 (N_12084,N_11501,N_11919);
xnor U12085 (N_12085,N_11637,N_11832);
nor U12086 (N_12086,N_11959,N_11625);
or U12087 (N_12087,N_11574,N_11713);
nor U12088 (N_12088,N_11865,N_11827);
or U12089 (N_12089,N_11569,N_11960);
nor U12090 (N_12090,N_11948,N_11744);
or U12091 (N_12091,N_11738,N_11863);
and U12092 (N_12092,N_11655,N_11693);
nor U12093 (N_12093,N_11822,N_11844);
xnor U12094 (N_12094,N_11888,N_11737);
or U12095 (N_12095,N_11506,N_11941);
and U12096 (N_12096,N_11521,N_11747);
or U12097 (N_12097,N_11963,N_11966);
nand U12098 (N_12098,N_11838,N_11641);
or U12099 (N_12099,N_11564,N_11926);
nand U12100 (N_12100,N_11669,N_11802);
xnor U12101 (N_12101,N_11940,N_11869);
and U12102 (N_12102,N_11554,N_11518);
nor U12103 (N_12103,N_11837,N_11808);
and U12104 (N_12104,N_11817,N_11921);
nand U12105 (N_12105,N_11629,N_11517);
nor U12106 (N_12106,N_11768,N_11652);
and U12107 (N_12107,N_11642,N_11656);
and U12108 (N_12108,N_11562,N_11780);
or U12109 (N_12109,N_11684,N_11531);
or U12110 (N_12110,N_11774,N_11534);
xnor U12111 (N_12111,N_11859,N_11849);
nor U12112 (N_12112,N_11529,N_11762);
nand U12113 (N_12113,N_11952,N_11771);
nor U12114 (N_12114,N_11603,N_11570);
nor U12115 (N_12115,N_11915,N_11732);
and U12116 (N_12116,N_11585,N_11828);
nor U12117 (N_12117,N_11830,N_11551);
and U12118 (N_12118,N_11638,N_11514);
nand U12119 (N_12119,N_11796,N_11834);
or U12120 (N_12120,N_11937,N_11923);
nand U12121 (N_12121,N_11965,N_11944);
nor U12122 (N_12122,N_11523,N_11612);
nand U12123 (N_12123,N_11654,N_11516);
and U12124 (N_12124,N_11677,N_11527);
or U12125 (N_12125,N_11867,N_11907);
and U12126 (N_12126,N_11770,N_11994);
and U12127 (N_12127,N_11789,N_11695);
nor U12128 (N_12128,N_11639,N_11912);
nor U12129 (N_12129,N_11573,N_11927);
xor U12130 (N_12130,N_11507,N_11895);
and U12131 (N_12131,N_11547,N_11709);
nand U12132 (N_12132,N_11906,N_11914);
nor U12133 (N_12133,N_11933,N_11601);
nor U12134 (N_12134,N_11619,N_11685);
or U12135 (N_12135,N_11908,N_11823);
nand U12136 (N_12136,N_11630,N_11646);
nand U12137 (N_12137,N_11776,N_11556);
xor U12138 (N_12138,N_11790,N_11903);
and U12139 (N_12139,N_11721,N_11528);
nand U12140 (N_12140,N_11861,N_11846);
nor U12141 (N_12141,N_11833,N_11751);
and U12142 (N_12142,N_11588,N_11997);
and U12143 (N_12143,N_11750,N_11767);
nor U12144 (N_12144,N_11633,N_11687);
nor U12145 (N_12145,N_11765,N_11678);
xor U12146 (N_12146,N_11884,N_11991);
nand U12147 (N_12147,N_11961,N_11784);
and U12148 (N_12148,N_11567,N_11565);
or U12149 (N_12149,N_11964,N_11977);
and U12150 (N_12150,N_11936,N_11798);
and U12151 (N_12151,N_11692,N_11584);
xor U12152 (N_12152,N_11811,N_11797);
nor U12153 (N_12153,N_11887,N_11525);
or U12154 (N_12154,N_11710,N_11726);
and U12155 (N_12155,N_11524,N_11975);
or U12156 (N_12156,N_11575,N_11731);
nor U12157 (N_12157,N_11831,N_11739);
nor U12158 (N_12158,N_11651,N_11756);
nand U12159 (N_12159,N_11886,N_11613);
nor U12160 (N_12160,N_11946,N_11552);
nor U12161 (N_12161,N_11520,N_11804);
nand U12162 (N_12162,N_11676,N_11871);
nor U12163 (N_12163,N_11999,N_11704);
or U12164 (N_12164,N_11985,N_11749);
nand U12165 (N_12165,N_11537,N_11807);
nor U12166 (N_12166,N_11852,N_11891);
nand U12167 (N_12167,N_11700,N_11868);
or U12168 (N_12168,N_11535,N_11578);
nand U12169 (N_12169,N_11794,N_11902);
and U12170 (N_12170,N_11775,N_11929);
xor U12171 (N_12171,N_11910,N_11740);
and U12172 (N_12172,N_11644,N_11862);
nor U12173 (N_12173,N_11978,N_11668);
xnor U12174 (N_12174,N_11943,N_11992);
nand U12175 (N_12175,N_11754,N_11689);
nor U12176 (N_12176,N_11636,N_11876);
and U12177 (N_12177,N_11995,N_11586);
nor U12178 (N_12178,N_11917,N_11674);
or U12179 (N_12179,N_11741,N_11665);
and U12180 (N_12180,N_11729,N_11611);
and U12181 (N_12181,N_11894,N_11589);
nor U12182 (N_12182,N_11968,N_11782);
xor U12183 (N_12183,N_11889,N_11924);
nor U12184 (N_12184,N_11773,N_11544);
and U12185 (N_12185,N_11882,N_11505);
nand U12186 (N_12186,N_11840,N_11663);
xor U12187 (N_12187,N_11628,N_11627);
and U12188 (N_12188,N_11820,N_11898);
nand U12189 (N_12189,N_11935,N_11864);
or U12190 (N_12190,N_11583,N_11631);
and U12191 (N_12191,N_11647,N_11785);
nand U12192 (N_12192,N_11786,N_11733);
xnor U12193 (N_12193,N_11974,N_11591);
nand U12194 (N_12194,N_11873,N_11673);
or U12195 (N_12195,N_11988,N_11596);
nand U12196 (N_12196,N_11679,N_11667);
nor U12197 (N_12197,N_11753,N_11723);
nor U12198 (N_12198,N_11870,N_11607);
xnor U12199 (N_12199,N_11841,N_11714);
and U12200 (N_12200,N_11620,N_11608);
and U12201 (N_12201,N_11900,N_11605);
nand U12202 (N_12202,N_11909,N_11519);
nor U12203 (N_12203,N_11899,N_11799);
or U12204 (N_12204,N_11725,N_11504);
xnor U12205 (N_12205,N_11509,N_11962);
and U12206 (N_12206,N_11814,N_11824);
and U12207 (N_12207,N_11920,N_11533);
nand U12208 (N_12208,N_11813,N_11839);
nand U12209 (N_12209,N_11795,N_11675);
and U12210 (N_12210,N_11691,N_11954);
and U12211 (N_12211,N_11649,N_11719);
nor U12212 (N_12212,N_11953,N_11510);
and U12213 (N_12213,N_11809,N_11855);
and U12214 (N_12214,N_11576,N_11511);
nand U12215 (N_12215,N_11947,N_11916);
xor U12216 (N_12216,N_11600,N_11980);
xor U12217 (N_12217,N_11660,N_11835);
nor U12218 (N_12218,N_11958,N_11653);
nor U12219 (N_12219,N_11829,N_11805);
or U12220 (N_12220,N_11686,N_11945);
or U12221 (N_12221,N_11853,N_11657);
and U12222 (N_12222,N_11622,N_11640);
xnor U12223 (N_12223,N_11752,N_11681);
nor U12224 (N_12224,N_11967,N_11793);
nor U12225 (N_12225,N_11905,N_11885);
nor U12226 (N_12226,N_11508,N_11616);
or U12227 (N_12227,N_11698,N_11680);
or U12228 (N_12228,N_11996,N_11806);
or U12229 (N_12229,N_11500,N_11901);
nor U12230 (N_12230,N_11724,N_11581);
nand U12231 (N_12231,N_11734,N_11810);
nor U12232 (N_12232,N_11623,N_11659);
and U12233 (N_12233,N_11913,N_11711);
and U12234 (N_12234,N_11896,N_11715);
xnor U12235 (N_12235,N_11939,N_11549);
or U12236 (N_12236,N_11541,N_11536);
nor U12237 (N_12237,N_11545,N_11857);
nand U12238 (N_12238,N_11559,N_11984);
or U12239 (N_12239,N_11664,N_11854);
or U12240 (N_12240,N_11728,N_11990);
nor U12241 (N_12241,N_11701,N_11890);
nand U12242 (N_12242,N_11557,N_11918);
nand U12243 (N_12243,N_11593,N_11763);
or U12244 (N_12244,N_11720,N_11986);
and U12245 (N_12245,N_11566,N_11818);
and U12246 (N_12246,N_11532,N_11602);
and U12247 (N_12247,N_11658,N_11690);
nor U12248 (N_12248,N_11736,N_11563);
nor U12249 (N_12249,N_11843,N_11540);
xor U12250 (N_12250,N_11904,N_11706);
nor U12251 (N_12251,N_11567,N_11543);
nor U12252 (N_12252,N_11647,N_11993);
or U12253 (N_12253,N_11763,N_11935);
nand U12254 (N_12254,N_11919,N_11954);
or U12255 (N_12255,N_11832,N_11908);
xnor U12256 (N_12256,N_11600,N_11937);
and U12257 (N_12257,N_11847,N_11987);
nand U12258 (N_12258,N_11590,N_11566);
xnor U12259 (N_12259,N_11529,N_11897);
or U12260 (N_12260,N_11543,N_11750);
nand U12261 (N_12261,N_11501,N_11888);
or U12262 (N_12262,N_11870,N_11950);
xor U12263 (N_12263,N_11811,N_11933);
or U12264 (N_12264,N_11695,N_11694);
and U12265 (N_12265,N_11961,N_11627);
nor U12266 (N_12266,N_11774,N_11675);
nor U12267 (N_12267,N_11638,N_11743);
or U12268 (N_12268,N_11753,N_11651);
and U12269 (N_12269,N_11768,N_11963);
nor U12270 (N_12270,N_11501,N_11939);
xnor U12271 (N_12271,N_11542,N_11627);
and U12272 (N_12272,N_11701,N_11911);
nor U12273 (N_12273,N_11993,N_11502);
nand U12274 (N_12274,N_11868,N_11577);
and U12275 (N_12275,N_11792,N_11704);
nand U12276 (N_12276,N_11994,N_11623);
xor U12277 (N_12277,N_11518,N_11664);
or U12278 (N_12278,N_11729,N_11817);
nand U12279 (N_12279,N_11756,N_11712);
nand U12280 (N_12280,N_11773,N_11823);
nor U12281 (N_12281,N_11955,N_11557);
nand U12282 (N_12282,N_11968,N_11519);
and U12283 (N_12283,N_11813,N_11938);
or U12284 (N_12284,N_11903,N_11942);
nand U12285 (N_12285,N_11578,N_11645);
and U12286 (N_12286,N_11732,N_11629);
nand U12287 (N_12287,N_11598,N_11719);
nand U12288 (N_12288,N_11615,N_11918);
nor U12289 (N_12289,N_11653,N_11707);
and U12290 (N_12290,N_11772,N_11840);
nand U12291 (N_12291,N_11625,N_11567);
and U12292 (N_12292,N_11505,N_11694);
xor U12293 (N_12293,N_11721,N_11846);
or U12294 (N_12294,N_11640,N_11923);
nand U12295 (N_12295,N_11739,N_11772);
nor U12296 (N_12296,N_11954,N_11735);
nor U12297 (N_12297,N_11735,N_11558);
nor U12298 (N_12298,N_11620,N_11827);
nor U12299 (N_12299,N_11588,N_11771);
nor U12300 (N_12300,N_11864,N_11887);
xnor U12301 (N_12301,N_11693,N_11672);
nor U12302 (N_12302,N_11565,N_11994);
nand U12303 (N_12303,N_11788,N_11611);
nand U12304 (N_12304,N_11554,N_11920);
nor U12305 (N_12305,N_11842,N_11627);
nand U12306 (N_12306,N_11950,N_11925);
or U12307 (N_12307,N_11567,N_11564);
nor U12308 (N_12308,N_11794,N_11586);
or U12309 (N_12309,N_11539,N_11664);
nor U12310 (N_12310,N_11928,N_11876);
or U12311 (N_12311,N_11736,N_11511);
nand U12312 (N_12312,N_11570,N_11572);
nor U12313 (N_12313,N_11506,N_11671);
nor U12314 (N_12314,N_11740,N_11742);
or U12315 (N_12315,N_11627,N_11737);
nor U12316 (N_12316,N_11862,N_11981);
and U12317 (N_12317,N_11820,N_11805);
nor U12318 (N_12318,N_11532,N_11827);
or U12319 (N_12319,N_11868,N_11982);
nor U12320 (N_12320,N_11685,N_11518);
and U12321 (N_12321,N_11753,N_11628);
nand U12322 (N_12322,N_11661,N_11711);
nand U12323 (N_12323,N_11569,N_11873);
nor U12324 (N_12324,N_11912,N_11649);
or U12325 (N_12325,N_11922,N_11602);
nand U12326 (N_12326,N_11724,N_11926);
nor U12327 (N_12327,N_11855,N_11796);
xor U12328 (N_12328,N_11937,N_11793);
nor U12329 (N_12329,N_11850,N_11632);
xnor U12330 (N_12330,N_11986,N_11575);
and U12331 (N_12331,N_11609,N_11621);
or U12332 (N_12332,N_11543,N_11885);
and U12333 (N_12333,N_11533,N_11856);
nor U12334 (N_12334,N_11761,N_11972);
and U12335 (N_12335,N_11667,N_11767);
nor U12336 (N_12336,N_11675,N_11645);
nand U12337 (N_12337,N_11758,N_11927);
or U12338 (N_12338,N_11599,N_11679);
and U12339 (N_12339,N_11892,N_11840);
nor U12340 (N_12340,N_11919,N_11517);
or U12341 (N_12341,N_11515,N_11588);
nand U12342 (N_12342,N_11762,N_11826);
and U12343 (N_12343,N_11673,N_11781);
nor U12344 (N_12344,N_11964,N_11854);
or U12345 (N_12345,N_11661,N_11983);
and U12346 (N_12346,N_11693,N_11871);
nand U12347 (N_12347,N_11676,N_11940);
nand U12348 (N_12348,N_11582,N_11760);
and U12349 (N_12349,N_11811,N_11982);
or U12350 (N_12350,N_11509,N_11516);
nand U12351 (N_12351,N_11848,N_11730);
or U12352 (N_12352,N_11619,N_11826);
xnor U12353 (N_12353,N_11890,N_11719);
nand U12354 (N_12354,N_11524,N_11712);
nand U12355 (N_12355,N_11507,N_11629);
nor U12356 (N_12356,N_11508,N_11935);
nand U12357 (N_12357,N_11586,N_11549);
or U12358 (N_12358,N_11816,N_11583);
and U12359 (N_12359,N_11638,N_11574);
nand U12360 (N_12360,N_11800,N_11986);
xor U12361 (N_12361,N_11594,N_11643);
xor U12362 (N_12362,N_11999,N_11762);
or U12363 (N_12363,N_11624,N_11577);
nand U12364 (N_12364,N_11632,N_11883);
or U12365 (N_12365,N_11892,N_11701);
and U12366 (N_12366,N_11618,N_11640);
nor U12367 (N_12367,N_11766,N_11558);
and U12368 (N_12368,N_11608,N_11634);
nor U12369 (N_12369,N_11802,N_11595);
or U12370 (N_12370,N_11892,N_11918);
and U12371 (N_12371,N_11927,N_11982);
xor U12372 (N_12372,N_11813,N_11739);
or U12373 (N_12373,N_11838,N_11551);
xnor U12374 (N_12374,N_11608,N_11700);
or U12375 (N_12375,N_11504,N_11663);
nand U12376 (N_12376,N_11516,N_11943);
or U12377 (N_12377,N_11579,N_11528);
or U12378 (N_12378,N_11606,N_11540);
or U12379 (N_12379,N_11879,N_11618);
nand U12380 (N_12380,N_11822,N_11571);
nor U12381 (N_12381,N_11571,N_11725);
nor U12382 (N_12382,N_11886,N_11888);
xor U12383 (N_12383,N_11583,N_11992);
and U12384 (N_12384,N_11520,N_11534);
and U12385 (N_12385,N_11630,N_11906);
nor U12386 (N_12386,N_11917,N_11801);
or U12387 (N_12387,N_11594,N_11931);
nand U12388 (N_12388,N_11869,N_11791);
or U12389 (N_12389,N_11994,N_11653);
nor U12390 (N_12390,N_11552,N_11846);
and U12391 (N_12391,N_11532,N_11865);
xor U12392 (N_12392,N_11947,N_11580);
or U12393 (N_12393,N_11568,N_11981);
nand U12394 (N_12394,N_11641,N_11914);
or U12395 (N_12395,N_11900,N_11549);
nand U12396 (N_12396,N_11529,N_11714);
xnor U12397 (N_12397,N_11662,N_11962);
and U12398 (N_12398,N_11964,N_11776);
nor U12399 (N_12399,N_11607,N_11861);
or U12400 (N_12400,N_11639,N_11894);
nand U12401 (N_12401,N_11590,N_11521);
nor U12402 (N_12402,N_11708,N_11731);
nand U12403 (N_12403,N_11847,N_11906);
nor U12404 (N_12404,N_11561,N_11719);
and U12405 (N_12405,N_11692,N_11813);
nand U12406 (N_12406,N_11558,N_11902);
or U12407 (N_12407,N_11800,N_11786);
nor U12408 (N_12408,N_11807,N_11938);
xor U12409 (N_12409,N_11950,N_11568);
and U12410 (N_12410,N_11843,N_11550);
or U12411 (N_12411,N_11885,N_11948);
nand U12412 (N_12412,N_11645,N_11889);
nor U12413 (N_12413,N_11728,N_11942);
or U12414 (N_12414,N_11610,N_11557);
and U12415 (N_12415,N_11657,N_11573);
or U12416 (N_12416,N_11651,N_11608);
and U12417 (N_12417,N_11628,N_11882);
nand U12418 (N_12418,N_11922,N_11523);
and U12419 (N_12419,N_11751,N_11978);
nor U12420 (N_12420,N_11940,N_11737);
nor U12421 (N_12421,N_11702,N_11959);
or U12422 (N_12422,N_11585,N_11974);
and U12423 (N_12423,N_11953,N_11848);
and U12424 (N_12424,N_11794,N_11630);
or U12425 (N_12425,N_11769,N_11741);
nor U12426 (N_12426,N_11858,N_11944);
xor U12427 (N_12427,N_11599,N_11856);
and U12428 (N_12428,N_11936,N_11857);
and U12429 (N_12429,N_11919,N_11816);
or U12430 (N_12430,N_11957,N_11741);
nand U12431 (N_12431,N_11840,N_11745);
xnor U12432 (N_12432,N_11538,N_11869);
xor U12433 (N_12433,N_11635,N_11686);
and U12434 (N_12434,N_11608,N_11998);
nor U12435 (N_12435,N_11739,N_11908);
or U12436 (N_12436,N_11687,N_11626);
nand U12437 (N_12437,N_11918,N_11905);
nand U12438 (N_12438,N_11751,N_11524);
nand U12439 (N_12439,N_11515,N_11782);
nand U12440 (N_12440,N_11645,N_11545);
nor U12441 (N_12441,N_11932,N_11715);
nor U12442 (N_12442,N_11503,N_11885);
nor U12443 (N_12443,N_11637,N_11799);
or U12444 (N_12444,N_11748,N_11978);
or U12445 (N_12445,N_11847,N_11522);
and U12446 (N_12446,N_11512,N_11696);
or U12447 (N_12447,N_11589,N_11509);
nor U12448 (N_12448,N_11544,N_11813);
and U12449 (N_12449,N_11908,N_11963);
nand U12450 (N_12450,N_11650,N_11988);
or U12451 (N_12451,N_11626,N_11922);
or U12452 (N_12452,N_11733,N_11875);
and U12453 (N_12453,N_11749,N_11557);
and U12454 (N_12454,N_11565,N_11837);
nor U12455 (N_12455,N_11611,N_11523);
or U12456 (N_12456,N_11751,N_11609);
nand U12457 (N_12457,N_11701,N_11638);
nor U12458 (N_12458,N_11759,N_11962);
nor U12459 (N_12459,N_11990,N_11863);
and U12460 (N_12460,N_11860,N_11807);
and U12461 (N_12461,N_11635,N_11681);
or U12462 (N_12462,N_11921,N_11927);
nand U12463 (N_12463,N_11909,N_11505);
or U12464 (N_12464,N_11661,N_11582);
or U12465 (N_12465,N_11967,N_11930);
or U12466 (N_12466,N_11731,N_11646);
or U12467 (N_12467,N_11718,N_11597);
or U12468 (N_12468,N_11629,N_11818);
and U12469 (N_12469,N_11998,N_11738);
nor U12470 (N_12470,N_11948,N_11596);
xnor U12471 (N_12471,N_11825,N_11719);
or U12472 (N_12472,N_11538,N_11979);
nor U12473 (N_12473,N_11773,N_11732);
or U12474 (N_12474,N_11958,N_11889);
or U12475 (N_12475,N_11766,N_11752);
nor U12476 (N_12476,N_11510,N_11545);
or U12477 (N_12477,N_11855,N_11833);
nor U12478 (N_12478,N_11711,N_11954);
or U12479 (N_12479,N_11707,N_11956);
nand U12480 (N_12480,N_11615,N_11673);
nor U12481 (N_12481,N_11978,N_11781);
nor U12482 (N_12482,N_11544,N_11617);
nor U12483 (N_12483,N_11792,N_11857);
nor U12484 (N_12484,N_11791,N_11853);
nand U12485 (N_12485,N_11693,N_11934);
or U12486 (N_12486,N_11648,N_11962);
and U12487 (N_12487,N_11600,N_11855);
nand U12488 (N_12488,N_11666,N_11755);
and U12489 (N_12489,N_11516,N_11658);
xnor U12490 (N_12490,N_11633,N_11744);
nor U12491 (N_12491,N_11787,N_11817);
and U12492 (N_12492,N_11647,N_11772);
nor U12493 (N_12493,N_11568,N_11953);
xnor U12494 (N_12494,N_11935,N_11601);
nand U12495 (N_12495,N_11984,N_11721);
or U12496 (N_12496,N_11517,N_11653);
and U12497 (N_12497,N_11502,N_11680);
nand U12498 (N_12498,N_11903,N_11999);
nand U12499 (N_12499,N_11705,N_11891);
and U12500 (N_12500,N_12148,N_12192);
nor U12501 (N_12501,N_12352,N_12254);
nand U12502 (N_12502,N_12472,N_12016);
nor U12503 (N_12503,N_12340,N_12443);
and U12504 (N_12504,N_12456,N_12180);
xnor U12505 (N_12505,N_12412,N_12074);
nor U12506 (N_12506,N_12140,N_12185);
nor U12507 (N_12507,N_12319,N_12250);
nor U12508 (N_12508,N_12142,N_12367);
and U12509 (N_12509,N_12124,N_12166);
nor U12510 (N_12510,N_12076,N_12360);
or U12511 (N_12511,N_12145,N_12290);
and U12512 (N_12512,N_12109,N_12117);
or U12513 (N_12513,N_12184,N_12435);
or U12514 (N_12514,N_12235,N_12343);
or U12515 (N_12515,N_12474,N_12050);
or U12516 (N_12516,N_12439,N_12302);
nand U12517 (N_12517,N_12197,N_12297);
xnor U12518 (N_12518,N_12287,N_12432);
xnor U12519 (N_12519,N_12133,N_12424);
and U12520 (N_12520,N_12332,N_12260);
nand U12521 (N_12521,N_12266,N_12431);
or U12522 (N_12522,N_12233,N_12425);
and U12523 (N_12523,N_12144,N_12452);
or U12524 (N_12524,N_12062,N_12314);
and U12525 (N_12525,N_12085,N_12331);
and U12526 (N_12526,N_12322,N_12155);
nand U12527 (N_12527,N_12103,N_12087);
and U12528 (N_12528,N_12017,N_12213);
or U12529 (N_12529,N_12131,N_12460);
nand U12530 (N_12530,N_12323,N_12027);
or U12531 (N_12531,N_12053,N_12168);
nor U12532 (N_12532,N_12129,N_12450);
nand U12533 (N_12533,N_12299,N_12348);
xor U12534 (N_12534,N_12318,N_12019);
nor U12535 (N_12535,N_12304,N_12191);
and U12536 (N_12536,N_12040,N_12153);
nor U12537 (N_12537,N_12335,N_12437);
and U12538 (N_12538,N_12020,N_12383);
nand U12539 (N_12539,N_12081,N_12210);
and U12540 (N_12540,N_12342,N_12363);
nand U12541 (N_12541,N_12276,N_12405);
and U12542 (N_12542,N_12253,N_12070);
nor U12543 (N_12543,N_12067,N_12284);
or U12544 (N_12544,N_12089,N_12402);
nand U12545 (N_12545,N_12337,N_12024);
or U12546 (N_12546,N_12061,N_12420);
nor U12547 (N_12547,N_12119,N_12313);
or U12548 (N_12548,N_12308,N_12088);
nor U12549 (N_12549,N_12098,N_12060);
xor U12550 (N_12550,N_12388,N_12277);
xnor U12551 (N_12551,N_12366,N_12118);
nor U12552 (N_12552,N_12411,N_12303);
nand U12553 (N_12553,N_12056,N_12384);
xor U12554 (N_12554,N_12032,N_12486);
and U12555 (N_12555,N_12465,N_12028);
xnor U12556 (N_12556,N_12039,N_12334);
nand U12557 (N_12557,N_12030,N_12436);
nor U12558 (N_12558,N_12414,N_12125);
nor U12559 (N_12559,N_12312,N_12479);
nor U12560 (N_12560,N_12264,N_12338);
and U12561 (N_12561,N_12374,N_12396);
and U12562 (N_12562,N_12451,N_12150);
or U12563 (N_12563,N_12400,N_12358);
nand U12564 (N_12564,N_12014,N_12218);
nor U12565 (N_12565,N_12245,N_12341);
or U12566 (N_12566,N_12347,N_12079);
nor U12567 (N_12567,N_12357,N_12296);
nand U12568 (N_12568,N_12438,N_12468);
or U12569 (N_12569,N_12012,N_12256);
or U12570 (N_12570,N_12283,N_12391);
nor U12571 (N_12571,N_12491,N_12442);
nor U12572 (N_12572,N_12049,N_12324);
or U12573 (N_12573,N_12077,N_12057);
or U12574 (N_12574,N_12490,N_12230);
or U12575 (N_12575,N_12301,N_12138);
nand U12576 (N_12576,N_12418,N_12105);
or U12577 (N_12577,N_12237,N_12499);
and U12578 (N_12578,N_12373,N_12033);
nor U12579 (N_12579,N_12082,N_12380);
and U12580 (N_12580,N_12196,N_12139);
or U12581 (N_12581,N_12395,N_12226);
or U12582 (N_12582,N_12493,N_12170);
nand U12583 (N_12583,N_12010,N_12289);
or U12584 (N_12584,N_12035,N_12398);
nand U12585 (N_12585,N_12257,N_12204);
and U12586 (N_12586,N_12488,N_12065);
or U12587 (N_12587,N_12280,N_12158);
and U12588 (N_12588,N_12116,N_12201);
xnor U12589 (N_12589,N_12227,N_12455);
nand U12590 (N_12590,N_12228,N_12446);
or U12591 (N_12591,N_12059,N_12477);
nand U12592 (N_12592,N_12307,N_12454);
or U12593 (N_12593,N_12325,N_12052);
and U12594 (N_12594,N_12419,N_12270);
nand U12595 (N_12595,N_12372,N_12128);
xnor U12596 (N_12596,N_12494,N_12362);
nand U12597 (N_12597,N_12149,N_12249);
and U12598 (N_12598,N_12369,N_12206);
and U12599 (N_12599,N_12200,N_12444);
nand U12600 (N_12600,N_12108,N_12328);
nor U12601 (N_12601,N_12422,N_12397);
or U12602 (N_12602,N_12350,N_12263);
xor U12603 (N_12603,N_12058,N_12497);
and U12604 (N_12604,N_12173,N_12262);
and U12605 (N_12605,N_12234,N_12464);
nand U12606 (N_12606,N_12072,N_12271);
nand U12607 (N_12607,N_12169,N_12489);
nor U12608 (N_12608,N_12484,N_12187);
nand U12609 (N_12609,N_12154,N_12445);
nor U12610 (N_12610,N_12247,N_12006);
and U12611 (N_12611,N_12386,N_12433);
xnor U12612 (N_12612,N_12048,N_12399);
nand U12613 (N_12613,N_12045,N_12475);
and U12614 (N_12614,N_12194,N_12416);
nand U12615 (N_12615,N_12447,N_12458);
nand U12616 (N_12616,N_12147,N_12137);
nand U12617 (N_12617,N_12075,N_12333);
nand U12618 (N_12618,N_12102,N_12410);
nand U12619 (N_12619,N_12320,N_12162);
or U12620 (N_12620,N_12151,N_12143);
and U12621 (N_12621,N_12498,N_12326);
nor U12622 (N_12622,N_12344,N_12495);
nand U12623 (N_12623,N_12214,N_12037);
or U12624 (N_12624,N_12258,N_12159);
and U12625 (N_12625,N_12375,N_12174);
nor U12626 (N_12626,N_12066,N_12188);
nand U12627 (N_12627,N_12240,N_12121);
and U12628 (N_12628,N_12164,N_12345);
nand U12629 (N_12629,N_12036,N_12292);
or U12630 (N_12630,N_12195,N_12034);
nor U12631 (N_12631,N_12078,N_12252);
or U12632 (N_12632,N_12161,N_12005);
and U12633 (N_12633,N_12208,N_12127);
xnor U12634 (N_12634,N_12093,N_12272);
xnor U12635 (N_12635,N_12483,N_12219);
nor U12636 (N_12636,N_12055,N_12141);
and U12637 (N_12637,N_12244,N_12293);
nor U12638 (N_12638,N_12298,N_12346);
nor U12639 (N_12639,N_12094,N_12220);
and U12640 (N_12640,N_12286,N_12099);
nor U12641 (N_12641,N_12091,N_12275);
and U12642 (N_12642,N_12107,N_12243);
nor U12643 (N_12643,N_12354,N_12481);
nor U12644 (N_12644,N_12023,N_12090);
and U12645 (N_12645,N_12259,N_12086);
or U12646 (N_12646,N_12216,N_12111);
and U12647 (N_12647,N_12248,N_12156);
or U12648 (N_12648,N_12356,N_12393);
and U12649 (N_12649,N_12361,N_12008);
xor U12650 (N_12650,N_12406,N_12370);
nand U12651 (N_12651,N_12011,N_12123);
and U12652 (N_12652,N_12064,N_12122);
nor U12653 (N_12653,N_12267,N_12231);
and U12654 (N_12654,N_12434,N_12069);
nand U12655 (N_12655,N_12279,N_12378);
nor U12656 (N_12656,N_12215,N_12316);
nand U12657 (N_12657,N_12047,N_12013);
nand U12658 (N_12658,N_12015,N_12135);
and U12659 (N_12659,N_12232,N_12476);
nor U12660 (N_12660,N_12110,N_12209);
xnor U12661 (N_12661,N_12415,N_12001);
xor U12662 (N_12662,N_12310,N_12291);
xnor U12663 (N_12663,N_12413,N_12177);
or U12664 (N_12664,N_12251,N_12198);
and U12665 (N_12665,N_12407,N_12329);
nand U12666 (N_12666,N_12294,N_12261);
xnor U12667 (N_12667,N_12221,N_12295);
nor U12668 (N_12668,N_12182,N_12043);
or U12669 (N_12669,N_12171,N_12080);
nand U12670 (N_12670,N_12470,N_12007);
and U12671 (N_12671,N_12430,N_12134);
or U12672 (N_12672,N_12379,N_12496);
xnor U12673 (N_12673,N_12190,N_12466);
and U12674 (N_12674,N_12467,N_12440);
nor U12675 (N_12675,N_12146,N_12273);
xor U12676 (N_12676,N_12176,N_12385);
nor U12677 (N_12677,N_12478,N_12183);
xor U12678 (N_12678,N_12364,N_12038);
nand U12679 (N_12679,N_12355,N_12368);
xor U12680 (N_12680,N_12471,N_12207);
nand U12681 (N_12681,N_12469,N_12448);
or U12682 (N_12682,N_12051,N_12175);
and U12683 (N_12683,N_12462,N_12031);
nor U12684 (N_12684,N_12202,N_12239);
or U12685 (N_12685,N_12315,N_12157);
or U12686 (N_12686,N_12113,N_12120);
or U12687 (N_12687,N_12381,N_12212);
xnor U12688 (N_12688,N_12371,N_12282);
and U12689 (N_12689,N_12441,N_12163);
xor U12690 (N_12690,N_12428,N_12178);
nand U12691 (N_12691,N_12321,N_12401);
or U12692 (N_12692,N_12041,N_12106);
or U12693 (N_12693,N_12054,N_12172);
and U12694 (N_12694,N_12009,N_12309);
nand U12695 (N_12695,N_12193,N_12417);
nor U12696 (N_12696,N_12288,N_12306);
nor U12697 (N_12697,N_12365,N_12042);
and U12698 (N_12698,N_12376,N_12222);
or U12699 (N_12699,N_12268,N_12026);
nand U12700 (N_12700,N_12274,N_12068);
nor U12701 (N_12701,N_12217,N_12097);
or U12702 (N_12702,N_12349,N_12255);
nand U12703 (N_12703,N_12387,N_12100);
and U12704 (N_12704,N_12160,N_12317);
and U12705 (N_12705,N_12492,N_12095);
xor U12706 (N_12706,N_12046,N_12104);
and U12707 (N_12707,N_12223,N_12165);
or U12708 (N_12708,N_12018,N_12327);
and U12709 (N_12709,N_12203,N_12000);
nand U12710 (N_12710,N_12463,N_12389);
or U12711 (N_12711,N_12473,N_12179);
or U12712 (N_12712,N_12453,N_12152);
xnor U12713 (N_12713,N_12403,N_12487);
nor U12714 (N_12714,N_12285,N_12073);
nor U12715 (N_12715,N_12377,N_12242);
and U12716 (N_12716,N_12281,N_12167);
nand U12717 (N_12717,N_12269,N_12096);
and U12718 (N_12718,N_12429,N_12485);
nand U12719 (N_12719,N_12063,N_12225);
nand U12720 (N_12720,N_12071,N_12330);
nor U12721 (N_12721,N_12003,N_12189);
nor U12722 (N_12722,N_12025,N_12421);
nor U12723 (N_12723,N_12351,N_12022);
nand U12724 (N_12724,N_12112,N_12339);
or U12725 (N_12725,N_12426,N_12390);
nor U12726 (N_12726,N_12427,N_12101);
or U12727 (N_12727,N_12246,N_12181);
or U12728 (N_12728,N_12392,N_12136);
nor U12729 (N_12729,N_12449,N_12353);
and U12730 (N_12730,N_12459,N_12457);
nand U12731 (N_12731,N_12482,N_12409);
nor U12732 (N_12732,N_12408,N_12004);
or U12733 (N_12733,N_12205,N_12404);
nand U12734 (N_12734,N_12002,N_12461);
or U12735 (N_12735,N_12126,N_12311);
nor U12736 (N_12736,N_12084,N_12092);
nor U12737 (N_12737,N_12199,N_12115);
nor U12738 (N_12738,N_12423,N_12336);
nor U12739 (N_12739,N_12229,N_12021);
or U12740 (N_12740,N_12186,N_12300);
xor U12741 (N_12741,N_12265,N_12044);
and U12742 (N_12742,N_12083,N_12029);
or U12743 (N_12743,N_12480,N_12236);
nand U12744 (N_12744,N_12224,N_12132);
or U12745 (N_12745,N_12305,N_12382);
or U12746 (N_12746,N_12359,N_12114);
or U12747 (N_12747,N_12278,N_12238);
xor U12748 (N_12748,N_12241,N_12394);
nor U12749 (N_12749,N_12130,N_12211);
nand U12750 (N_12750,N_12337,N_12404);
and U12751 (N_12751,N_12160,N_12389);
nor U12752 (N_12752,N_12232,N_12491);
nand U12753 (N_12753,N_12398,N_12400);
or U12754 (N_12754,N_12310,N_12498);
or U12755 (N_12755,N_12138,N_12041);
xnor U12756 (N_12756,N_12363,N_12322);
nor U12757 (N_12757,N_12047,N_12470);
or U12758 (N_12758,N_12366,N_12023);
nand U12759 (N_12759,N_12121,N_12275);
nor U12760 (N_12760,N_12078,N_12242);
nand U12761 (N_12761,N_12178,N_12226);
and U12762 (N_12762,N_12133,N_12384);
and U12763 (N_12763,N_12424,N_12312);
and U12764 (N_12764,N_12018,N_12171);
or U12765 (N_12765,N_12413,N_12354);
nor U12766 (N_12766,N_12029,N_12194);
nand U12767 (N_12767,N_12058,N_12270);
xnor U12768 (N_12768,N_12019,N_12336);
nand U12769 (N_12769,N_12273,N_12294);
or U12770 (N_12770,N_12130,N_12230);
nand U12771 (N_12771,N_12385,N_12489);
or U12772 (N_12772,N_12188,N_12141);
nor U12773 (N_12773,N_12157,N_12203);
xnor U12774 (N_12774,N_12362,N_12394);
nand U12775 (N_12775,N_12360,N_12403);
or U12776 (N_12776,N_12449,N_12482);
nand U12777 (N_12777,N_12197,N_12102);
and U12778 (N_12778,N_12385,N_12428);
xor U12779 (N_12779,N_12005,N_12079);
nand U12780 (N_12780,N_12042,N_12014);
nand U12781 (N_12781,N_12015,N_12387);
and U12782 (N_12782,N_12186,N_12131);
or U12783 (N_12783,N_12114,N_12318);
nor U12784 (N_12784,N_12074,N_12230);
nor U12785 (N_12785,N_12357,N_12115);
or U12786 (N_12786,N_12074,N_12487);
nor U12787 (N_12787,N_12154,N_12467);
or U12788 (N_12788,N_12250,N_12235);
nand U12789 (N_12789,N_12077,N_12448);
and U12790 (N_12790,N_12194,N_12207);
or U12791 (N_12791,N_12102,N_12029);
or U12792 (N_12792,N_12247,N_12488);
and U12793 (N_12793,N_12066,N_12476);
nor U12794 (N_12794,N_12233,N_12266);
nor U12795 (N_12795,N_12468,N_12404);
nor U12796 (N_12796,N_12417,N_12387);
nand U12797 (N_12797,N_12292,N_12167);
and U12798 (N_12798,N_12179,N_12219);
nand U12799 (N_12799,N_12469,N_12273);
and U12800 (N_12800,N_12108,N_12224);
xor U12801 (N_12801,N_12447,N_12294);
and U12802 (N_12802,N_12059,N_12153);
xnor U12803 (N_12803,N_12388,N_12014);
or U12804 (N_12804,N_12017,N_12306);
xnor U12805 (N_12805,N_12136,N_12236);
xor U12806 (N_12806,N_12465,N_12136);
and U12807 (N_12807,N_12110,N_12102);
and U12808 (N_12808,N_12450,N_12364);
and U12809 (N_12809,N_12197,N_12173);
or U12810 (N_12810,N_12448,N_12349);
nor U12811 (N_12811,N_12069,N_12288);
or U12812 (N_12812,N_12353,N_12248);
xnor U12813 (N_12813,N_12054,N_12117);
or U12814 (N_12814,N_12005,N_12025);
or U12815 (N_12815,N_12447,N_12040);
nand U12816 (N_12816,N_12027,N_12102);
nand U12817 (N_12817,N_12156,N_12433);
and U12818 (N_12818,N_12084,N_12325);
xnor U12819 (N_12819,N_12107,N_12341);
and U12820 (N_12820,N_12207,N_12460);
nor U12821 (N_12821,N_12312,N_12197);
or U12822 (N_12822,N_12356,N_12197);
nand U12823 (N_12823,N_12183,N_12105);
and U12824 (N_12824,N_12049,N_12457);
nor U12825 (N_12825,N_12171,N_12490);
or U12826 (N_12826,N_12089,N_12420);
xor U12827 (N_12827,N_12193,N_12458);
or U12828 (N_12828,N_12314,N_12497);
and U12829 (N_12829,N_12379,N_12369);
and U12830 (N_12830,N_12249,N_12471);
xor U12831 (N_12831,N_12422,N_12320);
and U12832 (N_12832,N_12257,N_12404);
xor U12833 (N_12833,N_12445,N_12196);
or U12834 (N_12834,N_12469,N_12298);
nand U12835 (N_12835,N_12480,N_12359);
or U12836 (N_12836,N_12211,N_12113);
nand U12837 (N_12837,N_12470,N_12113);
and U12838 (N_12838,N_12481,N_12195);
and U12839 (N_12839,N_12467,N_12095);
or U12840 (N_12840,N_12381,N_12442);
or U12841 (N_12841,N_12281,N_12188);
or U12842 (N_12842,N_12444,N_12410);
or U12843 (N_12843,N_12203,N_12245);
and U12844 (N_12844,N_12407,N_12012);
nand U12845 (N_12845,N_12213,N_12022);
nor U12846 (N_12846,N_12262,N_12073);
nor U12847 (N_12847,N_12137,N_12033);
xor U12848 (N_12848,N_12124,N_12135);
or U12849 (N_12849,N_12247,N_12357);
and U12850 (N_12850,N_12466,N_12323);
nand U12851 (N_12851,N_12071,N_12308);
and U12852 (N_12852,N_12263,N_12167);
nor U12853 (N_12853,N_12451,N_12234);
nor U12854 (N_12854,N_12046,N_12335);
nor U12855 (N_12855,N_12374,N_12360);
nor U12856 (N_12856,N_12396,N_12006);
nand U12857 (N_12857,N_12182,N_12203);
nand U12858 (N_12858,N_12228,N_12477);
xnor U12859 (N_12859,N_12367,N_12289);
and U12860 (N_12860,N_12485,N_12223);
nand U12861 (N_12861,N_12199,N_12324);
nor U12862 (N_12862,N_12291,N_12137);
nor U12863 (N_12863,N_12115,N_12038);
nor U12864 (N_12864,N_12169,N_12363);
xnor U12865 (N_12865,N_12483,N_12186);
nand U12866 (N_12866,N_12439,N_12398);
nand U12867 (N_12867,N_12303,N_12031);
nor U12868 (N_12868,N_12029,N_12224);
and U12869 (N_12869,N_12428,N_12378);
nor U12870 (N_12870,N_12099,N_12257);
nand U12871 (N_12871,N_12100,N_12152);
nand U12872 (N_12872,N_12358,N_12217);
and U12873 (N_12873,N_12229,N_12350);
and U12874 (N_12874,N_12254,N_12248);
and U12875 (N_12875,N_12330,N_12218);
and U12876 (N_12876,N_12277,N_12202);
nor U12877 (N_12877,N_12495,N_12276);
and U12878 (N_12878,N_12400,N_12224);
and U12879 (N_12879,N_12336,N_12210);
and U12880 (N_12880,N_12243,N_12114);
or U12881 (N_12881,N_12443,N_12086);
or U12882 (N_12882,N_12327,N_12238);
xnor U12883 (N_12883,N_12321,N_12017);
nand U12884 (N_12884,N_12114,N_12344);
or U12885 (N_12885,N_12029,N_12321);
and U12886 (N_12886,N_12301,N_12315);
or U12887 (N_12887,N_12449,N_12360);
xnor U12888 (N_12888,N_12356,N_12434);
nor U12889 (N_12889,N_12446,N_12319);
nand U12890 (N_12890,N_12060,N_12394);
nand U12891 (N_12891,N_12457,N_12319);
nor U12892 (N_12892,N_12477,N_12036);
nand U12893 (N_12893,N_12180,N_12433);
and U12894 (N_12894,N_12240,N_12222);
or U12895 (N_12895,N_12423,N_12246);
or U12896 (N_12896,N_12316,N_12006);
or U12897 (N_12897,N_12054,N_12214);
or U12898 (N_12898,N_12051,N_12328);
nor U12899 (N_12899,N_12152,N_12136);
xor U12900 (N_12900,N_12191,N_12034);
nor U12901 (N_12901,N_12215,N_12244);
and U12902 (N_12902,N_12007,N_12345);
or U12903 (N_12903,N_12265,N_12259);
nand U12904 (N_12904,N_12253,N_12191);
and U12905 (N_12905,N_12467,N_12124);
nor U12906 (N_12906,N_12233,N_12151);
and U12907 (N_12907,N_12420,N_12234);
nand U12908 (N_12908,N_12350,N_12113);
nand U12909 (N_12909,N_12387,N_12315);
nand U12910 (N_12910,N_12290,N_12117);
and U12911 (N_12911,N_12291,N_12033);
nor U12912 (N_12912,N_12240,N_12092);
and U12913 (N_12913,N_12102,N_12145);
and U12914 (N_12914,N_12173,N_12285);
and U12915 (N_12915,N_12257,N_12413);
nand U12916 (N_12916,N_12314,N_12447);
nand U12917 (N_12917,N_12357,N_12002);
nand U12918 (N_12918,N_12223,N_12319);
or U12919 (N_12919,N_12381,N_12240);
and U12920 (N_12920,N_12472,N_12205);
or U12921 (N_12921,N_12450,N_12005);
and U12922 (N_12922,N_12286,N_12487);
nor U12923 (N_12923,N_12160,N_12465);
and U12924 (N_12924,N_12124,N_12152);
or U12925 (N_12925,N_12473,N_12429);
or U12926 (N_12926,N_12208,N_12115);
nor U12927 (N_12927,N_12465,N_12366);
nor U12928 (N_12928,N_12402,N_12303);
nand U12929 (N_12929,N_12086,N_12381);
or U12930 (N_12930,N_12084,N_12408);
and U12931 (N_12931,N_12271,N_12159);
nor U12932 (N_12932,N_12306,N_12405);
nand U12933 (N_12933,N_12281,N_12375);
nor U12934 (N_12934,N_12461,N_12050);
nand U12935 (N_12935,N_12097,N_12359);
nand U12936 (N_12936,N_12411,N_12155);
nor U12937 (N_12937,N_12324,N_12204);
nand U12938 (N_12938,N_12026,N_12246);
nand U12939 (N_12939,N_12232,N_12115);
nor U12940 (N_12940,N_12462,N_12161);
and U12941 (N_12941,N_12216,N_12187);
or U12942 (N_12942,N_12217,N_12173);
nor U12943 (N_12943,N_12275,N_12083);
nor U12944 (N_12944,N_12045,N_12364);
nor U12945 (N_12945,N_12137,N_12043);
or U12946 (N_12946,N_12137,N_12245);
and U12947 (N_12947,N_12249,N_12170);
and U12948 (N_12948,N_12222,N_12466);
nand U12949 (N_12949,N_12359,N_12043);
or U12950 (N_12950,N_12396,N_12460);
or U12951 (N_12951,N_12423,N_12008);
nor U12952 (N_12952,N_12077,N_12074);
or U12953 (N_12953,N_12056,N_12196);
or U12954 (N_12954,N_12353,N_12356);
nand U12955 (N_12955,N_12404,N_12044);
and U12956 (N_12956,N_12163,N_12264);
nor U12957 (N_12957,N_12257,N_12006);
nand U12958 (N_12958,N_12380,N_12057);
or U12959 (N_12959,N_12116,N_12400);
or U12960 (N_12960,N_12260,N_12353);
and U12961 (N_12961,N_12324,N_12296);
nor U12962 (N_12962,N_12224,N_12001);
or U12963 (N_12963,N_12216,N_12021);
or U12964 (N_12964,N_12027,N_12101);
or U12965 (N_12965,N_12265,N_12130);
and U12966 (N_12966,N_12299,N_12232);
or U12967 (N_12967,N_12049,N_12399);
or U12968 (N_12968,N_12047,N_12020);
nor U12969 (N_12969,N_12141,N_12427);
nand U12970 (N_12970,N_12296,N_12005);
nand U12971 (N_12971,N_12451,N_12394);
and U12972 (N_12972,N_12190,N_12158);
and U12973 (N_12973,N_12424,N_12092);
xnor U12974 (N_12974,N_12098,N_12457);
nor U12975 (N_12975,N_12412,N_12382);
nand U12976 (N_12976,N_12039,N_12467);
nand U12977 (N_12977,N_12259,N_12274);
nor U12978 (N_12978,N_12069,N_12303);
nand U12979 (N_12979,N_12294,N_12198);
and U12980 (N_12980,N_12010,N_12216);
xnor U12981 (N_12981,N_12343,N_12163);
xor U12982 (N_12982,N_12069,N_12119);
and U12983 (N_12983,N_12119,N_12487);
and U12984 (N_12984,N_12078,N_12429);
nor U12985 (N_12985,N_12213,N_12112);
nor U12986 (N_12986,N_12030,N_12148);
or U12987 (N_12987,N_12109,N_12388);
nor U12988 (N_12988,N_12373,N_12029);
nand U12989 (N_12989,N_12139,N_12367);
or U12990 (N_12990,N_12277,N_12108);
and U12991 (N_12991,N_12293,N_12443);
or U12992 (N_12992,N_12457,N_12085);
xor U12993 (N_12993,N_12406,N_12070);
or U12994 (N_12994,N_12310,N_12325);
nor U12995 (N_12995,N_12407,N_12401);
xor U12996 (N_12996,N_12461,N_12009);
and U12997 (N_12997,N_12262,N_12245);
or U12998 (N_12998,N_12270,N_12008);
nand U12999 (N_12999,N_12401,N_12215);
xnor U13000 (N_13000,N_12772,N_12839);
nor U13001 (N_13001,N_12722,N_12926);
nor U13002 (N_13002,N_12723,N_12780);
nand U13003 (N_13003,N_12909,N_12822);
nor U13004 (N_13004,N_12762,N_12883);
nand U13005 (N_13005,N_12749,N_12713);
nor U13006 (N_13006,N_12715,N_12670);
or U13007 (N_13007,N_12934,N_12878);
nor U13008 (N_13008,N_12577,N_12704);
and U13009 (N_13009,N_12565,N_12532);
nand U13010 (N_13010,N_12785,N_12967);
or U13011 (N_13011,N_12993,N_12694);
and U13012 (N_13012,N_12553,N_12628);
and U13013 (N_13013,N_12684,N_12851);
or U13014 (N_13014,N_12793,N_12691);
xor U13015 (N_13015,N_12576,N_12736);
and U13016 (N_13016,N_12697,N_12900);
or U13017 (N_13017,N_12580,N_12719);
and U13018 (N_13018,N_12817,N_12929);
nand U13019 (N_13019,N_12591,N_12999);
nor U13020 (N_13020,N_12972,N_12585);
nand U13021 (N_13021,N_12826,N_12709);
xor U13022 (N_13022,N_12874,N_12703);
and U13023 (N_13023,N_12562,N_12796);
and U13024 (N_13024,N_12634,N_12862);
and U13025 (N_13025,N_12905,N_12799);
or U13026 (N_13026,N_12743,N_12931);
nand U13027 (N_13027,N_12551,N_12728);
xnor U13028 (N_13028,N_12604,N_12756);
and U13029 (N_13029,N_12849,N_12695);
or U13030 (N_13030,N_12998,N_12813);
nor U13031 (N_13031,N_12599,N_12659);
or U13032 (N_13032,N_12730,N_12942);
and U13033 (N_13033,N_12665,N_12525);
or U13034 (N_13034,N_12613,N_12920);
nand U13035 (N_13035,N_12600,N_12984);
and U13036 (N_13036,N_12584,N_12768);
nand U13037 (N_13037,N_12891,N_12877);
xnor U13038 (N_13038,N_12852,N_12579);
nor U13039 (N_13039,N_12540,N_12733);
nor U13040 (N_13040,N_12823,N_12569);
and U13041 (N_13041,N_12609,N_12753);
xnor U13042 (N_13042,N_12986,N_12821);
nand U13043 (N_13043,N_12507,N_12936);
or U13044 (N_13044,N_12661,N_12593);
or U13045 (N_13045,N_12519,N_12650);
nor U13046 (N_13046,N_12963,N_12624);
xnor U13047 (N_13047,N_12892,N_12524);
xor U13048 (N_13048,N_12872,N_12979);
nor U13049 (N_13049,N_12784,N_12549);
nand U13050 (N_13050,N_12649,N_12790);
or U13051 (N_13051,N_12651,N_12786);
nand U13052 (N_13052,N_12542,N_12607);
or U13053 (N_13053,N_12528,N_12969);
xnor U13054 (N_13054,N_12976,N_12810);
nand U13055 (N_13055,N_12829,N_12781);
and U13056 (N_13056,N_12667,N_12882);
nor U13057 (N_13057,N_12676,N_12933);
nand U13058 (N_13058,N_12958,N_12923);
nand U13059 (N_13059,N_12720,N_12671);
xnor U13060 (N_13060,N_12792,N_12721);
or U13061 (N_13061,N_12800,N_12991);
nand U13062 (N_13062,N_12625,N_12737);
xnor U13063 (N_13063,N_12603,N_12914);
xnor U13064 (N_13064,N_12505,N_12937);
nand U13065 (N_13065,N_12701,N_12775);
or U13066 (N_13066,N_12645,N_12702);
or U13067 (N_13067,N_12746,N_12765);
or U13068 (N_13068,N_12724,N_12951);
or U13069 (N_13069,N_12754,N_12961);
nand U13070 (N_13070,N_12994,N_12547);
or U13071 (N_13071,N_12825,N_12896);
nor U13072 (N_13072,N_12752,N_12601);
nand U13073 (N_13073,N_12582,N_12731);
and U13074 (N_13074,N_12848,N_12708);
and U13075 (N_13075,N_12666,N_12847);
and U13076 (N_13076,N_12949,N_12757);
nand U13077 (N_13077,N_12930,N_12558);
and U13078 (N_13078,N_12988,N_12578);
and U13079 (N_13079,N_12637,N_12857);
nand U13080 (N_13080,N_12870,N_12617);
nor U13081 (N_13081,N_12619,N_12801);
or U13082 (N_13082,N_12980,N_12924);
nor U13083 (N_13083,N_12554,N_12971);
and U13084 (N_13084,N_12621,N_12950);
and U13085 (N_13085,N_12606,N_12517);
or U13086 (N_13086,N_12560,N_12876);
and U13087 (N_13087,N_12598,N_12778);
nand U13088 (N_13088,N_12592,N_12614);
and U13089 (N_13089,N_12534,N_12710);
or U13090 (N_13090,N_12858,N_12777);
or U13091 (N_13091,N_12643,N_12788);
nor U13092 (N_13092,N_12831,N_12644);
and U13093 (N_13093,N_12654,N_12820);
and U13094 (N_13094,N_12818,N_12631);
or U13095 (N_13095,N_12873,N_12632);
xor U13096 (N_13096,N_12902,N_12764);
and U13097 (N_13097,N_12975,N_12866);
xor U13098 (N_13098,N_12843,N_12610);
or U13099 (N_13099,N_12575,N_12978);
nand U13100 (N_13100,N_12954,N_12875);
and U13101 (N_13101,N_12987,N_12732);
and U13102 (N_13102,N_12888,N_12716);
and U13103 (N_13103,N_12734,N_12544);
nand U13104 (N_13104,N_12660,N_12844);
and U13105 (N_13105,N_12537,N_12652);
nor U13106 (N_13106,N_12559,N_12539);
or U13107 (N_13107,N_12512,N_12895);
or U13108 (N_13108,N_12504,N_12804);
and U13109 (N_13109,N_12566,N_12726);
nor U13110 (N_13110,N_12769,N_12770);
nand U13111 (N_13111,N_12766,N_12612);
and U13112 (N_13112,N_12767,N_12911);
nor U13113 (N_13113,N_12832,N_12861);
or U13114 (N_13114,N_12518,N_12982);
and U13115 (N_13115,N_12912,N_12646);
nor U13116 (N_13116,N_12538,N_12906);
and U13117 (N_13117,N_12957,N_12513);
nand U13118 (N_13118,N_12570,N_12529);
or U13119 (N_13119,N_12618,N_12791);
and U13120 (N_13120,N_12620,N_12556);
or U13121 (N_13121,N_12572,N_12623);
or U13122 (N_13122,N_12904,N_12755);
xnor U13123 (N_13123,N_12997,N_12889);
nand U13124 (N_13124,N_12741,N_12630);
and U13125 (N_13125,N_12738,N_12992);
and U13126 (N_13126,N_12955,N_12776);
or U13127 (N_13127,N_12946,N_12700);
and U13128 (N_13128,N_12989,N_12927);
nor U13129 (N_13129,N_12859,N_12658);
or U13130 (N_13130,N_12536,N_12589);
nor U13131 (N_13131,N_12548,N_12583);
or U13132 (N_13132,N_12836,N_12869);
or U13133 (N_13133,N_12677,N_12587);
nor U13134 (N_13134,N_12729,N_12985);
nand U13135 (N_13135,N_12655,N_12674);
nand U13136 (N_13136,N_12952,N_12682);
nand U13137 (N_13137,N_12939,N_12595);
or U13138 (N_13138,N_12845,N_12712);
and U13139 (N_13139,N_12615,N_12932);
and U13140 (N_13140,N_12867,N_12835);
and U13141 (N_13141,N_12514,N_12626);
nor U13142 (N_13142,N_12675,N_12885);
or U13143 (N_13143,N_12699,N_12917);
and U13144 (N_13144,N_12500,N_12616);
nor U13145 (N_13145,N_12640,N_12627);
or U13146 (N_13146,N_12856,N_12956);
and U13147 (N_13147,N_12664,N_12501);
or U13148 (N_13148,N_12983,N_12838);
nor U13149 (N_13149,N_12725,N_12629);
xnor U13150 (N_13150,N_12745,N_12531);
and U13151 (N_13151,N_12890,N_12510);
nor U13152 (N_13152,N_12568,N_12879);
nor U13153 (N_13153,N_12899,N_12779);
or U13154 (N_13154,N_12901,N_12639);
nand U13155 (N_13155,N_12865,N_12760);
nand U13156 (N_13156,N_12802,N_12679);
nand U13157 (N_13157,N_12960,N_12990);
or U13158 (N_13158,N_12508,N_12968);
nor U13159 (N_13159,N_12657,N_12693);
and U13160 (N_13160,N_12594,N_12633);
nand U13161 (N_13161,N_12806,N_12515);
nand U13162 (N_13162,N_12893,N_12908);
xnor U13163 (N_13163,N_12506,N_12871);
nand U13164 (N_13164,N_12744,N_12509);
or U13165 (N_13165,N_12748,N_12868);
and U13166 (N_13166,N_12561,N_12855);
xor U13167 (N_13167,N_12688,N_12678);
or U13168 (N_13168,N_12663,N_12673);
or U13169 (N_13169,N_12550,N_12794);
nand U13170 (N_13170,N_12846,N_12530);
or U13171 (N_13171,N_12681,N_12687);
xor U13172 (N_13172,N_12842,N_12683);
nand U13173 (N_13173,N_12965,N_12668);
nor U13174 (N_13174,N_12915,N_12834);
nand U13175 (N_13175,N_12918,N_12742);
xnor U13176 (N_13176,N_12680,N_12763);
nand U13177 (N_13177,N_12921,N_12916);
or U13178 (N_13178,N_12840,N_12622);
and U13179 (N_13179,N_12546,N_12970);
or U13180 (N_13180,N_12789,N_12574);
or U13181 (N_13181,N_12773,N_12837);
nor U13182 (N_13182,N_12833,N_12698);
or U13183 (N_13183,N_12611,N_12692);
nand U13184 (N_13184,N_12907,N_12995);
nand U13185 (N_13185,N_12966,N_12656);
or U13186 (N_13186,N_12647,N_12642);
nor U13187 (N_13187,N_12805,N_12581);
or U13188 (N_13188,N_12571,N_12819);
and U13189 (N_13189,N_12555,N_12925);
nor U13190 (N_13190,N_12543,N_12814);
xnor U13191 (N_13191,N_12945,N_12567);
nor U13192 (N_13192,N_12535,N_12953);
xor U13193 (N_13193,N_12827,N_12783);
and U13194 (N_13194,N_12758,N_12830);
and U13195 (N_13195,N_12586,N_12897);
or U13196 (N_13196,N_12964,N_12850);
nand U13197 (N_13197,N_12520,N_12811);
and U13198 (N_13198,N_12863,N_12841);
or U13199 (N_13199,N_12941,N_12910);
nand U13200 (N_13200,N_12714,N_12761);
or U13201 (N_13201,N_12808,N_12884);
and U13202 (N_13202,N_12774,N_12935);
or U13203 (N_13203,N_12635,N_12602);
or U13204 (N_13204,N_12944,N_12854);
nor U13205 (N_13205,N_12913,N_12959);
nand U13206 (N_13206,N_12807,N_12686);
nand U13207 (N_13207,N_12798,N_12727);
or U13208 (N_13208,N_12689,N_12662);
nand U13209 (N_13209,N_12718,N_12669);
nor U13210 (N_13210,N_12881,N_12894);
nand U13211 (N_13211,N_12588,N_12564);
or U13212 (N_13212,N_12853,N_12545);
xor U13213 (N_13213,N_12739,N_12922);
or U13214 (N_13214,N_12809,N_12740);
and U13215 (N_13215,N_12940,N_12685);
xnor U13216 (N_13216,N_12563,N_12672);
and U13217 (N_13217,N_12973,N_12750);
nand U13218 (N_13218,N_12511,N_12747);
or U13219 (N_13219,N_12636,N_12977);
nand U13220 (N_13220,N_12717,N_12533);
or U13221 (N_13221,N_12596,N_12981);
or U13222 (N_13222,N_12597,N_12690);
nand U13223 (N_13223,N_12903,N_12938);
xor U13224 (N_13224,N_12557,N_12526);
or U13225 (N_13225,N_12735,N_12919);
nor U13226 (N_13226,N_12706,N_12797);
nand U13227 (N_13227,N_12523,N_12787);
nand U13228 (N_13228,N_12974,N_12962);
and U13229 (N_13229,N_12887,N_12608);
nand U13230 (N_13230,N_12812,N_12707);
nor U13231 (N_13231,N_12996,N_12880);
nor U13232 (N_13232,N_12816,N_12503);
xnor U13233 (N_13233,N_12527,N_12815);
and U13234 (N_13234,N_12541,N_12860);
or U13235 (N_13235,N_12521,N_12696);
or U13236 (N_13236,N_12947,N_12803);
or U13237 (N_13237,N_12552,N_12782);
nor U13238 (N_13238,N_12590,N_12898);
and U13239 (N_13239,N_12516,N_12864);
nand U13240 (N_13240,N_12573,N_12641);
and U13241 (N_13241,N_12522,N_12648);
or U13242 (N_13242,N_12928,N_12705);
and U13243 (N_13243,N_12638,N_12771);
xor U13244 (N_13244,N_12502,N_12824);
or U13245 (N_13245,N_12886,N_12605);
nor U13246 (N_13246,N_12828,N_12948);
nand U13247 (N_13247,N_12759,N_12943);
nor U13248 (N_13248,N_12653,N_12795);
xor U13249 (N_13249,N_12751,N_12711);
or U13250 (N_13250,N_12666,N_12539);
nor U13251 (N_13251,N_12920,N_12850);
and U13252 (N_13252,N_12537,N_12559);
nor U13253 (N_13253,N_12741,N_12895);
nand U13254 (N_13254,N_12936,N_12845);
and U13255 (N_13255,N_12512,N_12923);
nor U13256 (N_13256,N_12669,N_12986);
nor U13257 (N_13257,N_12523,N_12912);
nand U13258 (N_13258,N_12686,N_12991);
nor U13259 (N_13259,N_12908,N_12781);
nand U13260 (N_13260,N_12576,N_12503);
nand U13261 (N_13261,N_12619,N_12811);
nand U13262 (N_13262,N_12758,N_12614);
nor U13263 (N_13263,N_12778,N_12507);
or U13264 (N_13264,N_12662,N_12693);
nor U13265 (N_13265,N_12582,N_12889);
or U13266 (N_13266,N_12926,N_12622);
xnor U13267 (N_13267,N_12825,N_12778);
or U13268 (N_13268,N_12938,N_12968);
nand U13269 (N_13269,N_12980,N_12578);
or U13270 (N_13270,N_12953,N_12611);
nor U13271 (N_13271,N_12922,N_12528);
and U13272 (N_13272,N_12529,N_12644);
nor U13273 (N_13273,N_12840,N_12633);
and U13274 (N_13274,N_12847,N_12792);
xor U13275 (N_13275,N_12616,N_12745);
nand U13276 (N_13276,N_12505,N_12910);
or U13277 (N_13277,N_12813,N_12908);
nand U13278 (N_13278,N_12509,N_12587);
or U13279 (N_13279,N_12898,N_12587);
xor U13280 (N_13280,N_12787,N_12581);
and U13281 (N_13281,N_12831,N_12519);
nand U13282 (N_13282,N_12603,N_12755);
or U13283 (N_13283,N_12793,N_12960);
or U13284 (N_13284,N_12790,N_12954);
and U13285 (N_13285,N_12788,N_12688);
nand U13286 (N_13286,N_12529,N_12900);
xnor U13287 (N_13287,N_12879,N_12692);
nand U13288 (N_13288,N_12529,N_12987);
and U13289 (N_13289,N_12737,N_12890);
nor U13290 (N_13290,N_12538,N_12712);
nand U13291 (N_13291,N_12836,N_12961);
nand U13292 (N_13292,N_12517,N_12623);
nand U13293 (N_13293,N_12585,N_12547);
nand U13294 (N_13294,N_12620,N_12653);
and U13295 (N_13295,N_12728,N_12725);
and U13296 (N_13296,N_12944,N_12920);
nor U13297 (N_13297,N_12727,N_12693);
and U13298 (N_13298,N_12678,N_12532);
or U13299 (N_13299,N_12553,N_12905);
and U13300 (N_13300,N_12946,N_12565);
nor U13301 (N_13301,N_12784,N_12765);
or U13302 (N_13302,N_12941,N_12969);
and U13303 (N_13303,N_12562,N_12876);
and U13304 (N_13304,N_12990,N_12619);
nor U13305 (N_13305,N_12946,N_12504);
nor U13306 (N_13306,N_12861,N_12855);
or U13307 (N_13307,N_12958,N_12829);
and U13308 (N_13308,N_12822,N_12972);
and U13309 (N_13309,N_12900,N_12985);
and U13310 (N_13310,N_12517,N_12983);
or U13311 (N_13311,N_12879,N_12554);
and U13312 (N_13312,N_12723,N_12756);
and U13313 (N_13313,N_12603,N_12754);
nor U13314 (N_13314,N_12703,N_12559);
nor U13315 (N_13315,N_12509,N_12897);
and U13316 (N_13316,N_12668,N_12796);
or U13317 (N_13317,N_12696,N_12575);
and U13318 (N_13318,N_12569,N_12501);
or U13319 (N_13319,N_12510,N_12733);
nand U13320 (N_13320,N_12623,N_12858);
nand U13321 (N_13321,N_12907,N_12542);
xnor U13322 (N_13322,N_12825,N_12518);
or U13323 (N_13323,N_12639,N_12837);
nor U13324 (N_13324,N_12774,N_12561);
or U13325 (N_13325,N_12886,N_12816);
nor U13326 (N_13326,N_12795,N_12757);
or U13327 (N_13327,N_12818,N_12562);
and U13328 (N_13328,N_12527,N_12856);
or U13329 (N_13329,N_12881,N_12915);
nor U13330 (N_13330,N_12955,N_12555);
and U13331 (N_13331,N_12879,N_12998);
nand U13332 (N_13332,N_12859,N_12828);
nand U13333 (N_13333,N_12973,N_12783);
and U13334 (N_13334,N_12789,N_12591);
nor U13335 (N_13335,N_12862,N_12587);
nor U13336 (N_13336,N_12874,N_12513);
or U13337 (N_13337,N_12629,N_12914);
nand U13338 (N_13338,N_12810,N_12774);
nor U13339 (N_13339,N_12758,N_12619);
nor U13340 (N_13340,N_12669,N_12586);
nor U13341 (N_13341,N_12591,N_12858);
xnor U13342 (N_13342,N_12685,N_12760);
or U13343 (N_13343,N_12580,N_12838);
nand U13344 (N_13344,N_12896,N_12757);
xor U13345 (N_13345,N_12749,N_12902);
or U13346 (N_13346,N_12932,N_12514);
and U13347 (N_13347,N_12770,N_12536);
and U13348 (N_13348,N_12999,N_12811);
nor U13349 (N_13349,N_12506,N_12880);
nor U13350 (N_13350,N_12897,N_12759);
xnor U13351 (N_13351,N_12631,N_12974);
nand U13352 (N_13352,N_12795,N_12840);
nor U13353 (N_13353,N_12683,N_12694);
nand U13354 (N_13354,N_12601,N_12988);
and U13355 (N_13355,N_12966,N_12756);
nand U13356 (N_13356,N_12836,N_12658);
or U13357 (N_13357,N_12798,N_12559);
or U13358 (N_13358,N_12603,N_12996);
and U13359 (N_13359,N_12958,N_12613);
nor U13360 (N_13360,N_12613,N_12886);
nand U13361 (N_13361,N_12610,N_12713);
and U13362 (N_13362,N_12916,N_12583);
or U13363 (N_13363,N_12952,N_12944);
nor U13364 (N_13364,N_12504,N_12874);
or U13365 (N_13365,N_12513,N_12930);
and U13366 (N_13366,N_12516,N_12738);
nor U13367 (N_13367,N_12728,N_12623);
and U13368 (N_13368,N_12657,N_12627);
and U13369 (N_13369,N_12987,N_12867);
and U13370 (N_13370,N_12590,N_12966);
nand U13371 (N_13371,N_12920,N_12719);
and U13372 (N_13372,N_12992,N_12911);
and U13373 (N_13373,N_12912,N_12791);
or U13374 (N_13374,N_12728,N_12659);
and U13375 (N_13375,N_12502,N_12677);
nor U13376 (N_13376,N_12615,N_12622);
nand U13377 (N_13377,N_12865,N_12897);
nor U13378 (N_13378,N_12564,N_12967);
nand U13379 (N_13379,N_12879,N_12733);
or U13380 (N_13380,N_12728,N_12895);
and U13381 (N_13381,N_12693,N_12950);
or U13382 (N_13382,N_12605,N_12819);
nor U13383 (N_13383,N_12908,N_12792);
xor U13384 (N_13384,N_12612,N_12611);
nand U13385 (N_13385,N_12738,N_12880);
or U13386 (N_13386,N_12551,N_12954);
and U13387 (N_13387,N_12700,N_12768);
and U13388 (N_13388,N_12934,N_12955);
or U13389 (N_13389,N_12901,N_12882);
or U13390 (N_13390,N_12560,N_12634);
nor U13391 (N_13391,N_12894,N_12991);
or U13392 (N_13392,N_12666,N_12926);
or U13393 (N_13393,N_12759,N_12710);
nand U13394 (N_13394,N_12724,N_12709);
or U13395 (N_13395,N_12602,N_12826);
nand U13396 (N_13396,N_12858,N_12700);
nand U13397 (N_13397,N_12934,N_12954);
or U13398 (N_13398,N_12952,N_12780);
and U13399 (N_13399,N_12549,N_12595);
or U13400 (N_13400,N_12833,N_12581);
nor U13401 (N_13401,N_12938,N_12808);
nor U13402 (N_13402,N_12593,N_12834);
and U13403 (N_13403,N_12638,N_12858);
nor U13404 (N_13404,N_12579,N_12566);
and U13405 (N_13405,N_12985,N_12758);
and U13406 (N_13406,N_12663,N_12788);
and U13407 (N_13407,N_12986,N_12994);
nand U13408 (N_13408,N_12557,N_12517);
or U13409 (N_13409,N_12932,N_12638);
xnor U13410 (N_13410,N_12874,N_12752);
nand U13411 (N_13411,N_12559,N_12928);
nor U13412 (N_13412,N_12615,N_12575);
nor U13413 (N_13413,N_12742,N_12952);
nand U13414 (N_13414,N_12594,N_12934);
xnor U13415 (N_13415,N_12999,N_12832);
and U13416 (N_13416,N_12980,N_12527);
nor U13417 (N_13417,N_12526,N_12601);
xor U13418 (N_13418,N_12527,N_12970);
or U13419 (N_13419,N_12555,N_12978);
and U13420 (N_13420,N_12648,N_12958);
nand U13421 (N_13421,N_12816,N_12913);
and U13422 (N_13422,N_12659,N_12561);
nor U13423 (N_13423,N_12885,N_12629);
nor U13424 (N_13424,N_12544,N_12636);
nor U13425 (N_13425,N_12899,N_12675);
and U13426 (N_13426,N_12835,N_12695);
xor U13427 (N_13427,N_12703,N_12604);
and U13428 (N_13428,N_12866,N_12783);
nor U13429 (N_13429,N_12618,N_12697);
and U13430 (N_13430,N_12715,N_12578);
xor U13431 (N_13431,N_12503,N_12745);
or U13432 (N_13432,N_12718,N_12813);
and U13433 (N_13433,N_12652,N_12573);
or U13434 (N_13434,N_12880,N_12693);
or U13435 (N_13435,N_12634,N_12648);
nand U13436 (N_13436,N_12525,N_12791);
nor U13437 (N_13437,N_12865,N_12874);
nor U13438 (N_13438,N_12869,N_12871);
or U13439 (N_13439,N_12879,N_12653);
or U13440 (N_13440,N_12520,N_12609);
and U13441 (N_13441,N_12788,N_12539);
xnor U13442 (N_13442,N_12764,N_12540);
or U13443 (N_13443,N_12526,N_12826);
nor U13444 (N_13444,N_12816,N_12649);
or U13445 (N_13445,N_12791,N_12888);
xnor U13446 (N_13446,N_12549,N_12850);
nand U13447 (N_13447,N_12566,N_12899);
and U13448 (N_13448,N_12678,N_12514);
nor U13449 (N_13449,N_12829,N_12963);
nor U13450 (N_13450,N_12840,N_12863);
and U13451 (N_13451,N_12540,N_12736);
or U13452 (N_13452,N_12733,N_12729);
nor U13453 (N_13453,N_12574,N_12991);
nor U13454 (N_13454,N_12754,N_12602);
or U13455 (N_13455,N_12874,N_12819);
or U13456 (N_13456,N_12902,N_12551);
nand U13457 (N_13457,N_12984,N_12644);
nand U13458 (N_13458,N_12559,N_12602);
nand U13459 (N_13459,N_12744,N_12803);
nand U13460 (N_13460,N_12641,N_12824);
or U13461 (N_13461,N_12533,N_12620);
and U13462 (N_13462,N_12665,N_12746);
nand U13463 (N_13463,N_12911,N_12822);
nand U13464 (N_13464,N_12680,N_12574);
nor U13465 (N_13465,N_12836,N_12745);
and U13466 (N_13466,N_12566,N_12880);
nor U13467 (N_13467,N_12756,N_12835);
or U13468 (N_13468,N_12581,N_12685);
or U13469 (N_13469,N_12965,N_12948);
and U13470 (N_13470,N_12613,N_12948);
nor U13471 (N_13471,N_12684,N_12760);
and U13472 (N_13472,N_12799,N_12949);
xnor U13473 (N_13473,N_12829,N_12802);
and U13474 (N_13474,N_12716,N_12648);
xnor U13475 (N_13475,N_12645,N_12741);
nor U13476 (N_13476,N_12606,N_12747);
nor U13477 (N_13477,N_12575,N_12827);
nor U13478 (N_13478,N_12663,N_12918);
or U13479 (N_13479,N_12654,N_12763);
and U13480 (N_13480,N_12666,N_12902);
and U13481 (N_13481,N_12592,N_12716);
and U13482 (N_13482,N_12708,N_12692);
xor U13483 (N_13483,N_12948,N_12706);
nand U13484 (N_13484,N_12543,N_12794);
nor U13485 (N_13485,N_12715,N_12771);
nand U13486 (N_13486,N_12612,N_12575);
nand U13487 (N_13487,N_12929,N_12846);
nand U13488 (N_13488,N_12986,N_12918);
nor U13489 (N_13489,N_12949,N_12785);
or U13490 (N_13490,N_12628,N_12790);
or U13491 (N_13491,N_12875,N_12747);
nor U13492 (N_13492,N_12522,N_12632);
and U13493 (N_13493,N_12686,N_12774);
xnor U13494 (N_13494,N_12583,N_12925);
nand U13495 (N_13495,N_12619,N_12640);
and U13496 (N_13496,N_12904,N_12546);
or U13497 (N_13497,N_12898,N_12994);
nor U13498 (N_13498,N_12798,N_12761);
nand U13499 (N_13499,N_12511,N_12534);
and U13500 (N_13500,N_13354,N_13493);
nor U13501 (N_13501,N_13148,N_13463);
nand U13502 (N_13502,N_13486,N_13136);
and U13503 (N_13503,N_13280,N_13288);
xnor U13504 (N_13504,N_13081,N_13255);
and U13505 (N_13505,N_13012,N_13079);
xnor U13506 (N_13506,N_13004,N_13165);
and U13507 (N_13507,N_13097,N_13343);
or U13508 (N_13508,N_13202,N_13472);
or U13509 (N_13509,N_13241,N_13240);
nand U13510 (N_13510,N_13294,N_13145);
xnor U13511 (N_13511,N_13268,N_13398);
nor U13512 (N_13512,N_13428,N_13190);
and U13513 (N_13513,N_13408,N_13490);
or U13514 (N_13514,N_13159,N_13309);
nor U13515 (N_13515,N_13313,N_13312);
and U13516 (N_13516,N_13096,N_13266);
and U13517 (N_13517,N_13410,N_13073);
nand U13518 (N_13518,N_13456,N_13392);
and U13519 (N_13519,N_13495,N_13088);
or U13520 (N_13520,N_13386,N_13494);
nand U13521 (N_13521,N_13066,N_13361);
and U13522 (N_13522,N_13439,N_13427);
nor U13523 (N_13523,N_13483,N_13184);
and U13524 (N_13524,N_13417,N_13158);
and U13525 (N_13525,N_13450,N_13496);
or U13526 (N_13526,N_13037,N_13282);
and U13527 (N_13527,N_13185,N_13462);
nand U13528 (N_13528,N_13230,N_13247);
xnor U13529 (N_13529,N_13084,N_13388);
nand U13530 (N_13530,N_13470,N_13074);
and U13531 (N_13531,N_13090,N_13194);
nor U13532 (N_13532,N_13203,N_13444);
nand U13533 (N_13533,N_13337,N_13479);
xnor U13534 (N_13534,N_13039,N_13369);
nand U13535 (N_13535,N_13395,N_13347);
xor U13536 (N_13536,N_13429,N_13433);
nand U13537 (N_13537,N_13334,N_13476);
nor U13538 (N_13538,N_13305,N_13344);
nor U13539 (N_13539,N_13272,N_13466);
nor U13540 (N_13540,N_13061,N_13100);
nor U13541 (N_13541,N_13001,N_13289);
nand U13542 (N_13542,N_13278,N_13024);
xor U13543 (N_13543,N_13403,N_13436);
or U13544 (N_13544,N_13207,N_13359);
or U13545 (N_13545,N_13011,N_13155);
or U13546 (N_13546,N_13365,N_13364);
and U13547 (N_13547,N_13105,N_13258);
or U13548 (N_13548,N_13394,N_13426);
and U13549 (N_13549,N_13209,N_13254);
nand U13550 (N_13550,N_13380,N_13201);
and U13551 (N_13551,N_13414,N_13296);
nor U13552 (N_13552,N_13485,N_13446);
nand U13553 (N_13553,N_13242,N_13325);
xor U13554 (N_13554,N_13431,N_13409);
and U13555 (N_13555,N_13021,N_13089);
nand U13556 (N_13556,N_13250,N_13009);
nand U13557 (N_13557,N_13323,N_13251);
or U13558 (N_13558,N_13285,N_13437);
and U13559 (N_13559,N_13477,N_13357);
nand U13560 (N_13560,N_13176,N_13290);
nand U13561 (N_13561,N_13449,N_13143);
nor U13562 (N_13562,N_13453,N_13146);
or U13563 (N_13563,N_13306,N_13221);
nor U13564 (N_13564,N_13188,N_13179);
xnor U13565 (N_13565,N_13316,N_13162);
xor U13566 (N_13566,N_13082,N_13062);
or U13567 (N_13567,N_13101,N_13385);
or U13568 (N_13568,N_13459,N_13186);
nand U13569 (N_13569,N_13400,N_13461);
or U13570 (N_13570,N_13283,N_13275);
nor U13571 (N_13571,N_13413,N_13269);
and U13572 (N_13572,N_13064,N_13038);
nor U13573 (N_13573,N_13399,N_13396);
nand U13574 (N_13574,N_13141,N_13033);
and U13575 (N_13575,N_13475,N_13378);
xor U13576 (N_13576,N_13420,N_13134);
nor U13577 (N_13577,N_13180,N_13318);
xnor U13578 (N_13578,N_13457,N_13020);
nor U13579 (N_13579,N_13035,N_13326);
nand U13580 (N_13580,N_13416,N_13229);
nand U13581 (N_13581,N_13174,N_13065);
or U13582 (N_13582,N_13091,N_13224);
nor U13583 (N_13583,N_13451,N_13328);
nand U13584 (N_13584,N_13234,N_13198);
xnor U13585 (N_13585,N_13372,N_13440);
and U13586 (N_13586,N_13125,N_13467);
nand U13587 (N_13587,N_13482,N_13383);
nand U13588 (N_13588,N_13070,N_13358);
and U13589 (N_13589,N_13362,N_13214);
nor U13590 (N_13590,N_13235,N_13246);
nand U13591 (N_13591,N_13052,N_13126);
and U13592 (N_13592,N_13137,N_13128);
nor U13593 (N_13593,N_13259,N_13435);
and U13594 (N_13594,N_13333,N_13034);
nand U13595 (N_13595,N_13054,N_13161);
nand U13596 (N_13596,N_13103,N_13171);
or U13597 (N_13597,N_13406,N_13123);
and U13598 (N_13598,N_13048,N_13249);
or U13599 (N_13599,N_13366,N_13345);
xor U13600 (N_13600,N_13220,N_13032);
and U13601 (N_13601,N_13488,N_13481);
nand U13602 (N_13602,N_13338,N_13072);
or U13603 (N_13603,N_13412,N_13006);
nand U13604 (N_13604,N_13276,N_13114);
nor U13605 (N_13605,N_13492,N_13191);
or U13606 (N_13606,N_13121,N_13487);
or U13607 (N_13607,N_13122,N_13115);
xor U13608 (N_13608,N_13434,N_13225);
and U13609 (N_13609,N_13042,N_13215);
xnor U13610 (N_13610,N_13363,N_13212);
nand U13611 (N_13611,N_13469,N_13106);
or U13612 (N_13612,N_13014,N_13160);
nor U13613 (N_13613,N_13013,N_13098);
and U13614 (N_13614,N_13069,N_13330);
nand U13615 (N_13615,N_13017,N_13087);
nand U13616 (N_13616,N_13102,N_13175);
nand U13617 (N_13617,N_13418,N_13293);
nand U13618 (N_13618,N_13142,N_13007);
nor U13619 (N_13619,N_13057,N_13022);
xor U13620 (N_13620,N_13077,N_13029);
nand U13621 (N_13621,N_13382,N_13041);
and U13622 (N_13622,N_13206,N_13315);
nand U13623 (N_13623,N_13166,N_13473);
nand U13624 (N_13624,N_13292,N_13248);
nor U13625 (N_13625,N_13371,N_13132);
or U13626 (N_13626,N_13063,N_13302);
nand U13627 (N_13627,N_13441,N_13216);
nor U13628 (N_13628,N_13131,N_13055);
nor U13629 (N_13629,N_13425,N_13468);
nand U13630 (N_13630,N_13213,N_13404);
nor U13631 (N_13631,N_13231,N_13243);
or U13632 (N_13632,N_13197,N_13455);
nor U13633 (N_13633,N_13168,N_13445);
and U13634 (N_13634,N_13192,N_13262);
and U13635 (N_13635,N_13484,N_13442);
nor U13636 (N_13636,N_13182,N_13270);
nand U13637 (N_13637,N_13119,N_13265);
nor U13638 (N_13638,N_13238,N_13204);
or U13639 (N_13639,N_13295,N_13046);
and U13640 (N_13640,N_13411,N_13000);
nand U13641 (N_13641,N_13341,N_13257);
nor U13642 (N_13642,N_13005,N_13422);
or U13643 (N_13643,N_13443,N_13397);
nor U13644 (N_13644,N_13335,N_13018);
nor U13645 (N_13645,N_13419,N_13104);
and U13646 (N_13646,N_13164,N_13107);
and U13647 (N_13647,N_13044,N_13219);
or U13648 (N_13648,N_13068,N_13253);
or U13649 (N_13649,N_13298,N_13080);
and U13650 (N_13650,N_13112,N_13489);
nor U13651 (N_13651,N_13045,N_13150);
xor U13652 (N_13652,N_13120,N_13281);
nand U13653 (N_13653,N_13423,N_13163);
and U13654 (N_13654,N_13199,N_13391);
and U13655 (N_13655,N_13002,N_13353);
nand U13656 (N_13656,N_13332,N_13244);
nand U13657 (N_13657,N_13239,N_13223);
nand U13658 (N_13658,N_13177,N_13154);
or U13659 (N_13659,N_13284,N_13178);
nor U13660 (N_13660,N_13233,N_13458);
and U13661 (N_13661,N_13109,N_13195);
or U13662 (N_13662,N_13351,N_13093);
nand U13663 (N_13663,N_13497,N_13226);
nor U13664 (N_13664,N_13384,N_13355);
nor U13665 (N_13665,N_13390,N_13454);
and U13666 (N_13666,N_13060,N_13227);
or U13667 (N_13667,N_13217,N_13252);
xnor U13668 (N_13668,N_13036,N_13153);
and U13669 (N_13669,N_13379,N_13311);
or U13670 (N_13670,N_13169,N_13491);
or U13671 (N_13671,N_13321,N_13376);
nand U13672 (N_13672,N_13256,N_13236);
nand U13673 (N_13673,N_13085,N_13393);
nand U13674 (N_13674,N_13019,N_13360);
nor U13675 (N_13675,N_13200,N_13050);
and U13676 (N_13676,N_13499,N_13324);
nor U13677 (N_13677,N_13172,N_13049);
nor U13678 (N_13678,N_13067,N_13099);
nand U13679 (N_13679,N_13480,N_13308);
nand U13680 (N_13680,N_13151,N_13407);
and U13681 (N_13681,N_13023,N_13304);
nor U13682 (N_13682,N_13157,N_13314);
or U13683 (N_13683,N_13405,N_13196);
nor U13684 (N_13684,N_13300,N_13317);
and U13685 (N_13685,N_13352,N_13375);
or U13686 (N_13686,N_13015,N_13139);
nand U13687 (N_13687,N_13127,N_13310);
or U13688 (N_13688,N_13053,N_13075);
and U13689 (N_13689,N_13322,N_13144);
xnor U13690 (N_13690,N_13031,N_13346);
or U13691 (N_13691,N_13415,N_13076);
or U13692 (N_13692,N_13016,N_13350);
nor U13693 (N_13693,N_13028,N_13218);
xor U13694 (N_13694,N_13156,N_13078);
or U13695 (N_13695,N_13245,N_13320);
or U13696 (N_13696,N_13279,N_13263);
nand U13697 (N_13697,N_13183,N_13210);
nor U13698 (N_13698,N_13030,N_13432);
nor U13699 (N_13699,N_13271,N_13026);
or U13700 (N_13700,N_13430,N_13367);
nand U13701 (N_13701,N_13264,N_13474);
nand U13702 (N_13702,N_13083,N_13261);
nor U13703 (N_13703,N_13348,N_13349);
nand U13704 (N_13704,N_13149,N_13092);
nand U13705 (N_13705,N_13222,N_13059);
and U13706 (N_13706,N_13273,N_13111);
and U13707 (N_13707,N_13130,N_13086);
xnor U13708 (N_13708,N_13374,N_13116);
xor U13709 (N_13709,N_13368,N_13277);
and U13710 (N_13710,N_13170,N_13117);
and U13711 (N_13711,N_13274,N_13377);
nand U13712 (N_13712,N_13237,N_13402);
or U13713 (N_13713,N_13010,N_13135);
and U13714 (N_13714,N_13003,N_13452);
nand U13715 (N_13715,N_13299,N_13438);
nor U13716 (N_13716,N_13181,N_13303);
nor U13717 (N_13717,N_13339,N_13051);
and U13718 (N_13718,N_13327,N_13389);
nand U13719 (N_13719,N_13140,N_13370);
nand U13720 (N_13720,N_13056,N_13387);
nor U13721 (N_13721,N_13071,N_13401);
nand U13722 (N_13722,N_13286,N_13147);
and U13723 (N_13723,N_13208,N_13460);
nor U13724 (N_13724,N_13336,N_13498);
or U13725 (N_13725,N_13331,N_13448);
nand U13726 (N_13726,N_13108,N_13340);
or U13727 (N_13727,N_13027,N_13095);
and U13728 (N_13728,N_13187,N_13008);
nand U13729 (N_13729,N_13287,N_13118);
and U13730 (N_13730,N_13129,N_13047);
nor U13731 (N_13731,N_13167,N_13152);
nor U13732 (N_13732,N_13189,N_13291);
nand U13733 (N_13733,N_13319,N_13267);
xor U13734 (N_13734,N_13110,N_13356);
and U13735 (N_13735,N_13471,N_13228);
nand U13736 (N_13736,N_13138,N_13465);
or U13737 (N_13737,N_13232,N_13173);
or U13738 (N_13738,N_13040,N_13424);
and U13739 (N_13739,N_13211,N_13043);
nor U13740 (N_13740,N_13025,N_13478);
or U13741 (N_13741,N_13058,N_13301);
or U13742 (N_13742,N_13260,N_13094);
nand U13743 (N_13743,N_13464,N_13124);
nor U13744 (N_13744,N_13381,N_13329);
nand U13745 (N_13745,N_13193,N_13373);
nand U13746 (N_13746,N_13133,N_13342);
nand U13747 (N_13747,N_13113,N_13307);
nand U13748 (N_13748,N_13421,N_13205);
nor U13749 (N_13749,N_13297,N_13447);
and U13750 (N_13750,N_13044,N_13324);
or U13751 (N_13751,N_13159,N_13346);
or U13752 (N_13752,N_13172,N_13198);
and U13753 (N_13753,N_13096,N_13220);
xor U13754 (N_13754,N_13002,N_13383);
nor U13755 (N_13755,N_13241,N_13232);
and U13756 (N_13756,N_13414,N_13053);
xnor U13757 (N_13757,N_13490,N_13349);
or U13758 (N_13758,N_13275,N_13101);
nor U13759 (N_13759,N_13363,N_13147);
nand U13760 (N_13760,N_13214,N_13361);
or U13761 (N_13761,N_13184,N_13253);
nand U13762 (N_13762,N_13228,N_13243);
nand U13763 (N_13763,N_13397,N_13377);
xnor U13764 (N_13764,N_13332,N_13376);
nor U13765 (N_13765,N_13054,N_13261);
xor U13766 (N_13766,N_13106,N_13450);
nand U13767 (N_13767,N_13233,N_13312);
or U13768 (N_13768,N_13163,N_13424);
and U13769 (N_13769,N_13265,N_13455);
nand U13770 (N_13770,N_13023,N_13285);
nand U13771 (N_13771,N_13259,N_13477);
or U13772 (N_13772,N_13247,N_13300);
nand U13773 (N_13773,N_13052,N_13446);
xnor U13774 (N_13774,N_13337,N_13475);
nand U13775 (N_13775,N_13481,N_13188);
nand U13776 (N_13776,N_13090,N_13299);
and U13777 (N_13777,N_13407,N_13264);
nor U13778 (N_13778,N_13384,N_13153);
nand U13779 (N_13779,N_13333,N_13212);
nand U13780 (N_13780,N_13285,N_13101);
or U13781 (N_13781,N_13293,N_13181);
and U13782 (N_13782,N_13251,N_13464);
nor U13783 (N_13783,N_13050,N_13380);
and U13784 (N_13784,N_13460,N_13305);
nand U13785 (N_13785,N_13303,N_13260);
nand U13786 (N_13786,N_13435,N_13112);
nand U13787 (N_13787,N_13013,N_13242);
and U13788 (N_13788,N_13281,N_13196);
xor U13789 (N_13789,N_13276,N_13146);
and U13790 (N_13790,N_13274,N_13082);
nand U13791 (N_13791,N_13344,N_13292);
or U13792 (N_13792,N_13338,N_13153);
or U13793 (N_13793,N_13225,N_13082);
nor U13794 (N_13794,N_13026,N_13180);
xor U13795 (N_13795,N_13308,N_13326);
nand U13796 (N_13796,N_13292,N_13159);
and U13797 (N_13797,N_13071,N_13456);
or U13798 (N_13798,N_13158,N_13028);
or U13799 (N_13799,N_13134,N_13382);
nand U13800 (N_13800,N_13342,N_13420);
nor U13801 (N_13801,N_13283,N_13292);
and U13802 (N_13802,N_13057,N_13124);
and U13803 (N_13803,N_13457,N_13333);
nor U13804 (N_13804,N_13329,N_13051);
nor U13805 (N_13805,N_13143,N_13276);
xnor U13806 (N_13806,N_13027,N_13400);
and U13807 (N_13807,N_13124,N_13117);
nand U13808 (N_13808,N_13458,N_13093);
nand U13809 (N_13809,N_13467,N_13188);
or U13810 (N_13810,N_13315,N_13036);
nand U13811 (N_13811,N_13105,N_13194);
nor U13812 (N_13812,N_13185,N_13414);
and U13813 (N_13813,N_13385,N_13058);
xor U13814 (N_13814,N_13119,N_13271);
or U13815 (N_13815,N_13277,N_13464);
or U13816 (N_13816,N_13035,N_13212);
and U13817 (N_13817,N_13386,N_13418);
nor U13818 (N_13818,N_13071,N_13442);
nand U13819 (N_13819,N_13140,N_13285);
xor U13820 (N_13820,N_13176,N_13493);
xor U13821 (N_13821,N_13047,N_13251);
and U13822 (N_13822,N_13194,N_13122);
and U13823 (N_13823,N_13340,N_13096);
nor U13824 (N_13824,N_13269,N_13307);
and U13825 (N_13825,N_13309,N_13106);
or U13826 (N_13826,N_13357,N_13337);
nand U13827 (N_13827,N_13429,N_13035);
nand U13828 (N_13828,N_13486,N_13104);
or U13829 (N_13829,N_13241,N_13394);
nand U13830 (N_13830,N_13293,N_13459);
nor U13831 (N_13831,N_13415,N_13464);
and U13832 (N_13832,N_13032,N_13394);
nor U13833 (N_13833,N_13396,N_13132);
or U13834 (N_13834,N_13357,N_13481);
nor U13835 (N_13835,N_13114,N_13399);
and U13836 (N_13836,N_13052,N_13363);
nand U13837 (N_13837,N_13382,N_13006);
nor U13838 (N_13838,N_13000,N_13194);
nor U13839 (N_13839,N_13283,N_13231);
or U13840 (N_13840,N_13028,N_13256);
or U13841 (N_13841,N_13443,N_13148);
or U13842 (N_13842,N_13127,N_13137);
and U13843 (N_13843,N_13064,N_13332);
and U13844 (N_13844,N_13495,N_13338);
nand U13845 (N_13845,N_13318,N_13481);
or U13846 (N_13846,N_13230,N_13097);
or U13847 (N_13847,N_13294,N_13491);
nor U13848 (N_13848,N_13274,N_13329);
xnor U13849 (N_13849,N_13356,N_13350);
nand U13850 (N_13850,N_13430,N_13390);
nor U13851 (N_13851,N_13131,N_13012);
nand U13852 (N_13852,N_13119,N_13167);
and U13853 (N_13853,N_13418,N_13321);
nor U13854 (N_13854,N_13004,N_13001);
xnor U13855 (N_13855,N_13231,N_13469);
or U13856 (N_13856,N_13466,N_13456);
or U13857 (N_13857,N_13025,N_13290);
xor U13858 (N_13858,N_13192,N_13152);
xnor U13859 (N_13859,N_13421,N_13136);
or U13860 (N_13860,N_13438,N_13478);
and U13861 (N_13861,N_13480,N_13155);
nor U13862 (N_13862,N_13357,N_13151);
nand U13863 (N_13863,N_13046,N_13004);
nand U13864 (N_13864,N_13004,N_13232);
nand U13865 (N_13865,N_13352,N_13403);
or U13866 (N_13866,N_13331,N_13371);
and U13867 (N_13867,N_13108,N_13205);
and U13868 (N_13868,N_13098,N_13073);
nor U13869 (N_13869,N_13429,N_13056);
nor U13870 (N_13870,N_13236,N_13138);
nand U13871 (N_13871,N_13034,N_13236);
nand U13872 (N_13872,N_13159,N_13261);
and U13873 (N_13873,N_13331,N_13345);
nand U13874 (N_13874,N_13138,N_13361);
or U13875 (N_13875,N_13400,N_13454);
and U13876 (N_13876,N_13364,N_13316);
nand U13877 (N_13877,N_13091,N_13115);
and U13878 (N_13878,N_13024,N_13334);
xnor U13879 (N_13879,N_13269,N_13120);
nor U13880 (N_13880,N_13367,N_13136);
nand U13881 (N_13881,N_13024,N_13443);
or U13882 (N_13882,N_13263,N_13283);
nand U13883 (N_13883,N_13491,N_13336);
nor U13884 (N_13884,N_13447,N_13126);
nand U13885 (N_13885,N_13422,N_13176);
or U13886 (N_13886,N_13266,N_13252);
nand U13887 (N_13887,N_13090,N_13258);
nor U13888 (N_13888,N_13199,N_13450);
nand U13889 (N_13889,N_13292,N_13486);
nor U13890 (N_13890,N_13478,N_13430);
xnor U13891 (N_13891,N_13182,N_13002);
xor U13892 (N_13892,N_13364,N_13390);
or U13893 (N_13893,N_13134,N_13457);
or U13894 (N_13894,N_13055,N_13091);
and U13895 (N_13895,N_13246,N_13251);
xnor U13896 (N_13896,N_13313,N_13140);
or U13897 (N_13897,N_13193,N_13080);
or U13898 (N_13898,N_13167,N_13316);
nor U13899 (N_13899,N_13084,N_13272);
nand U13900 (N_13900,N_13488,N_13353);
nor U13901 (N_13901,N_13297,N_13046);
and U13902 (N_13902,N_13147,N_13008);
and U13903 (N_13903,N_13364,N_13226);
nor U13904 (N_13904,N_13207,N_13273);
nor U13905 (N_13905,N_13248,N_13451);
and U13906 (N_13906,N_13190,N_13362);
nor U13907 (N_13907,N_13462,N_13222);
or U13908 (N_13908,N_13001,N_13117);
or U13909 (N_13909,N_13414,N_13298);
nor U13910 (N_13910,N_13221,N_13330);
or U13911 (N_13911,N_13277,N_13420);
and U13912 (N_13912,N_13412,N_13257);
nor U13913 (N_13913,N_13351,N_13182);
or U13914 (N_13914,N_13346,N_13392);
nand U13915 (N_13915,N_13396,N_13049);
or U13916 (N_13916,N_13276,N_13126);
nor U13917 (N_13917,N_13141,N_13248);
or U13918 (N_13918,N_13055,N_13481);
or U13919 (N_13919,N_13061,N_13253);
nor U13920 (N_13920,N_13422,N_13171);
xnor U13921 (N_13921,N_13156,N_13063);
nand U13922 (N_13922,N_13037,N_13138);
and U13923 (N_13923,N_13398,N_13232);
nand U13924 (N_13924,N_13106,N_13163);
or U13925 (N_13925,N_13312,N_13111);
and U13926 (N_13926,N_13042,N_13057);
nor U13927 (N_13927,N_13401,N_13352);
and U13928 (N_13928,N_13423,N_13402);
and U13929 (N_13929,N_13425,N_13487);
and U13930 (N_13930,N_13325,N_13424);
nor U13931 (N_13931,N_13097,N_13334);
or U13932 (N_13932,N_13424,N_13042);
nor U13933 (N_13933,N_13029,N_13087);
nor U13934 (N_13934,N_13060,N_13044);
nand U13935 (N_13935,N_13053,N_13164);
xor U13936 (N_13936,N_13024,N_13480);
nor U13937 (N_13937,N_13279,N_13320);
and U13938 (N_13938,N_13189,N_13127);
nand U13939 (N_13939,N_13277,N_13347);
and U13940 (N_13940,N_13367,N_13211);
nand U13941 (N_13941,N_13177,N_13012);
nand U13942 (N_13942,N_13095,N_13182);
nand U13943 (N_13943,N_13483,N_13190);
and U13944 (N_13944,N_13291,N_13483);
xor U13945 (N_13945,N_13197,N_13068);
nor U13946 (N_13946,N_13328,N_13240);
and U13947 (N_13947,N_13211,N_13466);
nand U13948 (N_13948,N_13376,N_13020);
and U13949 (N_13949,N_13067,N_13482);
and U13950 (N_13950,N_13021,N_13012);
xor U13951 (N_13951,N_13324,N_13459);
nor U13952 (N_13952,N_13433,N_13242);
nor U13953 (N_13953,N_13187,N_13250);
nand U13954 (N_13954,N_13286,N_13158);
nand U13955 (N_13955,N_13439,N_13128);
nand U13956 (N_13956,N_13144,N_13050);
nand U13957 (N_13957,N_13211,N_13426);
and U13958 (N_13958,N_13031,N_13271);
xnor U13959 (N_13959,N_13480,N_13464);
xor U13960 (N_13960,N_13041,N_13429);
xnor U13961 (N_13961,N_13186,N_13146);
nand U13962 (N_13962,N_13351,N_13071);
and U13963 (N_13963,N_13023,N_13480);
and U13964 (N_13964,N_13007,N_13094);
and U13965 (N_13965,N_13283,N_13173);
nor U13966 (N_13966,N_13123,N_13274);
or U13967 (N_13967,N_13454,N_13327);
and U13968 (N_13968,N_13089,N_13095);
nor U13969 (N_13969,N_13060,N_13461);
or U13970 (N_13970,N_13473,N_13062);
and U13971 (N_13971,N_13441,N_13327);
nor U13972 (N_13972,N_13188,N_13173);
and U13973 (N_13973,N_13458,N_13339);
xor U13974 (N_13974,N_13315,N_13120);
or U13975 (N_13975,N_13314,N_13287);
or U13976 (N_13976,N_13089,N_13181);
or U13977 (N_13977,N_13401,N_13141);
nand U13978 (N_13978,N_13199,N_13216);
and U13979 (N_13979,N_13199,N_13294);
nor U13980 (N_13980,N_13417,N_13108);
nor U13981 (N_13981,N_13312,N_13157);
nand U13982 (N_13982,N_13268,N_13019);
xor U13983 (N_13983,N_13182,N_13146);
xor U13984 (N_13984,N_13250,N_13481);
nand U13985 (N_13985,N_13216,N_13159);
and U13986 (N_13986,N_13309,N_13052);
and U13987 (N_13987,N_13059,N_13203);
or U13988 (N_13988,N_13125,N_13359);
and U13989 (N_13989,N_13171,N_13457);
or U13990 (N_13990,N_13387,N_13196);
and U13991 (N_13991,N_13313,N_13028);
and U13992 (N_13992,N_13137,N_13085);
and U13993 (N_13993,N_13092,N_13357);
and U13994 (N_13994,N_13364,N_13413);
nand U13995 (N_13995,N_13334,N_13200);
nand U13996 (N_13996,N_13302,N_13379);
xnor U13997 (N_13997,N_13325,N_13480);
or U13998 (N_13998,N_13059,N_13204);
xor U13999 (N_13999,N_13336,N_13413);
nor U14000 (N_14000,N_13773,N_13629);
and U14001 (N_14001,N_13618,N_13876);
nor U14002 (N_14002,N_13502,N_13774);
and U14003 (N_14003,N_13881,N_13596);
xor U14004 (N_14004,N_13752,N_13790);
nand U14005 (N_14005,N_13849,N_13525);
and U14006 (N_14006,N_13980,N_13813);
or U14007 (N_14007,N_13555,N_13778);
or U14008 (N_14008,N_13583,N_13702);
xnor U14009 (N_14009,N_13852,N_13714);
nand U14010 (N_14010,N_13511,N_13522);
nor U14011 (N_14011,N_13788,N_13937);
and U14012 (N_14012,N_13893,N_13894);
and U14013 (N_14013,N_13756,N_13757);
or U14014 (N_14014,N_13973,N_13754);
and U14015 (N_14015,N_13805,N_13635);
or U14016 (N_14016,N_13895,N_13738);
xnor U14017 (N_14017,N_13559,N_13612);
nand U14018 (N_14018,N_13520,N_13642);
or U14019 (N_14019,N_13573,N_13939);
and U14020 (N_14020,N_13554,N_13724);
xnor U14021 (N_14021,N_13709,N_13720);
and U14022 (N_14022,N_13861,N_13965);
or U14023 (N_14023,N_13747,N_13935);
nand U14024 (N_14024,N_13515,N_13510);
nor U14025 (N_14025,N_13808,N_13683);
xnor U14026 (N_14026,N_13868,N_13769);
nand U14027 (N_14027,N_13964,N_13557);
or U14028 (N_14028,N_13674,N_13797);
nand U14029 (N_14029,N_13732,N_13562);
or U14030 (N_14030,N_13907,N_13827);
or U14031 (N_14031,N_13750,N_13706);
nand U14032 (N_14032,N_13666,N_13838);
and U14033 (N_14033,N_13902,N_13616);
nand U14034 (N_14034,N_13904,N_13682);
or U14035 (N_14035,N_13631,N_13696);
nand U14036 (N_14036,N_13829,N_13984);
nor U14037 (N_14037,N_13842,N_13770);
or U14038 (N_14038,N_13816,N_13719);
nand U14039 (N_14039,N_13560,N_13906);
xnor U14040 (N_14040,N_13780,N_13912);
and U14041 (N_14041,N_13675,N_13978);
nand U14042 (N_14042,N_13529,N_13872);
nand U14043 (N_14043,N_13803,N_13593);
and U14044 (N_14044,N_13843,N_13531);
and U14045 (N_14045,N_13755,N_13552);
nor U14046 (N_14046,N_13609,N_13691);
and U14047 (N_14047,N_13587,N_13979);
nand U14048 (N_14048,N_13753,N_13987);
nand U14049 (N_14049,N_13646,N_13685);
xnor U14050 (N_14050,N_13841,N_13763);
and U14051 (N_14051,N_13801,N_13657);
nor U14052 (N_14052,N_13862,N_13995);
or U14053 (N_14053,N_13684,N_13925);
nand U14054 (N_14054,N_13637,N_13940);
or U14055 (N_14055,N_13891,N_13837);
or U14056 (N_14056,N_13850,N_13716);
and U14057 (N_14057,N_13595,N_13951);
and U14058 (N_14058,N_13848,N_13544);
and U14059 (N_14059,N_13762,N_13539);
xnor U14060 (N_14060,N_13857,N_13699);
xor U14061 (N_14061,N_13556,N_13955);
or U14062 (N_14062,N_13880,N_13653);
nor U14063 (N_14063,N_13545,N_13630);
and U14064 (N_14064,N_13795,N_13644);
nor U14065 (N_14065,N_13865,N_13695);
and U14066 (N_14066,N_13929,N_13972);
xor U14067 (N_14067,N_13603,N_13892);
and U14068 (N_14068,N_13991,N_13664);
nor U14069 (N_14069,N_13711,N_13647);
or U14070 (N_14070,N_13659,N_13812);
or U14071 (N_14071,N_13731,N_13878);
nor U14072 (N_14072,N_13650,N_13598);
nand U14073 (N_14073,N_13981,N_13758);
or U14074 (N_14074,N_13864,N_13707);
or U14075 (N_14075,N_13798,N_13896);
nor U14076 (N_14076,N_13854,N_13915);
nand U14077 (N_14077,N_13638,N_13996);
nand U14078 (N_14078,N_13819,N_13890);
and U14079 (N_14079,N_13582,N_13748);
or U14080 (N_14080,N_13820,N_13810);
and U14081 (N_14081,N_13985,N_13503);
or U14082 (N_14082,N_13500,N_13986);
nor U14083 (N_14083,N_13610,N_13941);
and U14084 (N_14084,N_13645,N_13920);
or U14085 (N_14085,N_13883,N_13811);
and U14086 (N_14086,N_13949,N_13513);
nand U14087 (N_14087,N_13866,N_13831);
nor U14088 (N_14088,N_13938,N_13698);
nor U14089 (N_14089,N_13768,N_13885);
nand U14090 (N_14090,N_13739,N_13922);
nor U14091 (N_14091,N_13879,N_13835);
and U14092 (N_14092,N_13708,N_13670);
or U14093 (N_14093,N_13814,N_13537);
or U14094 (N_14094,N_13615,N_13967);
xor U14095 (N_14095,N_13626,N_13656);
or U14096 (N_14096,N_13688,N_13608);
nor U14097 (N_14097,N_13668,N_13833);
xor U14098 (N_14098,N_13992,N_13578);
nor U14099 (N_14099,N_13746,N_13860);
xnor U14100 (N_14100,N_13651,N_13575);
and U14101 (N_14101,N_13663,N_13667);
and U14102 (N_14102,N_13526,N_13577);
and U14103 (N_14103,N_13634,N_13782);
and U14104 (N_14104,N_13519,N_13607);
nand U14105 (N_14105,N_13749,N_13953);
or U14106 (N_14106,N_13553,N_13936);
nand U14107 (N_14107,N_13565,N_13740);
or U14108 (N_14108,N_13543,N_13793);
nand U14109 (N_14109,N_13734,N_13649);
or U14110 (N_14110,N_13926,N_13844);
or U14111 (N_14111,N_13789,N_13518);
or U14112 (N_14112,N_13761,N_13957);
and U14113 (N_14113,N_13558,N_13530);
and U14114 (N_14114,N_13825,N_13648);
nand U14115 (N_14115,N_13680,N_13867);
or U14116 (N_14116,N_13767,N_13580);
or U14117 (N_14117,N_13772,N_13786);
nor U14118 (N_14118,N_13942,N_13889);
nor U14119 (N_14119,N_13822,N_13845);
nand U14120 (N_14120,N_13660,N_13606);
nand U14121 (N_14121,N_13538,N_13821);
or U14122 (N_14122,N_13723,N_13547);
or U14123 (N_14123,N_13705,N_13976);
xnor U14124 (N_14124,N_13771,N_13540);
nand U14125 (N_14125,N_13585,N_13913);
and U14126 (N_14126,N_13548,N_13946);
or U14127 (N_14127,N_13990,N_13592);
or U14128 (N_14128,N_13870,N_13527);
nor U14129 (N_14129,N_13673,N_13561);
or U14130 (N_14130,N_13588,N_13799);
and U14131 (N_14131,N_13584,N_13514);
and U14132 (N_14132,N_13916,N_13509);
and U14133 (N_14133,N_13931,N_13806);
nor U14134 (N_14134,N_13785,N_13903);
nand U14135 (N_14135,N_13692,N_13943);
nand U14136 (N_14136,N_13818,N_13963);
and U14137 (N_14137,N_13690,N_13662);
and U14138 (N_14138,N_13546,N_13625);
nor U14139 (N_14139,N_13781,N_13947);
nand U14140 (N_14140,N_13742,N_13549);
and U14141 (N_14141,N_13735,N_13859);
nand U14142 (N_14142,N_13617,N_13970);
and U14143 (N_14143,N_13794,N_13960);
or U14144 (N_14144,N_13921,N_13505);
or U14145 (N_14145,N_13988,N_13792);
nor U14146 (N_14146,N_13877,N_13760);
or U14147 (N_14147,N_13777,N_13779);
nor U14148 (N_14148,N_13570,N_13873);
and U14149 (N_14149,N_13542,N_13874);
or U14150 (N_14150,N_13727,N_13804);
nor U14151 (N_14151,N_13506,N_13851);
nand U14152 (N_14152,N_13574,N_13600);
nor U14153 (N_14153,N_13982,N_13636);
nand U14154 (N_14154,N_13908,N_13744);
nor U14155 (N_14155,N_13839,N_13669);
nand U14156 (N_14156,N_13997,N_13655);
nand U14157 (N_14157,N_13932,N_13620);
or U14158 (N_14158,N_13954,N_13977);
and U14159 (N_14159,N_13501,N_13589);
nor U14160 (N_14160,N_13886,N_13897);
nand U14161 (N_14161,N_13639,N_13817);
and U14162 (N_14162,N_13604,N_13787);
or U14163 (N_14163,N_13571,N_13776);
or U14164 (N_14164,N_13581,N_13905);
nand U14165 (N_14165,N_13567,N_13534);
nand U14166 (N_14166,N_13871,N_13622);
or U14167 (N_14167,N_13627,N_13783);
or U14168 (N_14168,N_13703,N_13952);
or U14169 (N_14169,N_13633,N_13933);
or U14170 (N_14170,N_13909,N_13676);
and U14171 (N_14171,N_13875,N_13983);
and U14172 (N_14172,N_13614,N_13602);
and U14173 (N_14173,N_13678,N_13899);
and U14174 (N_14174,N_13715,N_13579);
nor U14175 (N_14175,N_13658,N_13728);
xnor U14176 (N_14176,N_13802,N_13784);
nor U14177 (N_14177,N_13536,N_13846);
or U14178 (N_14178,N_13971,N_13621);
nand U14179 (N_14179,N_13733,N_13856);
or U14180 (N_14180,N_13564,N_13517);
or U14181 (N_14181,N_13911,N_13928);
nor U14182 (N_14182,N_13751,N_13632);
or U14183 (N_14183,N_13853,N_13800);
or U14184 (N_14184,N_13605,N_13945);
or U14185 (N_14185,N_13550,N_13640);
nor U14186 (N_14186,N_13969,N_13791);
nand U14187 (N_14187,N_13665,N_13576);
nand U14188 (N_14188,N_13958,N_13591);
nor U14189 (N_14189,N_13834,N_13759);
and U14190 (N_14190,N_13590,N_13807);
and U14191 (N_14191,N_13741,N_13677);
or U14192 (N_14192,N_13840,N_13766);
nor U14193 (N_14193,N_13898,N_13775);
or U14194 (N_14194,N_13882,N_13701);
or U14195 (N_14195,N_13624,N_13764);
or U14196 (N_14196,N_13950,N_13924);
nor U14197 (N_14197,N_13729,N_13586);
nor U14198 (N_14198,N_13523,N_13796);
and U14199 (N_14199,N_13989,N_13974);
nor U14200 (N_14200,N_13919,N_13689);
and U14201 (N_14201,N_13830,N_13563);
nand U14202 (N_14202,N_13568,N_13994);
and U14203 (N_14203,N_13726,N_13934);
nor U14204 (N_14204,N_13836,N_13858);
and U14205 (N_14205,N_13679,N_13697);
or U14206 (N_14206,N_13504,N_13694);
and U14207 (N_14207,N_13999,N_13736);
xnor U14208 (N_14208,N_13661,N_13672);
or U14209 (N_14209,N_13532,N_13521);
nor U14210 (N_14210,N_13566,N_13823);
nor U14211 (N_14211,N_13809,N_13681);
nand U14212 (N_14212,N_13968,N_13737);
or U14213 (N_14213,N_13671,N_13717);
or U14214 (N_14214,N_13594,N_13826);
xnor U14215 (N_14215,N_13725,N_13914);
xnor U14216 (N_14216,N_13869,N_13628);
nand U14217 (N_14217,N_13745,N_13551);
nand U14218 (N_14218,N_13572,N_13828);
xnor U14219 (N_14219,N_13944,N_13765);
or U14220 (N_14220,N_13722,N_13930);
nor U14221 (N_14221,N_13961,N_13535);
nand U14222 (N_14222,N_13619,N_13884);
nand U14223 (N_14223,N_13693,N_13652);
and U14224 (N_14224,N_13641,N_13569);
and U14225 (N_14225,N_13832,N_13863);
xor U14226 (N_14226,N_13993,N_13541);
nand U14227 (N_14227,N_13713,N_13601);
nor U14228 (N_14228,N_13918,N_13512);
and U14229 (N_14229,N_13887,N_13948);
nand U14230 (N_14230,N_13998,N_13730);
or U14231 (N_14231,N_13597,N_13824);
or U14232 (N_14232,N_13528,N_13712);
or U14233 (N_14233,N_13611,N_13966);
xnor U14234 (N_14234,N_13900,N_13743);
and U14235 (N_14235,N_13815,N_13718);
and U14236 (N_14236,N_13888,N_13686);
nor U14237 (N_14237,N_13917,N_13956);
or U14238 (N_14238,N_13927,N_13599);
or U14239 (N_14239,N_13923,N_13710);
and U14240 (N_14240,N_13508,N_13700);
and U14241 (N_14241,N_13687,N_13855);
and U14242 (N_14242,N_13910,N_13721);
or U14243 (N_14243,N_13613,N_13533);
or U14244 (N_14244,N_13524,N_13654);
and U14245 (N_14245,N_13507,N_13623);
nand U14246 (N_14246,N_13643,N_13962);
nor U14247 (N_14247,N_13704,N_13847);
nand U14248 (N_14248,N_13901,N_13975);
and U14249 (N_14249,N_13959,N_13516);
nor U14250 (N_14250,N_13676,N_13887);
or U14251 (N_14251,N_13903,N_13977);
nor U14252 (N_14252,N_13542,N_13907);
or U14253 (N_14253,N_13757,N_13511);
xor U14254 (N_14254,N_13607,N_13639);
nor U14255 (N_14255,N_13621,N_13653);
and U14256 (N_14256,N_13680,N_13825);
or U14257 (N_14257,N_13612,N_13767);
and U14258 (N_14258,N_13952,N_13814);
or U14259 (N_14259,N_13905,N_13815);
or U14260 (N_14260,N_13948,N_13992);
and U14261 (N_14261,N_13580,N_13656);
nand U14262 (N_14262,N_13570,N_13809);
nand U14263 (N_14263,N_13871,N_13509);
and U14264 (N_14264,N_13886,N_13874);
or U14265 (N_14265,N_13649,N_13648);
or U14266 (N_14266,N_13856,N_13500);
nor U14267 (N_14267,N_13928,N_13852);
nand U14268 (N_14268,N_13756,N_13997);
nor U14269 (N_14269,N_13595,N_13673);
nor U14270 (N_14270,N_13581,N_13544);
or U14271 (N_14271,N_13941,N_13755);
nand U14272 (N_14272,N_13749,N_13805);
and U14273 (N_14273,N_13631,N_13534);
or U14274 (N_14274,N_13560,N_13919);
or U14275 (N_14275,N_13721,N_13525);
nor U14276 (N_14276,N_13848,N_13802);
nand U14277 (N_14277,N_13786,N_13780);
or U14278 (N_14278,N_13871,N_13630);
nor U14279 (N_14279,N_13966,N_13918);
and U14280 (N_14280,N_13909,N_13913);
nor U14281 (N_14281,N_13762,N_13742);
nor U14282 (N_14282,N_13802,N_13842);
nand U14283 (N_14283,N_13552,N_13867);
or U14284 (N_14284,N_13874,N_13719);
nand U14285 (N_14285,N_13726,N_13825);
or U14286 (N_14286,N_13531,N_13737);
and U14287 (N_14287,N_13503,N_13812);
nand U14288 (N_14288,N_13867,N_13996);
and U14289 (N_14289,N_13937,N_13759);
nor U14290 (N_14290,N_13591,N_13907);
nor U14291 (N_14291,N_13695,N_13885);
and U14292 (N_14292,N_13654,N_13836);
and U14293 (N_14293,N_13881,N_13829);
nand U14294 (N_14294,N_13931,N_13969);
or U14295 (N_14295,N_13784,N_13660);
nor U14296 (N_14296,N_13666,N_13703);
xnor U14297 (N_14297,N_13599,N_13565);
nor U14298 (N_14298,N_13957,N_13512);
and U14299 (N_14299,N_13716,N_13664);
and U14300 (N_14300,N_13512,N_13551);
xnor U14301 (N_14301,N_13901,N_13939);
nand U14302 (N_14302,N_13528,N_13665);
nand U14303 (N_14303,N_13833,N_13670);
nor U14304 (N_14304,N_13755,N_13954);
or U14305 (N_14305,N_13969,N_13771);
and U14306 (N_14306,N_13501,N_13643);
xor U14307 (N_14307,N_13916,N_13822);
or U14308 (N_14308,N_13662,N_13718);
and U14309 (N_14309,N_13588,N_13933);
nand U14310 (N_14310,N_13909,N_13891);
and U14311 (N_14311,N_13616,N_13976);
nand U14312 (N_14312,N_13940,N_13799);
nor U14313 (N_14313,N_13515,N_13652);
xor U14314 (N_14314,N_13817,N_13702);
xor U14315 (N_14315,N_13944,N_13851);
or U14316 (N_14316,N_13678,N_13851);
nand U14317 (N_14317,N_13535,N_13706);
or U14318 (N_14318,N_13713,N_13842);
and U14319 (N_14319,N_13536,N_13900);
xnor U14320 (N_14320,N_13873,N_13663);
nand U14321 (N_14321,N_13833,N_13581);
nand U14322 (N_14322,N_13767,N_13933);
nor U14323 (N_14323,N_13749,N_13849);
nand U14324 (N_14324,N_13525,N_13939);
xor U14325 (N_14325,N_13809,N_13687);
nand U14326 (N_14326,N_13697,N_13919);
and U14327 (N_14327,N_13544,N_13961);
nor U14328 (N_14328,N_13745,N_13810);
nand U14329 (N_14329,N_13889,N_13757);
and U14330 (N_14330,N_13572,N_13909);
xor U14331 (N_14331,N_13700,N_13926);
or U14332 (N_14332,N_13966,N_13736);
nor U14333 (N_14333,N_13641,N_13805);
nand U14334 (N_14334,N_13670,N_13965);
or U14335 (N_14335,N_13744,N_13550);
nor U14336 (N_14336,N_13553,N_13972);
nor U14337 (N_14337,N_13611,N_13672);
xnor U14338 (N_14338,N_13842,N_13926);
nand U14339 (N_14339,N_13797,N_13504);
nand U14340 (N_14340,N_13718,N_13881);
nor U14341 (N_14341,N_13951,N_13870);
nor U14342 (N_14342,N_13661,N_13866);
xnor U14343 (N_14343,N_13852,N_13518);
xor U14344 (N_14344,N_13828,N_13993);
xor U14345 (N_14345,N_13602,N_13660);
and U14346 (N_14346,N_13934,N_13709);
and U14347 (N_14347,N_13539,N_13773);
or U14348 (N_14348,N_13696,N_13594);
and U14349 (N_14349,N_13973,N_13960);
nand U14350 (N_14350,N_13941,N_13580);
xor U14351 (N_14351,N_13760,N_13863);
nand U14352 (N_14352,N_13740,N_13949);
nand U14353 (N_14353,N_13732,N_13997);
xnor U14354 (N_14354,N_13885,N_13769);
xnor U14355 (N_14355,N_13594,N_13576);
xnor U14356 (N_14356,N_13724,N_13601);
nand U14357 (N_14357,N_13718,N_13666);
or U14358 (N_14358,N_13632,N_13982);
or U14359 (N_14359,N_13931,N_13692);
xnor U14360 (N_14360,N_13571,N_13690);
nor U14361 (N_14361,N_13907,N_13647);
or U14362 (N_14362,N_13838,N_13669);
or U14363 (N_14363,N_13720,N_13591);
nor U14364 (N_14364,N_13661,N_13503);
nor U14365 (N_14365,N_13957,N_13758);
and U14366 (N_14366,N_13736,N_13711);
or U14367 (N_14367,N_13748,N_13928);
nand U14368 (N_14368,N_13761,N_13703);
and U14369 (N_14369,N_13547,N_13585);
xnor U14370 (N_14370,N_13956,N_13739);
or U14371 (N_14371,N_13780,N_13583);
nand U14372 (N_14372,N_13605,N_13798);
nor U14373 (N_14373,N_13779,N_13825);
nor U14374 (N_14374,N_13845,N_13919);
or U14375 (N_14375,N_13611,N_13749);
or U14376 (N_14376,N_13921,N_13881);
nor U14377 (N_14377,N_13580,N_13573);
nand U14378 (N_14378,N_13668,N_13658);
nor U14379 (N_14379,N_13913,N_13603);
or U14380 (N_14380,N_13912,N_13528);
nor U14381 (N_14381,N_13551,N_13755);
and U14382 (N_14382,N_13715,N_13889);
nor U14383 (N_14383,N_13779,N_13789);
nand U14384 (N_14384,N_13736,N_13570);
and U14385 (N_14385,N_13661,N_13541);
xnor U14386 (N_14386,N_13548,N_13783);
or U14387 (N_14387,N_13845,N_13936);
nor U14388 (N_14388,N_13604,N_13579);
or U14389 (N_14389,N_13829,N_13556);
nor U14390 (N_14390,N_13729,N_13909);
and U14391 (N_14391,N_13774,N_13823);
or U14392 (N_14392,N_13620,N_13761);
nor U14393 (N_14393,N_13667,N_13986);
or U14394 (N_14394,N_13940,N_13631);
xnor U14395 (N_14395,N_13592,N_13667);
xor U14396 (N_14396,N_13670,N_13770);
or U14397 (N_14397,N_13530,N_13926);
nand U14398 (N_14398,N_13917,N_13922);
nand U14399 (N_14399,N_13988,N_13772);
or U14400 (N_14400,N_13787,N_13830);
nor U14401 (N_14401,N_13540,N_13644);
nand U14402 (N_14402,N_13977,N_13533);
or U14403 (N_14403,N_13671,N_13989);
and U14404 (N_14404,N_13841,N_13630);
nor U14405 (N_14405,N_13755,N_13833);
or U14406 (N_14406,N_13999,N_13802);
nand U14407 (N_14407,N_13975,N_13718);
xnor U14408 (N_14408,N_13802,N_13940);
nor U14409 (N_14409,N_13758,N_13899);
or U14410 (N_14410,N_13567,N_13568);
nor U14411 (N_14411,N_13741,N_13833);
nand U14412 (N_14412,N_13630,N_13626);
nor U14413 (N_14413,N_13774,N_13916);
nand U14414 (N_14414,N_13954,N_13700);
and U14415 (N_14415,N_13975,N_13559);
and U14416 (N_14416,N_13948,N_13744);
nor U14417 (N_14417,N_13959,N_13884);
nor U14418 (N_14418,N_13814,N_13513);
nand U14419 (N_14419,N_13768,N_13569);
nand U14420 (N_14420,N_13585,N_13698);
or U14421 (N_14421,N_13512,N_13846);
and U14422 (N_14422,N_13649,N_13545);
and U14423 (N_14423,N_13551,N_13805);
nand U14424 (N_14424,N_13613,N_13989);
and U14425 (N_14425,N_13990,N_13521);
nor U14426 (N_14426,N_13587,N_13522);
nor U14427 (N_14427,N_13816,N_13822);
and U14428 (N_14428,N_13806,N_13964);
and U14429 (N_14429,N_13966,N_13923);
and U14430 (N_14430,N_13633,N_13926);
or U14431 (N_14431,N_13887,N_13783);
xor U14432 (N_14432,N_13733,N_13660);
xor U14433 (N_14433,N_13923,N_13519);
nor U14434 (N_14434,N_13687,N_13972);
or U14435 (N_14435,N_13706,N_13633);
xor U14436 (N_14436,N_13747,N_13898);
nand U14437 (N_14437,N_13569,N_13860);
nand U14438 (N_14438,N_13914,N_13882);
and U14439 (N_14439,N_13691,N_13719);
nor U14440 (N_14440,N_13643,N_13607);
or U14441 (N_14441,N_13644,N_13596);
and U14442 (N_14442,N_13750,N_13989);
or U14443 (N_14443,N_13759,N_13734);
nand U14444 (N_14444,N_13793,N_13598);
or U14445 (N_14445,N_13521,N_13887);
nor U14446 (N_14446,N_13813,N_13636);
and U14447 (N_14447,N_13533,N_13954);
nor U14448 (N_14448,N_13840,N_13843);
or U14449 (N_14449,N_13974,N_13867);
nor U14450 (N_14450,N_13958,N_13824);
xnor U14451 (N_14451,N_13708,N_13742);
or U14452 (N_14452,N_13642,N_13543);
nand U14453 (N_14453,N_13611,N_13788);
nand U14454 (N_14454,N_13535,N_13579);
or U14455 (N_14455,N_13622,N_13876);
and U14456 (N_14456,N_13833,N_13633);
and U14457 (N_14457,N_13549,N_13699);
or U14458 (N_14458,N_13612,N_13939);
xnor U14459 (N_14459,N_13532,N_13577);
nand U14460 (N_14460,N_13532,N_13548);
nand U14461 (N_14461,N_13897,N_13940);
nand U14462 (N_14462,N_13872,N_13869);
nand U14463 (N_14463,N_13942,N_13548);
nor U14464 (N_14464,N_13897,N_13585);
and U14465 (N_14465,N_13972,N_13847);
nand U14466 (N_14466,N_13518,N_13766);
or U14467 (N_14467,N_13529,N_13776);
and U14468 (N_14468,N_13979,N_13777);
and U14469 (N_14469,N_13982,N_13816);
and U14470 (N_14470,N_13601,N_13649);
nor U14471 (N_14471,N_13838,N_13830);
nor U14472 (N_14472,N_13721,N_13633);
xnor U14473 (N_14473,N_13993,N_13547);
nand U14474 (N_14474,N_13502,N_13611);
nor U14475 (N_14475,N_13756,N_13502);
nor U14476 (N_14476,N_13813,N_13654);
xnor U14477 (N_14477,N_13594,N_13870);
nor U14478 (N_14478,N_13822,N_13858);
or U14479 (N_14479,N_13908,N_13631);
nor U14480 (N_14480,N_13931,N_13825);
or U14481 (N_14481,N_13766,N_13758);
nor U14482 (N_14482,N_13726,N_13983);
or U14483 (N_14483,N_13838,N_13842);
and U14484 (N_14484,N_13941,N_13568);
or U14485 (N_14485,N_13841,N_13847);
or U14486 (N_14486,N_13914,N_13743);
nor U14487 (N_14487,N_13831,N_13892);
nand U14488 (N_14488,N_13970,N_13879);
nand U14489 (N_14489,N_13653,N_13964);
or U14490 (N_14490,N_13573,N_13814);
or U14491 (N_14491,N_13625,N_13756);
or U14492 (N_14492,N_13697,N_13777);
and U14493 (N_14493,N_13614,N_13652);
and U14494 (N_14494,N_13955,N_13957);
and U14495 (N_14495,N_13998,N_13517);
or U14496 (N_14496,N_13708,N_13892);
xnor U14497 (N_14497,N_13669,N_13758);
xor U14498 (N_14498,N_13993,N_13598);
and U14499 (N_14499,N_13675,N_13851);
and U14500 (N_14500,N_14207,N_14188);
nor U14501 (N_14501,N_14422,N_14144);
nor U14502 (N_14502,N_14299,N_14010);
nor U14503 (N_14503,N_14011,N_14113);
nor U14504 (N_14504,N_14298,N_14013);
nor U14505 (N_14505,N_14069,N_14140);
xnor U14506 (N_14506,N_14202,N_14258);
nand U14507 (N_14507,N_14018,N_14412);
nand U14508 (N_14508,N_14323,N_14187);
nor U14509 (N_14509,N_14428,N_14349);
or U14510 (N_14510,N_14189,N_14129);
or U14511 (N_14511,N_14200,N_14418);
and U14512 (N_14512,N_14364,N_14145);
and U14513 (N_14513,N_14467,N_14431);
nor U14514 (N_14514,N_14355,N_14173);
and U14515 (N_14515,N_14096,N_14139);
nor U14516 (N_14516,N_14109,N_14409);
and U14517 (N_14517,N_14333,N_14348);
nor U14518 (N_14518,N_14219,N_14047);
or U14519 (N_14519,N_14233,N_14192);
nor U14520 (N_14520,N_14407,N_14388);
xor U14521 (N_14521,N_14228,N_14122);
or U14522 (N_14522,N_14260,N_14120);
nand U14523 (N_14523,N_14420,N_14395);
and U14524 (N_14524,N_14161,N_14235);
nand U14525 (N_14525,N_14330,N_14148);
nand U14526 (N_14526,N_14170,N_14309);
xor U14527 (N_14527,N_14267,N_14004);
nor U14528 (N_14528,N_14157,N_14392);
or U14529 (N_14529,N_14034,N_14269);
nand U14530 (N_14530,N_14087,N_14117);
and U14531 (N_14531,N_14121,N_14015);
xnor U14532 (N_14532,N_14281,N_14459);
nor U14533 (N_14533,N_14376,N_14166);
and U14534 (N_14534,N_14190,N_14461);
nand U14535 (N_14535,N_14062,N_14284);
and U14536 (N_14536,N_14435,N_14186);
nor U14537 (N_14537,N_14012,N_14180);
nand U14538 (N_14538,N_14375,N_14068);
nand U14539 (N_14539,N_14093,N_14220);
or U14540 (N_14540,N_14071,N_14421);
or U14541 (N_14541,N_14266,N_14221);
xnor U14542 (N_14542,N_14019,N_14239);
and U14543 (N_14543,N_14240,N_14227);
or U14544 (N_14544,N_14027,N_14091);
nand U14545 (N_14545,N_14119,N_14110);
or U14546 (N_14546,N_14048,N_14063);
and U14547 (N_14547,N_14084,N_14445);
and U14548 (N_14548,N_14072,N_14454);
or U14549 (N_14549,N_14021,N_14230);
xnor U14550 (N_14550,N_14497,N_14413);
and U14551 (N_14551,N_14114,N_14329);
or U14552 (N_14552,N_14095,N_14059);
or U14553 (N_14553,N_14070,N_14378);
nand U14554 (N_14554,N_14316,N_14433);
and U14555 (N_14555,N_14404,N_14311);
nor U14556 (N_14556,N_14265,N_14271);
nand U14557 (N_14557,N_14137,N_14244);
nand U14558 (N_14558,N_14101,N_14029);
nor U14559 (N_14559,N_14451,N_14124);
nor U14560 (N_14560,N_14367,N_14424);
nand U14561 (N_14561,N_14369,N_14492);
or U14562 (N_14562,N_14256,N_14468);
nand U14563 (N_14563,N_14389,N_14469);
xnor U14564 (N_14564,N_14051,N_14257);
or U14565 (N_14565,N_14306,N_14074);
and U14566 (N_14566,N_14305,N_14464);
nand U14567 (N_14567,N_14481,N_14423);
nor U14568 (N_14568,N_14127,N_14462);
or U14569 (N_14569,N_14406,N_14112);
or U14570 (N_14570,N_14372,N_14055);
and U14571 (N_14571,N_14210,N_14253);
nor U14572 (N_14572,N_14303,N_14480);
nor U14573 (N_14573,N_14336,N_14106);
and U14574 (N_14574,N_14094,N_14044);
nand U14575 (N_14575,N_14479,N_14438);
or U14576 (N_14576,N_14211,N_14171);
nor U14577 (N_14577,N_14191,N_14273);
nand U14578 (N_14578,N_14030,N_14380);
nor U14579 (N_14579,N_14359,N_14485);
and U14580 (N_14580,N_14272,N_14098);
and U14581 (N_14581,N_14088,N_14143);
nor U14582 (N_14582,N_14429,N_14415);
and U14583 (N_14583,N_14146,N_14009);
or U14584 (N_14584,N_14286,N_14224);
and U14585 (N_14585,N_14308,N_14078);
nor U14586 (N_14586,N_14089,N_14496);
nand U14587 (N_14587,N_14107,N_14079);
or U14588 (N_14588,N_14172,N_14357);
or U14589 (N_14589,N_14000,N_14159);
and U14590 (N_14590,N_14342,N_14338);
nor U14591 (N_14591,N_14463,N_14123);
or U14592 (N_14592,N_14035,N_14322);
and U14593 (N_14593,N_14448,N_14394);
nand U14594 (N_14594,N_14458,N_14478);
xor U14595 (N_14595,N_14493,N_14393);
nand U14596 (N_14596,N_14195,N_14115);
nand U14597 (N_14597,N_14229,N_14152);
nor U14598 (N_14598,N_14215,N_14118);
nor U14599 (N_14599,N_14344,N_14066);
nor U14600 (N_14600,N_14208,N_14499);
nor U14601 (N_14601,N_14263,N_14136);
nor U14602 (N_14602,N_14169,N_14442);
xnor U14603 (N_14603,N_14248,N_14405);
or U14604 (N_14604,N_14432,N_14446);
or U14605 (N_14605,N_14167,N_14193);
nor U14606 (N_14606,N_14196,N_14434);
nor U14607 (N_14607,N_14197,N_14108);
xor U14608 (N_14608,N_14486,N_14377);
and U14609 (N_14609,N_14276,N_14222);
or U14610 (N_14610,N_14043,N_14384);
or U14611 (N_14611,N_14053,N_14391);
nand U14612 (N_14612,N_14155,N_14259);
or U14613 (N_14613,N_14437,N_14312);
or U14614 (N_14614,N_14040,N_14440);
xor U14615 (N_14615,N_14090,N_14282);
nor U14616 (N_14616,N_14007,N_14283);
nand U14617 (N_14617,N_14397,N_14277);
nand U14618 (N_14618,N_14076,N_14280);
or U14619 (N_14619,N_14472,N_14238);
xnor U14620 (N_14620,N_14016,N_14425);
and U14621 (N_14621,N_14453,N_14199);
nor U14622 (N_14622,N_14484,N_14223);
or U14623 (N_14623,N_14226,N_14134);
and U14624 (N_14624,N_14476,N_14082);
and U14625 (N_14625,N_14252,N_14494);
nor U14626 (N_14626,N_14061,N_14275);
or U14627 (N_14627,N_14443,N_14141);
or U14628 (N_14628,N_14455,N_14296);
and U14629 (N_14629,N_14046,N_14174);
nor U14630 (N_14630,N_14331,N_14313);
nor U14631 (N_14631,N_14017,N_14241);
and U14632 (N_14632,N_14396,N_14345);
xnor U14633 (N_14633,N_14450,N_14184);
and U14634 (N_14634,N_14335,N_14125);
xor U14635 (N_14635,N_14178,N_14149);
xnor U14636 (N_14636,N_14270,N_14102);
and U14637 (N_14637,N_14288,N_14441);
nand U14638 (N_14638,N_14483,N_14398);
and U14639 (N_14639,N_14411,N_14201);
nor U14640 (N_14640,N_14278,N_14028);
or U14641 (N_14641,N_14430,N_14319);
and U14642 (N_14642,N_14362,N_14156);
nor U14643 (N_14643,N_14482,N_14142);
or U14644 (N_14644,N_14328,N_14067);
xnor U14645 (N_14645,N_14163,N_14491);
or U14646 (N_14646,N_14225,N_14206);
nand U14647 (N_14647,N_14456,N_14132);
xor U14648 (N_14648,N_14343,N_14042);
nor U14649 (N_14649,N_14150,N_14387);
or U14650 (N_14650,N_14116,N_14085);
nor U14651 (N_14651,N_14250,N_14358);
nor U14652 (N_14652,N_14470,N_14179);
nand U14653 (N_14653,N_14317,N_14341);
or U14654 (N_14654,N_14056,N_14340);
or U14655 (N_14655,N_14293,N_14318);
or U14656 (N_14656,N_14465,N_14365);
nor U14657 (N_14657,N_14151,N_14247);
and U14658 (N_14658,N_14386,N_14334);
or U14659 (N_14659,N_14006,N_14041);
nor U14660 (N_14660,N_14243,N_14060);
xor U14661 (N_14661,N_14473,N_14399);
and U14662 (N_14662,N_14022,N_14057);
and U14663 (N_14663,N_14488,N_14374);
nand U14664 (N_14664,N_14401,N_14005);
nand U14665 (N_14665,N_14050,N_14254);
and U14666 (N_14666,N_14326,N_14054);
or U14667 (N_14667,N_14321,N_14194);
and U14668 (N_14668,N_14287,N_14354);
and U14669 (N_14669,N_14039,N_14036);
nand U14670 (N_14670,N_14315,N_14176);
or U14671 (N_14671,N_14177,N_14198);
and U14672 (N_14672,N_14217,N_14255);
or U14673 (N_14673,N_14495,N_14371);
xnor U14674 (N_14674,N_14291,N_14024);
nand U14675 (N_14675,N_14213,N_14182);
nand U14676 (N_14676,N_14353,N_14410);
and U14677 (N_14677,N_14408,N_14379);
and U14678 (N_14678,N_14460,N_14310);
nand U14679 (N_14679,N_14475,N_14332);
and U14680 (N_14680,N_14083,N_14268);
and U14681 (N_14681,N_14154,N_14400);
nand U14682 (N_14682,N_14444,N_14447);
and U14683 (N_14683,N_14264,N_14097);
nor U14684 (N_14684,N_14302,N_14204);
or U14685 (N_14685,N_14175,N_14471);
or U14686 (N_14686,N_14290,N_14350);
nand U14687 (N_14687,N_14160,N_14324);
nand U14688 (N_14688,N_14297,N_14477);
and U14689 (N_14689,N_14352,N_14138);
nand U14690 (N_14690,N_14383,N_14162);
and U14691 (N_14691,N_14131,N_14232);
and U14692 (N_14692,N_14274,N_14285);
nor U14693 (N_14693,N_14237,N_14295);
nand U14694 (N_14694,N_14158,N_14236);
and U14695 (N_14695,N_14203,N_14064);
or U14696 (N_14696,N_14382,N_14249);
and U14697 (N_14697,N_14346,N_14474);
and U14698 (N_14698,N_14426,N_14075);
nor U14699 (N_14699,N_14073,N_14103);
and U14700 (N_14700,N_14307,N_14077);
and U14701 (N_14701,N_14147,N_14449);
and U14702 (N_14702,N_14363,N_14279);
nor U14703 (N_14703,N_14314,N_14081);
or U14704 (N_14704,N_14419,N_14320);
nor U14705 (N_14705,N_14360,N_14402);
or U14706 (N_14706,N_14304,N_14020);
nand U14707 (N_14707,N_14032,N_14168);
and U14708 (N_14708,N_14153,N_14218);
nor U14709 (N_14709,N_14023,N_14104);
xnor U14710 (N_14710,N_14417,N_14294);
nor U14711 (N_14711,N_14300,N_14452);
nand U14712 (N_14712,N_14361,N_14133);
and U14713 (N_14713,N_14457,N_14065);
nand U14714 (N_14714,N_14181,N_14038);
nand U14715 (N_14715,N_14356,N_14183);
or U14716 (N_14716,N_14058,N_14246);
nor U14717 (N_14717,N_14111,N_14289);
xor U14718 (N_14718,N_14001,N_14086);
and U14719 (N_14719,N_14185,N_14351);
nand U14720 (N_14720,N_14366,N_14014);
or U14721 (N_14721,N_14214,N_14080);
nor U14722 (N_14722,N_14008,N_14165);
nor U14723 (N_14723,N_14261,N_14099);
or U14724 (N_14724,N_14031,N_14498);
nand U14725 (N_14725,N_14026,N_14052);
xor U14726 (N_14726,N_14164,N_14414);
or U14727 (N_14727,N_14416,N_14381);
and U14728 (N_14728,N_14037,N_14209);
nand U14729 (N_14729,N_14049,N_14403);
nor U14730 (N_14730,N_14347,N_14135);
or U14731 (N_14731,N_14339,N_14436);
and U14732 (N_14732,N_14466,N_14262);
nor U14733 (N_14733,N_14245,N_14128);
nor U14734 (N_14734,N_14216,N_14301);
nor U14735 (N_14735,N_14292,N_14325);
nand U14736 (N_14736,N_14105,N_14234);
nand U14737 (N_14737,N_14130,N_14427);
nor U14738 (N_14738,N_14100,N_14002);
nor U14739 (N_14739,N_14487,N_14390);
xor U14740 (N_14740,N_14368,N_14025);
nor U14741 (N_14741,N_14385,N_14092);
and U14742 (N_14742,N_14490,N_14370);
nor U14743 (N_14743,N_14033,N_14439);
nor U14744 (N_14744,N_14489,N_14126);
xor U14745 (N_14745,N_14242,N_14337);
nand U14746 (N_14746,N_14212,N_14327);
and U14747 (N_14747,N_14251,N_14205);
and U14748 (N_14748,N_14373,N_14231);
or U14749 (N_14749,N_14003,N_14045);
or U14750 (N_14750,N_14206,N_14274);
and U14751 (N_14751,N_14165,N_14485);
nor U14752 (N_14752,N_14220,N_14384);
nand U14753 (N_14753,N_14467,N_14310);
nor U14754 (N_14754,N_14119,N_14115);
nand U14755 (N_14755,N_14376,N_14428);
nor U14756 (N_14756,N_14258,N_14458);
or U14757 (N_14757,N_14283,N_14474);
nand U14758 (N_14758,N_14280,N_14265);
and U14759 (N_14759,N_14120,N_14335);
nor U14760 (N_14760,N_14060,N_14071);
and U14761 (N_14761,N_14364,N_14187);
nor U14762 (N_14762,N_14025,N_14135);
and U14763 (N_14763,N_14462,N_14086);
nand U14764 (N_14764,N_14106,N_14153);
and U14765 (N_14765,N_14323,N_14071);
nand U14766 (N_14766,N_14057,N_14342);
and U14767 (N_14767,N_14193,N_14116);
and U14768 (N_14768,N_14331,N_14094);
or U14769 (N_14769,N_14375,N_14152);
or U14770 (N_14770,N_14043,N_14213);
nand U14771 (N_14771,N_14175,N_14451);
and U14772 (N_14772,N_14069,N_14258);
xor U14773 (N_14773,N_14473,N_14371);
nor U14774 (N_14774,N_14301,N_14061);
and U14775 (N_14775,N_14441,N_14093);
or U14776 (N_14776,N_14137,N_14117);
or U14777 (N_14777,N_14100,N_14365);
nand U14778 (N_14778,N_14471,N_14401);
or U14779 (N_14779,N_14408,N_14129);
nor U14780 (N_14780,N_14475,N_14015);
nor U14781 (N_14781,N_14233,N_14263);
xor U14782 (N_14782,N_14125,N_14085);
and U14783 (N_14783,N_14460,N_14498);
or U14784 (N_14784,N_14334,N_14398);
or U14785 (N_14785,N_14362,N_14373);
nor U14786 (N_14786,N_14322,N_14242);
nand U14787 (N_14787,N_14395,N_14224);
nor U14788 (N_14788,N_14270,N_14187);
nor U14789 (N_14789,N_14014,N_14323);
nand U14790 (N_14790,N_14254,N_14044);
and U14791 (N_14791,N_14014,N_14127);
or U14792 (N_14792,N_14282,N_14432);
and U14793 (N_14793,N_14014,N_14200);
nand U14794 (N_14794,N_14256,N_14343);
and U14795 (N_14795,N_14433,N_14289);
and U14796 (N_14796,N_14042,N_14346);
nand U14797 (N_14797,N_14254,N_14295);
nor U14798 (N_14798,N_14217,N_14207);
or U14799 (N_14799,N_14079,N_14318);
and U14800 (N_14800,N_14491,N_14126);
nand U14801 (N_14801,N_14277,N_14317);
nor U14802 (N_14802,N_14472,N_14094);
or U14803 (N_14803,N_14073,N_14336);
nor U14804 (N_14804,N_14134,N_14178);
nand U14805 (N_14805,N_14474,N_14384);
nand U14806 (N_14806,N_14068,N_14157);
or U14807 (N_14807,N_14182,N_14112);
nand U14808 (N_14808,N_14470,N_14335);
nand U14809 (N_14809,N_14158,N_14490);
nand U14810 (N_14810,N_14249,N_14068);
nand U14811 (N_14811,N_14152,N_14227);
or U14812 (N_14812,N_14192,N_14384);
nand U14813 (N_14813,N_14228,N_14076);
and U14814 (N_14814,N_14269,N_14138);
and U14815 (N_14815,N_14161,N_14366);
nand U14816 (N_14816,N_14427,N_14147);
xor U14817 (N_14817,N_14370,N_14499);
nor U14818 (N_14818,N_14073,N_14299);
or U14819 (N_14819,N_14070,N_14412);
or U14820 (N_14820,N_14280,N_14059);
nand U14821 (N_14821,N_14476,N_14244);
nand U14822 (N_14822,N_14259,N_14082);
nor U14823 (N_14823,N_14490,N_14121);
nand U14824 (N_14824,N_14183,N_14456);
or U14825 (N_14825,N_14251,N_14354);
or U14826 (N_14826,N_14393,N_14060);
or U14827 (N_14827,N_14303,N_14354);
or U14828 (N_14828,N_14468,N_14215);
or U14829 (N_14829,N_14017,N_14311);
or U14830 (N_14830,N_14449,N_14066);
or U14831 (N_14831,N_14171,N_14076);
or U14832 (N_14832,N_14387,N_14129);
and U14833 (N_14833,N_14338,N_14249);
nand U14834 (N_14834,N_14050,N_14064);
or U14835 (N_14835,N_14327,N_14388);
nand U14836 (N_14836,N_14111,N_14133);
nor U14837 (N_14837,N_14015,N_14239);
or U14838 (N_14838,N_14376,N_14318);
or U14839 (N_14839,N_14288,N_14497);
and U14840 (N_14840,N_14352,N_14465);
or U14841 (N_14841,N_14407,N_14253);
or U14842 (N_14842,N_14001,N_14267);
xnor U14843 (N_14843,N_14485,N_14232);
nor U14844 (N_14844,N_14328,N_14275);
and U14845 (N_14845,N_14331,N_14494);
nand U14846 (N_14846,N_14339,N_14131);
nand U14847 (N_14847,N_14186,N_14100);
and U14848 (N_14848,N_14144,N_14267);
and U14849 (N_14849,N_14348,N_14072);
xnor U14850 (N_14850,N_14140,N_14438);
or U14851 (N_14851,N_14052,N_14469);
and U14852 (N_14852,N_14419,N_14234);
or U14853 (N_14853,N_14414,N_14451);
and U14854 (N_14854,N_14130,N_14278);
or U14855 (N_14855,N_14390,N_14063);
or U14856 (N_14856,N_14442,N_14186);
or U14857 (N_14857,N_14347,N_14247);
nand U14858 (N_14858,N_14235,N_14049);
or U14859 (N_14859,N_14147,N_14245);
or U14860 (N_14860,N_14127,N_14451);
nor U14861 (N_14861,N_14461,N_14469);
nor U14862 (N_14862,N_14365,N_14110);
and U14863 (N_14863,N_14171,N_14087);
nand U14864 (N_14864,N_14352,N_14124);
or U14865 (N_14865,N_14419,N_14104);
and U14866 (N_14866,N_14298,N_14243);
nor U14867 (N_14867,N_14272,N_14493);
and U14868 (N_14868,N_14261,N_14104);
nand U14869 (N_14869,N_14074,N_14143);
nor U14870 (N_14870,N_14073,N_14061);
and U14871 (N_14871,N_14210,N_14343);
nor U14872 (N_14872,N_14164,N_14141);
nor U14873 (N_14873,N_14269,N_14293);
nand U14874 (N_14874,N_14211,N_14113);
or U14875 (N_14875,N_14297,N_14089);
nand U14876 (N_14876,N_14082,N_14177);
nor U14877 (N_14877,N_14084,N_14198);
nor U14878 (N_14878,N_14392,N_14012);
or U14879 (N_14879,N_14445,N_14351);
or U14880 (N_14880,N_14413,N_14174);
or U14881 (N_14881,N_14458,N_14250);
or U14882 (N_14882,N_14100,N_14183);
or U14883 (N_14883,N_14424,N_14080);
or U14884 (N_14884,N_14391,N_14211);
and U14885 (N_14885,N_14081,N_14096);
or U14886 (N_14886,N_14218,N_14339);
or U14887 (N_14887,N_14088,N_14291);
or U14888 (N_14888,N_14416,N_14107);
xor U14889 (N_14889,N_14254,N_14238);
and U14890 (N_14890,N_14005,N_14120);
nor U14891 (N_14891,N_14156,N_14180);
nor U14892 (N_14892,N_14481,N_14496);
xor U14893 (N_14893,N_14407,N_14495);
nand U14894 (N_14894,N_14295,N_14306);
or U14895 (N_14895,N_14327,N_14347);
and U14896 (N_14896,N_14003,N_14380);
nand U14897 (N_14897,N_14454,N_14151);
and U14898 (N_14898,N_14396,N_14430);
or U14899 (N_14899,N_14252,N_14085);
or U14900 (N_14900,N_14365,N_14442);
nand U14901 (N_14901,N_14234,N_14187);
nor U14902 (N_14902,N_14322,N_14464);
xor U14903 (N_14903,N_14495,N_14449);
and U14904 (N_14904,N_14363,N_14330);
nor U14905 (N_14905,N_14121,N_14444);
nor U14906 (N_14906,N_14057,N_14143);
or U14907 (N_14907,N_14110,N_14472);
or U14908 (N_14908,N_14096,N_14483);
and U14909 (N_14909,N_14473,N_14321);
xor U14910 (N_14910,N_14326,N_14482);
and U14911 (N_14911,N_14489,N_14399);
or U14912 (N_14912,N_14092,N_14020);
and U14913 (N_14913,N_14185,N_14085);
nand U14914 (N_14914,N_14496,N_14448);
nor U14915 (N_14915,N_14068,N_14084);
nand U14916 (N_14916,N_14275,N_14489);
xnor U14917 (N_14917,N_14483,N_14144);
or U14918 (N_14918,N_14390,N_14019);
nand U14919 (N_14919,N_14490,N_14464);
nor U14920 (N_14920,N_14039,N_14353);
and U14921 (N_14921,N_14006,N_14035);
or U14922 (N_14922,N_14266,N_14128);
or U14923 (N_14923,N_14052,N_14437);
nor U14924 (N_14924,N_14158,N_14042);
nor U14925 (N_14925,N_14170,N_14236);
or U14926 (N_14926,N_14354,N_14221);
nand U14927 (N_14927,N_14347,N_14156);
nand U14928 (N_14928,N_14153,N_14395);
or U14929 (N_14929,N_14497,N_14062);
nand U14930 (N_14930,N_14134,N_14413);
nand U14931 (N_14931,N_14162,N_14359);
nor U14932 (N_14932,N_14389,N_14072);
or U14933 (N_14933,N_14067,N_14038);
and U14934 (N_14934,N_14383,N_14240);
and U14935 (N_14935,N_14134,N_14020);
xor U14936 (N_14936,N_14054,N_14444);
xor U14937 (N_14937,N_14221,N_14488);
or U14938 (N_14938,N_14053,N_14302);
or U14939 (N_14939,N_14372,N_14232);
and U14940 (N_14940,N_14118,N_14301);
nand U14941 (N_14941,N_14347,N_14391);
xnor U14942 (N_14942,N_14059,N_14395);
or U14943 (N_14943,N_14429,N_14447);
nor U14944 (N_14944,N_14482,N_14261);
and U14945 (N_14945,N_14073,N_14085);
nor U14946 (N_14946,N_14092,N_14375);
or U14947 (N_14947,N_14242,N_14296);
nand U14948 (N_14948,N_14314,N_14357);
and U14949 (N_14949,N_14474,N_14417);
or U14950 (N_14950,N_14355,N_14177);
nor U14951 (N_14951,N_14284,N_14182);
nand U14952 (N_14952,N_14024,N_14089);
nor U14953 (N_14953,N_14279,N_14496);
or U14954 (N_14954,N_14462,N_14120);
xor U14955 (N_14955,N_14306,N_14000);
or U14956 (N_14956,N_14159,N_14414);
nand U14957 (N_14957,N_14482,N_14246);
nor U14958 (N_14958,N_14066,N_14119);
nor U14959 (N_14959,N_14167,N_14402);
nor U14960 (N_14960,N_14279,N_14461);
nor U14961 (N_14961,N_14487,N_14282);
nand U14962 (N_14962,N_14448,N_14268);
and U14963 (N_14963,N_14454,N_14128);
and U14964 (N_14964,N_14124,N_14037);
nor U14965 (N_14965,N_14425,N_14304);
nand U14966 (N_14966,N_14191,N_14421);
or U14967 (N_14967,N_14485,N_14402);
or U14968 (N_14968,N_14076,N_14182);
or U14969 (N_14969,N_14109,N_14015);
or U14970 (N_14970,N_14166,N_14310);
nand U14971 (N_14971,N_14437,N_14324);
nor U14972 (N_14972,N_14218,N_14360);
and U14973 (N_14973,N_14084,N_14057);
nand U14974 (N_14974,N_14492,N_14065);
nand U14975 (N_14975,N_14461,N_14150);
or U14976 (N_14976,N_14487,N_14114);
nor U14977 (N_14977,N_14438,N_14271);
nor U14978 (N_14978,N_14069,N_14475);
or U14979 (N_14979,N_14452,N_14010);
nor U14980 (N_14980,N_14271,N_14289);
nor U14981 (N_14981,N_14128,N_14244);
nand U14982 (N_14982,N_14389,N_14009);
nand U14983 (N_14983,N_14470,N_14419);
nand U14984 (N_14984,N_14266,N_14220);
nand U14985 (N_14985,N_14379,N_14154);
nand U14986 (N_14986,N_14332,N_14223);
nand U14987 (N_14987,N_14163,N_14251);
or U14988 (N_14988,N_14470,N_14365);
xor U14989 (N_14989,N_14483,N_14256);
or U14990 (N_14990,N_14149,N_14284);
xor U14991 (N_14991,N_14075,N_14002);
and U14992 (N_14992,N_14284,N_14420);
nor U14993 (N_14993,N_14271,N_14000);
or U14994 (N_14994,N_14318,N_14423);
nor U14995 (N_14995,N_14451,N_14248);
nor U14996 (N_14996,N_14186,N_14310);
nand U14997 (N_14997,N_14370,N_14328);
or U14998 (N_14998,N_14476,N_14053);
nand U14999 (N_14999,N_14286,N_14237);
and UO_0 (O_0,N_14892,N_14806);
nand UO_1 (O_1,N_14962,N_14740);
and UO_2 (O_2,N_14929,N_14605);
nor UO_3 (O_3,N_14956,N_14875);
nor UO_4 (O_4,N_14969,N_14646);
nand UO_5 (O_5,N_14935,N_14586);
nand UO_6 (O_6,N_14871,N_14502);
nor UO_7 (O_7,N_14803,N_14743);
and UO_8 (O_8,N_14512,N_14642);
and UO_9 (O_9,N_14587,N_14556);
or UO_10 (O_10,N_14667,N_14887);
or UO_11 (O_11,N_14976,N_14736);
and UO_12 (O_12,N_14786,N_14568);
or UO_13 (O_13,N_14934,N_14999);
nor UO_14 (O_14,N_14614,N_14672);
nor UO_15 (O_15,N_14623,N_14581);
xnor UO_16 (O_16,N_14860,N_14737);
and UO_17 (O_17,N_14645,N_14615);
and UO_18 (O_18,N_14560,N_14886);
or UO_19 (O_19,N_14735,N_14977);
xor UO_20 (O_20,N_14703,N_14948);
nor UO_21 (O_21,N_14894,N_14798);
or UO_22 (O_22,N_14524,N_14611);
or UO_23 (O_23,N_14988,N_14778);
or UO_24 (O_24,N_14538,N_14507);
nand UO_25 (O_25,N_14692,N_14807);
nor UO_26 (O_26,N_14613,N_14527);
nor UO_27 (O_27,N_14591,N_14801);
nand UO_28 (O_28,N_14846,N_14525);
and UO_29 (O_29,N_14983,N_14598);
nand UO_30 (O_30,N_14684,N_14693);
or UO_31 (O_31,N_14734,N_14984);
or UO_32 (O_32,N_14987,N_14731);
nor UO_33 (O_33,N_14589,N_14767);
nand UO_34 (O_34,N_14809,N_14669);
nor UO_35 (O_35,N_14972,N_14583);
nor UO_36 (O_36,N_14794,N_14617);
or UO_37 (O_37,N_14608,N_14550);
or UO_38 (O_38,N_14784,N_14922);
and UO_39 (O_39,N_14503,N_14749);
xor UO_40 (O_40,N_14545,N_14931);
and UO_41 (O_41,N_14744,N_14594);
or UO_42 (O_42,N_14822,N_14723);
nor UO_43 (O_43,N_14989,N_14867);
nand UO_44 (O_44,N_14680,N_14604);
nand UO_45 (O_45,N_14795,N_14772);
xnor UO_46 (O_46,N_14810,N_14578);
xor UO_47 (O_47,N_14952,N_14547);
nor UO_48 (O_48,N_14982,N_14917);
or UO_49 (O_49,N_14730,N_14838);
nor UO_50 (O_50,N_14673,N_14814);
or UO_51 (O_51,N_14657,N_14928);
xor UO_52 (O_52,N_14592,N_14575);
and UO_53 (O_53,N_14571,N_14825);
nor UO_54 (O_54,N_14804,N_14762);
nor UO_55 (O_55,N_14517,N_14963);
nor UO_56 (O_56,N_14821,N_14812);
nor UO_57 (O_57,N_14661,N_14607);
nand UO_58 (O_58,N_14510,N_14920);
xor UO_59 (O_59,N_14558,N_14848);
and UO_60 (O_60,N_14792,N_14742);
nand UO_61 (O_61,N_14501,N_14873);
nand UO_62 (O_62,N_14946,N_14654);
or UO_63 (O_63,N_14633,N_14802);
nand UO_64 (O_64,N_14898,N_14745);
xnor UO_65 (O_65,N_14842,N_14981);
and UO_66 (O_66,N_14752,N_14576);
or UO_67 (O_67,N_14785,N_14820);
nand UO_68 (O_68,N_14997,N_14844);
or UO_69 (O_69,N_14921,N_14939);
or UO_70 (O_70,N_14632,N_14549);
nand UO_71 (O_71,N_14964,N_14683);
or UO_72 (O_72,N_14843,N_14659);
nand UO_73 (O_73,N_14521,N_14970);
xor UO_74 (O_74,N_14783,N_14841);
nand UO_75 (O_75,N_14790,N_14933);
and UO_76 (O_76,N_14559,N_14874);
nand UO_77 (O_77,N_14828,N_14665);
or UO_78 (O_78,N_14528,N_14513);
nor UO_79 (O_79,N_14811,N_14546);
nand UO_80 (O_80,N_14823,N_14722);
or UO_81 (O_81,N_14631,N_14638);
xnor UO_82 (O_82,N_14707,N_14971);
or UO_83 (O_83,N_14725,N_14602);
and UO_84 (O_84,N_14818,N_14567);
xnor UO_85 (O_85,N_14849,N_14833);
nor UO_86 (O_86,N_14597,N_14663);
or UO_87 (O_87,N_14616,N_14699);
xor UO_88 (O_88,N_14865,N_14534);
nand UO_89 (O_89,N_14685,N_14978);
nor UO_90 (O_90,N_14993,N_14697);
and UO_91 (O_91,N_14950,N_14557);
nand UO_92 (O_92,N_14688,N_14765);
nor UO_93 (O_93,N_14881,N_14796);
xor UO_94 (O_94,N_14915,N_14777);
or UO_95 (O_95,N_14516,N_14764);
and UO_96 (O_96,N_14855,N_14896);
nor UO_97 (O_97,N_14815,N_14694);
and UO_98 (O_98,N_14913,N_14554);
or UO_99 (O_99,N_14577,N_14544);
and UO_100 (O_100,N_14960,N_14756);
or UO_101 (O_101,N_14585,N_14717);
nor UO_102 (O_102,N_14603,N_14755);
or UO_103 (O_103,N_14961,N_14548);
xor UO_104 (O_104,N_14936,N_14720);
nand UO_105 (O_105,N_14690,N_14640);
nor UO_106 (O_106,N_14641,N_14564);
nand UO_107 (O_107,N_14543,N_14509);
nand UO_108 (O_108,N_14941,N_14979);
nor UO_109 (O_109,N_14870,N_14957);
and UO_110 (O_110,N_14940,N_14670);
nand UO_111 (O_111,N_14951,N_14845);
xnor UO_112 (O_112,N_14751,N_14553);
or UO_113 (O_113,N_14835,N_14671);
nor UO_114 (O_114,N_14907,N_14588);
and UO_115 (O_115,N_14862,N_14565);
or UO_116 (O_116,N_14562,N_14747);
or UO_117 (O_117,N_14884,N_14893);
nor UO_118 (O_118,N_14572,N_14912);
and UO_119 (O_119,N_14705,N_14709);
nor UO_120 (O_120,N_14901,N_14868);
and UO_121 (O_121,N_14781,N_14861);
and UO_122 (O_122,N_14609,N_14911);
nand UO_123 (O_123,N_14805,N_14955);
nor UO_124 (O_124,N_14771,N_14797);
and UO_125 (O_125,N_14746,N_14696);
or UO_126 (O_126,N_14698,N_14610);
or UO_127 (O_127,N_14628,N_14537);
or UO_128 (O_128,N_14953,N_14830);
nand UO_129 (O_129,N_14926,N_14569);
and UO_130 (O_130,N_14885,N_14664);
and UO_131 (O_131,N_14829,N_14891);
nand UO_132 (O_132,N_14662,N_14918);
and UO_133 (O_133,N_14506,N_14593);
and UO_134 (O_134,N_14721,N_14775);
and UO_135 (O_135,N_14500,N_14773);
nand UO_136 (O_136,N_14980,N_14863);
xor UO_137 (O_137,N_14619,N_14760);
nand UO_138 (O_138,N_14600,N_14561);
or UO_139 (O_139,N_14649,N_14768);
xnor UO_140 (O_140,N_14769,N_14504);
or UO_141 (O_141,N_14776,N_14715);
or UO_142 (O_142,N_14656,N_14679);
or UO_143 (O_143,N_14530,N_14650);
and UO_144 (O_144,N_14759,N_14895);
nor UO_145 (O_145,N_14714,N_14878);
nand UO_146 (O_146,N_14973,N_14741);
or UO_147 (O_147,N_14655,N_14630);
nor UO_148 (O_148,N_14853,N_14748);
nor UO_149 (O_149,N_14858,N_14750);
or UO_150 (O_150,N_14648,N_14716);
or UO_151 (O_151,N_14508,N_14541);
nor UO_152 (O_152,N_14519,N_14925);
or UO_153 (O_153,N_14943,N_14582);
and UO_154 (O_154,N_14618,N_14724);
nor UO_155 (O_155,N_14859,N_14729);
and UO_156 (O_156,N_14555,N_14954);
nand UO_157 (O_157,N_14949,N_14854);
or UO_158 (O_158,N_14622,N_14727);
nand UO_159 (O_159,N_14579,N_14994);
xor UO_160 (O_160,N_14678,N_14791);
nand UO_161 (O_161,N_14540,N_14682);
and UO_162 (O_162,N_14832,N_14932);
or UO_163 (O_163,N_14601,N_14563);
nand UO_164 (O_164,N_14728,N_14856);
xor UO_165 (O_165,N_14816,N_14651);
nand UO_166 (O_166,N_14942,N_14847);
xor UO_167 (O_167,N_14706,N_14869);
and UO_168 (O_168,N_14904,N_14552);
xnor UO_169 (O_169,N_14701,N_14910);
xnor UO_170 (O_170,N_14647,N_14542);
nor UO_171 (O_171,N_14520,N_14888);
nand UO_172 (O_172,N_14627,N_14686);
or UO_173 (O_173,N_14840,N_14634);
nand UO_174 (O_174,N_14580,N_14660);
nor UO_175 (O_175,N_14839,N_14643);
xor UO_176 (O_176,N_14629,N_14890);
nor UO_177 (O_177,N_14924,N_14836);
and UO_178 (O_178,N_14674,N_14566);
or UO_179 (O_179,N_14695,N_14880);
or UO_180 (O_180,N_14908,N_14787);
nor UO_181 (O_181,N_14713,N_14626);
nor UO_182 (O_182,N_14808,N_14532);
and UO_183 (O_183,N_14711,N_14905);
or UO_184 (O_184,N_14570,N_14710);
nand UO_185 (O_185,N_14995,N_14526);
nor UO_186 (O_186,N_14906,N_14573);
nor UO_187 (O_187,N_14927,N_14621);
nor UO_188 (O_188,N_14857,N_14712);
or UO_189 (O_189,N_14719,N_14852);
or UO_190 (O_190,N_14531,N_14937);
nor UO_191 (O_191,N_14819,N_14947);
and UO_192 (O_192,N_14511,N_14788);
nand UO_193 (O_193,N_14899,N_14606);
and UO_194 (O_194,N_14687,N_14866);
nand UO_195 (O_195,N_14584,N_14533);
nor UO_196 (O_196,N_14799,N_14945);
and UO_197 (O_197,N_14919,N_14996);
nor UO_198 (O_198,N_14824,N_14831);
and UO_199 (O_199,N_14636,N_14872);
and UO_200 (O_200,N_14535,N_14635);
and UO_201 (O_201,N_14739,N_14770);
nor UO_202 (O_202,N_14691,N_14826);
and UO_203 (O_203,N_14738,N_14595);
xor UO_204 (O_204,N_14596,N_14914);
nor UO_205 (O_205,N_14668,N_14992);
or UO_206 (O_206,N_14681,N_14726);
nand UO_207 (O_207,N_14652,N_14529);
nand UO_208 (O_208,N_14864,N_14612);
nand UO_209 (O_209,N_14902,N_14704);
nor UO_210 (O_210,N_14967,N_14644);
or UO_211 (O_211,N_14985,N_14625);
and UO_212 (O_212,N_14718,N_14998);
xnor UO_213 (O_213,N_14518,N_14774);
xor UO_214 (O_214,N_14900,N_14817);
nor UO_215 (O_215,N_14761,N_14990);
and UO_216 (O_216,N_14758,N_14599);
nand UO_217 (O_217,N_14732,N_14879);
nand UO_218 (O_218,N_14624,N_14965);
or UO_219 (O_219,N_14974,N_14780);
nor UO_220 (O_220,N_14676,N_14837);
and UO_221 (O_221,N_14909,N_14733);
and UO_222 (O_222,N_14782,N_14515);
xor UO_223 (O_223,N_14708,N_14958);
and UO_224 (O_224,N_14700,N_14986);
nor UO_225 (O_225,N_14930,N_14551);
or UO_226 (O_226,N_14505,N_14658);
or UO_227 (O_227,N_14763,N_14675);
and UO_228 (O_228,N_14813,N_14923);
and UO_229 (O_229,N_14689,N_14959);
and UO_230 (O_230,N_14882,N_14834);
nand UO_231 (O_231,N_14702,N_14620);
xnor UO_232 (O_232,N_14938,N_14539);
nand UO_233 (O_233,N_14827,N_14889);
nor UO_234 (O_234,N_14850,N_14975);
or UO_235 (O_235,N_14800,N_14753);
or UO_236 (O_236,N_14522,N_14991);
or UO_237 (O_237,N_14916,N_14944);
xor UO_238 (O_238,N_14536,N_14789);
or UO_239 (O_239,N_14876,N_14883);
and UO_240 (O_240,N_14779,N_14766);
and UO_241 (O_241,N_14793,N_14757);
nand UO_242 (O_242,N_14754,N_14677);
and UO_243 (O_243,N_14968,N_14639);
and UO_244 (O_244,N_14637,N_14966);
nor UO_245 (O_245,N_14523,N_14903);
and UO_246 (O_246,N_14574,N_14653);
and UO_247 (O_247,N_14851,N_14897);
nor UO_248 (O_248,N_14666,N_14514);
nor UO_249 (O_249,N_14590,N_14877);
nand UO_250 (O_250,N_14825,N_14829);
or UO_251 (O_251,N_14615,N_14583);
and UO_252 (O_252,N_14756,N_14532);
or UO_253 (O_253,N_14950,N_14792);
nor UO_254 (O_254,N_14632,N_14890);
nor UO_255 (O_255,N_14549,N_14735);
nand UO_256 (O_256,N_14894,N_14532);
or UO_257 (O_257,N_14785,N_14722);
and UO_258 (O_258,N_14930,N_14700);
nor UO_259 (O_259,N_14905,N_14539);
nor UO_260 (O_260,N_14508,N_14972);
nand UO_261 (O_261,N_14777,N_14556);
and UO_262 (O_262,N_14991,N_14894);
nand UO_263 (O_263,N_14516,N_14819);
nand UO_264 (O_264,N_14756,N_14894);
nor UO_265 (O_265,N_14980,N_14810);
or UO_266 (O_266,N_14871,N_14742);
nor UO_267 (O_267,N_14625,N_14703);
or UO_268 (O_268,N_14663,N_14905);
nor UO_269 (O_269,N_14795,N_14915);
xnor UO_270 (O_270,N_14990,N_14661);
and UO_271 (O_271,N_14727,N_14788);
xnor UO_272 (O_272,N_14540,N_14910);
xor UO_273 (O_273,N_14536,N_14908);
nand UO_274 (O_274,N_14819,N_14872);
and UO_275 (O_275,N_14742,N_14866);
xnor UO_276 (O_276,N_14977,N_14921);
or UO_277 (O_277,N_14952,N_14732);
nor UO_278 (O_278,N_14844,N_14662);
and UO_279 (O_279,N_14902,N_14965);
xor UO_280 (O_280,N_14780,N_14612);
or UO_281 (O_281,N_14876,N_14604);
nand UO_282 (O_282,N_14726,N_14956);
nand UO_283 (O_283,N_14876,N_14846);
nand UO_284 (O_284,N_14535,N_14600);
and UO_285 (O_285,N_14893,N_14514);
nand UO_286 (O_286,N_14714,N_14901);
or UO_287 (O_287,N_14729,N_14931);
and UO_288 (O_288,N_14799,N_14769);
nand UO_289 (O_289,N_14858,N_14553);
nor UO_290 (O_290,N_14648,N_14564);
and UO_291 (O_291,N_14886,N_14753);
or UO_292 (O_292,N_14826,N_14610);
nor UO_293 (O_293,N_14906,N_14585);
or UO_294 (O_294,N_14984,N_14638);
nand UO_295 (O_295,N_14526,N_14908);
or UO_296 (O_296,N_14602,N_14972);
nor UO_297 (O_297,N_14833,N_14699);
and UO_298 (O_298,N_14810,N_14954);
or UO_299 (O_299,N_14777,N_14994);
nand UO_300 (O_300,N_14734,N_14920);
nand UO_301 (O_301,N_14857,N_14826);
nor UO_302 (O_302,N_14817,N_14512);
nand UO_303 (O_303,N_14571,N_14507);
nor UO_304 (O_304,N_14811,N_14531);
and UO_305 (O_305,N_14776,N_14938);
nand UO_306 (O_306,N_14818,N_14762);
or UO_307 (O_307,N_14852,N_14713);
and UO_308 (O_308,N_14747,N_14660);
nor UO_309 (O_309,N_14651,N_14642);
nand UO_310 (O_310,N_14864,N_14622);
xnor UO_311 (O_311,N_14736,N_14994);
xor UO_312 (O_312,N_14666,N_14782);
or UO_313 (O_313,N_14897,N_14761);
nor UO_314 (O_314,N_14768,N_14896);
or UO_315 (O_315,N_14788,N_14928);
or UO_316 (O_316,N_14742,N_14586);
or UO_317 (O_317,N_14640,N_14749);
nor UO_318 (O_318,N_14999,N_14875);
xnor UO_319 (O_319,N_14781,N_14904);
and UO_320 (O_320,N_14977,N_14826);
xnor UO_321 (O_321,N_14689,N_14875);
nor UO_322 (O_322,N_14856,N_14829);
nor UO_323 (O_323,N_14937,N_14665);
or UO_324 (O_324,N_14940,N_14961);
or UO_325 (O_325,N_14697,N_14646);
and UO_326 (O_326,N_14943,N_14652);
nor UO_327 (O_327,N_14804,N_14942);
xor UO_328 (O_328,N_14596,N_14793);
and UO_329 (O_329,N_14741,N_14771);
or UO_330 (O_330,N_14548,N_14578);
nand UO_331 (O_331,N_14667,N_14635);
nor UO_332 (O_332,N_14655,N_14707);
or UO_333 (O_333,N_14919,N_14947);
nor UO_334 (O_334,N_14954,N_14859);
or UO_335 (O_335,N_14799,N_14919);
or UO_336 (O_336,N_14951,N_14803);
xor UO_337 (O_337,N_14612,N_14932);
nand UO_338 (O_338,N_14966,N_14806);
nor UO_339 (O_339,N_14807,N_14769);
nor UO_340 (O_340,N_14978,N_14588);
or UO_341 (O_341,N_14824,N_14880);
nor UO_342 (O_342,N_14543,N_14553);
nor UO_343 (O_343,N_14762,N_14622);
and UO_344 (O_344,N_14977,N_14630);
xnor UO_345 (O_345,N_14592,N_14503);
or UO_346 (O_346,N_14671,N_14655);
xor UO_347 (O_347,N_14561,N_14908);
nor UO_348 (O_348,N_14948,N_14533);
and UO_349 (O_349,N_14950,N_14816);
and UO_350 (O_350,N_14881,N_14906);
xnor UO_351 (O_351,N_14826,N_14889);
nand UO_352 (O_352,N_14890,N_14762);
and UO_353 (O_353,N_14924,N_14921);
nand UO_354 (O_354,N_14949,N_14562);
and UO_355 (O_355,N_14801,N_14533);
or UO_356 (O_356,N_14550,N_14559);
or UO_357 (O_357,N_14729,N_14664);
nor UO_358 (O_358,N_14915,N_14762);
or UO_359 (O_359,N_14515,N_14613);
nand UO_360 (O_360,N_14796,N_14774);
xnor UO_361 (O_361,N_14785,N_14910);
nand UO_362 (O_362,N_14853,N_14866);
xnor UO_363 (O_363,N_14587,N_14768);
and UO_364 (O_364,N_14764,N_14695);
nor UO_365 (O_365,N_14625,N_14548);
nand UO_366 (O_366,N_14845,N_14886);
xnor UO_367 (O_367,N_14952,N_14924);
and UO_368 (O_368,N_14866,N_14737);
nor UO_369 (O_369,N_14968,N_14819);
or UO_370 (O_370,N_14522,N_14902);
and UO_371 (O_371,N_14775,N_14705);
and UO_372 (O_372,N_14683,N_14903);
nor UO_373 (O_373,N_14860,N_14524);
xnor UO_374 (O_374,N_14874,N_14926);
nor UO_375 (O_375,N_14820,N_14881);
nand UO_376 (O_376,N_14676,N_14641);
nand UO_377 (O_377,N_14934,N_14705);
nand UO_378 (O_378,N_14912,N_14840);
xor UO_379 (O_379,N_14764,N_14792);
nand UO_380 (O_380,N_14696,N_14649);
nor UO_381 (O_381,N_14909,N_14750);
and UO_382 (O_382,N_14559,N_14829);
or UO_383 (O_383,N_14691,N_14612);
nand UO_384 (O_384,N_14710,N_14705);
and UO_385 (O_385,N_14652,N_14679);
and UO_386 (O_386,N_14909,N_14893);
nand UO_387 (O_387,N_14733,N_14564);
nor UO_388 (O_388,N_14714,N_14506);
and UO_389 (O_389,N_14872,N_14765);
nor UO_390 (O_390,N_14877,N_14752);
or UO_391 (O_391,N_14811,N_14998);
and UO_392 (O_392,N_14758,N_14552);
nor UO_393 (O_393,N_14534,N_14853);
or UO_394 (O_394,N_14683,N_14658);
or UO_395 (O_395,N_14708,N_14598);
and UO_396 (O_396,N_14582,N_14687);
and UO_397 (O_397,N_14813,N_14895);
nand UO_398 (O_398,N_14904,N_14678);
nor UO_399 (O_399,N_14773,N_14514);
and UO_400 (O_400,N_14708,N_14562);
nor UO_401 (O_401,N_14587,N_14981);
nand UO_402 (O_402,N_14681,N_14678);
nor UO_403 (O_403,N_14653,N_14983);
nor UO_404 (O_404,N_14951,N_14549);
nor UO_405 (O_405,N_14817,N_14788);
nor UO_406 (O_406,N_14753,N_14501);
or UO_407 (O_407,N_14774,N_14847);
nand UO_408 (O_408,N_14672,N_14701);
nor UO_409 (O_409,N_14665,N_14575);
nor UO_410 (O_410,N_14589,N_14718);
or UO_411 (O_411,N_14898,N_14577);
nand UO_412 (O_412,N_14668,N_14985);
or UO_413 (O_413,N_14990,N_14587);
and UO_414 (O_414,N_14693,N_14893);
nor UO_415 (O_415,N_14987,N_14519);
and UO_416 (O_416,N_14832,N_14520);
and UO_417 (O_417,N_14711,N_14516);
nand UO_418 (O_418,N_14869,N_14656);
or UO_419 (O_419,N_14949,N_14896);
nor UO_420 (O_420,N_14590,N_14964);
nand UO_421 (O_421,N_14548,N_14723);
or UO_422 (O_422,N_14921,N_14538);
or UO_423 (O_423,N_14883,N_14502);
and UO_424 (O_424,N_14596,N_14750);
or UO_425 (O_425,N_14687,N_14573);
and UO_426 (O_426,N_14940,N_14720);
and UO_427 (O_427,N_14876,N_14845);
and UO_428 (O_428,N_14563,N_14645);
xnor UO_429 (O_429,N_14633,N_14768);
or UO_430 (O_430,N_14715,N_14734);
or UO_431 (O_431,N_14800,N_14618);
and UO_432 (O_432,N_14843,N_14722);
and UO_433 (O_433,N_14955,N_14678);
or UO_434 (O_434,N_14801,N_14670);
and UO_435 (O_435,N_14927,N_14856);
and UO_436 (O_436,N_14843,N_14881);
nor UO_437 (O_437,N_14804,N_14586);
nor UO_438 (O_438,N_14663,N_14866);
and UO_439 (O_439,N_14807,N_14980);
nor UO_440 (O_440,N_14617,N_14869);
and UO_441 (O_441,N_14653,N_14844);
and UO_442 (O_442,N_14710,N_14881);
and UO_443 (O_443,N_14743,N_14967);
nand UO_444 (O_444,N_14854,N_14996);
or UO_445 (O_445,N_14865,N_14709);
xor UO_446 (O_446,N_14797,N_14741);
xnor UO_447 (O_447,N_14517,N_14696);
nand UO_448 (O_448,N_14582,N_14897);
and UO_449 (O_449,N_14659,N_14645);
and UO_450 (O_450,N_14566,N_14809);
nand UO_451 (O_451,N_14893,N_14595);
xnor UO_452 (O_452,N_14964,N_14661);
or UO_453 (O_453,N_14949,N_14976);
or UO_454 (O_454,N_14661,N_14888);
xnor UO_455 (O_455,N_14640,N_14604);
nor UO_456 (O_456,N_14794,N_14944);
or UO_457 (O_457,N_14706,N_14961);
and UO_458 (O_458,N_14589,N_14991);
or UO_459 (O_459,N_14826,N_14983);
and UO_460 (O_460,N_14866,N_14580);
xnor UO_461 (O_461,N_14842,N_14504);
nand UO_462 (O_462,N_14795,N_14646);
xnor UO_463 (O_463,N_14766,N_14554);
nand UO_464 (O_464,N_14931,N_14556);
or UO_465 (O_465,N_14755,N_14840);
xnor UO_466 (O_466,N_14990,N_14575);
or UO_467 (O_467,N_14849,N_14937);
and UO_468 (O_468,N_14689,N_14590);
nand UO_469 (O_469,N_14738,N_14690);
and UO_470 (O_470,N_14951,N_14672);
nand UO_471 (O_471,N_14854,N_14897);
xnor UO_472 (O_472,N_14861,N_14995);
nor UO_473 (O_473,N_14604,N_14571);
or UO_474 (O_474,N_14703,N_14818);
nor UO_475 (O_475,N_14759,N_14552);
nor UO_476 (O_476,N_14986,N_14531);
or UO_477 (O_477,N_14631,N_14619);
nand UO_478 (O_478,N_14631,N_14780);
nand UO_479 (O_479,N_14966,N_14676);
nor UO_480 (O_480,N_14920,N_14924);
xor UO_481 (O_481,N_14742,N_14552);
nand UO_482 (O_482,N_14891,N_14539);
nor UO_483 (O_483,N_14778,N_14533);
nand UO_484 (O_484,N_14622,N_14707);
nand UO_485 (O_485,N_14866,N_14625);
or UO_486 (O_486,N_14745,N_14780);
and UO_487 (O_487,N_14711,N_14848);
nor UO_488 (O_488,N_14959,N_14930);
and UO_489 (O_489,N_14831,N_14602);
and UO_490 (O_490,N_14845,N_14628);
nor UO_491 (O_491,N_14612,N_14866);
nand UO_492 (O_492,N_14796,N_14600);
nand UO_493 (O_493,N_14716,N_14680);
or UO_494 (O_494,N_14785,N_14716);
and UO_495 (O_495,N_14551,N_14704);
or UO_496 (O_496,N_14881,N_14775);
or UO_497 (O_497,N_14505,N_14699);
and UO_498 (O_498,N_14766,N_14772);
or UO_499 (O_499,N_14781,N_14854);
nand UO_500 (O_500,N_14673,N_14906);
nor UO_501 (O_501,N_14544,N_14580);
nand UO_502 (O_502,N_14771,N_14673);
nand UO_503 (O_503,N_14668,N_14873);
nor UO_504 (O_504,N_14677,N_14532);
and UO_505 (O_505,N_14775,N_14523);
nor UO_506 (O_506,N_14716,N_14909);
nor UO_507 (O_507,N_14527,N_14949);
nor UO_508 (O_508,N_14744,N_14810);
nor UO_509 (O_509,N_14724,N_14762);
nor UO_510 (O_510,N_14873,N_14944);
and UO_511 (O_511,N_14555,N_14706);
nor UO_512 (O_512,N_14942,N_14953);
or UO_513 (O_513,N_14794,N_14815);
and UO_514 (O_514,N_14917,N_14909);
nand UO_515 (O_515,N_14634,N_14818);
or UO_516 (O_516,N_14680,N_14624);
or UO_517 (O_517,N_14623,N_14546);
and UO_518 (O_518,N_14533,N_14694);
nand UO_519 (O_519,N_14519,N_14888);
nor UO_520 (O_520,N_14625,N_14781);
and UO_521 (O_521,N_14614,N_14611);
and UO_522 (O_522,N_14640,N_14990);
xnor UO_523 (O_523,N_14742,N_14708);
nor UO_524 (O_524,N_14915,N_14972);
nor UO_525 (O_525,N_14620,N_14831);
nand UO_526 (O_526,N_14694,N_14918);
nand UO_527 (O_527,N_14853,N_14972);
nand UO_528 (O_528,N_14612,N_14555);
and UO_529 (O_529,N_14651,N_14939);
nand UO_530 (O_530,N_14534,N_14929);
xnor UO_531 (O_531,N_14688,N_14984);
or UO_532 (O_532,N_14637,N_14986);
or UO_533 (O_533,N_14954,N_14856);
and UO_534 (O_534,N_14729,N_14565);
nor UO_535 (O_535,N_14873,N_14649);
and UO_536 (O_536,N_14889,N_14987);
or UO_537 (O_537,N_14808,N_14668);
or UO_538 (O_538,N_14784,N_14800);
or UO_539 (O_539,N_14921,N_14853);
nand UO_540 (O_540,N_14733,N_14520);
or UO_541 (O_541,N_14943,N_14860);
or UO_542 (O_542,N_14595,N_14536);
or UO_543 (O_543,N_14509,N_14634);
nand UO_544 (O_544,N_14562,N_14543);
nor UO_545 (O_545,N_14833,N_14674);
xor UO_546 (O_546,N_14916,N_14553);
nor UO_547 (O_547,N_14592,N_14680);
nor UO_548 (O_548,N_14506,N_14824);
or UO_549 (O_549,N_14695,N_14719);
xnor UO_550 (O_550,N_14970,N_14777);
or UO_551 (O_551,N_14751,N_14554);
or UO_552 (O_552,N_14666,N_14992);
xnor UO_553 (O_553,N_14989,N_14711);
nand UO_554 (O_554,N_14568,N_14750);
or UO_555 (O_555,N_14501,N_14747);
nand UO_556 (O_556,N_14782,N_14972);
nand UO_557 (O_557,N_14991,N_14673);
and UO_558 (O_558,N_14638,N_14830);
xnor UO_559 (O_559,N_14616,N_14868);
or UO_560 (O_560,N_14511,N_14935);
or UO_561 (O_561,N_14680,N_14647);
nand UO_562 (O_562,N_14614,N_14581);
nand UO_563 (O_563,N_14984,N_14588);
nand UO_564 (O_564,N_14744,N_14896);
nand UO_565 (O_565,N_14628,N_14830);
nand UO_566 (O_566,N_14636,N_14789);
xnor UO_567 (O_567,N_14795,N_14530);
and UO_568 (O_568,N_14583,N_14913);
nand UO_569 (O_569,N_14766,N_14759);
nor UO_570 (O_570,N_14654,N_14848);
and UO_571 (O_571,N_14692,N_14771);
xor UO_572 (O_572,N_14995,N_14822);
and UO_573 (O_573,N_14778,N_14935);
nor UO_574 (O_574,N_14688,N_14997);
nor UO_575 (O_575,N_14784,N_14632);
or UO_576 (O_576,N_14978,N_14751);
nor UO_577 (O_577,N_14959,N_14788);
nand UO_578 (O_578,N_14753,N_14955);
or UO_579 (O_579,N_14893,N_14673);
and UO_580 (O_580,N_14563,N_14642);
nand UO_581 (O_581,N_14945,N_14925);
or UO_582 (O_582,N_14513,N_14711);
and UO_583 (O_583,N_14542,N_14759);
and UO_584 (O_584,N_14727,N_14661);
nor UO_585 (O_585,N_14622,N_14674);
or UO_586 (O_586,N_14863,N_14670);
nor UO_587 (O_587,N_14505,N_14742);
nor UO_588 (O_588,N_14761,N_14768);
and UO_589 (O_589,N_14860,N_14910);
nor UO_590 (O_590,N_14998,N_14846);
nor UO_591 (O_591,N_14603,N_14812);
and UO_592 (O_592,N_14937,N_14858);
and UO_593 (O_593,N_14707,N_14834);
and UO_594 (O_594,N_14618,N_14514);
nor UO_595 (O_595,N_14846,N_14619);
nor UO_596 (O_596,N_14641,N_14640);
and UO_597 (O_597,N_14890,N_14611);
or UO_598 (O_598,N_14957,N_14601);
xor UO_599 (O_599,N_14835,N_14698);
or UO_600 (O_600,N_14956,N_14977);
or UO_601 (O_601,N_14601,N_14695);
and UO_602 (O_602,N_14555,N_14710);
nor UO_603 (O_603,N_14554,N_14720);
and UO_604 (O_604,N_14652,N_14658);
nand UO_605 (O_605,N_14823,N_14960);
nand UO_606 (O_606,N_14767,N_14741);
and UO_607 (O_607,N_14743,N_14501);
nor UO_608 (O_608,N_14714,N_14833);
and UO_609 (O_609,N_14824,N_14731);
nor UO_610 (O_610,N_14541,N_14577);
nor UO_611 (O_611,N_14917,N_14981);
nor UO_612 (O_612,N_14964,N_14856);
xor UO_613 (O_613,N_14503,N_14941);
nor UO_614 (O_614,N_14759,N_14826);
and UO_615 (O_615,N_14716,N_14888);
nor UO_616 (O_616,N_14968,N_14891);
xor UO_617 (O_617,N_14825,N_14975);
nand UO_618 (O_618,N_14923,N_14897);
nor UO_619 (O_619,N_14781,N_14749);
nor UO_620 (O_620,N_14784,N_14541);
or UO_621 (O_621,N_14799,N_14843);
and UO_622 (O_622,N_14990,N_14930);
or UO_623 (O_623,N_14700,N_14894);
nand UO_624 (O_624,N_14876,N_14857);
or UO_625 (O_625,N_14873,N_14886);
nor UO_626 (O_626,N_14559,N_14709);
nand UO_627 (O_627,N_14679,N_14810);
and UO_628 (O_628,N_14925,N_14611);
nand UO_629 (O_629,N_14528,N_14649);
and UO_630 (O_630,N_14822,N_14828);
and UO_631 (O_631,N_14742,N_14901);
nand UO_632 (O_632,N_14626,N_14685);
and UO_633 (O_633,N_14651,N_14946);
nand UO_634 (O_634,N_14644,N_14649);
nor UO_635 (O_635,N_14945,N_14718);
or UO_636 (O_636,N_14704,N_14745);
or UO_637 (O_637,N_14916,N_14899);
nand UO_638 (O_638,N_14937,N_14971);
and UO_639 (O_639,N_14675,N_14968);
and UO_640 (O_640,N_14620,N_14517);
nor UO_641 (O_641,N_14809,N_14569);
nor UO_642 (O_642,N_14719,N_14578);
and UO_643 (O_643,N_14657,N_14707);
nand UO_644 (O_644,N_14996,N_14926);
and UO_645 (O_645,N_14972,N_14652);
and UO_646 (O_646,N_14895,N_14733);
or UO_647 (O_647,N_14591,N_14686);
nor UO_648 (O_648,N_14874,N_14875);
nor UO_649 (O_649,N_14953,N_14706);
or UO_650 (O_650,N_14778,N_14823);
nor UO_651 (O_651,N_14764,N_14844);
nand UO_652 (O_652,N_14887,N_14677);
nand UO_653 (O_653,N_14667,N_14724);
and UO_654 (O_654,N_14688,N_14763);
nand UO_655 (O_655,N_14671,N_14946);
or UO_656 (O_656,N_14550,N_14670);
or UO_657 (O_657,N_14681,N_14724);
nand UO_658 (O_658,N_14633,N_14763);
nand UO_659 (O_659,N_14974,N_14513);
and UO_660 (O_660,N_14848,N_14912);
nand UO_661 (O_661,N_14752,N_14686);
nor UO_662 (O_662,N_14915,N_14527);
nor UO_663 (O_663,N_14667,N_14706);
xor UO_664 (O_664,N_14981,N_14918);
xor UO_665 (O_665,N_14970,N_14843);
or UO_666 (O_666,N_14666,N_14801);
or UO_667 (O_667,N_14736,N_14989);
nand UO_668 (O_668,N_14961,N_14944);
nand UO_669 (O_669,N_14979,N_14772);
nor UO_670 (O_670,N_14504,N_14615);
nand UO_671 (O_671,N_14592,N_14730);
and UO_672 (O_672,N_14960,N_14870);
nand UO_673 (O_673,N_14580,N_14953);
nand UO_674 (O_674,N_14750,N_14528);
and UO_675 (O_675,N_14722,N_14959);
nand UO_676 (O_676,N_14870,N_14649);
nor UO_677 (O_677,N_14618,N_14625);
nand UO_678 (O_678,N_14734,N_14817);
xor UO_679 (O_679,N_14837,N_14598);
or UO_680 (O_680,N_14972,N_14687);
or UO_681 (O_681,N_14751,N_14878);
nor UO_682 (O_682,N_14604,N_14563);
and UO_683 (O_683,N_14631,N_14733);
and UO_684 (O_684,N_14926,N_14557);
and UO_685 (O_685,N_14649,N_14666);
nand UO_686 (O_686,N_14630,N_14742);
nand UO_687 (O_687,N_14918,N_14845);
nor UO_688 (O_688,N_14661,N_14688);
xor UO_689 (O_689,N_14732,N_14789);
nor UO_690 (O_690,N_14736,N_14735);
and UO_691 (O_691,N_14626,N_14957);
and UO_692 (O_692,N_14825,N_14818);
nand UO_693 (O_693,N_14750,N_14815);
and UO_694 (O_694,N_14612,N_14970);
or UO_695 (O_695,N_14506,N_14670);
nand UO_696 (O_696,N_14925,N_14791);
nor UO_697 (O_697,N_14635,N_14675);
nand UO_698 (O_698,N_14943,N_14823);
nor UO_699 (O_699,N_14959,N_14965);
or UO_700 (O_700,N_14687,N_14708);
nand UO_701 (O_701,N_14869,N_14885);
and UO_702 (O_702,N_14555,N_14944);
or UO_703 (O_703,N_14859,N_14944);
or UO_704 (O_704,N_14956,N_14971);
or UO_705 (O_705,N_14679,N_14951);
and UO_706 (O_706,N_14723,N_14583);
and UO_707 (O_707,N_14982,N_14592);
or UO_708 (O_708,N_14861,N_14624);
and UO_709 (O_709,N_14524,N_14793);
nor UO_710 (O_710,N_14672,N_14517);
nor UO_711 (O_711,N_14949,N_14807);
xor UO_712 (O_712,N_14993,N_14704);
or UO_713 (O_713,N_14776,N_14771);
xnor UO_714 (O_714,N_14548,N_14945);
nand UO_715 (O_715,N_14771,N_14522);
or UO_716 (O_716,N_14837,N_14584);
or UO_717 (O_717,N_14930,N_14718);
or UO_718 (O_718,N_14733,N_14612);
and UO_719 (O_719,N_14961,N_14819);
xor UO_720 (O_720,N_14716,N_14892);
nand UO_721 (O_721,N_14518,N_14523);
or UO_722 (O_722,N_14690,N_14660);
nor UO_723 (O_723,N_14840,N_14604);
or UO_724 (O_724,N_14996,N_14945);
or UO_725 (O_725,N_14791,N_14795);
nor UO_726 (O_726,N_14869,N_14712);
and UO_727 (O_727,N_14993,N_14839);
and UO_728 (O_728,N_14980,N_14531);
nand UO_729 (O_729,N_14878,N_14815);
xor UO_730 (O_730,N_14603,N_14665);
nand UO_731 (O_731,N_14806,N_14556);
nor UO_732 (O_732,N_14645,N_14783);
or UO_733 (O_733,N_14671,N_14653);
nor UO_734 (O_734,N_14778,N_14986);
nand UO_735 (O_735,N_14551,N_14851);
and UO_736 (O_736,N_14551,N_14958);
and UO_737 (O_737,N_14811,N_14517);
and UO_738 (O_738,N_14765,N_14819);
or UO_739 (O_739,N_14970,N_14685);
nor UO_740 (O_740,N_14690,N_14832);
nor UO_741 (O_741,N_14827,N_14590);
nand UO_742 (O_742,N_14803,N_14908);
nand UO_743 (O_743,N_14594,N_14522);
nand UO_744 (O_744,N_14879,N_14814);
nand UO_745 (O_745,N_14692,N_14916);
nand UO_746 (O_746,N_14643,N_14704);
nor UO_747 (O_747,N_14574,N_14781);
or UO_748 (O_748,N_14854,N_14542);
nand UO_749 (O_749,N_14858,N_14601);
xnor UO_750 (O_750,N_14689,N_14589);
and UO_751 (O_751,N_14865,N_14536);
nor UO_752 (O_752,N_14592,N_14643);
nand UO_753 (O_753,N_14747,N_14940);
xor UO_754 (O_754,N_14904,N_14955);
or UO_755 (O_755,N_14563,N_14612);
and UO_756 (O_756,N_14602,N_14715);
and UO_757 (O_757,N_14684,N_14755);
nor UO_758 (O_758,N_14965,N_14642);
or UO_759 (O_759,N_14626,N_14808);
nand UO_760 (O_760,N_14730,N_14683);
nor UO_761 (O_761,N_14515,N_14966);
and UO_762 (O_762,N_14767,N_14638);
nand UO_763 (O_763,N_14895,N_14724);
nor UO_764 (O_764,N_14760,N_14772);
nor UO_765 (O_765,N_14694,N_14916);
nor UO_766 (O_766,N_14799,N_14745);
or UO_767 (O_767,N_14940,N_14624);
nand UO_768 (O_768,N_14870,N_14966);
or UO_769 (O_769,N_14809,N_14756);
and UO_770 (O_770,N_14867,N_14909);
or UO_771 (O_771,N_14679,N_14914);
or UO_772 (O_772,N_14618,N_14727);
nor UO_773 (O_773,N_14601,N_14770);
and UO_774 (O_774,N_14826,N_14650);
or UO_775 (O_775,N_14737,N_14877);
or UO_776 (O_776,N_14700,N_14852);
nand UO_777 (O_777,N_14724,N_14841);
nand UO_778 (O_778,N_14965,N_14659);
or UO_779 (O_779,N_14628,N_14804);
nor UO_780 (O_780,N_14850,N_14616);
nor UO_781 (O_781,N_14875,N_14513);
nor UO_782 (O_782,N_14918,N_14850);
nand UO_783 (O_783,N_14692,N_14867);
or UO_784 (O_784,N_14792,N_14514);
or UO_785 (O_785,N_14960,N_14686);
and UO_786 (O_786,N_14968,N_14628);
nand UO_787 (O_787,N_14734,N_14591);
xor UO_788 (O_788,N_14562,N_14654);
and UO_789 (O_789,N_14872,N_14681);
nor UO_790 (O_790,N_14870,N_14734);
nor UO_791 (O_791,N_14954,N_14538);
nor UO_792 (O_792,N_14927,N_14989);
or UO_793 (O_793,N_14862,N_14820);
nand UO_794 (O_794,N_14860,N_14881);
nand UO_795 (O_795,N_14704,N_14947);
or UO_796 (O_796,N_14723,N_14827);
and UO_797 (O_797,N_14557,N_14854);
and UO_798 (O_798,N_14729,N_14607);
and UO_799 (O_799,N_14748,N_14821);
nand UO_800 (O_800,N_14645,N_14800);
nand UO_801 (O_801,N_14637,N_14953);
xnor UO_802 (O_802,N_14962,N_14917);
and UO_803 (O_803,N_14524,N_14641);
xnor UO_804 (O_804,N_14599,N_14775);
xor UO_805 (O_805,N_14969,N_14689);
or UO_806 (O_806,N_14771,N_14529);
nor UO_807 (O_807,N_14823,N_14501);
and UO_808 (O_808,N_14738,N_14643);
and UO_809 (O_809,N_14933,N_14847);
nand UO_810 (O_810,N_14740,N_14689);
or UO_811 (O_811,N_14967,N_14557);
or UO_812 (O_812,N_14851,N_14590);
nor UO_813 (O_813,N_14771,N_14611);
nor UO_814 (O_814,N_14707,N_14654);
or UO_815 (O_815,N_14543,N_14944);
xor UO_816 (O_816,N_14861,N_14733);
nand UO_817 (O_817,N_14909,N_14842);
nand UO_818 (O_818,N_14899,N_14832);
nor UO_819 (O_819,N_14844,N_14947);
and UO_820 (O_820,N_14937,N_14786);
nand UO_821 (O_821,N_14730,N_14976);
nand UO_822 (O_822,N_14820,N_14931);
nand UO_823 (O_823,N_14952,N_14916);
nor UO_824 (O_824,N_14681,N_14613);
xnor UO_825 (O_825,N_14653,N_14878);
and UO_826 (O_826,N_14612,N_14723);
or UO_827 (O_827,N_14729,N_14832);
xnor UO_828 (O_828,N_14508,N_14731);
or UO_829 (O_829,N_14918,N_14649);
xnor UO_830 (O_830,N_14593,N_14667);
nor UO_831 (O_831,N_14516,N_14958);
nand UO_832 (O_832,N_14620,N_14727);
or UO_833 (O_833,N_14873,N_14566);
nand UO_834 (O_834,N_14785,N_14702);
and UO_835 (O_835,N_14756,N_14806);
and UO_836 (O_836,N_14509,N_14809);
nor UO_837 (O_837,N_14547,N_14826);
and UO_838 (O_838,N_14956,N_14729);
nor UO_839 (O_839,N_14973,N_14958);
or UO_840 (O_840,N_14840,N_14616);
xnor UO_841 (O_841,N_14902,N_14872);
and UO_842 (O_842,N_14571,N_14874);
nor UO_843 (O_843,N_14631,N_14669);
nor UO_844 (O_844,N_14555,N_14672);
xnor UO_845 (O_845,N_14735,N_14837);
and UO_846 (O_846,N_14769,N_14919);
and UO_847 (O_847,N_14692,N_14662);
or UO_848 (O_848,N_14986,N_14530);
nand UO_849 (O_849,N_14660,N_14796);
or UO_850 (O_850,N_14544,N_14774);
or UO_851 (O_851,N_14820,N_14636);
nor UO_852 (O_852,N_14951,N_14650);
and UO_853 (O_853,N_14752,N_14666);
and UO_854 (O_854,N_14774,N_14853);
nand UO_855 (O_855,N_14747,N_14727);
or UO_856 (O_856,N_14608,N_14808);
or UO_857 (O_857,N_14615,N_14808);
and UO_858 (O_858,N_14648,N_14921);
xor UO_859 (O_859,N_14803,N_14848);
or UO_860 (O_860,N_14719,N_14532);
nor UO_861 (O_861,N_14927,N_14948);
nor UO_862 (O_862,N_14896,N_14951);
xor UO_863 (O_863,N_14537,N_14502);
nor UO_864 (O_864,N_14898,N_14802);
xnor UO_865 (O_865,N_14530,N_14725);
nand UO_866 (O_866,N_14550,N_14934);
or UO_867 (O_867,N_14738,N_14776);
and UO_868 (O_868,N_14547,N_14638);
and UO_869 (O_869,N_14607,N_14875);
nor UO_870 (O_870,N_14838,N_14922);
nand UO_871 (O_871,N_14772,N_14690);
or UO_872 (O_872,N_14767,N_14993);
xnor UO_873 (O_873,N_14802,N_14924);
xor UO_874 (O_874,N_14601,N_14644);
nor UO_875 (O_875,N_14813,N_14768);
and UO_876 (O_876,N_14640,N_14718);
or UO_877 (O_877,N_14910,N_14510);
nor UO_878 (O_878,N_14523,N_14507);
or UO_879 (O_879,N_14890,N_14962);
nand UO_880 (O_880,N_14621,N_14635);
xnor UO_881 (O_881,N_14974,N_14601);
xnor UO_882 (O_882,N_14940,N_14893);
nand UO_883 (O_883,N_14927,N_14528);
or UO_884 (O_884,N_14519,N_14608);
nor UO_885 (O_885,N_14936,N_14907);
xnor UO_886 (O_886,N_14612,N_14757);
and UO_887 (O_887,N_14655,N_14962);
or UO_888 (O_888,N_14753,N_14566);
nand UO_889 (O_889,N_14529,N_14685);
or UO_890 (O_890,N_14670,N_14953);
nor UO_891 (O_891,N_14917,N_14733);
and UO_892 (O_892,N_14819,N_14913);
nor UO_893 (O_893,N_14881,N_14597);
and UO_894 (O_894,N_14940,N_14600);
nor UO_895 (O_895,N_14705,N_14915);
nor UO_896 (O_896,N_14617,N_14830);
nor UO_897 (O_897,N_14638,N_14529);
and UO_898 (O_898,N_14583,N_14805);
and UO_899 (O_899,N_14574,N_14758);
nand UO_900 (O_900,N_14804,N_14714);
or UO_901 (O_901,N_14892,N_14511);
and UO_902 (O_902,N_14981,N_14974);
nand UO_903 (O_903,N_14604,N_14683);
and UO_904 (O_904,N_14788,N_14774);
nor UO_905 (O_905,N_14727,N_14816);
nand UO_906 (O_906,N_14769,N_14580);
and UO_907 (O_907,N_14821,N_14540);
nand UO_908 (O_908,N_14773,N_14512);
nor UO_909 (O_909,N_14716,N_14873);
and UO_910 (O_910,N_14760,N_14674);
and UO_911 (O_911,N_14787,N_14641);
nor UO_912 (O_912,N_14702,N_14764);
or UO_913 (O_913,N_14881,N_14575);
nand UO_914 (O_914,N_14843,N_14828);
or UO_915 (O_915,N_14988,N_14744);
or UO_916 (O_916,N_14909,N_14787);
nand UO_917 (O_917,N_14844,N_14839);
nor UO_918 (O_918,N_14565,N_14991);
and UO_919 (O_919,N_14920,N_14620);
and UO_920 (O_920,N_14807,N_14926);
nand UO_921 (O_921,N_14875,N_14925);
nor UO_922 (O_922,N_14916,N_14930);
xor UO_923 (O_923,N_14729,N_14828);
nor UO_924 (O_924,N_14549,N_14925);
or UO_925 (O_925,N_14901,N_14893);
nand UO_926 (O_926,N_14851,N_14670);
nor UO_927 (O_927,N_14544,N_14978);
and UO_928 (O_928,N_14714,N_14739);
or UO_929 (O_929,N_14970,N_14529);
nand UO_930 (O_930,N_14849,N_14906);
nand UO_931 (O_931,N_14503,N_14813);
xor UO_932 (O_932,N_14699,N_14876);
or UO_933 (O_933,N_14616,N_14760);
nor UO_934 (O_934,N_14622,N_14825);
nor UO_935 (O_935,N_14719,N_14929);
nand UO_936 (O_936,N_14894,N_14581);
xor UO_937 (O_937,N_14644,N_14635);
nand UO_938 (O_938,N_14936,N_14595);
xnor UO_939 (O_939,N_14570,N_14674);
nand UO_940 (O_940,N_14932,N_14822);
and UO_941 (O_941,N_14840,N_14693);
and UO_942 (O_942,N_14794,N_14720);
nand UO_943 (O_943,N_14953,N_14999);
or UO_944 (O_944,N_14997,N_14629);
and UO_945 (O_945,N_14590,N_14637);
and UO_946 (O_946,N_14881,N_14598);
or UO_947 (O_947,N_14633,N_14782);
xnor UO_948 (O_948,N_14911,N_14743);
nand UO_949 (O_949,N_14512,N_14722);
nor UO_950 (O_950,N_14714,N_14579);
nor UO_951 (O_951,N_14820,N_14919);
and UO_952 (O_952,N_14855,N_14970);
xnor UO_953 (O_953,N_14568,N_14888);
or UO_954 (O_954,N_14770,N_14801);
and UO_955 (O_955,N_14620,N_14588);
nor UO_956 (O_956,N_14878,N_14957);
xnor UO_957 (O_957,N_14801,N_14809);
or UO_958 (O_958,N_14719,N_14892);
or UO_959 (O_959,N_14650,N_14656);
and UO_960 (O_960,N_14765,N_14559);
and UO_961 (O_961,N_14776,N_14653);
nand UO_962 (O_962,N_14941,N_14947);
nand UO_963 (O_963,N_14620,N_14859);
nor UO_964 (O_964,N_14533,N_14836);
and UO_965 (O_965,N_14899,N_14626);
nor UO_966 (O_966,N_14611,N_14906);
nor UO_967 (O_967,N_14514,N_14901);
nor UO_968 (O_968,N_14825,N_14827);
or UO_969 (O_969,N_14636,N_14868);
nand UO_970 (O_970,N_14870,N_14824);
or UO_971 (O_971,N_14738,N_14808);
and UO_972 (O_972,N_14628,N_14591);
nand UO_973 (O_973,N_14654,N_14818);
or UO_974 (O_974,N_14814,N_14539);
nor UO_975 (O_975,N_14987,N_14838);
nand UO_976 (O_976,N_14780,N_14914);
xor UO_977 (O_977,N_14931,N_14690);
xor UO_978 (O_978,N_14711,N_14724);
nor UO_979 (O_979,N_14590,N_14889);
nor UO_980 (O_980,N_14963,N_14525);
or UO_981 (O_981,N_14982,N_14674);
nor UO_982 (O_982,N_14929,N_14934);
nor UO_983 (O_983,N_14841,N_14556);
or UO_984 (O_984,N_14767,N_14611);
and UO_985 (O_985,N_14922,N_14714);
and UO_986 (O_986,N_14538,N_14772);
xor UO_987 (O_987,N_14543,N_14994);
or UO_988 (O_988,N_14720,N_14839);
or UO_989 (O_989,N_14569,N_14543);
and UO_990 (O_990,N_14616,N_14785);
or UO_991 (O_991,N_14519,N_14713);
xnor UO_992 (O_992,N_14500,N_14930);
nand UO_993 (O_993,N_14755,N_14885);
and UO_994 (O_994,N_14975,N_14833);
nand UO_995 (O_995,N_14618,N_14844);
nor UO_996 (O_996,N_14813,N_14805);
nand UO_997 (O_997,N_14833,N_14900);
nor UO_998 (O_998,N_14951,N_14660);
or UO_999 (O_999,N_14851,N_14639);
or UO_1000 (O_1000,N_14728,N_14687);
nand UO_1001 (O_1001,N_14548,N_14717);
or UO_1002 (O_1002,N_14808,N_14958);
nor UO_1003 (O_1003,N_14798,N_14794);
nor UO_1004 (O_1004,N_14872,N_14907);
and UO_1005 (O_1005,N_14682,N_14694);
xor UO_1006 (O_1006,N_14618,N_14511);
and UO_1007 (O_1007,N_14765,N_14921);
and UO_1008 (O_1008,N_14609,N_14656);
nor UO_1009 (O_1009,N_14680,N_14623);
nor UO_1010 (O_1010,N_14734,N_14623);
nand UO_1011 (O_1011,N_14876,N_14770);
nand UO_1012 (O_1012,N_14974,N_14911);
nor UO_1013 (O_1013,N_14819,N_14541);
and UO_1014 (O_1014,N_14820,N_14964);
nand UO_1015 (O_1015,N_14992,N_14730);
nand UO_1016 (O_1016,N_14807,N_14628);
xor UO_1017 (O_1017,N_14570,N_14996);
and UO_1018 (O_1018,N_14812,N_14847);
nor UO_1019 (O_1019,N_14628,N_14853);
xnor UO_1020 (O_1020,N_14727,N_14784);
xor UO_1021 (O_1021,N_14914,N_14513);
nor UO_1022 (O_1022,N_14820,N_14822);
nand UO_1023 (O_1023,N_14555,N_14870);
and UO_1024 (O_1024,N_14538,N_14637);
or UO_1025 (O_1025,N_14792,N_14672);
nor UO_1026 (O_1026,N_14790,N_14830);
nor UO_1027 (O_1027,N_14678,N_14829);
nand UO_1028 (O_1028,N_14743,N_14515);
or UO_1029 (O_1029,N_14776,N_14937);
and UO_1030 (O_1030,N_14988,N_14708);
and UO_1031 (O_1031,N_14626,N_14639);
nor UO_1032 (O_1032,N_14882,N_14531);
and UO_1033 (O_1033,N_14674,N_14980);
and UO_1034 (O_1034,N_14945,N_14889);
nand UO_1035 (O_1035,N_14863,N_14962);
nor UO_1036 (O_1036,N_14843,N_14501);
nand UO_1037 (O_1037,N_14907,N_14923);
and UO_1038 (O_1038,N_14541,N_14888);
nor UO_1039 (O_1039,N_14562,N_14571);
or UO_1040 (O_1040,N_14875,N_14717);
and UO_1041 (O_1041,N_14636,N_14923);
nor UO_1042 (O_1042,N_14717,N_14703);
nor UO_1043 (O_1043,N_14710,N_14765);
nand UO_1044 (O_1044,N_14760,N_14885);
nor UO_1045 (O_1045,N_14525,N_14798);
nand UO_1046 (O_1046,N_14856,N_14868);
nand UO_1047 (O_1047,N_14927,N_14533);
and UO_1048 (O_1048,N_14672,N_14809);
nand UO_1049 (O_1049,N_14631,N_14757);
or UO_1050 (O_1050,N_14673,N_14812);
nand UO_1051 (O_1051,N_14907,N_14979);
nor UO_1052 (O_1052,N_14835,N_14848);
or UO_1053 (O_1053,N_14869,N_14605);
nor UO_1054 (O_1054,N_14837,N_14712);
or UO_1055 (O_1055,N_14579,N_14815);
xnor UO_1056 (O_1056,N_14611,N_14818);
nand UO_1057 (O_1057,N_14632,N_14814);
nor UO_1058 (O_1058,N_14989,N_14719);
xor UO_1059 (O_1059,N_14590,N_14736);
and UO_1060 (O_1060,N_14934,N_14646);
and UO_1061 (O_1061,N_14601,N_14833);
or UO_1062 (O_1062,N_14594,N_14802);
or UO_1063 (O_1063,N_14889,N_14904);
or UO_1064 (O_1064,N_14841,N_14917);
nand UO_1065 (O_1065,N_14741,N_14935);
nand UO_1066 (O_1066,N_14647,N_14798);
xnor UO_1067 (O_1067,N_14521,N_14855);
nand UO_1068 (O_1068,N_14532,N_14943);
or UO_1069 (O_1069,N_14870,N_14518);
and UO_1070 (O_1070,N_14877,N_14978);
nand UO_1071 (O_1071,N_14847,N_14702);
or UO_1072 (O_1072,N_14993,N_14912);
or UO_1073 (O_1073,N_14765,N_14594);
or UO_1074 (O_1074,N_14984,N_14799);
nand UO_1075 (O_1075,N_14816,N_14841);
nand UO_1076 (O_1076,N_14658,N_14839);
nand UO_1077 (O_1077,N_14997,N_14858);
or UO_1078 (O_1078,N_14858,N_14668);
nor UO_1079 (O_1079,N_14759,N_14538);
xor UO_1080 (O_1080,N_14855,N_14808);
and UO_1081 (O_1081,N_14935,N_14604);
xor UO_1082 (O_1082,N_14567,N_14823);
nand UO_1083 (O_1083,N_14568,N_14834);
nor UO_1084 (O_1084,N_14748,N_14697);
and UO_1085 (O_1085,N_14692,N_14617);
nor UO_1086 (O_1086,N_14826,N_14523);
xor UO_1087 (O_1087,N_14673,N_14871);
nand UO_1088 (O_1088,N_14504,N_14894);
nor UO_1089 (O_1089,N_14892,N_14550);
nand UO_1090 (O_1090,N_14788,N_14845);
or UO_1091 (O_1091,N_14814,N_14906);
and UO_1092 (O_1092,N_14984,N_14808);
xor UO_1093 (O_1093,N_14690,N_14788);
and UO_1094 (O_1094,N_14513,N_14862);
and UO_1095 (O_1095,N_14591,N_14975);
xnor UO_1096 (O_1096,N_14608,N_14799);
and UO_1097 (O_1097,N_14557,N_14630);
nand UO_1098 (O_1098,N_14718,N_14680);
nand UO_1099 (O_1099,N_14588,N_14821);
xor UO_1100 (O_1100,N_14624,N_14990);
and UO_1101 (O_1101,N_14526,N_14640);
and UO_1102 (O_1102,N_14759,N_14583);
or UO_1103 (O_1103,N_14807,N_14510);
and UO_1104 (O_1104,N_14603,N_14994);
or UO_1105 (O_1105,N_14847,N_14834);
or UO_1106 (O_1106,N_14786,N_14734);
or UO_1107 (O_1107,N_14855,N_14943);
nand UO_1108 (O_1108,N_14929,N_14656);
and UO_1109 (O_1109,N_14926,N_14820);
or UO_1110 (O_1110,N_14835,N_14571);
and UO_1111 (O_1111,N_14634,N_14862);
nand UO_1112 (O_1112,N_14820,N_14551);
xnor UO_1113 (O_1113,N_14836,N_14669);
nor UO_1114 (O_1114,N_14630,N_14785);
and UO_1115 (O_1115,N_14890,N_14622);
and UO_1116 (O_1116,N_14774,N_14733);
and UO_1117 (O_1117,N_14874,N_14714);
xor UO_1118 (O_1118,N_14998,N_14545);
or UO_1119 (O_1119,N_14605,N_14531);
nor UO_1120 (O_1120,N_14948,N_14601);
or UO_1121 (O_1121,N_14557,N_14586);
and UO_1122 (O_1122,N_14780,N_14641);
or UO_1123 (O_1123,N_14845,N_14799);
or UO_1124 (O_1124,N_14548,N_14694);
nand UO_1125 (O_1125,N_14805,N_14983);
or UO_1126 (O_1126,N_14973,N_14705);
or UO_1127 (O_1127,N_14729,N_14973);
nor UO_1128 (O_1128,N_14523,N_14921);
nand UO_1129 (O_1129,N_14727,N_14561);
and UO_1130 (O_1130,N_14595,N_14972);
nand UO_1131 (O_1131,N_14580,N_14948);
or UO_1132 (O_1132,N_14520,N_14663);
nand UO_1133 (O_1133,N_14652,N_14984);
nor UO_1134 (O_1134,N_14582,N_14807);
or UO_1135 (O_1135,N_14911,N_14805);
or UO_1136 (O_1136,N_14778,N_14701);
nor UO_1137 (O_1137,N_14534,N_14651);
or UO_1138 (O_1138,N_14558,N_14799);
or UO_1139 (O_1139,N_14865,N_14849);
nand UO_1140 (O_1140,N_14563,N_14627);
and UO_1141 (O_1141,N_14628,N_14510);
nand UO_1142 (O_1142,N_14851,N_14855);
or UO_1143 (O_1143,N_14697,N_14544);
nor UO_1144 (O_1144,N_14990,N_14902);
and UO_1145 (O_1145,N_14997,N_14790);
nor UO_1146 (O_1146,N_14655,N_14916);
or UO_1147 (O_1147,N_14903,N_14539);
and UO_1148 (O_1148,N_14777,N_14675);
and UO_1149 (O_1149,N_14686,N_14995);
xor UO_1150 (O_1150,N_14532,N_14915);
xor UO_1151 (O_1151,N_14806,N_14596);
and UO_1152 (O_1152,N_14872,N_14894);
and UO_1153 (O_1153,N_14627,N_14985);
nor UO_1154 (O_1154,N_14685,N_14611);
and UO_1155 (O_1155,N_14827,N_14744);
xor UO_1156 (O_1156,N_14709,N_14921);
xor UO_1157 (O_1157,N_14600,N_14800);
and UO_1158 (O_1158,N_14564,N_14542);
nor UO_1159 (O_1159,N_14981,N_14944);
or UO_1160 (O_1160,N_14572,N_14728);
nor UO_1161 (O_1161,N_14962,N_14884);
and UO_1162 (O_1162,N_14901,N_14992);
and UO_1163 (O_1163,N_14761,N_14585);
nor UO_1164 (O_1164,N_14594,N_14663);
and UO_1165 (O_1165,N_14940,N_14858);
and UO_1166 (O_1166,N_14521,N_14625);
nand UO_1167 (O_1167,N_14763,N_14640);
and UO_1168 (O_1168,N_14514,N_14818);
xnor UO_1169 (O_1169,N_14666,N_14697);
and UO_1170 (O_1170,N_14536,N_14969);
nor UO_1171 (O_1171,N_14652,N_14866);
nand UO_1172 (O_1172,N_14547,N_14816);
nor UO_1173 (O_1173,N_14634,N_14700);
nand UO_1174 (O_1174,N_14693,N_14740);
and UO_1175 (O_1175,N_14501,N_14551);
xnor UO_1176 (O_1176,N_14550,N_14681);
nand UO_1177 (O_1177,N_14699,N_14828);
and UO_1178 (O_1178,N_14727,N_14500);
nor UO_1179 (O_1179,N_14907,N_14842);
nand UO_1180 (O_1180,N_14662,N_14638);
and UO_1181 (O_1181,N_14834,N_14548);
nand UO_1182 (O_1182,N_14876,N_14725);
or UO_1183 (O_1183,N_14542,N_14511);
nor UO_1184 (O_1184,N_14563,N_14797);
or UO_1185 (O_1185,N_14866,N_14805);
and UO_1186 (O_1186,N_14887,N_14589);
nor UO_1187 (O_1187,N_14865,N_14704);
nor UO_1188 (O_1188,N_14836,N_14713);
and UO_1189 (O_1189,N_14607,N_14554);
and UO_1190 (O_1190,N_14987,N_14815);
nand UO_1191 (O_1191,N_14979,N_14554);
and UO_1192 (O_1192,N_14630,N_14970);
or UO_1193 (O_1193,N_14920,N_14557);
nor UO_1194 (O_1194,N_14708,N_14986);
xor UO_1195 (O_1195,N_14805,N_14778);
or UO_1196 (O_1196,N_14680,N_14712);
nand UO_1197 (O_1197,N_14740,N_14592);
and UO_1198 (O_1198,N_14818,N_14546);
xnor UO_1199 (O_1199,N_14524,N_14874);
and UO_1200 (O_1200,N_14751,N_14520);
nand UO_1201 (O_1201,N_14503,N_14890);
nor UO_1202 (O_1202,N_14671,N_14689);
or UO_1203 (O_1203,N_14533,N_14522);
nand UO_1204 (O_1204,N_14803,N_14927);
nor UO_1205 (O_1205,N_14545,N_14811);
nor UO_1206 (O_1206,N_14562,N_14554);
nor UO_1207 (O_1207,N_14745,N_14988);
nor UO_1208 (O_1208,N_14505,N_14522);
nor UO_1209 (O_1209,N_14921,N_14598);
nand UO_1210 (O_1210,N_14999,N_14905);
and UO_1211 (O_1211,N_14556,N_14824);
nand UO_1212 (O_1212,N_14999,N_14992);
and UO_1213 (O_1213,N_14605,N_14924);
nor UO_1214 (O_1214,N_14764,N_14567);
and UO_1215 (O_1215,N_14983,N_14584);
nand UO_1216 (O_1216,N_14946,N_14625);
nand UO_1217 (O_1217,N_14710,N_14529);
nor UO_1218 (O_1218,N_14910,N_14682);
and UO_1219 (O_1219,N_14604,N_14645);
nor UO_1220 (O_1220,N_14521,N_14501);
nand UO_1221 (O_1221,N_14732,N_14618);
or UO_1222 (O_1222,N_14864,N_14903);
nand UO_1223 (O_1223,N_14610,N_14956);
nand UO_1224 (O_1224,N_14605,N_14648);
or UO_1225 (O_1225,N_14876,N_14569);
nand UO_1226 (O_1226,N_14625,N_14626);
or UO_1227 (O_1227,N_14790,N_14927);
nor UO_1228 (O_1228,N_14514,N_14836);
nor UO_1229 (O_1229,N_14889,N_14808);
or UO_1230 (O_1230,N_14504,N_14770);
nor UO_1231 (O_1231,N_14803,N_14816);
or UO_1232 (O_1232,N_14564,N_14682);
and UO_1233 (O_1233,N_14501,N_14795);
nand UO_1234 (O_1234,N_14912,N_14917);
or UO_1235 (O_1235,N_14773,N_14885);
and UO_1236 (O_1236,N_14968,N_14601);
and UO_1237 (O_1237,N_14893,N_14883);
xor UO_1238 (O_1238,N_14816,N_14584);
and UO_1239 (O_1239,N_14918,N_14767);
nand UO_1240 (O_1240,N_14932,N_14594);
nand UO_1241 (O_1241,N_14884,N_14650);
nand UO_1242 (O_1242,N_14746,N_14711);
or UO_1243 (O_1243,N_14597,N_14622);
and UO_1244 (O_1244,N_14733,N_14869);
xnor UO_1245 (O_1245,N_14559,N_14603);
or UO_1246 (O_1246,N_14981,N_14851);
nand UO_1247 (O_1247,N_14782,N_14891);
nor UO_1248 (O_1248,N_14814,N_14918);
nor UO_1249 (O_1249,N_14762,N_14675);
nand UO_1250 (O_1250,N_14766,N_14783);
or UO_1251 (O_1251,N_14742,N_14930);
or UO_1252 (O_1252,N_14855,N_14504);
xnor UO_1253 (O_1253,N_14553,N_14500);
nor UO_1254 (O_1254,N_14573,N_14628);
and UO_1255 (O_1255,N_14688,N_14779);
nor UO_1256 (O_1256,N_14891,N_14520);
nor UO_1257 (O_1257,N_14881,N_14939);
nor UO_1258 (O_1258,N_14922,N_14727);
nand UO_1259 (O_1259,N_14631,N_14961);
nor UO_1260 (O_1260,N_14501,N_14844);
or UO_1261 (O_1261,N_14734,N_14849);
and UO_1262 (O_1262,N_14535,N_14931);
or UO_1263 (O_1263,N_14590,N_14663);
nand UO_1264 (O_1264,N_14635,N_14649);
nand UO_1265 (O_1265,N_14701,N_14877);
nand UO_1266 (O_1266,N_14609,N_14720);
nor UO_1267 (O_1267,N_14922,N_14902);
and UO_1268 (O_1268,N_14779,N_14733);
and UO_1269 (O_1269,N_14976,N_14705);
nand UO_1270 (O_1270,N_14857,N_14513);
or UO_1271 (O_1271,N_14731,N_14950);
or UO_1272 (O_1272,N_14656,N_14530);
nand UO_1273 (O_1273,N_14869,N_14888);
nand UO_1274 (O_1274,N_14865,N_14754);
nand UO_1275 (O_1275,N_14859,N_14705);
xor UO_1276 (O_1276,N_14662,N_14839);
nand UO_1277 (O_1277,N_14770,N_14675);
or UO_1278 (O_1278,N_14821,N_14543);
or UO_1279 (O_1279,N_14839,N_14989);
nand UO_1280 (O_1280,N_14619,N_14604);
nand UO_1281 (O_1281,N_14861,N_14945);
and UO_1282 (O_1282,N_14639,N_14811);
nor UO_1283 (O_1283,N_14689,N_14822);
nor UO_1284 (O_1284,N_14802,N_14790);
nand UO_1285 (O_1285,N_14828,N_14892);
or UO_1286 (O_1286,N_14835,N_14927);
and UO_1287 (O_1287,N_14510,N_14849);
nand UO_1288 (O_1288,N_14771,N_14681);
and UO_1289 (O_1289,N_14699,N_14737);
nand UO_1290 (O_1290,N_14535,N_14973);
nand UO_1291 (O_1291,N_14998,N_14771);
or UO_1292 (O_1292,N_14944,N_14648);
and UO_1293 (O_1293,N_14633,N_14583);
nor UO_1294 (O_1294,N_14508,N_14933);
and UO_1295 (O_1295,N_14871,N_14931);
nand UO_1296 (O_1296,N_14808,N_14717);
nor UO_1297 (O_1297,N_14602,N_14552);
nor UO_1298 (O_1298,N_14805,N_14678);
nand UO_1299 (O_1299,N_14524,N_14994);
or UO_1300 (O_1300,N_14845,N_14973);
or UO_1301 (O_1301,N_14954,N_14868);
and UO_1302 (O_1302,N_14911,N_14673);
nand UO_1303 (O_1303,N_14741,N_14764);
nand UO_1304 (O_1304,N_14928,N_14777);
nand UO_1305 (O_1305,N_14740,N_14606);
nor UO_1306 (O_1306,N_14611,N_14540);
xnor UO_1307 (O_1307,N_14503,N_14571);
xor UO_1308 (O_1308,N_14516,N_14696);
nand UO_1309 (O_1309,N_14756,N_14985);
nor UO_1310 (O_1310,N_14537,N_14570);
and UO_1311 (O_1311,N_14709,N_14546);
and UO_1312 (O_1312,N_14952,N_14907);
and UO_1313 (O_1313,N_14949,N_14537);
xnor UO_1314 (O_1314,N_14553,N_14952);
xor UO_1315 (O_1315,N_14661,N_14811);
and UO_1316 (O_1316,N_14864,N_14959);
nor UO_1317 (O_1317,N_14519,N_14927);
nor UO_1318 (O_1318,N_14967,N_14875);
nand UO_1319 (O_1319,N_14508,N_14877);
nand UO_1320 (O_1320,N_14504,N_14697);
or UO_1321 (O_1321,N_14856,N_14732);
or UO_1322 (O_1322,N_14507,N_14864);
and UO_1323 (O_1323,N_14538,N_14554);
and UO_1324 (O_1324,N_14680,N_14787);
and UO_1325 (O_1325,N_14619,N_14674);
or UO_1326 (O_1326,N_14701,N_14832);
or UO_1327 (O_1327,N_14731,N_14542);
nor UO_1328 (O_1328,N_14868,N_14614);
nand UO_1329 (O_1329,N_14939,N_14780);
or UO_1330 (O_1330,N_14698,N_14995);
xnor UO_1331 (O_1331,N_14527,N_14874);
and UO_1332 (O_1332,N_14692,N_14956);
xnor UO_1333 (O_1333,N_14522,N_14852);
nand UO_1334 (O_1334,N_14903,N_14990);
nand UO_1335 (O_1335,N_14714,N_14754);
and UO_1336 (O_1336,N_14682,N_14890);
and UO_1337 (O_1337,N_14958,N_14735);
nor UO_1338 (O_1338,N_14592,N_14997);
nand UO_1339 (O_1339,N_14635,N_14671);
and UO_1340 (O_1340,N_14750,N_14995);
xnor UO_1341 (O_1341,N_14507,N_14881);
or UO_1342 (O_1342,N_14679,N_14796);
nand UO_1343 (O_1343,N_14697,N_14536);
nand UO_1344 (O_1344,N_14815,N_14714);
or UO_1345 (O_1345,N_14657,N_14998);
or UO_1346 (O_1346,N_14580,N_14595);
or UO_1347 (O_1347,N_14600,N_14754);
and UO_1348 (O_1348,N_14541,N_14830);
and UO_1349 (O_1349,N_14785,N_14803);
nand UO_1350 (O_1350,N_14600,N_14643);
or UO_1351 (O_1351,N_14893,N_14978);
nor UO_1352 (O_1352,N_14737,N_14788);
and UO_1353 (O_1353,N_14609,N_14716);
nand UO_1354 (O_1354,N_14649,N_14612);
or UO_1355 (O_1355,N_14983,N_14611);
nor UO_1356 (O_1356,N_14707,N_14993);
nor UO_1357 (O_1357,N_14706,N_14884);
xor UO_1358 (O_1358,N_14556,N_14668);
xor UO_1359 (O_1359,N_14913,N_14851);
nand UO_1360 (O_1360,N_14618,N_14659);
xor UO_1361 (O_1361,N_14853,N_14576);
nand UO_1362 (O_1362,N_14935,N_14856);
nand UO_1363 (O_1363,N_14805,N_14636);
or UO_1364 (O_1364,N_14909,N_14851);
nor UO_1365 (O_1365,N_14852,N_14919);
nand UO_1366 (O_1366,N_14540,N_14877);
and UO_1367 (O_1367,N_14776,N_14572);
nand UO_1368 (O_1368,N_14571,N_14822);
nor UO_1369 (O_1369,N_14617,N_14877);
nor UO_1370 (O_1370,N_14810,N_14732);
nor UO_1371 (O_1371,N_14717,N_14658);
nand UO_1372 (O_1372,N_14772,N_14956);
nor UO_1373 (O_1373,N_14980,N_14592);
and UO_1374 (O_1374,N_14725,N_14953);
or UO_1375 (O_1375,N_14986,N_14540);
nand UO_1376 (O_1376,N_14757,N_14639);
and UO_1377 (O_1377,N_14709,N_14595);
nand UO_1378 (O_1378,N_14503,N_14756);
and UO_1379 (O_1379,N_14734,N_14799);
or UO_1380 (O_1380,N_14559,N_14707);
nand UO_1381 (O_1381,N_14928,N_14518);
nand UO_1382 (O_1382,N_14656,N_14585);
nor UO_1383 (O_1383,N_14628,N_14675);
or UO_1384 (O_1384,N_14674,N_14624);
and UO_1385 (O_1385,N_14896,N_14909);
and UO_1386 (O_1386,N_14860,N_14793);
or UO_1387 (O_1387,N_14716,N_14710);
nand UO_1388 (O_1388,N_14614,N_14670);
nand UO_1389 (O_1389,N_14804,N_14592);
nand UO_1390 (O_1390,N_14978,N_14692);
nand UO_1391 (O_1391,N_14615,N_14536);
or UO_1392 (O_1392,N_14839,N_14625);
nand UO_1393 (O_1393,N_14951,N_14627);
and UO_1394 (O_1394,N_14783,N_14743);
or UO_1395 (O_1395,N_14794,N_14793);
or UO_1396 (O_1396,N_14838,N_14920);
nor UO_1397 (O_1397,N_14946,N_14505);
or UO_1398 (O_1398,N_14835,N_14590);
nor UO_1399 (O_1399,N_14810,N_14843);
or UO_1400 (O_1400,N_14667,N_14955);
nand UO_1401 (O_1401,N_14594,N_14525);
and UO_1402 (O_1402,N_14633,N_14899);
nor UO_1403 (O_1403,N_14937,N_14518);
or UO_1404 (O_1404,N_14576,N_14730);
and UO_1405 (O_1405,N_14833,N_14831);
nor UO_1406 (O_1406,N_14598,N_14530);
or UO_1407 (O_1407,N_14503,N_14752);
nand UO_1408 (O_1408,N_14982,N_14728);
nor UO_1409 (O_1409,N_14874,N_14693);
xnor UO_1410 (O_1410,N_14791,N_14851);
xor UO_1411 (O_1411,N_14940,N_14767);
nor UO_1412 (O_1412,N_14767,N_14723);
nor UO_1413 (O_1413,N_14588,N_14602);
nand UO_1414 (O_1414,N_14748,N_14689);
nor UO_1415 (O_1415,N_14907,N_14974);
nand UO_1416 (O_1416,N_14866,N_14843);
nor UO_1417 (O_1417,N_14909,N_14680);
xor UO_1418 (O_1418,N_14815,N_14939);
nor UO_1419 (O_1419,N_14724,N_14784);
nand UO_1420 (O_1420,N_14698,N_14790);
and UO_1421 (O_1421,N_14694,N_14615);
or UO_1422 (O_1422,N_14671,N_14695);
nor UO_1423 (O_1423,N_14749,N_14974);
nand UO_1424 (O_1424,N_14739,N_14950);
nor UO_1425 (O_1425,N_14743,N_14860);
and UO_1426 (O_1426,N_14976,N_14766);
or UO_1427 (O_1427,N_14694,N_14530);
or UO_1428 (O_1428,N_14516,N_14892);
nand UO_1429 (O_1429,N_14890,N_14938);
nor UO_1430 (O_1430,N_14976,N_14722);
or UO_1431 (O_1431,N_14684,N_14511);
xnor UO_1432 (O_1432,N_14763,N_14919);
and UO_1433 (O_1433,N_14755,N_14812);
nand UO_1434 (O_1434,N_14756,N_14582);
and UO_1435 (O_1435,N_14801,N_14818);
nor UO_1436 (O_1436,N_14595,N_14888);
or UO_1437 (O_1437,N_14949,N_14993);
nor UO_1438 (O_1438,N_14816,N_14615);
and UO_1439 (O_1439,N_14581,N_14609);
nand UO_1440 (O_1440,N_14578,N_14948);
nand UO_1441 (O_1441,N_14958,N_14950);
or UO_1442 (O_1442,N_14779,N_14581);
nor UO_1443 (O_1443,N_14625,N_14726);
xnor UO_1444 (O_1444,N_14752,N_14840);
nor UO_1445 (O_1445,N_14557,N_14695);
nand UO_1446 (O_1446,N_14821,N_14509);
nand UO_1447 (O_1447,N_14502,N_14780);
nor UO_1448 (O_1448,N_14837,N_14873);
nor UO_1449 (O_1449,N_14698,N_14941);
or UO_1450 (O_1450,N_14565,N_14756);
nor UO_1451 (O_1451,N_14544,N_14933);
nor UO_1452 (O_1452,N_14574,N_14557);
xnor UO_1453 (O_1453,N_14991,N_14667);
nor UO_1454 (O_1454,N_14737,N_14661);
or UO_1455 (O_1455,N_14595,N_14547);
nand UO_1456 (O_1456,N_14652,N_14569);
nand UO_1457 (O_1457,N_14685,N_14591);
or UO_1458 (O_1458,N_14597,N_14550);
and UO_1459 (O_1459,N_14570,N_14859);
nor UO_1460 (O_1460,N_14640,N_14978);
and UO_1461 (O_1461,N_14760,N_14818);
and UO_1462 (O_1462,N_14645,N_14654);
nor UO_1463 (O_1463,N_14951,N_14601);
nand UO_1464 (O_1464,N_14898,N_14993);
or UO_1465 (O_1465,N_14594,N_14917);
and UO_1466 (O_1466,N_14599,N_14735);
nor UO_1467 (O_1467,N_14589,N_14584);
nor UO_1468 (O_1468,N_14963,N_14917);
and UO_1469 (O_1469,N_14950,N_14821);
xor UO_1470 (O_1470,N_14543,N_14742);
xor UO_1471 (O_1471,N_14779,N_14981);
and UO_1472 (O_1472,N_14982,N_14972);
or UO_1473 (O_1473,N_14860,N_14855);
or UO_1474 (O_1474,N_14848,N_14512);
nand UO_1475 (O_1475,N_14849,N_14516);
or UO_1476 (O_1476,N_14919,N_14816);
nand UO_1477 (O_1477,N_14662,N_14985);
or UO_1478 (O_1478,N_14859,N_14549);
nor UO_1479 (O_1479,N_14634,N_14766);
and UO_1480 (O_1480,N_14607,N_14578);
nor UO_1481 (O_1481,N_14839,N_14509);
nand UO_1482 (O_1482,N_14598,N_14601);
nor UO_1483 (O_1483,N_14572,N_14961);
and UO_1484 (O_1484,N_14993,N_14640);
nor UO_1485 (O_1485,N_14516,N_14921);
xor UO_1486 (O_1486,N_14632,N_14621);
xor UO_1487 (O_1487,N_14874,N_14811);
nand UO_1488 (O_1488,N_14752,N_14890);
or UO_1489 (O_1489,N_14695,N_14783);
nor UO_1490 (O_1490,N_14681,N_14581);
nor UO_1491 (O_1491,N_14621,N_14581);
and UO_1492 (O_1492,N_14928,N_14728);
or UO_1493 (O_1493,N_14705,N_14552);
nor UO_1494 (O_1494,N_14852,N_14994);
or UO_1495 (O_1495,N_14661,N_14610);
nor UO_1496 (O_1496,N_14561,N_14757);
and UO_1497 (O_1497,N_14592,N_14959);
nand UO_1498 (O_1498,N_14923,N_14619);
nor UO_1499 (O_1499,N_14918,N_14664);
nor UO_1500 (O_1500,N_14935,N_14986);
nor UO_1501 (O_1501,N_14717,N_14763);
nor UO_1502 (O_1502,N_14854,N_14621);
and UO_1503 (O_1503,N_14618,N_14842);
nand UO_1504 (O_1504,N_14542,N_14908);
nand UO_1505 (O_1505,N_14983,N_14935);
nand UO_1506 (O_1506,N_14883,N_14581);
or UO_1507 (O_1507,N_14726,N_14578);
and UO_1508 (O_1508,N_14680,N_14583);
nand UO_1509 (O_1509,N_14827,N_14649);
nor UO_1510 (O_1510,N_14999,N_14733);
nor UO_1511 (O_1511,N_14929,N_14981);
or UO_1512 (O_1512,N_14733,N_14929);
nor UO_1513 (O_1513,N_14783,N_14719);
nand UO_1514 (O_1514,N_14949,N_14708);
or UO_1515 (O_1515,N_14634,N_14521);
xnor UO_1516 (O_1516,N_14656,N_14533);
or UO_1517 (O_1517,N_14536,N_14531);
and UO_1518 (O_1518,N_14796,N_14752);
and UO_1519 (O_1519,N_14873,N_14990);
and UO_1520 (O_1520,N_14501,N_14960);
or UO_1521 (O_1521,N_14660,N_14581);
nand UO_1522 (O_1522,N_14633,N_14675);
or UO_1523 (O_1523,N_14502,N_14882);
and UO_1524 (O_1524,N_14924,N_14699);
nor UO_1525 (O_1525,N_14523,N_14895);
nand UO_1526 (O_1526,N_14506,N_14976);
nor UO_1527 (O_1527,N_14626,N_14855);
or UO_1528 (O_1528,N_14984,N_14502);
nor UO_1529 (O_1529,N_14666,N_14644);
and UO_1530 (O_1530,N_14692,N_14849);
or UO_1531 (O_1531,N_14826,N_14651);
nor UO_1532 (O_1532,N_14566,N_14932);
or UO_1533 (O_1533,N_14665,N_14998);
and UO_1534 (O_1534,N_14597,N_14870);
nor UO_1535 (O_1535,N_14634,N_14915);
and UO_1536 (O_1536,N_14909,N_14565);
nor UO_1537 (O_1537,N_14940,N_14924);
nor UO_1538 (O_1538,N_14608,N_14522);
nand UO_1539 (O_1539,N_14581,N_14718);
nand UO_1540 (O_1540,N_14870,N_14641);
or UO_1541 (O_1541,N_14510,N_14826);
or UO_1542 (O_1542,N_14771,N_14846);
nor UO_1543 (O_1543,N_14572,N_14791);
nor UO_1544 (O_1544,N_14542,N_14844);
and UO_1545 (O_1545,N_14584,N_14925);
nor UO_1546 (O_1546,N_14978,N_14858);
and UO_1547 (O_1547,N_14949,N_14735);
and UO_1548 (O_1548,N_14873,N_14697);
xnor UO_1549 (O_1549,N_14780,N_14912);
or UO_1550 (O_1550,N_14634,N_14639);
and UO_1551 (O_1551,N_14767,N_14773);
nand UO_1552 (O_1552,N_14601,N_14891);
and UO_1553 (O_1553,N_14858,N_14888);
or UO_1554 (O_1554,N_14831,N_14978);
nor UO_1555 (O_1555,N_14889,N_14613);
and UO_1556 (O_1556,N_14605,N_14565);
nor UO_1557 (O_1557,N_14510,N_14656);
nor UO_1558 (O_1558,N_14658,N_14635);
nor UO_1559 (O_1559,N_14809,N_14851);
nor UO_1560 (O_1560,N_14665,N_14880);
xnor UO_1561 (O_1561,N_14708,N_14686);
nor UO_1562 (O_1562,N_14887,N_14501);
or UO_1563 (O_1563,N_14843,N_14570);
and UO_1564 (O_1564,N_14628,N_14597);
or UO_1565 (O_1565,N_14981,N_14522);
or UO_1566 (O_1566,N_14599,N_14977);
nand UO_1567 (O_1567,N_14704,N_14639);
nor UO_1568 (O_1568,N_14636,N_14581);
nand UO_1569 (O_1569,N_14839,N_14925);
nor UO_1570 (O_1570,N_14847,N_14527);
and UO_1571 (O_1571,N_14799,N_14547);
nor UO_1572 (O_1572,N_14521,N_14788);
xnor UO_1573 (O_1573,N_14898,N_14819);
nand UO_1574 (O_1574,N_14898,N_14930);
nand UO_1575 (O_1575,N_14981,N_14844);
nand UO_1576 (O_1576,N_14559,N_14746);
xnor UO_1577 (O_1577,N_14896,N_14543);
and UO_1578 (O_1578,N_14684,N_14775);
nand UO_1579 (O_1579,N_14830,N_14554);
or UO_1580 (O_1580,N_14623,N_14869);
xor UO_1581 (O_1581,N_14852,N_14711);
and UO_1582 (O_1582,N_14756,N_14667);
nand UO_1583 (O_1583,N_14754,N_14954);
nor UO_1584 (O_1584,N_14732,N_14737);
and UO_1585 (O_1585,N_14874,N_14568);
xor UO_1586 (O_1586,N_14663,N_14930);
and UO_1587 (O_1587,N_14562,N_14764);
xnor UO_1588 (O_1588,N_14611,N_14736);
and UO_1589 (O_1589,N_14618,N_14686);
and UO_1590 (O_1590,N_14987,N_14714);
or UO_1591 (O_1591,N_14992,N_14868);
or UO_1592 (O_1592,N_14965,N_14991);
nor UO_1593 (O_1593,N_14826,N_14504);
and UO_1594 (O_1594,N_14847,N_14809);
nor UO_1595 (O_1595,N_14799,N_14671);
nor UO_1596 (O_1596,N_14784,N_14606);
nand UO_1597 (O_1597,N_14971,N_14617);
and UO_1598 (O_1598,N_14532,N_14964);
nand UO_1599 (O_1599,N_14709,N_14628);
and UO_1600 (O_1600,N_14572,N_14788);
or UO_1601 (O_1601,N_14524,N_14550);
nand UO_1602 (O_1602,N_14884,N_14838);
nand UO_1603 (O_1603,N_14828,N_14630);
and UO_1604 (O_1604,N_14776,N_14656);
nand UO_1605 (O_1605,N_14827,N_14851);
or UO_1606 (O_1606,N_14638,N_14870);
nor UO_1607 (O_1607,N_14574,N_14689);
or UO_1608 (O_1608,N_14765,N_14663);
nand UO_1609 (O_1609,N_14553,N_14657);
and UO_1610 (O_1610,N_14625,N_14550);
and UO_1611 (O_1611,N_14696,N_14831);
xor UO_1612 (O_1612,N_14911,N_14786);
nand UO_1613 (O_1613,N_14651,N_14559);
or UO_1614 (O_1614,N_14905,N_14624);
nand UO_1615 (O_1615,N_14729,N_14611);
and UO_1616 (O_1616,N_14844,N_14741);
or UO_1617 (O_1617,N_14955,N_14789);
or UO_1618 (O_1618,N_14673,N_14813);
and UO_1619 (O_1619,N_14680,N_14713);
and UO_1620 (O_1620,N_14504,N_14943);
xnor UO_1621 (O_1621,N_14738,N_14608);
nor UO_1622 (O_1622,N_14871,N_14745);
and UO_1623 (O_1623,N_14901,N_14780);
or UO_1624 (O_1624,N_14681,N_14504);
nor UO_1625 (O_1625,N_14748,N_14891);
nand UO_1626 (O_1626,N_14627,N_14587);
nor UO_1627 (O_1627,N_14969,N_14590);
and UO_1628 (O_1628,N_14784,N_14821);
nand UO_1629 (O_1629,N_14697,N_14785);
or UO_1630 (O_1630,N_14543,N_14547);
xor UO_1631 (O_1631,N_14657,N_14632);
and UO_1632 (O_1632,N_14983,N_14528);
nand UO_1633 (O_1633,N_14907,N_14587);
nor UO_1634 (O_1634,N_14967,N_14847);
and UO_1635 (O_1635,N_14739,N_14818);
and UO_1636 (O_1636,N_14500,N_14725);
or UO_1637 (O_1637,N_14674,N_14639);
nand UO_1638 (O_1638,N_14820,N_14951);
xnor UO_1639 (O_1639,N_14580,N_14975);
nand UO_1640 (O_1640,N_14912,N_14829);
nor UO_1641 (O_1641,N_14637,N_14585);
and UO_1642 (O_1642,N_14502,N_14506);
and UO_1643 (O_1643,N_14890,N_14709);
nand UO_1644 (O_1644,N_14750,N_14621);
nor UO_1645 (O_1645,N_14674,N_14906);
nand UO_1646 (O_1646,N_14719,N_14673);
nand UO_1647 (O_1647,N_14880,N_14746);
nand UO_1648 (O_1648,N_14621,N_14514);
or UO_1649 (O_1649,N_14776,N_14963);
and UO_1650 (O_1650,N_14894,N_14957);
nor UO_1651 (O_1651,N_14658,N_14994);
and UO_1652 (O_1652,N_14641,N_14858);
nor UO_1653 (O_1653,N_14883,N_14555);
nand UO_1654 (O_1654,N_14903,N_14875);
nand UO_1655 (O_1655,N_14917,N_14855);
and UO_1656 (O_1656,N_14959,N_14903);
nand UO_1657 (O_1657,N_14782,N_14698);
nand UO_1658 (O_1658,N_14559,N_14597);
or UO_1659 (O_1659,N_14933,N_14872);
nor UO_1660 (O_1660,N_14693,N_14581);
or UO_1661 (O_1661,N_14687,N_14775);
and UO_1662 (O_1662,N_14773,N_14704);
nor UO_1663 (O_1663,N_14796,N_14993);
nor UO_1664 (O_1664,N_14563,N_14898);
and UO_1665 (O_1665,N_14528,N_14878);
and UO_1666 (O_1666,N_14836,N_14826);
nor UO_1667 (O_1667,N_14890,N_14608);
nand UO_1668 (O_1668,N_14579,N_14593);
nand UO_1669 (O_1669,N_14784,N_14996);
nor UO_1670 (O_1670,N_14685,N_14872);
nor UO_1671 (O_1671,N_14915,N_14988);
or UO_1672 (O_1672,N_14604,N_14570);
nand UO_1673 (O_1673,N_14749,N_14775);
nor UO_1674 (O_1674,N_14782,N_14512);
or UO_1675 (O_1675,N_14968,N_14621);
nor UO_1676 (O_1676,N_14837,N_14663);
and UO_1677 (O_1677,N_14794,N_14872);
nor UO_1678 (O_1678,N_14734,N_14981);
and UO_1679 (O_1679,N_14715,N_14793);
xnor UO_1680 (O_1680,N_14750,N_14530);
or UO_1681 (O_1681,N_14586,N_14767);
nor UO_1682 (O_1682,N_14973,N_14952);
nand UO_1683 (O_1683,N_14804,N_14525);
nand UO_1684 (O_1684,N_14653,N_14857);
or UO_1685 (O_1685,N_14580,N_14942);
nor UO_1686 (O_1686,N_14691,N_14568);
or UO_1687 (O_1687,N_14717,N_14862);
nand UO_1688 (O_1688,N_14820,N_14630);
xor UO_1689 (O_1689,N_14856,N_14881);
and UO_1690 (O_1690,N_14586,N_14791);
nand UO_1691 (O_1691,N_14719,N_14858);
and UO_1692 (O_1692,N_14673,N_14973);
xnor UO_1693 (O_1693,N_14942,N_14654);
nand UO_1694 (O_1694,N_14757,N_14786);
nor UO_1695 (O_1695,N_14851,N_14679);
and UO_1696 (O_1696,N_14657,N_14884);
nor UO_1697 (O_1697,N_14955,N_14637);
nand UO_1698 (O_1698,N_14947,N_14952);
or UO_1699 (O_1699,N_14520,N_14689);
nor UO_1700 (O_1700,N_14630,N_14759);
and UO_1701 (O_1701,N_14549,N_14796);
xnor UO_1702 (O_1702,N_14884,N_14864);
and UO_1703 (O_1703,N_14505,N_14536);
and UO_1704 (O_1704,N_14681,N_14695);
and UO_1705 (O_1705,N_14630,N_14911);
or UO_1706 (O_1706,N_14534,N_14906);
and UO_1707 (O_1707,N_14699,N_14827);
nor UO_1708 (O_1708,N_14597,N_14755);
or UO_1709 (O_1709,N_14660,N_14537);
nand UO_1710 (O_1710,N_14639,N_14555);
nor UO_1711 (O_1711,N_14972,N_14814);
nor UO_1712 (O_1712,N_14718,N_14884);
and UO_1713 (O_1713,N_14559,N_14769);
and UO_1714 (O_1714,N_14799,N_14617);
nand UO_1715 (O_1715,N_14637,N_14600);
nand UO_1716 (O_1716,N_14770,N_14682);
nor UO_1717 (O_1717,N_14822,N_14657);
nor UO_1718 (O_1718,N_14753,N_14938);
and UO_1719 (O_1719,N_14794,N_14987);
nor UO_1720 (O_1720,N_14528,N_14963);
nand UO_1721 (O_1721,N_14984,N_14887);
nand UO_1722 (O_1722,N_14579,N_14858);
nor UO_1723 (O_1723,N_14822,N_14927);
nor UO_1724 (O_1724,N_14523,N_14645);
nand UO_1725 (O_1725,N_14585,N_14667);
nand UO_1726 (O_1726,N_14859,N_14890);
xor UO_1727 (O_1727,N_14952,N_14661);
nor UO_1728 (O_1728,N_14614,N_14794);
or UO_1729 (O_1729,N_14870,N_14621);
nor UO_1730 (O_1730,N_14892,N_14804);
and UO_1731 (O_1731,N_14506,N_14738);
or UO_1732 (O_1732,N_14823,N_14967);
nor UO_1733 (O_1733,N_14865,N_14950);
nor UO_1734 (O_1734,N_14642,N_14592);
nand UO_1735 (O_1735,N_14759,N_14878);
and UO_1736 (O_1736,N_14902,N_14786);
nand UO_1737 (O_1737,N_14784,N_14522);
or UO_1738 (O_1738,N_14732,N_14751);
nand UO_1739 (O_1739,N_14538,N_14865);
xor UO_1740 (O_1740,N_14560,N_14933);
or UO_1741 (O_1741,N_14560,N_14839);
or UO_1742 (O_1742,N_14629,N_14889);
and UO_1743 (O_1743,N_14837,N_14591);
and UO_1744 (O_1744,N_14926,N_14978);
nand UO_1745 (O_1745,N_14782,N_14599);
nand UO_1746 (O_1746,N_14547,N_14889);
nor UO_1747 (O_1747,N_14831,N_14713);
nand UO_1748 (O_1748,N_14629,N_14612);
nand UO_1749 (O_1749,N_14920,N_14592);
nor UO_1750 (O_1750,N_14968,N_14630);
or UO_1751 (O_1751,N_14709,N_14926);
and UO_1752 (O_1752,N_14671,N_14613);
and UO_1753 (O_1753,N_14762,N_14791);
and UO_1754 (O_1754,N_14563,N_14587);
nand UO_1755 (O_1755,N_14585,N_14635);
or UO_1756 (O_1756,N_14875,N_14564);
or UO_1757 (O_1757,N_14986,N_14714);
nand UO_1758 (O_1758,N_14770,N_14815);
xnor UO_1759 (O_1759,N_14823,N_14907);
or UO_1760 (O_1760,N_14694,N_14600);
nand UO_1761 (O_1761,N_14794,N_14530);
or UO_1762 (O_1762,N_14981,N_14506);
or UO_1763 (O_1763,N_14605,N_14980);
nor UO_1764 (O_1764,N_14975,N_14715);
nor UO_1765 (O_1765,N_14751,N_14857);
nand UO_1766 (O_1766,N_14869,N_14961);
nand UO_1767 (O_1767,N_14672,N_14929);
or UO_1768 (O_1768,N_14556,N_14669);
nand UO_1769 (O_1769,N_14727,N_14803);
and UO_1770 (O_1770,N_14562,N_14941);
or UO_1771 (O_1771,N_14814,N_14868);
nand UO_1772 (O_1772,N_14703,N_14759);
nand UO_1773 (O_1773,N_14893,N_14802);
and UO_1774 (O_1774,N_14691,N_14660);
and UO_1775 (O_1775,N_14979,N_14559);
nor UO_1776 (O_1776,N_14684,N_14598);
or UO_1777 (O_1777,N_14839,N_14781);
nand UO_1778 (O_1778,N_14997,N_14661);
nand UO_1779 (O_1779,N_14828,N_14620);
nor UO_1780 (O_1780,N_14735,N_14983);
or UO_1781 (O_1781,N_14566,N_14505);
nor UO_1782 (O_1782,N_14592,N_14819);
or UO_1783 (O_1783,N_14538,N_14901);
xor UO_1784 (O_1784,N_14628,N_14639);
nor UO_1785 (O_1785,N_14517,N_14635);
xor UO_1786 (O_1786,N_14675,N_14525);
or UO_1787 (O_1787,N_14653,N_14616);
or UO_1788 (O_1788,N_14533,N_14852);
nor UO_1789 (O_1789,N_14550,N_14882);
nor UO_1790 (O_1790,N_14571,N_14811);
nand UO_1791 (O_1791,N_14792,N_14686);
nand UO_1792 (O_1792,N_14667,N_14901);
and UO_1793 (O_1793,N_14597,N_14695);
nand UO_1794 (O_1794,N_14845,N_14535);
nand UO_1795 (O_1795,N_14926,N_14738);
nand UO_1796 (O_1796,N_14754,N_14800);
xnor UO_1797 (O_1797,N_14658,N_14821);
nor UO_1798 (O_1798,N_14642,N_14628);
nand UO_1799 (O_1799,N_14808,N_14703);
nor UO_1800 (O_1800,N_14687,N_14753);
xor UO_1801 (O_1801,N_14646,N_14912);
nand UO_1802 (O_1802,N_14560,N_14617);
nand UO_1803 (O_1803,N_14814,N_14535);
nand UO_1804 (O_1804,N_14866,N_14741);
nor UO_1805 (O_1805,N_14740,N_14757);
or UO_1806 (O_1806,N_14606,N_14643);
or UO_1807 (O_1807,N_14777,N_14688);
nand UO_1808 (O_1808,N_14774,N_14702);
or UO_1809 (O_1809,N_14898,N_14863);
nor UO_1810 (O_1810,N_14799,N_14766);
nor UO_1811 (O_1811,N_14924,N_14664);
or UO_1812 (O_1812,N_14930,N_14518);
or UO_1813 (O_1813,N_14907,N_14651);
nand UO_1814 (O_1814,N_14775,N_14799);
nor UO_1815 (O_1815,N_14791,N_14626);
nand UO_1816 (O_1816,N_14574,N_14693);
and UO_1817 (O_1817,N_14523,N_14617);
nor UO_1818 (O_1818,N_14596,N_14567);
nor UO_1819 (O_1819,N_14876,N_14806);
and UO_1820 (O_1820,N_14807,N_14600);
and UO_1821 (O_1821,N_14583,N_14672);
or UO_1822 (O_1822,N_14571,N_14621);
xnor UO_1823 (O_1823,N_14968,N_14531);
nand UO_1824 (O_1824,N_14577,N_14545);
and UO_1825 (O_1825,N_14771,N_14667);
and UO_1826 (O_1826,N_14690,N_14645);
nand UO_1827 (O_1827,N_14668,N_14614);
nand UO_1828 (O_1828,N_14729,N_14592);
nor UO_1829 (O_1829,N_14674,N_14819);
nor UO_1830 (O_1830,N_14889,N_14777);
nand UO_1831 (O_1831,N_14919,N_14823);
or UO_1832 (O_1832,N_14625,N_14631);
and UO_1833 (O_1833,N_14826,N_14624);
nor UO_1834 (O_1834,N_14874,N_14531);
xor UO_1835 (O_1835,N_14706,N_14887);
or UO_1836 (O_1836,N_14865,N_14514);
and UO_1837 (O_1837,N_14644,N_14902);
nor UO_1838 (O_1838,N_14624,N_14641);
or UO_1839 (O_1839,N_14600,N_14524);
and UO_1840 (O_1840,N_14511,N_14523);
and UO_1841 (O_1841,N_14674,N_14994);
and UO_1842 (O_1842,N_14843,N_14530);
and UO_1843 (O_1843,N_14868,N_14813);
nor UO_1844 (O_1844,N_14862,N_14711);
nor UO_1845 (O_1845,N_14725,N_14918);
nor UO_1846 (O_1846,N_14901,N_14942);
nand UO_1847 (O_1847,N_14813,N_14810);
and UO_1848 (O_1848,N_14831,N_14650);
nor UO_1849 (O_1849,N_14859,N_14531);
or UO_1850 (O_1850,N_14978,N_14803);
nand UO_1851 (O_1851,N_14963,N_14687);
nand UO_1852 (O_1852,N_14715,N_14993);
nor UO_1853 (O_1853,N_14927,N_14961);
and UO_1854 (O_1854,N_14619,N_14824);
xnor UO_1855 (O_1855,N_14970,N_14814);
and UO_1856 (O_1856,N_14975,N_14804);
nor UO_1857 (O_1857,N_14543,N_14927);
or UO_1858 (O_1858,N_14589,N_14966);
and UO_1859 (O_1859,N_14780,N_14923);
and UO_1860 (O_1860,N_14998,N_14952);
and UO_1861 (O_1861,N_14749,N_14676);
xnor UO_1862 (O_1862,N_14506,N_14969);
nand UO_1863 (O_1863,N_14788,N_14575);
or UO_1864 (O_1864,N_14578,N_14674);
nor UO_1865 (O_1865,N_14543,N_14590);
and UO_1866 (O_1866,N_14711,N_14598);
nor UO_1867 (O_1867,N_14522,N_14907);
nand UO_1868 (O_1868,N_14606,N_14661);
nor UO_1869 (O_1869,N_14683,N_14608);
nor UO_1870 (O_1870,N_14867,N_14549);
xor UO_1871 (O_1871,N_14973,N_14979);
or UO_1872 (O_1872,N_14866,N_14545);
and UO_1873 (O_1873,N_14995,N_14949);
nand UO_1874 (O_1874,N_14984,N_14578);
or UO_1875 (O_1875,N_14747,N_14618);
or UO_1876 (O_1876,N_14687,N_14755);
and UO_1877 (O_1877,N_14585,N_14618);
nor UO_1878 (O_1878,N_14660,N_14559);
or UO_1879 (O_1879,N_14899,N_14886);
or UO_1880 (O_1880,N_14982,N_14755);
nand UO_1881 (O_1881,N_14506,N_14733);
xor UO_1882 (O_1882,N_14781,N_14611);
xnor UO_1883 (O_1883,N_14597,N_14537);
nor UO_1884 (O_1884,N_14663,N_14629);
nor UO_1885 (O_1885,N_14545,N_14767);
nand UO_1886 (O_1886,N_14977,N_14761);
xor UO_1887 (O_1887,N_14588,N_14755);
nor UO_1888 (O_1888,N_14730,N_14562);
and UO_1889 (O_1889,N_14638,N_14731);
or UO_1890 (O_1890,N_14683,N_14778);
nor UO_1891 (O_1891,N_14734,N_14647);
nand UO_1892 (O_1892,N_14757,N_14552);
or UO_1893 (O_1893,N_14653,N_14502);
and UO_1894 (O_1894,N_14689,N_14931);
nand UO_1895 (O_1895,N_14899,N_14639);
and UO_1896 (O_1896,N_14649,N_14984);
xor UO_1897 (O_1897,N_14955,N_14864);
and UO_1898 (O_1898,N_14567,N_14645);
and UO_1899 (O_1899,N_14968,N_14858);
or UO_1900 (O_1900,N_14816,N_14720);
nand UO_1901 (O_1901,N_14978,N_14522);
or UO_1902 (O_1902,N_14964,N_14954);
nand UO_1903 (O_1903,N_14770,N_14993);
nor UO_1904 (O_1904,N_14627,N_14501);
and UO_1905 (O_1905,N_14947,N_14850);
or UO_1906 (O_1906,N_14714,N_14963);
or UO_1907 (O_1907,N_14671,N_14656);
or UO_1908 (O_1908,N_14866,N_14870);
or UO_1909 (O_1909,N_14970,N_14714);
nand UO_1910 (O_1910,N_14635,N_14781);
or UO_1911 (O_1911,N_14705,N_14764);
or UO_1912 (O_1912,N_14945,N_14609);
nand UO_1913 (O_1913,N_14824,N_14694);
or UO_1914 (O_1914,N_14874,N_14519);
nand UO_1915 (O_1915,N_14907,N_14701);
nor UO_1916 (O_1916,N_14715,N_14739);
and UO_1917 (O_1917,N_14678,N_14795);
nor UO_1918 (O_1918,N_14995,N_14854);
nor UO_1919 (O_1919,N_14843,N_14859);
or UO_1920 (O_1920,N_14790,N_14701);
nand UO_1921 (O_1921,N_14534,N_14539);
nand UO_1922 (O_1922,N_14621,N_14644);
nor UO_1923 (O_1923,N_14884,N_14663);
xor UO_1924 (O_1924,N_14995,N_14938);
nand UO_1925 (O_1925,N_14719,N_14556);
or UO_1926 (O_1926,N_14923,N_14848);
and UO_1927 (O_1927,N_14801,N_14755);
and UO_1928 (O_1928,N_14874,N_14937);
nor UO_1929 (O_1929,N_14884,N_14621);
nor UO_1930 (O_1930,N_14812,N_14973);
nor UO_1931 (O_1931,N_14553,N_14685);
nor UO_1932 (O_1932,N_14547,N_14563);
nor UO_1933 (O_1933,N_14993,N_14790);
nor UO_1934 (O_1934,N_14832,N_14835);
or UO_1935 (O_1935,N_14590,N_14914);
and UO_1936 (O_1936,N_14998,N_14770);
nand UO_1937 (O_1937,N_14811,N_14781);
and UO_1938 (O_1938,N_14697,N_14806);
xnor UO_1939 (O_1939,N_14988,N_14759);
and UO_1940 (O_1940,N_14914,N_14843);
or UO_1941 (O_1941,N_14586,N_14594);
and UO_1942 (O_1942,N_14983,N_14928);
nor UO_1943 (O_1943,N_14789,N_14912);
nor UO_1944 (O_1944,N_14938,N_14861);
nand UO_1945 (O_1945,N_14837,N_14512);
nor UO_1946 (O_1946,N_14501,N_14571);
or UO_1947 (O_1947,N_14677,N_14908);
nor UO_1948 (O_1948,N_14593,N_14997);
or UO_1949 (O_1949,N_14680,N_14828);
or UO_1950 (O_1950,N_14916,N_14790);
or UO_1951 (O_1951,N_14955,N_14818);
or UO_1952 (O_1952,N_14807,N_14791);
or UO_1953 (O_1953,N_14568,N_14702);
nor UO_1954 (O_1954,N_14897,N_14930);
nor UO_1955 (O_1955,N_14955,N_14662);
nand UO_1956 (O_1956,N_14672,N_14545);
xnor UO_1957 (O_1957,N_14962,N_14693);
nand UO_1958 (O_1958,N_14947,N_14653);
and UO_1959 (O_1959,N_14525,N_14896);
nor UO_1960 (O_1960,N_14890,N_14917);
nor UO_1961 (O_1961,N_14639,N_14828);
and UO_1962 (O_1962,N_14693,N_14702);
or UO_1963 (O_1963,N_14841,N_14932);
xnor UO_1964 (O_1964,N_14710,N_14898);
and UO_1965 (O_1965,N_14772,N_14555);
and UO_1966 (O_1966,N_14802,N_14917);
and UO_1967 (O_1967,N_14991,N_14947);
nand UO_1968 (O_1968,N_14945,N_14777);
and UO_1969 (O_1969,N_14828,N_14610);
nor UO_1970 (O_1970,N_14920,N_14669);
nor UO_1971 (O_1971,N_14925,N_14741);
nor UO_1972 (O_1972,N_14643,N_14691);
or UO_1973 (O_1973,N_14720,N_14737);
and UO_1974 (O_1974,N_14649,N_14510);
nor UO_1975 (O_1975,N_14887,N_14517);
and UO_1976 (O_1976,N_14563,N_14705);
nor UO_1977 (O_1977,N_14605,N_14940);
xor UO_1978 (O_1978,N_14535,N_14683);
and UO_1979 (O_1979,N_14672,N_14775);
and UO_1980 (O_1980,N_14642,N_14690);
and UO_1981 (O_1981,N_14749,N_14773);
nand UO_1982 (O_1982,N_14888,N_14524);
or UO_1983 (O_1983,N_14937,N_14967);
xnor UO_1984 (O_1984,N_14893,N_14672);
nor UO_1985 (O_1985,N_14548,N_14567);
nor UO_1986 (O_1986,N_14799,N_14834);
nand UO_1987 (O_1987,N_14567,N_14804);
or UO_1988 (O_1988,N_14929,N_14802);
nand UO_1989 (O_1989,N_14922,N_14708);
and UO_1990 (O_1990,N_14962,N_14627);
and UO_1991 (O_1991,N_14919,N_14588);
nand UO_1992 (O_1992,N_14963,N_14946);
nor UO_1993 (O_1993,N_14534,N_14684);
and UO_1994 (O_1994,N_14638,N_14747);
xor UO_1995 (O_1995,N_14504,N_14853);
nand UO_1996 (O_1996,N_14944,N_14828);
nor UO_1997 (O_1997,N_14997,N_14864);
nand UO_1998 (O_1998,N_14736,N_14544);
nor UO_1999 (O_1999,N_14699,N_14808);
endmodule