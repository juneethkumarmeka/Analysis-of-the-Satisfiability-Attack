module basic_2000_20000_2500_20_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nor U0 (N_0,In_1265,In_123);
and U1 (N_1,In_1938,In_696);
nand U2 (N_2,In_191,In_1645);
or U3 (N_3,In_85,In_1154);
nand U4 (N_4,In_572,In_1443);
nor U5 (N_5,In_1200,In_1041);
xor U6 (N_6,In_927,In_517);
nand U7 (N_7,In_308,In_44);
xor U8 (N_8,In_86,In_1741);
and U9 (N_9,In_299,In_1233);
or U10 (N_10,In_364,In_1906);
xnor U11 (N_11,In_1398,In_377);
nand U12 (N_12,In_1325,In_983);
or U13 (N_13,In_1329,In_1498);
and U14 (N_14,In_8,In_1499);
and U15 (N_15,In_1139,In_1280);
xnor U16 (N_16,In_38,In_962);
or U17 (N_17,In_1298,In_1977);
nor U18 (N_18,In_940,In_1501);
nor U19 (N_19,In_1581,In_180);
or U20 (N_20,In_1259,In_627);
nor U21 (N_21,In_617,In_807);
nor U22 (N_22,In_1919,In_45);
or U23 (N_23,In_1676,In_1295);
nand U24 (N_24,In_944,In_839);
nand U25 (N_25,In_501,In_1624);
nand U26 (N_26,In_24,In_272);
xor U27 (N_27,In_888,In_1143);
and U28 (N_28,In_1273,In_1455);
nor U29 (N_29,In_1383,In_1758);
nand U30 (N_30,In_1330,In_1453);
nand U31 (N_31,In_1195,In_535);
xnor U32 (N_32,In_1544,In_613);
nand U33 (N_33,In_217,In_757);
or U34 (N_34,In_1721,In_1780);
nand U35 (N_35,In_1769,In_1983);
nor U36 (N_36,In_656,In_523);
nand U37 (N_37,In_1971,In_1696);
or U38 (N_38,In_285,In_374);
and U39 (N_39,In_1700,In_1852);
xnor U40 (N_40,In_150,In_245);
or U41 (N_41,In_1836,In_1223);
nor U42 (N_42,In_826,In_1937);
xnor U43 (N_43,In_271,In_1691);
and U44 (N_44,In_1240,In_1601);
and U45 (N_45,In_867,In_662);
nor U46 (N_46,In_231,In_1221);
and U47 (N_47,In_718,In_1803);
or U48 (N_48,In_844,In_371);
nor U49 (N_49,In_280,In_1880);
and U50 (N_50,In_225,In_505);
nand U51 (N_51,In_861,In_887);
and U52 (N_52,In_1933,In_152);
xor U53 (N_53,In_636,In_243);
and U54 (N_54,In_83,In_1970);
nand U55 (N_55,In_1695,In_256);
nand U56 (N_56,In_1133,In_1214);
or U57 (N_57,In_904,In_1297);
nand U58 (N_58,In_712,In_1620);
or U59 (N_59,In_520,In_866);
nor U60 (N_60,In_1538,In_65);
nand U61 (N_61,In_604,In_946);
nand U62 (N_62,In_63,In_1738);
nand U63 (N_63,In_71,In_976);
xnor U64 (N_64,In_500,In_898);
nor U65 (N_65,In_1351,In_561);
nand U66 (N_66,In_1791,In_1377);
or U67 (N_67,In_970,In_129);
nand U68 (N_68,In_184,In_1136);
nor U69 (N_69,In_193,In_1596);
and U70 (N_70,In_1343,In_833);
nand U71 (N_71,In_1323,In_1177);
xor U72 (N_72,In_558,In_1489);
nor U73 (N_73,In_282,In_1110);
nand U74 (N_74,In_610,In_507);
nor U75 (N_75,In_682,In_229);
or U76 (N_76,In_390,In_711);
nand U77 (N_77,In_1333,In_1788);
or U78 (N_78,In_676,In_880);
and U79 (N_79,In_1679,In_705);
or U80 (N_80,In_434,In_480);
nand U81 (N_81,In_289,In_1754);
and U82 (N_82,In_1943,In_792);
xnor U83 (N_83,In_1226,In_1474);
nor U84 (N_84,In_619,In_1213);
nor U85 (N_85,In_127,In_1219);
nor U86 (N_86,In_296,In_1655);
nor U87 (N_87,In_1617,In_1135);
and U88 (N_88,In_1885,In_61);
xnor U89 (N_89,In_1484,In_1775);
nand U90 (N_90,In_1465,In_1032);
and U91 (N_91,In_1235,In_181);
or U92 (N_92,In_1089,In_1193);
and U93 (N_93,In_514,In_939);
nand U94 (N_94,In_1069,In_798);
or U95 (N_95,In_665,In_1402);
or U96 (N_96,In_1653,In_144);
nor U97 (N_97,In_1429,In_1868);
and U98 (N_98,In_1512,In_1876);
xnor U99 (N_99,In_7,In_108);
or U100 (N_100,In_1814,In_873);
and U101 (N_101,In_173,In_1988);
xor U102 (N_102,In_1486,In_462);
and U103 (N_103,In_131,In_1423);
nor U104 (N_104,In_226,In_1495);
or U105 (N_105,In_1161,In_725);
or U106 (N_106,In_330,In_418);
nor U107 (N_107,In_550,In_1187);
nor U108 (N_108,In_1610,In_160);
or U109 (N_109,In_1790,In_760);
and U110 (N_110,In_1730,In_466);
nor U111 (N_111,In_835,In_649);
or U112 (N_112,In_1327,In_1651);
or U113 (N_113,In_1397,In_1349);
nand U114 (N_114,In_343,In_993);
nor U115 (N_115,In_1237,In_583);
xor U116 (N_116,In_742,In_1989);
nand U117 (N_117,In_941,In_167);
nor U118 (N_118,In_1516,In_1412);
and U119 (N_119,In_1199,In_1204);
nor U120 (N_120,In_1254,In_305);
xor U121 (N_121,In_1042,In_1153);
nand U122 (N_122,In_1019,In_1766);
xnor U123 (N_123,In_1660,In_774);
nor U124 (N_124,In_1583,In_1144);
nor U125 (N_125,In_1787,In_1936);
xor U126 (N_126,In_128,In_1736);
nand U127 (N_127,In_1373,In_1865);
nand U128 (N_128,In_452,In_678);
xor U129 (N_129,In_761,In_148);
nand U130 (N_130,In_1698,In_1578);
nand U131 (N_131,In_234,In_1785);
or U132 (N_132,In_338,In_9);
nor U133 (N_133,In_259,In_263);
xor U134 (N_134,In_1863,In_879);
and U135 (N_135,In_692,In_1198);
nor U136 (N_136,In_872,In_1071);
nand U137 (N_137,In_1063,In_641);
xnor U138 (N_138,In_821,In_1815);
and U139 (N_139,In_1543,In_97);
or U140 (N_140,In_1682,In_1080);
xnor U141 (N_141,In_281,In_1737);
and U142 (N_142,In_618,In_1843);
or U143 (N_143,In_29,In_1652);
nand U144 (N_144,In_1889,In_727);
xnor U145 (N_145,In_155,In_153);
xnor U146 (N_146,In_413,In_1291);
nor U147 (N_147,In_1001,In_235);
xnor U148 (N_148,In_111,In_415);
xor U149 (N_149,In_936,In_1684);
or U150 (N_150,In_135,In_1269);
nand U151 (N_151,In_1012,In_669);
nand U152 (N_152,In_1091,In_1629);
xor U153 (N_153,In_357,In_1407);
nand U154 (N_154,In_1955,In_776);
and U155 (N_155,In_1303,In_526);
nand U156 (N_156,In_437,In_533);
nand U157 (N_157,In_1656,In_412);
or U158 (N_158,In_713,In_1621);
xnor U159 (N_159,In_52,In_1597);
nor U160 (N_160,In_633,In_901);
and U161 (N_161,In_494,In_1463);
nor U162 (N_162,In_1304,In_102);
nand U163 (N_163,In_1229,In_1745);
nor U164 (N_164,In_1522,In_811);
and U165 (N_165,In_704,In_929);
xnor U166 (N_166,In_699,In_924);
nor U167 (N_167,In_1085,In_1473);
or U168 (N_168,In_1916,In_1371);
xnor U169 (N_169,In_349,In_92);
xor U170 (N_170,In_1793,In_1904);
and U171 (N_171,In_758,In_1644);
or U172 (N_172,In_270,In_744);
and U173 (N_173,In_477,In_1637);
xnor U174 (N_174,In_450,In_841);
or U175 (N_175,In_1894,In_1967);
nor U176 (N_176,In_1452,In_23);
xor U177 (N_177,In_1598,In_333);
nand U178 (N_178,In_1494,In_1996);
xor U179 (N_179,In_883,In_1382);
nor U180 (N_180,In_732,In_1387);
nand U181 (N_181,In_1664,In_518);
or U182 (N_182,In_1277,In_1764);
and U183 (N_183,In_588,In_1215);
xnor U184 (N_184,In_361,In_1432);
or U185 (N_185,In_64,In_1768);
nor U186 (N_186,In_571,In_1286);
xnor U187 (N_187,In_75,In_224);
and U188 (N_188,In_1266,In_47);
or U189 (N_189,In_1997,In_298);
nor U190 (N_190,In_1207,In_1282);
and U191 (N_191,In_15,In_1920);
nand U192 (N_192,In_1564,In_870);
nand U193 (N_193,In_857,In_2);
or U194 (N_194,In_1175,In_750);
xnor U195 (N_195,In_1987,In_239);
nand U196 (N_196,In_1990,In_1514);
or U197 (N_197,In_306,In_88);
xnor U198 (N_198,In_913,In_607);
nor U199 (N_199,In_762,In_1687);
nor U200 (N_200,In_1994,In_141);
nand U201 (N_201,In_765,In_1324);
nand U202 (N_202,In_379,In_1449);
xor U203 (N_203,In_1874,In_287);
nand U204 (N_204,In_1546,In_809);
nand U205 (N_205,In_468,In_1417);
or U206 (N_206,In_1427,In_1929);
and U207 (N_207,In_1444,In_566);
nor U208 (N_208,In_320,In_508);
nor U209 (N_209,In_1457,In_1061);
and U210 (N_210,In_1164,In_815);
nand U211 (N_211,In_1435,In_408);
xor U212 (N_212,In_1934,In_1993);
and U213 (N_213,In_1060,In_1064);
and U214 (N_214,In_50,In_549);
nand U215 (N_215,In_286,In_481);
or U216 (N_216,In_1582,In_174);
and U217 (N_217,In_1833,In_1928);
nand U218 (N_218,In_325,In_441);
or U219 (N_219,In_118,In_1609);
and U220 (N_220,In_892,In_1419);
or U221 (N_221,In_708,In_1886);
xor U222 (N_222,In_852,In_965);
xnor U223 (N_223,In_1249,In_1973);
or U224 (N_224,In_1530,In_1281);
or U225 (N_225,In_159,In_1878);
xor U226 (N_226,In_1718,In_1328);
and U227 (N_227,In_1013,In_130);
xor U228 (N_228,In_474,In_543);
or U229 (N_229,In_1520,In_400);
or U230 (N_230,In_579,In_1146);
and U231 (N_231,In_548,In_856);
xnor U232 (N_232,In_104,In_706);
nor U233 (N_233,In_1563,In_1710);
nor U234 (N_234,In_113,In_1663);
and U235 (N_235,In_733,In_824);
and U236 (N_236,In_1539,In_76);
nand U237 (N_237,In_211,In_1202);
nor U238 (N_238,In_985,In_1336);
nand U239 (N_239,In_1574,In_996);
nand U240 (N_240,In_1572,In_1232);
or U241 (N_241,In_1410,In_10);
nand U242 (N_242,In_989,In_593);
xor U243 (N_243,In_1095,In_203);
and U244 (N_244,In_16,In_1999);
nand U245 (N_245,In_419,In_1593);
nand U246 (N_246,In_56,In_120);
nor U247 (N_247,In_444,In_1339);
nand U248 (N_248,In_176,In_1571);
xnor U249 (N_249,In_464,In_810);
and U250 (N_250,In_915,In_1467);
nor U251 (N_251,In_378,In_1168);
nand U252 (N_252,In_1258,In_726);
nor U253 (N_253,In_254,In_1132);
or U254 (N_254,In_1873,In_1807);
xnor U255 (N_255,In_1116,In_1093);
or U256 (N_256,In_172,In_1600);
and U257 (N_257,In_304,In_398);
and U258 (N_258,In_1121,In_385);
or U259 (N_259,In_1079,In_1702);
nand U260 (N_260,In_1699,In_1912);
nor U261 (N_261,In_1851,In_1502);
nand U262 (N_262,In_1331,In_589);
nor U263 (N_263,In_801,In_802);
and U264 (N_264,In_19,In_43);
and U265 (N_265,In_746,In_1309);
nor U266 (N_266,In_319,In_1547);
xor U267 (N_267,In_1211,In_1005);
xnor U268 (N_268,In_1503,In_1666);
nand U269 (N_269,In_1023,In_1228);
xnor U270 (N_270,In_1421,In_1742);
and U271 (N_271,In_1954,In_580);
nand U272 (N_272,In_958,In_564);
xnor U273 (N_273,In_1713,In_1027);
nand U274 (N_274,In_1898,In_534);
nand U275 (N_275,In_1035,In_592);
or U276 (N_276,In_1853,In_553);
and U277 (N_277,In_702,In_1466);
or U278 (N_278,In_568,In_1065);
and U279 (N_279,In_1350,In_66);
or U280 (N_280,In_685,In_1033);
nand U281 (N_281,In_823,In_647);
nor U282 (N_282,In_205,In_1872);
and U283 (N_283,In_612,In_1053);
nor U284 (N_284,In_1401,In_731);
or U285 (N_285,In_1513,In_206);
nand U286 (N_286,In_322,In_1956);
nor U287 (N_287,In_1585,In_198);
xnor U288 (N_288,In_318,In_640);
nand U289 (N_289,In_1356,In_1589);
nor U290 (N_290,In_1284,In_486);
xnor U291 (N_291,In_1584,In_310);
and U292 (N_292,In_1527,In_1000);
nor U293 (N_293,In_70,In_1756);
xor U294 (N_294,In_295,In_869);
nor U295 (N_295,In_652,In_313);
nand U296 (N_296,In_275,In_1976);
and U297 (N_297,In_812,In_753);
xnor U298 (N_298,In_1267,In_171);
nand U299 (N_299,In_22,In_957);
nor U300 (N_300,In_430,In_951);
nor U301 (N_301,In_1386,In_797);
nor U302 (N_302,In_1839,In_1480);
xnor U303 (N_303,In_1603,In_1818);
nand U304 (N_304,In_1140,In_110);
xor U305 (N_305,In_663,In_1073);
nand U306 (N_306,In_1220,In_1082);
xnor U307 (N_307,In_12,In_825);
nor U308 (N_308,In_1622,In_736);
xor U309 (N_309,In_903,In_264);
nor U310 (N_310,In_445,In_659);
and U311 (N_311,In_1460,In_411);
nor U312 (N_312,In_1899,In_384);
or U313 (N_313,In_1316,In_502);
nor U314 (N_314,In_575,In_1366);
and U315 (N_315,In_701,In_845);
or U316 (N_316,In_294,In_238);
nor U317 (N_317,In_690,In_1347);
or U318 (N_318,In_1641,In_1557);
nor U319 (N_319,In_1192,In_383);
or U320 (N_320,In_541,In_1813);
nor U321 (N_321,In_767,In_233);
nand U322 (N_322,In_747,In_1523);
nand U323 (N_323,In_794,In_1487);
and U324 (N_324,In_1074,In_1831);
xnor U325 (N_325,In_829,In_981);
nor U326 (N_326,In_143,In_1517);
nand U327 (N_327,In_804,In_513);
nand U328 (N_328,In_1126,In_1832);
xnor U329 (N_329,In_563,In_789);
nand U330 (N_330,In_122,In_328);
or U331 (N_331,In_1208,In_1072);
xnor U332 (N_332,In_297,In_849);
or U333 (N_333,In_202,In_1375);
xnor U334 (N_334,In_373,In_1558);
or U335 (N_335,In_599,In_847);
or U336 (N_336,In_1313,In_42);
and U337 (N_337,In_218,In_1978);
nand U338 (N_338,In_168,In_145);
nor U339 (N_339,In_1902,In_1526);
xor U340 (N_340,In_365,In_771);
xor U341 (N_341,In_1828,In_1104);
and U342 (N_342,In_1358,In_1887);
nand U343 (N_343,In_1740,In_1757);
and U344 (N_344,In_695,In_459);
or U345 (N_345,In_1078,In_1850);
and U346 (N_346,In_14,In_414);
and U347 (N_347,In_921,In_854);
xnor U348 (N_348,In_1595,In_1068);
xor U349 (N_349,In_860,In_355);
xor U350 (N_350,In_538,In_600);
nand U351 (N_351,In_1170,In_1521);
xnor U352 (N_352,In_1472,In_269);
or U353 (N_353,In_1234,In_1877);
and U354 (N_354,In_1114,In_1846);
or U355 (N_355,In_625,In_1840);
nand U356 (N_356,In_473,In_995);
xnor U357 (N_357,In_674,In_1210);
xnor U358 (N_358,In_536,In_230);
or U359 (N_359,In_654,In_162);
xor U360 (N_360,In_573,In_782);
nand U361 (N_361,In_142,In_1812);
and U362 (N_362,In_154,In_1418);
nand U363 (N_363,In_734,In_817);
nor U364 (N_364,In_213,In_158);
or U365 (N_365,In_576,In_200);
or U366 (N_366,In_201,In_1657);
nand U367 (N_367,In_999,In_1537);
nor U368 (N_368,In_863,In_27);
xnor U369 (N_369,In_1606,In_209);
nor U370 (N_370,In_114,In_585);
nand U371 (N_371,In_214,In_1364);
and U372 (N_372,In_425,In_1545);
xnor U373 (N_373,In_1442,In_1250);
nor U374 (N_374,In_1,In_1196);
xor U375 (N_375,In_1714,In_342);
xnor U376 (N_376,In_274,In_945);
and U377 (N_377,In_475,In_99);
and U378 (N_378,In_886,In_1026);
and U379 (N_379,In_504,In_1562);
nor U380 (N_380,In_1275,In_1772);
xor U381 (N_381,In_1491,In_1626);
nor U382 (N_382,In_793,In_315);
xor U383 (N_383,In_309,In_1551);
xnor U384 (N_384,In_1142,In_717);
nand U385 (N_385,In_1824,In_1396);
or U386 (N_386,In_442,In_41);
nor U387 (N_387,In_1131,In_994);
nand U388 (N_388,In_1296,In_1554);
nand U389 (N_389,In_1752,In_1774);
nand U390 (N_390,In_1307,In_1561);
nor U391 (N_391,In_1122,In_1524);
or U392 (N_392,In_881,In_1608);
nand U393 (N_393,In_928,In_1395);
xnor U394 (N_394,In_1290,In_1690);
or U395 (N_395,In_1145,In_1535);
and U396 (N_396,In_1166,In_1062);
xnor U397 (N_397,In_1206,In_426);
nand U398 (N_398,In_178,In_1124);
or U399 (N_399,In_1471,In_855);
and U400 (N_400,In_1723,In_407);
and U401 (N_401,In_897,In_116);
nor U402 (N_402,In_766,In_1991);
nor U403 (N_403,In_529,In_1819);
nor U404 (N_404,In_1947,In_1311);
or U405 (N_405,In_1342,In_183);
xnor U406 (N_406,In_133,In_1932);
and U407 (N_407,In_643,In_1217);
nor U408 (N_408,In_488,In_1010);
and U409 (N_409,In_1782,In_1334);
or U410 (N_410,In_843,In_1370);
nand U411 (N_411,In_1454,In_1654);
and U412 (N_412,In_545,In_525);
xnor U413 (N_413,In_1070,In_117);
nand U414 (N_414,In_1761,In_420);
nor U415 (N_415,In_1367,In_257);
or U416 (N_416,In_1119,In_163);
xor U417 (N_417,In_323,In_1821);
nor U418 (N_418,In_1820,In_1972);
nand U419 (N_419,In_859,In_449);
nor U420 (N_420,In_555,In_716);
xor U421 (N_421,In_1568,In_603);
xor U422 (N_422,In_220,In_554);
and U423 (N_423,In_1125,In_1150);
or U424 (N_424,In_1411,In_498);
xor U425 (N_425,In_1239,In_986);
nand U426 (N_426,In_755,In_1923);
or U427 (N_427,In_1209,In_1744);
xnor U428 (N_428,In_1340,In_1577);
or U429 (N_429,In_1504,In_1555);
nand U430 (N_430,In_1279,In_1492);
nor U431 (N_431,In_741,In_650);
nand U432 (N_432,In_1711,In_1260);
nand U433 (N_433,In_5,In_237);
or U434 (N_434,In_1924,In_1253);
nand U435 (N_435,In_1008,In_1525);
or U436 (N_436,In_1216,In_806);
or U437 (N_437,In_1014,In_614);
or U438 (N_438,In_1362,In_1141);
nand U439 (N_439,In_1860,In_1709);
or U440 (N_440,In_925,In_780);
and U441 (N_441,In_1227,In_1246);
or U442 (N_442,In_1058,In_1167);
nor U443 (N_443,In_346,In_1649);
nor U444 (N_444,In_1674,In_288);
or U445 (N_445,In_1570,In_1384);
nor U446 (N_446,In_190,In_165);
or U447 (N_447,In_1188,In_1755);
nor U448 (N_448,In_493,In_611);
and U449 (N_449,In_1909,In_1245);
and U450 (N_450,In_822,In_138);
nor U451 (N_451,In_963,In_1045);
nand U452 (N_452,In_1592,In_1784);
nor U453 (N_453,In_1392,In_1834);
or U454 (N_454,In_1077,In_1781);
and U455 (N_455,In_46,In_703);
and U456 (N_456,In_340,In_341);
nand U457 (N_457,In_1619,In_1779);
and U458 (N_458,In_889,In_503);
or U459 (N_459,In_316,In_1986);
xnor U460 (N_460,In_937,In_516);
or U461 (N_461,In_495,In_393);
nor U462 (N_462,In_509,In_1826);
nor U463 (N_463,In_187,In_1178);
or U464 (N_464,In_483,In_637);
nand U465 (N_465,In_62,In_3);
and U466 (N_466,In_359,In_1565);
nor U467 (N_467,In_952,In_394);
and U468 (N_468,In_1155,In_1439);
nand U469 (N_469,In_1127,In_1952);
or U470 (N_470,In_1390,In_606);
xor U471 (N_471,In_763,In_478);
and U472 (N_472,In_1862,In_1294);
xor U473 (N_473,In_32,In_651);
nand U474 (N_474,In_998,In_506);
and U475 (N_475,In_1433,In_714);
or U476 (N_476,In_1201,In_1315);
nor U477 (N_477,In_101,In_1385);
xnor U478 (N_478,In_1092,In_891);
nand U479 (N_479,In_1369,In_1532);
or U480 (N_480,In_973,In_95);
nand U481 (N_481,In_1067,In_431);
xor U482 (N_482,In_1638,In_1586);
nand U483 (N_483,In_906,In_1083);
and U484 (N_484,In_1515,In_813);
xor U485 (N_485,In_1055,In_842);
or U486 (N_486,In_1251,In_1647);
xnor U487 (N_487,In_1845,In_764);
and U488 (N_488,In_646,In_926);
nand U489 (N_489,In_247,In_730);
and U490 (N_490,In_1891,In_1102);
nor U491 (N_491,In_876,In_689);
or U492 (N_492,In_1770,In_836);
or U493 (N_493,In_1935,In_1478);
xnor U494 (N_494,In_78,In_519);
nor U495 (N_495,In_302,In_1729);
nand U496 (N_496,In_882,In_634);
or U497 (N_497,In_1047,In_490);
xnor U498 (N_498,In_1796,In_1205);
and U499 (N_499,In_1966,In_1022);
nor U500 (N_500,In_253,In_910);
nor U501 (N_501,In_942,In_1255);
nor U502 (N_502,In_1194,In_124);
nand U503 (N_503,In_832,In_1365);
xor U504 (N_504,In_916,In_620);
and U505 (N_505,In_447,In_1483);
and U506 (N_506,In_1300,In_628);
nand U507 (N_507,In_770,In_1725);
or U508 (N_508,In_458,In_1913);
nand U509 (N_509,In_348,In_410);
nand U510 (N_510,In_1158,In_1533);
nand U511 (N_511,In_1485,In_1841);
xor U512 (N_512,In_1867,In_671);
and U513 (N_513,In_1591,In_756);
xnor U514 (N_514,In_1614,In_1389);
and U515 (N_515,In_1859,In_485);
nand U516 (N_516,In_598,In_1426);
xnor U517 (N_517,In_707,In_284);
nand U518 (N_518,In_1482,In_1149);
xor U519 (N_519,In_1271,In_48);
or U520 (N_520,In_984,In_1391);
or U521 (N_521,In_632,In_687);
and U522 (N_522,In_1726,In_820);
and U523 (N_523,In_1917,In_1276);
nor U524 (N_524,In_248,In_1944);
xnor U525 (N_525,In_1939,In_37);
xnor U526 (N_526,In_808,In_20);
nor U527 (N_527,In_1088,In_805);
and U528 (N_528,In_1152,In_814);
and U529 (N_529,In_1009,In_1942);
and U530 (N_530,In_1958,In_1461);
nand U531 (N_531,In_1950,In_1475);
or U532 (N_532,In_642,In_693);
nor U533 (N_533,In_1882,In_356);
xor U534 (N_534,In_666,In_1106);
xnor U535 (N_535,In_956,In_1931);
and U536 (N_536,In_1172,In_1712);
xor U537 (N_537,In_968,In_1985);
xor U538 (N_538,In_551,In_1848);
and U539 (N_539,In_1580,In_51);
nor U540 (N_540,In_1798,In_1907);
nand U541 (N_541,In_1635,In_864);
nor U542 (N_542,In_786,In_1665);
xor U543 (N_543,In_960,In_1308);
xnor U544 (N_544,In_1048,In_236);
or U545 (N_545,In_878,In_595);
nand U546 (N_546,In_1100,In_1021);
nand U547 (N_547,In_546,In_1440);
and U548 (N_548,In_911,In_1029);
nand U549 (N_549,In_1575,In_268);
and U550 (N_550,In_1016,In_743);
nor U551 (N_551,In_376,In_1084);
and U552 (N_552,In_366,In_1688);
or U553 (N_553,In_1184,In_1186);
nand U554 (N_554,In_386,In_653);
and U555 (N_555,In_98,In_453);
nor U556 (N_556,In_82,In_721);
xnor U557 (N_557,In_1030,In_1926);
nand U558 (N_558,In_1374,In_339);
nor U559 (N_559,In_1642,In_1567);
and U560 (N_560,In_1914,In_1951);
nand U561 (N_561,In_997,In_1804);
and U562 (N_562,In_1278,In_1552);
nor U563 (N_563,In_1359,In_719);
or U564 (N_564,In_1922,In_577);
or U565 (N_565,In_1322,In_1668);
nor U566 (N_566,In_277,In_1675);
and U567 (N_567,In_422,In_1372);
xor U568 (N_568,In_250,In_954);
nor U569 (N_569,In_629,In_918);
nand U570 (N_570,In_1871,In_1879);
and U571 (N_571,In_1314,In_739);
or U572 (N_572,In_1101,In_1111);
and U573 (N_573,In_905,In_276);
nand U574 (N_574,In_358,In_871);
nand U575 (N_575,In_1464,In_709);
nand U576 (N_576,In_1884,In_803);
nor U577 (N_577,In_161,In_1236);
and U578 (N_578,In_1505,In_1587);
xnor U579 (N_579,In_421,In_1633);
xor U580 (N_580,In_399,In_1667);
nand U581 (N_581,In_896,In_510);
nand U582 (N_582,In_1519,In_283);
and U583 (N_583,In_935,In_582);
xor U584 (N_584,In_635,In_992);
nand U585 (N_585,In_715,In_428);
nand U586 (N_586,In_1112,In_112);
xnor U587 (N_587,In_179,In_1773);
and U588 (N_588,In_1238,In_1404);
xnor U589 (N_589,In_221,In_93);
xnor U590 (N_590,In_1628,In_1783);
and U591 (N_591,In_1719,In_1961);
and U592 (N_592,In_406,In_18);
xnor U593 (N_593,In_680,In_197);
nand U594 (N_594,In_694,In_748);
nand U595 (N_595,In_1957,In_1908);
xor U596 (N_596,In_1953,In_775);
or U597 (N_597,In_1469,In_991);
or U598 (N_598,In_28,In_436);
and U599 (N_599,In_207,In_1566);
and U600 (N_600,In_433,In_1031);
nand U601 (N_601,In_301,In_397);
or U602 (N_602,In_222,In_1611);
nand U603 (N_603,In_608,In_865);
xor U604 (N_604,In_955,In_948);
nor U605 (N_605,In_1191,In_1960);
or U606 (N_606,In_1827,In_828);
nor U607 (N_607,In_1403,In_1760);
xor U608 (N_608,In_1670,In_1968);
nand U609 (N_609,In_175,In_597);
nor U610 (N_610,In_1794,In_511);
nor U611 (N_611,In_971,In_1844);
or U612 (N_612,In_1648,In_932);
nand U613 (N_613,In_681,In_1735);
and U614 (N_614,In_1422,In_25);
nor U615 (N_615,In_395,In_188);
xnor U616 (N_616,In_1542,In_1076);
nor U617 (N_617,In_1335,In_1470);
and U618 (N_618,In_1293,In_1094);
nor U619 (N_619,In_626,In_858);
xor U620 (N_620,In_499,In_1256);
nand U621 (N_621,In_252,In_1039);
nand U622 (N_622,In_368,In_427);
xnor U623 (N_623,In_964,In_885);
nor U624 (N_624,In_800,In_204);
nand U625 (N_625,In_1056,In_84);
nand U626 (N_626,In_1701,In_1639);
nand U627 (N_627,In_1995,In_1910);
xnor U628 (N_628,In_677,In_1646);
nand U629 (N_629,In_601,In_1394);
and U630 (N_630,In_544,In_1612);
nor U631 (N_631,In_375,In_539);
or U632 (N_632,In_465,In_1376);
xor U633 (N_633,In_125,In_1618);
xnor U634 (N_634,In_291,In_700);
and U635 (N_635,In_1749,In_1531);
xor U636 (N_636,In_210,In_327);
and U637 (N_637,In_773,In_851);
nand U638 (N_638,In_899,In_105);
nor U639 (N_639,In_1751,In_1107);
nand U640 (N_640,In_1715,In_1451);
or U641 (N_641,In_818,In_1822);
or U642 (N_642,In_1559,In_1044);
or U643 (N_643,In_1753,In_265);
nand U644 (N_644,In_482,In_1087);
nor U645 (N_645,In_1345,In_1795);
nand U646 (N_646,In_609,In_470);
xor U647 (N_647,In_664,In_1508);
or U648 (N_648,In_1003,In_369);
xor U649 (N_649,In_581,In_667);
xor U650 (N_650,In_784,In_1534);
nor U651 (N_651,In_1448,In_212);
xnor U652 (N_652,In_1148,In_1805);
or U653 (N_653,In_515,In_121);
nor U654 (N_654,In_260,In_91);
or U655 (N_655,In_1098,In_1911);
or U656 (N_656,In_1979,In_1965);
nand U657 (N_657,In_1855,In_324);
and U658 (N_658,In_1317,In_1147);
nor U659 (N_659,In_391,In_1802);
xor U660 (N_660,In_648,In_1015);
or U661 (N_661,In_1038,In_644);
nor U662 (N_662,In_1707,In_1299);
or U663 (N_663,In_1222,In_846);
and U664 (N_664,In_1692,In_487);
and U665 (N_665,In_1248,In_69);
nand U666 (N_666,In_382,In_68);
or U667 (N_667,In_868,In_219);
and U668 (N_668,In_1103,In_1703);
nand U669 (N_669,In_1890,In_569);
nor U670 (N_670,In_594,In_1927);
and U671 (N_671,In_621,In_1767);
or U672 (N_672,In_830,In_258);
and U673 (N_673,In_273,In_73);
and U674 (N_674,In_1789,In_389);
and U675 (N_675,In_1594,In_722);
xnor U676 (N_676,In_1731,In_759);
nor U677 (N_677,In_132,In_1799);
and U678 (N_678,In_853,In_266);
xnor U679 (N_679,In_920,In_1406);
xor U680 (N_680,In_17,In_1549);
nor U681 (N_681,In_943,In_768);
or U682 (N_682,In_1099,In_166);
nand U683 (N_683,In_360,In_1173);
nand U684 (N_684,In_1728,In_67);
or U685 (N_685,In_1462,In_1497);
nand U686 (N_686,In_908,In_912);
nor U687 (N_687,In_1634,In_909);
and U688 (N_688,In_961,In_317);
or U689 (N_689,In_1287,In_1108);
or U690 (N_690,In_1326,In_1786);
nor U691 (N_691,In_1903,In_454);
or U692 (N_692,In_1881,In_479);
nand U693 (N_693,In_435,In_1430);
and U694 (N_694,In_216,In_1964);
and U695 (N_695,In_1959,In_1476);
and U696 (N_696,In_751,In_720);
nor U697 (N_697,In_326,In_311);
or U698 (N_698,In_403,In_1708);
or U699 (N_699,In_1244,In_424);
or U700 (N_700,In_1312,In_1683);
nand U701 (N_701,In_4,In_1733);
xnor U702 (N_702,In_1837,In_697);
xor U703 (N_703,In_1409,In_1252);
xor U704 (N_704,In_670,In_244);
nand U705 (N_705,In_136,In_79);
or U706 (N_706,In_36,In_931);
nor U707 (N_707,In_1212,In_1134);
or U708 (N_708,In_615,In_30);
and U709 (N_709,In_586,In_416);
xnor U710 (N_710,In_347,In_1866);
or U711 (N_711,In_574,In_1261);
nand U712 (N_712,In_1414,In_87);
or U713 (N_713,In_1176,In_1225);
and U714 (N_714,In_769,In_1050);
nor U715 (N_715,In_1183,In_781);
nor U716 (N_716,In_1732,In_978);
nand U717 (N_717,In_77,In_1579);
and U718 (N_718,In_1727,In_785);
and U719 (N_719,In_89,In_1921);
and U720 (N_720,In_1130,In_1888);
or U721 (N_721,In_1974,In_1247);
or U722 (N_722,In_1096,In_1105);
nor U723 (N_723,In_39,In_907);
xnor U724 (N_724,In_1416,In_1777);
nand U725 (N_725,In_438,In_1590);
nor U726 (N_726,In_914,In_1459);
nand U727 (N_727,In_331,In_969);
xor U728 (N_728,In_31,In_630);
nor U729 (N_729,In_489,In_684);
xnor U730 (N_730,In_1825,In_1477);
nand U731 (N_731,In_698,In_1658);
or U732 (N_732,In_1662,In_557);
nand U733 (N_733,In_950,In_396);
nand U734 (N_734,In_151,In_1129);
nor U735 (N_735,In_605,In_1344);
and U736 (N_736,In_1716,In_1869);
xor U737 (N_737,In_1159,In_1673);
and U738 (N_738,In_215,In_1829);
nand U739 (N_739,In_1722,In_923);
or U740 (N_740,In_409,In_1425);
nand U741 (N_741,In_1493,In_401);
nor U742 (N_742,In_668,In_1174);
nor U743 (N_743,In_1998,In_1607);
and U744 (N_744,In_312,In_570);
and U745 (N_745,In_1036,In_1857);
and U746 (N_746,In_107,In_279);
nand U747 (N_747,In_58,In_1694);
nand U748 (N_748,In_177,In_1066);
or U749 (N_749,In_1361,In_439);
nand U750 (N_750,In_947,In_1685);
or U751 (N_751,In_1569,In_749);
or U752 (N_752,In_1017,In_194);
or U753 (N_753,In_1490,In_537);
nand U754 (N_754,In_779,In_1636);
nand U755 (N_755,In_54,In_1861);
nor U756 (N_756,In_1081,In_1378);
nand U757 (N_757,In_1004,In_33);
or U758 (N_758,In_1338,In_1900);
nor U759 (N_759,In_293,In_1875);
or U760 (N_760,In_457,In_1241);
xnor U761 (N_761,In_1980,In_388);
nor U762 (N_762,In_850,In_816);
nand U763 (N_763,In_1984,In_1856);
and U764 (N_764,In_1588,In_623);
nor U765 (N_765,In_1801,In_1630);
or U766 (N_766,In_837,In_1940);
nor U767 (N_767,In_1858,In_638);
nand U768 (N_768,In_1625,In_189);
nand U769 (N_769,In_1034,In_1059);
and U770 (N_770,In_1759,In_169);
nand U771 (N_771,In_1488,In_754);
and U772 (N_772,In_967,In_522);
and U773 (N_773,In_660,In_890);
nor U774 (N_774,In_21,In_185);
and U775 (N_775,In_922,In_100);
and U776 (N_776,In_1778,In_1550);
xnor U777 (N_777,In_1669,In_1305);
or U778 (N_778,In_448,In_1337);
nand U779 (N_779,In_381,In_156);
nor U780 (N_780,In_241,In_469);
nand U781 (N_781,In_1268,In_772);
and U782 (N_782,In_959,In_367);
xor U783 (N_783,In_884,In_559);
and U784 (N_784,In_332,In_917);
nand U785 (N_785,In_1925,In_1536);
xor U786 (N_786,In_1399,In_1157);
nand U787 (N_787,In_195,In_0);
nor U788 (N_788,In_1018,In_1496);
nand U789 (N_789,In_1816,In_974);
xnor U790 (N_790,In_988,In_1289);
nand U791 (N_791,In_933,In_737);
or U792 (N_792,In_455,In_423);
nor U793 (N_793,In_139,In_1963);
or U794 (N_794,In_1123,In_157);
xor U795 (N_795,In_1156,In_1671);
or U796 (N_796,In_1941,In_1352);
xor U797 (N_797,In_796,In_1128);
and U798 (N_798,In_1697,In_1051);
or U799 (N_799,In_1632,In_895);
and U800 (N_800,In_831,In_930);
nand U801 (N_801,In_686,In_1264);
nor U802 (N_802,In_1540,In_1054);
xnor U803 (N_803,In_26,In_679);
nor U804 (N_804,In_60,In_1842);
or U805 (N_805,In_1945,In_1446);
xnor U806 (N_806,In_1746,In_1434);
nand U807 (N_807,In_1905,In_1037);
nor U808 (N_808,In_673,In_1864);
or U809 (N_809,In_261,In_777);
or U810 (N_810,In_1118,In_1541);
xnor U811 (N_811,In_1481,In_336);
xnor U812 (N_812,In_1203,In_255);
xor U813 (N_813,In_1808,In_838);
and U814 (N_814,In_1318,In_227);
or U815 (N_815,In_1441,In_729);
xor U816 (N_816,In_1509,In_1800);
or U817 (N_817,In_1171,In_392);
nor U818 (N_818,In_1897,In_147);
or U819 (N_819,In_471,In_13);
nand U820 (N_820,In_1830,In_980);
nand U821 (N_821,In_1763,In_990);
xnor U822 (N_822,In_109,In_1981);
nand U823 (N_823,In_303,In_1292);
and U824 (N_824,In_432,In_57);
nand U825 (N_825,In_1163,In_1823);
nor U826 (N_826,In_1776,In_1151);
xor U827 (N_827,In_1704,In_1043);
xor U828 (N_828,In_496,In_476);
nor U829 (N_829,In_875,In_1346);
nand U830 (N_830,In_639,In_1230);
xnor U831 (N_831,In_840,In_1115);
xor U832 (N_832,In_567,In_1388);
nand U833 (N_833,In_446,In_560);
nor U834 (N_834,In_344,In_1189);
or U835 (N_835,In_59,In_710);
xnor U836 (N_836,In_146,In_1243);
nand U837 (N_837,In_405,In_484);
xor U838 (N_838,In_591,In_467);
nor U839 (N_839,In_1901,In_1354);
nand U840 (N_840,In_790,In_34);
nor U841 (N_841,In_1992,In_1306);
nor U842 (N_842,In_1605,In_1854);
and U843 (N_843,In_1659,In_1028);
xor U844 (N_844,In_1348,In_228);
or U845 (N_845,In_1810,In_1479);
nand U846 (N_846,In_1797,In_1762);
nor U847 (N_847,In_350,In_351);
xor U848 (N_848,In_463,In_186);
and U849 (N_849,In_1573,In_1405);
or U850 (N_850,In_1456,In_240);
nand U851 (N_851,In_1379,In_137);
nand U852 (N_852,In_848,In_1870);
nor U853 (N_853,In_1661,In_1020);
nor U854 (N_854,In_1353,In_96);
nand U855 (N_855,In_795,In_1218);
nand U856 (N_856,In_35,In_1368);
or U857 (N_857,In_1893,In_532);
nand U858 (N_858,In_1507,In_1090);
or U859 (N_859,In_372,In_1918);
nand U860 (N_860,In_1892,In_292);
nand U861 (N_861,In_631,In_1915);
nand U862 (N_862,In_352,In_6);
or U863 (N_863,In_1319,In_1556);
and U864 (N_864,In_1310,In_724);
and U865 (N_865,In_745,In_691);
or U866 (N_866,In_1057,In_1182);
nor U867 (N_867,In_80,In_1002);
and U868 (N_868,In_1320,In_1160);
xor U869 (N_869,In_1242,In_672);
or U870 (N_870,In_893,In_752);
or U871 (N_871,In_1458,In_934);
xnor U872 (N_872,In_1982,In_1049);
nor U873 (N_873,In_1678,In_472);
nand U874 (N_874,In_370,In_683);
xnor U875 (N_875,In_440,In_491);
xor U876 (N_876,In_460,In_531);
nor U877 (N_877,In_246,In_81);
and U878 (N_878,In_149,In_1224);
and U879 (N_879,In_267,In_1724);
and U880 (N_880,In_1528,In_979);
or U881 (N_881,In_1748,In_547);
and U882 (N_882,In_307,In_657);
xor U883 (N_883,In_1616,In_223);
xor U884 (N_884,In_874,In_1946);
nand U885 (N_885,In_1285,In_11);
nor U886 (N_886,In_735,In_688);
nor U887 (N_887,In_1190,In_552);
and U888 (N_888,In_1693,In_1720);
or U889 (N_889,In_262,In_1734);
or U890 (N_890,In_354,In_1500);
xnor U891 (N_891,In_1355,In_938);
or U892 (N_892,In_1640,In_1162);
and U893 (N_893,In_1436,In_655);
xor U894 (N_894,In_1809,In_1849);
nand U895 (N_895,In_1270,In_1681);
nand U896 (N_896,In_1896,In_1025);
or U897 (N_897,In_1332,In_1739);
nand U898 (N_898,In_658,In_787);
or U899 (N_899,In_192,In_590);
nor U900 (N_900,In_40,In_1445);
and U901 (N_901,In_126,In_966);
and U902 (N_902,In_987,In_512);
xor U903 (N_903,In_1321,In_1181);
xnor U904 (N_904,In_1949,In_723);
or U905 (N_905,In_791,In_451);
nand U906 (N_906,In_788,In_1302);
and U907 (N_907,In_249,In_778);
nor U908 (N_908,In_1415,In_1506);
xnor U909 (N_909,In_1560,In_456);
nor U910 (N_910,In_1883,In_242);
nor U911 (N_911,In_1180,In_528);
and U912 (N_912,In_1838,In_1717);
or U913 (N_913,In_1510,In_1185);
nand U914 (N_914,In_49,In_1930);
or U915 (N_915,In_94,In_337);
nor U916 (N_916,In_362,In_380);
nand U917 (N_917,In_119,In_1437);
xor U918 (N_918,In_596,In_1447);
xnor U919 (N_919,In_1806,In_1613);
and U920 (N_920,In_170,In_587);
and U921 (N_921,In_1086,In_1381);
nor U922 (N_922,In_740,In_834);
nand U923 (N_923,In_1288,In_602);
or U924 (N_924,In_1962,In_1120);
nand U925 (N_925,In_1529,In_953);
and U926 (N_926,In_1011,In_624);
nand U927 (N_927,In_1518,In_1283);
and U928 (N_928,In_74,In_1046);
or U929 (N_929,In_1771,In_645);
or U930 (N_930,In_1602,In_1792);
nor U931 (N_931,In_53,In_1705);
or U932 (N_932,In_1615,In_562);
xor U933 (N_933,In_461,In_1257);
nor U934 (N_934,In_199,In_1975);
or U935 (N_935,In_1969,In_1274);
nor U936 (N_936,In_1895,In_1847);
xor U937 (N_937,In_232,In_140);
nor U938 (N_938,In_321,In_1075);
nor U939 (N_939,In_675,In_334);
nand U940 (N_940,In_1169,In_497);
or U941 (N_941,In_1599,In_1263);
xor U942 (N_942,In_1817,In_103);
nand U943 (N_943,In_1650,In_819);
nor U944 (N_944,In_182,In_134);
xor U945 (N_945,In_1231,In_1393);
or U946 (N_946,In_1511,In_345);
or U947 (N_947,In_1138,In_977);
and U948 (N_948,In_314,In_877);
nor U949 (N_949,In_975,In_1677);
nand U950 (N_950,In_1631,In_1689);
and U951 (N_951,In_728,In_1413);
or U952 (N_952,In_1007,In_1627);
xor U953 (N_953,In_300,In_530);
nor U954 (N_954,In_542,In_1024);
or U955 (N_955,In_429,In_738);
or U956 (N_956,In_1548,In_1835);
or U957 (N_957,In_164,In_556);
or U958 (N_958,In_949,In_55);
nand U959 (N_959,In_1428,In_1706);
nor U960 (N_960,In_1363,In_919);
nand U961 (N_961,In_894,In_402);
and U962 (N_962,In_115,In_1301);
and U963 (N_963,In_72,In_404);
nor U964 (N_964,In_1109,In_1262);
xnor U965 (N_965,In_278,In_1747);
nand U966 (N_966,In_1137,In_1468);
nor U967 (N_967,In_329,In_1643);
and U968 (N_968,In_616,In_578);
or U969 (N_969,In_1360,In_1006);
xor U970 (N_970,In_208,In_196);
or U971 (N_971,In_1765,In_1686);
or U972 (N_972,In_1623,In_1400);
nor U973 (N_973,In_524,In_862);
xor U974 (N_974,In_1553,In_1811);
or U975 (N_975,In_622,In_902);
or U976 (N_976,In_1948,In_1743);
and U977 (N_977,In_900,In_1576);
or U978 (N_978,In_799,In_1113);
nor U979 (N_979,In_1424,In_565);
nor U980 (N_980,In_1357,In_1680);
or U981 (N_981,In_972,In_1117);
nand U982 (N_982,In_335,In_387);
nor U983 (N_983,In_363,In_1672);
and U984 (N_984,In_353,In_1420);
and U985 (N_985,In_1097,In_1052);
or U986 (N_986,In_584,In_1272);
nand U987 (N_987,In_1438,In_1380);
or U988 (N_988,In_1040,In_521);
or U989 (N_989,In_827,In_290);
nand U990 (N_990,In_251,In_1197);
and U991 (N_991,In_540,In_1750);
or U992 (N_992,In_982,In_1165);
or U993 (N_993,In_90,In_1179);
nand U994 (N_994,In_1341,In_1431);
xor U995 (N_995,In_661,In_783);
xor U996 (N_996,In_527,In_106);
nand U997 (N_997,In_492,In_1408);
xor U998 (N_998,In_1450,In_1604);
xor U999 (N_999,In_443,In_417);
or U1000 (N_1000,N_557,N_854);
nand U1001 (N_1001,N_878,N_542);
nand U1002 (N_1002,N_797,N_720);
nand U1003 (N_1003,N_832,N_287);
and U1004 (N_1004,N_267,N_409);
and U1005 (N_1005,N_957,N_348);
nor U1006 (N_1006,N_572,N_990);
and U1007 (N_1007,N_412,N_15);
nand U1008 (N_1008,N_458,N_440);
nand U1009 (N_1009,N_177,N_326);
xnor U1010 (N_1010,N_928,N_959);
nand U1011 (N_1011,N_489,N_4);
nor U1012 (N_1012,N_783,N_59);
and U1013 (N_1013,N_510,N_951);
xor U1014 (N_1014,N_317,N_387);
xor U1015 (N_1015,N_689,N_104);
nor U1016 (N_1016,N_973,N_723);
nor U1017 (N_1017,N_149,N_869);
xnor U1018 (N_1018,N_618,N_593);
nand U1019 (N_1019,N_891,N_532);
and U1020 (N_1020,N_242,N_760);
xnor U1021 (N_1021,N_987,N_761);
nor U1022 (N_1022,N_327,N_286);
xnor U1023 (N_1023,N_288,N_465);
or U1024 (N_1024,N_230,N_470);
nor U1025 (N_1025,N_768,N_155);
xnor U1026 (N_1026,N_915,N_405);
or U1027 (N_1027,N_274,N_211);
or U1028 (N_1028,N_0,N_164);
xor U1029 (N_1029,N_377,N_328);
and U1030 (N_1030,N_578,N_560);
nand U1031 (N_1031,N_147,N_140);
and U1032 (N_1032,N_993,N_830);
or U1033 (N_1033,N_507,N_715);
nor U1034 (N_1034,N_30,N_127);
nor U1035 (N_1035,N_185,N_635);
nand U1036 (N_1036,N_129,N_918);
and U1037 (N_1037,N_124,N_197);
or U1038 (N_1038,N_673,N_645);
or U1039 (N_1039,N_144,N_693);
xor U1040 (N_1040,N_887,N_270);
xor U1041 (N_1041,N_485,N_240);
xor U1042 (N_1042,N_269,N_17);
or U1043 (N_1043,N_820,N_852);
and U1044 (N_1044,N_904,N_469);
and U1045 (N_1045,N_210,N_359);
nand U1046 (N_1046,N_639,N_498);
and U1047 (N_1047,N_162,N_863);
xnor U1048 (N_1048,N_529,N_655);
xnor U1049 (N_1049,N_91,N_468);
nor U1050 (N_1050,N_422,N_716);
nor U1051 (N_1051,N_912,N_664);
nor U1052 (N_1052,N_259,N_365);
or U1053 (N_1053,N_448,N_695);
and U1054 (N_1054,N_337,N_800);
and U1055 (N_1055,N_674,N_315);
and U1056 (N_1056,N_838,N_116);
and U1057 (N_1057,N_478,N_853);
nor U1058 (N_1058,N_152,N_913);
xnor U1059 (N_1059,N_480,N_921);
nor U1060 (N_1060,N_861,N_748);
nand U1061 (N_1061,N_602,N_681);
or U1062 (N_1062,N_974,N_581);
xnor U1063 (N_1063,N_705,N_61);
xor U1064 (N_1064,N_640,N_552);
nor U1065 (N_1065,N_893,N_601);
or U1066 (N_1066,N_594,N_133);
nor U1067 (N_1067,N_880,N_848);
nand U1068 (N_1068,N_889,N_976);
xnor U1069 (N_1069,N_428,N_879);
or U1070 (N_1070,N_636,N_927);
xnor U1071 (N_1071,N_20,N_989);
nand U1072 (N_1072,N_729,N_86);
xor U1073 (N_1073,N_383,N_855);
nand U1074 (N_1074,N_785,N_910);
nor U1075 (N_1075,N_576,N_379);
or U1076 (N_1076,N_430,N_719);
xnor U1077 (N_1077,N_305,N_410);
nand U1078 (N_1078,N_707,N_517);
or U1079 (N_1079,N_514,N_434);
nand U1080 (N_1080,N_738,N_109);
and U1081 (N_1081,N_427,N_728);
nor U1082 (N_1082,N_805,N_679);
and U1083 (N_1083,N_262,N_304);
nand U1084 (N_1084,N_652,N_93);
nand U1085 (N_1085,N_660,N_174);
nor U1086 (N_1086,N_841,N_402);
nor U1087 (N_1087,N_996,N_416);
nand U1088 (N_1088,N_179,N_366);
nor U1089 (N_1089,N_83,N_876);
nand U1090 (N_1090,N_672,N_318);
and U1091 (N_1091,N_214,N_323);
nand U1092 (N_1092,N_455,N_970);
nor U1093 (N_1093,N_450,N_403);
and U1094 (N_1094,N_226,N_237);
or U1095 (N_1095,N_73,N_435);
nand U1096 (N_1096,N_63,N_941);
nor U1097 (N_1097,N_567,N_68);
nor U1098 (N_1098,N_895,N_49);
xnor U1099 (N_1099,N_90,N_393);
or U1100 (N_1100,N_678,N_342);
nand U1101 (N_1101,N_611,N_914);
nand U1102 (N_1102,N_801,N_472);
xor U1103 (N_1103,N_603,N_616);
or U1104 (N_1104,N_739,N_438);
nand U1105 (N_1105,N_633,N_400);
nand U1106 (N_1106,N_505,N_592);
or U1107 (N_1107,N_453,N_299);
nand U1108 (N_1108,N_96,N_656);
or U1109 (N_1109,N_967,N_630);
and U1110 (N_1110,N_824,N_24);
xor U1111 (N_1111,N_444,N_621);
and U1112 (N_1112,N_826,N_186);
nor U1113 (N_1113,N_734,N_370);
and U1114 (N_1114,N_436,N_141);
xnor U1115 (N_1115,N_559,N_385);
or U1116 (N_1116,N_481,N_721);
and U1117 (N_1117,N_657,N_632);
and U1118 (N_1118,N_971,N_932);
and U1119 (N_1119,N_661,N_651);
nor U1120 (N_1120,N_950,N_804);
nand U1121 (N_1121,N_969,N_421);
and U1122 (N_1122,N_619,N_81);
nor U1123 (N_1123,N_527,N_113);
nor U1124 (N_1124,N_835,N_122);
and U1125 (N_1125,N_992,N_628);
nand U1126 (N_1126,N_271,N_770);
and U1127 (N_1127,N_117,N_997);
and U1128 (N_1128,N_199,N_28);
nor U1129 (N_1129,N_943,N_500);
xnor U1130 (N_1130,N_585,N_683);
and U1131 (N_1131,N_404,N_173);
xor U1132 (N_1132,N_982,N_239);
xnor U1133 (N_1133,N_952,N_35);
and U1134 (N_1134,N_789,N_341);
nor U1135 (N_1135,N_769,N_972);
and U1136 (N_1136,N_154,N_75);
xor U1137 (N_1137,N_792,N_201);
xnor U1138 (N_1138,N_330,N_870);
or U1139 (N_1139,N_846,N_840);
or U1140 (N_1140,N_819,N_871);
nand U1141 (N_1141,N_503,N_419);
nand U1142 (N_1142,N_495,N_775);
xor U1143 (N_1143,N_145,N_136);
and U1144 (N_1144,N_439,N_528);
nor U1145 (N_1145,N_471,N_442);
and U1146 (N_1146,N_275,N_429);
xnor U1147 (N_1147,N_386,N_261);
nand U1148 (N_1148,N_663,N_638);
nor U1149 (N_1149,N_132,N_614);
nand U1150 (N_1150,N_224,N_77);
nand U1151 (N_1151,N_954,N_827);
nor U1152 (N_1152,N_986,N_190);
and U1153 (N_1153,N_725,N_675);
nand U1154 (N_1154,N_196,N_546);
and U1155 (N_1155,N_248,N_361);
or U1156 (N_1156,N_961,N_277);
nor U1157 (N_1157,N_708,N_191);
xor U1158 (N_1158,N_446,N_176);
and U1159 (N_1159,N_965,N_260);
nor U1160 (N_1160,N_968,N_41);
nor U1161 (N_1161,N_977,N_25);
xnor U1162 (N_1162,N_676,N_441);
and U1163 (N_1163,N_245,N_825);
and U1164 (N_1164,N_780,N_53);
xnor U1165 (N_1165,N_839,N_266);
or U1166 (N_1166,N_349,N_713);
nand U1167 (N_1167,N_620,N_740);
or U1168 (N_1168,N_699,N_920);
or U1169 (N_1169,N_169,N_384);
nor U1170 (N_1170,N_627,N_47);
or U1171 (N_1171,N_108,N_733);
nor U1172 (N_1172,N_206,N_903);
xnor U1173 (N_1173,N_212,N_216);
and U1174 (N_1174,N_781,N_795);
or U1175 (N_1175,N_418,N_942);
nor U1176 (N_1176,N_255,N_747);
or U1177 (N_1177,N_979,N_798);
xor U1178 (N_1178,N_231,N_479);
or U1179 (N_1179,N_623,N_896);
and U1180 (N_1180,N_408,N_431);
xor U1181 (N_1181,N_909,N_571);
and U1182 (N_1182,N_555,N_566);
xnor U1183 (N_1183,N_5,N_818);
nand U1184 (N_1184,N_953,N_16);
nand U1185 (N_1185,N_811,N_380);
xor U1186 (N_1186,N_14,N_452);
nor U1187 (N_1187,N_634,N_771);
nand U1188 (N_1188,N_101,N_36);
nand U1189 (N_1189,N_204,N_360);
and U1190 (N_1190,N_29,N_533);
and U1191 (N_1191,N_282,N_238);
nor U1192 (N_1192,N_70,N_934);
or U1193 (N_1193,N_589,N_449);
nand U1194 (N_1194,N_964,N_929);
xnor U1195 (N_1195,N_45,N_232);
nor U1196 (N_1196,N_843,N_935);
nor U1197 (N_1197,N_178,N_482);
xnor U1198 (N_1198,N_369,N_432);
and U1199 (N_1199,N_872,N_494);
and U1200 (N_1200,N_550,N_937);
nand U1201 (N_1201,N_586,N_19);
or U1202 (N_1202,N_121,N_499);
xnor U1203 (N_1203,N_755,N_697);
and U1204 (N_1204,N_849,N_868);
nand U1205 (N_1205,N_900,N_536);
nor U1206 (N_1206,N_724,N_189);
or U1207 (N_1207,N_252,N_72);
xnor U1208 (N_1208,N_40,N_146);
nand U1209 (N_1209,N_44,N_98);
xor U1210 (N_1210,N_235,N_736);
xnor U1211 (N_1211,N_730,N_228);
or U1212 (N_1212,N_765,N_411);
nand U1213 (N_1213,N_549,N_31);
or U1214 (N_1214,N_649,N_758);
nand U1215 (N_1215,N_998,N_847);
or U1216 (N_1216,N_65,N_7);
nor U1217 (N_1217,N_845,N_160);
and U1218 (N_1218,N_751,N_741);
nand U1219 (N_1219,N_57,N_234);
or U1220 (N_1220,N_926,N_375);
nor U1221 (N_1221,N_99,N_873);
or U1222 (N_1222,N_790,N_492);
xnor U1223 (N_1223,N_389,N_391);
nand U1224 (N_1224,N_220,N_772);
nor U1225 (N_1225,N_42,N_281);
nand U1226 (N_1226,N_312,N_483);
nor U1227 (N_1227,N_131,N_322);
or U1228 (N_1228,N_609,N_574);
and U1229 (N_1229,N_130,N_320);
xor U1230 (N_1230,N_960,N_488);
nand U1231 (N_1231,N_850,N_193);
nand U1232 (N_1232,N_423,N_249);
and U1233 (N_1233,N_539,N_62);
and U1234 (N_1234,N_82,N_78);
or U1235 (N_1235,N_321,N_808);
nand U1236 (N_1236,N_759,N_219);
and U1237 (N_1237,N_646,N_749);
nand U1238 (N_1238,N_426,N_491);
nand U1239 (N_1239,N_598,N_666);
xnor U1240 (N_1240,N_222,N_984);
or U1241 (N_1241,N_788,N_263);
or U1242 (N_1242,N_867,N_607);
nand U1243 (N_1243,N_311,N_866);
and U1244 (N_1244,N_744,N_233);
and U1245 (N_1245,N_486,N_936);
and U1246 (N_1246,N_637,N_938);
or U1247 (N_1247,N_278,N_350);
nand U1248 (N_1248,N_991,N_837);
nor U1249 (N_1249,N_540,N_583);
or U1250 (N_1250,N_829,N_244);
or U1251 (N_1251,N_735,N_148);
nor U1252 (N_1252,N_570,N_115);
or U1253 (N_1253,N_836,N_339);
nand U1254 (N_1254,N_816,N_112);
and U1255 (N_1255,N_170,N_163);
nor U1256 (N_1256,N_183,N_156);
xnor U1257 (N_1257,N_851,N_496);
and U1258 (N_1258,N_454,N_319);
nand U1259 (N_1259,N_135,N_258);
and U1260 (N_1260,N_626,N_726);
and U1261 (N_1261,N_347,N_786);
xnor U1262 (N_1262,N_625,N_182);
or U1263 (N_1263,N_21,N_551);
or U1264 (N_1264,N_310,N_84);
nor U1265 (N_1265,N_670,N_501);
xnor U1266 (N_1266,N_512,N_764);
nand U1267 (N_1267,N_906,N_949);
nor U1268 (N_1268,N_692,N_802);
nand U1269 (N_1269,N_324,N_665);
nor U1270 (N_1270,N_3,N_159);
and U1271 (N_1271,N_743,N_945);
xnor U1272 (N_1272,N_213,N_737);
nand U1273 (N_1273,N_296,N_161);
xor U1274 (N_1274,N_300,N_700);
and U1275 (N_1275,N_18,N_823);
and U1276 (N_1276,N_754,N_329);
xor U1277 (N_1277,N_103,N_881);
or U1278 (N_1278,N_886,N_703);
xor U1279 (N_1279,N_158,N_944);
and U1280 (N_1280,N_460,N_834);
or U1281 (N_1281,N_401,N_396);
xor U1282 (N_1282,N_357,N_985);
nor U1283 (N_1283,N_126,N_752);
nand U1284 (N_1284,N_515,N_207);
nor U1285 (N_1285,N_654,N_294);
nand U1286 (N_1286,N_939,N_352);
or U1287 (N_1287,N_487,N_128);
and U1288 (N_1288,N_803,N_92);
nand U1289 (N_1289,N_209,N_413);
nand U1290 (N_1290,N_433,N_898);
nand U1291 (N_1291,N_680,N_958);
nand U1292 (N_1292,N_668,N_691);
and U1293 (N_1293,N_612,N_822);
xnor U1294 (N_1294,N_704,N_604);
nor U1295 (N_1295,N_509,N_995);
nand U1296 (N_1296,N_451,N_882);
nand U1297 (N_1297,N_981,N_208);
and U1298 (N_1298,N_813,N_530);
nand U1299 (N_1299,N_198,N_285);
nor U1300 (N_1300,N_659,N_87);
nand U1301 (N_1301,N_289,N_554);
or U1302 (N_1302,N_476,N_526);
or U1303 (N_1303,N_291,N_301);
or U1304 (N_1304,N_392,N_706);
and U1305 (N_1305,N_746,N_279);
or U1306 (N_1306,N_864,N_605);
and U1307 (N_1307,N_80,N_157);
or U1308 (N_1308,N_187,N_883);
or U1309 (N_1309,N_902,N_241);
and U1310 (N_1310,N_622,N_573);
or U1311 (N_1311,N_946,N_732);
or U1312 (N_1312,N_221,N_246);
xnor U1313 (N_1313,N_38,N_316);
nand U1314 (N_1314,N_22,N_66);
nor U1315 (N_1315,N_833,N_456);
or U1316 (N_1316,N_64,N_667);
and U1317 (N_1317,N_856,N_95);
or U1318 (N_1318,N_363,N_756);
or U1319 (N_1319,N_821,N_71);
xor U1320 (N_1320,N_745,N_37);
nand U1321 (N_1321,N_709,N_26);
and U1322 (N_1322,N_650,N_181);
nor U1323 (N_1323,N_580,N_685);
nor U1324 (N_1324,N_894,N_766);
nor U1325 (N_1325,N_520,N_466);
nand U1326 (N_1326,N_606,N_888);
xor U1327 (N_1327,N_138,N_215);
nor U1328 (N_1328,N_343,N_56);
nor U1329 (N_1329,N_809,N_516);
or U1330 (N_1330,N_50,N_314);
and U1331 (N_1331,N_975,N_857);
and U1332 (N_1332,N_55,N_51);
or U1333 (N_1333,N_710,N_669);
or U1334 (N_1334,N_273,N_257);
nor U1335 (N_1335,N_335,N_265);
and U1336 (N_1336,N_687,N_356);
nor U1337 (N_1337,N_963,N_139);
and U1338 (N_1338,N_79,N_763);
or U1339 (N_1339,N_579,N_1);
nor U1340 (N_1340,N_523,N_338);
or U1341 (N_1341,N_643,N_897);
and U1342 (N_1342,N_791,N_548);
or U1343 (N_1343,N_297,N_563);
and U1344 (N_1344,N_647,N_497);
and U1345 (N_1345,N_123,N_955);
and U1346 (N_1346,N_617,N_194);
nand U1347 (N_1347,N_569,N_223);
and U1348 (N_1348,N_437,N_52);
nand U1349 (N_1349,N_877,N_597);
nand U1350 (N_1350,N_653,N_899);
or U1351 (N_1351,N_308,N_97);
and U1352 (N_1352,N_599,N_94);
nor U1353 (N_1353,N_12,N_376);
nor U1354 (N_1354,N_462,N_671);
nor U1355 (N_1355,N_587,N_544);
nand U1356 (N_1356,N_718,N_925);
or U1357 (N_1357,N_556,N_908);
or U1358 (N_1358,N_812,N_168);
or U1359 (N_1359,N_388,N_577);
nand U1360 (N_1360,N_662,N_43);
and U1361 (N_1361,N_511,N_331);
and U1362 (N_1362,N_205,N_373);
nand U1363 (N_1363,N_293,N_782);
nand U1364 (N_1364,N_200,N_796);
nand U1365 (N_1365,N_742,N_842);
nor U1366 (N_1366,N_537,N_506);
nor U1367 (N_1367,N_398,N_309);
xnor U1368 (N_1368,N_930,N_793);
or U1369 (N_1369,N_2,N_844);
nor U1370 (N_1370,N_484,N_336);
nand U1371 (N_1371,N_712,N_966);
and U1372 (N_1372,N_447,N_333);
nand U1373 (N_1373,N_727,N_568);
and U1374 (N_1374,N_415,N_931);
and U1375 (N_1375,N_947,N_890);
nand U1376 (N_1376,N_23,N_541);
or U1377 (N_1377,N_151,N_777);
nor U1378 (N_1378,N_58,N_615);
nor U1379 (N_1379,N_48,N_688);
xor U1380 (N_1380,N_106,N_773);
and U1381 (N_1381,N_831,N_648);
or U1382 (N_1382,N_558,N_518);
nand U1383 (N_1383,N_88,N_332);
or U1384 (N_1384,N_767,N_280);
nand U1385 (N_1385,N_610,N_254);
nand U1386 (N_1386,N_394,N_407);
or U1387 (N_1387,N_828,N_111);
xnor U1388 (N_1388,N_988,N_283);
or U1389 (N_1389,N_702,N_74);
nor U1390 (N_1390,N_717,N_658);
and U1391 (N_1391,N_776,N_247);
and U1392 (N_1392,N_757,N_67);
nand U1393 (N_1393,N_120,N_420);
nor U1394 (N_1394,N_862,N_504);
nor U1395 (N_1395,N_980,N_46);
or U1396 (N_1396,N_368,N_325);
nor U1397 (N_1397,N_60,N_100);
xor U1398 (N_1398,N_39,N_217);
xor U1399 (N_1399,N_250,N_358);
or U1400 (N_1400,N_110,N_166);
xor U1401 (N_1401,N_694,N_810);
nor U1402 (N_1402,N_817,N_543);
or U1403 (N_1403,N_519,N_613);
nor U1404 (N_1404,N_701,N_295);
nor U1405 (N_1405,N_521,N_11);
and U1406 (N_1406,N_445,N_753);
xnor U1407 (N_1407,N_180,N_364);
nor U1408 (N_1408,N_171,N_414);
nand U1409 (N_1409,N_531,N_784);
and U1410 (N_1410,N_268,N_397);
and U1411 (N_1411,N_584,N_714);
xnor U1412 (N_1412,N_535,N_892);
xnor U1413 (N_1413,N_962,N_994);
nand U1414 (N_1414,N_901,N_188);
and U1415 (N_1415,N_778,N_983);
nand U1416 (N_1416,N_565,N_334);
xnor U1417 (N_1417,N_195,N_313);
xnor U1418 (N_1418,N_225,N_229);
nor U1419 (N_1419,N_192,N_682);
nand U1420 (N_1420,N_134,N_371);
xor U1421 (N_1421,N_590,N_424);
nor U1422 (N_1422,N_911,N_362);
nor U1423 (N_1423,N_490,N_508);
nor U1424 (N_1424,N_545,N_165);
nand U1425 (N_1425,N_919,N_306);
nand U1426 (N_1426,N_474,N_54);
nand U1427 (N_1427,N_762,N_473);
or U1428 (N_1428,N_390,N_76);
nor U1429 (N_1429,N_524,N_464);
or U1430 (N_1430,N_354,N_292);
nand U1431 (N_1431,N_6,N_722);
and U1432 (N_1432,N_562,N_32);
nand U1433 (N_1433,N_395,N_353);
and U1434 (N_1434,N_114,N_779);
nand U1435 (N_1435,N_600,N_696);
nand U1436 (N_1436,N_493,N_10);
nand U1437 (N_1437,N_582,N_107);
nand U1438 (N_1438,N_502,N_874);
nor U1439 (N_1439,N_875,N_642);
xnor U1440 (N_1440,N_561,N_253);
nand U1441 (N_1441,N_340,N_34);
or U1442 (N_1442,N_102,N_806);
or U1443 (N_1443,N_443,N_956);
nand U1444 (N_1444,N_425,N_774);
and U1445 (N_1445,N_203,N_89);
nor U1446 (N_1446,N_463,N_351);
nor U1447 (N_1447,N_142,N_538);
and U1448 (N_1448,N_399,N_475);
nor U1449 (N_1449,N_940,N_547);
nor U1450 (N_1450,N_588,N_553);
nand U1451 (N_1451,N_302,N_251);
nand U1452 (N_1452,N_923,N_284);
xor U1453 (N_1453,N_907,N_513);
xnor U1454 (N_1454,N_346,N_807);
nor U1455 (N_1455,N_9,N_884);
nand U1456 (N_1456,N_641,N_125);
xor U1457 (N_1457,N_264,N_175);
or U1458 (N_1458,N_406,N_885);
nor U1459 (N_1459,N_218,N_167);
nand U1460 (N_1460,N_999,N_13);
nand U1461 (N_1461,N_644,N_150);
or U1462 (N_1462,N_303,N_794);
nor U1463 (N_1463,N_202,N_137);
and U1464 (N_1464,N_243,N_374);
nor U1465 (N_1465,N_917,N_85);
and U1466 (N_1466,N_978,N_69);
nor U1467 (N_1467,N_924,N_272);
and U1468 (N_1468,N_859,N_417);
or U1469 (N_1469,N_677,N_564);
nand U1470 (N_1470,N_236,N_172);
nand U1471 (N_1471,N_459,N_575);
nand U1472 (N_1472,N_276,N_372);
xor U1473 (N_1473,N_345,N_461);
xor U1474 (N_1474,N_905,N_698);
nand U1475 (N_1475,N_184,N_534);
nor U1476 (N_1476,N_922,N_378);
or U1477 (N_1477,N_256,N_686);
or U1478 (N_1478,N_799,N_948);
nor U1479 (N_1479,N_153,N_814);
and U1480 (N_1480,N_631,N_355);
nand U1481 (N_1481,N_457,N_624);
nor U1482 (N_1482,N_27,N_8);
xor U1483 (N_1483,N_731,N_467);
and U1484 (N_1484,N_787,N_119);
xnor U1485 (N_1485,N_382,N_858);
xor U1486 (N_1486,N_381,N_815);
nand U1487 (N_1487,N_629,N_227);
and U1488 (N_1488,N_298,N_307);
nor U1489 (N_1489,N_608,N_860);
nor U1490 (N_1490,N_290,N_367);
xnor U1491 (N_1491,N_933,N_750);
nor U1492 (N_1492,N_477,N_690);
and U1493 (N_1493,N_591,N_865);
nand U1494 (N_1494,N_711,N_105);
and U1495 (N_1495,N_684,N_143);
and U1496 (N_1496,N_118,N_525);
nand U1497 (N_1497,N_916,N_522);
nor U1498 (N_1498,N_344,N_33);
nand U1499 (N_1499,N_595,N_596);
or U1500 (N_1500,N_660,N_989);
or U1501 (N_1501,N_308,N_635);
nand U1502 (N_1502,N_671,N_773);
or U1503 (N_1503,N_266,N_480);
xor U1504 (N_1504,N_563,N_234);
or U1505 (N_1505,N_941,N_192);
nor U1506 (N_1506,N_414,N_672);
nor U1507 (N_1507,N_803,N_417);
nor U1508 (N_1508,N_165,N_907);
and U1509 (N_1509,N_508,N_395);
xor U1510 (N_1510,N_614,N_757);
or U1511 (N_1511,N_964,N_797);
nand U1512 (N_1512,N_816,N_282);
nand U1513 (N_1513,N_966,N_138);
or U1514 (N_1514,N_479,N_255);
nor U1515 (N_1515,N_401,N_883);
nand U1516 (N_1516,N_344,N_493);
and U1517 (N_1517,N_790,N_876);
or U1518 (N_1518,N_662,N_25);
nand U1519 (N_1519,N_295,N_157);
nor U1520 (N_1520,N_200,N_117);
nand U1521 (N_1521,N_445,N_124);
nor U1522 (N_1522,N_167,N_295);
xnor U1523 (N_1523,N_850,N_503);
or U1524 (N_1524,N_63,N_31);
or U1525 (N_1525,N_876,N_244);
nand U1526 (N_1526,N_188,N_532);
nand U1527 (N_1527,N_435,N_181);
and U1528 (N_1528,N_301,N_587);
and U1529 (N_1529,N_450,N_249);
xor U1530 (N_1530,N_503,N_651);
nand U1531 (N_1531,N_28,N_733);
xor U1532 (N_1532,N_491,N_535);
nor U1533 (N_1533,N_904,N_108);
and U1534 (N_1534,N_820,N_222);
xnor U1535 (N_1535,N_876,N_72);
and U1536 (N_1536,N_258,N_949);
and U1537 (N_1537,N_7,N_295);
nand U1538 (N_1538,N_566,N_870);
or U1539 (N_1539,N_791,N_140);
and U1540 (N_1540,N_537,N_25);
nor U1541 (N_1541,N_6,N_82);
nor U1542 (N_1542,N_227,N_165);
and U1543 (N_1543,N_28,N_689);
or U1544 (N_1544,N_727,N_691);
xor U1545 (N_1545,N_166,N_268);
and U1546 (N_1546,N_970,N_755);
or U1547 (N_1547,N_75,N_270);
xor U1548 (N_1548,N_392,N_337);
or U1549 (N_1549,N_534,N_574);
xnor U1550 (N_1550,N_831,N_606);
and U1551 (N_1551,N_649,N_271);
nand U1552 (N_1552,N_693,N_410);
xnor U1553 (N_1553,N_926,N_891);
xnor U1554 (N_1554,N_466,N_895);
nor U1555 (N_1555,N_570,N_385);
xnor U1556 (N_1556,N_860,N_803);
and U1557 (N_1557,N_486,N_69);
nor U1558 (N_1558,N_103,N_329);
nand U1559 (N_1559,N_92,N_363);
nor U1560 (N_1560,N_57,N_925);
or U1561 (N_1561,N_469,N_797);
xnor U1562 (N_1562,N_661,N_0);
xor U1563 (N_1563,N_610,N_117);
and U1564 (N_1564,N_45,N_957);
xor U1565 (N_1565,N_803,N_142);
and U1566 (N_1566,N_603,N_871);
xnor U1567 (N_1567,N_545,N_813);
and U1568 (N_1568,N_454,N_668);
nand U1569 (N_1569,N_783,N_916);
or U1570 (N_1570,N_585,N_705);
nand U1571 (N_1571,N_844,N_685);
nor U1572 (N_1572,N_994,N_799);
and U1573 (N_1573,N_628,N_108);
or U1574 (N_1574,N_368,N_311);
xor U1575 (N_1575,N_505,N_457);
nor U1576 (N_1576,N_210,N_271);
or U1577 (N_1577,N_284,N_483);
xor U1578 (N_1578,N_597,N_695);
nor U1579 (N_1579,N_375,N_486);
nand U1580 (N_1580,N_613,N_715);
or U1581 (N_1581,N_391,N_989);
xnor U1582 (N_1582,N_312,N_947);
xnor U1583 (N_1583,N_907,N_868);
nand U1584 (N_1584,N_800,N_470);
xnor U1585 (N_1585,N_549,N_597);
xor U1586 (N_1586,N_280,N_662);
nand U1587 (N_1587,N_907,N_171);
nand U1588 (N_1588,N_0,N_833);
xor U1589 (N_1589,N_796,N_551);
nor U1590 (N_1590,N_384,N_379);
and U1591 (N_1591,N_56,N_467);
or U1592 (N_1592,N_522,N_873);
and U1593 (N_1593,N_249,N_823);
nand U1594 (N_1594,N_768,N_433);
nor U1595 (N_1595,N_772,N_750);
or U1596 (N_1596,N_111,N_442);
xnor U1597 (N_1597,N_261,N_913);
xnor U1598 (N_1598,N_809,N_683);
or U1599 (N_1599,N_277,N_598);
nand U1600 (N_1600,N_645,N_476);
or U1601 (N_1601,N_831,N_712);
or U1602 (N_1602,N_766,N_329);
and U1603 (N_1603,N_957,N_602);
nand U1604 (N_1604,N_908,N_865);
nand U1605 (N_1605,N_151,N_452);
or U1606 (N_1606,N_140,N_203);
and U1607 (N_1607,N_431,N_552);
nor U1608 (N_1608,N_319,N_224);
or U1609 (N_1609,N_677,N_674);
or U1610 (N_1610,N_898,N_110);
or U1611 (N_1611,N_881,N_807);
nand U1612 (N_1612,N_381,N_433);
nor U1613 (N_1613,N_805,N_3);
xnor U1614 (N_1614,N_116,N_909);
xnor U1615 (N_1615,N_386,N_959);
nand U1616 (N_1616,N_624,N_839);
or U1617 (N_1617,N_333,N_823);
or U1618 (N_1618,N_869,N_593);
or U1619 (N_1619,N_548,N_293);
or U1620 (N_1620,N_504,N_258);
nand U1621 (N_1621,N_387,N_38);
xor U1622 (N_1622,N_186,N_760);
or U1623 (N_1623,N_217,N_265);
nand U1624 (N_1624,N_85,N_807);
xor U1625 (N_1625,N_90,N_98);
and U1626 (N_1626,N_27,N_616);
xor U1627 (N_1627,N_146,N_975);
and U1628 (N_1628,N_798,N_731);
nor U1629 (N_1629,N_85,N_967);
nor U1630 (N_1630,N_906,N_951);
and U1631 (N_1631,N_975,N_779);
nor U1632 (N_1632,N_296,N_26);
nor U1633 (N_1633,N_180,N_745);
or U1634 (N_1634,N_316,N_34);
nor U1635 (N_1635,N_726,N_644);
nor U1636 (N_1636,N_458,N_977);
nand U1637 (N_1637,N_671,N_41);
or U1638 (N_1638,N_213,N_517);
and U1639 (N_1639,N_636,N_869);
xor U1640 (N_1640,N_649,N_200);
xnor U1641 (N_1641,N_981,N_656);
and U1642 (N_1642,N_379,N_77);
or U1643 (N_1643,N_213,N_913);
nor U1644 (N_1644,N_182,N_335);
nor U1645 (N_1645,N_132,N_49);
or U1646 (N_1646,N_128,N_669);
and U1647 (N_1647,N_973,N_824);
nand U1648 (N_1648,N_701,N_449);
or U1649 (N_1649,N_497,N_307);
or U1650 (N_1650,N_681,N_527);
nand U1651 (N_1651,N_300,N_566);
and U1652 (N_1652,N_646,N_686);
xnor U1653 (N_1653,N_517,N_677);
nand U1654 (N_1654,N_376,N_131);
nand U1655 (N_1655,N_136,N_198);
or U1656 (N_1656,N_398,N_235);
nor U1657 (N_1657,N_800,N_699);
xnor U1658 (N_1658,N_512,N_92);
or U1659 (N_1659,N_989,N_105);
or U1660 (N_1660,N_419,N_126);
nor U1661 (N_1661,N_439,N_163);
nor U1662 (N_1662,N_264,N_598);
xnor U1663 (N_1663,N_787,N_473);
and U1664 (N_1664,N_629,N_432);
and U1665 (N_1665,N_571,N_308);
and U1666 (N_1666,N_754,N_981);
nor U1667 (N_1667,N_588,N_233);
or U1668 (N_1668,N_383,N_534);
or U1669 (N_1669,N_404,N_766);
nor U1670 (N_1670,N_783,N_950);
xor U1671 (N_1671,N_227,N_5);
xor U1672 (N_1672,N_305,N_40);
nor U1673 (N_1673,N_844,N_904);
and U1674 (N_1674,N_364,N_550);
nand U1675 (N_1675,N_426,N_966);
and U1676 (N_1676,N_287,N_943);
xnor U1677 (N_1677,N_47,N_134);
nor U1678 (N_1678,N_475,N_348);
nand U1679 (N_1679,N_715,N_704);
xnor U1680 (N_1680,N_348,N_716);
xnor U1681 (N_1681,N_899,N_169);
nand U1682 (N_1682,N_404,N_376);
xnor U1683 (N_1683,N_530,N_198);
nand U1684 (N_1684,N_280,N_240);
or U1685 (N_1685,N_153,N_823);
nand U1686 (N_1686,N_950,N_535);
nand U1687 (N_1687,N_426,N_251);
or U1688 (N_1688,N_202,N_652);
nand U1689 (N_1689,N_316,N_508);
nand U1690 (N_1690,N_30,N_503);
nor U1691 (N_1691,N_294,N_820);
nand U1692 (N_1692,N_815,N_501);
or U1693 (N_1693,N_98,N_215);
and U1694 (N_1694,N_601,N_941);
nor U1695 (N_1695,N_351,N_8);
xor U1696 (N_1696,N_528,N_90);
or U1697 (N_1697,N_832,N_147);
and U1698 (N_1698,N_968,N_50);
or U1699 (N_1699,N_45,N_280);
or U1700 (N_1700,N_24,N_115);
or U1701 (N_1701,N_963,N_18);
nand U1702 (N_1702,N_14,N_153);
and U1703 (N_1703,N_948,N_84);
nor U1704 (N_1704,N_984,N_625);
xor U1705 (N_1705,N_282,N_720);
nand U1706 (N_1706,N_31,N_258);
xor U1707 (N_1707,N_707,N_297);
nor U1708 (N_1708,N_580,N_782);
or U1709 (N_1709,N_959,N_759);
nor U1710 (N_1710,N_84,N_745);
or U1711 (N_1711,N_257,N_970);
nor U1712 (N_1712,N_342,N_815);
nand U1713 (N_1713,N_521,N_150);
nor U1714 (N_1714,N_142,N_564);
or U1715 (N_1715,N_402,N_418);
xnor U1716 (N_1716,N_856,N_764);
xnor U1717 (N_1717,N_224,N_256);
nand U1718 (N_1718,N_740,N_48);
nor U1719 (N_1719,N_90,N_278);
xor U1720 (N_1720,N_674,N_350);
nor U1721 (N_1721,N_884,N_15);
and U1722 (N_1722,N_248,N_32);
and U1723 (N_1723,N_354,N_334);
nand U1724 (N_1724,N_1,N_720);
nor U1725 (N_1725,N_792,N_878);
nand U1726 (N_1726,N_12,N_298);
and U1727 (N_1727,N_691,N_292);
and U1728 (N_1728,N_530,N_306);
and U1729 (N_1729,N_718,N_749);
nor U1730 (N_1730,N_448,N_602);
or U1731 (N_1731,N_708,N_797);
and U1732 (N_1732,N_538,N_107);
or U1733 (N_1733,N_16,N_642);
nor U1734 (N_1734,N_328,N_327);
nor U1735 (N_1735,N_672,N_828);
or U1736 (N_1736,N_954,N_592);
nor U1737 (N_1737,N_508,N_411);
xnor U1738 (N_1738,N_37,N_909);
or U1739 (N_1739,N_436,N_361);
or U1740 (N_1740,N_43,N_269);
nor U1741 (N_1741,N_936,N_745);
and U1742 (N_1742,N_568,N_264);
xor U1743 (N_1743,N_273,N_607);
or U1744 (N_1744,N_408,N_413);
or U1745 (N_1745,N_832,N_796);
nor U1746 (N_1746,N_317,N_418);
or U1747 (N_1747,N_738,N_758);
xnor U1748 (N_1748,N_889,N_998);
or U1749 (N_1749,N_571,N_23);
nor U1750 (N_1750,N_496,N_990);
and U1751 (N_1751,N_462,N_740);
xnor U1752 (N_1752,N_178,N_565);
nor U1753 (N_1753,N_310,N_909);
xor U1754 (N_1754,N_140,N_804);
and U1755 (N_1755,N_163,N_671);
xnor U1756 (N_1756,N_545,N_489);
or U1757 (N_1757,N_729,N_824);
xnor U1758 (N_1758,N_903,N_795);
nand U1759 (N_1759,N_7,N_802);
or U1760 (N_1760,N_319,N_776);
and U1761 (N_1761,N_175,N_749);
nand U1762 (N_1762,N_171,N_628);
and U1763 (N_1763,N_507,N_924);
and U1764 (N_1764,N_177,N_847);
nor U1765 (N_1765,N_923,N_717);
nor U1766 (N_1766,N_969,N_720);
nor U1767 (N_1767,N_270,N_665);
or U1768 (N_1768,N_875,N_855);
nand U1769 (N_1769,N_561,N_817);
and U1770 (N_1770,N_192,N_69);
nand U1771 (N_1771,N_530,N_648);
nor U1772 (N_1772,N_228,N_740);
and U1773 (N_1773,N_629,N_290);
nor U1774 (N_1774,N_619,N_613);
and U1775 (N_1775,N_455,N_289);
or U1776 (N_1776,N_978,N_821);
xnor U1777 (N_1777,N_242,N_182);
xor U1778 (N_1778,N_300,N_679);
or U1779 (N_1779,N_496,N_769);
nor U1780 (N_1780,N_388,N_192);
nor U1781 (N_1781,N_350,N_941);
nand U1782 (N_1782,N_85,N_926);
or U1783 (N_1783,N_208,N_32);
and U1784 (N_1784,N_137,N_615);
nand U1785 (N_1785,N_931,N_145);
and U1786 (N_1786,N_375,N_238);
nand U1787 (N_1787,N_197,N_89);
nor U1788 (N_1788,N_656,N_300);
xnor U1789 (N_1789,N_477,N_967);
nor U1790 (N_1790,N_365,N_53);
xor U1791 (N_1791,N_977,N_513);
nor U1792 (N_1792,N_836,N_353);
nand U1793 (N_1793,N_189,N_991);
xnor U1794 (N_1794,N_7,N_433);
nand U1795 (N_1795,N_100,N_77);
xnor U1796 (N_1796,N_485,N_130);
and U1797 (N_1797,N_740,N_963);
nor U1798 (N_1798,N_680,N_329);
and U1799 (N_1799,N_487,N_585);
nor U1800 (N_1800,N_838,N_84);
or U1801 (N_1801,N_784,N_673);
nor U1802 (N_1802,N_837,N_868);
and U1803 (N_1803,N_985,N_306);
or U1804 (N_1804,N_743,N_763);
or U1805 (N_1805,N_647,N_532);
nor U1806 (N_1806,N_726,N_942);
nand U1807 (N_1807,N_860,N_92);
and U1808 (N_1808,N_87,N_402);
xor U1809 (N_1809,N_322,N_241);
and U1810 (N_1810,N_211,N_135);
nor U1811 (N_1811,N_541,N_504);
and U1812 (N_1812,N_747,N_691);
xnor U1813 (N_1813,N_512,N_590);
nand U1814 (N_1814,N_298,N_574);
nor U1815 (N_1815,N_397,N_379);
and U1816 (N_1816,N_570,N_890);
nor U1817 (N_1817,N_41,N_467);
nor U1818 (N_1818,N_22,N_747);
and U1819 (N_1819,N_753,N_234);
xor U1820 (N_1820,N_172,N_304);
and U1821 (N_1821,N_395,N_384);
or U1822 (N_1822,N_33,N_629);
and U1823 (N_1823,N_813,N_918);
nor U1824 (N_1824,N_146,N_636);
nor U1825 (N_1825,N_496,N_666);
nand U1826 (N_1826,N_686,N_575);
xor U1827 (N_1827,N_69,N_738);
xor U1828 (N_1828,N_866,N_589);
nand U1829 (N_1829,N_432,N_880);
xnor U1830 (N_1830,N_346,N_44);
nor U1831 (N_1831,N_10,N_903);
xnor U1832 (N_1832,N_765,N_384);
or U1833 (N_1833,N_364,N_604);
xnor U1834 (N_1834,N_598,N_497);
or U1835 (N_1835,N_553,N_369);
nand U1836 (N_1836,N_532,N_816);
xnor U1837 (N_1837,N_205,N_398);
nand U1838 (N_1838,N_49,N_105);
and U1839 (N_1839,N_333,N_530);
or U1840 (N_1840,N_331,N_28);
and U1841 (N_1841,N_712,N_107);
xnor U1842 (N_1842,N_797,N_602);
or U1843 (N_1843,N_764,N_804);
or U1844 (N_1844,N_5,N_67);
and U1845 (N_1845,N_818,N_786);
nor U1846 (N_1846,N_536,N_366);
nand U1847 (N_1847,N_399,N_915);
nor U1848 (N_1848,N_368,N_440);
and U1849 (N_1849,N_472,N_551);
xnor U1850 (N_1850,N_110,N_492);
nand U1851 (N_1851,N_492,N_107);
and U1852 (N_1852,N_928,N_455);
nor U1853 (N_1853,N_977,N_667);
nand U1854 (N_1854,N_665,N_841);
nand U1855 (N_1855,N_724,N_324);
nor U1856 (N_1856,N_524,N_969);
nand U1857 (N_1857,N_207,N_648);
xor U1858 (N_1858,N_709,N_273);
nand U1859 (N_1859,N_551,N_7);
and U1860 (N_1860,N_357,N_689);
xor U1861 (N_1861,N_239,N_72);
and U1862 (N_1862,N_125,N_317);
and U1863 (N_1863,N_435,N_339);
or U1864 (N_1864,N_806,N_931);
nor U1865 (N_1865,N_489,N_311);
nand U1866 (N_1866,N_184,N_131);
and U1867 (N_1867,N_436,N_968);
and U1868 (N_1868,N_785,N_704);
nand U1869 (N_1869,N_857,N_925);
nor U1870 (N_1870,N_367,N_123);
nand U1871 (N_1871,N_552,N_59);
nand U1872 (N_1872,N_132,N_600);
nor U1873 (N_1873,N_537,N_583);
nor U1874 (N_1874,N_475,N_793);
nor U1875 (N_1875,N_227,N_192);
and U1876 (N_1876,N_294,N_206);
nor U1877 (N_1877,N_968,N_433);
nor U1878 (N_1878,N_840,N_844);
nand U1879 (N_1879,N_63,N_190);
or U1880 (N_1880,N_360,N_820);
and U1881 (N_1881,N_406,N_224);
nor U1882 (N_1882,N_334,N_289);
or U1883 (N_1883,N_30,N_116);
nand U1884 (N_1884,N_766,N_429);
nand U1885 (N_1885,N_417,N_948);
nor U1886 (N_1886,N_289,N_612);
or U1887 (N_1887,N_699,N_431);
nor U1888 (N_1888,N_625,N_513);
or U1889 (N_1889,N_107,N_618);
or U1890 (N_1890,N_764,N_862);
or U1891 (N_1891,N_378,N_903);
xor U1892 (N_1892,N_418,N_642);
xnor U1893 (N_1893,N_252,N_367);
xor U1894 (N_1894,N_469,N_465);
or U1895 (N_1895,N_755,N_668);
xor U1896 (N_1896,N_503,N_531);
nand U1897 (N_1897,N_174,N_863);
nand U1898 (N_1898,N_70,N_210);
xnor U1899 (N_1899,N_795,N_534);
and U1900 (N_1900,N_939,N_479);
nand U1901 (N_1901,N_524,N_933);
nor U1902 (N_1902,N_246,N_572);
nor U1903 (N_1903,N_348,N_754);
xnor U1904 (N_1904,N_824,N_880);
and U1905 (N_1905,N_428,N_568);
nor U1906 (N_1906,N_399,N_602);
nor U1907 (N_1907,N_633,N_707);
and U1908 (N_1908,N_109,N_997);
nand U1909 (N_1909,N_161,N_693);
or U1910 (N_1910,N_589,N_847);
nand U1911 (N_1911,N_687,N_3);
nand U1912 (N_1912,N_259,N_182);
nor U1913 (N_1913,N_322,N_672);
nand U1914 (N_1914,N_429,N_238);
nand U1915 (N_1915,N_172,N_598);
or U1916 (N_1916,N_511,N_422);
nor U1917 (N_1917,N_59,N_683);
xor U1918 (N_1918,N_979,N_151);
nor U1919 (N_1919,N_108,N_462);
or U1920 (N_1920,N_199,N_600);
xor U1921 (N_1921,N_444,N_694);
or U1922 (N_1922,N_299,N_284);
or U1923 (N_1923,N_116,N_961);
nand U1924 (N_1924,N_442,N_495);
nor U1925 (N_1925,N_773,N_384);
or U1926 (N_1926,N_503,N_190);
nand U1927 (N_1927,N_402,N_438);
or U1928 (N_1928,N_283,N_654);
nand U1929 (N_1929,N_610,N_827);
xor U1930 (N_1930,N_725,N_328);
nor U1931 (N_1931,N_514,N_620);
xnor U1932 (N_1932,N_187,N_279);
and U1933 (N_1933,N_362,N_916);
nor U1934 (N_1934,N_448,N_941);
and U1935 (N_1935,N_176,N_525);
and U1936 (N_1936,N_658,N_945);
nand U1937 (N_1937,N_396,N_154);
xor U1938 (N_1938,N_779,N_613);
xor U1939 (N_1939,N_741,N_369);
nor U1940 (N_1940,N_121,N_862);
xnor U1941 (N_1941,N_415,N_962);
and U1942 (N_1942,N_894,N_563);
xnor U1943 (N_1943,N_761,N_223);
or U1944 (N_1944,N_612,N_936);
xor U1945 (N_1945,N_276,N_47);
or U1946 (N_1946,N_923,N_897);
and U1947 (N_1947,N_552,N_220);
and U1948 (N_1948,N_293,N_969);
nand U1949 (N_1949,N_422,N_696);
or U1950 (N_1950,N_134,N_549);
nand U1951 (N_1951,N_571,N_46);
and U1952 (N_1952,N_289,N_151);
nand U1953 (N_1953,N_150,N_279);
or U1954 (N_1954,N_772,N_147);
nor U1955 (N_1955,N_762,N_460);
and U1956 (N_1956,N_568,N_769);
and U1957 (N_1957,N_48,N_507);
nand U1958 (N_1958,N_602,N_418);
xor U1959 (N_1959,N_883,N_91);
or U1960 (N_1960,N_795,N_7);
xnor U1961 (N_1961,N_745,N_228);
nor U1962 (N_1962,N_673,N_787);
nor U1963 (N_1963,N_130,N_423);
nor U1964 (N_1964,N_337,N_816);
nand U1965 (N_1965,N_927,N_790);
and U1966 (N_1966,N_425,N_483);
or U1967 (N_1967,N_416,N_758);
nor U1968 (N_1968,N_673,N_822);
nor U1969 (N_1969,N_607,N_216);
and U1970 (N_1970,N_476,N_221);
xor U1971 (N_1971,N_807,N_284);
xnor U1972 (N_1972,N_874,N_23);
xnor U1973 (N_1973,N_294,N_72);
nor U1974 (N_1974,N_895,N_727);
or U1975 (N_1975,N_369,N_895);
nor U1976 (N_1976,N_245,N_648);
nor U1977 (N_1977,N_514,N_117);
xnor U1978 (N_1978,N_874,N_558);
nand U1979 (N_1979,N_658,N_828);
nor U1980 (N_1980,N_64,N_632);
nor U1981 (N_1981,N_179,N_746);
nand U1982 (N_1982,N_972,N_396);
and U1983 (N_1983,N_760,N_706);
nor U1984 (N_1984,N_104,N_256);
and U1985 (N_1985,N_609,N_25);
or U1986 (N_1986,N_667,N_653);
or U1987 (N_1987,N_795,N_135);
or U1988 (N_1988,N_915,N_845);
and U1989 (N_1989,N_914,N_890);
xnor U1990 (N_1990,N_817,N_134);
xor U1991 (N_1991,N_57,N_580);
nor U1992 (N_1992,N_516,N_343);
and U1993 (N_1993,N_498,N_217);
nor U1994 (N_1994,N_226,N_342);
and U1995 (N_1995,N_462,N_467);
nor U1996 (N_1996,N_837,N_6);
xor U1997 (N_1997,N_381,N_688);
nor U1998 (N_1998,N_886,N_469);
nor U1999 (N_1999,N_299,N_608);
and U2000 (N_2000,N_1416,N_1493);
or U2001 (N_2001,N_1239,N_1485);
or U2002 (N_2002,N_1055,N_1097);
xor U2003 (N_2003,N_1506,N_1192);
or U2004 (N_2004,N_1842,N_1821);
nand U2005 (N_2005,N_1965,N_1788);
xor U2006 (N_2006,N_1618,N_1566);
nand U2007 (N_2007,N_1004,N_1305);
nand U2008 (N_2008,N_1530,N_1881);
and U2009 (N_2009,N_1740,N_1407);
xnor U2010 (N_2010,N_1406,N_1456);
nor U2011 (N_2011,N_1068,N_1054);
nand U2012 (N_2012,N_1830,N_1536);
and U2013 (N_2013,N_1392,N_1575);
or U2014 (N_2014,N_1016,N_1169);
xnor U2015 (N_2015,N_1621,N_1430);
or U2016 (N_2016,N_1084,N_1771);
and U2017 (N_2017,N_1252,N_1633);
xor U2018 (N_2018,N_1237,N_1165);
nor U2019 (N_2019,N_1547,N_1543);
and U2020 (N_2020,N_1094,N_1580);
nand U2021 (N_2021,N_1974,N_1149);
or U2022 (N_2022,N_1310,N_1177);
nor U2023 (N_2023,N_1729,N_1394);
and U2024 (N_2024,N_1675,N_1926);
xnor U2025 (N_2025,N_1998,N_1155);
nand U2026 (N_2026,N_1044,N_1510);
and U2027 (N_2027,N_1541,N_1253);
xor U2028 (N_2028,N_1997,N_1971);
nor U2029 (N_2029,N_1369,N_1791);
xnor U2030 (N_2030,N_1098,N_1442);
xnor U2031 (N_2031,N_1495,N_1435);
and U2032 (N_2032,N_1304,N_1377);
or U2033 (N_2033,N_1993,N_1433);
and U2034 (N_2034,N_1587,N_1714);
nand U2035 (N_2035,N_1003,N_1031);
nand U2036 (N_2036,N_1801,N_1307);
xor U2037 (N_2037,N_1662,N_1123);
nand U2038 (N_2038,N_1522,N_1851);
and U2039 (N_2039,N_1035,N_1915);
or U2040 (N_2040,N_1591,N_1319);
nand U2041 (N_2041,N_1255,N_1475);
or U2042 (N_2042,N_1298,N_1519);
nand U2043 (N_2043,N_1563,N_1589);
or U2044 (N_2044,N_1507,N_1374);
nand U2045 (N_2045,N_1057,N_1183);
nor U2046 (N_2046,N_1725,N_1758);
nand U2047 (N_2047,N_1138,N_1599);
nor U2048 (N_2048,N_1635,N_1898);
xnor U2049 (N_2049,N_1620,N_1478);
and U2050 (N_2050,N_1835,N_1415);
xnor U2051 (N_2051,N_1204,N_1963);
nand U2052 (N_2052,N_1611,N_1245);
nand U2053 (N_2053,N_1903,N_1362);
xor U2054 (N_2054,N_1875,N_1989);
nand U2055 (N_2055,N_1007,N_1327);
and U2056 (N_2056,N_1778,N_1048);
and U2057 (N_2057,N_1349,N_1460);
nand U2058 (N_2058,N_1070,N_1689);
and U2059 (N_2059,N_1405,N_1013);
nor U2060 (N_2060,N_1655,N_1968);
xor U2061 (N_2061,N_1562,N_1122);
nor U2062 (N_2062,N_1347,N_1303);
or U2063 (N_2063,N_1592,N_1212);
and U2064 (N_2064,N_1657,N_1700);
nand U2065 (N_2065,N_1900,N_1776);
and U2066 (N_2066,N_1756,N_1353);
and U2067 (N_2067,N_1453,N_1019);
nand U2068 (N_2068,N_1140,N_1271);
xor U2069 (N_2069,N_1528,N_1373);
nor U2070 (N_2070,N_1560,N_1841);
nor U2071 (N_2071,N_1499,N_1557);
or U2072 (N_2072,N_1201,N_1170);
or U2073 (N_2073,N_1315,N_1627);
or U2074 (N_2074,N_1500,N_1059);
or U2075 (N_2075,N_1247,N_1262);
xor U2076 (N_2076,N_1669,N_1189);
xnor U2077 (N_2077,N_1833,N_1371);
xor U2078 (N_2078,N_1643,N_1737);
or U2079 (N_2079,N_1784,N_1261);
or U2080 (N_2080,N_1780,N_1660);
and U2081 (N_2081,N_1947,N_1082);
xnor U2082 (N_2082,N_1981,N_1857);
and U2083 (N_2083,N_1930,N_1151);
and U2084 (N_2084,N_1697,N_1158);
and U2085 (N_2085,N_1559,N_1814);
and U2086 (N_2086,N_1739,N_1424);
xnor U2087 (N_2087,N_1918,N_1847);
xnor U2088 (N_2088,N_1622,N_1120);
xnor U2089 (N_2089,N_1205,N_1412);
or U2090 (N_2090,N_1157,N_1939);
or U2091 (N_2091,N_1295,N_1532);
or U2092 (N_2092,N_1064,N_1273);
xor U2093 (N_2093,N_1086,N_1066);
or U2094 (N_2094,N_1916,N_1326);
or U2095 (N_2095,N_1039,N_1108);
or U2096 (N_2096,N_1889,N_1703);
or U2097 (N_2097,N_1710,N_1984);
nor U2098 (N_2098,N_1376,N_1584);
or U2099 (N_2099,N_1713,N_1921);
nor U2100 (N_2100,N_1036,N_1886);
and U2101 (N_2101,N_1095,N_1153);
nand U2102 (N_2102,N_1985,N_1053);
or U2103 (N_2103,N_1463,N_1490);
xor U2104 (N_2104,N_1839,N_1173);
nand U2105 (N_2105,N_1292,N_1929);
and U2106 (N_2106,N_1227,N_1366);
or U2107 (N_2107,N_1508,N_1001);
xor U2108 (N_2108,N_1026,N_1146);
nand U2109 (N_2109,N_1300,N_1755);
nand U2110 (N_2110,N_1504,N_1159);
nand U2111 (N_2111,N_1800,N_1333);
xnor U2112 (N_2112,N_1017,N_1029);
nor U2113 (N_2113,N_1777,N_1786);
or U2114 (N_2114,N_1494,N_1783);
and U2115 (N_2115,N_1595,N_1753);
nand U2116 (N_2116,N_1815,N_1678);
xor U2117 (N_2117,N_1311,N_1822);
or U2118 (N_2118,N_1744,N_1583);
xor U2119 (N_2119,N_1260,N_1395);
nand U2120 (N_2120,N_1705,N_1887);
xor U2121 (N_2121,N_1874,N_1264);
nor U2122 (N_2122,N_1040,N_1280);
and U2123 (N_2123,N_1859,N_1397);
or U2124 (N_2124,N_1336,N_1950);
xor U2125 (N_2125,N_1518,N_1888);
or U2126 (N_2126,N_1243,N_1846);
and U2127 (N_2127,N_1897,N_1542);
nor U2128 (N_2128,N_1109,N_1308);
or U2129 (N_2129,N_1883,N_1820);
or U2130 (N_2130,N_1905,N_1471);
and U2131 (N_2131,N_1681,N_1992);
xor U2132 (N_2132,N_1079,N_1661);
nand U2133 (N_2133,N_1287,N_1021);
xor U2134 (N_2134,N_1706,N_1938);
nor U2135 (N_2135,N_1578,N_1860);
and U2136 (N_2136,N_1286,N_1512);
xor U2137 (N_2137,N_1167,N_1411);
nand U2138 (N_2138,N_1297,N_1025);
nor U2139 (N_2139,N_1870,N_1221);
xor U2140 (N_2140,N_1537,N_1607);
nand U2141 (N_2141,N_1955,N_1624);
and U2142 (N_2142,N_1524,N_1346);
or U2143 (N_2143,N_1555,N_1717);
nand U2144 (N_2144,N_1638,N_1680);
and U2145 (N_2145,N_1919,N_1914);
nand U2146 (N_2146,N_1840,N_1999);
nor U2147 (N_2147,N_1861,N_1266);
nand U2148 (N_2148,N_1663,N_1853);
xor U2149 (N_2149,N_1795,N_1879);
or U2150 (N_2150,N_1722,N_1849);
nand U2151 (N_2151,N_1571,N_1693);
nand U2152 (N_2152,N_1630,N_1350);
xor U2153 (N_2153,N_1804,N_1650);
nor U2154 (N_2154,N_1690,N_1610);
and U2155 (N_2155,N_1937,N_1338);
nand U2156 (N_2156,N_1639,N_1642);
and U2157 (N_2157,N_1698,N_1579);
and U2158 (N_2158,N_1958,N_1793);
xnor U2159 (N_2159,N_1182,N_1345);
or U2160 (N_2160,N_1552,N_1249);
xnor U2161 (N_2161,N_1976,N_1145);
xnor U2162 (N_2162,N_1278,N_1439);
or U2163 (N_2163,N_1360,N_1332);
xor U2164 (N_2164,N_1535,N_1426);
xnor U2165 (N_2165,N_1190,N_1389);
nand U2166 (N_2166,N_1275,N_1090);
nor U2167 (N_2167,N_1745,N_1634);
nor U2168 (N_2168,N_1175,N_1802);
and U2169 (N_2169,N_1723,N_1083);
xor U2170 (N_2170,N_1144,N_1343);
nor U2171 (N_2171,N_1796,N_1482);
xnor U2172 (N_2172,N_1012,N_1730);
or U2173 (N_2173,N_1604,N_1534);
xor U2174 (N_2174,N_1142,N_1114);
nor U2175 (N_2175,N_1850,N_1826);
and U2176 (N_2176,N_1464,N_1445);
and U2177 (N_2177,N_1402,N_1948);
xnor U2178 (N_2178,N_1166,N_1876);
and U2179 (N_2179,N_1076,N_1092);
nand U2180 (N_2180,N_1827,N_1299);
xor U2181 (N_2181,N_1113,N_1588);
xor U2182 (N_2182,N_1441,N_1837);
and U2183 (N_2183,N_1431,N_1609);
or U2184 (N_2184,N_1746,N_1052);
nand U2185 (N_2185,N_1276,N_1051);
nand U2186 (N_2186,N_1207,N_1427);
xnor U2187 (N_2187,N_1891,N_1174);
nand U2188 (N_2188,N_1654,N_1568);
xor U2189 (N_2189,N_1263,N_1787);
xor U2190 (N_2190,N_1523,N_1188);
or U2191 (N_2191,N_1231,N_1503);
or U2192 (N_2192,N_1909,N_1488);
nor U2193 (N_2193,N_1359,N_1752);
xnor U2194 (N_2194,N_1226,N_1404);
nand U2195 (N_2195,N_1421,N_1790);
and U2196 (N_2196,N_1973,N_1131);
nand U2197 (N_2197,N_1284,N_1996);
or U2198 (N_2198,N_1472,N_1325);
and U2199 (N_2199,N_1553,N_1080);
xnor U2200 (N_2200,N_1682,N_1372);
nand U2201 (N_2201,N_1110,N_1664);
or U2202 (N_2202,N_1761,N_1465);
nand U2203 (N_2203,N_1202,N_1838);
nor U2204 (N_2204,N_1133,N_1486);
and U2205 (N_2205,N_1648,N_1436);
nor U2206 (N_2206,N_1018,N_1000);
and U2207 (N_2207,N_1546,N_1674);
or U2208 (N_2208,N_1818,N_1330);
nand U2209 (N_2209,N_1124,N_1767);
xor U2210 (N_2210,N_1961,N_1569);
and U2211 (N_2211,N_1843,N_1550);
xnor U2212 (N_2212,N_1210,N_1008);
nor U2213 (N_2213,N_1731,N_1922);
xor U2214 (N_2214,N_1715,N_1208);
and U2215 (N_2215,N_1342,N_1880);
nor U2216 (N_2216,N_1854,N_1257);
and U2217 (N_2217,N_1625,N_1775);
and U2218 (N_2218,N_1565,N_1483);
nand U2219 (N_2219,N_1816,N_1699);
xor U2220 (N_2220,N_1198,N_1015);
nand U2221 (N_2221,N_1251,N_1712);
nand U2222 (N_2222,N_1873,N_1458);
or U2223 (N_2223,N_1214,N_1509);
xor U2224 (N_2224,N_1281,N_1502);
nor U2225 (N_2225,N_1331,N_1196);
xor U2226 (N_2226,N_1932,N_1195);
xor U2227 (N_2227,N_1228,N_1668);
or U2228 (N_2228,N_1960,N_1869);
and U2229 (N_2229,N_1732,N_1748);
nand U2230 (N_2230,N_1238,N_1005);
nor U2231 (N_2231,N_1893,N_1945);
nand U2232 (N_2232,N_1259,N_1455);
nand U2233 (N_2233,N_1213,N_1708);
nand U2234 (N_2234,N_1477,N_1152);
or U2235 (N_2235,N_1267,N_1106);
nand U2236 (N_2236,N_1967,N_1282);
nand U2237 (N_2237,N_1056,N_1832);
or U2238 (N_2238,N_1254,N_1063);
and U2239 (N_2239,N_1696,N_1768);
nor U2240 (N_2240,N_1823,N_1970);
nor U2241 (N_2241,N_1258,N_1378);
or U2242 (N_2242,N_1387,N_1692);
xor U2243 (N_2243,N_1549,N_1707);
nand U2244 (N_2244,N_1572,N_1679);
nand U2245 (N_2245,N_1551,N_1983);
xor U2246 (N_2246,N_1619,N_1803);
and U2247 (N_2247,N_1529,N_1577);
or U2248 (N_2248,N_1812,N_1323);
xnor U2249 (N_2249,N_1521,N_1806);
nor U2250 (N_2250,N_1002,N_1462);
or U2251 (N_2251,N_1250,N_1913);
nor U2252 (N_2252,N_1694,N_1593);
and U2253 (N_2253,N_1720,N_1269);
nor U2254 (N_2254,N_1774,N_1043);
nor U2255 (N_2255,N_1450,N_1337);
or U2256 (N_2256,N_1162,N_1759);
nand U2257 (N_2257,N_1199,N_1209);
xor U2258 (N_2258,N_1576,N_1398);
and U2259 (N_2259,N_1107,N_1096);
or U2260 (N_2260,N_1322,N_1115);
nor U2261 (N_2261,N_1469,N_1283);
nor U2262 (N_2262,N_1651,N_1561);
nand U2263 (N_2263,N_1573,N_1949);
or U2264 (N_2264,N_1491,N_1187);
nand U2265 (N_2265,N_1071,N_1101);
and U2266 (N_2266,N_1061,N_1119);
xnor U2267 (N_2267,N_1799,N_1487);
and U2268 (N_2268,N_1234,N_1480);
nand U2269 (N_2269,N_1733,N_1367);
or U2270 (N_2270,N_1836,N_1390);
xor U2271 (N_2271,N_1074,N_1809);
nor U2272 (N_2272,N_1341,N_1652);
or U2273 (N_2273,N_1912,N_1470);
or U2274 (N_2274,N_1316,N_1320);
nand U2275 (N_2275,N_1134,N_1721);
or U2276 (N_2276,N_1088,N_1193);
xor U2277 (N_2277,N_1928,N_1220);
or U2278 (N_2278,N_1099,N_1348);
or U2279 (N_2279,N_1747,N_1824);
nor U2280 (N_2280,N_1130,N_1764);
xnor U2281 (N_2281,N_1798,N_1329);
and U2282 (N_2282,N_1454,N_1409);
xor U2283 (N_2283,N_1856,N_1093);
and U2284 (N_2284,N_1184,N_1489);
xor U2285 (N_2285,N_1978,N_1894);
and U2286 (N_2286,N_1538,N_1075);
and U2287 (N_2287,N_1147,N_1139);
nor U2288 (N_2288,N_1515,N_1218);
nor U2289 (N_2289,N_1709,N_1590);
xnor U2290 (N_2290,N_1539,N_1011);
nor U2291 (N_2291,N_1864,N_1437);
xor U2292 (N_2292,N_1296,N_1137);
or U2293 (N_2293,N_1024,N_1741);
or U2294 (N_2294,N_1381,N_1511);
nor U2295 (N_2295,N_1461,N_1265);
nor U2296 (N_2296,N_1628,N_1194);
or U2297 (N_2297,N_1449,N_1884);
and U2298 (N_2298,N_1046,N_1224);
and U2299 (N_2299,N_1766,N_1363);
nor U2300 (N_2300,N_1423,N_1616);
xor U2301 (N_2301,N_1863,N_1907);
nand U2302 (N_2302,N_1656,N_1819);
or U2303 (N_2303,N_1274,N_1288);
xnor U2304 (N_2304,N_1779,N_1375);
nand U2305 (N_2305,N_1042,N_1641);
or U2306 (N_2306,N_1531,N_1314);
nor U2307 (N_2307,N_1126,N_1762);
and U2308 (N_2308,N_1111,N_1977);
nand U2309 (N_2309,N_1041,N_1647);
xnor U2310 (N_2310,N_1339,N_1940);
nor U2311 (N_2311,N_1476,N_1871);
xor U2312 (N_2312,N_1022,N_1223);
or U2313 (N_2313,N_1865,N_1558);
or U2314 (N_2314,N_1936,N_1601);
xor U2315 (N_2315,N_1062,N_1726);
and U2316 (N_2316,N_1760,N_1200);
nand U2317 (N_2317,N_1023,N_1959);
nand U2318 (N_2318,N_1391,N_1902);
nand U2319 (N_2319,N_1517,N_1232);
and U2320 (N_2320,N_1683,N_1279);
nand U2321 (N_2321,N_1581,N_1073);
or U2322 (N_2322,N_1781,N_1605);
nor U2323 (N_2323,N_1540,N_1516);
xnor U2324 (N_2324,N_1751,N_1085);
and U2325 (N_2325,N_1216,N_1782);
nand U2326 (N_2326,N_1688,N_1217);
or U2327 (N_2327,N_1178,N_1340);
nand U2328 (N_2328,N_1154,N_1117);
xnor U2329 (N_2329,N_1701,N_1136);
nand U2330 (N_2330,N_1161,N_1105);
or U2331 (N_2331,N_1582,N_1908);
nand U2332 (N_2332,N_1100,N_1666);
xnor U2333 (N_2333,N_1727,N_1990);
or U2334 (N_2334,N_1614,N_1617);
nand U2335 (N_2335,N_1236,N_1684);
and U2336 (N_2336,N_1289,N_1087);
and U2337 (N_2337,N_1736,N_1129);
nand U2338 (N_2338,N_1225,N_1479);
or U2339 (N_2339,N_1933,N_1246);
and U2340 (N_2340,N_1986,N_1355);
and U2341 (N_2341,N_1185,N_1241);
xnor U2342 (N_2342,N_1829,N_1270);
and U2343 (N_2343,N_1396,N_1385);
or U2344 (N_2344,N_1808,N_1148);
nor U2345 (N_2345,N_1277,N_1498);
nor U2346 (N_2346,N_1899,N_1743);
xor U2347 (N_2347,N_1452,N_1334);
xnor U2348 (N_2348,N_1368,N_1230);
and U2349 (N_2349,N_1203,N_1934);
nor U2350 (N_2350,N_1403,N_1248);
nand U2351 (N_2351,N_1112,N_1716);
or U2352 (N_2352,N_1527,N_1969);
and U2353 (N_2353,N_1393,N_1691);
nor U2354 (N_2354,N_1467,N_1451);
xor U2355 (N_2355,N_1567,N_1554);
or U2356 (N_2356,N_1176,N_1980);
nor U2357 (N_2357,N_1687,N_1670);
and U2358 (N_2358,N_1006,N_1636);
nor U2359 (N_2359,N_1388,N_1150);
xor U2360 (N_2360,N_1291,N_1877);
xnor U2361 (N_2361,N_1078,N_1895);
and U2362 (N_2362,N_1659,N_1302);
nand U2363 (N_2363,N_1324,N_1724);
nor U2364 (N_2364,N_1233,N_1769);
xnor U2365 (N_2365,N_1944,N_1585);
nand U2366 (N_2366,N_1370,N_1676);
or U2367 (N_2367,N_1598,N_1594);
or U2368 (N_2368,N_1020,N_1408);
nor U2369 (N_2369,N_1972,N_1317);
xor U2370 (N_2370,N_1734,N_1364);
or U2371 (N_2371,N_1906,N_1718);
or U2372 (N_2372,N_1501,N_1410);
or U2373 (N_2373,N_1457,N_1352);
xor U2374 (N_2374,N_1030,N_1418);
xor U2375 (N_2375,N_1321,N_1520);
nand U2376 (N_2376,N_1077,N_1866);
nor U2377 (N_2377,N_1135,N_1091);
xnor U2378 (N_2378,N_1072,N_1496);
nor U2379 (N_2379,N_1982,N_1514);
or U2380 (N_2380,N_1586,N_1844);
or U2381 (N_2381,N_1757,N_1702);
and U2382 (N_2382,N_1831,N_1941);
nor U2383 (N_2383,N_1602,N_1646);
xnor U2384 (N_2384,N_1952,N_1285);
and U2385 (N_2385,N_1414,N_1644);
nor U2386 (N_2386,N_1067,N_1991);
and U2387 (N_2387,N_1448,N_1867);
xnor U2388 (N_2388,N_1600,N_1645);
xnor U2389 (N_2389,N_1789,N_1313);
and U2390 (N_2390,N_1294,N_1596);
nand U2391 (N_2391,N_1637,N_1141);
nor U2392 (N_2392,N_1711,N_1034);
and U2393 (N_2393,N_1825,N_1956);
or U2394 (N_2394,N_1738,N_1492);
nor U2395 (N_2395,N_1807,N_1828);
and U2396 (N_2396,N_1413,N_1419);
nor U2397 (N_2397,N_1268,N_1810);
nor U2398 (N_2398,N_1858,N_1658);
xnor U2399 (N_2399,N_1354,N_1058);
or U2400 (N_2400,N_1817,N_1719);
xnor U2401 (N_2401,N_1910,N_1047);
nor U2402 (N_2402,N_1763,N_1923);
or U2403 (N_2403,N_1770,N_1878);
xor U2404 (N_2404,N_1848,N_1060);
or U2405 (N_2405,N_1222,N_1672);
nor U2406 (N_2406,N_1966,N_1446);
and U2407 (N_2407,N_1612,N_1631);
nor U2408 (N_2408,N_1069,N_1027);
or U2409 (N_2409,N_1163,N_1386);
nand U2410 (N_2410,N_1191,N_1197);
nand U2411 (N_2411,N_1365,N_1885);
and U2412 (N_2412,N_1953,N_1862);
nand U2413 (N_2413,N_1422,N_1811);
or U2414 (N_2414,N_1420,N_1957);
or U2415 (N_2415,N_1975,N_1399);
nor U2416 (N_2416,N_1132,N_1868);
nor U2417 (N_2417,N_1328,N_1765);
and U2418 (N_2418,N_1242,N_1855);
or U2419 (N_2419,N_1384,N_1168);
or U2420 (N_2420,N_1235,N_1946);
xnor U2421 (N_2421,N_1852,N_1603);
nor U2422 (N_2422,N_1104,N_1361);
nor U2423 (N_2423,N_1290,N_1116);
xnor U2424 (N_2424,N_1009,N_1049);
nand U2425 (N_2425,N_1673,N_1935);
and U2426 (N_2426,N_1211,N_1028);
nand U2427 (N_2427,N_1608,N_1749);
nor U2428 (N_2428,N_1033,N_1964);
and U2429 (N_2429,N_1671,N_1813);
and U2430 (N_2430,N_1089,N_1979);
or U2431 (N_2431,N_1653,N_1309);
nand U2432 (N_2432,N_1497,N_1545);
and U2433 (N_2433,N_1038,N_1570);
nand U2434 (N_2434,N_1754,N_1574);
xor U2435 (N_2435,N_1065,N_1306);
xnor U2436 (N_2436,N_1613,N_1351);
nor U2437 (N_2437,N_1911,N_1925);
nor U2438 (N_2438,N_1102,N_1901);
nor U2439 (N_2439,N_1443,N_1256);
or U2440 (N_2440,N_1335,N_1677);
xnor U2441 (N_2441,N_1121,N_1440);
or U2442 (N_2442,N_1244,N_1417);
xor U2443 (N_2443,N_1037,N_1081);
and U2444 (N_2444,N_1143,N_1533);
and U2445 (N_2445,N_1206,N_1942);
or U2446 (N_2446,N_1240,N_1229);
nor U2447 (N_2447,N_1954,N_1181);
nor U2448 (N_2448,N_1103,N_1665);
nor U2449 (N_2449,N_1344,N_1513);
nand U2450 (N_2450,N_1773,N_1400);
nand U2451 (N_2451,N_1272,N_1606);
or U2452 (N_2452,N_1380,N_1526);
xor U2453 (N_2453,N_1805,N_1032);
and U2454 (N_2454,N_1357,N_1615);
xnor U2455 (N_2455,N_1164,N_1797);
xor U2456 (N_2456,N_1125,N_1728);
and U2457 (N_2457,N_1994,N_1704);
nor U2458 (N_2458,N_1924,N_1735);
and U2459 (N_2459,N_1312,N_1010);
nand U2460 (N_2460,N_1474,N_1951);
xnor U2461 (N_2461,N_1525,N_1318);
xor U2462 (N_2462,N_1872,N_1548);
or U2463 (N_2463,N_1379,N_1127);
and U2464 (N_2464,N_1995,N_1626);
xor U2465 (N_2465,N_1383,N_1050);
and U2466 (N_2466,N_1564,N_1505);
and U2467 (N_2467,N_1425,N_1845);
and U2468 (N_2468,N_1118,N_1927);
nor U2469 (N_2469,N_1401,N_1962);
and U2470 (N_2470,N_1186,N_1667);
nand U2471 (N_2471,N_1356,N_1160);
or U2472 (N_2472,N_1171,N_1447);
xor U2473 (N_2473,N_1484,N_1597);
and U2474 (N_2474,N_1468,N_1179);
xor U2475 (N_2475,N_1215,N_1632);
nand U2476 (N_2476,N_1785,N_1649);
and U2477 (N_2477,N_1180,N_1988);
and U2478 (N_2478,N_1834,N_1014);
nor U2479 (N_2479,N_1750,N_1890);
nand U2480 (N_2480,N_1473,N_1428);
nor U2481 (N_2481,N_1943,N_1987);
xor U2482 (N_2482,N_1432,N_1544);
nor U2483 (N_2483,N_1466,N_1792);
or U2484 (N_2484,N_1429,N_1358);
or U2485 (N_2485,N_1434,N_1896);
or U2486 (N_2486,N_1459,N_1882);
nor U2487 (N_2487,N_1920,N_1629);
xor U2488 (N_2488,N_1444,N_1301);
or U2489 (N_2489,N_1904,N_1382);
and U2490 (N_2490,N_1172,N_1128);
or U2491 (N_2491,N_1794,N_1640);
xnor U2492 (N_2492,N_1892,N_1686);
or U2493 (N_2493,N_1045,N_1742);
nor U2494 (N_2494,N_1556,N_1219);
nand U2495 (N_2495,N_1931,N_1772);
nand U2496 (N_2496,N_1623,N_1293);
or U2497 (N_2497,N_1917,N_1685);
and U2498 (N_2498,N_1156,N_1438);
nor U2499 (N_2499,N_1695,N_1481);
xor U2500 (N_2500,N_1291,N_1300);
nor U2501 (N_2501,N_1067,N_1984);
nor U2502 (N_2502,N_1167,N_1059);
xnor U2503 (N_2503,N_1426,N_1442);
or U2504 (N_2504,N_1752,N_1575);
nor U2505 (N_2505,N_1801,N_1560);
and U2506 (N_2506,N_1107,N_1412);
xor U2507 (N_2507,N_1356,N_1872);
or U2508 (N_2508,N_1190,N_1755);
xor U2509 (N_2509,N_1761,N_1353);
and U2510 (N_2510,N_1220,N_1529);
or U2511 (N_2511,N_1359,N_1891);
and U2512 (N_2512,N_1637,N_1621);
or U2513 (N_2513,N_1239,N_1360);
and U2514 (N_2514,N_1415,N_1052);
or U2515 (N_2515,N_1395,N_1178);
nor U2516 (N_2516,N_1998,N_1434);
and U2517 (N_2517,N_1683,N_1742);
and U2518 (N_2518,N_1629,N_1359);
xor U2519 (N_2519,N_1606,N_1004);
and U2520 (N_2520,N_1062,N_1346);
and U2521 (N_2521,N_1918,N_1239);
and U2522 (N_2522,N_1317,N_1888);
and U2523 (N_2523,N_1468,N_1338);
nor U2524 (N_2524,N_1244,N_1441);
and U2525 (N_2525,N_1671,N_1454);
nor U2526 (N_2526,N_1887,N_1558);
or U2527 (N_2527,N_1333,N_1080);
xor U2528 (N_2528,N_1510,N_1407);
xor U2529 (N_2529,N_1717,N_1204);
and U2530 (N_2530,N_1466,N_1455);
nand U2531 (N_2531,N_1880,N_1701);
nor U2532 (N_2532,N_1119,N_1260);
or U2533 (N_2533,N_1667,N_1873);
or U2534 (N_2534,N_1347,N_1761);
xor U2535 (N_2535,N_1751,N_1449);
nand U2536 (N_2536,N_1499,N_1597);
and U2537 (N_2537,N_1380,N_1833);
and U2538 (N_2538,N_1569,N_1660);
and U2539 (N_2539,N_1411,N_1807);
and U2540 (N_2540,N_1388,N_1929);
nand U2541 (N_2541,N_1084,N_1171);
nand U2542 (N_2542,N_1269,N_1689);
or U2543 (N_2543,N_1257,N_1302);
nand U2544 (N_2544,N_1444,N_1373);
and U2545 (N_2545,N_1367,N_1323);
xor U2546 (N_2546,N_1878,N_1257);
and U2547 (N_2547,N_1934,N_1161);
nor U2548 (N_2548,N_1980,N_1255);
xnor U2549 (N_2549,N_1198,N_1533);
nor U2550 (N_2550,N_1895,N_1916);
xnor U2551 (N_2551,N_1723,N_1064);
xnor U2552 (N_2552,N_1113,N_1228);
xor U2553 (N_2553,N_1044,N_1641);
and U2554 (N_2554,N_1221,N_1283);
nand U2555 (N_2555,N_1753,N_1040);
or U2556 (N_2556,N_1964,N_1542);
and U2557 (N_2557,N_1509,N_1542);
nor U2558 (N_2558,N_1350,N_1493);
or U2559 (N_2559,N_1668,N_1301);
or U2560 (N_2560,N_1496,N_1111);
or U2561 (N_2561,N_1208,N_1429);
and U2562 (N_2562,N_1306,N_1809);
nor U2563 (N_2563,N_1756,N_1029);
and U2564 (N_2564,N_1000,N_1162);
nand U2565 (N_2565,N_1475,N_1613);
nand U2566 (N_2566,N_1224,N_1519);
nand U2567 (N_2567,N_1802,N_1896);
and U2568 (N_2568,N_1710,N_1537);
nand U2569 (N_2569,N_1909,N_1711);
nor U2570 (N_2570,N_1891,N_1191);
nor U2571 (N_2571,N_1878,N_1499);
nand U2572 (N_2572,N_1066,N_1833);
nand U2573 (N_2573,N_1149,N_1095);
nand U2574 (N_2574,N_1700,N_1835);
nand U2575 (N_2575,N_1961,N_1728);
and U2576 (N_2576,N_1061,N_1682);
nor U2577 (N_2577,N_1795,N_1406);
xor U2578 (N_2578,N_1906,N_1768);
nand U2579 (N_2579,N_1267,N_1736);
nand U2580 (N_2580,N_1391,N_1787);
nor U2581 (N_2581,N_1196,N_1884);
xor U2582 (N_2582,N_1137,N_1713);
or U2583 (N_2583,N_1324,N_1002);
nand U2584 (N_2584,N_1269,N_1353);
xor U2585 (N_2585,N_1480,N_1658);
nand U2586 (N_2586,N_1919,N_1677);
xnor U2587 (N_2587,N_1678,N_1791);
nor U2588 (N_2588,N_1838,N_1251);
and U2589 (N_2589,N_1210,N_1994);
and U2590 (N_2590,N_1775,N_1074);
nor U2591 (N_2591,N_1267,N_1456);
and U2592 (N_2592,N_1081,N_1587);
nand U2593 (N_2593,N_1073,N_1622);
nor U2594 (N_2594,N_1569,N_1947);
or U2595 (N_2595,N_1227,N_1855);
and U2596 (N_2596,N_1908,N_1885);
and U2597 (N_2597,N_1438,N_1781);
or U2598 (N_2598,N_1725,N_1651);
nor U2599 (N_2599,N_1663,N_1329);
nand U2600 (N_2600,N_1664,N_1761);
or U2601 (N_2601,N_1141,N_1271);
xor U2602 (N_2602,N_1250,N_1671);
and U2603 (N_2603,N_1437,N_1946);
nand U2604 (N_2604,N_1728,N_1880);
nand U2605 (N_2605,N_1606,N_1131);
and U2606 (N_2606,N_1921,N_1077);
nor U2607 (N_2607,N_1568,N_1837);
nand U2608 (N_2608,N_1175,N_1099);
nor U2609 (N_2609,N_1500,N_1593);
and U2610 (N_2610,N_1125,N_1848);
and U2611 (N_2611,N_1005,N_1145);
nor U2612 (N_2612,N_1844,N_1280);
nor U2613 (N_2613,N_1518,N_1059);
nand U2614 (N_2614,N_1824,N_1343);
xor U2615 (N_2615,N_1941,N_1194);
nand U2616 (N_2616,N_1243,N_1071);
nor U2617 (N_2617,N_1196,N_1904);
or U2618 (N_2618,N_1970,N_1119);
or U2619 (N_2619,N_1678,N_1919);
or U2620 (N_2620,N_1046,N_1805);
nor U2621 (N_2621,N_1285,N_1569);
xnor U2622 (N_2622,N_1338,N_1602);
and U2623 (N_2623,N_1359,N_1534);
nor U2624 (N_2624,N_1622,N_1466);
xor U2625 (N_2625,N_1381,N_1003);
nor U2626 (N_2626,N_1262,N_1154);
and U2627 (N_2627,N_1639,N_1158);
and U2628 (N_2628,N_1417,N_1817);
nand U2629 (N_2629,N_1000,N_1891);
nand U2630 (N_2630,N_1428,N_1964);
xnor U2631 (N_2631,N_1017,N_1084);
xnor U2632 (N_2632,N_1468,N_1979);
or U2633 (N_2633,N_1812,N_1738);
xnor U2634 (N_2634,N_1187,N_1024);
xnor U2635 (N_2635,N_1727,N_1687);
and U2636 (N_2636,N_1869,N_1601);
xor U2637 (N_2637,N_1772,N_1159);
nor U2638 (N_2638,N_1979,N_1551);
nand U2639 (N_2639,N_1762,N_1841);
and U2640 (N_2640,N_1897,N_1988);
nand U2641 (N_2641,N_1986,N_1567);
and U2642 (N_2642,N_1193,N_1655);
xnor U2643 (N_2643,N_1118,N_1419);
and U2644 (N_2644,N_1542,N_1776);
or U2645 (N_2645,N_1368,N_1452);
or U2646 (N_2646,N_1182,N_1073);
xor U2647 (N_2647,N_1098,N_1305);
nor U2648 (N_2648,N_1801,N_1136);
nor U2649 (N_2649,N_1353,N_1969);
or U2650 (N_2650,N_1964,N_1617);
xor U2651 (N_2651,N_1876,N_1277);
and U2652 (N_2652,N_1144,N_1083);
and U2653 (N_2653,N_1861,N_1598);
nand U2654 (N_2654,N_1517,N_1876);
nand U2655 (N_2655,N_1992,N_1753);
or U2656 (N_2656,N_1807,N_1732);
or U2657 (N_2657,N_1080,N_1493);
or U2658 (N_2658,N_1805,N_1427);
nor U2659 (N_2659,N_1549,N_1171);
or U2660 (N_2660,N_1406,N_1684);
nor U2661 (N_2661,N_1522,N_1036);
xor U2662 (N_2662,N_1901,N_1491);
or U2663 (N_2663,N_1248,N_1097);
xnor U2664 (N_2664,N_1170,N_1009);
or U2665 (N_2665,N_1810,N_1674);
and U2666 (N_2666,N_1658,N_1853);
and U2667 (N_2667,N_1965,N_1706);
and U2668 (N_2668,N_1964,N_1571);
nor U2669 (N_2669,N_1188,N_1583);
or U2670 (N_2670,N_1463,N_1901);
or U2671 (N_2671,N_1098,N_1532);
and U2672 (N_2672,N_1522,N_1347);
or U2673 (N_2673,N_1709,N_1514);
and U2674 (N_2674,N_1942,N_1303);
nand U2675 (N_2675,N_1846,N_1019);
or U2676 (N_2676,N_1180,N_1730);
nand U2677 (N_2677,N_1506,N_1686);
nor U2678 (N_2678,N_1765,N_1219);
nand U2679 (N_2679,N_1453,N_1074);
nand U2680 (N_2680,N_1975,N_1279);
nor U2681 (N_2681,N_1244,N_1311);
and U2682 (N_2682,N_1821,N_1538);
nand U2683 (N_2683,N_1401,N_1826);
nand U2684 (N_2684,N_1299,N_1999);
and U2685 (N_2685,N_1684,N_1865);
nor U2686 (N_2686,N_1451,N_1993);
xnor U2687 (N_2687,N_1433,N_1485);
xor U2688 (N_2688,N_1787,N_1051);
or U2689 (N_2689,N_1776,N_1585);
xnor U2690 (N_2690,N_1493,N_1371);
or U2691 (N_2691,N_1378,N_1645);
nand U2692 (N_2692,N_1441,N_1454);
and U2693 (N_2693,N_1660,N_1247);
nand U2694 (N_2694,N_1526,N_1116);
or U2695 (N_2695,N_1350,N_1352);
nor U2696 (N_2696,N_1465,N_1192);
nand U2697 (N_2697,N_1368,N_1769);
or U2698 (N_2698,N_1758,N_1572);
nor U2699 (N_2699,N_1635,N_1968);
nand U2700 (N_2700,N_1174,N_1002);
xor U2701 (N_2701,N_1307,N_1868);
and U2702 (N_2702,N_1844,N_1295);
and U2703 (N_2703,N_1003,N_1437);
and U2704 (N_2704,N_1408,N_1879);
xor U2705 (N_2705,N_1518,N_1463);
xor U2706 (N_2706,N_1226,N_1159);
or U2707 (N_2707,N_1048,N_1598);
nand U2708 (N_2708,N_1158,N_1732);
xnor U2709 (N_2709,N_1072,N_1220);
or U2710 (N_2710,N_1492,N_1990);
and U2711 (N_2711,N_1280,N_1588);
and U2712 (N_2712,N_1963,N_1336);
or U2713 (N_2713,N_1868,N_1276);
nand U2714 (N_2714,N_1402,N_1080);
or U2715 (N_2715,N_1970,N_1405);
nor U2716 (N_2716,N_1130,N_1008);
nand U2717 (N_2717,N_1366,N_1923);
or U2718 (N_2718,N_1639,N_1036);
nand U2719 (N_2719,N_1388,N_1951);
or U2720 (N_2720,N_1889,N_1333);
xor U2721 (N_2721,N_1861,N_1425);
and U2722 (N_2722,N_1583,N_1281);
nor U2723 (N_2723,N_1079,N_1700);
and U2724 (N_2724,N_1773,N_1806);
nor U2725 (N_2725,N_1853,N_1604);
and U2726 (N_2726,N_1589,N_1076);
or U2727 (N_2727,N_1289,N_1291);
nor U2728 (N_2728,N_1839,N_1521);
xor U2729 (N_2729,N_1385,N_1554);
xnor U2730 (N_2730,N_1972,N_1322);
nand U2731 (N_2731,N_1798,N_1461);
and U2732 (N_2732,N_1745,N_1155);
nand U2733 (N_2733,N_1400,N_1155);
nor U2734 (N_2734,N_1319,N_1015);
nand U2735 (N_2735,N_1099,N_1064);
nand U2736 (N_2736,N_1916,N_1679);
and U2737 (N_2737,N_1889,N_1207);
nor U2738 (N_2738,N_1266,N_1207);
or U2739 (N_2739,N_1120,N_1462);
and U2740 (N_2740,N_1946,N_1103);
nand U2741 (N_2741,N_1341,N_1491);
xnor U2742 (N_2742,N_1964,N_1157);
nand U2743 (N_2743,N_1842,N_1017);
xnor U2744 (N_2744,N_1384,N_1921);
or U2745 (N_2745,N_1275,N_1801);
xnor U2746 (N_2746,N_1283,N_1317);
and U2747 (N_2747,N_1802,N_1217);
or U2748 (N_2748,N_1696,N_1021);
nor U2749 (N_2749,N_1980,N_1673);
xnor U2750 (N_2750,N_1326,N_1636);
or U2751 (N_2751,N_1753,N_1496);
xnor U2752 (N_2752,N_1182,N_1276);
xnor U2753 (N_2753,N_1618,N_1400);
nand U2754 (N_2754,N_1641,N_1753);
xnor U2755 (N_2755,N_1345,N_1529);
xor U2756 (N_2756,N_1235,N_1940);
nand U2757 (N_2757,N_1632,N_1360);
xor U2758 (N_2758,N_1703,N_1963);
or U2759 (N_2759,N_1413,N_1931);
nor U2760 (N_2760,N_1816,N_1696);
nor U2761 (N_2761,N_1919,N_1369);
or U2762 (N_2762,N_1625,N_1461);
xor U2763 (N_2763,N_1665,N_1995);
or U2764 (N_2764,N_1634,N_1271);
nand U2765 (N_2765,N_1622,N_1710);
nor U2766 (N_2766,N_1039,N_1556);
xor U2767 (N_2767,N_1193,N_1172);
xnor U2768 (N_2768,N_1490,N_1404);
nor U2769 (N_2769,N_1264,N_1251);
and U2770 (N_2770,N_1398,N_1401);
nand U2771 (N_2771,N_1281,N_1971);
nor U2772 (N_2772,N_1617,N_1881);
and U2773 (N_2773,N_1278,N_1252);
nor U2774 (N_2774,N_1072,N_1676);
nor U2775 (N_2775,N_1911,N_1101);
and U2776 (N_2776,N_1076,N_1306);
nand U2777 (N_2777,N_1440,N_1899);
nor U2778 (N_2778,N_1589,N_1141);
nand U2779 (N_2779,N_1722,N_1706);
nor U2780 (N_2780,N_1453,N_1814);
and U2781 (N_2781,N_1945,N_1822);
nand U2782 (N_2782,N_1589,N_1579);
nand U2783 (N_2783,N_1489,N_1738);
and U2784 (N_2784,N_1259,N_1924);
nor U2785 (N_2785,N_1384,N_1313);
nand U2786 (N_2786,N_1520,N_1030);
nand U2787 (N_2787,N_1732,N_1245);
xor U2788 (N_2788,N_1116,N_1377);
or U2789 (N_2789,N_1124,N_1914);
nor U2790 (N_2790,N_1354,N_1667);
or U2791 (N_2791,N_1751,N_1584);
and U2792 (N_2792,N_1820,N_1353);
nand U2793 (N_2793,N_1081,N_1878);
nor U2794 (N_2794,N_1596,N_1170);
xnor U2795 (N_2795,N_1489,N_1340);
or U2796 (N_2796,N_1157,N_1067);
xnor U2797 (N_2797,N_1931,N_1035);
and U2798 (N_2798,N_1430,N_1396);
or U2799 (N_2799,N_1270,N_1124);
or U2800 (N_2800,N_1244,N_1912);
nand U2801 (N_2801,N_1605,N_1265);
or U2802 (N_2802,N_1863,N_1906);
and U2803 (N_2803,N_1847,N_1703);
and U2804 (N_2804,N_1351,N_1395);
xnor U2805 (N_2805,N_1851,N_1862);
and U2806 (N_2806,N_1387,N_1066);
xor U2807 (N_2807,N_1297,N_1876);
nand U2808 (N_2808,N_1646,N_1783);
or U2809 (N_2809,N_1052,N_1693);
nor U2810 (N_2810,N_1961,N_1223);
or U2811 (N_2811,N_1577,N_1613);
and U2812 (N_2812,N_1440,N_1842);
nor U2813 (N_2813,N_1260,N_1182);
nand U2814 (N_2814,N_1070,N_1646);
or U2815 (N_2815,N_1819,N_1201);
or U2816 (N_2816,N_1920,N_1135);
and U2817 (N_2817,N_1191,N_1748);
nand U2818 (N_2818,N_1986,N_1735);
and U2819 (N_2819,N_1468,N_1735);
xnor U2820 (N_2820,N_1793,N_1387);
nor U2821 (N_2821,N_1819,N_1249);
nor U2822 (N_2822,N_1946,N_1638);
nand U2823 (N_2823,N_1654,N_1664);
xor U2824 (N_2824,N_1715,N_1479);
nor U2825 (N_2825,N_1092,N_1476);
or U2826 (N_2826,N_1953,N_1155);
nor U2827 (N_2827,N_1863,N_1137);
or U2828 (N_2828,N_1612,N_1795);
nand U2829 (N_2829,N_1529,N_1107);
nand U2830 (N_2830,N_1873,N_1473);
xor U2831 (N_2831,N_1219,N_1187);
nor U2832 (N_2832,N_1920,N_1428);
or U2833 (N_2833,N_1544,N_1844);
and U2834 (N_2834,N_1455,N_1412);
nand U2835 (N_2835,N_1182,N_1150);
nand U2836 (N_2836,N_1571,N_1590);
nor U2837 (N_2837,N_1145,N_1281);
nor U2838 (N_2838,N_1567,N_1984);
and U2839 (N_2839,N_1878,N_1636);
and U2840 (N_2840,N_1745,N_1983);
nand U2841 (N_2841,N_1885,N_1828);
nand U2842 (N_2842,N_1003,N_1572);
or U2843 (N_2843,N_1335,N_1803);
xnor U2844 (N_2844,N_1285,N_1621);
and U2845 (N_2845,N_1340,N_1172);
or U2846 (N_2846,N_1586,N_1759);
nand U2847 (N_2847,N_1883,N_1490);
nor U2848 (N_2848,N_1609,N_1908);
and U2849 (N_2849,N_1446,N_1604);
nand U2850 (N_2850,N_1402,N_1335);
or U2851 (N_2851,N_1737,N_1781);
nor U2852 (N_2852,N_1283,N_1038);
and U2853 (N_2853,N_1341,N_1838);
nor U2854 (N_2854,N_1944,N_1375);
or U2855 (N_2855,N_1371,N_1578);
nand U2856 (N_2856,N_1989,N_1262);
and U2857 (N_2857,N_1532,N_1575);
nor U2858 (N_2858,N_1284,N_1722);
xnor U2859 (N_2859,N_1960,N_1667);
or U2860 (N_2860,N_1138,N_1776);
or U2861 (N_2861,N_1068,N_1008);
or U2862 (N_2862,N_1637,N_1851);
nor U2863 (N_2863,N_1823,N_1941);
nand U2864 (N_2864,N_1554,N_1510);
or U2865 (N_2865,N_1200,N_1180);
xnor U2866 (N_2866,N_1341,N_1383);
nor U2867 (N_2867,N_1415,N_1391);
nor U2868 (N_2868,N_1762,N_1000);
xnor U2869 (N_2869,N_1841,N_1797);
and U2870 (N_2870,N_1120,N_1878);
nor U2871 (N_2871,N_1206,N_1360);
nor U2872 (N_2872,N_1098,N_1966);
nand U2873 (N_2873,N_1108,N_1742);
and U2874 (N_2874,N_1419,N_1574);
xor U2875 (N_2875,N_1947,N_1575);
nor U2876 (N_2876,N_1459,N_1359);
nor U2877 (N_2877,N_1007,N_1999);
or U2878 (N_2878,N_1865,N_1574);
xnor U2879 (N_2879,N_1077,N_1920);
or U2880 (N_2880,N_1845,N_1523);
and U2881 (N_2881,N_1305,N_1078);
nand U2882 (N_2882,N_1577,N_1889);
nor U2883 (N_2883,N_1008,N_1894);
xnor U2884 (N_2884,N_1266,N_1470);
nand U2885 (N_2885,N_1509,N_1230);
nand U2886 (N_2886,N_1767,N_1401);
nor U2887 (N_2887,N_1752,N_1845);
and U2888 (N_2888,N_1060,N_1049);
nand U2889 (N_2889,N_1738,N_1796);
xor U2890 (N_2890,N_1081,N_1235);
and U2891 (N_2891,N_1760,N_1497);
or U2892 (N_2892,N_1924,N_1047);
and U2893 (N_2893,N_1813,N_1342);
xnor U2894 (N_2894,N_1300,N_1616);
xnor U2895 (N_2895,N_1161,N_1228);
nor U2896 (N_2896,N_1147,N_1549);
or U2897 (N_2897,N_1311,N_1812);
nand U2898 (N_2898,N_1411,N_1926);
nand U2899 (N_2899,N_1118,N_1739);
xnor U2900 (N_2900,N_1028,N_1753);
xor U2901 (N_2901,N_1501,N_1371);
or U2902 (N_2902,N_1948,N_1496);
or U2903 (N_2903,N_1289,N_1042);
xor U2904 (N_2904,N_1471,N_1581);
and U2905 (N_2905,N_1593,N_1729);
xnor U2906 (N_2906,N_1567,N_1519);
nand U2907 (N_2907,N_1385,N_1983);
and U2908 (N_2908,N_1865,N_1878);
or U2909 (N_2909,N_1218,N_1762);
nor U2910 (N_2910,N_1348,N_1870);
or U2911 (N_2911,N_1582,N_1774);
xor U2912 (N_2912,N_1693,N_1528);
xnor U2913 (N_2913,N_1866,N_1225);
nor U2914 (N_2914,N_1380,N_1959);
nor U2915 (N_2915,N_1464,N_1328);
nand U2916 (N_2916,N_1587,N_1842);
and U2917 (N_2917,N_1075,N_1769);
nand U2918 (N_2918,N_1448,N_1027);
nand U2919 (N_2919,N_1370,N_1507);
nand U2920 (N_2920,N_1191,N_1094);
and U2921 (N_2921,N_1461,N_1359);
or U2922 (N_2922,N_1845,N_1292);
xnor U2923 (N_2923,N_1717,N_1706);
or U2924 (N_2924,N_1454,N_1935);
nor U2925 (N_2925,N_1601,N_1843);
nand U2926 (N_2926,N_1618,N_1354);
and U2927 (N_2927,N_1234,N_1335);
xor U2928 (N_2928,N_1887,N_1280);
xor U2929 (N_2929,N_1310,N_1840);
nor U2930 (N_2930,N_1190,N_1733);
and U2931 (N_2931,N_1653,N_1205);
and U2932 (N_2932,N_1350,N_1677);
or U2933 (N_2933,N_1184,N_1318);
nand U2934 (N_2934,N_1877,N_1726);
and U2935 (N_2935,N_1069,N_1429);
or U2936 (N_2936,N_1049,N_1042);
nor U2937 (N_2937,N_1735,N_1942);
xor U2938 (N_2938,N_1990,N_1369);
xor U2939 (N_2939,N_1872,N_1974);
and U2940 (N_2940,N_1083,N_1907);
or U2941 (N_2941,N_1722,N_1237);
nand U2942 (N_2942,N_1060,N_1265);
or U2943 (N_2943,N_1767,N_1509);
xnor U2944 (N_2944,N_1400,N_1012);
nor U2945 (N_2945,N_1793,N_1883);
nor U2946 (N_2946,N_1803,N_1679);
or U2947 (N_2947,N_1121,N_1426);
nor U2948 (N_2948,N_1378,N_1840);
and U2949 (N_2949,N_1026,N_1705);
nand U2950 (N_2950,N_1911,N_1658);
nor U2951 (N_2951,N_1781,N_1468);
xnor U2952 (N_2952,N_1786,N_1876);
nor U2953 (N_2953,N_1669,N_1252);
and U2954 (N_2954,N_1268,N_1988);
or U2955 (N_2955,N_1450,N_1061);
or U2956 (N_2956,N_1673,N_1745);
nand U2957 (N_2957,N_1175,N_1857);
nand U2958 (N_2958,N_1227,N_1754);
nor U2959 (N_2959,N_1531,N_1726);
xor U2960 (N_2960,N_1784,N_1058);
or U2961 (N_2961,N_1407,N_1233);
and U2962 (N_2962,N_1181,N_1521);
nand U2963 (N_2963,N_1216,N_1345);
or U2964 (N_2964,N_1804,N_1836);
nand U2965 (N_2965,N_1365,N_1487);
xnor U2966 (N_2966,N_1458,N_1852);
nand U2967 (N_2967,N_1839,N_1279);
xnor U2968 (N_2968,N_1387,N_1186);
nand U2969 (N_2969,N_1670,N_1901);
or U2970 (N_2970,N_1829,N_1765);
nor U2971 (N_2971,N_1923,N_1941);
or U2972 (N_2972,N_1669,N_1106);
or U2973 (N_2973,N_1995,N_1600);
or U2974 (N_2974,N_1374,N_1217);
and U2975 (N_2975,N_1720,N_1061);
xor U2976 (N_2976,N_1286,N_1339);
or U2977 (N_2977,N_1669,N_1035);
or U2978 (N_2978,N_1824,N_1427);
nor U2979 (N_2979,N_1332,N_1005);
nand U2980 (N_2980,N_1324,N_1300);
nor U2981 (N_2981,N_1688,N_1017);
nand U2982 (N_2982,N_1607,N_1295);
or U2983 (N_2983,N_1668,N_1732);
or U2984 (N_2984,N_1419,N_1141);
and U2985 (N_2985,N_1263,N_1107);
xnor U2986 (N_2986,N_1122,N_1457);
nand U2987 (N_2987,N_1893,N_1179);
xnor U2988 (N_2988,N_1749,N_1053);
xnor U2989 (N_2989,N_1849,N_1002);
nand U2990 (N_2990,N_1098,N_1935);
and U2991 (N_2991,N_1209,N_1615);
and U2992 (N_2992,N_1595,N_1955);
or U2993 (N_2993,N_1651,N_1592);
nand U2994 (N_2994,N_1584,N_1869);
xnor U2995 (N_2995,N_1328,N_1052);
or U2996 (N_2996,N_1454,N_1977);
xnor U2997 (N_2997,N_1811,N_1498);
nand U2998 (N_2998,N_1813,N_1709);
or U2999 (N_2999,N_1351,N_1727);
or U3000 (N_3000,N_2052,N_2769);
nor U3001 (N_3001,N_2643,N_2698);
nor U3002 (N_3002,N_2898,N_2558);
xor U3003 (N_3003,N_2192,N_2340);
nand U3004 (N_3004,N_2519,N_2156);
nor U3005 (N_3005,N_2064,N_2116);
and U3006 (N_3006,N_2183,N_2754);
nand U3007 (N_3007,N_2756,N_2590);
and U3008 (N_3008,N_2556,N_2843);
xnor U3009 (N_3009,N_2215,N_2013);
and U3010 (N_3010,N_2806,N_2456);
or U3011 (N_3011,N_2933,N_2567);
nand U3012 (N_3012,N_2951,N_2150);
and U3013 (N_3013,N_2853,N_2303);
nor U3014 (N_3014,N_2483,N_2328);
xor U3015 (N_3015,N_2321,N_2514);
nand U3016 (N_3016,N_2286,N_2316);
or U3017 (N_3017,N_2784,N_2538);
xor U3018 (N_3018,N_2135,N_2385);
nand U3019 (N_3019,N_2731,N_2677);
nand U3020 (N_3020,N_2145,N_2568);
xnor U3021 (N_3021,N_2096,N_2256);
xor U3022 (N_3022,N_2720,N_2804);
xor U3023 (N_3023,N_2608,N_2897);
nand U3024 (N_3024,N_2219,N_2870);
or U3025 (N_3025,N_2840,N_2586);
xnor U3026 (N_3026,N_2393,N_2300);
nand U3027 (N_3027,N_2403,N_2924);
nand U3028 (N_3028,N_2553,N_2847);
and U3029 (N_3029,N_2450,N_2092);
nor U3030 (N_3030,N_2954,N_2195);
and U3031 (N_3031,N_2762,N_2005);
and U3032 (N_3032,N_2277,N_2711);
and U3033 (N_3033,N_2622,N_2181);
or U3034 (N_3034,N_2324,N_2065);
xor U3035 (N_3035,N_2260,N_2470);
or U3036 (N_3036,N_2548,N_2780);
or U3037 (N_3037,N_2845,N_2705);
and U3038 (N_3038,N_2902,N_2903);
nor U3039 (N_3039,N_2476,N_2722);
xnor U3040 (N_3040,N_2326,N_2571);
or U3041 (N_3041,N_2123,N_2048);
or U3042 (N_3042,N_2108,N_2199);
nor U3043 (N_3043,N_2111,N_2376);
nand U3044 (N_3044,N_2383,N_2703);
nor U3045 (N_3045,N_2889,N_2280);
xnor U3046 (N_3046,N_2288,N_2886);
and U3047 (N_3047,N_2752,N_2479);
or U3048 (N_3048,N_2344,N_2781);
and U3049 (N_3049,N_2066,N_2615);
xor U3050 (N_3050,N_2671,N_2121);
or U3051 (N_3051,N_2059,N_2103);
nand U3052 (N_3052,N_2075,N_2319);
and U3053 (N_3053,N_2070,N_2651);
nor U3054 (N_3054,N_2496,N_2530);
and U3055 (N_3055,N_2139,N_2390);
nand U3056 (N_3056,N_2320,N_2982);
nor U3057 (N_3057,N_2387,N_2373);
or U3058 (N_3058,N_2291,N_2161);
or U3059 (N_3059,N_2492,N_2855);
and U3060 (N_3060,N_2351,N_2824);
nand U3061 (N_3061,N_2576,N_2517);
nand U3062 (N_3062,N_2991,N_2407);
xnor U3063 (N_3063,N_2910,N_2415);
nor U3064 (N_3064,N_2687,N_2079);
xnor U3065 (N_3065,N_2660,N_2396);
nor U3066 (N_3066,N_2544,N_2697);
nand U3067 (N_3067,N_2680,N_2453);
and U3068 (N_3068,N_2871,N_2078);
nand U3069 (N_3069,N_2799,N_2063);
nand U3070 (N_3070,N_2274,N_2743);
or U3071 (N_3071,N_2733,N_2644);
nand U3072 (N_3072,N_2433,N_2691);
nand U3073 (N_3073,N_2253,N_2023);
and U3074 (N_3074,N_2186,N_2829);
nor U3075 (N_3075,N_2466,N_2893);
or U3076 (N_3076,N_2685,N_2931);
nor U3077 (N_3077,N_2487,N_2489);
nand U3078 (N_3078,N_2707,N_2750);
xor U3079 (N_3079,N_2400,N_2346);
nand U3080 (N_3080,N_2867,N_2439);
nand U3081 (N_3081,N_2729,N_2170);
nor U3082 (N_3082,N_2266,N_2412);
nor U3083 (N_3083,N_2455,N_2936);
xnor U3084 (N_3084,N_2234,N_2832);
xor U3085 (N_3085,N_2823,N_2222);
nor U3086 (N_3086,N_2033,N_2899);
or U3087 (N_3087,N_2881,N_2540);
and U3088 (N_3088,N_2332,N_2503);
xor U3089 (N_3089,N_2034,N_2989);
nor U3090 (N_3090,N_2746,N_2378);
nand U3091 (N_3091,N_2649,N_2996);
nor U3092 (N_3092,N_2647,N_2485);
or U3093 (N_3093,N_2993,N_2411);
or U3094 (N_3094,N_2419,N_2448);
nor U3095 (N_3095,N_2721,N_2499);
or U3096 (N_3096,N_2976,N_2603);
nand U3097 (N_3097,N_2361,N_2205);
nor U3098 (N_3098,N_2481,N_2851);
and U3099 (N_3099,N_2408,N_2473);
or U3100 (N_3100,N_2301,N_2375);
and U3101 (N_3101,N_2279,N_2238);
nor U3102 (N_3102,N_2778,N_2157);
nor U3103 (N_3103,N_2024,N_2020);
nor U3104 (N_3104,N_2113,N_2213);
nor U3105 (N_3105,N_2038,N_2755);
nand U3106 (N_3106,N_2307,N_2016);
nand U3107 (N_3107,N_2826,N_2596);
and U3108 (N_3108,N_2188,N_2665);
nand U3109 (N_3109,N_2774,N_2626);
or U3110 (N_3110,N_2146,N_2144);
or U3111 (N_3111,N_2668,N_2381);
and U3112 (N_3112,N_2354,N_2735);
nand U3113 (N_3113,N_2475,N_2726);
or U3114 (N_3114,N_2527,N_2153);
xnor U3115 (N_3115,N_2552,N_2682);
xnor U3116 (N_3116,N_2347,N_2086);
nor U3117 (N_3117,N_2045,N_2230);
or U3118 (N_3118,N_2271,N_2179);
or U3119 (N_3119,N_2012,N_2771);
and U3120 (N_3120,N_2399,N_2001);
or U3121 (N_3121,N_2563,N_2652);
nand U3122 (N_3122,N_2290,N_2640);
nor U3123 (N_3123,N_2437,N_2624);
and U3124 (N_3124,N_2357,N_2427);
and U3125 (N_3125,N_2609,N_2734);
xor U3126 (N_3126,N_2147,N_2151);
xor U3127 (N_3127,N_2356,N_2678);
and U3128 (N_3128,N_2262,N_2040);
and U3129 (N_3129,N_2670,N_2801);
or U3130 (N_3130,N_2792,N_2573);
and U3131 (N_3131,N_2463,N_2287);
and U3132 (N_3132,N_2039,N_2180);
xor U3133 (N_3133,N_2152,N_2493);
nand U3134 (N_3134,N_2486,N_2133);
nor U3135 (N_3135,N_2459,N_2283);
and U3136 (N_3136,N_2642,N_2629);
nand U3137 (N_3137,N_2768,N_2782);
xnor U3138 (N_3138,N_2969,N_2441);
and U3139 (N_3139,N_2429,N_2424);
nand U3140 (N_3140,N_2334,N_2964);
xnor U3141 (N_3141,N_2716,N_2593);
nand U3142 (N_3142,N_2035,N_2841);
nor U3143 (N_3143,N_2068,N_2862);
xor U3144 (N_3144,N_2817,N_2606);
or U3145 (N_3145,N_2641,N_2158);
nand U3146 (N_3146,N_2732,N_2822);
nor U3147 (N_3147,N_2342,N_2686);
or U3148 (N_3148,N_2592,N_2074);
nor U3149 (N_3149,N_2474,N_2598);
nor U3150 (N_3150,N_2082,N_2767);
nor U3151 (N_3151,N_2143,N_2120);
and U3152 (N_3152,N_2241,N_2060);
xnor U3153 (N_3153,N_2207,N_2449);
nor U3154 (N_3154,N_2249,N_2512);
xnor U3155 (N_3155,N_2115,N_2118);
or U3156 (N_3156,N_2027,N_2591);
nand U3157 (N_3157,N_2839,N_2008);
nor U3158 (N_3158,N_2397,N_2764);
nand U3159 (N_3159,N_2923,N_2257);
nor U3160 (N_3160,N_2416,N_2259);
nand U3161 (N_3161,N_2384,N_2509);
nor U3162 (N_3162,N_2233,N_2715);
xor U3163 (N_3163,N_2236,N_2193);
or U3164 (N_3164,N_2560,N_2638);
xor U3165 (N_3165,N_2612,N_2173);
nand U3166 (N_3166,N_2919,N_2907);
and U3167 (N_3167,N_2329,N_2901);
xnor U3168 (N_3168,N_2928,N_2825);
xnor U3169 (N_3169,N_2442,N_2635);
or U3170 (N_3170,N_2171,N_2104);
xor U3171 (N_3171,N_2404,N_2607);
and U3172 (N_3172,N_2659,N_2110);
and U3173 (N_3173,N_2454,N_2551);
and U3174 (N_3174,N_2892,N_2088);
nand U3175 (N_3175,N_2701,N_2336);
nor U3176 (N_3176,N_2564,N_2258);
xnor U3177 (N_3177,N_2337,N_2718);
xor U3178 (N_3178,N_2895,N_2873);
nand U3179 (N_3179,N_2816,N_2107);
nand U3180 (N_3180,N_2223,N_2683);
and U3181 (N_3181,N_2263,N_2681);
or U3182 (N_3182,N_2748,N_2136);
or U3183 (N_3183,N_2468,N_2330);
and U3184 (N_3184,N_2141,N_2490);
nor U3185 (N_3185,N_2878,N_2518);
and U3186 (N_3186,N_2112,N_2003);
nand U3187 (N_3187,N_2478,N_2057);
nand U3188 (N_3188,N_2946,N_2968);
nor U3189 (N_3189,N_2246,N_2401);
or U3190 (N_3190,N_2973,N_2655);
and U3191 (N_3191,N_2852,N_2206);
and U3192 (N_3192,N_2975,N_2338);
xnor U3193 (N_3193,N_2155,N_2842);
nor U3194 (N_3194,N_2937,N_2235);
nand U3195 (N_3195,N_2838,N_2597);
xnor U3196 (N_3196,N_2406,N_2138);
xor U3197 (N_3197,N_2097,N_2917);
xor U3198 (N_3198,N_2741,N_2377);
or U3199 (N_3199,N_2605,N_2498);
xnor U3200 (N_3200,N_2243,N_2617);
nor U3201 (N_3201,N_2394,N_2916);
or U3202 (N_3202,N_2464,N_2539);
and U3203 (N_3203,N_2327,N_2696);
or U3204 (N_3204,N_2046,N_2363);
nor U3205 (N_3205,N_2986,N_2245);
or U3206 (N_3206,N_2458,N_2938);
or U3207 (N_3207,N_2998,N_2572);
nor U3208 (N_3208,N_2710,N_2389);
nor U3209 (N_3209,N_2550,N_2861);
nand U3210 (N_3210,N_2943,N_2542);
or U3211 (N_3211,N_2737,N_2105);
nor U3212 (N_3212,N_2164,N_2929);
nand U3213 (N_3213,N_2240,N_2983);
and U3214 (N_3214,N_2443,N_2160);
nor U3215 (N_3215,N_2315,N_2508);
or U3216 (N_3216,N_2927,N_2805);
or U3217 (N_3217,N_2252,N_2744);
xnor U3218 (N_3218,N_2457,N_2728);
and U3219 (N_3219,N_2106,N_2083);
xor U3220 (N_3220,N_2058,N_2440);
or U3221 (N_3221,N_2545,N_2913);
and U3222 (N_3222,N_2358,N_2312);
or U3223 (N_3223,N_2758,N_2030);
xor U3224 (N_3224,N_2472,N_2264);
xor U3225 (N_3225,N_2438,N_2294);
xor U3226 (N_3226,N_2694,N_2885);
xor U3227 (N_3227,N_2275,N_2981);
or U3228 (N_3228,N_2452,N_2790);
xor U3229 (N_3229,N_2185,N_2557);
nand U3230 (N_3230,N_2882,N_2430);
and U3231 (N_3231,N_2634,N_2080);
nor U3232 (N_3232,N_2465,N_2584);
xor U3233 (N_3233,N_2350,N_2071);
or U3234 (N_3234,N_2210,N_2887);
nor U3235 (N_3235,N_2537,N_2611);
and U3236 (N_3236,N_2434,N_2610);
nand U3237 (N_3237,N_2579,N_2272);
nand U3238 (N_3238,N_2248,N_2765);
or U3239 (N_3239,N_2190,N_2979);
nand U3240 (N_3240,N_2226,N_2021);
and U3241 (N_3241,N_2884,N_2445);
nor U3242 (N_3242,N_2119,N_2239);
nand U3243 (N_3243,N_2006,N_2601);
or U3244 (N_3244,N_2796,N_2997);
xnor U3245 (N_3245,N_2322,N_2041);
and U3246 (N_3246,N_2793,N_2727);
xnor U3247 (N_3247,N_2658,N_2967);
and U3248 (N_3248,N_2410,N_2561);
nand U3249 (N_3249,N_2507,N_2614);
or U3250 (N_3250,N_2331,N_2093);
xnor U3251 (N_3251,N_2977,N_2753);
xnor U3252 (N_3252,N_2896,N_2175);
nand U3253 (N_3253,N_2522,N_2395);
xnor U3254 (N_3254,N_2094,N_2432);
or U3255 (N_3255,N_2846,N_2723);
and U3256 (N_3256,N_2761,N_2566);
nor U3257 (N_3257,N_2374,N_2906);
xnor U3258 (N_3258,N_2305,N_2345);
or U3259 (N_3259,N_2461,N_2621);
and U3260 (N_3260,N_2879,N_2314);
nand U3261 (N_3261,N_2061,N_2420);
or U3262 (N_3262,N_2306,N_2676);
and U3263 (N_3263,N_2883,N_2015);
nor U3264 (N_3264,N_2541,N_2877);
xnor U3265 (N_3265,N_2688,N_2124);
xnor U3266 (N_3266,N_2127,N_2036);
or U3267 (N_3267,N_2209,N_2516);
nand U3268 (N_3268,N_2055,N_2911);
nand U3269 (N_3269,N_2828,N_2582);
or U3270 (N_3270,N_2662,N_2630);
nor U3271 (N_3271,N_2405,N_2081);
nand U3272 (N_3272,N_2578,N_2747);
nand U3273 (N_3273,N_2856,N_2679);
nor U3274 (N_3274,N_2142,N_2335);
nand U3275 (N_3275,N_2864,N_2914);
or U3276 (N_3276,N_2921,N_2978);
nor U3277 (N_3277,N_2858,N_2802);
xor U3278 (N_3278,N_2304,N_2296);
or U3279 (N_3279,N_2289,N_2776);
xnor U3280 (N_3280,N_2216,N_2625);
or U3281 (N_3281,N_2325,N_2000);
or U3282 (N_3282,N_2201,N_2085);
or U3283 (N_3283,N_2369,N_2787);
nand U3284 (N_3284,N_2505,N_2043);
nor U3285 (N_3285,N_2599,N_2834);
or U3286 (N_3286,N_2689,N_2912);
or U3287 (N_3287,N_2785,N_2925);
and U3288 (N_3288,N_2953,N_2724);
or U3289 (N_3289,N_2706,N_2469);
or U3290 (N_3290,N_2583,N_2242);
nor U3291 (N_3291,N_2821,N_2848);
nor U3292 (N_3292,N_2225,N_2506);
and U3293 (N_3293,N_2663,N_2820);
nand U3294 (N_3294,N_2313,N_2056);
nand U3295 (N_3295,N_2451,N_2182);
and U3296 (N_3296,N_2019,N_2631);
nand U3297 (N_3297,N_2809,N_2247);
nand U3298 (N_3298,N_2007,N_2178);
nand U3299 (N_3299,N_2779,N_2684);
or U3300 (N_3300,N_2084,N_2494);
xor U3301 (N_3301,N_2637,N_2211);
nand U3302 (N_3302,N_2053,N_2690);
nor U3303 (N_3303,N_2276,N_2069);
nand U3304 (N_3304,N_2231,N_2428);
nand U3305 (N_3305,N_2212,N_2543);
nor U3306 (N_3306,N_2585,N_2117);
or U3307 (N_3307,N_2446,N_2054);
nor U3308 (N_3308,N_2218,N_2109);
or U3309 (N_3309,N_2844,N_2292);
or U3310 (N_3310,N_2772,N_2431);
and U3311 (N_3311,N_2866,N_2187);
nor U3312 (N_3312,N_2812,N_2391);
nand U3313 (N_3313,N_2920,N_2942);
xor U3314 (N_3314,N_2382,N_2278);
xor U3315 (N_3315,N_2890,N_2815);
xnor U3316 (N_3316,N_2952,N_2200);
nor U3317 (N_3317,N_2589,N_2777);
or U3318 (N_3318,N_2992,N_2860);
and U3319 (N_3319,N_2282,N_2130);
nand U3320 (N_3320,N_2224,N_2559);
nand U3321 (N_3321,N_2939,N_2126);
xor U3322 (N_3322,N_2380,N_2909);
nor U3323 (N_3323,N_2738,N_2051);
nand U3324 (N_3324,N_2196,N_2497);
nand U3325 (N_3325,N_2349,N_2368);
nor U3326 (N_3326,N_2203,N_2669);
nand U3327 (N_3327,N_2859,N_2810);
xor U3328 (N_3328,N_2162,N_2632);
and U3329 (N_3329,N_2818,N_2011);
xor U3330 (N_3330,N_2739,N_2653);
nor U3331 (N_3331,N_2700,N_2129);
nand U3332 (N_3332,N_2032,N_2797);
xnor U3333 (N_3333,N_2740,N_2017);
nor U3334 (N_3334,N_2414,N_2409);
nor U3335 (N_3335,N_2656,N_2674);
and U3336 (N_3336,N_2714,N_2513);
and U3337 (N_3337,N_2667,N_2044);
and U3338 (N_3338,N_2984,N_2900);
xor U3339 (N_3339,N_2837,N_2220);
nand U3340 (N_3340,N_2819,N_2602);
or U3341 (N_3341,N_2491,N_2811);
nand U3342 (N_3342,N_2177,N_2095);
xnor U3343 (N_3343,N_2214,N_2298);
nor U3344 (N_3344,N_2713,N_2348);
nor U3345 (N_3345,N_2891,N_2831);
xnor U3346 (N_3346,N_2229,N_2184);
nor U3347 (N_3347,N_2128,N_2388);
nand U3348 (N_3348,N_2999,N_2029);
and U3349 (N_3349,N_2482,N_2645);
nor U3350 (N_3350,N_2595,N_2398);
and U3351 (N_3351,N_2009,N_2339);
and U3352 (N_3352,N_2786,N_2633);
nor U3353 (N_3353,N_2132,N_2309);
nor U3354 (N_3354,N_2962,N_2392);
xor U3355 (N_3355,N_2562,N_2956);
xor U3356 (N_3356,N_2959,N_2198);
nor U3357 (N_3357,N_2308,N_2908);
nor U3358 (N_3358,N_2874,N_2935);
nand U3359 (N_3359,N_2050,N_2789);
xor U3360 (N_3360,N_2835,N_2894);
nand U3361 (N_3361,N_2159,N_2073);
nand U3362 (N_3362,N_2857,N_2049);
xnor U3363 (N_3363,N_2089,N_2619);
and U3364 (N_3364,N_2646,N_2830);
xor U3365 (N_3365,N_2934,N_2208);
nor U3366 (N_3366,N_2704,N_2949);
xor U3367 (N_3367,N_2987,N_2194);
nor U3368 (N_3368,N_2569,N_2323);
or U3369 (N_3369,N_2849,N_2281);
nor U3370 (N_3370,N_2520,N_2947);
xnor U3371 (N_3371,N_2620,N_2444);
xnor U3372 (N_3372,N_2504,N_2114);
xor U3373 (N_3373,N_2966,N_2985);
nor U3374 (N_3374,N_2317,N_2709);
xor U3375 (N_3375,N_2355,N_2730);
xnor U3376 (N_3376,N_2791,N_2269);
or U3377 (N_3377,N_2604,N_2672);
and U3378 (N_3378,N_2627,N_2367);
xor U3379 (N_3379,N_2770,N_2421);
or U3380 (N_3380,N_2963,N_2875);
or U3381 (N_3381,N_2546,N_2197);
or U3382 (N_3382,N_2650,N_2510);
and U3383 (N_3383,N_2836,N_2125);
nor U3384 (N_3384,N_2462,N_2788);
xor U3385 (N_3385,N_2692,N_2702);
nand U3386 (N_3386,N_2359,N_2850);
and U3387 (N_3387,N_2808,N_2751);
nor U3388 (N_3388,N_2166,N_2501);
xnor U3389 (N_3389,N_2531,N_2090);
nor U3390 (N_3390,N_2028,N_2783);
nor U3391 (N_3391,N_2423,N_2958);
nand U3392 (N_3392,N_2863,N_2955);
xor U3393 (N_3393,N_2961,N_2948);
xnor U3394 (N_3394,N_2775,N_2371);
and U3395 (N_3395,N_2763,N_2310);
nor U3396 (N_3396,N_2915,N_2265);
nand U3397 (N_3397,N_2418,N_2575);
or U3398 (N_3398,N_2719,N_2343);
or U3399 (N_3399,N_2965,N_2759);
and U3400 (N_3400,N_2435,N_2268);
or U3401 (N_3401,N_2189,N_2945);
nor U3402 (N_3402,N_2425,N_2022);
nor U3403 (N_3403,N_2285,N_2749);
nand U3404 (N_3404,N_2072,N_2639);
or U3405 (N_3405,N_2417,N_2467);
nand U3406 (N_3406,N_2944,N_2480);
and U3407 (N_3407,N_2657,N_2244);
or U3408 (N_3408,N_2666,N_2854);
nor U3409 (N_3409,N_2654,N_2010);
or U3410 (N_3410,N_2379,N_2102);
or U3411 (N_3411,N_2302,N_2352);
nand U3412 (N_3412,N_2869,N_2026);
and U3413 (N_3413,N_2365,N_2536);
nor U3414 (N_3414,N_2284,N_2648);
xor U3415 (N_3415,N_2814,N_2970);
xnor U3416 (N_3416,N_2098,N_2270);
or U3417 (N_3417,N_2581,N_2436);
or U3418 (N_3418,N_2370,N_2717);
and U3419 (N_3419,N_2957,N_2994);
or U3420 (N_3420,N_2712,N_2413);
nor U3421 (N_3421,N_2031,N_2594);
nor U3422 (N_3422,N_2255,N_2535);
or U3423 (N_3423,N_2293,N_2077);
and U3424 (N_3424,N_2267,N_2515);
and U3425 (N_3425,N_2299,N_2251);
nand U3426 (N_3426,N_2447,N_2980);
and U3427 (N_3427,N_2795,N_2695);
nand U3428 (N_3428,N_2693,N_2311);
nor U3429 (N_3429,N_2484,N_2636);
and U3430 (N_3430,N_2827,N_2760);
xnor U3431 (N_3431,N_2148,N_2757);
nand U3432 (N_3432,N_2002,N_2426);
nor U3433 (N_3433,N_2122,N_2524);
nor U3434 (N_3434,N_2523,N_2167);
or U3435 (N_3435,N_2295,N_2872);
nand U3436 (N_3436,N_2364,N_2025);
or U3437 (N_3437,N_2067,N_2237);
xnor U3438 (N_3438,N_2333,N_2580);
and U3439 (N_3439,N_2922,N_2725);
nor U3440 (N_3440,N_2154,N_2100);
xor U3441 (N_3441,N_2554,N_2047);
nand U3442 (N_3442,N_2460,N_2880);
nand U3443 (N_3443,N_2533,N_2528);
or U3444 (N_3444,N_2570,N_2773);
nor U3445 (N_3445,N_2500,N_2169);
xor U3446 (N_3446,N_2076,N_2091);
nand U3447 (N_3447,N_2547,N_2062);
or U3448 (N_3448,N_2163,N_2742);
nand U3449 (N_3449,N_2477,N_2587);
xor U3450 (N_3450,N_2675,N_2661);
nor U3451 (N_3451,N_2988,N_2664);
xnor U3452 (N_3452,N_2174,N_2521);
nor U3453 (N_3453,N_2261,N_2618);
nand U3454 (N_3454,N_2227,N_2574);
xor U3455 (N_3455,N_2736,N_2960);
nor U3456 (N_3456,N_2932,N_2488);
xnor U3457 (N_3457,N_2565,N_2708);
nand U3458 (N_3458,N_2250,N_2888);
or U3459 (N_3459,N_2204,N_2534);
or U3460 (N_3460,N_2588,N_2004);
nor U3461 (N_3461,N_2803,N_2613);
nor U3462 (N_3462,N_2273,N_2876);
nand U3463 (N_3463,N_2532,N_2940);
nor U3464 (N_3464,N_2037,N_2918);
xor U3465 (N_3465,N_2502,N_2623);
nor U3466 (N_3466,N_2529,N_2318);
or U3467 (N_3467,N_2577,N_2168);
xnor U3468 (N_3468,N_2549,N_2087);
nor U3469 (N_3469,N_2926,N_2228);
nor U3470 (N_3470,N_2995,N_2353);
nor U3471 (N_3471,N_2254,N_2149);
xnor U3472 (N_3472,N_2865,N_2018);
nand U3473 (N_3473,N_2341,N_2191);
or U3474 (N_3474,N_2386,N_2099);
nor U3475 (N_3475,N_2101,N_2555);
or U3476 (N_3476,N_2833,N_2794);
or U3477 (N_3477,N_2798,N_2673);
or U3478 (N_3478,N_2950,N_2366);
or U3479 (N_3479,N_2766,N_2176);
and U3480 (N_3480,N_2202,N_2525);
or U3481 (N_3481,N_2990,N_2165);
and U3482 (N_3482,N_2905,N_2471);
nand U3483 (N_3483,N_2042,N_2495);
and U3484 (N_3484,N_2699,N_2232);
nand U3485 (N_3485,N_2297,N_2813);
nor U3486 (N_3486,N_2974,N_2600);
or U3487 (N_3487,N_2360,N_2526);
and U3488 (N_3488,N_2134,N_2941);
nor U3489 (N_3489,N_2422,N_2014);
nor U3490 (N_3490,N_2807,N_2402);
or U3491 (N_3491,N_2971,N_2172);
and U3492 (N_3492,N_2972,N_2362);
nor U3493 (N_3493,N_2904,N_2131);
xor U3494 (N_3494,N_2628,N_2511);
and U3495 (N_3495,N_2745,N_2140);
nor U3496 (N_3496,N_2137,N_2217);
or U3497 (N_3497,N_2930,N_2372);
nor U3498 (N_3498,N_2616,N_2868);
and U3499 (N_3499,N_2800,N_2221);
nand U3500 (N_3500,N_2720,N_2058);
and U3501 (N_3501,N_2070,N_2598);
nor U3502 (N_3502,N_2569,N_2069);
or U3503 (N_3503,N_2996,N_2870);
nor U3504 (N_3504,N_2749,N_2429);
and U3505 (N_3505,N_2052,N_2656);
nand U3506 (N_3506,N_2978,N_2404);
nand U3507 (N_3507,N_2973,N_2352);
nand U3508 (N_3508,N_2266,N_2055);
nor U3509 (N_3509,N_2664,N_2627);
xor U3510 (N_3510,N_2949,N_2122);
nor U3511 (N_3511,N_2178,N_2118);
nand U3512 (N_3512,N_2214,N_2427);
xnor U3513 (N_3513,N_2024,N_2529);
nand U3514 (N_3514,N_2208,N_2467);
or U3515 (N_3515,N_2174,N_2537);
xnor U3516 (N_3516,N_2630,N_2705);
and U3517 (N_3517,N_2378,N_2527);
or U3518 (N_3518,N_2875,N_2100);
or U3519 (N_3519,N_2222,N_2972);
xnor U3520 (N_3520,N_2455,N_2582);
nand U3521 (N_3521,N_2455,N_2721);
nor U3522 (N_3522,N_2578,N_2386);
nand U3523 (N_3523,N_2772,N_2663);
and U3524 (N_3524,N_2897,N_2109);
nor U3525 (N_3525,N_2017,N_2179);
and U3526 (N_3526,N_2474,N_2721);
or U3527 (N_3527,N_2410,N_2786);
and U3528 (N_3528,N_2041,N_2786);
nand U3529 (N_3529,N_2235,N_2722);
xnor U3530 (N_3530,N_2772,N_2370);
nor U3531 (N_3531,N_2524,N_2507);
or U3532 (N_3532,N_2221,N_2169);
or U3533 (N_3533,N_2299,N_2872);
nand U3534 (N_3534,N_2893,N_2673);
or U3535 (N_3535,N_2317,N_2133);
xor U3536 (N_3536,N_2681,N_2841);
nor U3537 (N_3537,N_2244,N_2493);
and U3538 (N_3538,N_2334,N_2434);
xnor U3539 (N_3539,N_2191,N_2763);
nor U3540 (N_3540,N_2453,N_2973);
xor U3541 (N_3541,N_2311,N_2179);
nand U3542 (N_3542,N_2194,N_2757);
and U3543 (N_3543,N_2045,N_2761);
and U3544 (N_3544,N_2774,N_2195);
nand U3545 (N_3545,N_2623,N_2627);
xnor U3546 (N_3546,N_2366,N_2382);
and U3547 (N_3547,N_2211,N_2417);
and U3548 (N_3548,N_2771,N_2163);
nand U3549 (N_3549,N_2423,N_2808);
nand U3550 (N_3550,N_2978,N_2897);
nor U3551 (N_3551,N_2648,N_2317);
xor U3552 (N_3552,N_2282,N_2487);
and U3553 (N_3553,N_2040,N_2945);
nand U3554 (N_3554,N_2484,N_2212);
nor U3555 (N_3555,N_2965,N_2005);
xor U3556 (N_3556,N_2141,N_2249);
and U3557 (N_3557,N_2168,N_2548);
or U3558 (N_3558,N_2247,N_2926);
nand U3559 (N_3559,N_2824,N_2309);
nand U3560 (N_3560,N_2815,N_2612);
nor U3561 (N_3561,N_2523,N_2425);
xor U3562 (N_3562,N_2720,N_2937);
or U3563 (N_3563,N_2681,N_2604);
and U3564 (N_3564,N_2924,N_2477);
and U3565 (N_3565,N_2913,N_2440);
xor U3566 (N_3566,N_2145,N_2627);
and U3567 (N_3567,N_2284,N_2807);
xnor U3568 (N_3568,N_2751,N_2908);
and U3569 (N_3569,N_2997,N_2017);
and U3570 (N_3570,N_2786,N_2045);
nand U3571 (N_3571,N_2202,N_2132);
nor U3572 (N_3572,N_2363,N_2392);
nor U3573 (N_3573,N_2872,N_2727);
nand U3574 (N_3574,N_2425,N_2479);
xor U3575 (N_3575,N_2764,N_2460);
or U3576 (N_3576,N_2726,N_2894);
nand U3577 (N_3577,N_2647,N_2334);
xnor U3578 (N_3578,N_2739,N_2055);
or U3579 (N_3579,N_2341,N_2746);
xnor U3580 (N_3580,N_2152,N_2278);
nor U3581 (N_3581,N_2308,N_2815);
and U3582 (N_3582,N_2201,N_2495);
and U3583 (N_3583,N_2009,N_2344);
nand U3584 (N_3584,N_2523,N_2269);
nand U3585 (N_3585,N_2036,N_2279);
nor U3586 (N_3586,N_2710,N_2199);
xnor U3587 (N_3587,N_2088,N_2887);
nand U3588 (N_3588,N_2151,N_2850);
xnor U3589 (N_3589,N_2991,N_2761);
nor U3590 (N_3590,N_2305,N_2280);
and U3591 (N_3591,N_2475,N_2801);
or U3592 (N_3592,N_2990,N_2601);
nor U3593 (N_3593,N_2023,N_2745);
nand U3594 (N_3594,N_2673,N_2258);
and U3595 (N_3595,N_2177,N_2441);
xor U3596 (N_3596,N_2471,N_2683);
xor U3597 (N_3597,N_2888,N_2238);
nand U3598 (N_3598,N_2593,N_2207);
nor U3599 (N_3599,N_2563,N_2457);
nand U3600 (N_3600,N_2194,N_2758);
or U3601 (N_3601,N_2529,N_2135);
and U3602 (N_3602,N_2551,N_2500);
and U3603 (N_3603,N_2896,N_2397);
xnor U3604 (N_3604,N_2792,N_2556);
or U3605 (N_3605,N_2798,N_2390);
or U3606 (N_3606,N_2860,N_2305);
xor U3607 (N_3607,N_2106,N_2745);
or U3608 (N_3608,N_2217,N_2957);
nor U3609 (N_3609,N_2934,N_2585);
nand U3610 (N_3610,N_2411,N_2236);
or U3611 (N_3611,N_2712,N_2128);
or U3612 (N_3612,N_2079,N_2005);
and U3613 (N_3613,N_2983,N_2073);
and U3614 (N_3614,N_2363,N_2420);
or U3615 (N_3615,N_2807,N_2995);
xnor U3616 (N_3616,N_2798,N_2739);
nor U3617 (N_3617,N_2254,N_2064);
nand U3618 (N_3618,N_2487,N_2605);
xnor U3619 (N_3619,N_2811,N_2047);
nor U3620 (N_3620,N_2749,N_2826);
nand U3621 (N_3621,N_2557,N_2426);
xor U3622 (N_3622,N_2340,N_2616);
nor U3623 (N_3623,N_2444,N_2214);
nor U3624 (N_3624,N_2387,N_2581);
nor U3625 (N_3625,N_2895,N_2582);
nor U3626 (N_3626,N_2659,N_2017);
nand U3627 (N_3627,N_2652,N_2004);
or U3628 (N_3628,N_2832,N_2809);
xnor U3629 (N_3629,N_2178,N_2413);
xnor U3630 (N_3630,N_2612,N_2726);
and U3631 (N_3631,N_2155,N_2369);
and U3632 (N_3632,N_2358,N_2348);
nor U3633 (N_3633,N_2531,N_2067);
nand U3634 (N_3634,N_2116,N_2226);
nand U3635 (N_3635,N_2266,N_2437);
and U3636 (N_3636,N_2564,N_2333);
and U3637 (N_3637,N_2726,N_2372);
nand U3638 (N_3638,N_2960,N_2823);
xnor U3639 (N_3639,N_2810,N_2904);
nand U3640 (N_3640,N_2707,N_2886);
and U3641 (N_3641,N_2807,N_2698);
or U3642 (N_3642,N_2222,N_2080);
nor U3643 (N_3643,N_2716,N_2184);
and U3644 (N_3644,N_2767,N_2741);
and U3645 (N_3645,N_2804,N_2824);
xor U3646 (N_3646,N_2746,N_2674);
xnor U3647 (N_3647,N_2293,N_2277);
nand U3648 (N_3648,N_2441,N_2360);
nand U3649 (N_3649,N_2860,N_2635);
xnor U3650 (N_3650,N_2064,N_2251);
nor U3651 (N_3651,N_2148,N_2077);
xor U3652 (N_3652,N_2574,N_2929);
xnor U3653 (N_3653,N_2201,N_2907);
and U3654 (N_3654,N_2623,N_2541);
or U3655 (N_3655,N_2113,N_2060);
or U3656 (N_3656,N_2486,N_2260);
nor U3657 (N_3657,N_2577,N_2873);
and U3658 (N_3658,N_2623,N_2898);
and U3659 (N_3659,N_2346,N_2876);
nor U3660 (N_3660,N_2245,N_2465);
nand U3661 (N_3661,N_2885,N_2913);
or U3662 (N_3662,N_2856,N_2934);
nor U3663 (N_3663,N_2343,N_2523);
nand U3664 (N_3664,N_2848,N_2629);
nand U3665 (N_3665,N_2264,N_2701);
nor U3666 (N_3666,N_2195,N_2342);
nand U3667 (N_3667,N_2521,N_2161);
or U3668 (N_3668,N_2952,N_2576);
xnor U3669 (N_3669,N_2261,N_2109);
or U3670 (N_3670,N_2194,N_2435);
nand U3671 (N_3671,N_2087,N_2687);
xnor U3672 (N_3672,N_2682,N_2767);
and U3673 (N_3673,N_2172,N_2484);
nor U3674 (N_3674,N_2638,N_2181);
nor U3675 (N_3675,N_2817,N_2993);
nor U3676 (N_3676,N_2907,N_2835);
nand U3677 (N_3677,N_2896,N_2200);
and U3678 (N_3678,N_2935,N_2255);
nor U3679 (N_3679,N_2090,N_2030);
and U3680 (N_3680,N_2307,N_2440);
or U3681 (N_3681,N_2851,N_2134);
xor U3682 (N_3682,N_2972,N_2013);
nand U3683 (N_3683,N_2161,N_2609);
nor U3684 (N_3684,N_2599,N_2516);
nand U3685 (N_3685,N_2685,N_2734);
nor U3686 (N_3686,N_2528,N_2527);
xor U3687 (N_3687,N_2927,N_2572);
nand U3688 (N_3688,N_2687,N_2096);
or U3689 (N_3689,N_2569,N_2973);
or U3690 (N_3690,N_2785,N_2461);
and U3691 (N_3691,N_2024,N_2422);
or U3692 (N_3692,N_2997,N_2442);
nor U3693 (N_3693,N_2558,N_2773);
or U3694 (N_3694,N_2710,N_2219);
xnor U3695 (N_3695,N_2158,N_2167);
and U3696 (N_3696,N_2312,N_2343);
or U3697 (N_3697,N_2776,N_2656);
nor U3698 (N_3698,N_2767,N_2372);
nand U3699 (N_3699,N_2382,N_2232);
xnor U3700 (N_3700,N_2204,N_2056);
nor U3701 (N_3701,N_2269,N_2982);
xor U3702 (N_3702,N_2593,N_2519);
nand U3703 (N_3703,N_2872,N_2132);
nor U3704 (N_3704,N_2243,N_2886);
xor U3705 (N_3705,N_2102,N_2440);
or U3706 (N_3706,N_2635,N_2931);
or U3707 (N_3707,N_2368,N_2515);
or U3708 (N_3708,N_2033,N_2726);
nor U3709 (N_3709,N_2952,N_2406);
xnor U3710 (N_3710,N_2897,N_2823);
nand U3711 (N_3711,N_2081,N_2696);
or U3712 (N_3712,N_2362,N_2685);
nor U3713 (N_3713,N_2552,N_2488);
xnor U3714 (N_3714,N_2437,N_2509);
xor U3715 (N_3715,N_2775,N_2996);
nand U3716 (N_3716,N_2322,N_2079);
nand U3717 (N_3717,N_2976,N_2113);
and U3718 (N_3718,N_2281,N_2932);
nand U3719 (N_3719,N_2713,N_2033);
and U3720 (N_3720,N_2935,N_2981);
xnor U3721 (N_3721,N_2318,N_2637);
and U3722 (N_3722,N_2556,N_2559);
or U3723 (N_3723,N_2038,N_2745);
xnor U3724 (N_3724,N_2074,N_2195);
xor U3725 (N_3725,N_2474,N_2787);
or U3726 (N_3726,N_2263,N_2730);
or U3727 (N_3727,N_2826,N_2685);
xor U3728 (N_3728,N_2912,N_2833);
xor U3729 (N_3729,N_2205,N_2178);
and U3730 (N_3730,N_2768,N_2300);
nor U3731 (N_3731,N_2978,N_2501);
or U3732 (N_3732,N_2166,N_2024);
nor U3733 (N_3733,N_2214,N_2649);
xor U3734 (N_3734,N_2408,N_2742);
xnor U3735 (N_3735,N_2104,N_2997);
nor U3736 (N_3736,N_2472,N_2991);
nand U3737 (N_3737,N_2545,N_2756);
nand U3738 (N_3738,N_2598,N_2173);
or U3739 (N_3739,N_2838,N_2200);
nand U3740 (N_3740,N_2822,N_2330);
xor U3741 (N_3741,N_2463,N_2414);
or U3742 (N_3742,N_2737,N_2102);
and U3743 (N_3743,N_2118,N_2187);
xnor U3744 (N_3744,N_2350,N_2863);
or U3745 (N_3745,N_2964,N_2398);
nor U3746 (N_3746,N_2827,N_2931);
and U3747 (N_3747,N_2110,N_2114);
xor U3748 (N_3748,N_2184,N_2273);
nand U3749 (N_3749,N_2781,N_2732);
nor U3750 (N_3750,N_2119,N_2616);
xnor U3751 (N_3751,N_2459,N_2259);
xor U3752 (N_3752,N_2312,N_2589);
or U3753 (N_3753,N_2779,N_2534);
and U3754 (N_3754,N_2255,N_2004);
nor U3755 (N_3755,N_2891,N_2753);
and U3756 (N_3756,N_2751,N_2261);
nand U3757 (N_3757,N_2469,N_2716);
or U3758 (N_3758,N_2755,N_2948);
xnor U3759 (N_3759,N_2943,N_2459);
or U3760 (N_3760,N_2911,N_2314);
or U3761 (N_3761,N_2420,N_2141);
nor U3762 (N_3762,N_2649,N_2577);
nor U3763 (N_3763,N_2693,N_2909);
and U3764 (N_3764,N_2498,N_2780);
and U3765 (N_3765,N_2500,N_2985);
xor U3766 (N_3766,N_2440,N_2539);
or U3767 (N_3767,N_2551,N_2812);
nor U3768 (N_3768,N_2895,N_2074);
xor U3769 (N_3769,N_2401,N_2006);
nand U3770 (N_3770,N_2504,N_2172);
nor U3771 (N_3771,N_2222,N_2228);
xnor U3772 (N_3772,N_2544,N_2561);
or U3773 (N_3773,N_2686,N_2954);
xnor U3774 (N_3774,N_2998,N_2466);
and U3775 (N_3775,N_2684,N_2475);
xnor U3776 (N_3776,N_2005,N_2072);
xor U3777 (N_3777,N_2172,N_2364);
and U3778 (N_3778,N_2975,N_2156);
and U3779 (N_3779,N_2251,N_2111);
and U3780 (N_3780,N_2804,N_2964);
nand U3781 (N_3781,N_2889,N_2508);
or U3782 (N_3782,N_2936,N_2751);
nand U3783 (N_3783,N_2549,N_2645);
xnor U3784 (N_3784,N_2945,N_2435);
xor U3785 (N_3785,N_2710,N_2519);
xor U3786 (N_3786,N_2362,N_2727);
nor U3787 (N_3787,N_2938,N_2041);
and U3788 (N_3788,N_2802,N_2778);
and U3789 (N_3789,N_2814,N_2359);
nand U3790 (N_3790,N_2786,N_2846);
or U3791 (N_3791,N_2179,N_2445);
nor U3792 (N_3792,N_2728,N_2275);
nand U3793 (N_3793,N_2257,N_2736);
nor U3794 (N_3794,N_2352,N_2966);
or U3795 (N_3795,N_2807,N_2480);
and U3796 (N_3796,N_2856,N_2724);
or U3797 (N_3797,N_2857,N_2745);
and U3798 (N_3798,N_2700,N_2166);
or U3799 (N_3799,N_2686,N_2589);
nand U3800 (N_3800,N_2528,N_2942);
or U3801 (N_3801,N_2155,N_2120);
and U3802 (N_3802,N_2737,N_2880);
xnor U3803 (N_3803,N_2229,N_2978);
and U3804 (N_3804,N_2843,N_2424);
xnor U3805 (N_3805,N_2511,N_2165);
nand U3806 (N_3806,N_2020,N_2927);
xnor U3807 (N_3807,N_2821,N_2014);
nand U3808 (N_3808,N_2462,N_2970);
or U3809 (N_3809,N_2684,N_2757);
and U3810 (N_3810,N_2723,N_2821);
xnor U3811 (N_3811,N_2147,N_2285);
nor U3812 (N_3812,N_2624,N_2216);
xor U3813 (N_3813,N_2518,N_2410);
nor U3814 (N_3814,N_2684,N_2017);
nor U3815 (N_3815,N_2433,N_2095);
or U3816 (N_3816,N_2632,N_2393);
nor U3817 (N_3817,N_2194,N_2003);
or U3818 (N_3818,N_2993,N_2428);
nand U3819 (N_3819,N_2690,N_2169);
or U3820 (N_3820,N_2611,N_2122);
or U3821 (N_3821,N_2199,N_2029);
nor U3822 (N_3822,N_2040,N_2061);
nand U3823 (N_3823,N_2109,N_2892);
and U3824 (N_3824,N_2688,N_2380);
nand U3825 (N_3825,N_2232,N_2319);
nand U3826 (N_3826,N_2235,N_2252);
xor U3827 (N_3827,N_2608,N_2498);
xor U3828 (N_3828,N_2399,N_2702);
xor U3829 (N_3829,N_2712,N_2533);
nand U3830 (N_3830,N_2458,N_2612);
and U3831 (N_3831,N_2714,N_2735);
xnor U3832 (N_3832,N_2782,N_2593);
nor U3833 (N_3833,N_2103,N_2212);
nor U3834 (N_3834,N_2673,N_2175);
xor U3835 (N_3835,N_2251,N_2421);
and U3836 (N_3836,N_2526,N_2970);
nor U3837 (N_3837,N_2077,N_2494);
nand U3838 (N_3838,N_2468,N_2091);
nand U3839 (N_3839,N_2847,N_2885);
or U3840 (N_3840,N_2353,N_2312);
or U3841 (N_3841,N_2305,N_2828);
and U3842 (N_3842,N_2489,N_2039);
or U3843 (N_3843,N_2724,N_2525);
xnor U3844 (N_3844,N_2264,N_2989);
and U3845 (N_3845,N_2312,N_2108);
nor U3846 (N_3846,N_2357,N_2304);
nor U3847 (N_3847,N_2423,N_2912);
nor U3848 (N_3848,N_2121,N_2131);
or U3849 (N_3849,N_2380,N_2611);
nor U3850 (N_3850,N_2118,N_2491);
nor U3851 (N_3851,N_2622,N_2288);
nand U3852 (N_3852,N_2839,N_2710);
and U3853 (N_3853,N_2661,N_2852);
nand U3854 (N_3854,N_2413,N_2490);
or U3855 (N_3855,N_2932,N_2016);
nor U3856 (N_3856,N_2067,N_2234);
and U3857 (N_3857,N_2584,N_2738);
nor U3858 (N_3858,N_2485,N_2936);
nand U3859 (N_3859,N_2552,N_2105);
nor U3860 (N_3860,N_2981,N_2525);
and U3861 (N_3861,N_2308,N_2197);
or U3862 (N_3862,N_2154,N_2692);
and U3863 (N_3863,N_2667,N_2656);
xor U3864 (N_3864,N_2128,N_2937);
xor U3865 (N_3865,N_2611,N_2685);
or U3866 (N_3866,N_2784,N_2666);
and U3867 (N_3867,N_2134,N_2030);
or U3868 (N_3868,N_2515,N_2813);
and U3869 (N_3869,N_2634,N_2490);
and U3870 (N_3870,N_2929,N_2460);
and U3871 (N_3871,N_2544,N_2689);
nand U3872 (N_3872,N_2464,N_2835);
nor U3873 (N_3873,N_2796,N_2661);
nand U3874 (N_3874,N_2744,N_2120);
xor U3875 (N_3875,N_2698,N_2644);
or U3876 (N_3876,N_2960,N_2308);
or U3877 (N_3877,N_2532,N_2760);
xor U3878 (N_3878,N_2899,N_2796);
and U3879 (N_3879,N_2573,N_2225);
nor U3880 (N_3880,N_2787,N_2714);
nor U3881 (N_3881,N_2976,N_2310);
and U3882 (N_3882,N_2594,N_2545);
or U3883 (N_3883,N_2269,N_2624);
xnor U3884 (N_3884,N_2249,N_2023);
xnor U3885 (N_3885,N_2847,N_2195);
or U3886 (N_3886,N_2575,N_2796);
nor U3887 (N_3887,N_2280,N_2657);
nor U3888 (N_3888,N_2544,N_2629);
xor U3889 (N_3889,N_2959,N_2791);
nand U3890 (N_3890,N_2813,N_2822);
or U3891 (N_3891,N_2437,N_2604);
or U3892 (N_3892,N_2509,N_2179);
nor U3893 (N_3893,N_2789,N_2083);
xnor U3894 (N_3894,N_2684,N_2798);
or U3895 (N_3895,N_2073,N_2121);
or U3896 (N_3896,N_2462,N_2083);
or U3897 (N_3897,N_2057,N_2806);
nor U3898 (N_3898,N_2749,N_2283);
xor U3899 (N_3899,N_2757,N_2446);
nand U3900 (N_3900,N_2529,N_2969);
nand U3901 (N_3901,N_2622,N_2473);
xnor U3902 (N_3902,N_2092,N_2884);
and U3903 (N_3903,N_2095,N_2066);
nand U3904 (N_3904,N_2727,N_2170);
and U3905 (N_3905,N_2703,N_2966);
and U3906 (N_3906,N_2139,N_2299);
or U3907 (N_3907,N_2616,N_2377);
and U3908 (N_3908,N_2503,N_2124);
or U3909 (N_3909,N_2453,N_2744);
nor U3910 (N_3910,N_2239,N_2577);
and U3911 (N_3911,N_2042,N_2372);
nand U3912 (N_3912,N_2910,N_2933);
and U3913 (N_3913,N_2182,N_2356);
and U3914 (N_3914,N_2482,N_2048);
and U3915 (N_3915,N_2372,N_2635);
nand U3916 (N_3916,N_2362,N_2795);
nand U3917 (N_3917,N_2691,N_2778);
and U3918 (N_3918,N_2146,N_2961);
nand U3919 (N_3919,N_2839,N_2049);
nor U3920 (N_3920,N_2976,N_2049);
or U3921 (N_3921,N_2340,N_2874);
xnor U3922 (N_3922,N_2841,N_2437);
and U3923 (N_3923,N_2490,N_2089);
nor U3924 (N_3924,N_2532,N_2777);
nand U3925 (N_3925,N_2985,N_2626);
xor U3926 (N_3926,N_2565,N_2818);
and U3927 (N_3927,N_2592,N_2600);
or U3928 (N_3928,N_2124,N_2011);
xor U3929 (N_3929,N_2430,N_2600);
nor U3930 (N_3930,N_2995,N_2692);
nor U3931 (N_3931,N_2876,N_2503);
nand U3932 (N_3932,N_2918,N_2837);
or U3933 (N_3933,N_2736,N_2981);
nand U3934 (N_3934,N_2298,N_2778);
nand U3935 (N_3935,N_2527,N_2857);
xor U3936 (N_3936,N_2724,N_2972);
nand U3937 (N_3937,N_2432,N_2044);
xor U3938 (N_3938,N_2804,N_2458);
nor U3939 (N_3939,N_2257,N_2625);
or U3940 (N_3940,N_2823,N_2064);
and U3941 (N_3941,N_2998,N_2190);
or U3942 (N_3942,N_2127,N_2106);
and U3943 (N_3943,N_2903,N_2716);
or U3944 (N_3944,N_2345,N_2744);
nand U3945 (N_3945,N_2064,N_2461);
and U3946 (N_3946,N_2365,N_2457);
nand U3947 (N_3947,N_2862,N_2125);
xor U3948 (N_3948,N_2533,N_2093);
and U3949 (N_3949,N_2651,N_2454);
xor U3950 (N_3950,N_2587,N_2037);
and U3951 (N_3951,N_2796,N_2269);
xnor U3952 (N_3952,N_2645,N_2867);
and U3953 (N_3953,N_2679,N_2648);
xnor U3954 (N_3954,N_2227,N_2270);
or U3955 (N_3955,N_2048,N_2071);
and U3956 (N_3956,N_2643,N_2320);
nand U3957 (N_3957,N_2647,N_2718);
nor U3958 (N_3958,N_2241,N_2207);
xnor U3959 (N_3959,N_2478,N_2458);
nand U3960 (N_3960,N_2124,N_2276);
xor U3961 (N_3961,N_2987,N_2600);
xor U3962 (N_3962,N_2464,N_2798);
xnor U3963 (N_3963,N_2357,N_2015);
nor U3964 (N_3964,N_2841,N_2467);
and U3965 (N_3965,N_2165,N_2036);
or U3966 (N_3966,N_2097,N_2678);
nand U3967 (N_3967,N_2930,N_2012);
or U3968 (N_3968,N_2773,N_2153);
or U3969 (N_3969,N_2960,N_2524);
and U3970 (N_3970,N_2903,N_2374);
or U3971 (N_3971,N_2235,N_2223);
and U3972 (N_3972,N_2694,N_2700);
nand U3973 (N_3973,N_2781,N_2774);
nand U3974 (N_3974,N_2432,N_2620);
xnor U3975 (N_3975,N_2979,N_2610);
nand U3976 (N_3976,N_2750,N_2464);
xnor U3977 (N_3977,N_2282,N_2178);
nor U3978 (N_3978,N_2103,N_2465);
and U3979 (N_3979,N_2458,N_2764);
nand U3980 (N_3980,N_2289,N_2915);
or U3981 (N_3981,N_2266,N_2554);
and U3982 (N_3982,N_2150,N_2556);
or U3983 (N_3983,N_2619,N_2983);
nand U3984 (N_3984,N_2654,N_2722);
nand U3985 (N_3985,N_2090,N_2991);
and U3986 (N_3986,N_2627,N_2251);
or U3987 (N_3987,N_2247,N_2144);
nand U3988 (N_3988,N_2199,N_2140);
or U3989 (N_3989,N_2198,N_2556);
xnor U3990 (N_3990,N_2182,N_2868);
nand U3991 (N_3991,N_2613,N_2283);
and U3992 (N_3992,N_2892,N_2262);
and U3993 (N_3993,N_2273,N_2951);
nand U3994 (N_3994,N_2843,N_2995);
and U3995 (N_3995,N_2789,N_2905);
or U3996 (N_3996,N_2700,N_2915);
nor U3997 (N_3997,N_2140,N_2864);
and U3998 (N_3998,N_2935,N_2192);
or U3999 (N_3999,N_2120,N_2336);
or U4000 (N_4000,N_3791,N_3476);
or U4001 (N_4001,N_3351,N_3815);
xnor U4002 (N_4002,N_3172,N_3730);
or U4003 (N_4003,N_3054,N_3403);
or U4004 (N_4004,N_3915,N_3685);
or U4005 (N_4005,N_3038,N_3466);
nand U4006 (N_4006,N_3604,N_3629);
nand U4007 (N_4007,N_3439,N_3027);
nand U4008 (N_4008,N_3876,N_3931);
nor U4009 (N_4009,N_3602,N_3847);
or U4010 (N_4010,N_3621,N_3872);
nand U4011 (N_4011,N_3966,N_3643);
and U4012 (N_4012,N_3025,N_3248);
nor U4013 (N_4013,N_3456,N_3808);
and U4014 (N_4014,N_3222,N_3976);
nor U4015 (N_4015,N_3048,N_3180);
nand U4016 (N_4016,N_3593,N_3071);
xor U4017 (N_4017,N_3680,N_3686);
nor U4018 (N_4018,N_3672,N_3842);
or U4019 (N_4019,N_3990,N_3104);
or U4020 (N_4020,N_3015,N_3102);
or U4021 (N_4021,N_3851,N_3067);
xnor U4022 (N_4022,N_3312,N_3000);
nand U4023 (N_4023,N_3418,N_3070);
and U4024 (N_4024,N_3941,N_3215);
xor U4025 (N_4025,N_3368,N_3066);
and U4026 (N_4026,N_3261,N_3028);
nand U4027 (N_4027,N_3073,N_3463);
nor U4028 (N_4028,N_3665,N_3991);
and U4029 (N_4029,N_3989,N_3706);
and U4030 (N_4030,N_3677,N_3828);
and U4031 (N_4031,N_3378,N_3252);
nor U4032 (N_4032,N_3986,N_3412);
nor U4033 (N_4033,N_3764,N_3540);
or U4034 (N_4034,N_3265,N_3902);
xnor U4035 (N_4035,N_3831,N_3366);
nor U4036 (N_4036,N_3678,N_3575);
and U4037 (N_4037,N_3085,N_3447);
and U4038 (N_4038,N_3005,N_3820);
and U4039 (N_4039,N_3186,N_3794);
and U4040 (N_4040,N_3585,N_3910);
nand U4041 (N_4041,N_3218,N_3525);
nand U4042 (N_4042,N_3074,N_3957);
and U4043 (N_4043,N_3765,N_3532);
nand U4044 (N_4044,N_3722,N_3316);
nand U4045 (N_4045,N_3635,N_3410);
and U4046 (N_4046,N_3296,N_3736);
xnor U4047 (N_4047,N_3224,N_3938);
nor U4048 (N_4048,N_3922,N_3354);
nand U4049 (N_4049,N_3277,N_3996);
and U4050 (N_4050,N_3513,N_3987);
or U4051 (N_4051,N_3472,N_3026);
nand U4052 (N_4052,N_3813,N_3689);
xor U4053 (N_4053,N_3504,N_3283);
xnor U4054 (N_4054,N_3272,N_3345);
nor U4055 (N_4055,N_3647,N_3414);
nor U4056 (N_4056,N_3519,N_3502);
nor U4057 (N_4057,N_3666,N_3599);
nand U4058 (N_4058,N_3276,N_3803);
and U4059 (N_4059,N_3759,N_3405);
and U4060 (N_4060,N_3959,N_3857);
xnor U4061 (N_4061,N_3006,N_3649);
nor U4062 (N_4062,N_3698,N_3386);
and U4063 (N_4063,N_3511,N_3162);
nor U4064 (N_4064,N_3630,N_3696);
or U4065 (N_4065,N_3520,N_3858);
nand U4066 (N_4066,N_3928,N_3233);
xor U4067 (N_4067,N_3792,N_3041);
or U4068 (N_4068,N_3595,N_3716);
nand U4069 (N_4069,N_3760,N_3578);
nor U4070 (N_4070,N_3369,N_3181);
or U4071 (N_4071,N_3388,N_3427);
and U4072 (N_4072,N_3691,N_3505);
nor U4073 (N_4073,N_3954,N_3302);
xnor U4074 (N_4074,N_3442,N_3622);
or U4075 (N_4075,N_3546,N_3245);
nor U4076 (N_4076,N_3583,N_3772);
xnor U4077 (N_4077,N_3281,N_3559);
xor U4078 (N_4078,N_3601,N_3538);
nor U4079 (N_4079,N_3790,N_3392);
and U4080 (N_4080,N_3165,N_3419);
nand U4081 (N_4081,N_3898,N_3873);
nor U4082 (N_4082,N_3499,N_3570);
nor U4083 (N_4083,N_3099,N_3079);
nand U4084 (N_4084,N_3637,N_3206);
xor U4085 (N_4085,N_3503,N_3133);
xor U4086 (N_4086,N_3752,N_3367);
nand U4087 (N_4087,N_3337,N_3607);
nor U4088 (N_4088,N_3269,N_3718);
nand U4089 (N_4089,N_3865,N_3664);
and U4090 (N_4090,N_3921,N_3747);
nor U4091 (N_4091,N_3982,N_3271);
nand U4092 (N_4092,N_3867,N_3154);
xnor U4093 (N_4093,N_3868,N_3690);
nand U4094 (N_4094,N_3527,N_3613);
nor U4095 (N_4095,N_3241,N_3783);
or U4096 (N_4096,N_3913,N_3125);
xnor U4097 (N_4097,N_3655,N_3217);
and U4098 (N_4098,N_3491,N_3209);
nand U4099 (N_4099,N_3662,N_3623);
xnor U4100 (N_4100,N_3160,N_3648);
and U4101 (N_4101,N_3156,N_3169);
nand U4102 (N_4102,N_3558,N_3237);
nand U4103 (N_4103,N_3116,N_3311);
or U4104 (N_4104,N_3045,N_3983);
nor U4105 (N_4105,N_3140,N_3018);
nor U4106 (N_4106,N_3817,N_3906);
nand U4107 (N_4107,N_3106,N_3756);
xnor U4108 (N_4108,N_3979,N_3053);
nand U4109 (N_4109,N_3138,N_3549);
or U4110 (N_4110,N_3565,N_3158);
nor U4111 (N_4111,N_3397,N_3946);
nor U4112 (N_4112,N_3908,N_3839);
nand U4113 (N_4113,N_3200,N_3609);
nand U4114 (N_4114,N_3615,N_3874);
nand U4115 (N_4115,N_3901,N_3882);
or U4116 (N_4116,N_3614,N_3624);
nand U4117 (N_4117,N_3961,N_3055);
or U4118 (N_4118,N_3278,N_3192);
xnor U4119 (N_4119,N_3379,N_3807);
xor U4120 (N_4120,N_3596,N_3660);
and U4121 (N_4121,N_3458,N_3349);
or U4122 (N_4122,N_3744,N_3346);
and U4123 (N_4123,N_3232,N_3030);
and U4124 (N_4124,N_3632,N_3462);
and U4125 (N_4125,N_3560,N_3421);
xor U4126 (N_4126,N_3460,N_3425);
xnor U4127 (N_4127,N_3885,N_3268);
nor U4128 (N_4128,N_3471,N_3521);
and U4129 (N_4129,N_3658,N_3184);
xnor U4130 (N_4130,N_3295,N_3709);
nand U4131 (N_4131,N_3582,N_3951);
or U4132 (N_4132,N_3897,N_3016);
nand U4133 (N_4133,N_3358,N_3082);
and U4134 (N_4134,N_3947,N_3416);
and U4135 (N_4135,N_3309,N_3597);
nand U4136 (N_4136,N_3308,N_3667);
or U4137 (N_4137,N_3802,N_3211);
nor U4138 (N_4138,N_3299,N_3487);
nand U4139 (N_4139,N_3816,N_3275);
or U4140 (N_4140,N_3720,N_3919);
xnor U4141 (N_4141,N_3444,N_3088);
or U4142 (N_4142,N_3291,N_3288);
nand U4143 (N_4143,N_3574,N_3687);
and U4144 (N_4144,N_3330,N_3579);
xnor U4145 (N_4145,N_3301,N_3924);
xor U4146 (N_4146,N_3568,N_3797);
nor U4147 (N_4147,N_3199,N_3547);
or U4148 (N_4148,N_3830,N_3773);
or U4149 (N_4149,N_3904,N_3262);
nor U4150 (N_4150,N_3167,N_3201);
nand U4151 (N_4151,N_3377,N_3250);
nand U4152 (N_4152,N_3229,N_3393);
or U4153 (N_4153,N_3004,N_3977);
xnor U4154 (N_4154,N_3469,N_3284);
and U4155 (N_4155,N_3436,N_3255);
nand U4156 (N_4156,N_3327,N_3374);
xnor U4157 (N_4157,N_3282,N_3900);
nand U4158 (N_4158,N_3431,N_3130);
or U4159 (N_4159,N_3888,N_3370);
or U4160 (N_4160,N_3193,N_3395);
and U4161 (N_4161,N_3213,N_3178);
nor U4162 (N_4162,N_3091,N_3702);
nand U4163 (N_4163,N_3955,N_3812);
nor U4164 (N_4164,N_3932,N_3605);
or U4165 (N_4165,N_3577,N_3497);
nor U4166 (N_4166,N_3714,N_3770);
xor U4167 (N_4167,N_3408,N_3117);
nor U4168 (N_4168,N_3474,N_3246);
or U4169 (N_4169,N_3749,N_3539);
xor U4170 (N_4170,N_3611,N_3226);
nor U4171 (N_4171,N_3550,N_3486);
and U4172 (N_4172,N_3884,N_3183);
xor U4173 (N_4173,N_3257,N_3925);
xor U4174 (N_4174,N_3653,N_3929);
or U4175 (N_4175,N_3953,N_3049);
and U4176 (N_4176,N_3533,N_3717);
nor U4177 (N_4177,N_3995,N_3542);
nor U4178 (N_4178,N_3318,N_3112);
xor U4179 (N_4179,N_3190,N_3185);
xnor U4180 (N_4180,N_3259,N_3132);
nand U4181 (N_4181,N_3965,N_3705);
nor U4182 (N_4182,N_3479,N_3103);
nand U4183 (N_4183,N_3153,N_3740);
nor U4184 (N_4184,N_3968,N_3887);
nor U4185 (N_4185,N_3774,N_3043);
and U4186 (N_4186,N_3422,N_3126);
or U4187 (N_4187,N_3177,N_3811);
nand U4188 (N_4188,N_3509,N_3506);
and U4189 (N_4189,N_3748,N_3173);
nand U4190 (N_4190,N_3974,N_3093);
nor U4191 (N_4191,N_3095,N_3789);
or U4192 (N_4192,N_3258,N_3600);
and U4193 (N_4193,N_3062,N_3659);
nor U4194 (N_4194,N_3610,N_3952);
nor U4195 (N_4195,N_3937,N_3734);
or U4196 (N_4196,N_3650,N_3762);
or U4197 (N_4197,N_3014,N_3775);
xor U4198 (N_4198,N_3451,N_3866);
and U4199 (N_4199,N_3267,N_3033);
nor U4200 (N_4200,N_3118,N_3700);
nor U4201 (N_4201,N_3371,N_3424);
nand U4202 (N_4202,N_3668,N_3052);
nand U4203 (N_4203,N_3478,N_3128);
xor U4204 (N_4204,N_3881,N_3473);
or U4205 (N_4205,N_3781,N_3287);
and U4206 (N_4206,N_3875,N_3776);
or U4207 (N_4207,N_3111,N_3676);
xnor U4208 (N_4208,N_3715,N_3712);
and U4209 (N_4209,N_3735,N_3244);
xor U4210 (N_4210,N_3844,N_3123);
and U4211 (N_4211,N_3013,N_3833);
xnor U4212 (N_4212,N_3068,N_3355);
and U4213 (N_4213,N_3544,N_3342);
xnor U4214 (N_4214,N_3840,N_3423);
or U4215 (N_4215,N_3090,N_3950);
nand U4216 (N_4216,N_3084,N_3654);
xnor U4217 (N_4217,N_3020,N_3120);
and U4218 (N_4218,N_3507,N_3510);
nand U4219 (N_4219,N_3806,N_3134);
nand U4220 (N_4220,N_3948,N_3795);
and U4221 (N_4221,N_3683,N_3394);
and U4222 (N_4222,N_3935,N_3854);
nor U4223 (N_4223,N_3305,N_3892);
nor U4224 (N_4224,N_3554,N_3303);
xor U4225 (N_4225,N_3530,N_3315);
nand U4226 (N_4226,N_3586,N_3646);
nor U4227 (N_4227,N_3127,N_3673);
xor U4228 (N_4228,N_3761,N_3352);
nor U4229 (N_4229,N_3981,N_3435);
or U4230 (N_4230,N_3149,N_3100);
nand U4231 (N_4231,N_3157,N_3603);
and U4232 (N_4232,N_3809,N_3307);
nor U4233 (N_4233,N_3823,N_3174);
and U4234 (N_4234,N_3306,N_3798);
and U4235 (N_4235,N_3835,N_3855);
nand U4236 (N_4236,N_3270,N_3264);
and U4237 (N_4237,N_3086,N_3779);
or U4238 (N_4238,N_3553,N_3001);
and U4239 (N_4239,N_3023,N_3861);
nand U4240 (N_4240,N_3956,N_3194);
nor U4241 (N_4241,N_3168,N_3407);
xnor U4242 (N_4242,N_3310,N_3485);
xnor U4243 (N_4243,N_3230,N_3555);
and U4244 (N_4244,N_3064,N_3286);
nor U4245 (N_4245,N_3640,N_3682);
xor U4246 (N_4246,N_3777,N_3385);
xnor U4247 (N_4247,N_3496,N_3707);
xor U4248 (N_4248,N_3383,N_3693);
and U4249 (N_4249,N_3348,N_3122);
xor U4250 (N_4250,N_3202,N_3638);
and U4251 (N_4251,N_3893,N_3606);
nand U4252 (N_4252,N_3446,N_3515);
nand U4253 (N_4253,N_3468,N_3273);
xor U4254 (N_4254,N_3988,N_3663);
and U4255 (N_4255,N_3899,N_3508);
nand U4256 (N_4256,N_3189,N_3007);
and U4257 (N_4257,N_3101,N_3300);
nand U4258 (N_4258,N_3022,N_3031);
nand U4259 (N_4259,N_3778,N_3978);
or U4260 (N_4260,N_3591,N_3060);
and U4261 (N_4261,N_3905,N_3588);
or U4262 (N_4262,N_3459,N_3853);
nor U4263 (N_4263,N_3290,N_3108);
xnor U4264 (N_4264,N_3482,N_3843);
nand U4265 (N_4265,N_3917,N_3896);
or U4266 (N_4266,N_3862,N_3821);
or U4267 (N_4267,N_3652,N_3280);
nor U4268 (N_4268,N_3399,N_3841);
and U4269 (N_4269,N_3389,N_3625);
or U4270 (N_4270,N_3390,N_3869);
nor U4271 (N_4271,N_3719,N_3512);
and U4272 (N_4272,N_3617,N_3836);
xnor U4273 (N_4273,N_3044,N_3498);
and U4274 (N_4274,N_3187,N_3518);
xnor U4275 (N_4275,N_3243,N_3036);
and U4276 (N_4276,N_3457,N_3175);
nand U4277 (N_4277,N_3782,N_3204);
xnor U4278 (N_4278,N_3256,N_3163);
or U4279 (N_4279,N_3531,N_3699);
nand U4280 (N_4280,N_3944,N_3263);
and U4281 (N_4281,N_3047,N_3235);
nand U4282 (N_4282,N_3238,N_3825);
nand U4283 (N_4283,N_3115,N_3801);
xnor U4284 (N_4284,N_3046,N_3590);
nor U4285 (N_4285,N_3159,N_3285);
nand U4286 (N_4286,N_3708,N_3037);
nor U4287 (N_4287,N_3384,N_3768);
xnor U4288 (N_4288,N_3753,N_3059);
and U4289 (N_4289,N_3751,N_3826);
and U4290 (N_4290,N_3434,N_3240);
xnor U4291 (N_4291,N_3490,N_3517);
xnor U4292 (N_4292,N_3837,N_3289);
xor U4293 (N_4293,N_3151,N_3894);
xor U4294 (N_4294,N_3065,N_3077);
nand U4295 (N_4295,N_3480,N_3694);
or U4296 (N_4296,N_3973,N_3526);
nand U4297 (N_4297,N_3985,N_3992);
or U4298 (N_4298,N_3196,N_3148);
or U4299 (N_4299,N_3972,N_3608);
or U4300 (N_4300,N_3092,N_3701);
or U4301 (N_4301,N_3721,N_3247);
nor U4302 (N_4302,N_3920,N_3804);
xor U4303 (N_4303,N_3710,N_3564);
or U4304 (N_4304,N_3338,N_3484);
nor U4305 (N_4305,N_3317,N_3143);
nand U4306 (N_4306,N_3771,N_3353);
or U4307 (N_4307,N_3832,N_3131);
nor U4308 (N_4308,N_3584,N_3819);
and U4309 (N_4309,N_3669,N_3347);
nand U4310 (N_4310,N_3642,N_3083);
xor U4311 (N_4311,N_3139,N_3713);
xnor U4312 (N_4312,N_3228,N_3332);
nand U4313 (N_4313,N_3380,N_3766);
nor U4314 (N_4314,N_3566,N_3911);
and U4315 (N_4315,N_3253,N_3936);
or U4316 (N_4316,N_3113,N_3877);
or U4317 (N_4317,N_3381,N_3814);
nand U4318 (N_4318,N_3061,N_3799);
xor U4319 (N_4319,N_3063,N_3207);
nand U4320 (N_4320,N_3145,N_3975);
xnor U4321 (N_4321,N_3333,N_3545);
or U4322 (N_4322,N_3889,N_3994);
nor U4323 (N_4323,N_3155,N_3003);
or U4324 (N_4324,N_3688,N_3440);
nor U4325 (N_4325,N_3227,N_3329);
and U4326 (N_4326,N_3428,N_3891);
nor U4327 (N_4327,N_3619,N_3800);
nand U4328 (N_4328,N_3930,N_3914);
nor U4329 (N_4329,N_3592,N_3171);
nand U4330 (N_4330,N_3949,N_3754);
nand U4331 (N_4331,N_3029,N_3012);
and U4332 (N_4332,N_3357,N_3081);
and U4333 (N_4333,N_3537,N_3274);
and U4334 (N_4334,N_3557,N_3021);
nor U4335 (N_4335,N_3058,N_3704);
xor U4336 (N_4336,N_3628,N_3633);
nand U4337 (N_4337,N_3890,N_3737);
and U4338 (N_4338,N_3960,N_3382);
nor U4339 (N_4339,N_3942,N_3860);
nor U4340 (N_4340,N_3725,N_3724);
and U4341 (N_4341,N_3136,N_3017);
nor U4342 (N_4342,N_3152,N_3109);
nand U4343 (N_4343,N_3684,N_3293);
nor U4344 (N_4344,N_3328,N_3089);
nand U4345 (N_4345,N_3135,N_3331);
nor U4346 (N_4346,N_3094,N_3675);
and U4347 (N_4347,N_3849,N_3846);
nand U4348 (N_4348,N_3144,N_3404);
or U4349 (N_4349,N_3529,N_3580);
and U4350 (N_4350,N_3406,N_3958);
xnor U4351 (N_4351,N_3341,N_3692);
nand U4352 (N_4352,N_3703,N_3326);
nor U4353 (N_4353,N_3373,N_3571);
and U4354 (N_4354,N_3411,N_3343);
and U4355 (N_4355,N_3645,N_3208);
nand U4356 (N_4356,N_3644,N_3522);
xnor U4357 (N_4357,N_3114,N_3572);
or U4358 (N_4358,N_3254,N_3481);
nor U4359 (N_4359,N_3344,N_3980);
xnor U4360 (N_4360,N_3695,N_3050);
nor U4361 (N_4361,N_3618,N_3780);
and U4362 (N_4362,N_3524,N_3733);
nand U4363 (N_4363,N_3119,N_3757);
xnor U4364 (N_4364,N_3438,N_3916);
or U4365 (N_4365,N_3137,N_3998);
nand U4366 (N_4366,N_3489,N_3923);
or U4367 (N_4367,N_3829,N_3032);
nand U4368 (N_4368,N_3969,N_3573);
or U4369 (N_4369,N_3594,N_3728);
and U4370 (N_4370,N_3445,N_3750);
nand U4371 (N_4371,N_3010,N_3039);
nand U4372 (N_4372,N_3477,N_3612);
or U4373 (N_4373,N_3964,N_3164);
and U4374 (N_4374,N_3170,N_3105);
nand U4375 (N_4375,N_3051,N_3926);
or U4376 (N_4376,N_3984,N_3726);
and U4377 (N_4377,N_3361,N_3219);
or U4378 (N_4378,N_3195,N_3651);
nor U4379 (N_4379,N_3784,N_3656);
xnor U4380 (N_4380,N_3587,N_3631);
nand U4381 (N_4381,N_3755,N_3729);
nand U4382 (N_4382,N_3501,N_3616);
or U4383 (N_4383,N_3743,N_3210);
and U4384 (N_4384,N_3516,N_3129);
or U4385 (N_4385,N_3786,N_3997);
nand U4386 (N_4386,N_3176,N_3731);
nand U4387 (N_4387,N_3671,N_3581);
nor U4388 (N_4388,N_3220,N_3339);
nor U4389 (N_4389,N_3417,N_3008);
nand U4390 (N_4390,N_3562,N_3034);
xnor U4391 (N_4391,N_3372,N_3805);
nand U4392 (N_4392,N_3075,N_3161);
xor U4393 (N_4393,N_3543,N_3249);
and U4394 (N_4394,N_3567,N_3824);
or U4395 (N_4395,N_3657,N_3465);
nand U4396 (N_4396,N_3767,N_3681);
or U4397 (N_4397,N_3727,N_3360);
or U4398 (N_4398,N_3294,N_3788);
nor U4399 (N_4399,N_3236,N_3551);
nand U4400 (N_4400,N_3298,N_3297);
and U4401 (N_4401,N_3069,N_3097);
xnor U4402 (N_4402,N_3182,N_3918);
xnor U4403 (N_4403,N_3963,N_3320);
xnor U4404 (N_4404,N_3493,N_3415);
or U4405 (N_4405,N_3970,N_3166);
or U4406 (N_4406,N_3437,N_3903);
nand U4407 (N_4407,N_3746,N_3711);
and U4408 (N_4408,N_3818,N_3321);
and U4409 (N_4409,N_3319,N_3124);
nor U4410 (N_4410,N_3535,N_3852);
nand U4411 (N_4411,N_3500,N_3895);
and U4412 (N_4412,N_3528,N_3314);
xor U4413 (N_4413,N_3912,N_3121);
or U4414 (N_4414,N_3212,N_3002);
nand U4415 (N_4415,N_3098,N_3534);
and U4416 (N_4416,N_3536,N_3433);
and U4417 (N_4417,N_3279,N_3464);
xnor U4418 (N_4418,N_3340,N_3461);
nor U4419 (N_4419,N_3492,N_3322);
and U4420 (N_4420,N_3864,N_3409);
nor U4421 (N_4421,N_3335,N_3494);
or U4422 (N_4422,N_3364,N_3198);
and U4423 (N_4423,N_3943,N_3455);
or U4424 (N_4424,N_3810,N_3110);
nor U4425 (N_4425,N_3880,N_3620);
nand U4426 (N_4426,N_3732,N_3639);
nor U4427 (N_4427,N_3879,N_3179);
nor U4428 (N_4428,N_3313,N_3871);
and U4429 (N_4429,N_3569,N_3292);
xor U4430 (N_4430,N_3376,N_3598);
nor U4431 (N_4431,N_3441,N_3999);
nand U4432 (N_4432,N_3769,N_3056);
xor U4433 (N_4433,N_3225,N_3350);
nand U4434 (N_4434,N_3362,N_3375);
and U4435 (N_4435,N_3334,N_3763);
nor U4436 (N_4436,N_3356,N_3907);
xnor U4437 (N_4437,N_3266,N_3856);
nand U4438 (N_4438,N_3679,N_3443);
or U4439 (N_4439,N_3723,N_3323);
nand U4440 (N_4440,N_3470,N_3787);
nand U4441 (N_4441,N_3514,N_3636);
or U4442 (N_4442,N_3214,N_3009);
xor U4443 (N_4443,N_3548,N_3739);
nand U4444 (N_4444,N_3216,N_3072);
nor U4445 (N_4445,N_3971,N_3838);
nor U4446 (N_4446,N_3231,N_3758);
xor U4447 (N_4447,N_3626,N_3845);
and U4448 (N_4448,N_3561,N_3848);
nand U4449 (N_4449,N_3042,N_3142);
xnor U4450 (N_4450,N_3391,N_3454);
xnor U4451 (N_4451,N_3429,N_3670);
xor U4452 (N_4452,N_3863,N_3745);
and U4453 (N_4453,N_3933,N_3398);
nor U4454 (N_4454,N_3413,N_3078);
nand U4455 (N_4455,N_3859,N_3822);
nand U4456 (N_4456,N_3934,N_3420);
or U4457 (N_4457,N_3107,N_3035);
and U4458 (N_4458,N_3827,N_3661);
and U4459 (N_4459,N_3742,N_3223);
xor U4460 (N_4460,N_3205,N_3495);
nor U4461 (N_4461,N_3239,N_3785);
nor U4462 (N_4462,N_3962,N_3304);
nand U4463 (N_4463,N_3945,N_3221);
or U4464 (N_4464,N_3426,N_3336);
xor U4465 (N_4465,N_3040,N_3191);
or U4466 (N_4466,N_3878,N_3401);
nor U4467 (N_4467,N_3641,N_3251);
or U4468 (N_4468,N_3448,N_3096);
and U4469 (N_4469,N_3576,N_3396);
nor U4470 (N_4470,N_3741,N_3365);
xnor U4471 (N_4471,N_3488,N_3467);
and U4472 (N_4472,N_3087,N_3674);
or U4473 (N_4473,N_3523,N_3150);
nand U4474 (N_4474,N_3197,N_3363);
nand U4475 (N_4475,N_3563,N_3738);
or U4476 (N_4476,N_3796,N_3634);
xor U4477 (N_4477,N_3483,N_3870);
nor U4478 (N_4478,N_3260,N_3402);
xor U4479 (N_4479,N_3057,N_3993);
xnor U4480 (N_4480,N_3541,N_3556);
nor U4481 (N_4481,N_3147,N_3387);
xnor U4482 (N_4482,N_3450,N_3432);
nand U4483 (N_4483,N_3011,N_3834);
nand U4484 (N_4484,N_3927,N_3400);
nor U4485 (N_4485,N_3203,N_3452);
nor U4486 (N_4486,N_3793,N_3453);
nor U4487 (N_4487,N_3234,N_3850);
and U4488 (N_4488,N_3627,N_3449);
nand U4489 (N_4489,N_3325,N_3188);
and U4490 (N_4490,N_3019,N_3024);
and U4491 (N_4491,N_3909,N_3967);
nand U4492 (N_4492,N_3080,N_3939);
nand U4493 (N_4493,N_3359,N_3940);
nand U4494 (N_4494,N_3697,N_3883);
or U4495 (N_4495,N_3886,N_3076);
nand U4496 (N_4496,N_3475,N_3430);
nand U4497 (N_4497,N_3324,N_3589);
and U4498 (N_4498,N_3552,N_3141);
or U4499 (N_4499,N_3242,N_3146);
and U4500 (N_4500,N_3370,N_3852);
nor U4501 (N_4501,N_3697,N_3885);
nand U4502 (N_4502,N_3727,N_3082);
or U4503 (N_4503,N_3757,N_3458);
and U4504 (N_4504,N_3525,N_3959);
nand U4505 (N_4505,N_3596,N_3673);
xor U4506 (N_4506,N_3590,N_3627);
nor U4507 (N_4507,N_3649,N_3095);
or U4508 (N_4508,N_3791,N_3562);
nor U4509 (N_4509,N_3694,N_3603);
and U4510 (N_4510,N_3540,N_3014);
nand U4511 (N_4511,N_3051,N_3095);
nand U4512 (N_4512,N_3697,N_3005);
xor U4513 (N_4513,N_3315,N_3324);
nor U4514 (N_4514,N_3172,N_3571);
and U4515 (N_4515,N_3627,N_3154);
nand U4516 (N_4516,N_3281,N_3629);
and U4517 (N_4517,N_3557,N_3006);
xnor U4518 (N_4518,N_3667,N_3791);
nor U4519 (N_4519,N_3247,N_3991);
xor U4520 (N_4520,N_3011,N_3582);
or U4521 (N_4521,N_3727,N_3681);
nand U4522 (N_4522,N_3698,N_3768);
and U4523 (N_4523,N_3224,N_3960);
and U4524 (N_4524,N_3122,N_3030);
and U4525 (N_4525,N_3162,N_3928);
or U4526 (N_4526,N_3603,N_3597);
nand U4527 (N_4527,N_3370,N_3893);
nand U4528 (N_4528,N_3876,N_3374);
nor U4529 (N_4529,N_3721,N_3444);
and U4530 (N_4530,N_3733,N_3910);
nand U4531 (N_4531,N_3728,N_3206);
xnor U4532 (N_4532,N_3756,N_3337);
nand U4533 (N_4533,N_3392,N_3999);
nor U4534 (N_4534,N_3873,N_3986);
nand U4535 (N_4535,N_3824,N_3248);
and U4536 (N_4536,N_3041,N_3117);
xnor U4537 (N_4537,N_3272,N_3577);
and U4538 (N_4538,N_3525,N_3988);
and U4539 (N_4539,N_3483,N_3554);
nand U4540 (N_4540,N_3595,N_3020);
and U4541 (N_4541,N_3969,N_3078);
or U4542 (N_4542,N_3613,N_3628);
nor U4543 (N_4543,N_3703,N_3243);
nor U4544 (N_4544,N_3449,N_3307);
or U4545 (N_4545,N_3279,N_3912);
nand U4546 (N_4546,N_3187,N_3614);
nand U4547 (N_4547,N_3862,N_3263);
or U4548 (N_4548,N_3215,N_3915);
xnor U4549 (N_4549,N_3101,N_3281);
and U4550 (N_4550,N_3527,N_3562);
or U4551 (N_4551,N_3288,N_3238);
nand U4552 (N_4552,N_3496,N_3791);
nand U4553 (N_4553,N_3520,N_3011);
and U4554 (N_4554,N_3984,N_3399);
or U4555 (N_4555,N_3406,N_3934);
nor U4556 (N_4556,N_3684,N_3876);
nand U4557 (N_4557,N_3657,N_3250);
nor U4558 (N_4558,N_3796,N_3567);
nor U4559 (N_4559,N_3499,N_3299);
nand U4560 (N_4560,N_3044,N_3613);
nand U4561 (N_4561,N_3629,N_3588);
or U4562 (N_4562,N_3160,N_3453);
nand U4563 (N_4563,N_3341,N_3359);
and U4564 (N_4564,N_3507,N_3393);
or U4565 (N_4565,N_3257,N_3305);
nand U4566 (N_4566,N_3229,N_3614);
nor U4567 (N_4567,N_3799,N_3820);
xor U4568 (N_4568,N_3979,N_3165);
or U4569 (N_4569,N_3900,N_3703);
nand U4570 (N_4570,N_3316,N_3947);
nand U4571 (N_4571,N_3420,N_3433);
nor U4572 (N_4572,N_3203,N_3786);
or U4573 (N_4573,N_3514,N_3886);
or U4574 (N_4574,N_3630,N_3381);
nand U4575 (N_4575,N_3732,N_3841);
nand U4576 (N_4576,N_3662,N_3505);
nand U4577 (N_4577,N_3100,N_3853);
nand U4578 (N_4578,N_3651,N_3206);
and U4579 (N_4579,N_3816,N_3959);
nor U4580 (N_4580,N_3714,N_3348);
or U4581 (N_4581,N_3313,N_3144);
xor U4582 (N_4582,N_3090,N_3994);
or U4583 (N_4583,N_3129,N_3606);
nand U4584 (N_4584,N_3210,N_3438);
nor U4585 (N_4585,N_3953,N_3352);
and U4586 (N_4586,N_3841,N_3686);
nand U4587 (N_4587,N_3841,N_3989);
nor U4588 (N_4588,N_3792,N_3934);
or U4589 (N_4589,N_3548,N_3125);
nor U4590 (N_4590,N_3239,N_3936);
nor U4591 (N_4591,N_3509,N_3649);
nand U4592 (N_4592,N_3851,N_3799);
and U4593 (N_4593,N_3352,N_3402);
nor U4594 (N_4594,N_3063,N_3951);
nand U4595 (N_4595,N_3316,N_3699);
xor U4596 (N_4596,N_3816,N_3839);
and U4597 (N_4597,N_3743,N_3957);
or U4598 (N_4598,N_3326,N_3607);
or U4599 (N_4599,N_3207,N_3162);
nand U4600 (N_4600,N_3265,N_3779);
and U4601 (N_4601,N_3836,N_3929);
nand U4602 (N_4602,N_3029,N_3515);
nor U4603 (N_4603,N_3055,N_3583);
xnor U4604 (N_4604,N_3914,N_3131);
or U4605 (N_4605,N_3576,N_3005);
or U4606 (N_4606,N_3574,N_3334);
xor U4607 (N_4607,N_3654,N_3301);
nand U4608 (N_4608,N_3249,N_3149);
or U4609 (N_4609,N_3215,N_3400);
nand U4610 (N_4610,N_3905,N_3257);
xor U4611 (N_4611,N_3355,N_3772);
xnor U4612 (N_4612,N_3991,N_3500);
nor U4613 (N_4613,N_3907,N_3930);
and U4614 (N_4614,N_3209,N_3871);
or U4615 (N_4615,N_3535,N_3709);
nor U4616 (N_4616,N_3112,N_3764);
nand U4617 (N_4617,N_3928,N_3575);
and U4618 (N_4618,N_3123,N_3368);
xnor U4619 (N_4619,N_3214,N_3754);
and U4620 (N_4620,N_3508,N_3047);
xor U4621 (N_4621,N_3322,N_3317);
and U4622 (N_4622,N_3514,N_3600);
and U4623 (N_4623,N_3322,N_3037);
nand U4624 (N_4624,N_3747,N_3157);
and U4625 (N_4625,N_3180,N_3389);
and U4626 (N_4626,N_3105,N_3681);
nor U4627 (N_4627,N_3286,N_3029);
nand U4628 (N_4628,N_3946,N_3652);
and U4629 (N_4629,N_3642,N_3370);
xnor U4630 (N_4630,N_3210,N_3037);
and U4631 (N_4631,N_3236,N_3843);
or U4632 (N_4632,N_3941,N_3625);
and U4633 (N_4633,N_3721,N_3179);
xor U4634 (N_4634,N_3203,N_3958);
nand U4635 (N_4635,N_3807,N_3698);
or U4636 (N_4636,N_3990,N_3055);
nor U4637 (N_4637,N_3453,N_3948);
or U4638 (N_4638,N_3738,N_3106);
xnor U4639 (N_4639,N_3940,N_3307);
nor U4640 (N_4640,N_3539,N_3756);
and U4641 (N_4641,N_3252,N_3152);
nor U4642 (N_4642,N_3765,N_3565);
nand U4643 (N_4643,N_3342,N_3078);
or U4644 (N_4644,N_3030,N_3515);
or U4645 (N_4645,N_3779,N_3414);
or U4646 (N_4646,N_3590,N_3049);
xor U4647 (N_4647,N_3915,N_3232);
nor U4648 (N_4648,N_3517,N_3140);
nor U4649 (N_4649,N_3455,N_3731);
xor U4650 (N_4650,N_3033,N_3571);
nand U4651 (N_4651,N_3266,N_3833);
and U4652 (N_4652,N_3720,N_3119);
nor U4653 (N_4653,N_3672,N_3196);
nor U4654 (N_4654,N_3910,N_3638);
nor U4655 (N_4655,N_3306,N_3933);
nor U4656 (N_4656,N_3049,N_3673);
or U4657 (N_4657,N_3542,N_3080);
or U4658 (N_4658,N_3336,N_3834);
and U4659 (N_4659,N_3615,N_3305);
nor U4660 (N_4660,N_3607,N_3275);
and U4661 (N_4661,N_3293,N_3736);
or U4662 (N_4662,N_3406,N_3589);
and U4663 (N_4663,N_3951,N_3744);
or U4664 (N_4664,N_3777,N_3276);
or U4665 (N_4665,N_3927,N_3864);
or U4666 (N_4666,N_3521,N_3414);
xor U4667 (N_4667,N_3395,N_3003);
nor U4668 (N_4668,N_3048,N_3457);
xnor U4669 (N_4669,N_3402,N_3238);
xor U4670 (N_4670,N_3121,N_3017);
and U4671 (N_4671,N_3488,N_3276);
or U4672 (N_4672,N_3331,N_3549);
xnor U4673 (N_4673,N_3648,N_3058);
or U4674 (N_4674,N_3689,N_3864);
or U4675 (N_4675,N_3159,N_3265);
and U4676 (N_4676,N_3189,N_3531);
xor U4677 (N_4677,N_3251,N_3564);
nand U4678 (N_4678,N_3818,N_3416);
or U4679 (N_4679,N_3725,N_3642);
xnor U4680 (N_4680,N_3342,N_3827);
or U4681 (N_4681,N_3299,N_3767);
xnor U4682 (N_4682,N_3181,N_3630);
xor U4683 (N_4683,N_3374,N_3204);
nor U4684 (N_4684,N_3778,N_3719);
xor U4685 (N_4685,N_3468,N_3116);
and U4686 (N_4686,N_3634,N_3239);
nor U4687 (N_4687,N_3871,N_3675);
or U4688 (N_4688,N_3065,N_3555);
nor U4689 (N_4689,N_3508,N_3726);
and U4690 (N_4690,N_3800,N_3325);
or U4691 (N_4691,N_3374,N_3469);
and U4692 (N_4692,N_3316,N_3291);
and U4693 (N_4693,N_3111,N_3268);
and U4694 (N_4694,N_3262,N_3096);
xnor U4695 (N_4695,N_3953,N_3906);
xnor U4696 (N_4696,N_3684,N_3441);
or U4697 (N_4697,N_3234,N_3105);
nand U4698 (N_4698,N_3628,N_3215);
xor U4699 (N_4699,N_3524,N_3365);
and U4700 (N_4700,N_3632,N_3148);
nor U4701 (N_4701,N_3916,N_3587);
nor U4702 (N_4702,N_3722,N_3634);
nor U4703 (N_4703,N_3880,N_3452);
and U4704 (N_4704,N_3184,N_3255);
xor U4705 (N_4705,N_3518,N_3533);
nor U4706 (N_4706,N_3977,N_3525);
nand U4707 (N_4707,N_3088,N_3496);
and U4708 (N_4708,N_3063,N_3285);
nor U4709 (N_4709,N_3253,N_3597);
and U4710 (N_4710,N_3144,N_3176);
nand U4711 (N_4711,N_3964,N_3366);
xnor U4712 (N_4712,N_3007,N_3058);
and U4713 (N_4713,N_3625,N_3587);
and U4714 (N_4714,N_3272,N_3232);
and U4715 (N_4715,N_3222,N_3615);
xor U4716 (N_4716,N_3535,N_3826);
and U4717 (N_4717,N_3042,N_3442);
and U4718 (N_4718,N_3329,N_3673);
nor U4719 (N_4719,N_3222,N_3183);
nand U4720 (N_4720,N_3891,N_3676);
and U4721 (N_4721,N_3541,N_3633);
xor U4722 (N_4722,N_3362,N_3395);
xor U4723 (N_4723,N_3779,N_3433);
or U4724 (N_4724,N_3449,N_3229);
or U4725 (N_4725,N_3999,N_3888);
xor U4726 (N_4726,N_3868,N_3160);
and U4727 (N_4727,N_3497,N_3399);
and U4728 (N_4728,N_3745,N_3151);
nor U4729 (N_4729,N_3969,N_3201);
nor U4730 (N_4730,N_3568,N_3116);
or U4731 (N_4731,N_3367,N_3017);
or U4732 (N_4732,N_3161,N_3235);
or U4733 (N_4733,N_3192,N_3778);
xnor U4734 (N_4734,N_3303,N_3381);
and U4735 (N_4735,N_3284,N_3506);
or U4736 (N_4736,N_3162,N_3580);
or U4737 (N_4737,N_3260,N_3886);
nor U4738 (N_4738,N_3744,N_3961);
nor U4739 (N_4739,N_3999,N_3477);
nand U4740 (N_4740,N_3043,N_3328);
nor U4741 (N_4741,N_3987,N_3936);
or U4742 (N_4742,N_3545,N_3944);
xnor U4743 (N_4743,N_3470,N_3772);
nand U4744 (N_4744,N_3106,N_3056);
and U4745 (N_4745,N_3809,N_3325);
or U4746 (N_4746,N_3772,N_3050);
nand U4747 (N_4747,N_3961,N_3906);
xnor U4748 (N_4748,N_3346,N_3767);
or U4749 (N_4749,N_3403,N_3025);
xor U4750 (N_4750,N_3791,N_3932);
nor U4751 (N_4751,N_3733,N_3094);
xor U4752 (N_4752,N_3214,N_3016);
nor U4753 (N_4753,N_3303,N_3220);
nand U4754 (N_4754,N_3400,N_3031);
nor U4755 (N_4755,N_3342,N_3525);
and U4756 (N_4756,N_3736,N_3916);
nand U4757 (N_4757,N_3331,N_3694);
or U4758 (N_4758,N_3384,N_3032);
nor U4759 (N_4759,N_3387,N_3447);
nand U4760 (N_4760,N_3509,N_3188);
nor U4761 (N_4761,N_3433,N_3084);
nor U4762 (N_4762,N_3226,N_3222);
xnor U4763 (N_4763,N_3761,N_3479);
or U4764 (N_4764,N_3496,N_3918);
nor U4765 (N_4765,N_3391,N_3801);
nor U4766 (N_4766,N_3710,N_3015);
nor U4767 (N_4767,N_3957,N_3362);
nor U4768 (N_4768,N_3066,N_3547);
and U4769 (N_4769,N_3134,N_3135);
xnor U4770 (N_4770,N_3548,N_3885);
xor U4771 (N_4771,N_3712,N_3288);
nand U4772 (N_4772,N_3819,N_3269);
and U4773 (N_4773,N_3967,N_3223);
nor U4774 (N_4774,N_3967,N_3352);
and U4775 (N_4775,N_3938,N_3720);
or U4776 (N_4776,N_3792,N_3499);
nor U4777 (N_4777,N_3346,N_3247);
and U4778 (N_4778,N_3489,N_3456);
nor U4779 (N_4779,N_3237,N_3231);
xnor U4780 (N_4780,N_3052,N_3911);
nand U4781 (N_4781,N_3889,N_3018);
nor U4782 (N_4782,N_3448,N_3708);
or U4783 (N_4783,N_3689,N_3047);
or U4784 (N_4784,N_3128,N_3415);
and U4785 (N_4785,N_3216,N_3117);
nand U4786 (N_4786,N_3380,N_3239);
nor U4787 (N_4787,N_3529,N_3095);
xor U4788 (N_4788,N_3604,N_3452);
and U4789 (N_4789,N_3570,N_3835);
xnor U4790 (N_4790,N_3438,N_3897);
xor U4791 (N_4791,N_3506,N_3058);
or U4792 (N_4792,N_3736,N_3013);
or U4793 (N_4793,N_3778,N_3620);
and U4794 (N_4794,N_3298,N_3885);
nand U4795 (N_4795,N_3383,N_3662);
or U4796 (N_4796,N_3448,N_3250);
nand U4797 (N_4797,N_3202,N_3712);
xnor U4798 (N_4798,N_3408,N_3480);
nor U4799 (N_4799,N_3491,N_3102);
or U4800 (N_4800,N_3702,N_3258);
or U4801 (N_4801,N_3011,N_3766);
and U4802 (N_4802,N_3826,N_3600);
xor U4803 (N_4803,N_3468,N_3790);
xor U4804 (N_4804,N_3161,N_3799);
or U4805 (N_4805,N_3113,N_3043);
xor U4806 (N_4806,N_3842,N_3085);
and U4807 (N_4807,N_3223,N_3851);
xnor U4808 (N_4808,N_3667,N_3995);
nor U4809 (N_4809,N_3403,N_3757);
or U4810 (N_4810,N_3464,N_3938);
xor U4811 (N_4811,N_3999,N_3502);
xor U4812 (N_4812,N_3053,N_3688);
nor U4813 (N_4813,N_3332,N_3779);
nand U4814 (N_4814,N_3818,N_3291);
xnor U4815 (N_4815,N_3292,N_3600);
nor U4816 (N_4816,N_3246,N_3457);
and U4817 (N_4817,N_3335,N_3665);
or U4818 (N_4818,N_3966,N_3240);
nand U4819 (N_4819,N_3057,N_3947);
and U4820 (N_4820,N_3975,N_3853);
and U4821 (N_4821,N_3407,N_3249);
nand U4822 (N_4822,N_3542,N_3126);
or U4823 (N_4823,N_3414,N_3731);
nor U4824 (N_4824,N_3051,N_3613);
nor U4825 (N_4825,N_3486,N_3928);
xor U4826 (N_4826,N_3561,N_3287);
nor U4827 (N_4827,N_3861,N_3578);
or U4828 (N_4828,N_3255,N_3732);
xnor U4829 (N_4829,N_3037,N_3713);
nor U4830 (N_4830,N_3266,N_3443);
or U4831 (N_4831,N_3573,N_3401);
and U4832 (N_4832,N_3647,N_3843);
xnor U4833 (N_4833,N_3224,N_3119);
nor U4834 (N_4834,N_3469,N_3147);
and U4835 (N_4835,N_3661,N_3458);
and U4836 (N_4836,N_3227,N_3152);
nor U4837 (N_4837,N_3840,N_3160);
and U4838 (N_4838,N_3128,N_3606);
xor U4839 (N_4839,N_3790,N_3512);
or U4840 (N_4840,N_3428,N_3934);
or U4841 (N_4841,N_3186,N_3993);
or U4842 (N_4842,N_3643,N_3829);
and U4843 (N_4843,N_3177,N_3157);
xor U4844 (N_4844,N_3529,N_3409);
nor U4845 (N_4845,N_3874,N_3633);
or U4846 (N_4846,N_3841,N_3906);
nand U4847 (N_4847,N_3268,N_3076);
xor U4848 (N_4848,N_3337,N_3887);
or U4849 (N_4849,N_3096,N_3590);
and U4850 (N_4850,N_3490,N_3599);
xnor U4851 (N_4851,N_3127,N_3730);
nand U4852 (N_4852,N_3099,N_3808);
nand U4853 (N_4853,N_3632,N_3723);
and U4854 (N_4854,N_3159,N_3301);
xor U4855 (N_4855,N_3533,N_3596);
xnor U4856 (N_4856,N_3456,N_3244);
or U4857 (N_4857,N_3504,N_3747);
or U4858 (N_4858,N_3434,N_3271);
xor U4859 (N_4859,N_3104,N_3212);
nor U4860 (N_4860,N_3014,N_3597);
or U4861 (N_4861,N_3621,N_3632);
or U4862 (N_4862,N_3546,N_3293);
xnor U4863 (N_4863,N_3126,N_3944);
and U4864 (N_4864,N_3243,N_3565);
xnor U4865 (N_4865,N_3725,N_3390);
nor U4866 (N_4866,N_3702,N_3132);
nand U4867 (N_4867,N_3230,N_3436);
or U4868 (N_4868,N_3844,N_3745);
xor U4869 (N_4869,N_3985,N_3748);
and U4870 (N_4870,N_3620,N_3394);
and U4871 (N_4871,N_3533,N_3806);
or U4872 (N_4872,N_3626,N_3449);
nand U4873 (N_4873,N_3433,N_3663);
or U4874 (N_4874,N_3268,N_3663);
xnor U4875 (N_4875,N_3521,N_3849);
xnor U4876 (N_4876,N_3845,N_3740);
nor U4877 (N_4877,N_3998,N_3443);
and U4878 (N_4878,N_3763,N_3690);
nand U4879 (N_4879,N_3149,N_3225);
and U4880 (N_4880,N_3258,N_3620);
xor U4881 (N_4881,N_3763,N_3817);
and U4882 (N_4882,N_3830,N_3377);
nand U4883 (N_4883,N_3972,N_3103);
xor U4884 (N_4884,N_3797,N_3526);
and U4885 (N_4885,N_3282,N_3846);
nor U4886 (N_4886,N_3775,N_3904);
and U4887 (N_4887,N_3596,N_3997);
nand U4888 (N_4888,N_3244,N_3882);
nand U4889 (N_4889,N_3598,N_3036);
and U4890 (N_4890,N_3026,N_3606);
xnor U4891 (N_4891,N_3518,N_3064);
and U4892 (N_4892,N_3559,N_3042);
nand U4893 (N_4893,N_3443,N_3873);
xnor U4894 (N_4894,N_3671,N_3437);
nand U4895 (N_4895,N_3079,N_3569);
nand U4896 (N_4896,N_3931,N_3499);
or U4897 (N_4897,N_3968,N_3326);
xor U4898 (N_4898,N_3173,N_3878);
or U4899 (N_4899,N_3704,N_3398);
and U4900 (N_4900,N_3201,N_3774);
and U4901 (N_4901,N_3960,N_3770);
xnor U4902 (N_4902,N_3573,N_3645);
and U4903 (N_4903,N_3275,N_3196);
or U4904 (N_4904,N_3339,N_3465);
nor U4905 (N_4905,N_3963,N_3360);
and U4906 (N_4906,N_3811,N_3693);
nand U4907 (N_4907,N_3890,N_3464);
nand U4908 (N_4908,N_3172,N_3839);
and U4909 (N_4909,N_3163,N_3001);
or U4910 (N_4910,N_3465,N_3590);
nor U4911 (N_4911,N_3672,N_3511);
and U4912 (N_4912,N_3089,N_3207);
and U4913 (N_4913,N_3560,N_3918);
or U4914 (N_4914,N_3184,N_3997);
and U4915 (N_4915,N_3442,N_3736);
nor U4916 (N_4916,N_3794,N_3702);
and U4917 (N_4917,N_3722,N_3565);
nand U4918 (N_4918,N_3792,N_3065);
and U4919 (N_4919,N_3243,N_3580);
xnor U4920 (N_4920,N_3775,N_3257);
and U4921 (N_4921,N_3597,N_3909);
or U4922 (N_4922,N_3110,N_3821);
and U4923 (N_4923,N_3946,N_3284);
and U4924 (N_4924,N_3679,N_3242);
xor U4925 (N_4925,N_3231,N_3789);
nor U4926 (N_4926,N_3916,N_3194);
nor U4927 (N_4927,N_3468,N_3010);
and U4928 (N_4928,N_3600,N_3218);
and U4929 (N_4929,N_3219,N_3964);
and U4930 (N_4930,N_3010,N_3429);
xor U4931 (N_4931,N_3595,N_3875);
or U4932 (N_4932,N_3293,N_3261);
nor U4933 (N_4933,N_3741,N_3450);
xor U4934 (N_4934,N_3126,N_3678);
and U4935 (N_4935,N_3093,N_3626);
and U4936 (N_4936,N_3062,N_3795);
and U4937 (N_4937,N_3912,N_3914);
and U4938 (N_4938,N_3163,N_3167);
or U4939 (N_4939,N_3333,N_3445);
or U4940 (N_4940,N_3103,N_3141);
or U4941 (N_4941,N_3047,N_3052);
and U4942 (N_4942,N_3407,N_3441);
nand U4943 (N_4943,N_3695,N_3029);
nor U4944 (N_4944,N_3900,N_3080);
nor U4945 (N_4945,N_3084,N_3026);
and U4946 (N_4946,N_3807,N_3131);
nor U4947 (N_4947,N_3733,N_3975);
or U4948 (N_4948,N_3911,N_3557);
nand U4949 (N_4949,N_3804,N_3796);
and U4950 (N_4950,N_3562,N_3895);
nand U4951 (N_4951,N_3794,N_3052);
xnor U4952 (N_4952,N_3445,N_3193);
nor U4953 (N_4953,N_3918,N_3574);
or U4954 (N_4954,N_3945,N_3394);
nor U4955 (N_4955,N_3471,N_3879);
or U4956 (N_4956,N_3636,N_3188);
or U4957 (N_4957,N_3146,N_3876);
nor U4958 (N_4958,N_3883,N_3209);
or U4959 (N_4959,N_3009,N_3040);
and U4960 (N_4960,N_3215,N_3547);
and U4961 (N_4961,N_3846,N_3640);
or U4962 (N_4962,N_3987,N_3220);
xnor U4963 (N_4963,N_3771,N_3003);
nor U4964 (N_4964,N_3408,N_3018);
or U4965 (N_4965,N_3298,N_3671);
xor U4966 (N_4966,N_3369,N_3436);
or U4967 (N_4967,N_3320,N_3172);
nor U4968 (N_4968,N_3302,N_3419);
or U4969 (N_4969,N_3566,N_3228);
nor U4970 (N_4970,N_3566,N_3309);
or U4971 (N_4971,N_3989,N_3058);
or U4972 (N_4972,N_3501,N_3665);
nand U4973 (N_4973,N_3068,N_3985);
or U4974 (N_4974,N_3288,N_3465);
nand U4975 (N_4975,N_3511,N_3782);
nor U4976 (N_4976,N_3620,N_3798);
nand U4977 (N_4977,N_3347,N_3071);
or U4978 (N_4978,N_3623,N_3256);
and U4979 (N_4979,N_3539,N_3857);
or U4980 (N_4980,N_3528,N_3142);
or U4981 (N_4981,N_3661,N_3905);
or U4982 (N_4982,N_3768,N_3968);
or U4983 (N_4983,N_3170,N_3178);
nand U4984 (N_4984,N_3994,N_3196);
xnor U4985 (N_4985,N_3346,N_3996);
nor U4986 (N_4986,N_3496,N_3563);
and U4987 (N_4987,N_3849,N_3794);
nor U4988 (N_4988,N_3614,N_3156);
or U4989 (N_4989,N_3090,N_3475);
xor U4990 (N_4990,N_3767,N_3052);
nand U4991 (N_4991,N_3958,N_3664);
or U4992 (N_4992,N_3073,N_3309);
nor U4993 (N_4993,N_3210,N_3343);
nand U4994 (N_4994,N_3190,N_3881);
xor U4995 (N_4995,N_3957,N_3868);
nor U4996 (N_4996,N_3745,N_3761);
nor U4997 (N_4997,N_3879,N_3685);
nand U4998 (N_4998,N_3672,N_3820);
or U4999 (N_4999,N_3335,N_3723);
nand U5000 (N_5000,N_4535,N_4751);
or U5001 (N_5001,N_4542,N_4488);
or U5002 (N_5002,N_4564,N_4607);
nor U5003 (N_5003,N_4243,N_4261);
nor U5004 (N_5004,N_4846,N_4916);
nor U5005 (N_5005,N_4735,N_4606);
and U5006 (N_5006,N_4239,N_4913);
or U5007 (N_5007,N_4779,N_4965);
and U5008 (N_5008,N_4932,N_4926);
and U5009 (N_5009,N_4794,N_4126);
xnor U5010 (N_5010,N_4331,N_4734);
nand U5011 (N_5011,N_4221,N_4283);
nand U5012 (N_5012,N_4543,N_4176);
nor U5013 (N_5013,N_4130,N_4000);
or U5014 (N_5014,N_4536,N_4904);
nand U5015 (N_5015,N_4765,N_4228);
nor U5016 (N_5016,N_4417,N_4274);
and U5017 (N_5017,N_4848,N_4737);
or U5018 (N_5018,N_4882,N_4335);
and U5019 (N_5019,N_4077,N_4871);
or U5020 (N_5020,N_4634,N_4299);
or U5021 (N_5021,N_4079,N_4850);
xnor U5022 (N_5022,N_4797,N_4592);
and U5023 (N_5023,N_4340,N_4747);
and U5024 (N_5024,N_4520,N_4367);
or U5025 (N_5025,N_4081,N_4329);
nand U5026 (N_5026,N_4103,N_4609);
xor U5027 (N_5027,N_4514,N_4674);
nor U5028 (N_5028,N_4008,N_4654);
nand U5029 (N_5029,N_4512,N_4333);
or U5030 (N_5030,N_4143,N_4045);
xnor U5031 (N_5031,N_4697,N_4825);
and U5032 (N_5032,N_4772,N_4391);
nor U5033 (N_5033,N_4027,N_4432);
and U5034 (N_5034,N_4442,N_4475);
nor U5035 (N_5035,N_4059,N_4234);
or U5036 (N_5036,N_4866,N_4999);
nand U5037 (N_5037,N_4852,N_4682);
or U5038 (N_5038,N_4863,N_4807);
xor U5039 (N_5039,N_4286,N_4260);
or U5040 (N_5040,N_4516,N_4446);
and U5041 (N_5041,N_4470,N_4736);
or U5042 (N_5042,N_4328,N_4337);
and U5043 (N_5043,N_4139,N_4481);
xor U5044 (N_5044,N_4209,N_4468);
nor U5045 (N_5045,N_4531,N_4281);
xor U5046 (N_5046,N_4048,N_4411);
xor U5047 (N_5047,N_4409,N_4502);
xor U5048 (N_5048,N_4907,N_4146);
xnor U5049 (N_5049,N_4256,N_4742);
nor U5050 (N_5050,N_4269,N_4111);
nand U5051 (N_5051,N_4067,N_4085);
nand U5052 (N_5052,N_4738,N_4461);
and U5053 (N_5053,N_4345,N_4722);
nor U5054 (N_5054,N_4716,N_4853);
nor U5055 (N_5055,N_4847,N_4587);
and U5056 (N_5056,N_4421,N_4912);
nand U5057 (N_5057,N_4011,N_4202);
nand U5058 (N_5058,N_4496,N_4030);
or U5059 (N_5059,N_4350,N_4346);
xor U5060 (N_5060,N_4249,N_4230);
nor U5061 (N_5061,N_4185,N_4074);
and U5062 (N_5062,N_4289,N_4184);
xnor U5063 (N_5063,N_4359,N_4672);
nor U5064 (N_5064,N_4678,N_4268);
nor U5065 (N_5065,N_4135,N_4719);
xor U5066 (N_5066,N_4441,N_4616);
or U5067 (N_5067,N_4725,N_4201);
and U5068 (N_5068,N_4589,N_4972);
xor U5069 (N_5069,N_4998,N_4036);
or U5070 (N_5070,N_4472,N_4386);
or U5071 (N_5071,N_4830,N_4348);
nand U5072 (N_5072,N_4508,N_4180);
and U5073 (N_5073,N_4692,N_4608);
nand U5074 (N_5074,N_4696,N_4219);
or U5075 (N_5075,N_4207,N_4903);
or U5076 (N_5076,N_4068,N_4887);
nor U5077 (N_5077,N_4562,N_4877);
nand U5078 (N_5078,N_4941,N_4881);
nand U5079 (N_5079,N_4856,N_4790);
and U5080 (N_5080,N_4050,N_4947);
or U5081 (N_5081,N_4250,N_4691);
or U5082 (N_5082,N_4694,N_4651);
nor U5083 (N_5083,N_4977,N_4650);
and U5084 (N_5084,N_4600,N_4473);
and U5085 (N_5085,N_4844,N_4604);
and U5086 (N_5086,N_4583,N_4192);
xnor U5087 (N_5087,N_4458,N_4643);
or U5088 (N_5088,N_4010,N_4099);
or U5089 (N_5089,N_4954,N_4084);
xor U5090 (N_5090,N_4205,N_4767);
nand U5091 (N_5091,N_4360,N_4172);
nand U5092 (N_5092,N_4664,N_4246);
and U5093 (N_5093,N_4768,N_4232);
nor U5094 (N_5094,N_4310,N_4482);
xnor U5095 (N_5095,N_4715,N_4297);
xor U5096 (N_5096,N_4880,N_4558);
or U5097 (N_5097,N_4223,N_4469);
and U5098 (N_5098,N_4132,N_4906);
or U5099 (N_5099,N_4053,N_4471);
nor U5100 (N_5100,N_4686,N_4293);
and U5101 (N_5101,N_4819,N_4814);
and U5102 (N_5102,N_4875,N_4620);
or U5103 (N_5103,N_4817,N_4955);
and U5104 (N_5104,N_4104,N_4673);
or U5105 (N_5105,N_4801,N_4624);
nor U5106 (N_5106,N_4319,N_4981);
or U5107 (N_5107,N_4330,N_4802);
and U5108 (N_5108,N_4950,N_4304);
nor U5109 (N_5109,N_4298,N_4518);
or U5110 (N_5110,N_4775,N_4506);
or U5111 (N_5111,N_4901,N_4653);
or U5112 (N_5112,N_4623,N_4290);
nor U5113 (N_5113,N_4191,N_4021);
and U5114 (N_5114,N_4138,N_4829);
xnor U5115 (N_5115,N_4167,N_4037);
nand U5116 (N_5116,N_4440,N_4748);
nand U5117 (N_5117,N_4773,N_4425);
and U5118 (N_5118,N_4480,N_4364);
xor U5119 (N_5119,N_4733,N_4428);
nor U5120 (N_5120,N_4646,N_4905);
or U5121 (N_5121,N_4115,N_4979);
nor U5122 (N_5122,N_4820,N_4296);
or U5123 (N_5123,N_4140,N_4336);
and U5124 (N_5124,N_4540,N_4983);
and U5125 (N_5125,N_4133,N_4776);
and U5126 (N_5126,N_4054,N_4888);
xnor U5127 (N_5127,N_4534,N_4577);
nor U5128 (N_5128,N_4484,N_4042);
and U5129 (N_5129,N_4033,N_4170);
xor U5130 (N_5130,N_4769,N_4395);
nor U5131 (N_5131,N_4575,N_4665);
xnor U5132 (N_5132,N_4056,N_4365);
nor U5133 (N_5133,N_4247,N_4810);
and U5134 (N_5134,N_4464,N_4612);
or U5135 (N_5135,N_4016,N_4766);
and U5136 (N_5136,N_4402,N_4164);
nor U5137 (N_5137,N_4334,N_4619);
nor U5138 (N_5138,N_4181,N_4519);
and U5139 (N_5139,N_4574,N_4559);
or U5140 (N_5140,N_4515,N_4277);
xnor U5141 (N_5141,N_4525,N_4640);
nor U5142 (N_5142,N_4029,N_4570);
nand U5143 (N_5143,N_4291,N_4509);
xnor U5144 (N_5144,N_4366,N_4422);
xor U5145 (N_5145,N_4278,N_4960);
xnor U5146 (N_5146,N_4724,N_4946);
nor U5147 (N_5147,N_4430,N_4627);
and U5148 (N_5148,N_4971,N_4656);
or U5149 (N_5149,N_4248,N_4460);
nor U5150 (N_5150,N_4320,N_4655);
xor U5151 (N_5151,N_4677,N_4339);
or U5152 (N_5152,N_4154,N_4936);
xor U5153 (N_5153,N_4821,N_4097);
nor U5154 (N_5154,N_4980,N_4265);
xnor U5155 (N_5155,N_4282,N_4770);
xnor U5156 (N_5156,N_4159,N_4136);
nand U5157 (N_5157,N_4034,N_4567);
xor U5158 (N_5158,N_4240,N_4521);
nor U5159 (N_5159,N_4098,N_4833);
xnor U5160 (N_5160,N_4996,N_4874);
or U5161 (N_5161,N_4726,N_4303);
and U5162 (N_5162,N_4668,N_4857);
nor U5163 (N_5163,N_4206,N_4476);
nand U5164 (N_5164,N_4595,N_4550);
or U5165 (N_5165,N_4593,N_4803);
or U5166 (N_5166,N_4675,N_4970);
nor U5167 (N_5167,N_4670,N_4704);
or U5168 (N_5168,N_4295,N_4617);
and U5169 (N_5169,N_4865,N_4727);
and U5170 (N_5170,N_4992,N_4944);
xor U5171 (N_5171,N_4233,N_4114);
nor U5172 (N_5172,N_4071,N_4973);
nor U5173 (N_5173,N_4862,N_4208);
nor U5174 (N_5174,N_4312,N_4193);
nand U5175 (N_5175,N_4003,N_4683);
xnor U5176 (N_5176,N_4487,N_4622);
or U5177 (N_5177,N_4764,N_4405);
xor U5178 (N_5178,N_4465,N_4910);
and U5179 (N_5179,N_4072,N_4958);
or U5180 (N_5180,N_4721,N_4571);
or U5181 (N_5181,N_4444,N_4047);
or U5182 (N_5182,N_4493,N_4568);
nand U5183 (N_5183,N_4501,N_4255);
nand U5184 (N_5184,N_4579,N_4511);
nor U5185 (N_5185,N_4919,N_4591);
xor U5186 (N_5186,N_4147,N_4080);
and U5187 (N_5187,N_4148,N_4435);
nor U5188 (N_5188,N_4922,N_4459);
and U5189 (N_5189,N_4566,N_4178);
nor U5190 (N_5190,N_4368,N_4541);
or U5191 (N_5191,N_4161,N_4210);
nand U5192 (N_5192,N_4194,N_4707);
nor U5193 (N_5193,N_4762,N_4043);
and U5194 (N_5194,N_4049,N_4845);
nor U5195 (N_5195,N_4284,N_4752);
xor U5196 (N_5196,N_4614,N_4083);
or U5197 (N_5197,N_4279,N_4717);
xor U5198 (N_5198,N_4401,N_4545);
and U5199 (N_5199,N_4106,N_4078);
and U5200 (N_5200,N_4065,N_4602);
and U5201 (N_5201,N_4244,N_4382);
and U5202 (N_5202,N_4700,N_4022);
nand U5203 (N_5203,N_4522,N_4920);
and U5204 (N_5204,N_4051,N_4058);
xor U5205 (N_5205,N_4870,N_4573);
xor U5206 (N_5206,N_4006,N_4175);
xnor U5207 (N_5207,N_4952,N_4578);
nand U5208 (N_5208,N_4393,N_4179);
nand U5209 (N_5209,N_4356,N_4272);
nor U5210 (N_5210,N_4069,N_4964);
nand U5211 (N_5211,N_4548,N_4093);
or U5212 (N_5212,N_4528,N_4236);
nor U5213 (N_5213,N_4537,N_4057);
and U5214 (N_5214,N_4757,N_4419);
or U5215 (N_5215,N_4145,N_4500);
nor U5216 (N_5216,N_4834,N_4288);
and U5217 (N_5217,N_4266,N_4226);
and U5218 (N_5218,N_4855,N_4137);
nor U5219 (N_5219,N_4533,N_4112);
nand U5220 (N_5220,N_4394,N_4584);
nand U5221 (N_5221,N_4371,N_4925);
nor U5222 (N_5222,N_4885,N_4787);
nand U5223 (N_5223,N_4427,N_4276);
nand U5224 (N_5224,N_4990,N_4526);
or U5225 (N_5225,N_4594,N_4743);
nor U5226 (N_5226,N_4759,N_4532);
xnor U5227 (N_5227,N_4215,N_4557);
and U5228 (N_5228,N_4235,N_4756);
or U5229 (N_5229,N_4495,N_4693);
or U5230 (N_5230,N_4914,N_4959);
and U5231 (N_5231,N_4598,N_4760);
or U5232 (N_5232,N_4529,N_4315);
or U5233 (N_5233,N_4553,N_4341);
nor U5234 (N_5234,N_4991,N_4659);
nand U5235 (N_5235,N_4387,N_4546);
nand U5236 (N_5236,N_4997,N_4032);
nor U5237 (N_5237,N_4153,N_4257);
xor U5238 (N_5238,N_4811,N_4373);
or U5239 (N_5239,N_4060,N_4252);
xnor U5240 (N_5240,N_4306,N_4188);
nor U5241 (N_5241,N_4549,N_4687);
xor U5242 (N_5242,N_4122,N_4489);
xnor U5243 (N_5243,N_4129,N_4052);
and U5244 (N_5244,N_4062,N_4791);
nand U5245 (N_5245,N_4452,N_4507);
and U5246 (N_5246,N_4151,N_4101);
and U5247 (N_5247,N_4889,N_4438);
and U5248 (N_5248,N_4615,N_4307);
xor U5249 (N_5249,N_4158,N_4504);
nor U5250 (N_5250,N_4636,N_4186);
and U5251 (N_5251,N_4777,N_4793);
and U5252 (N_5252,N_4923,N_4200);
xor U5253 (N_5253,N_4357,N_4224);
xor U5254 (N_5254,N_4799,N_4771);
nor U5255 (N_5255,N_4780,N_4864);
xor U5256 (N_5256,N_4899,N_4688);
and U5257 (N_5257,N_4044,N_4878);
and U5258 (N_5258,N_4826,N_4018);
nand U5259 (N_5259,N_4741,N_4258);
xor U5260 (N_5260,N_4629,N_4551);
nor U5261 (N_5261,N_4942,N_4978);
or U5262 (N_5262,N_4218,N_4915);
nor U5263 (N_5263,N_4822,N_4642);
nand U5264 (N_5264,N_4007,N_4993);
xor U5265 (N_5265,N_4462,N_4301);
xnor U5266 (N_5266,N_4217,N_4416);
nand U5267 (N_5267,N_4969,N_4927);
xor U5268 (N_5268,N_4563,N_4177);
and U5269 (N_5269,N_4711,N_4892);
nor U5270 (N_5270,N_4004,N_4648);
and U5271 (N_5271,N_4374,N_4828);
and U5272 (N_5272,N_4841,N_4705);
or U5273 (N_5273,N_4009,N_4220);
xnor U5274 (N_5274,N_4424,N_4182);
or U5275 (N_5275,N_4505,N_4613);
and U5276 (N_5276,N_4975,N_4835);
and U5277 (N_5277,N_4372,N_4581);
and U5278 (N_5278,N_4203,N_4994);
or U5279 (N_5279,N_4431,N_4398);
nor U5280 (N_5280,N_4381,N_4089);
nor U5281 (N_5281,N_4131,N_4038);
nor U5282 (N_5282,N_4527,N_4679);
and U5283 (N_5283,N_4831,N_4443);
nand U5284 (N_5284,N_4861,N_4890);
and U5285 (N_5285,N_4753,N_4453);
xor U5286 (N_5286,N_4805,N_4897);
and U5287 (N_5287,N_4872,N_4127);
nor U5288 (N_5288,N_4869,N_4690);
xor U5289 (N_5289,N_4397,N_4031);
xor U5290 (N_5290,N_4843,N_4091);
nor U5291 (N_5291,N_4204,N_4001);
nand U5292 (N_5292,N_4588,N_4412);
and U5293 (N_5293,N_4778,N_4370);
xor U5294 (N_5294,N_4755,N_4580);
nand U5295 (N_5295,N_4349,N_4597);
and U5296 (N_5296,N_4389,N_4924);
and U5297 (N_5297,N_4763,N_4241);
xnor U5298 (N_5298,N_4966,N_4723);
nand U5299 (N_5299,N_4168,N_4681);
or U5300 (N_5300,N_4292,N_4585);
and U5301 (N_5301,N_4860,N_4023);
xnor U5302 (N_5302,N_4781,N_4456);
xor U5303 (N_5303,N_4657,N_4949);
nor U5304 (N_5304,N_4216,N_4940);
xnor U5305 (N_5305,N_4020,N_4699);
nand U5306 (N_5306,N_4676,N_4183);
nand U5307 (N_5307,N_4404,N_4451);
nor U5308 (N_5308,N_4390,N_4714);
nand U5309 (N_5309,N_4231,N_4254);
xnor U5310 (N_5310,N_4426,N_4784);
nand U5311 (N_5311,N_4943,N_4963);
nand U5312 (N_5312,N_4423,N_4709);
nand U5313 (N_5313,N_4611,N_4322);
and U5314 (N_5314,N_4355,N_4728);
and U5315 (N_5315,N_4840,N_4197);
and U5316 (N_5316,N_4795,N_4087);
and U5317 (N_5317,N_4406,N_4832);
xor U5318 (N_5318,N_4895,N_4450);
and U5319 (N_5319,N_4929,N_4663);
and U5320 (N_5320,N_4174,N_4893);
or U5321 (N_5321,N_4447,N_4317);
nand U5322 (N_5322,N_4478,N_4930);
nor U5323 (N_5323,N_4666,N_4107);
nor U5324 (N_5324,N_4433,N_4075);
nand U5325 (N_5325,N_4908,N_4859);
and U5326 (N_5326,N_4227,N_4720);
and U5327 (N_5327,N_4938,N_4544);
or U5328 (N_5328,N_4073,N_4812);
xnor U5329 (N_5329,N_4539,N_4156);
nand U5330 (N_5330,N_4886,N_4891);
nand U5331 (N_5331,N_4917,N_4785);
or U5332 (N_5332,N_4400,N_4806);
xor U5333 (N_5333,N_4403,N_4851);
and U5334 (N_5334,N_4094,N_4524);
xnor U5335 (N_5335,N_4141,N_4530);
and U5336 (N_5336,N_4420,N_4647);
xor U5337 (N_5337,N_4909,N_4379);
nand U5338 (N_5338,N_4739,N_4900);
and U5339 (N_5339,N_4576,N_4935);
nand U5340 (N_5340,N_4198,N_4449);
nand U5341 (N_5341,N_4457,N_4351);
or U5342 (N_5342,N_4552,N_4933);
xnor U5343 (N_5343,N_4731,N_4652);
and U5344 (N_5344,N_4110,N_4454);
nand U5345 (N_5345,N_4347,N_4160);
nor U5346 (N_5346,N_4002,N_4984);
and U5347 (N_5347,N_4750,N_4327);
nor U5348 (N_5348,N_4212,N_4109);
xor U5349 (N_5349,N_4013,N_4867);
nand U5350 (N_5350,N_4123,N_4499);
nand U5351 (N_5351,N_4961,N_4565);
nand U5352 (N_5352,N_4633,N_4934);
nor U5353 (N_5353,N_4300,N_4637);
and U5354 (N_5354,N_4388,N_4586);
nor U5355 (N_5355,N_4928,N_4582);
xor U5356 (N_5356,N_4354,N_4105);
or U5357 (N_5357,N_4754,N_4658);
nand U5358 (N_5358,N_4618,N_4786);
xnor U5359 (N_5359,N_4155,N_4572);
nor U5360 (N_5360,N_4884,N_4989);
and U5361 (N_5361,N_4976,N_4641);
xor U5362 (N_5362,N_4792,N_4931);
or U5363 (N_5363,N_4245,N_4490);
xor U5364 (N_5364,N_4066,N_4015);
nor U5365 (N_5365,N_4196,N_4662);
nor U5366 (N_5366,N_4560,N_4090);
xor U5367 (N_5367,N_4119,N_4649);
and U5368 (N_5368,N_4157,N_4621);
and U5369 (N_5369,N_4171,N_4092);
and U5370 (N_5370,N_4342,N_4815);
nor U5371 (N_5371,N_4352,N_4494);
xor U5372 (N_5372,N_4684,N_4804);
nor U5373 (N_5373,N_4408,N_4967);
xnor U5374 (N_5374,N_4410,N_4418);
xnor U5375 (N_5375,N_4173,N_4635);
nand U5376 (N_5376,N_4353,N_4024);
nand U5377 (N_5377,N_4474,N_4986);
and U5378 (N_5378,N_4150,N_4894);
and U5379 (N_5379,N_4399,N_4323);
and U5380 (N_5380,N_4873,N_4842);
xor U5381 (N_5381,N_4921,N_4225);
nand U5382 (N_5382,N_4556,N_4729);
or U5383 (N_5383,N_4957,N_4713);
or U5384 (N_5384,N_4685,N_4344);
and U5385 (N_5385,N_4237,N_4788);
or U5386 (N_5386,N_4603,N_4088);
or U5387 (N_5387,N_4626,N_4325);
xnor U5388 (N_5388,N_4055,N_4166);
or U5389 (N_5389,N_4267,N_4937);
nand U5390 (N_5390,N_4982,N_4086);
nor U5391 (N_5391,N_4280,N_4305);
xnor U5392 (N_5392,N_4632,N_4375);
xnor U5393 (N_5393,N_4695,N_4968);
or U5394 (N_5394,N_4117,N_4761);
nor U5395 (N_5395,N_4270,N_4898);
nand U5396 (N_5396,N_4745,N_4229);
and U5397 (N_5397,N_4988,N_4439);
or U5398 (N_5398,N_4638,N_4321);
xor U5399 (N_5399,N_4590,N_4477);
nor U5400 (N_5400,N_4383,N_4839);
nor U5401 (N_5401,N_4945,N_4076);
xor U5402 (N_5402,N_4096,N_4195);
or U5403 (N_5403,N_4547,N_4144);
nor U5404 (N_5404,N_4703,N_4601);
and U5405 (N_5405,N_4378,N_4498);
xor U5406 (N_5406,N_4214,N_4596);
xor U5407 (N_5407,N_4689,N_4466);
nand U5408 (N_5408,N_4165,N_4318);
xnor U5409 (N_5409,N_4818,N_4035);
xnor U5410 (N_5410,N_4854,N_4262);
and U5411 (N_5411,N_4486,N_4702);
or U5412 (N_5412,N_4012,N_4883);
and U5413 (N_5413,N_4120,N_4377);
or U5414 (N_5414,N_4149,N_4463);
and U5415 (N_5415,N_4385,N_4605);
nand U5416 (N_5416,N_4287,N_4163);
nor U5417 (N_5417,N_4523,N_4902);
xor U5418 (N_5418,N_4273,N_4680);
nand U5419 (N_5419,N_4796,N_4956);
nand U5420 (N_5420,N_4698,N_4706);
or U5421 (N_5421,N_4479,N_4407);
xor U5422 (N_5422,N_4100,N_4644);
and U5423 (N_5423,N_4251,N_4491);
or U5424 (N_5424,N_4599,N_4974);
xor U5425 (N_5425,N_4314,N_4701);
or U5426 (N_5426,N_4669,N_4836);
and U5427 (N_5427,N_4610,N_4730);
nor U5428 (N_5428,N_4660,N_4774);
or U5429 (N_5429,N_4798,N_4896);
or U5430 (N_5430,N_4948,N_4800);
nand U5431 (N_5431,N_4628,N_4124);
or U5432 (N_5432,N_4162,N_4911);
and U5433 (N_5433,N_4121,N_4671);
nand U5434 (N_5434,N_4561,N_4190);
nand U5435 (N_5435,N_4253,N_4485);
nand U5436 (N_5436,N_4275,N_4823);
and U5437 (N_5437,N_4362,N_4413);
nor U5438 (N_5438,N_4187,N_4436);
and U5439 (N_5439,N_4061,N_4063);
nand U5440 (N_5440,N_4858,N_4712);
xnor U5441 (N_5441,N_4782,N_4434);
and U5442 (N_5442,N_4285,N_4169);
xnor U5443 (N_5443,N_4046,N_4108);
nor U5444 (N_5444,N_4376,N_4510);
or U5445 (N_5445,N_4455,N_4808);
nand U5446 (N_5446,N_4758,N_4789);
nor U5447 (N_5447,N_4316,N_4639);
or U5448 (N_5448,N_4102,N_4538);
nor U5449 (N_5449,N_4744,N_4326);
xor U5450 (N_5450,N_4467,N_4437);
and U5451 (N_5451,N_4302,N_4879);
and U5452 (N_5452,N_4838,N_4311);
and U5453 (N_5453,N_4040,N_4294);
xor U5454 (N_5454,N_4503,N_4661);
xnor U5455 (N_5455,N_4019,N_4953);
xor U5456 (N_5456,N_4497,N_4630);
or U5457 (N_5457,N_4363,N_4918);
nor U5458 (N_5458,N_4645,N_4308);
nand U5459 (N_5459,N_4824,N_4026);
or U5460 (N_5460,N_4849,N_4492);
or U5461 (N_5461,N_4569,N_4445);
or U5462 (N_5462,N_4962,N_4142);
nand U5463 (N_5463,N_4396,N_4039);
and U5464 (N_5464,N_4116,N_4813);
or U5465 (N_5465,N_4783,N_4816);
nand U5466 (N_5466,N_4554,N_4025);
nand U5467 (N_5467,N_4082,N_4513);
xnor U5468 (N_5468,N_4732,N_4837);
nor U5469 (N_5469,N_4199,N_4749);
nor U5470 (N_5470,N_4343,N_4118);
and U5471 (N_5471,N_4271,N_4392);
xor U5472 (N_5472,N_4876,N_4222);
nor U5473 (N_5473,N_4987,N_4995);
and U5474 (N_5474,N_4555,N_4369);
nor U5475 (N_5475,N_4710,N_4361);
and U5476 (N_5476,N_4189,N_4309);
and U5477 (N_5477,N_4868,N_4358);
or U5478 (N_5478,N_4985,N_4827);
xor U5479 (N_5479,N_4028,N_4667);
or U5480 (N_5480,N_4740,N_4631);
and U5481 (N_5481,N_4242,N_4070);
nand U5482 (N_5482,N_4125,N_4414);
and U5483 (N_5483,N_4809,N_4005);
nor U5484 (N_5484,N_4064,N_4017);
nor U5485 (N_5485,N_4211,N_4380);
xnor U5486 (N_5486,N_4014,N_4746);
or U5487 (N_5487,N_4625,N_4429);
and U5488 (N_5488,N_4384,N_4718);
and U5489 (N_5489,N_4095,N_4238);
xnor U5490 (N_5490,N_4448,N_4939);
nor U5491 (N_5491,N_4338,N_4324);
nor U5492 (N_5492,N_4152,N_4313);
or U5493 (N_5493,N_4517,N_4708);
or U5494 (N_5494,N_4259,N_4263);
and U5495 (N_5495,N_4415,N_4041);
and U5496 (N_5496,N_4483,N_4128);
nand U5497 (N_5497,N_4951,N_4264);
xor U5498 (N_5498,N_4134,N_4332);
xnor U5499 (N_5499,N_4213,N_4113);
and U5500 (N_5500,N_4286,N_4017);
and U5501 (N_5501,N_4161,N_4169);
nor U5502 (N_5502,N_4436,N_4517);
nor U5503 (N_5503,N_4612,N_4423);
xor U5504 (N_5504,N_4739,N_4244);
nor U5505 (N_5505,N_4244,N_4301);
and U5506 (N_5506,N_4888,N_4571);
nor U5507 (N_5507,N_4350,N_4116);
xor U5508 (N_5508,N_4289,N_4072);
xor U5509 (N_5509,N_4411,N_4276);
xnor U5510 (N_5510,N_4029,N_4973);
or U5511 (N_5511,N_4477,N_4351);
nor U5512 (N_5512,N_4443,N_4224);
nand U5513 (N_5513,N_4988,N_4348);
nand U5514 (N_5514,N_4521,N_4686);
nand U5515 (N_5515,N_4275,N_4369);
and U5516 (N_5516,N_4451,N_4532);
or U5517 (N_5517,N_4072,N_4319);
nor U5518 (N_5518,N_4556,N_4757);
nor U5519 (N_5519,N_4344,N_4023);
and U5520 (N_5520,N_4640,N_4781);
nor U5521 (N_5521,N_4654,N_4281);
nor U5522 (N_5522,N_4218,N_4592);
xnor U5523 (N_5523,N_4549,N_4622);
nand U5524 (N_5524,N_4645,N_4525);
nor U5525 (N_5525,N_4036,N_4068);
and U5526 (N_5526,N_4573,N_4213);
nand U5527 (N_5527,N_4500,N_4320);
and U5528 (N_5528,N_4246,N_4408);
nor U5529 (N_5529,N_4069,N_4652);
and U5530 (N_5530,N_4836,N_4120);
nor U5531 (N_5531,N_4260,N_4107);
nor U5532 (N_5532,N_4637,N_4812);
xnor U5533 (N_5533,N_4958,N_4314);
xor U5534 (N_5534,N_4283,N_4257);
xnor U5535 (N_5535,N_4368,N_4339);
and U5536 (N_5536,N_4345,N_4625);
xor U5537 (N_5537,N_4723,N_4615);
and U5538 (N_5538,N_4814,N_4585);
nand U5539 (N_5539,N_4671,N_4710);
nor U5540 (N_5540,N_4354,N_4189);
and U5541 (N_5541,N_4603,N_4680);
nor U5542 (N_5542,N_4474,N_4919);
and U5543 (N_5543,N_4755,N_4878);
or U5544 (N_5544,N_4535,N_4776);
nand U5545 (N_5545,N_4623,N_4925);
nand U5546 (N_5546,N_4350,N_4974);
and U5547 (N_5547,N_4089,N_4810);
xor U5548 (N_5548,N_4537,N_4885);
xor U5549 (N_5549,N_4601,N_4003);
xnor U5550 (N_5550,N_4376,N_4293);
xor U5551 (N_5551,N_4280,N_4895);
nand U5552 (N_5552,N_4978,N_4627);
or U5553 (N_5553,N_4932,N_4392);
or U5554 (N_5554,N_4040,N_4714);
nand U5555 (N_5555,N_4949,N_4281);
nor U5556 (N_5556,N_4333,N_4732);
nor U5557 (N_5557,N_4899,N_4810);
nor U5558 (N_5558,N_4174,N_4026);
xnor U5559 (N_5559,N_4606,N_4697);
xor U5560 (N_5560,N_4629,N_4660);
or U5561 (N_5561,N_4739,N_4895);
and U5562 (N_5562,N_4746,N_4691);
nand U5563 (N_5563,N_4108,N_4154);
nor U5564 (N_5564,N_4934,N_4829);
nor U5565 (N_5565,N_4989,N_4323);
nor U5566 (N_5566,N_4899,N_4235);
nand U5567 (N_5567,N_4104,N_4484);
or U5568 (N_5568,N_4896,N_4390);
or U5569 (N_5569,N_4603,N_4506);
and U5570 (N_5570,N_4526,N_4600);
or U5571 (N_5571,N_4318,N_4350);
nor U5572 (N_5572,N_4648,N_4300);
or U5573 (N_5573,N_4409,N_4495);
xor U5574 (N_5574,N_4183,N_4466);
nor U5575 (N_5575,N_4833,N_4630);
and U5576 (N_5576,N_4212,N_4090);
nor U5577 (N_5577,N_4562,N_4069);
and U5578 (N_5578,N_4546,N_4139);
xnor U5579 (N_5579,N_4751,N_4571);
nand U5580 (N_5580,N_4097,N_4852);
xor U5581 (N_5581,N_4791,N_4603);
or U5582 (N_5582,N_4454,N_4403);
or U5583 (N_5583,N_4850,N_4377);
and U5584 (N_5584,N_4015,N_4770);
and U5585 (N_5585,N_4717,N_4657);
nand U5586 (N_5586,N_4098,N_4365);
and U5587 (N_5587,N_4781,N_4311);
nand U5588 (N_5588,N_4554,N_4018);
or U5589 (N_5589,N_4787,N_4435);
nand U5590 (N_5590,N_4680,N_4894);
xnor U5591 (N_5591,N_4862,N_4358);
xor U5592 (N_5592,N_4183,N_4289);
and U5593 (N_5593,N_4445,N_4329);
xor U5594 (N_5594,N_4701,N_4141);
xnor U5595 (N_5595,N_4569,N_4423);
xnor U5596 (N_5596,N_4281,N_4630);
nor U5597 (N_5597,N_4815,N_4724);
nand U5598 (N_5598,N_4632,N_4266);
nand U5599 (N_5599,N_4660,N_4225);
nor U5600 (N_5600,N_4779,N_4427);
nand U5601 (N_5601,N_4054,N_4256);
xor U5602 (N_5602,N_4800,N_4040);
nor U5603 (N_5603,N_4025,N_4849);
nor U5604 (N_5604,N_4191,N_4265);
or U5605 (N_5605,N_4666,N_4888);
and U5606 (N_5606,N_4424,N_4351);
nor U5607 (N_5607,N_4274,N_4243);
nand U5608 (N_5608,N_4944,N_4677);
and U5609 (N_5609,N_4164,N_4242);
or U5610 (N_5610,N_4154,N_4582);
nand U5611 (N_5611,N_4368,N_4909);
nand U5612 (N_5612,N_4004,N_4145);
nor U5613 (N_5613,N_4199,N_4070);
or U5614 (N_5614,N_4296,N_4670);
or U5615 (N_5615,N_4288,N_4344);
nand U5616 (N_5616,N_4600,N_4223);
and U5617 (N_5617,N_4878,N_4632);
nor U5618 (N_5618,N_4910,N_4277);
nor U5619 (N_5619,N_4164,N_4029);
nor U5620 (N_5620,N_4428,N_4357);
and U5621 (N_5621,N_4188,N_4812);
xor U5622 (N_5622,N_4519,N_4980);
nor U5623 (N_5623,N_4691,N_4391);
nor U5624 (N_5624,N_4944,N_4805);
and U5625 (N_5625,N_4552,N_4563);
nor U5626 (N_5626,N_4775,N_4534);
or U5627 (N_5627,N_4481,N_4102);
and U5628 (N_5628,N_4046,N_4775);
and U5629 (N_5629,N_4563,N_4446);
nand U5630 (N_5630,N_4450,N_4062);
and U5631 (N_5631,N_4855,N_4994);
or U5632 (N_5632,N_4445,N_4273);
and U5633 (N_5633,N_4684,N_4195);
xor U5634 (N_5634,N_4376,N_4970);
xnor U5635 (N_5635,N_4136,N_4887);
xor U5636 (N_5636,N_4660,N_4282);
nand U5637 (N_5637,N_4193,N_4156);
xor U5638 (N_5638,N_4042,N_4799);
nand U5639 (N_5639,N_4234,N_4042);
and U5640 (N_5640,N_4271,N_4960);
xor U5641 (N_5641,N_4300,N_4659);
and U5642 (N_5642,N_4127,N_4422);
nor U5643 (N_5643,N_4573,N_4422);
and U5644 (N_5644,N_4538,N_4237);
nor U5645 (N_5645,N_4606,N_4287);
xor U5646 (N_5646,N_4893,N_4622);
nand U5647 (N_5647,N_4756,N_4218);
nor U5648 (N_5648,N_4149,N_4627);
or U5649 (N_5649,N_4296,N_4504);
or U5650 (N_5650,N_4977,N_4012);
nor U5651 (N_5651,N_4015,N_4272);
or U5652 (N_5652,N_4703,N_4889);
or U5653 (N_5653,N_4642,N_4930);
nor U5654 (N_5654,N_4503,N_4624);
nor U5655 (N_5655,N_4314,N_4876);
and U5656 (N_5656,N_4532,N_4494);
xor U5657 (N_5657,N_4342,N_4978);
and U5658 (N_5658,N_4639,N_4066);
nor U5659 (N_5659,N_4754,N_4927);
nor U5660 (N_5660,N_4740,N_4414);
xnor U5661 (N_5661,N_4661,N_4858);
nand U5662 (N_5662,N_4236,N_4419);
and U5663 (N_5663,N_4939,N_4485);
nand U5664 (N_5664,N_4833,N_4414);
nand U5665 (N_5665,N_4205,N_4958);
or U5666 (N_5666,N_4238,N_4345);
or U5667 (N_5667,N_4496,N_4379);
xnor U5668 (N_5668,N_4669,N_4696);
nor U5669 (N_5669,N_4484,N_4253);
and U5670 (N_5670,N_4703,N_4411);
nor U5671 (N_5671,N_4942,N_4495);
or U5672 (N_5672,N_4674,N_4084);
and U5673 (N_5673,N_4578,N_4976);
or U5674 (N_5674,N_4294,N_4796);
and U5675 (N_5675,N_4458,N_4123);
nor U5676 (N_5676,N_4476,N_4918);
nor U5677 (N_5677,N_4791,N_4476);
and U5678 (N_5678,N_4991,N_4748);
nand U5679 (N_5679,N_4662,N_4414);
nand U5680 (N_5680,N_4030,N_4882);
nand U5681 (N_5681,N_4503,N_4030);
xnor U5682 (N_5682,N_4360,N_4578);
and U5683 (N_5683,N_4891,N_4733);
or U5684 (N_5684,N_4741,N_4181);
xnor U5685 (N_5685,N_4095,N_4865);
xor U5686 (N_5686,N_4002,N_4262);
and U5687 (N_5687,N_4644,N_4829);
or U5688 (N_5688,N_4480,N_4769);
xnor U5689 (N_5689,N_4585,N_4829);
nand U5690 (N_5690,N_4312,N_4936);
or U5691 (N_5691,N_4084,N_4419);
or U5692 (N_5692,N_4532,N_4655);
and U5693 (N_5693,N_4116,N_4854);
and U5694 (N_5694,N_4627,N_4721);
xor U5695 (N_5695,N_4108,N_4304);
nand U5696 (N_5696,N_4072,N_4472);
nor U5697 (N_5697,N_4792,N_4417);
and U5698 (N_5698,N_4580,N_4874);
xor U5699 (N_5699,N_4200,N_4189);
nand U5700 (N_5700,N_4952,N_4373);
nor U5701 (N_5701,N_4017,N_4473);
nor U5702 (N_5702,N_4240,N_4269);
or U5703 (N_5703,N_4073,N_4582);
nor U5704 (N_5704,N_4280,N_4311);
and U5705 (N_5705,N_4801,N_4130);
or U5706 (N_5706,N_4677,N_4513);
nand U5707 (N_5707,N_4238,N_4101);
nand U5708 (N_5708,N_4581,N_4992);
nand U5709 (N_5709,N_4094,N_4885);
and U5710 (N_5710,N_4179,N_4356);
nor U5711 (N_5711,N_4784,N_4119);
nor U5712 (N_5712,N_4531,N_4204);
xor U5713 (N_5713,N_4913,N_4055);
nor U5714 (N_5714,N_4404,N_4663);
or U5715 (N_5715,N_4855,N_4449);
and U5716 (N_5716,N_4098,N_4514);
nand U5717 (N_5717,N_4599,N_4063);
nand U5718 (N_5718,N_4495,N_4207);
nand U5719 (N_5719,N_4856,N_4480);
nand U5720 (N_5720,N_4060,N_4157);
and U5721 (N_5721,N_4904,N_4923);
nor U5722 (N_5722,N_4236,N_4199);
or U5723 (N_5723,N_4514,N_4390);
and U5724 (N_5724,N_4658,N_4389);
nor U5725 (N_5725,N_4287,N_4054);
xor U5726 (N_5726,N_4027,N_4158);
nor U5727 (N_5727,N_4187,N_4556);
or U5728 (N_5728,N_4944,N_4858);
xor U5729 (N_5729,N_4636,N_4827);
and U5730 (N_5730,N_4056,N_4153);
and U5731 (N_5731,N_4861,N_4903);
nand U5732 (N_5732,N_4876,N_4691);
xor U5733 (N_5733,N_4972,N_4875);
or U5734 (N_5734,N_4773,N_4898);
nand U5735 (N_5735,N_4534,N_4222);
and U5736 (N_5736,N_4348,N_4369);
or U5737 (N_5737,N_4175,N_4500);
nor U5738 (N_5738,N_4082,N_4894);
nor U5739 (N_5739,N_4230,N_4329);
nor U5740 (N_5740,N_4611,N_4745);
nor U5741 (N_5741,N_4687,N_4395);
nand U5742 (N_5742,N_4090,N_4226);
or U5743 (N_5743,N_4219,N_4103);
nor U5744 (N_5744,N_4341,N_4775);
and U5745 (N_5745,N_4629,N_4769);
nor U5746 (N_5746,N_4321,N_4352);
nand U5747 (N_5747,N_4283,N_4439);
nor U5748 (N_5748,N_4259,N_4325);
nor U5749 (N_5749,N_4314,N_4290);
xor U5750 (N_5750,N_4789,N_4857);
nor U5751 (N_5751,N_4786,N_4309);
nor U5752 (N_5752,N_4193,N_4674);
xnor U5753 (N_5753,N_4008,N_4699);
nand U5754 (N_5754,N_4342,N_4879);
and U5755 (N_5755,N_4251,N_4137);
nand U5756 (N_5756,N_4787,N_4463);
nor U5757 (N_5757,N_4746,N_4074);
and U5758 (N_5758,N_4965,N_4434);
xnor U5759 (N_5759,N_4052,N_4013);
or U5760 (N_5760,N_4980,N_4450);
nand U5761 (N_5761,N_4030,N_4491);
xnor U5762 (N_5762,N_4400,N_4273);
nor U5763 (N_5763,N_4821,N_4290);
nand U5764 (N_5764,N_4098,N_4316);
xnor U5765 (N_5765,N_4190,N_4500);
or U5766 (N_5766,N_4530,N_4889);
nand U5767 (N_5767,N_4777,N_4359);
and U5768 (N_5768,N_4246,N_4056);
and U5769 (N_5769,N_4886,N_4808);
nor U5770 (N_5770,N_4998,N_4416);
nor U5771 (N_5771,N_4107,N_4772);
xnor U5772 (N_5772,N_4593,N_4806);
or U5773 (N_5773,N_4470,N_4154);
or U5774 (N_5774,N_4387,N_4884);
and U5775 (N_5775,N_4412,N_4859);
nand U5776 (N_5776,N_4567,N_4662);
or U5777 (N_5777,N_4464,N_4459);
nand U5778 (N_5778,N_4829,N_4667);
xnor U5779 (N_5779,N_4950,N_4370);
xor U5780 (N_5780,N_4943,N_4262);
nand U5781 (N_5781,N_4229,N_4384);
or U5782 (N_5782,N_4044,N_4982);
and U5783 (N_5783,N_4870,N_4557);
or U5784 (N_5784,N_4277,N_4089);
xor U5785 (N_5785,N_4854,N_4119);
nand U5786 (N_5786,N_4617,N_4816);
xor U5787 (N_5787,N_4269,N_4715);
xnor U5788 (N_5788,N_4289,N_4712);
nor U5789 (N_5789,N_4186,N_4586);
or U5790 (N_5790,N_4668,N_4388);
or U5791 (N_5791,N_4911,N_4353);
or U5792 (N_5792,N_4794,N_4951);
xnor U5793 (N_5793,N_4098,N_4484);
nand U5794 (N_5794,N_4007,N_4440);
and U5795 (N_5795,N_4470,N_4255);
and U5796 (N_5796,N_4343,N_4769);
or U5797 (N_5797,N_4518,N_4772);
or U5798 (N_5798,N_4215,N_4432);
nor U5799 (N_5799,N_4735,N_4813);
xor U5800 (N_5800,N_4852,N_4283);
xnor U5801 (N_5801,N_4259,N_4297);
nor U5802 (N_5802,N_4248,N_4883);
or U5803 (N_5803,N_4450,N_4914);
nand U5804 (N_5804,N_4492,N_4531);
nor U5805 (N_5805,N_4305,N_4908);
nor U5806 (N_5806,N_4725,N_4866);
or U5807 (N_5807,N_4173,N_4112);
xor U5808 (N_5808,N_4720,N_4430);
or U5809 (N_5809,N_4594,N_4189);
nand U5810 (N_5810,N_4754,N_4770);
and U5811 (N_5811,N_4978,N_4340);
nor U5812 (N_5812,N_4070,N_4498);
nor U5813 (N_5813,N_4276,N_4183);
and U5814 (N_5814,N_4902,N_4862);
or U5815 (N_5815,N_4950,N_4989);
xnor U5816 (N_5816,N_4438,N_4488);
or U5817 (N_5817,N_4000,N_4902);
and U5818 (N_5818,N_4504,N_4407);
nor U5819 (N_5819,N_4155,N_4076);
nand U5820 (N_5820,N_4754,N_4164);
xnor U5821 (N_5821,N_4314,N_4996);
xor U5822 (N_5822,N_4665,N_4271);
or U5823 (N_5823,N_4632,N_4662);
xor U5824 (N_5824,N_4373,N_4017);
or U5825 (N_5825,N_4969,N_4054);
nand U5826 (N_5826,N_4183,N_4932);
nor U5827 (N_5827,N_4993,N_4886);
xor U5828 (N_5828,N_4549,N_4788);
nor U5829 (N_5829,N_4306,N_4762);
nor U5830 (N_5830,N_4949,N_4968);
nand U5831 (N_5831,N_4036,N_4296);
or U5832 (N_5832,N_4503,N_4542);
nand U5833 (N_5833,N_4595,N_4948);
or U5834 (N_5834,N_4226,N_4261);
or U5835 (N_5835,N_4645,N_4872);
xnor U5836 (N_5836,N_4248,N_4222);
nand U5837 (N_5837,N_4964,N_4054);
or U5838 (N_5838,N_4008,N_4117);
and U5839 (N_5839,N_4435,N_4108);
and U5840 (N_5840,N_4395,N_4899);
nand U5841 (N_5841,N_4951,N_4808);
xnor U5842 (N_5842,N_4450,N_4904);
and U5843 (N_5843,N_4604,N_4815);
and U5844 (N_5844,N_4395,N_4368);
nor U5845 (N_5845,N_4977,N_4080);
and U5846 (N_5846,N_4532,N_4184);
xor U5847 (N_5847,N_4170,N_4185);
nor U5848 (N_5848,N_4761,N_4276);
xnor U5849 (N_5849,N_4286,N_4820);
and U5850 (N_5850,N_4775,N_4904);
and U5851 (N_5851,N_4103,N_4567);
xnor U5852 (N_5852,N_4637,N_4460);
xor U5853 (N_5853,N_4261,N_4098);
nand U5854 (N_5854,N_4168,N_4714);
nand U5855 (N_5855,N_4376,N_4142);
xnor U5856 (N_5856,N_4224,N_4190);
nand U5857 (N_5857,N_4930,N_4108);
xnor U5858 (N_5858,N_4842,N_4476);
and U5859 (N_5859,N_4408,N_4393);
or U5860 (N_5860,N_4499,N_4114);
nand U5861 (N_5861,N_4205,N_4980);
nor U5862 (N_5862,N_4258,N_4097);
nor U5863 (N_5863,N_4554,N_4944);
nor U5864 (N_5864,N_4099,N_4828);
nand U5865 (N_5865,N_4433,N_4371);
xnor U5866 (N_5866,N_4596,N_4685);
nor U5867 (N_5867,N_4636,N_4428);
nor U5868 (N_5868,N_4903,N_4304);
and U5869 (N_5869,N_4154,N_4721);
nand U5870 (N_5870,N_4621,N_4038);
xnor U5871 (N_5871,N_4553,N_4426);
nor U5872 (N_5872,N_4028,N_4632);
or U5873 (N_5873,N_4688,N_4270);
nor U5874 (N_5874,N_4439,N_4217);
xnor U5875 (N_5875,N_4918,N_4112);
xor U5876 (N_5876,N_4481,N_4162);
and U5877 (N_5877,N_4987,N_4852);
nor U5878 (N_5878,N_4449,N_4699);
or U5879 (N_5879,N_4406,N_4678);
xor U5880 (N_5880,N_4694,N_4128);
or U5881 (N_5881,N_4755,N_4298);
or U5882 (N_5882,N_4934,N_4453);
and U5883 (N_5883,N_4386,N_4315);
nor U5884 (N_5884,N_4906,N_4455);
xor U5885 (N_5885,N_4258,N_4129);
xor U5886 (N_5886,N_4059,N_4588);
xor U5887 (N_5887,N_4380,N_4888);
nand U5888 (N_5888,N_4623,N_4634);
nand U5889 (N_5889,N_4265,N_4876);
xnor U5890 (N_5890,N_4373,N_4449);
xnor U5891 (N_5891,N_4877,N_4703);
nor U5892 (N_5892,N_4982,N_4850);
nor U5893 (N_5893,N_4171,N_4266);
or U5894 (N_5894,N_4440,N_4891);
and U5895 (N_5895,N_4505,N_4227);
or U5896 (N_5896,N_4833,N_4199);
nand U5897 (N_5897,N_4949,N_4571);
nand U5898 (N_5898,N_4087,N_4365);
nand U5899 (N_5899,N_4005,N_4752);
nor U5900 (N_5900,N_4572,N_4262);
and U5901 (N_5901,N_4209,N_4386);
or U5902 (N_5902,N_4927,N_4632);
nand U5903 (N_5903,N_4960,N_4642);
nand U5904 (N_5904,N_4442,N_4782);
and U5905 (N_5905,N_4864,N_4775);
and U5906 (N_5906,N_4779,N_4414);
and U5907 (N_5907,N_4366,N_4451);
nor U5908 (N_5908,N_4007,N_4796);
nor U5909 (N_5909,N_4180,N_4664);
and U5910 (N_5910,N_4019,N_4177);
xnor U5911 (N_5911,N_4599,N_4442);
or U5912 (N_5912,N_4620,N_4455);
or U5913 (N_5913,N_4355,N_4289);
nor U5914 (N_5914,N_4956,N_4287);
or U5915 (N_5915,N_4772,N_4227);
nand U5916 (N_5916,N_4284,N_4149);
xor U5917 (N_5917,N_4445,N_4414);
and U5918 (N_5918,N_4500,N_4309);
nand U5919 (N_5919,N_4369,N_4882);
xnor U5920 (N_5920,N_4249,N_4271);
nor U5921 (N_5921,N_4192,N_4903);
xor U5922 (N_5922,N_4899,N_4960);
nand U5923 (N_5923,N_4593,N_4972);
or U5924 (N_5924,N_4944,N_4193);
nand U5925 (N_5925,N_4389,N_4809);
nand U5926 (N_5926,N_4209,N_4250);
xor U5927 (N_5927,N_4767,N_4176);
or U5928 (N_5928,N_4754,N_4317);
xnor U5929 (N_5929,N_4011,N_4279);
nand U5930 (N_5930,N_4428,N_4723);
or U5931 (N_5931,N_4462,N_4218);
or U5932 (N_5932,N_4364,N_4158);
or U5933 (N_5933,N_4970,N_4465);
or U5934 (N_5934,N_4166,N_4754);
nand U5935 (N_5935,N_4498,N_4795);
and U5936 (N_5936,N_4863,N_4314);
or U5937 (N_5937,N_4099,N_4992);
xnor U5938 (N_5938,N_4405,N_4596);
and U5939 (N_5939,N_4736,N_4959);
and U5940 (N_5940,N_4203,N_4180);
and U5941 (N_5941,N_4756,N_4123);
nor U5942 (N_5942,N_4811,N_4196);
xor U5943 (N_5943,N_4730,N_4706);
nand U5944 (N_5944,N_4168,N_4820);
or U5945 (N_5945,N_4909,N_4168);
and U5946 (N_5946,N_4470,N_4561);
or U5947 (N_5947,N_4289,N_4654);
nor U5948 (N_5948,N_4020,N_4971);
and U5949 (N_5949,N_4554,N_4809);
and U5950 (N_5950,N_4486,N_4807);
nor U5951 (N_5951,N_4445,N_4325);
xnor U5952 (N_5952,N_4737,N_4133);
or U5953 (N_5953,N_4343,N_4666);
xor U5954 (N_5954,N_4756,N_4797);
nor U5955 (N_5955,N_4861,N_4195);
nand U5956 (N_5956,N_4553,N_4250);
nand U5957 (N_5957,N_4749,N_4195);
or U5958 (N_5958,N_4202,N_4734);
or U5959 (N_5959,N_4222,N_4547);
nand U5960 (N_5960,N_4596,N_4669);
or U5961 (N_5961,N_4068,N_4489);
and U5962 (N_5962,N_4980,N_4525);
xnor U5963 (N_5963,N_4416,N_4936);
nor U5964 (N_5964,N_4166,N_4848);
xor U5965 (N_5965,N_4551,N_4730);
nand U5966 (N_5966,N_4117,N_4472);
xnor U5967 (N_5967,N_4617,N_4188);
nor U5968 (N_5968,N_4196,N_4663);
nand U5969 (N_5969,N_4374,N_4125);
and U5970 (N_5970,N_4473,N_4260);
nor U5971 (N_5971,N_4502,N_4589);
xnor U5972 (N_5972,N_4586,N_4009);
nor U5973 (N_5973,N_4786,N_4598);
and U5974 (N_5974,N_4022,N_4102);
xnor U5975 (N_5975,N_4126,N_4873);
nor U5976 (N_5976,N_4936,N_4482);
xor U5977 (N_5977,N_4638,N_4119);
nand U5978 (N_5978,N_4187,N_4122);
and U5979 (N_5979,N_4099,N_4375);
and U5980 (N_5980,N_4156,N_4336);
nor U5981 (N_5981,N_4810,N_4523);
xnor U5982 (N_5982,N_4127,N_4214);
xnor U5983 (N_5983,N_4979,N_4290);
and U5984 (N_5984,N_4825,N_4327);
nor U5985 (N_5985,N_4691,N_4358);
xor U5986 (N_5986,N_4001,N_4284);
and U5987 (N_5987,N_4003,N_4583);
xnor U5988 (N_5988,N_4773,N_4042);
and U5989 (N_5989,N_4978,N_4085);
nor U5990 (N_5990,N_4493,N_4571);
or U5991 (N_5991,N_4226,N_4099);
and U5992 (N_5992,N_4834,N_4205);
nand U5993 (N_5993,N_4351,N_4863);
nor U5994 (N_5994,N_4658,N_4568);
nor U5995 (N_5995,N_4913,N_4623);
xor U5996 (N_5996,N_4960,N_4238);
or U5997 (N_5997,N_4063,N_4168);
nor U5998 (N_5998,N_4316,N_4160);
and U5999 (N_5999,N_4079,N_4967);
or U6000 (N_6000,N_5750,N_5026);
or U6001 (N_6001,N_5855,N_5652);
nor U6002 (N_6002,N_5924,N_5837);
nand U6003 (N_6003,N_5226,N_5304);
and U6004 (N_6004,N_5248,N_5442);
nand U6005 (N_6005,N_5786,N_5046);
xor U6006 (N_6006,N_5053,N_5806);
nor U6007 (N_6007,N_5292,N_5421);
or U6008 (N_6008,N_5963,N_5899);
xor U6009 (N_6009,N_5504,N_5894);
nand U6010 (N_6010,N_5734,N_5940);
or U6011 (N_6011,N_5757,N_5383);
nor U6012 (N_6012,N_5577,N_5542);
nand U6013 (N_6013,N_5038,N_5281);
xor U6014 (N_6014,N_5785,N_5277);
nor U6015 (N_6015,N_5232,N_5264);
and U6016 (N_6016,N_5994,N_5533);
nand U6017 (N_6017,N_5209,N_5238);
nand U6018 (N_6018,N_5736,N_5344);
nor U6019 (N_6019,N_5787,N_5817);
and U6020 (N_6020,N_5491,N_5326);
nand U6021 (N_6021,N_5562,N_5741);
nor U6022 (N_6022,N_5278,N_5354);
nor U6023 (N_6023,N_5000,N_5916);
and U6024 (N_6024,N_5716,N_5477);
nand U6025 (N_6025,N_5879,N_5372);
and U6026 (N_6026,N_5431,N_5641);
nor U6027 (N_6027,N_5095,N_5211);
and U6028 (N_6028,N_5512,N_5018);
and U6029 (N_6029,N_5833,N_5931);
and U6030 (N_6030,N_5193,N_5124);
nand U6031 (N_6031,N_5460,N_5656);
or U6032 (N_6032,N_5585,N_5358);
xor U6033 (N_6033,N_5721,N_5132);
xnor U6034 (N_6034,N_5195,N_5932);
xor U6035 (N_6035,N_5423,N_5608);
nand U6036 (N_6036,N_5489,N_5543);
nor U6037 (N_6037,N_5307,N_5986);
or U6038 (N_6038,N_5649,N_5265);
nand U6039 (N_6039,N_5328,N_5197);
nand U6040 (N_6040,N_5041,N_5789);
xnor U6041 (N_6041,N_5137,N_5271);
xor U6042 (N_6042,N_5123,N_5602);
nand U6043 (N_6043,N_5039,N_5223);
and U6044 (N_6044,N_5581,N_5591);
nor U6045 (N_6045,N_5346,N_5715);
nor U6046 (N_6046,N_5766,N_5969);
or U6047 (N_6047,N_5306,N_5767);
xnor U6048 (N_6048,N_5490,N_5746);
xnor U6049 (N_6049,N_5037,N_5125);
nand U6050 (N_6050,N_5364,N_5361);
nand U6051 (N_6051,N_5954,N_5952);
or U6052 (N_6052,N_5783,N_5029);
nand U6053 (N_6053,N_5239,N_5711);
nand U6054 (N_6054,N_5389,N_5913);
nand U6055 (N_6055,N_5162,N_5249);
xnor U6056 (N_6056,N_5812,N_5398);
and U6057 (N_6057,N_5973,N_5164);
xor U6058 (N_6058,N_5353,N_5291);
nand U6059 (N_6059,N_5207,N_5293);
or U6060 (N_6060,N_5133,N_5637);
nand U6061 (N_6061,N_5409,N_5866);
nor U6062 (N_6062,N_5513,N_5152);
xnor U6063 (N_6063,N_5296,N_5476);
or U6064 (N_6064,N_5115,N_5961);
nand U6065 (N_6065,N_5544,N_5779);
and U6066 (N_6066,N_5023,N_5747);
or U6067 (N_6067,N_5534,N_5501);
nor U6068 (N_6068,N_5295,N_5206);
nand U6069 (N_6069,N_5427,N_5217);
xor U6070 (N_6070,N_5257,N_5625);
nand U6071 (N_6071,N_5813,N_5836);
xor U6072 (N_6072,N_5488,N_5673);
nand U6073 (N_6073,N_5486,N_5188);
nand U6074 (N_6074,N_5511,N_5834);
nand U6075 (N_6075,N_5025,N_5397);
nor U6076 (N_6076,N_5118,N_5370);
xor U6077 (N_6077,N_5576,N_5844);
xor U6078 (N_6078,N_5689,N_5283);
and U6079 (N_6079,N_5568,N_5998);
nor U6080 (N_6080,N_5744,N_5106);
xnor U6081 (N_6081,N_5301,N_5572);
nand U6082 (N_6082,N_5502,N_5943);
nand U6083 (N_6083,N_5246,N_5791);
or U6084 (N_6084,N_5600,N_5347);
nand U6085 (N_6085,N_5001,N_5237);
or U6086 (N_6086,N_5885,N_5097);
or U6087 (N_6087,N_5334,N_5492);
nor U6088 (N_6088,N_5191,N_5285);
nand U6089 (N_6089,N_5556,N_5500);
nand U6090 (N_6090,N_5590,N_5019);
or U6091 (N_6091,N_5907,N_5739);
or U6092 (N_6092,N_5467,N_5827);
nand U6093 (N_6093,N_5737,N_5979);
xnor U6094 (N_6094,N_5545,N_5064);
or U6095 (N_6095,N_5731,N_5977);
or U6096 (N_6096,N_5129,N_5540);
or U6097 (N_6097,N_5906,N_5367);
and U6098 (N_6098,N_5388,N_5623);
nand U6099 (N_6099,N_5550,N_5377);
or U6100 (N_6100,N_5144,N_5484);
xnor U6101 (N_6101,N_5374,N_5570);
and U6102 (N_6102,N_5036,N_5272);
nand U6103 (N_6103,N_5178,N_5674);
nor U6104 (N_6104,N_5089,N_5874);
or U6105 (N_6105,N_5816,N_5938);
and U6106 (N_6106,N_5901,N_5033);
xor U6107 (N_6107,N_5384,N_5158);
nand U6108 (N_6108,N_5310,N_5840);
nand U6109 (N_6109,N_5098,N_5989);
and U6110 (N_6110,N_5999,N_5558);
or U6111 (N_6111,N_5227,N_5345);
and U6112 (N_6112,N_5267,N_5273);
xnor U6113 (N_6113,N_5761,N_5063);
nand U6114 (N_6114,N_5742,N_5515);
nand U6115 (N_6115,N_5796,N_5980);
nand U6116 (N_6116,N_5122,N_5892);
nand U6117 (N_6117,N_5798,N_5280);
xnor U6118 (N_6118,N_5647,N_5159);
xor U6119 (N_6119,N_5003,N_5831);
nor U6120 (N_6120,N_5128,N_5432);
or U6121 (N_6121,N_5603,N_5911);
and U6122 (N_6122,N_5988,N_5758);
or U6123 (N_6123,N_5915,N_5302);
nor U6124 (N_6124,N_5012,N_5244);
or U6125 (N_6125,N_5852,N_5664);
nor U6126 (N_6126,N_5339,N_5927);
or U6127 (N_6127,N_5470,N_5365);
nand U6128 (N_6128,N_5262,N_5688);
nand U6129 (N_6129,N_5092,N_5618);
and U6130 (N_6130,N_5260,N_5690);
nor U6131 (N_6131,N_5522,N_5803);
xor U6132 (N_6132,N_5100,N_5478);
nand U6133 (N_6133,N_5182,N_5253);
xnor U6134 (N_6134,N_5371,N_5016);
and U6135 (N_6135,N_5826,N_5006);
and U6136 (N_6136,N_5459,N_5946);
or U6137 (N_6137,N_5828,N_5422);
xor U6138 (N_6138,N_5775,N_5765);
nor U6139 (N_6139,N_5996,N_5538);
and U6140 (N_6140,N_5677,N_5331);
and U6141 (N_6141,N_5043,N_5040);
nand U6142 (N_6142,N_5447,N_5536);
or U6143 (N_6143,N_5517,N_5587);
nand U6144 (N_6144,N_5663,N_5241);
and U6145 (N_6145,N_5546,N_5103);
or U6146 (N_6146,N_5763,N_5903);
xnor U6147 (N_6147,N_5982,N_5058);
xnor U6148 (N_6148,N_5069,N_5628);
nand U6149 (N_6149,N_5311,N_5658);
nor U6150 (N_6150,N_5090,N_5465);
nand U6151 (N_6151,N_5781,N_5147);
xor U6152 (N_6152,N_5096,N_5975);
nor U6153 (N_6153,N_5612,N_5030);
xor U6154 (N_6154,N_5774,N_5532);
nor U6155 (N_6155,N_5771,N_5926);
xnor U6156 (N_6156,N_5059,N_5263);
nand U6157 (N_6157,N_5357,N_5843);
and U6158 (N_6158,N_5565,N_5528);
nand U6159 (N_6159,N_5596,N_5194);
and U6160 (N_6160,N_5024,N_5413);
nor U6161 (N_6161,N_5317,N_5846);
and U6162 (N_6162,N_5450,N_5127);
nand U6163 (N_6163,N_5126,N_5896);
nand U6164 (N_6164,N_5314,N_5464);
nor U6165 (N_6165,N_5107,N_5212);
xor U6166 (N_6166,N_5718,N_5589);
xnor U6167 (N_6167,N_5245,N_5156);
or U6168 (N_6168,N_5815,N_5939);
or U6169 (N_6169,N_5017,N_5050);
and U6170 (N_6170,N_5526,N_5898);
nand U6171 (N_6171,N_5480,N_5325);
and U6172 (N_6172,N_5804,N_5385);
nand U6173 (N_6173,N_5944,N_5738);
or U6174 (N_6174,N_5108,N_5112);
xnor U6175 (N_6175,N_5205,N_5120);
nand U6176 (N_6176,N_5160,N_5379);
xor U6177 (N_6177,N_5167,N_5613);
or U6178 (N_6178,N_5466,N_5706);
xor U6179 (N_6179,N_5527,N_5822);
nand U6180 (N_6180,N_5407,N_5093);
nand U6181 (N_6181,N_5079,N_5266);
and U6182 (N_6182,N_5857,N_5682);
or U6183 (N_6183,N_5675,N_5609);
xnor U6184 (N_6184,N_5957,N_5258);
nor U6185 (N_6185,N_5644,N_5199);
xor U6186 (N_6186,N_5552,N_5729);
nor U6187 (N_6187,N_5131,N_5770);
nand U6188 (N_6188,N_5010,N_5936);
and U6189 (N_6189,N_5055,N_5062);
or U6190 (N_6190,N_5710,N_5506);
and U6191 (N_6191,N_5672,N_5780);
nor U6192 (N_6192,N_5387,N_5453);
or U6193 (N_6193,N_5066,N_5700);
nand U6194 (N_6194,N_5446,N_5820);
nor U6195 (N_6195,N_5308,N_5028);
and U6196 (N_6196,N_5851,N_5567);
nand U6197 (N_6197,N_5768,N_5743);
or U6198 (N_6198,N_5825,N_5784);
and U6199 (N_6199,N_5524,N_5138);
nand U6200 (N_6200,N_5369,N_5027);
nor U6201 (N_6201,N_5523,N_5376);
nand U6202 (N_6202,N_5518,N_5005);
or U6203 (N_6203,N_5252,N_5145);
nand U6204 (N_6204,N_5276,N_5286);
and U6205 (N_6205,N_5493,N_5454);
and U6206 (N_6206,N_5760,N_5720);
nand U6207 (N_6207,N_5222,N_5275);
nand U6208 (N_6208,N_5510,N_5990);
or U6209 (N_6209,N_5707,N_5274);
nand U6210 (N_6210,N_5614,N_5751);
xor U6211 (N_6211,N_5337,N_5897);
or U6212 (N_6212,N_5333,N_5404);
and U6213 (N_6213,N_5799,N_5714);
xor U6214 (N_6214,N_5964,N_5693);
nand U6215 (N_6215,N_5660,N_5261);
xnor U6216 (N_6216,N_5196,N_5335);
nor U6217 (N_6217,N_5149,N_5597);
nor U6218 (N_6218,N_5947,N_5918);
xnor U6219 (N_6219,N_5330,N_5582);
or U6220 (N_6220,N_5400,N_5895);
nor U6221 (N_6221,N_5588,N_5074);
and U6222 (N_6222,N_5636,N_5171);
nor U6223 (N_6223,N_5514,N_5200);
nor U6224 (N_6224,N_5179,N_5800);
nand U6225 (N_6225,N_5111,N_5529);
nand U6226 (N_6226,N_5322,N_5153);
nor U6227 (N_6227,N_5060,N_5724);
xor U6228 (N_6228,N_5324,N_5551);
nand U6229 (N_6229,N_5651,N_5399);
nor U6230 (N_6230,N_5530,N_5920);
nor U6231 (N_6231,N_5805,N_5284);
xor U6232 (N_6232,N_5181,N_5495);
or U6233 (N_6233,N_5878,N_5829);
nor U6234 (N_6234,N_5250,N_5270);
and U6235 (N_6235,N_5554,N_5624);
and U6236 (N_6236,N_5441,N_5221);
nand U6237 (N_6237,N_5329,N_5049);
xor U6238 (N_6238,N_5104,N_5881);
nor U6239 (N_6239,N_5219,N_5792);
nor U6240 (N_6240,N_5359,N_5838);
nand U6241 (N_6241,N_5189,N_5289);
and U6242 (N_6242,N_5279,N_5015);
and U6243 (N_6243,N_5726,N_5633);
nand U6244 (N_6244,N_5452,N_5368);
xor U6245 (N_6245,N_5653,N_5935);
xnor U6246 (N_6246,N_5841,N_5659);
nand U6247 (N_6247,N_5891,N_5919);
or U6248 (N_6248,N_5474,N_5229);
nor U6249 (N_6249,N_5605,N_5893);
or U6250 (N_6250,N_5198,N_5864);
xnor U6251 (N_6251,N_5351,N_5818);
and U6252 (N_6252,N_5186,N_5071);
or U6253 (N_6253,N_5748,N_5076);
nand U6254 (N_6254,N_5615,N_5457);
xor U6255 (N_6255,N_5349,N_5627);
nor U6256 (N_6256,N_5394,N_5231);
nor U6257 (N_6257,N_5290,N_5356);
and U6258 (N_6258,N_5561,N_5797);
and U6259 (N_6259,N_5436,N_5886);
or U6260 (N_6260,N_5665,N_5061);
and U6261 (N_6261,N_5643,N_5642);
xor U6262 (N_6262,N_5418,N_5560);
nand U6263 (N_6263,N_5119,N_5190);
xnor U6264 (N_6264,N_5044,N_5856);
xor U6265 (N_6265,N_5469,N_5676);
and U6266 (N_6266,N_5396,N_5505);
xnor U6267 (N_6267,N_5472,N_5539);
nor U6268 (N_6268,N_5704,N_5146);
xor U6269 (N_6269,N_5233,N_5516);
xnor U6270 (N_6270,N_5599,N_5109);
nand U6271 (N_6271,N_5553,N_5574);
xnor U6272 (N_6272,N_5559,N_5811);
nor U6273 (N_6273,N_5788,N_5686);
or U6274 (N_6274,N_5719,N_5121);
or U6275 (N_6275,N_5875,N_5177);
and U6276 (N_6276,N_5860,N_5993);
nor U6277 (N_6277,N_5052,N_5419);
and U6278 (N_6278,N_5320,N_5773);
and U6279 (N_6279,N_5303,N_5315);
or U6280 (N_6280,N_5762,N_5141);
or U6281 (N_6281,N_5616,N_5619);
xor U6282 (N_6282,N_5639,N_5795);
nand U6283 (N_6283,N_5575,N_5392);
nor U6284 (N_6284,N_5657,N_5976);
and U6285 (N_6285,N_5360,N_5862);
or U6286 (N_6286,N_5509,N_5908);
and U6287 (N_6287,N_5338,N_5687);
xor U6288 (N_6288,N_5201,N_5620);
or U6289 (N_6289,N_5921,N_5953);
and U6290 (N_6290,N_5905,N_5378);
xnor U6291 (N_6291,N_5978,N_5727);
or U6292 (N_6292,N_5228,N_5630);
nor U6293 (N_6293,N_5814,N_5685);
nand U6294 (N_6294,N_5631,N_5402);
xor U6295 (N_6295,N_5494,N_5305);
or U6296 (N_6296,N_5410,N_5547);
or U6297 (N_6297,N_5849,N_5697);
xor U6298 (N_6298,N_5088,N_5117);
nand U6299 (N_6299,N_5548,N_5184);
nand U6300 (N_6300,N_5332,N_5202);
and U6301 (N_6301,N_5832,N_5793);
or U6302 (N_6302,N_5081,N_5535);
xor U6303 (N_6303,N_5669,N_5667);
and U6304 (N_6304,N_5342,N_5435);
nand U6305 (N_6305,N_5150,N_5065);
nor U6306 (N_6306,N_5225,N_5116);
nor U6307 (N_6307,N_5080,N_5888);
and U6308 (N_6308,N_5958,N_5395);
nand U6309 (N_6309,N_5949,N_5297);
xor U6310 (N_6310,N_5702,N_5809);
and U6311 (N_6311,N_5728,N_5531);
or U6312 (N_6312,N_5443,N_5777);
nor U6313 (N_6313,N_5845,N_5869);
nor U6314 (N_6314,N_5414,N_5113);
xnor U6315 (N_6315,N_5403,N_5287);
or U6316 (N_6316,N_5580,N_5573);
or U6317 (N_6317,N_5730,N_5269);
or U6318 (N_6318,N_5316,N_5722);
or U6319 (N_6319,N_5645,N_5887);
and U6320 (N_6320,N_5853,N_5444);
or U6321 (N_6321,N_5481,N_5890);
nor U6322 (N_6322,N_5135,N_5930);
nor U6323 (N_6323,N_5130,N_5406);
or U6324 (N_6324,N_5482,N_5327);
xnor U6325 (N_6325,N_5366,N_5699);
nand U6326 (N_6326,N_5723,N_5604);
and U6327 (N_6327,N_5870,N_5503);
nor U6328 (N_6328,N_5070,N_5756);
and U6329 (N_6329,N_5009,N_5067);
xnor U6330 (N_6330,N_5230,N_5912);
nor U6331 (N_6331,N_5057,N_5640);
xor U6332 (N_6332,N_5312,N_5725);
xnor U6333 (N_6333,N_5499,N_5696);
nor U6334 (N_6334,N_5210,N_5584);
nand U6335 (N_6335,N_5821,N_5967);
nor U6336 (N_6336,N_5752,N_5951);
and U6337 (N_6337,N_5078,N_5790);
nor U6338 (N_6338,N_5968,N_5703);
or U6339 (N_6339,N_5684,N_5749);
and U6340 (N_6340,N_5175,N_5995);
or U6341 (N_6341,N_5610,N_5085);
xnor U6342 (N_6342,N_5110,N_5847);
or U6343 (N_6343,N_5617,N_5169);
or U6344 (N_6344,N_5165,N_5498);
xor U6345 (N_6345,N_5075,N_5634);
or U6346 (N_6346,N_5426,N_5022);
or U6347 (N_6347,N_5084,N_5835);
or U6348 (N_6348,N_5013,N_5872);
xor U6349 (N_6349,N_5754,N_5068);
or U6350 (N_6350,N_5868,N_5321);
or U6351 (N_6351,N_5842,N_5794);
and U6352 (N_6352,N_5479,N_5678);
xor U6353 (N_6353,N_5401,N_5655);
nor U6354 (N_6354,N_5965,N_5519);
nand U6355 (N_6355,N_5091,N_5031);
or U6356 (N_6356,N_5288,N_5143);
nand U6357 (N_6357,N_5923,N_5801);
or U6358 (N_6358,N_5213,N_5654);
nor U6359 (N_6359,N_5858,N_5298);
or U6360 (N_6360,N_5440,N_5668);
and U6361 (N_6361,N_5214,N_5701);
nor U6362 (N_6362,N_5176,N_5411);
nand U6363 (N_6363,N_5139,N_5564);
nand U6364 (N_6364,N_5830,N_5437);
or U6365 (N_6365,N_5309,N_5082);
nand U6366 (N_6366,N_5772,N_5808);
nor U6367 (N_6367,N_5537,N_5487);
nor U6368 (N_6368,N_5224,N_5373);
or U6369 (N_6369,N_5451,N_5984);
nand U6370 (N_6370,N_5236,N_5823);
nor U6371 (N_6371,N_5099,N_5987);
or U6372 (N_6372,N_5174,N_5424);
and U6373 (N_6373,N_5047,N_5635);
nand U6374 (N_6374,N_5735,N_5740);
nor U6375 (N_6375,N_5569,N_5458);
nor U6376 (N_6376,N_5319,N_5971);
nand U6377 (N_6377,N_5042,N_5732);
xor U6378 (N_6378,N_5733,N_5712);
and U6379 (N_6379,N_5077,N_5889);
nor U6380 (N_6380,N_5172,N_5708);
nor U6381 (N_6381,N_5363,N_5632);
xor U6382 (N_6382,N_5242,N_5004);
xor U6383 (N_6383,N_5698,N_5168);
and U6384 (N_6384,N_5592,N_5045);
nand U6385 (N_6385,N_5382,N_5336);
nand U6386 (N_6386,N_5883,N_5863);
and U6387 (N_6387,N_5586,N_5170);
and U6388 (N_6388,N_5094,N_5475);
nand U6389 (N_6389,N_5166,N_5163);
xor U6390 (N_6390,N_5782,N_5180);
nand U6391 (N_6391,N_5646,N_5429);
or U6392 (N_6392,N_5463,N_5549);
nor U6393 (N_6393,N_5848,N_5350);
nor U6394 (N_6394,N_5914,N_5933);
nor U6395 (N_6395,N_5393,N_5854);
nor U6396 (N_6396,N_5216,N_5520);
nor U6397 (N_6397,N_5485,N_5680);
nand U6398 (N_6398,N_5871,N_5102);
xor U6399 (N_6399,N_5900,N_5681);
nand U6400 (N_6400,N_5611,N_5405);
xor U6401 (N_6401,N_5629,N_5415);
xor U6402 (N_6402,N_5694,N_5254);
nand U6403 (N_6403,N_5034,N_5850);
and U6404 (N_6404,N_5755,N_5557);
xnor U6405 (N_6405,N_5861,N_5621);
nor U6406 (N_6406,N_5234,N_5622);
xnor U6407 (N_6407,N_5997,N_5884);
and U6408 (N_6408,N_5243,N_5445);
and U6409 (N_6409,N_5220,N_5648);
nand U6410 (N_6410,N_5962,N_5521);
nand U6411 (N_6411,N_5937,N_5929);
nand U6412 (N_6412,N_5456,N_5934);
and U6413 (N_6413,N_5764,N_5268);
and U6414 (N_6414,N_5666,N_5048);
or U6415 (N_6415,N_5140,N_5300);
nor U6416 (N_6416,N_5497,N_5468);
nand U6417 (N_6417,N_5555,N_5776);
xor U6418 (N_6418,N_5105,N_5192);
nand U6419 (N_6419,N_5101,N_5991);
nand U6420 (N_6420,N_5380,N_5318);
or U6421 (N_6421,N_5679,N_5683);
nor U6422 (N_6422,N_5910,N_5461);
nand U6423 (N_6423,N_5525,N_5972);
and U6424 (N_6424,N_5218,N_5807);
xor U6425 (N_6425,N_5208,N_5970);
xnor U6426 (N_6426,N_5087,N_5425);
or U6427 (N_6427,N_5769,N_5839);
xnor U6428 (N_6428,N_5626,N_5985);
or U6429 (N_6429,N_5428,N_5709);
and U6430 (N_6430,N_5873,N_5661);
xor U6431 (N_6431,N_5434,N_5928);
nand U6432 (N_6432,N_5313,N_5439);
and U6433 (N_6433,N_5323,N_5607);
xor U6434 (N_6434,N_5416,N_5578);
or U6435 (N_6435,N_5011,N_5981);
nor U6436 (N_6436,N_5114,N_5593);
nand U6437 (N_6437,N_5391,N_5902);
or U6438 (N_6438,N_5183,N_5185);
nor U6439 (N_6439,N_5598,N_5083);
nand U6440 (N_6440,N_5959,N_5705);
or U6441 (N_6441,N_5381,N_5983);
xor U6442 (N_6442,N_5072,N_5375);
or U6443 (N_6443,N_5922,N_5571);
nand U6444 (N_6444,N_5778,N_5294);
nor U6445 (N_6445,N_5007,N_5151);
and U6446 (N_6446,N_5204,N_5215);
and U6447 (N_6447,N_5235,N_5362);
or U6448 (N_6448,N_5203,N_5819);
nor U6449 (N_6449,N_5438,N_5867);
or U6450 (N_6450,N_5073,N_5240);
and U6451 (N_6451,N_5810,N_5148);
nand U6452 (N_6452,N_5054,N_5154);
xor U6453 (N_6453,N_5904,N_5247);
nand U6454 (N_6454,N_5021,N_5355);
and U6455 (N_6455,N_5594,N_5541);
or U6456 (N_6456,N_5691,N_5753);
nor U6457 (N_6457,N_5941,N_5256);
nor U6458 (N_6458,N_5483,N_5601);
xnor U6459 (N_6459,N_5759,N_5909);
and U6460 (N_6460,N_5950,N_5865);
and U6461 (N_6461,N_5448,N_5882);
nor U6462 (N_6462,N_5161,N_5086);
nand U6463 (N_6463,N_5255,N_5583);
nand U6464 (N_6464,N_5142,N_5638);
nor U6465 (N_6465,N_5917,N_5449);
or U6466 (N_6466,N_5251,N_5157);
or U6467 (N_6467,N_5455,N_5876);
nor U6468 (N_6468,N_5948,N_5430);
xor U6469 (N_6469,N_5992,N_5408);
and U6470 (N_6470,N_5173,N_5566);
nor U6471 (N_6471,N_5462,N_5956);
nor U6472 (N_6472,N_5877,N_5299);
or U6473 (N_6473,N_5051,N_5966);
and U6474 (N_6474,N_5341,N_5348);
nor U6475 (N_6475,N_5420,N_5670);
and U6476 (N_6476,N_5859,N_5745);
nor U6477 (N_6477,N_5134,N_5925);
xnor U6478 (N_6478,N_5671,N_5136);
or U6479 (N_6479,N_5945,N_5717);
or U6480 (N_6480,N_5650,N_5417);
or U6481 (N_6481,N_5433,N_5032);
or U6482 (N_6482,N_5386,N_5606);
or U6483 (N_6483,N_5187,N_5802);
or U6484 (N_6484,N_5960,N_5390);
nor U6485 (N_6485,N_5955,N_5496);
xnor U6486 (N_6486,N_5020,N_5352);
nor U6487 (N_6487,N_5259,N_5014);
or U6488 (N_6488,N_5595,N_5008);
xnor U6489 (N_6489,N_5579,N_5056);
xor U6490 (N_6490,N_5002,N_5035);
or U6491 (N_6491,N_5880,N_5507);
xnor U6492 (N_6492,N_5282,N_5563);
nand U6493 (N_6493,N_5824,N_5412);
nand U6494 (N_6494,N_5662,N_5942);
or U6495 (N_6495,N_5155,N_5473);
xor U6496 (N_6496,N_5713,N_5343);
xnor U6497 (N_6497,N_5692,N_5340);
nor U6498 (N_6498,N_5471,N_5695);
nor U6499 (N_6499,N_5508,N_5974);
nand U6500 (N_6500,N_5196,N_5798);
xor U6501 (N_6501,N_5171,N_5384);
xor U6502 (N_6502,N_5524,N_5750);
or U6503 (N_6503,N_5823,N_5321);
or U6504 (N_6504,N_5020,N_5082);
and U6505 (N_6505,N_5317,N_5965);
nand U6506 (N_6506,N_5348,N_5768);
nor U6507 (N_6507,N_5281,N_5070);
or U6508 (N_6508,N_5977,N_5324);
xor U6509 (N_6509,N_5685,N_5290);
nor U6510 (N_6510,N_5222,N_5985);
and U6511 (N_6511,N_5823,N_5929);
nand U6512 (N_6512,N_5162,N_5966);
and U6513 (N_6513,N_5778,N_5187);
and U6514 (N_6514,N_5147,N_5211);
and U6515 (N_6515,N_5766,N_5917);
xnor U6516 (N_6516,N_5672,N_5294);
nand U6517 (N_6517,N_5120,N_5506);
or U6518 (N_6518,N_5316,N_5647);
nand U6519 (N_6519,N_5321,N_5714);
or U6520 (N_6520,N_5975,N_5016);
and U6521 (N_6521,N_5318,N_5546);
nand U6522 (N_6522,N_5635,N_5928);
nor U6523 (N_6523,N_5192,N_5770);
nand U6524 (N_6524,N_5130,N_5876);
and U6525 (N_6525,N_5842,N_5719);
and U6526 (N_6526,N_5083,N_5299);
nor U6527 (N_6527,N_5433,N_5161);
nand U6528 (N_6528,N_5383,N_5631);
and U6529 (N_6529,N_5152,N_5201);
xnor U6530 (N_6530,N_5953,N_5470);
nand U6531 (N_6531,N_5918,N_5073);
xnor U6532 (N_6532,N_5496,N_5609);
nor U6533 (N_6533,N_5879,N_5522);
nand U6534 (N_6534,N_5267,N_5593);
nor U6535 (N_6535,N_5155,N_5811);
xnor U6536 (N_6536,N_5389,N_5664);
nand U6537 (N_6537,N_5634,N_5172);
nor U6538 (N_6538,N_5451,N_5847);
or U6539 (N_6539,N_5146,N_5545);
and U6540 (N_6540,N_5479,N_5882);
or U6541 (N_6541,N_5478,N_5295);
and U6542 (N_6542,N_5296,N_5069);
nand U6543 (N_6543,N_5913,N_5859);
xnor U6544 (N_6544,N_5013,N_5342);
xnor U6545 (N_6545,N_5960,N_5236);
nor U6546 (N_6546,N_5692,N_5558);
and U6547 (N_6547,N_5658,N_5594);
and U6548 (N_6548,N_5207,N_5560);
or U6549 (N_6549,N_5661,N_5503);
or U6550 (N_6550,N_5575,N_5098);
and U6551 (N_6551,N_5733,N_5729);
nand U6552 (N_6552,N_5120,N_5648);
xor U6553 (N_6553,N_5432,N_5237);
nor U6554 (N_6554,N_5143,N_5692);
nand U6555 (N_6555,N_5604,N_5889);
and U6556 (N_6556,N_5006,N_5855);
xor U6557 (N_6557,N_5165,N_5904);
and U6558 (N_6558,N_5103,N_5289);
nor U6559 (N_6559,N_5265,N_5692);
xor U6560 (N_6560,N_5110,N_5313);
and U6561 (N_6561,N_5495,N_5246);
or U6562 (N_6562,N_5867,N_5140);
or U6563 (N_6563,N_5869,N_5635);
nand U6564 (N_6564,N_5437,N_5396);
and U6565 (N_6565,N_5756,N_5550);
nor U6566 (N_6566,N_5813,N_5657);
and U6567 (N_6567,N_5157,N_5518);
xnor U6568 (N_6568,N_5163,N_5915);
xnor U6569 (N_6569,N_5608,N_5882);
or U6570 (N_6570,N_5192,N_5432);
and U6571 (N_6571,N_5133,N_5311);
xnor U6572 (N_6572,N_5409,N_5271);
or U6573 (N_6573,N_5933,N_5196);
and U6574 (N_6574,N_5972,N_5416);
nor U6575 (N_6575,N_5074,N_5683);
nand U6576 (N_6576,N_5959,N_5950);
and U6577 (N_6577,N_5248,N_5293);
nand U6578 (N_6578,N_5496,N_5182);
or U6579 (N_6579,N_5188,N_5717);
nor U6580 (N_6580,N_5604,N_5975);
and U6581 (N_6581,N_5096,N_5036);
and U6582 (N_6582,N_5488,N_5306);
nor U6583 (N_6583,N_5423,N_5599);
xor U6584 (N_6584,N_5417,N_5209);
nand U6585 (N_6585,N_5418,N_5626);
nor U6586 (N_6586,N_5793,N_5813);
and U6587 (N_6587,N_5369,N_5332);
nand U6588 (N_6588,N_5974,N_5904);
xor U6589 (N_6589,N_5715,N_5358);
and U6590 (N_6590,N_5209,N_5005);
and U6591 (N_6591,N_5489,N_5479);
and U6592 (N_6592,N_5686,N_5051);
xor U6593 (N_6593,N_5269,N_5417);
and U6594 (N_6594,N_5438,N_5372);
nand U6595 (N_6595,N_5485,N_5389);
xor U6596 (N_6596,N_5477,N_5366);
and U6597 (N_6597,N_5937,N_5691);
or U6598 (N_6598,N_5779,N_5576);
nor U6599 (N_6599,N_5557,N_5842);
nor U6600 (N_6600,N_5172,N_5980);
nand U6601 (N_6601,N_5678,N_5448);
nand U6602 (N_6602,N_5943,N_5554);
nor U6603 (N_6603,N_5678,N_5852);
nand U6604 (N_6604,N_5631,N_5087);
nor U6605 (N_6605,N_5371,N_5715);
and U6606 (N_6606,N_5788,N_5044);
nand U6607 (N_6607,N_5225,N_5189);
nand U6608 (N_6608,N_5867,N_5806);
xnor U6609 (N_6609,N_5937,N_5515);
nand U6610 (N_6610,N_5206,N_5181);
nor U6611 (N_6611,N_5173,N_5672);
nor U6612 (N_6612,N_5238,N_5461);
and U6613 (N_6613,N_5571,N_5980);
nand U6614 (N_6614,N_5932,N_5789);
and U6615 (N_6615,N_5325,N_5429);
nor U6616 (N_6616,N_5563,N_5300);
nor U6617 (N_6617,N_5232,N_5362);
nor U6618 (N_6618,N_5872,N_5787);
xnor U6619 (N_6619,N_5911,N_5860);
nand U6620 (N_6620,N_5783,N_5983);
and U6621 (N_6621,N_5262,N_5551);
xor U6622 (N_6622,N_5050,N_5574);
or U6623 (N_6623,N_5914,N_5928);
xnor U6624 (N_6624,N_5209,N_5415);
xnor U6625 (N_6625,N_5110,N_5929);
and U6626 (N_6626,N_5739,N_5839);
and U6627 (N_6627,N_5535,N_5967);
or U6628 (N_6628,N_5791,N_5011);
or U6629 (N_6629,N_5653,N_5964);
xor U6630 (N_6630,N_5317,N_5474);
or U6631 (N_6631,N_5636,N_5290);
and U6632 (N_6632,N_5565,N_5504);
nand U6633 (N_6633,N_5307,N_5170);
nand U6634 (N_6634,N_5884,N_5996);
or U6635 (N_6635,N_5581,N_5536);
or U6636 (N_6636,N_5028,N_5738);
nor U6637 (N_6637,N_5751,N_5961);
or U6638 (N_6638,N_5205,N_5513);
or U6639 (N_6639,N_5891,N_5214);
and U6640 (N_6640,N_5933,N_5663);
and U6641 (N_6641,N_5931,N_5839);
nand U6642 (N_6642,N_5297,N_5577);
nand U6643 (N_6643,N_5737,N_5354);
xnor U6644 (N_6644,N_5387,N_5842);
and U6645 (N_6645,N_5709,N_5009);
and U6646 (N_6646,N_5222,N_5870);
nor U6647 (N_6647,N_5728,N_5614);
or U6648 (N_6648,N_5003,N_5463);
and U6649 (N_6649,N_5118,N_5685);
nand U6650 (N_6650,N_5073,N_5657);
or U6651 (N_6651,N_5255,N_5575);
nand U6652 (N_6652,N_5795,N_5652);
xor U6653 (N_6653,N_5574,N_5345);
xor U6654 (N_6654,N_5324,N_5745);
nand U6655 (N_6655,N_5421,N_5669);
and U6656 (N_6656,N_5109,N_5143);
xor U6657 (N_6657,N_5024,N_5517);
nand U6658 (N_6658,N_5643,N_5388);
xor U6659 (N_6659,N_5916,N_5983);
nand U6660 (N_6660,N_5405,N_5152);
or U6661 (N_6661,N_5943,N_5410);
nand U6662 (N_6662,N_5743,N_5140);
xnor U6663 (N_6663,N_5425,N_5118);
or U6664 (N_6664,N_5810,N_5348);
nand U6665 (N_6665,N_5189,N_5371);
and U6666 (N_6666,N_5009,N_5493);
nor U6667 (N_6667,N_5235,N_5250);
nand U6668 (N_6668,N_5050,N_5620);
nand U6669 (N_6669,N_5782,N_5486);
nor U6670 (N_6670,N_5131,N_5287);
and U6671 (N_6671,N_5801,N_5764);
nand U6672 (N_6672,N_5871,N_5904);
xnor U6673 (N_6673,N_5866,N_5622);
and U6674 (N_6674,N_5586,N_5656);
and U6675 (N_6675,N_5081,N_5096);
or U6676 (N_6676,N_5172,N_5480);
and U6677 (N_6677,N_5500,N_5820);
xor U6678 (N_6678,N_5653,N_5956);
or U6679 (N_6679,N_5814,N_5686);
nand U6680 (N_6680,N_5096,N_5297);
and U6681 (N_6681,N_5674,N_5363);
and U6682 (N_6682,N_5431,N_5609);
and U6683 (N_6683,N_5128,N_5902);
nand U6684 (N_6684,N_5455,N_5173);
nand U6685 (N_6685,N_5181,N_5266);
and U6686 (N_6686,N_5319,N_5659);
nand U6687 (N_6687,N_5895,N_5872);
nand U6688 (N_6688,N_5100,N_5675);
nand U6689 (N_6689,N_5467,N_5440);
nor U6690 (N_6690,N_5344,N_5638);
and U6691 (N_6691,N_5316,N_5552);
and U6692 (N_6692,N_5853,N_5955);
xor U6693 (N_6693,N_5901,N_5790);
nand U6694 (N_6694,N_5032,N_5542);
xnor U6695 (N_6695,N_5961,N_5462);
xor U6696 (N_6696,N_5999,N_5696);
and U6697 (N_6697,N_5321,N_5810);
or U6698 (N_6698,N_5806,N_5086);
and U6699 (N_6699,N_5083,N_5636);
nand U6700 (N_6700,N_5920,N_5103);
xor U6701 (N_6701,N_5385,N_5122);
and U6702 (N_6702,N_5748,N_5747);
nor U6703 (N_6703,N_5976,N_5337);
nand U6704 (N_6704,N_5512,N_5867);
xor U6705 (N_6705,N_5351,N_5417);
nand U6706 (N_6706,N_5427,N_5627);
and U6707 (N_6707,N_5076,N_5200);
nor U6708 (N_6708,N_5540,N_5178);
nor U6709 (N_6709,N_5972,N_5681);
or U6710 (N_6710,N_5492,N_5944);
or U6711 (N_6711,N_5951,N_5083);
nor U6712 (N_6712,N_5111,N_5562);
and U6713 (N_6713,N_5093,N_5042);
or U6714 (N_6714,N_5090,N_5538);
or U6715 (N_6715,N_5108,N_5722);
nand U6716 (N_6716,N_5789,N_5649);
or U6717 (N_6717,N_5607,N_5582);
nor U6718 (N_6718,N_5247,N_5541);
xnor U6719 (N_6719,N_5332,N_5198);
or U6720 (N_6720,N_5144,N_5887);
nor U6721 (N_6721,N_5755,N_5935);
nand U6722 (N_6722,N_5185,N_5148);
xnor U6723 (N_6723,N_5005,N_5166);
nand U6724 (N_6724,N_5691,N_5101);
nand U6725 (N_6725,N_5551,N_5507);
or U6726 (N_6726,N_5564,N_5762);
nor U6727 (N_6727,N_5169,N_5847);
nand U6728 (N_6728,N_5667,N_5082);
or U6729 (N_6729,N_5825,N_5713);
xnor U6730 (N_6730,N_5368,N_5614);
xnor U6731 (N_6731,N_5315,N_5058);
nor U6732 (N_6732,N_5889,N_5905);
nand U6733 (N_6733,N_5361,N_5672);
and U6734 (N_6734,N_5828,N_5796);
nand U6735 (N_6735,N_5448,N_5245);
xnor U6736 (N_6736,N_5404,N_5294);
nor U6737 (N_6737,N_5771,N_5628);
and U6738 (N_6738,N_5624,N_5779);
nand U6739 (N_6739,N_5824,N_5426);
or U6740 (N_6740,N_5366,N_5687);
nand U6741 (N_6741,N_5994,N_5957);
nor U6742 (N_6742,N_5290,N_5697);
nand U6743 (N_6743,N_5188,N_5226);
nand U6744 (N_6744,N_5224,N_5848);
nor U6745 (N_6745,N_5160,N_5139);
or U6746 (N_6746,N_5464,N_5129);
nor U6747 (N_6747,N_5856,N_5693);
or U6748 (N_6748,N_5989,N_5084);
nor U6749 (N_6749,N_5643,N_5711);
or U6750 (N_6750,N_5787,N_5656);
xnor U6751 (N_6751,N_5596,N_5024);
nand U6752 (N_6752,N_5306,N_5558);
or U6753 (N_6753,N_5567,N_5960);
or U6754 (N_6754,N_5104,N_5405);
xnor U6755 (N_6755,N_5621,N_5180);
nor U6756 (N_6756,N_5852,N_5218);
nor U6757 (N_6757,N_5954,N_5249);
and U6758 (N_6758,N_5121,N_5400);
xnor U6759 (N_6759,N_5823,N_5162);
nor U6760 (N_6760,N_5356,N_5624);
and U6761 (N_6761,N_5952,N_5936);
or U6762 (N_6762,N_5193,N_5108);
and U6763 (N_6763,N_5365,N_5082);
nor U6764 (N_6764,N_5035,N_5813);
nand U6765 (N_6765,N_5725,N_5184);
and U6766 (N_6766,N_5413,N_5756);
xnor U6767 (N_6767,N_5944,N_5826);
or U6768 (N_6768,N_5012,N_5993);
xnor U6769 (N_6769,N_5709,N_5311);
and U6770 (N_6770,N_5912,N_5811);
xnor U6771 (N_6771,N_5970,N_5474);
and U6772 (N_6772,N_5832,N_5115);
xnor U6773 (N_6773,N_5681,N_5421);
xor U6774 (N_6774,N_5089,N_5201);
and U6775 (N_6775,N_5587,N_5077);
or U6776 (N_6776,N_5624,N_5718);
nor U6777 (N_6777,N_5676,N_5285);
nor U6778 (N_6778,N_5076,N_5082);
nor U6779 (N_6779,N_5596,N_5965);
nand U6780 (N_6780,N_5198,N_5329);
or U6781 (N_6781,N_5091,N_5117);
nand U6782 (N_6782,N_5290,N_5450);
or U6783 (N_6783,N_5582,N_5618);
nor U6784 (N_6784,N_5194,N_5329);
nand U6785 (N_6785,N_5738,N_5718);
nand U6786 (N_6786,N_5066,N_5743);
or U6787 (N_6787,N_5879,N_5186);
or U6788 (N_6788,N_5684,N_5584);
nand U6789 (N_6789,N_5619,N_5383);
nor U6790 (N_6790,N_5099,N_5904);
or U6791 (N_6791,N_5396,N_5207);
and U6792 (N_6792,N_5002,N_5206);
or U6793 (N_6793,N_5893,N_5689);
and U6794 (N_6794,N_5178,N_5986);
nor U6795 (N_6795,N_5396,N_5008);
or U6796 (N_6796,N_5935,N_5236);
or U6797 (N_6797,N_5511,N_5072);
xnor U6798 (N_6798,N_5330,N_5781);
nand U6799 (N_6799,N_5429,N_5205);
nor U6800 (N_6800,N_5531,N_5365);
xnor U6801 (N_6801,N_5342,N_5027);
xor U6802 (N_6802,N_5317,N_5647);
or U6803 (N_6803,N_5290,N_5068);
nand U6804 (N_6804,N_5080,N_5064);
and U6805 (N_6805,N_5794,N_5445);
nand U6806 (N_6806,N_5963,N_5071);
nor U6807 (N_6807,N_5551,N_5756);
nand U6808 (N_6808,N_5935,N_5583);
xor U6809 (N_6809,N_5317,N_5522);
or U6810 (N_6810,N_5436,N_5247);
nand U6811 (N_6811,N_5296,N_5749);
and U6812 (N_6812,N_5003,N_5712);
nand U6813 (N_6813,N_5217,N_5350);
nor U6814 (N_6814,N_5700,N_5636);
nand U6815 (N_6815,N_5106,N_5927);
or U6816 (N_6816,N_5935,N_5362);
or U6817 (N_6817,N_5764,N_5336);
nor U6818 (N_6818,N_5146,N_5007);
nor U6819 (N_6819,N_5595,N_5960);
or U6820 (N_6820,N_5019,N_5562);
and U6821 (N_6821,N_5169,N_5256);
nand U6822 (N_6822,N_5510,N_5358);
nor U6823 (N_6823,N_5684,N_5841);
nand U6824 (N_6824,N_5701,N_5008);
or U6825 (N_6825,N_5568,N_5311);
or U6826 (N_6826,N_5965,N_5817);
nand U6827 (N_6827,N_5012,N_5528);
and U6828 (N_6828,N_5219,N_5274);
nor U6829 (N_6829,N_5697,N_5147);
or U6830 (N_6830,N_5856,N_5696);
or U6831 (N_6831,N_5469,N_5560);
xor U6832 (N_6832,N_5664,N_5228);
nor U6833 (N_6833,N_5992,N_5083);
or U6834 (N_6834,N_5871,N_5931);
nor U6835 (N_6835,N_5750,N_5237);
xnor U6836 (N_6836,N_5989,N_5898);
or U6837 (N_6837,N_5037,N_5632);
nor U6838 (N_6838,N_5603,N_5058);
nor U6839 (N_6839,N_5365,N_5963);
nor U6840 (N_6840,N_5354,N_5914);
nor U6841 (N_6841,N_5770,N_5870);
and U6842 (N_6842,N_5057,N_5854);
and U6843 (N_6843,N_5849,N_5475);
or U6844 (N_6844,N_5719,N_5048);
nor U6845 (N_6845,N_5109,N_5898);
xnor U6846 (N_6846,N_5864,N_5209);
nand U6847 (N_6847,N_5592,N_5267);
nor U6848 (N_6848,N_5213,N_5559);
xnor U6849 (N_6849,N_5753,N_5300);
xor U6850 (N_6850,N_5380,N_5979);
nand U6851 (N_6851,N_5991,N_5106);
or U6852 (N_6852,N_5301,N_5737);
nand U6853 (N_6853,N_5926,N_5311);
nand U6854 (N_6854,N_5153,N_5416);
nand U6855 (N_6855,N_5667,N_5364);
nand U6856 (N_6856,N_5776,N_5911);
xnor U6857 (N_6857,N_5363,N_5275);
nand U6858 (N_6858,N_5723,N_5293);
nor U6859 (N_6859,N_5724,N_5059);
nand U6860 (N_6860,N_5057,N_5285);
or U6861 (N_6861,N_5994,N_5368);
nand U6862 (N_6862,N_5501,N_5835);
nor U6863 (N_6863,N_5182,N_5034);
or U6864 (N_6864,N_5289,N_5203);
xnor U6865 (N_6865,N_5759,N_5893);
nand U6866 (N_6866,N_5153,N_5398);
nor U6867 (N_6867,N_5128,N_5076);
nor U6868 (N_6868,N_5826,N_5445);
nand U6869 (N_6869,N_5295,N_5632);
or U6870 (N_6870,N_5196,N_5801);
xor U6871 (N_6871,N_5713,N_5638);
nand U6872 (N_6872,N_5421,N_5257);
nor U6873 (N_6873,N_5068,N_5585);
and U6874 (N_6874,N_5962,N_5790);
nor U6875 (N_6875,N_5154,N_5141);
and U6876 (N_6876,N_5155,N_5404);
nand U6877 (N_6877,N_5235,N_5434);
xnor U6878 (N_6878,N_5943,N_5486);
and U6879 (N_6879,N_5895,N_5059);
nand U6880 (N_6880,N_5494,N_5007);
xnor U6881 (N_6881,N_5314,N_5970);
nand U6882 (N_6882,N_5564,N_5351);
nand U6883 (N_6883,N_5138,N_5207);
or U6884 (N_6884,N_5945,N_5828);
or U6885 (N_6885,N_5341,N_5029);
and U6886 (N_6886,N_5731,N_5742);
nor U6887 (N_6887,N_5155,N_5421);
xnor U6888 (N_6888,N_5632,N_5140);
nand U6889 (N_6889,N_5347,N_5445);
or U6890 (N_6890,N_5812,N_5147);
and U6891 (N_6891,N_5818,N_5726);
xnor U6892 (N_6892,N_5191,N_5202);
and U6893 (N_6893,N_5943,N_5413);
or U6894 (N_6894,N_5251,N_5647);
and U6895 (N_6895,N_5958,N_5925);
nor U6896 (N_6896,N_5933,N_5722);
or U6897 (N_6897,N_5909,N_5739);
nand U6898 (N_6898,N_5613,N_5434);
or U6899 (N_6899,N_5134,N_5880);
nor U6900 (N_6900,N_5890,N_5778);
nand U6901 (N_6901,N_5106,N_5599);
nand U6902 (N_6902,N_5761,N_5677);
xor U6903 (N_6903,N_5187,N_5922);
xor U6904 (N_6904,N_5037,N_5309);
and U6905 (N_6905,N_5387,N_5992);
nand U6906 (N_6906,N_5286,N_5355);
nand U6907 (N_6907,N_5843,N_5599);
xnor U6908 (N_6908,N_5045,N_5479);
and U6909 (N_6909,N_5359,N_5858);
xor U6910 (N_6910,N_5540,N_5533);
or U6911 (N_6911,N_5202,N_5189);
xor U6912 (N_6912,N_5799,N_5702);
or U6913 (N_6913,N_5638,N_5284);
or U6914 (N_6914,N_5112,N_5497);
nor U6915 (N_6915,N_5723,N_5825);
nor U6916 (N_6916,N_5933,N_5112);
and U6917 (N_6917,N_5923,N_5741);
or U6918 (N_6918,N_5503,N_5079);
or U6919 (N_6919,N_5762,N_5032);
nor U6920 (N_6920,N_5446,N_5626);
or U6921 (N_6921,N_5256,N_5527);
xnor U6922 (N_6922,N_5516,N_5718);
and U6923 (N_6923,N_5535,N_5588);
and U6924 (N_6924,N_5147,N_5359);
and U6925 (N_6925,N_5904,N_5278);
nor U6926 (N_6926,N_5759,N_5874);
xnor U6927 (N_6927,N_5682,N_5157);
or U6928 (N_6928,N_5534,N_5014);
and U6929 (N_6929,N_5600,N_5125);
nor U6930 (N_6930,N_5082,N_5600);
xor U6931 (N_6931,N_5303,N_5273);
nor U6932 (N_6932,N_5027,N_5596);
or U6933 (N_6933,N_5333,N_5390);
nand U6934 (N_6934,N_5595,N_5497);
and U6935 (N_6935,N_5996,N_5002);
and U6936 (N_6936,N_5336,N_5375);
or U6937 (N_6937,N_5293,N_5295);
and U6938 (N_6938,N_5526,N_5477);
or U6939 (N_6939,N_5060,N_5681);
xor U6940 (N_6940,N_5370,N_5018);
xnor U6941 (N_6941,N_5766,N_5683);
nor U6942 (N_6942,N_5851,N_5700);
xnor U6943 (N_6943,N_5319,N_5027);
nor U6944 (N_6944,N_5521,N_5808);
and U6945 (N_6945,N_5541,N_5056);
or U6946 (N_6946,N_5521,N_5876);
nand U6947 (N_6947,N_5595,N_5967);
nor U6948 (N_6948,N_5792,N_5805);
and U6949 (N_6949,N_5163,N_5624);
nand U6950 (N_6950,N_5580,N_5624);
or U6951 (N_6951,N_5974,N_5497);
and U6952 (N_6952,N_5622,N_5395);
and U6953 (N_6953,N_5954,N_5188);
or U6954 (N_6954,N_5823,N_5484);
nor U6955 (N_6955,N_5998,N_5213);
xnor U6956 (N_6956,N_5749,N_5432);
xnor U6957 (N_6957,N_5141,N_5639);
xor U6958 (N_6958,N_5233,N_5514);
nor U6959 (N_6959,N_5195,N_5439);
or U6960 (N_6960,N_5023,N_5574);
xor U6961 (N_6961,N_5491,N_5718);
or U6962 (N_6962,N_5745,N_5249);
nand U6963 (N_6963,N_5922,N_5420);
nand U6964 (N_6964,N_5449,N_5843);
xor U6965 (N_6965,N_5783,N_5322);
or U6966 (N_6966,N_5172,N_5792);
nor U6967 (N_6967,N_5500,N_5149);
nor U6968 (N_6968,N_5673,N_5921);
nor U6969 (N_6969,N_5174,N_5032);
xor U6970 (N_6970,N_5790,N_5699);
or U6971 (N_6971,N_5978,N_5324);
and U6972 (N_6972,N_5319,N_5029);
nand U6973 (N_6973,N_5322,N_5990);
and U6974 (N_6974,N_5212,N_5827);
xnor U6975 (N_6975,N_5119,N_5410);
nand U6976 (N_6976,N_5042,N_5205);
and U6977 (N_6977,N_5009,N_5252);
nand U6978 (N_6978,N_5201,N_5651);
or U6979 (N_6979,N_5634,N_5266);
and U6980 (N_6980,N_5225,N_5178);
or U6981 (N_6981,N_5926,N_5855);
and U6982 (N_6982,N_5368,N_5426);
nor U6983 (N_6983,N_5643,N_5135);
or U6984 (N_6984,N_5479,N_5993);
nor U6985 (N_6985,N_5824,N_5905);
nor U6986 (N_6986,N_5866,N_5378);
and U6987 (N_6987,N_5062,N_5752);
or U6988 (N_6988,N_5841,N_5068);
or U6989 (N_6989,N_5366,N_5459);
nor U6990 (N_6990,N_5905,N_5788);
nand U6991 (N_6991,N_5142,N_5055);
or U6992 (N_6992,N_5285,N_5389);
nand U6993 (N_6993,N_5230,N_5488);
xnor U6994 (N_6994,N_5161,N_5237);
or U6995 (N_6995,N_5222,N_5428);
nand U6996 (N_6996,N_5930,N_5758);
or U6997 (N_6997,N_5008,N_5891);
or U6998 (N_6998,N_5411,N_5298);
nor U6999 (N_6999,N_5727,N_5078);
and U7000 (N_7000,N_6295,N_6313);
nor U7001 (N_7001,N_6112,N_6994);
nand U7002 (N_7002,N_6944,N_6069);
xnor U7003 (N_7003,N_6446,N_6523);
nand U7004 (N_7004,N_6336,N_6596);
or U7005 (N_7005,N_6632,N_6009);
xor U7006 (N_7006,N_6582,N_6160);
xnor U7007 (N_7007,N_6146,N_6440);
and U7008 (N_7008,N_6049,N_6846);
nand U7009 (N_7009,N_6294,N_6766);
or U7010 (N_7010,N_6122,N_6171);
nor U7011 (N_7011,N_6188,N_6547);
and U7012 (N_7012,N_6000,N_6803);
xnor U7013 (N_7013,N_6284,N_6301);
and U7014 (N_7014,N_6155,N_6512);
nand U7015 (N_7015,N_6731,N_6159);
and U7016 (N_7016,N_6973,N_6256);
and U7017 (N_7017,N_6214,N_6922);
nor U7018 (N_7018,N_6535,N_6511);
or U7019 (N_7019,N_6283,N_6402);
nor U7020 (N_7020,N_6267,N_6299);
nor U7021 (N_7021,N_6437,N_6269);
nor U7022 (N_7022,N_6891,N_6292);
nand U7023 (N_7023,N_6379,N_6829);
nand U7024 (N_7024,N_6491,N_6821);
or U7025 (N_7025,N_6908,N_6770);
or U7026 (N_7026,N_6241,N_6854);
nor U7027 (N_7027,N_6985,N_6033);
xnor U7028 (N_7028,N_6149,N_6881);
nand U7029 (N_7029,N_6273,N_6842);
xor U7030 (N_7030,N_6137,N_6763);
nand U7031 (N_7031,N_6430,N_6442);
nand U7032 (N_7032,N_6579,N_6817);
nand U7033 (N_7033,N_6485,N_6525);
nor U7034 (N_7034,N_6066,N_6427);
and U7035 (N_7035,N_6056,N_6712);
xor U7036 (N_7036,N_6342,N_6786);
xnor U7037 (N_7037,N_6691,N_6627);
or U7038 (N_7038,N_6896,N_6978);
and U7039 (N_7039,N_6309,N_6096);
xor U7040 (N_7040,N_6239,N_6259);
nand U7041 (N_7041,N_6539,N_6948);
nor U7042 (N_7042,N_6135,N_6420);
nand U7043 (N_7043,N_6394,N_6813);
nor U7044 (N_7044,N_6277,N_6290);
xor U7045 (N_7045,N_6411,N_6010);
and U7046 (N_7046,N_6199,N_6477);
or U7047 (N_7047,N_6240,N_6963);
and U7048 (N_7048,N_6074,N_6636);
and U7049 (N_7049,N_6676,N_6460);
and U7050 (N_7050,N_6100,N_6822);
nor U7051 (N_7051,N_6193,N_6794);
or U7052 (N_7052,N_6017,N_6625);
nor U7053 (N_7053,N_6031,N_6417);
nand U7054 (N_7054,N_6787,N_6459);
nand U7055 (N_7055,N_6654,N_6971);
nand U7056 (N_7056,N_6436,N_6153);
xnor U7057 (N_7057,N_6716,N_6921);
or U7058 (N_7058,N_6097,N_6736);
xnor U7059 (N_7059,N_6601,N_6263);
and U7060 (N_7060,N_6289,N_6138);
or U7061 (N_7061,N_6217,N_6139);
nand U7062 (N_7062,N_6197,N_6665);
nand U7063 (N_7063,N_6573,N_6004);
nand U7064 (N_7064,N_6529,N_6707);
xor U7065 (N_7065,N_6488,N_6245);
and U7066 (N_7066,N_6564,N_6690);
nand U7067 (N_7067,N_6509,N_6725);
and U7068 (N_7068,N_6989,N_6492);
xor U7069 (N_7069,N_6917,N_6605);
or U7070 (N_7070,N_6611,N_6330);
and U7071 (N_7071,N_6649,N_6723);
and U7072 (N_7072,N_6385,N_6623);
xnor U7073 (N_7073,N_6494,N_6077);
nor U7074 (N_7074,N_6435,N_6785);
nand U7075 (N_7075,N_6775,N_6237);
nor U7076 (N_7076,N_6520,N_6085);
or U7077 (N_7077,N_6316,N_6132);
nor U7078 (N_7078,N_6063,N_6484);
or U7079 (N_7079,N_6373,N_6161);
and U7080 (N_7080,N_6319,N_6646);
xor U7081 (N_7081,N_6013,N_6044);
xor U7082 (N_7082,N_6081,N_6694);
xor U7083 (N_7083,N_6659,N_6195);
xor U7084 (N_7084,N_6234,N_6769);
nor U7085 (N_7085,N_6489,N_6597);
nand U7086 (N_7086,N_6550,N_6473);
xor U7087 (N_7087,N_6230,N_6183);
nand U7088 (N_7088,N_6305,N_6522);
nor U7089 (N_7089,N_6997,N_6203);
or U7090 (N_7090,N_6895,N_6006);
xor U7091 (N_7091,N_6588,N_6567);
and U7092 (N_7092,N_6622,N_6128);
xnor U7093 (N_7093,N_6873,N_6101);
nand U7094 (N_7094,N_6984,N_6875);
xnor U7095 (N_7095,N_6657,N_6118);
or U7096 (N_7096,N_6426,N_6415);
xnor U7097 (N_7097,N_6923,N_6496);
nand U7098 (N_7098,N_6508,N_6023);
or U7099 (N_7099,N_6324,N_6951);
nand U7100 (N_7100,N_6840,N_6943);
and U7101 (N_7101,N_6253,N_6860);
and U7102 (N_7102,N_6483,N_6897);
xnor U7103 (N_7103,N_6104,N_6030);
or U7104 (N_7104,N_6879,N_6278);
or U7105 (N_7105,N_6580,N_6397);
or U7106 (N_7106,N_6924,N_6920);
nor U7107 (N_7107,N_6872,N_6852);
and U7108 (N_7108,N_6062,N_6046);
and U7109 (N_7109,N_6124,N_6647);
xor U7110 (N_7110,N_6850,N_6094);
nor U7111 (N_7111,N_6679,N_6447);
xor U7112 (N_7112,N_6747,N_6981);
nor U7113 (N_7113,N_6003,N_6047);
xor U7114 (N_7114,N_6403,N_6025);
xor U7115 (N_7115,N_6705,N_6334);
and U7116 (N_7116,N_6793,N_6629);
xnor U7117 (N_7117,N_6753,N_6838);
xnor U7118 (N_7118,N_6482,N_6699);
xnor U7119 (N_7119,N_6113,N_6857);
nor U7120 (N_7120,N_6453,N_6162);
nand U7121 (N_7121,N_6792,N_6359);
nor U7122 (N_7122,N_6142,N_6586);
xnor U7123 (N_7123,N_6158,N_6350);
xor U7124 (N_7124,N_6804,N_6515);
nor U7125 (N_7125,N_6396,N_6519);
or U7126 (N_7126,N_6714,N_6980);
xnor U7127 (N_7127,N_6765,N_6903);
or U7128 (N_7128,N_6381,N_6734);
nand U7129 (N_7129,N_6789,N_6377);
or U7130 (N_7130,N_6530,N_6667);
and U7131 (N_7131,N_6185,N_6098);
and U7132 (N_7132,N_6560,N_6035);
nor U7133 (N_7133,N_6554,N_6826);
nor U7134 (N_7134,N_6858,N_6021);
or U7135 (N_7135,N_6628,N_6036);
nor U7136 (N_7136,N_6678,N_6120);
xnor U7137 (N_7137,N_6938,N_6772);
or U7138 (N_7138,N_6189,N_6900);
nand U7139 (N_7139,N_6907,N_6246);
or U7140 (N_7140,N_6758,N_6005);
xnor U7141 (N_7141,N_6020,N_6653);
and U7142 (N_7142,N_6929,N_6585);
nand U7143 (N_7143,N_6507,N_6320);
or U7144 (N_7144,N_6754,N_6387);
xnor U7145 (N_7145,N_6422,N_6904);
nor U7146 (N_7146,N_6784,N_6285);
xnor U7147 (N_7147,N_6696,N_6177);
nand U7148 (N_7148,N_6052,N_6574);
xor U7149 (N_7149,N_6556,N_6869);
xor U7150 (N_7150,N_6429,N_6503);
nand U7151 (N_7151,N_6527,N_6602);
and U7152 (N_7152,N_6048,N_6455);
nand U7153 (N_7153,N_6079,N_6007);
or U7154 (N_7154,N_6669,N_6034);
nand U7155 (N_7155,N_6764,N_6448);
nand U7156 (N_7156,N_6834,N_6167);
nand U7157 (N_7157,N_6932,N_6075);
nand U7158 (N_7158,N_6478,N_6972);
or U7159 (N_7159,N_6011,N_6966);
xor U7160 (N_7160,N_6143,N_6552);
and U7161 (N_7161,N_6053,N_6721);
xor U7162 (N_7162,N_6480,N_6412);
and U7163 (N_7163,N_6687,N_6641);
xor U7164 (N_7164,N_6252,N_6670);
and U7165 (N_7165,N_6180,N_6768);
nor U7166 (N_7166,N_6068,N_6406);
nand U7167 (N_7167,N_6986,N_6959);
or U7168 (N_7168,N_6992,N_6909);
and U7169 (N_7169,N_6534,N_6443);
nand U7170 (N_7170,N_6391,N_6370);
nand U7171 (N_7171,N_6867,N_6376);
nand U7172 (N_7172,N_6014,N_6713);
and U7173 (N_7173,N_6710,N_6968);
nand U7174 (N_7174,N_6839,N_6783);
nand U7175 (N_7175,N_6619,N_6414);
nor U7176 (N_7176,N_6626,N_6178);
xor U7177 (N_7177,N_6365,N_6836);
nand U7178 (N_7178,N_6913,N_6543);
nor U7179 (N_7179,N_6516,N_6592);
or U7180 (N_7180,N_6463,N_6991);
nand U7181 (N_7181,N_6756,N_6998);
nand U7182 (N_7182,N_6828,N_6206);
or U7183 (N_7183,N_6018,N_6421);
nand U7184 (N_7184,N_6045,N_6987);
xor U7185 (N_7185,N_6321,N_6739);
xor U7186 (N_7186,N_6136,N_6732);
or U7187 (N_7187,N_6400,N_6250);
xnor U7188 (N_7188,N_6419,N_6911);
xor U7189 (N_7189,N_6957,N_6235);
and U7190 (N_7190,N_6399,N_6255);
or U7191 (N_7191,N_6759,N_6486);
nor U7192 (N_7192,N_6367,N_6902);
nor U7193 (N_7193,N_6498,N_6983);
xnor U7194 (N_7194,N_6060,N_6565);
xor U7195 (N_7195,N_6578,N_6233);
and U7196 (N_7196,N_6102,N_6608);
nor U7197 (N_7197,N_6272,N_6302);
xnor U7198 (N_7198,N_6815,N_6607);
and U7199 (N_7199,N_6868,N_6589);
nand U7200 (N_7200,N_6466,N_6563);
and U7201 (N_7201,N_6729,N_6244);
xor U7202 (N_7202,N_6660,N_6280);
nor U7203 (N_7203,N_6479,N_6261);
xnor U7204 (N_7204,N_6490,N_6746);
or U7205 (N_7205,N_6859,N_6349);
and U7206 (N_7206,N_6374,N_6054);
xor U7207 (N_7207,N_6404,N_6595);
nor U7208 (N_7208,N_6974,N_6371);
nor U7209 (N_7209,N_6121,N_6856);
or U7210 (N_7210,N_6548,N_6791);
xnor U7211 (N_7211,N_6688,N_6117);
nand U7212 (N_7212,N_6166,N_6340);
and U7213 (N_7213,N_6941,N_6057);
nor U7214 (N_7214,N_6827,N_6092);
xor U7215 (N_7215,N_6843,N_6639);
xnor U7216 (N_7216,N_6767,N_6878);
or U7217 (N_7217,N_6439,N_6172);
nor U7218 (N_7218,N_6999,N_6979);
or U7219 (N_7219,N_6493,N_6502);
nand U7220 (N_7220,N_6845,N_6583);
xor U7221 (N_7221,N_6975,N_6735);
nand U7222 (N_7222,N_6949,N_6886);
and U7223 (N_7223,N_6888,N_6300);
nand U7224 (N_7224,N_6610,N_6876);
or U7225 (N_7225,N_6219,N_6617);
xor U7226 (N_7226,N_6618,N_6742);
nor U7227 (N_7227,N_6820,N_6380);
or U7228 (N_7228,N_6545,N_6078);
and U7229 (N_7229,N_6952,N_6147);
xnor U7230 (N_7230,N_6884,N_6083);
and U7231 (N_7231,N_6870,N_6717);
or U7232 (N_7232,N_6029,N_6022);
nand U7233 (N_7233,N_6606,N_6914);
or U7234 (N_7234,N_6107,N_6964);
xnor U7235 (N_7235,N_6110,N_6111);
and U7236 (N_7236,N_6635,N_6012);
xor U7237 (N_7237,N_6559,N_6231);
xor U7238 (N_7238,N_6940,N_6835);
nand U7239 (N_7239,N_6740,N_6788);
and U7240 (N_7240,N_6645,N_6528);
nand U7241 (N_7241,N_6631,N_6418);
nand U7242 (N_7242,N_6312,N_6621);
and U7243 (N_7243,N_6894,N_6348);
and U7244 (N_7244,N_6222,N_6663);
xnor U7245 (N_7245,N_6366,N_6157);
nor U7246 (N_7246,N_6750,N_6115);
or U7247 (N_7247,N_6861,N_6282);
and U7248 (N_7248,N_6598,N_6039);
and U7249 (N_7249,N_6616,N_6795);
xor U7250 (N_7250,N_6613,N_6774);
nand U7251 (N_7251,N_6229,N_6849);
xor U7252 (N_7252,N_6880,N_6258);
or U7253 (N_7253,N_6848,N_6844);
xnor U7254 (N_7254,N_6883,N_6458);
xnor U7255 (N_7255,N_6433,N_6898);
and U7256 (N_7256,N_6428,N_6262);
and U7257 (N_7257,N_6958,N_6542);
and U7258 (N_7258,N_6333,N_6939);
nand U7259 (N_7259,N_6425,N_6378);
and U7260 (N_7260,N_6182,N_6450);
xor U7261 (N_7261,N_6257,N_6454);
nor U7262 (N_7262,N_6072,N_6771);
nor U7263 (N_7263,N_6877,N_6893);
or U7264 (N_7264,N_6401,N_6393);
nand U7265 (N_7265,N_6549,N_6593);
xor U7266 (N_7266,N_6851,N_6733);
nor U7267 (N_7267,N_6469,N_6906);
or U7268 (N_7268,N_6487,N_6633);
nor U7269 (N_7269,N_6109,N_6467);
xor U7270 (N_7270,N_6328,N_6051);
and U7271 (N_7271,N_6743,N_6925);
or U7272 (N_7272,N_6500,N_6087);
nand U7273 (N_7273,N_6561,N_6651);
nor U7274 (N_7274,N_6457,N_6223);
nor U7275 (N_7275,N_6431,N_6002);
or U7276 (N_7276,N_6346,N_6232);
nand U7277 (N_7277,N_6581,N_6163);
nand U7278 (N_7278,N_6040,N_6615);
or U7279 (N_7279,N_6495,N_6499);
xnor U7280 (N_7280,N_6709,N_6553);
or U7281 (N_7281,N_6584,N_6778);
nand U7282 (N_7282,N_6684,N_6095);
xnor U7283 (N_7283,N_6557,N_6027);
xnor U7284 (N_7284,N_6726,N_6315);
nor U7285 (N_7285,N_6945,N_6953);
and U7286 (N_7286,N_6700,N_6314);
nor U7287 (N_7287,N_6644,N_6600);
and U7288 (N_7288,N_6781,N_6474);
nor U7289 (N_7289,N_6354,N_6541);
or U7290 (N_7290,N_6666,N_6703);
xnor U7291 (N_7291,N_6970,N_6782);
xnor U7292 (N_7292,N_6064,N_6291);
nand U7293 (N_7293,N_6026,N_6363);
xor U7294 (N_7294,N_6720,N_6745);
or U7295 (N_7295,N_6501,N_6326);
nand U7296 (N_7296,N_6140,N_6073);
xnor U7297 (N_7297,N_6192,N_6755);
nand U7298 (N_7298,N_6928,N_6360);
nand U7299 (N_7299,N_6200,N_6650);
and U7300 (N_7300,N_6995,N_6386);
and U7301 (N_7301,N_6930,N_6042);
nand U7302 (N_7302,N_6347,N_6701);
or U7303 (N_7303,N_6942,N_6505);
nand U7304 (N_7304,N_6179,N_6853);
and U7305 (N_7305,N_6802,N_6086);
nor U7306 (N_7306,N_6213,N_6668);
nand U7307 (N_7307,N_6369,N_6801);
nand U7308 (N_7308,N_6198,N_6796);
nor U7309 (N_7309,N_6572,N_6551);
nand U7310 (N_7310,N_6620,N_6962);
nor U7311 (N_7311,N_6212,N_6812);
nor U7312 (N_7312,N_6531,N_6915);
and U7313 (N_7313,N_6260,N_6916);
nor U7314 (N_7314,N_6969,N_6016);
or U7315 (N_7315,N_6090,N_6693);
or U7316 (N_7316,N_6043,N_6797);
or U7317 (N_7317,N_6341,N_6905);
or U7318 (N_7318,N_6640,N_6566);
nor U7319 (N_7319,N_6224,N_6536);
xnor U7320 (N_7320,N_6744,N_6780);
xnor U7321 (N_7321,N_6936,N_6228);
and U7322 (N_7322,N_6874,N_6708);
nor U7323 (N_7323,N_6424,N_6175);
xnor U7324 (N_7324,N_6254,N_6151);
nor U7325 (N_7325,N_6332,N_6187);
xnor U7326 (N_7326,N_6306,N_6226);
or U7327 (N_7327,N_6497,N_6238);
nor U7328 (N_7328,N_6704,N_6298);
nand U7329 (N_7329,N_6960,N_6819);
or U7330 (N_7330,N_6521,N_6337);
and U7331 (N_7331,N_6242,N_6407);
nand U7332 (N_7332,N_6555,N_6624);
or U7333 (N_7333,N_6355,N_6977);
xnor U7334 (N_7334,N_6630,N_6329);
nor U7335 (N_7335,N_6697,N_6304);
nor U7336 (N_7336,N_6470,N_6270);
nor U7337 (N_7337,N_6777,N_6871);
or U7338 (N_7338,N_6130,N_6032);
nand U7339 (N_7339,N_6818,N_6382);
or U7340 (N_7340,N_6674,N_6296);
nor U7341 (N_7341,N_6410,N_6976);
and U7342 (N_7342,N_6445,N_6331);
and U7343 (N_7343,N_6275,N_6384);
nor U7344 (N_7344,N_6954,N_6558);
or U7345 (N_7345,N_6288,N_6220);
nand U7346 (N_7346,N_6706,N_6760);
and U7347 (N_7347,N_6946,N_6824);
nor U7348 (N_7348,N_6024,N_6207);
and U7349 (N_7349,N_6912,N_6800);
xor U7350 (N_7350,N_6015,N_6395);
and U7351 (N_7351,N_6279,N_6372);
nor U7352 (N_7352,N_6236,N_6510);
xor U7353 (N_7353,N_6388,N_6173);
xor U7354 (N_7354,N_6779,N_6215);
xnor U7355 (N_7355,N_6456,N_6808);
nand U7356 (N_7356,N_6191,N_6170);
or U7357 (N_7357,N_6672,N_6310);
nand U7358 (N_7358,N_6658,N_6449);
nor U7359 (N_7359,N_6937,N_6737);
nor U7360 (N_7360,N_6125,N_6037);
and U7361 (N_7361,N_6680,N_6356);
or U7362 (N_7362,N_6686,N_6965);
nand U7363 (N_7363,N_6947,N_6677);
xor U7364 (N_7364,N_6345,N_6416);
and U7365 (N_7365,N_6671,N_6001);
xor U7366 (N_7366,N_6196,N_6210);
nand U7367 (N_7367,N_6741,N_6145);
and U7368 (N_7368,N_6209,N_6591);
nor U7369 (N_7369,N_6790,N_6517);
nor U7370 (N_7370,N_6899,N_6481);
nand U7371 (N_7371,N_6643,N_6599);
or U7372 (N_7372,N_6216,N_6218);
xnor U7373 (N_7373,N_6807,N_6637);
xnor U7374 (N_7374,N_6357,N_6882);
nand U7375 (N_7375,N_6506,N_6127);
and U7376 (N_7376,N_6368,N_6243);
nand U7377 (N_7377,N_6988,N_6833);
nand U7378 (N_7378,N_6587,N_6855);
xnor U7379 (N_7379,N_6082,N_6451);
or U7380 (N_7380,N_6810,N_6084);
or U7381 (N_7381,N_6123,N_6168);
nor U7382 (N_7382,N_6061,N_6204);
or U7383 (N_7383,N_6661,N_6863);
xnor U7384 (N_7384,N_6106,N_6748);
nor U7385 (N_7385,N_6773,N_6413);
nor U7386 (N_7386,N_6268,N_6533);
and U7387 (N_7387,N_6752,N_6089);
and U7388 (N_7388,N_6405,N_6830);
and U7389 (N_7389,N_6832,N_6652);
xor U7390 (N_7390,N_6464,N_6814);
nand U7391 (N_7391,N_6603,N_6303);
or U7392 (N_7392,N_6919,N_6514);
nand U7393 (N_7393,N_6642,N_6311);
xnor U7394 (N_7394,N_6325,N_6664);
and U7395 (N_7395,N_6156,N_6809);
and U7396 (N_7396,N_6577,N_6546);
or U7397 (N_7397,N_6108,N_6675);
nand U7398 (N_7398,N_6080,N_6264);
and U7399 (N_7399,N_6926,N_6961);
and U7400 (N_7400,N_6339,N_6776);
xnor U7401 (N_7401,N_6841,N_6059);
nand U7402 (N_7402,N_6638,N_6996);
xnor U7403 (N_7403,N_6569,N_6141);
and U7404 (N_7404,N_6266,N_6575);
nor U7405 (N_7405,N_6343,N_6805);
xor U7406 (N_7406,N_6685,N_6297);
xor U7407 (N_7407,N_6901,N_6811);
and U7408 (N_7408,N_6544,N_6576);
xor U7409 (N_7409,N_6662,N_6184);
or U7410 (N_7410,N_6186,N_6590);
and U7411 (N_7411,N_6967,N_6148);
or U7412 (N_7412,N_6462,N_6344);
xnor U7413 (N_7413,N_6798,N_6648);
nand U7414 (N_7414,N_6119,N_6181);
nand U7415 (N_7415,N_6950,N_6008);
xnor U7416 (N_7416,N_6208,N_6927);
xor U7417 (N_7417,N_6890,N_6317);
or U7418 (N_7418,N_6067,N_6562);
and U7419 (N_7419,N_6114,N_6065);
and U7420 (N_7420,N_6276,N_6169);
nand U7421 (N_7421,N_6571,N_6823);
xor U7422 (N_7422,N_6211,N_6472);
and U7423 (N_7423,N_6715,N_6041);
xnor U7424 (N_7424,N_6831,N_6935);
nand U7425 (N_7425,N_6934,N_6538);
xnor U7426 (N_7426,N_6205,N_6799);
and U7427 (N_7427,N_6614,N_6308);
nor U7428 (N_7428,N_6126,N_6982);
or U7429 (N_7429,N_6892,N_6461);
nand U7430 (N_7430,N_6910,N_6055);
xnor U7431 (N_7431,N_6202,N_6749);
xor U7432 (N_7432,N_6116,N_6362);
nor U7433 (N_7433,N_6375,N_6174);
nor U7434 (N_7434,N_6129,N_6471);
and U7435 (N_7435,N_6133,N_6718);
nor U7436 (N_7436,N_6438,N_6570);
nor U7437 (N_7437,N_6933,N_6757);
and U7438 (N_7438,N_6383,N_6164);
nand U7439 (N_7439,N_6221,N_6955);
or U7440 (N_7440,N_6656,N_6327);
xnor U7441 (N_7441,N_6287,N_6609);
or U7442 (N_7442,N_6398,N_6751);
xnor U7443 (N_7443,N_6103,N_6389);
and U7444 (N_7444,N_6468,N_6692);
xor U7445 (N_7445,N_6190,N_6227);
or U7446 (N_7446,N_6058,N_6475);
and U7447 (N_7447,N_6201,N_6423);
nand U7448 (N_7448,N_6816,N_6038);
xor U7449 (N_7449,N_6719,N_6150);
or U7450 (N_7450,N_6131,N_6351);
and U7451 (N_7451,N_6722,N_6866);
nor U7452 (N_7452,N_6322,N_6634);
nand U7453 (N_7453,N_6409,N_6837);
nand U7454 (N_7454,N_6318,N_6465);
nor U7455 (N_7455,N_6825,N_6353);
nand U7456 (N_7456,N_6071,N_6165);
xnor U7457 (N_7457,N_6526,N_6728);
xnor U7458 (N_7458,N_6918,N_6931);
nand U7459 (N_7459,N_6682,N_6673);
nand U7460 (N_7460,N_6099,N_6956);
and U7461 (N_7461,N_6612,N_6540);
or U7462 (N_7462,N_6513,N_6738);
and U7463 (N_7463,N_6247,N_6154);
nand U7464 (N_7464,N_6885,N_6028);
nor U7465 (N_7465,N_6286,N_6249);
xor U7466 (N_7466,N_6352,N_6864);
nor U7467 (N_7467,N_6070,N_6358);
nor U7468 (N_7468,N_6093,N_6091);
nor U7469 (N_7469,N_6361,N_6307);
or U7470 (N_7470,N_6727,N_6144);
nand U7471 (N_7471,N_6476,N_6293);
xnor U7472 (N_7472,N_6225,N_6762);
nand U7473 (N_7473,N_6338,N_6702);
nor U7474 (N_7474,N_6452,N_6444);
and U7475 (N_7475,N_6862,N_6271);
and U7476 (N_7476,N_6281,N_6134);
nand U7477 (N_7477,N_6604,N_6990);
xnor U7478 (N_7478,N_6847,N_6176);
and U7479 (N_7479,N_6537,N_6806);
and U7480 (N_7480,N_6323,N_6019);
xnor U7481 (N_7481,N_6655,N_6152);
or U7482 (N_7482,N_6698,N_6724);
xor U7483 (N_7483,N_6689,N_6248);
or U7484 (N_7484,N_6050,N_6434);
xnor U7485 (N_7485,N_6887,N_6695);
xnor U7486 (N_7486,N_6594,N_6194);
nand U7487 (N_7487,N_6432,N_6251);
and U7488 (N_7488,N_6335,N_6568);
or U7489 (N_7489,N_6088,N_6265);
xor U7490 (N_7490,N_6711,N_6524);
xor U7491 (N_7491,N_6504,N_6681);
xor U7492 (N_7492,N_6274,N_6865);
nor U7493 (N_7493,N_6364,N_6532);
or U7494 (N_7494,N_6518,N_6076);
xnor U7495 (N_7495,N_6105,N_6408);
xor U7496 (N_7496,N_6993,N_6441);
nand U7497 (N_7497,N_6889,N_6392);
and U7498 (N_7498,N_6730,N_6390);
or U7499 (N_7499,N_6683,N_6761);
or U7500 (N_7500,N_6645,N_6297);
and U7501 (N_7501,N_6424,N_6372);
or U7502 (N_7502,N_6696,N_6237);
and U7503 (N_7503,N_6372,N_6878);
nand U7504 (N_7504,N_6077,N_6788);
nor U7505 (N_7505,N_6804,N_6541);
or U7506 (N_7506,N_6922,N_6438);
xnor U7507 (N_7507,N_6288,N_6976);
or U7508 (N_7508,N_6319,N_6804);
nand U7509 (N_7509,N_6065,N_6044);
and U7510 (N_7510,N_6530,N_6637);
or U7511 (N_7511,N_6063,N_6756);
nor U7512 (N_7512,N_6861,N_6686);
nor U7513 (N_7513,N_6428,N_6324);
or U7514 (N_7514,N_6577,N_6102);
nand U7515 (N_7515,N_6625,N_6815);
or U7516 (N_7516,N_6049,N_6080);
nand U7517 (N_7517,N_6577,N_6336);
or U7518 (N_7518,N_6072,N_6462);
or U7519 (N_7519,N_6236,N_6886);
nor U7520 (N_7520,N_6457,N_6357);
nand U7521 (N_7521,N_6520,N_6594);
and U7522 (N_7522,N_6711,N_6255);
xnor U7523 (N_7523,N_6504,N_6026);
nor U7524 (N_7524,N_6304,N_6106);
and U7525 (N_7525,N_6324,N_6980);
and U7526 (N_7526,N_6851,N_6518);
nand U7527 (N_7527,N_6781,N_6943);
nand U7528 (N_7528,N_6868,N_6056);
or U7529 (N_7529,N_6877,N_6731);
xnor U7530 (N_7530,N_6320,N_6156);
xnor U7531 (N_7531,N_6078,N_6996);
xnor U7532 (N_7532,N_6265,N_6875);
nor U7533 (N_7533,N_6539,N_6511);
xnor U7534 (N_7534,N_6427,N_6016);
and U7535 (N_7535,N_6125,N_6844);
nor U7536 (N_7536,N_6545,N_6315);
or U7537 (N_7537,N_6822,N_6386);
nor U7538 (N_7538,N_6863,N_6444);
nor U7539 (N_7539,N_6081,N_6217);
or U7540 (N_7540,N_6711,N_6324);
and U7541 (N_7541,N_6322,N_6223);
xor U7542 (N_7542,N_6707,N_6790);
nor U7543 (N_7543,N_6532,N_6041);
xnor U7544 (N_7544,N_6257,N_6819);
xnor U7545 (N_7545,N_6495,N_6522);
nand U7546 (N_7546,N_6111,N_6792);
nor U7547 (N_7547,N_6007,N_6755);
xor U7548 (N_7548,N_6755,N_6300);
and U7549 (N_7549,N_6465,N_6118);
nor U7550 (N_7550,N_6301,N_6769);
nor U7551 (N_7551,N_6400,N_6898);
xnor U7552 (N_7552,N_6060,N_6100);
nor U7553 (N_7553,N_6381,N_6265);
or U7554 (N_7554,N_6842,N_6351);
nor U7555 (N_7555,N_6187,N_6673);
or U7556 (N_7556,N_6928,N_6786);
nand U7557 (N_7557,N_6166,N_6948);
or U7558 (N_7558,N_6503,N_6336);
xor U7559 (N_7559,N_6334,N_6389);
nand U7560 (N_7560,N_6943,N_6853);
or U7561 (N_7561,N_6238,N_6401);
and U7562 (N_7562,N_6220,N_6823);
and U7563 (N_7563,N_6478,N_6170);
or U7564 (N_7564,N_6300,N_6308);
nand U7565 (N_7565,N_6430,N_6147);
and U7566 (N_7566,N_6442,N_6846);
and U7567 (N_7567,N_6622,N_6003);
or U7568 (N_7568,N_6672,N_6090);
or U7569 (N_7569,N_6938,N_6881);
or U7570 (N_7570,N_6381,N_6091);
and U7571 (N_7571,N_6252,N_6257);
or U7572 (N_7572,N_6251,N_6143);
nor U7573 (N_7573,N_6974,N_6171);
xor U7574 (N_7574,N_6670,N_6146);
nor U7575 (N_7575,N_6291,N_6712);
nor U7576 (N_7576,N_6896,N_6637);
xnor U7577 (N_7577,N_6059,N_6007);
and U7578 (N_7578,N_6398,N_6287);
xor U7579 (N_7579,N_6054,N_6287);
nor U7580 (N_7580,N_6180,N_6536);
or U7581 (N_7581,N_6506,N_6270);
xor U7582 (N_7582,N_6128,N_6870);
or U7583 (N_7583,N_6525,N_6705);
or U7584 (N_7584,N_6008,N_6649);
nor U7585 (N_7585,N_6616,N_6294);
and U7586 (N_7586,N_6588,N_6363);
xnor U7587 (N_7587,N_6566,N_6362);
and U7588 (N_7588,N_6459,N_6866);
and U7589 (N_7589,N_6300,N_6507);
nand U7590 (N_7590,N_6287,N_6713);
nand U7591 (N_7591,N_6949,N_6507);
nor U7592 (N_7592,N_6589,N_6055);
nand U7593 (N_7593,N_6386,N_6573);
nand U7594 (N_7594,N_6720,N_6977);
nor U7595 (N_7595,N_6083,N_6165);
nand U7596 (N_7596,N_6061,N_6832);
nor U7597 (N_7597,N_6785,N_6217);
and U7598 (N_7598,N_6309,N_6105);
or U7599 (N_7599,N_6397,N_6443);
nor U7600 (N_7600,N_6694,N_6298);
and U7601 (N_7601,N_6351,N_6805);
and U7602 (N_7602,N_6105,N_6649);
or U7603 (N_7603,N_6701,N_6206);
xnor U7604 (N_7604,N_6705,N_6396);
nand U7605 (N_7605,N_6967,N_6458);
and U7606 (N_7606,N_6003,N_6358);
xor U7607 (N_7607,N_6079,N_6463);
nand U7608 (N_7608,N_6098,N_6645);
xor U7609 (N_7609,N_6843,N_6111);
xor U7610 (N_7610,N_6052,N_6774);
and U7611 (N_7611,N_6331,N_6677);
and U7612 (N_7612,N_6142,N_6672);
xnor U7613 (N_7613,N_6145,N_6182);
or U7614 (N_7614,N_6618,N_6802);
nor U7615 (N_7615,N_6606,N_6096);
nor U7616 (N_7616,N_6144,N_6545);
xnor U7617 (N_7617,N_6032,N_6047);
nand U7618 (N_7618,N_6454,N_6274);
nor U7619 (N_7619,N_6455,N_6988);
nor U7620 (N_7620,N_6244,N_6616);
xor U7621 (N_7621,N_6200,N_6904);
nand U7622 (N_7622,N_6177,N_6047);
xor U7623 (N_7623,N_6199,N_6664);
xnor U7624 (N_7624,N_6553,N_6448);
xor U7625 (N_7625,N_6838,N_6301);
nand U7626 (N_7626,N_6128,N_6418);
nor U7627 (N_7627,N_6597,N_6652);
and U7628 (N_7628,N_6569,N_6959);
or U7629 (N_7629,N_6894,N_6195);
and U7630 (N_7630,N_6471,N_6117);
nor U7631 (N_7631,N_6919,N_6250);
nand U7632 (N_7632,N_6269,N_6672);
nor U7633 (N_7633,N_6208,N_6104);
nand U7634 (N_7634,N_6923,N_6627);
nor U7635 (N_7635,N_6411,N_6860);
nand U7636 (N_7636,N_6117,N_6150);
nand U7637 (N_7637,N_6487,N_6327);
nand U7638 (N_7638,N_6362,N_6644);
nand U7639 (N_7639,N_6531,N_6823);
nor U7640 (N_7640,N_6141,N_6732);
nand U7641 (N_7641,N_6717,N_6442);
and U7642 (N_7642,N_6335,N_6392);
or U7643 (N_7643,N_6881,N_6116);
nor U7644 (N_7644,N_6771,N_6051);
or U7645 (N_7645,N_6479,N_6138);
or U7646 (N_7646,N_6183,N_6362);
nor U7647 (N_7647,N_6198,N_6566);
and U7648 (N_7648,N_6321,N_6618);
nand U7649 (N_7649,N_6452,N_6823);
nand U7650 (N_7650,N_6598,N_6434);
and U7651 (N_7651,N_6456,N_6291);
or U7652 (N_7652,N_6918,N_6704);
nor U7653 (N_7653,N_6319,N_6140);
and U7654 (N_7654,N_6233,N_6784);
or U7655 (N_7655,N_6616,N_6221);
or U7656 (N_7656,N_6936,N_6900);
or U7657 (N_7657,N_6211,N_6021);
and U7658 (N_7658,N_6387,N_6408);
nor U7659 (N_7659,N_6349,N_6978);
and U7660 (N_7660,N_6286,N_6695);
or U7661 (N_7661,N_6755,N_6040);
or U7662 (N_7662,N_6183,N_6952);
or U7663 (N_7663,N_6025,N_6547);
or U7664 (N_7664,N_6145,N_6571);
nor U7665 (N_7665,N_6305,N_6991);
or U7666 (N_7666,N_6150,N_6421);
and U7667 (N_7667,N_6198,N_6281);
nand U7668 (N_7668,N_6580,N_6404);
nand U7669 (N_7669,N_6708,N_6414);
xor U7670 (N_7670,N_6030,N_6182);
and U7671 (N_7671,N_6031,N_6395);
or U7672 (N_7672,N_6549,N_6873);
nand U7673 (N_7673,N_6844,N_6415);
nand U7674 (N_7674,N_6149,N_6322);
or U7675 (N_7675,N_6528,N_6136);
nand U7676 (N_7676,N_6555,N_6630);
nor U7677 (N_7677,N_6369,N_6753);
nand U7678 (N_7678,N_6142,N_6376);
xor U7679 (N_7679,N_6977,N_6497);
and U7680 (N_7680,N_6673,N_6902);
nor U7681 (N_7681,N_6567,N_6159);
nand U7682 (N_7682,N_6319,N_6407);
nor U7683 (N_7683,N_6754,N_6621);
xor U7684 (N_7684,N_6509,N_6429);
and U7685 (N_7685,N_6183,N_6736);
nor U7686 (N_7686,N_6557,N_6731);
and U7687 (N_7687,N_6793,N_6823);
and U7688 (N_7688,N_6880,N_6474);
xor U7689 (N_7689,N_6764,N_6688);
nand U7690 (N_7690,N_6016,N_6096);
nand U7691 (N_7691,N_6941,N_6593);
nor U7692 (N_7692,N_6190,N_6311);
and U7693 (N_7693,N_6370,N_6234);
and U7694 (N_7694,N_6259,N_6738);
nand U7695 (N_7695,N_6273,N_6120);
or U7696 (N_7696,N_6807,N_6822);
nor U7697 (N_7697,N_6072,N_6724);
nand U7698 (N_7698,N_6752,N_6921);
and U7699 (N_7699,N_6234,N_6721);
nor U7700 (N_7700,N_6966,N_6317);
xnor U7701 (N_7701,N_6833,N_6226);
nor U7702 (N_7702,N_6093,N_6243);
or U7703 (N_7703,N_6577,N_6504);
or U7704 (N_7704,N_6167,N_6472);
xnor U7705 (N_7705,N_6890,N_6146);
nor U7706 (N_7706,N_6921,N_6396);
and U7707 (N_7707,N_6950,N_6883);
or U7708 (N_7708,N_6997,N_6256);
xnor U7709 (N_7709,N_6696,N_6262);
and U7710 (N_7710,N_6343,N_6997);
and U7711 (N_7711,N_6843,N_6113);
or U7712 (N_7712,N_6511,N_6724);
and U7713 (N_7713,N_6232,N_6914);
nand U7714 (N_7714,N_6231,N_6503);
nand U7715 (N_7715,N_6012,N_6499);
nand U7716 (N_7716,N_6321,N_6908);
or U7717 (N_7717,N_6845,N_6182);
or U7718 (N_7718,N_6838,N_6599);
nor U7719 (N_7719,N_6491,N_6991);
nor U7720 (N_7720,N_6783,N_6891);
or U7721 (N_7721,N_6543,N_6231);
xnor U7722 (N_7722,N_6317,N_6901);
nor U7723 (N_7723,N_6897,N_6991);
nor U7724 (N_7724,N_6438,N_6175);
nand U7725 (N_7725,N_6650,N_6089);
xnor U7726 (N_7726,N_6104,N_6209);
or U7727 (N_7727,N_6381,N_6154);
nand U7728 (N_7728,N_6417,N_6203);
and U7729 (N_7729,N_6173,N_6893);
or U7730 (N_7730,N_6797,N_6946);
nor U7731 (N_7731,N_6659,N_6691);
nand U7732 (N_7732,N_6456,N_6177);
and U7733 (N_7733,N_6843,N_6359);
and U7734 (N_7734,N_6463,N_6709);
nor U7735 (N_7735,N_6707,N_6075);
and U7736 (N_7736,N_6761,N_6892);
and U7737 (N_7737,N_6400,N_6706);
or U7738 (N_7738,N_6872,N_6475);
nand U7739 (N_7739,N_6980,N_6677);
nand U7740 (N_7740,N_6786,N_6519);
nand U7741 (N_7741,N_6299,N_6151);
xor U7742 (N_7742,N_6899,N_6573);
xor U7743 (N_7743,N_6152,N_6476);
and U7744 (N_7744,N_6884,N_6428);
or U7745 (N_7745,N_6789,N_6956);
nor U7746 (N_7746,N_6591,N_6734);
nor U7747 (N_7747,N_6061,N_6170);
nand U7748 (N_7748,N_6003,N_6713);
nand U7749 (N_7749,N_6037,N_6669);
nand U7750 (N_7750,N_6190,N_6730);
xnor U7751 (N_7751,N_6043,N_6469);
or U7752 (N_7752,N_6512,N_6815);
nand U7753 (N_7753,N_6796,N_6983);
and U7754 (N_7754,N_6456,N_6865);
and U7755 (N_7755,N_6232,N_6615);
or U7756 (N_7756,N_6547,N_6915);
nand U7757 (N_7757,N_6241,N_6874);
and U7758 (N_7758,N_6466,N_6476);
or U7759 (N_7759,N_6415,N_6610);
nor U7760 (N_7760,N_6093,N_6505);
xnor U7761 (N_7761,N_6691,N_6879);
and U7762 (N_7762,N_6620,N_6709);
and U7763 (N_7763,N_6389,N_6518);
xnor U7764 (N_7764,N_6238,N_6171);
nor U7765 (N_7765,N_6984,N_6121);
nand U7766 (N_7766,N_6862,N_6112);
and U7767 (N_7767,N_6392,N_6155);
nor U7768 (N_7768,N_6605,N_6256);
or U7769 (N_7769,N_6652,N_6821);
nor U7770 (N_7770,N_6347,N_6792);
nand U7771 (N_7771,N_6336,N_6005);
nor U7772 (N_7772,N_6907,N_6911);
or U7773 (N_7773,N_6722,N_6894);
and U7774 (N_7774,N_6318,N_6407);
and U7775 (N_7775,N_6897,N_6407);
and U7776 (N_7776,N_6062,N_6200);
nand U7777 (N_7777,N_6137,N_6460);
and U7778 (N_7778,N_6964,N_6697);
and U7779 (N_7779,N_6666,N_6082);
nand U7780 (N_7780,N_6707,N_6499);
nand U7781 (N_7781,N_6696,N_6036);
xnor U7782 (N_7782,N_6012,N_6478);
nand U7783 (N_7783,N_6703,N_6638);
nor U7784 (N_7784,N_6434,N_6237);
nand U7785 (N_7785,N_6570,N_6221);
nor U7786 (N_7786,N_6080,N_6350);
or U7787 (N_7787,N_6575,N_6742);
nor U7788 (N_7788,N_6692,N_6499);
or U7789 (N_7789,N_6553,N_6127);
nor U7790 (N_7790,N_6400,N_6938);
nand U7791 (N_7791,N_6484,N_6023);
nor U7792 (N_7792,N_6180,N_6914);
nand U7793 (N_7793,N_6731,N_6209);
xnor U7794 (N_7794,N_6811,N_6268);
xnor U7795 (N_7795,N_6801,N_6854);
nand U7796 (N_7796,N_6283,N_6275);
xnor U7797 (N_7797,N_6247,N_6726);
xor U7798 (N_7798,N_6525,N_6629);
nor U7799 (N_7799,N_6269,N_6996);
xor U7800 (N_7800,N_6094,N_6903);
nand U7801 (N_7801,N_6464,N_6325);
xnor U7802 (N_7802,N_6629,N_6548);
nor U7803 (N_7803,N_6195,N_6080);
and U7804 (N_7804,N_6833,N_6811);
nand U7805 (N_7805,N_6595,N_6991);
and U7806 (N_7806,N_6216,N_6677);
and U7807 (N_7807,N_6139,N_6049);
xor U7808 (N_7808,N_6642,N_6548);
or U7809 (N_7809,N_6317,N_6870);
nand U7810 (N_7810,N_6728,N_6538);
xor U7811 (N_7811,N_6329,N_6830);
nand U7812 (N_7812,N_6642,N_6288);
nand U7813 (N_7813,N_6628,N_6031);
nor U7814 (N_7814,N_6392,N_6398);
nand U7815 (N_7815,N_6733,N_6093);
xor U7816 (N_7816,N_6160,N_6780);
nand U7817 (N_7817,N_6791,N_6991);
nor U7818 (N_7818,N_6440,N_6413);
nand U7819 (N_7819,N_6461,N_6161);
xor U7820 (N_7820,N_6494,N_6825);
or U7821 (N_7821,N_6778,N_6341);
and U7822 (N_7822,N_6410,N_6456);
and U7823 (N_7823,N_6184,N_6466);
nand U7824 (N_7824,N_6797,N_6992);
and U7825 (N_7825,N_6215,N_6433);
nand U7826 (N_7826,N_6671,N_6592);
or U7827 (N_7827,N_6198,N_6152);
or U7828 (N_7828,N_6195,N_6724);
or U7829 (N_7829,N_6174,N_6841);
and U7830 (N_7830,N_6691,N_6933);
nor U7831 (N_7831,N_6415,N_6849);
and U7832 (N_7832,N_6547,N_6023);
nor U7833 (N_7833,N_6763,N_6403);
and U7834 (N_7834,N_6264,N_6597);
and U7835 (N_7835,N_6802,N_6093);
nand U7836 (N_7836,N_6678,N_6271);
xnor U7837 (N_7837,N_6799,N_6221);
nor U7838 (N_7838,N_6545,N_6739);
and U7839 (N_7839,N_6369,N_6206);
xnor U7840 (N_7840,N_6171,N_6325);
and U7841 (N_7841,N_6873,N_6896);
and U7842 (N_7842,N_6816,N_6089);
or U7843 (N_7843,N_6530,N_6576);
nor U7844 (N_7844,N_6532,N_6908);
and U7845 (N_7845,N_6409,N_6963);
nor U7846 (N_7846,N_6847,N_6309);
or U7847 (N_7847,N_6130,N_6498);
xnor U7848 (N_7848,N_6883,N_6834);
nand U7849 (N_7849,N_6313,N_6422);
xor U7850 (N_7850,N_6254,N_6435);
and U7851 (N_7851,N_6782,N_6228);
xor U7852 (N_7852,N_6961,N_6706);
xnor U7853 (N_7853,N_6905,N_6833);
xnor U7854 (N_7854,N_6129,N_6380);
nand U7855 (N_7855,N_6617,N_6566);
or U7856 (N_7856,N_6293,N_6944);
and U7857 (N_7857,N_6365,N_6061);
or U7858 (N_7858,N_6917,N_6180);
xnor U7859 (N_7859,N_6767,N_6173);
xnor U7860 (N_7860,N_6984,N_6230);
and U7861 (N_7861,N_6117,N_6171);
nand U7862 (N_7862,N_6733,N_6130);
nand U7863 (N_7863,N_6003,N_6185);
nand U7864 (N_7864,N_6801,N_6101);
and U7865 (N_7865,N_6420,N_6688);
and U7866 (N_7866,N_6814,N_6894);
and U7867 (N_7867,N_6936,N_6640);
or U7868 (N_7868,N_6937,N_6047);
nand U7869 (N_7869,N_6276,N_6338);
nand U7870 (N_7870,N_6609,N_6508);
and U7871 (N_7871,N_6958,N_6384);
nand U7872 (N_7872,N_6502,N_6267);
or U7873 (N_7873,N_6502,N_6595);
and U7874 (N_7874,N_6648,N_6543);
and U7875 (N_7875,N_6000,N_6238);
nand U7876 (N_7876,N_6412,N_6227);
nor U7877 (N_7877,N_6859,N_6465);
xor U7878 (N_7878,N_6487,N_6429);
xor U7879 (N_7879,N_6773,N_6499);
or U7880 (N_7880,N_6580,N_6046);
nor U7881 (N_7881,N_6541,N_6999);
nand U7882 (N_7882,N_6715,N_6265);
and U7883 (N_7883,N_6921,N_6596);
nand U7884 (N_7884,N_6412,N_6034);
xnor U7885 (N_7885,N_6924,N_6586);
nand U7886 (N_7886,N_6348,N_6430);
nor U7887 (N_7887,N_6151,N_6214);
or U7888 (N_7888,N_6030,N_6914);
and U7889 (N_7889,N_6977,N_6797);
nand U7890 (N_7890,N_6562,N_6973);
or U7891 (N_7891,N_6487,N_6712);
and U7892 (N_7892,N_6611,N_6255);
nand U7893 (N_7893,N_6449,N_6953);
or U7894 (N_7894,N_6989,N_6977);
xor U7895 (N_7895,N_6969,N_6165);
xor U7896 (N_7896,N_6209,N_6080);
xnor U7897 (N_7897,N_6849,N_6857);
and U7898 (N_7898,N_6548,N_6951);
xnor U7899 (N_7899,N_6667,N_6229);
nor U7900 (N_7900,N_6553,N_6945);
xor U7901 (N_7901,N_6218,N_6965);
nand U7902 (N_7902,N_6171,N_6873);
nand U7903 (N_7903,N_6898,N_6088);
xnor U7904 (N_7904,N_6953,N_6790);
and U7905 (N_7905,N_6618,N_6547);
nor U7906 (N_7906,N_6781,N_6279);
nor U7907 (N_7907,N_6096,N_6027);
and U7908 (N_7908,N_6359,N_6816);
and U7909 (N_7909,N_6071,N_6942);
and U7910 (N_7910,N_6213,N_6569);
and U7911 (N_7911,N_6831,N_6450);
nor U7912 (N_7912,N_6639,N_6099);
nor U7913 (N_7913,N_6711,N_6012);
and U7914 (N_7914,N_6069,N_6613);
xor U7915 (N_7915,N_6424,N_6609);
and U7916 (N_7916,N_6692,N_6418);
or U7917 (N_7917,N_6923,N_6839);
nand U7918 (N_7918,N_6913,N_6449);
or U7919 (N_7919,N_6784,N_6755);
nand U7920 (N_7920,N_6405,N_6627);
and U7921 (N_7921,N_6150,N_6606);
and U7922 (N_7922,N_6148,N_6300);
or U7923 (N_7923,N_6520,N_6296);
nor U7924 (N_7924,N_6709,N_6283);
or U7925 (N_7925,N_6075,N_6684);
nor U7926 (N_7926,N_6742,N_6552);
or U7927 (N_7927,N_6299,N_6324);
or U7928 (N_7928,N_6715,N_6412);
xnor U7929 (N_7929,N_6423,N_6632);
xor U7930 (N_7930,N_6011,N_6049);
or U7931 (N_7931,N_6963,N_6503);
nor U7932 (N_7932,N_6841,N_6120);
and U7933 (N_7933,N_6512,N_6130);
and U7934 (N_7934,N_6858,N_6869);
and U7935 (N_7935,N_6078,N_6543);
xnor U7936 (N_7936,N_6289,N_6732);
nand U7937 (N_7937,N_6062,N_6456);
xor U7938 (N_7938,N_6673,N_6367);
and U7939 (N_7939,N_6774,N_6508);
nor U7940 (N_7940,N_6416,N_6517);
nand U7941 (N_7941,N_6916,N_6719);
and U7942 (N_7942,N_6392,N_6110);
nor U7943 (N_7943,N_6707,N_6777);
xnor U7944 (N_7944,N_6715,N_6448);
or U7945 (N_7945,N_6004,N_6541);
nor U7946 (N_7946,N_6244,N_6165);
xnor U7947 (N_7947,N_6977,N_6844);
or U7948 (N_7948,N_6557,N_6501);
and U7949 (N_7949,N_6435,N_6554);
and U7950 (N_7950,N_6482,N_6479);
nor U7951 (N_7951,N_6511,N_6630);
or U7952 (N_7952,N_6725,N_6023);
xnor U7953 (N_7953,N_6046,N_6956);
xor U7954 (N_7954,N_6704,N_6642);
nand U7955 (N_7955,N_6006,N_6029);
xor U7956 (N_7956,N_6317,N_6608);
or U7957 (N_7957,N_6657,N_6718);
nor U7958 (N_7958,N_6251,N_6782);
xor U7959 (N_7959,N_6506,N_6246);
and U7960 (N_7960,N_6347,N_6579);
xor U7961 (N_7961,N_6332,N_6581);
and U7962 (N_7962,N_6864,N_6033);
nand U7963 (N_7963,N_6597,N_6334);
nand U7964 (N_7964,N_6647,N_6935);
or U7965 (N_7965,N_6084,N_6190);
and U7966 (N_7966,N_6768,N_6748);
xnor U7967 (N_7967,N_6234,N_6921);
and U7968 (N_7968,N_6945,N_6430);
nand U7969 (N_7969,N_6974,N_6893);
nand U7970 (N_7970,N_6328,N_6042);
or U7971 (N_7971,N_6377,N_6901);
xnor U7972 (N_7972,N_6299,N_6169);
xnor U7973 (N_7973,N_6948,N_6389);
nand U7974 (N_7974,N_6869,N_6251);
nand U7975 (N_7975,N_6480,N_6644);
xor U7976 (N_7976,N_6083,N_6769);
nand U7977 (N_7977,N_6606,N_6246);
or U7978 (N_7978,N_6774,N_6529);
and U7979 (N_7979,N_6162,N_6873);
nand U7980 (N_7980,N_6468,N_6613);
nand U7981 (N_7981,N_6222,N_6255);
xnor U7982 (N_7982,N_6526,N_6614);
or U7983 (N_7983,N_6976,N_6020);
or U7984 (N_7984,N_6965,N_6316);
nor U7985 (N_7985,N_6473,N_6512);
nand U7986 (N_7986,N_6110,N_6577);
nor U7987 (N_7987,N_6555,N_6561);
nand U7988 (N_7988,N_6253,N_6669);
nor U7989 (N_7989,N_6807,N_6318);
nand U7990 (N_7990,N_6431,N_6382);
or U7991 (N_7991,N_6213,N_6214);
nand U7992 (N_7992,N_6439,N_6186);
and U7993 (N_7993,N_6444,N_6456);
nor U7994 (N_7994,N_6220,N_6759);
and U7995 (N_7995,N_6557,N_6121);
and U7996 (N_7996,N_6869,N_6288);
xor U7997 (N_7997,N_6208,N_6654);
nor U7998 (N_7998,N_6880,N_6416);
or U7999 (N_7999,N_6046,N_6022);
nor U8000 (N_8000,N_7305,N_7799);
nor U8001 (N_8001,N_7037,N_7947);
and U8002 (N_8002,N_7998,N_7743);
and U8003 (N_8003,N_7185,N_7670);
nand U8004 (N_8004,N_7414,N_7661);
xnor U8005 (N_8005,N_7088,N_7957);
or U8006 (N_8006,N_7331,N_7677);
nor U8007 (N_8007,N_7004,N_7736);
xor U8008 (N_8008,N_7649,N_7558);
or U8009 (N_8009,N_7692,N_7653);
and U8010 (N_8010,N_7448,N_7808);
xor U8011 (N_8011,N_7800,N_7499);
xor U8012 (N_8012,N_7474,N_7607);
or U8013 (N_8013,N_7408,N_7481);
nand U8014 (N_8014,N_7456,N_7547);
or U8015 (N_8015,N_7500,N_7564);
nor U8016 (N_8016,N_7232,N_7893);
and U8017 (N_8017,N_7503,N_7440);
nand U8018 (N_8018,N_7156,N_7952);
and U8019 (N_8019,N_7642,N_7300);
and U8020 (N_8020,N_7195,N_7626);
or U8021 (N_8021,N_7805,N_7086);
nand U8022 (N_8022,N_7052,N_7497);
nand U8023 (N_8023,N_7719,N_7676);
and U8024 (N_8024,N_7884,N_7298);
nand U8025 (N_8025,N_7940,N_7760);
nor U8026 (N_8026,N_7355,N_7202);
nor U8027 (N_8027,N_7365,N_7748);
and U8028 (N_8028,N_7010,N_7686);
xor U8029 (N_8029,N_7096,N_7917);
nor U8030 (N_8030,N_7356,N_7269);
nor U8031 (N_8031,N_7629,N_7941);
or U8032 (N_8032,N_7991,N_7498);
nand U8033 (N_8033,N_7566,N_7031);
nand U8034 (N_8034,N_7048,N_7915);
or U8035 (N_8035,N_7410,N_7039);
xor U8036 (N_8036,N_7099,N_7869);
nor U8037 (N_8037,N_7621,N_7726);
nor U8038 (N_8038,N_7264,N_7696);
xor U8039 (N_8039,N_7506,N_7775);
or U8040 (N_8040,N_7371,N_7296);
nor U8041 (N_8041,N_7703,N_7336);
nor U8042 (N_8042,N_7059,N_7971);
nand U8043 (N_8043,N_7055,N_7938);
and U8044 (N_8044,N_7276,N_7322);
xor U8045 (N_8045,N_7681,N_7081);
nor U8046 (N_8046,N_7572,N_7043);
and U8047 (N_8047,N_7975,N_7773);
and U8048 (N_8048,N_7718,N_7482);
nor U8049 (N_8049,N_7980,N_7426);
nand U8050 (N_8050,N_7476,N_7458);
or U8051 (N_8051,N_7981,N_7928);
or U8052 (N_8052,N_7823,N_7578);
and U8053 (N_8053,N_7142,N_7892);
nor U8054 (N_8054,N_7242,N_7575);
xor U8055 (N_8055,N_7285,N_7400);
xnor U8056 (N_8056,N_7449,N_7491);
nand U8057 (N_8057,N_7749,N_7699);
nor U8058 (N_8058,N_7279,N_7023);
nand U8059 (N_8059,N_7071,N_7047);
nor U8060 (N_8060,N_7544,N_7453);
nor U8061 (N_8061,N_7271,N_7493);
xor U8062 (N_8062,N_7148,N_7781);
and U8063 (N_8063,N_7916,N_7537);
xor U8064 (N_8064,N_7252,N_7559);
xnor U8065 (N_8065,N_7581,N_7118);
nand U8066 (N_8066,N_7469,N_7442);
and U8067 (N_8067,N_7890,N_7046);
and U8068 (N_8068,N_7894,N_7600);
and U8069 (N_8069,N_7309,N_7223);
xnor U8070 (N_8070,N_7210,N_7967);
or U8071 (N_8071,N_7423,N_7465);
or U8072 (N_8072,N_7119,N_7635);
or U8073 (N_8073,N_7644,N_7138);
nor U8074 (N_8074,N_7652,N_7831);
and U8075 (N_8075,N_7092,N_7791);
nor U8076 (N_8076,N_7253,N_7844);
and U8077 (N_8077,N_7974,N_7204);
nor U8078 (N_8078,N_7530,N_7602);
xnor U8079 (N_8079,N_7539,N_7714);
xnor U8080 (N_8080,N_7648,N_7673);
nor U8081 (N_8081,N_7970,N_7401);
and U8082 (N_8082,N_7815,N_7872);
nand U8083 (N_8083,N_7058,N_7238);
nand U8084 (N_8084,N_7294,N_7307);
or U8085 (N_8085,N_7066,N_7394);
nand U8086 (N_8086,N_7814,N_7067);
nand U8087 (N_8087,N_7985,N_7885);
nand U8088 (N_8088,N_7467,N_7295);
nor U8089 (N_8089,N_7793,N_7550);
nor U8090 (N_8090,N_7524,N_7083);
and U8091 (N_8091,N_7640,N_7461);
xor U8092 (N_8092,N_7505,N_7116);
xor U8093 (N_8093,N_7929,N_7728);
nor U8094 (N_8094,N_7310,N_7430);
xnor U8095 (N_8095,N_7669,N_7839);
nand U8096 (N_8096,N_7645,N_7035);
nor U8097 (N_8097,N_7886,N_7016);
and U8098 (N_8098,N_7569,N_7533);
or U8099 (N_8099,N_7989,N_7175);
xnor U8100 (N_8100,N_7447,N_7567);
xnor U8101 (N_8101,N_7209,N_7361);
nand U8102 (N_8102,N_7756,N_7965);
or U8103 (N_8103,N_7996,N_7406);
nor U8104 (N_8104,N_7571,N_7211);
nand U8105 (N_8105,N_7326,N_7995);
xnor U8106 (N_8106,N_7802,N_7022);
and U8107 (N_8107,N_7437,N_7806);
nor U8108 (N_8108,N_7056,N_7552);
nand U8109 (N_8109,N_7249,N_7381);
nor U8110 (N_8110,N_7280,N_7742);
and U8111 (N_8111,N_7289,N_7450);
and U8112 (N_8112,N_7932,N_7688);
or U8113 (N_8113,N_7427,N_7701);
nor U8114 (N_8114,N_7656,N_7638);
or U8115 (N_8115,N_7105,N_7784);
and U8116 (N_8116,N_7866,N_7883);
xor U8117 (N_8117,N_7245,N_7093);
and U8118 (N_8118,N_7032,N_7360);
xnor U8119 (N_8119,N_7944,N_7682);
nor U8120 (N_8120,N_7036,N_7299);
xnor U8121 (N_8121,N_7608,N_7378);
and U8122 (N_8122,N_7939,N_7191);
nand U8123 (N_8123,N_7573,N_7794);
nand U8124 (N_8124,N_7949,N_7910);
and U8125 (N_8125,N_7229,N_7856);
nand U8126 (N_8126,N_7315,N_7766);
or U8127 (N_8127,N_7759,N_7895);
or U8128 (N_8128,N_7170,N_7704);
nor U8129 (N_8129,N_7841,N_7412);
or U8130 (N_8130,N_7472,N_7553);
and U8131 (N_8131,N_7897,N_7542);
and U8132 (N_8132,N_7934,N_7377);
nand U8133 (N_8133,N_7863,N_7405);
xnor U8134 (N_8134,N_7370,N_7404);
or U8135 (N_8135,N_7950,N_7040);
nand U8136 (N_8136,N_7145,N_7616);
or U8137 (N_8137,N_7327,N_7140);
or U8138 (N_8138,N_7876,N_7376);
nand U8139 (N_8139,N_7297,N_7843);
xnor U8140 (N_8140,N_7065,N_7132);
and U8141 (N_8141,N_7134,N_7684);
nand U8142 (N_8142,N_7538,N_7987);
nand U8143 (N_8143,N_7250,N_7108);
xor U8144 (N_8144,N_7333,N_7512);
nand U8145 (N_8145,N_7804,N_7779);
xor U8146 (N_8146,N_7477,N_7655);
nand U8147 (N_8147,N_7842,N_7109);
nand U8148 (N_8148,N_7254,N_7918);
nor U8149 (N_8149,N_7772,N_7617);
or U8150 (N_8150,N_7694,N_7343);
nand U8151 (N_8151,N_7601,N_7339);
xor U8152 (N_8152,N_7903,N_7671);
or U8153 (N_8153,N_7383,N_7597);
and U8154 (N_8154,N_7479,N_7992);
and U8155 (N_8155,N_7787,N_7041);
xnor U8156 (N_8156,N_7531,N_7197);
or U8157 (N_8157,N_7536,N_7064);
and U8158 (N_8158,N_7292,N_7741);
xor U8159 (N_8159,N_7125,N_7785);
nand U8160 (N_8160,N_7735,N_7180);
nand U8161 (N_8161,N_7758,N_7009);
xor U8162 (N_8162,N_7389,N_7062);
and U8163 (N_8163,N_7146,N_7015);
nand U8164 (N_8164,N_7877,N_7751);
or U8165 (N_8165,N_7433,N_7402);
nand U8166 (N_8166,N_7359,N_7001);
nand U8167 (N_8167,N_7962,N_7727);
xnor U8168 (N_8168,N_7155,N_7979);
and U8169 (N_8169,N_7659,N_7786);
nor U8170 (N_8170,N_7364,N_7446);
or U8171 (N_8171,N_7907,N_7958);
nand U8172 (N_8172,N_7610,N_7809);
nand U8173 (N_8173,N_7258,N_7077);
or U8174 (N_8174,N_7836,N_7501);
or U8175 (N_8175,N_7054,N_7328);
nand U8176 (N_8176,N_7923,N_7392);
nor U8177 (N_8177,N_7922,N_7205);
and U8178 (N_8178,N_7122,N_7545);
and U8179 (N_8179,N_7919,N_7921);
nand U8180 (N_8180,N_7619,N_7777);
or U8181 (N_8181,N_7018,N_7445);
and U8182 (N_8182,N_7582,N_7455);
nor U8183 (N_8183,N_7367,N_7709);
nor U8184 (N_8184,N_7591,N_7434);
nor U8185 (N_8185,N_7137,N_7090);
nand U8186 (N_8186,N_7261,N_7424);
and U8187 (N_8187,N_7340,N_7335);
nor U8188 (N_8188,N_7854,N_7855);
xnor U8189 (N_8189,N_7259,N_7675);
and U8190 (N_8190,N_7691,N_7990);
xnor U8191 (N_8191,N_7165,N_7945);
or U8192 (N_8192,N_7960,N_7951);
xor U8193 (N_8193,N_7080,N_7959);
nor U8194 (N_8194,N_7768,N_7126);
and U8195 (N_8195,N_7710,N_7592);
and U8196 (N_8196,N_7935,N_7061);
or U8197 (N_8197,N_7235,N_7650);
xnor U8198 (N_8198,N_7002,N_7632);
xnor U8199 (N_8199,N_7633,N_7901);
and U8200 (N_8200,N_7613,N_7593);
or U8201 (N_8201,N_7218,N_7618);
nor U8202 (N_8202,N_7221,N_7712);
nor U8203 (N_8203,N_7820,N_7395);
or U8204 (N_8204,N_7143,N_7576);
or U8205 (N_8205,N_7764,N_7986);
nand U8206 (N_8206,N_7407,N_7312);
and U8207 (N_8207,N_7366,N_7875);
and U8208 (N_8208,N_7717,N_7154);
or U8209 (N_8209,N_7466,N_7181);
nor U8210 (N_8210,N_7308,N_7079);
nand U8211 (N_8211,N_7549,N_7795);
or U8212 (N_8212,N_7111,N_7888);
or U8213 (N_8213,N_7438,N_7347);
nand U8214 (N_8214,N_7139,N_7858);
and U8215 (N_8215,N_7283,N_7431);
and U8216 (N_8216,N_7471,N_7730);
xnor U8217 (N_8217,N_7946,N_7878);
xor U8218 (N_8218,N_7144,N_7612);
or U8219 (N_8219,N_7899,N_7349);
and U8220 (N_8220,N_7630,N_7548);
nor U8221 (N_8221,N_7473,N_7329);
xor U8222 (N_8222,N_7754,N_7291);
or U8223 (N_8223,N_7912,N_7207);
nor U8224 (N_8224,N_7044,N_7783);
xor U8225 (N_8225,N_7818,N_7240);
or U8226 (N_8226,N_7429,N_7819);
nor U8227 (N_8227,N_7487,N_7087);
and U8228 (N_8228,N_7171,N_7006);
xnor U8229 (N_8229,N_7812,N_7273);
xor U8230 (N_8230,N_7925,N_7379);
nand U8231 (N_8231,N_7270,N_7829);
nand U8232 (N_8232,N_7095,N_7492);
xnor U8233 (N_8233,N_7107,N_7237);
xnor U8234 (N_8234,N_7443,N_7849);
or U8235 (N_8235,N_7382,N_7320);
or U8236 (N_8236,N_7225,N_7561);
and U8237 (N_8237,N_7973,N_7452);
xor U8238 (N_8238,N_7346,N_7007);
nor U8239 (N_8239,N_7847,N_7091);
and U8240 (N_8240,N_7387,N_7076);
nor U8241 (N_8241,N_7590,N_7924);
or U8242 (N_8242,N_7603,N_7121);
or U8243 (N_8243,N_7070,N_7464);
and U8244 (N_8244,N_7149,N_7520);
xor U8245 (N_8245,N_7821,N_7129);
xnor U8246 (N_8246,N_7341,N_7337);
or U8247 (N_8247,N_7074,N_7332);
or U8248 (N_8248,N_7789,N_7803);
nand U8249 (N_8249,N_7509,N_7663);
nor U8250 (N_8250,N_7029,N_7599);
and U8251 (N_8251,N_7457,N_7906);
and U8252 (N_8252,N_7374,N_7737);
xor U8253 (N_8253,N_7306,N_7390);
nor U8254 (N_8254,N_7515,N_7828);
nor U8255 (N_8255,N_7200,N_7643);
nor U8256 (N_8256,N_7683,N_7324);
or U8257 (N_8257,N_7051,N_7323);
and U8258 (N_8258,N_7373,N_7516);
nand U8259 (N_8259,N_7215,N_7152);
xor U8260 (N_8260,N_7598,N_7358);
or U8261 (N_8261,N_7075,N_7792);
or U8262 (N_8262,N_7348,N_7251);
xor U8263 (N_8263,N_7428,N_7247);
nand U8264 (N_8264,N_7021,N_7738);
or U8265 (N_8265,N_7117,N_7705);
xnor U8266 (N_8266,N_7848,N_7744);
xor U8267 (N_8267,N_7830,N_7003);
nand U8268 (N_8268,N_7227,N_7120);
xor U8269 (N_8269,N_7089,N_7868);
nor U8270 (N_8270,N_7840,N_7110);
and U8271 (N_8271,N_7199,N_7311);
nor U8272 (N_8272,N_7711,N_7810);
xnor U8273 (N_8273,N_7268,N_7551);
or U8274 (N_8274,N_7005,N_7920);
nor U8275 (N_8275,N_7807,N_7563);
or U8276 (N_8276,N_7303,N_7725);
and U8277 (N_8277,N_7865,N_7475);
nor U8278 (N_8278,N_7033,N_7668);
nor U8279 (N_8279,N_7972,N_7518);
nor U8280 (N_8280,N_7415,N_7679);
and U8281 (N_8281,N_7160,N_7522);
nor U8282 (N_8282,N_7060,N_7157);
or U8283 (N_8283,N_7579,N_7664);
and U8284 (N_8284,N_7565,N_7769);
or U8285 (N_8285,N_7672,N_7724);
xnor U8286 (N_8286,N_7909,N_7931);
and U8287 (N_8287,N_7027,N_7123);
or U8288 (N_8288,N_7186,N_7860);
nor U8289 (N_8289,N_7050,N_7028);
nor U8290 (N_8290,N_7695,N_7462);
or U8291 (N_8291,N_7017,N_7595);
and U8292 (N_8292,N_7720,N_7141);
nor U8293 (N_8293,N_7713,N_7483);
or U8294 (N_8294,N_7024,N_7375);
and U8295 (N_8295,N_7835,N_7263);
xnor U8296 (N_8296,N_7556,N_7274);
nor U8297 (N_8297,N_7224,N_7898);
xor U8298 (N_8298,N_7813,N_7494);
nor U8299 (N_8299,N_7510,N_7338);
xor U8300 (N_8300,N_7167,N_7997);
xnor U8301 (N_8301,N_7179,N_7073);
xnor U8302 (N_8302,N_7385,N_7135);
and U8303 (N_8303,N_7723,N_7441);
or U8304 (N_8304,N_7236,N_7666);
xnor U8305 (N_8305,N_7034,N_7478);
or U8306 (N_8306,N_7063,N_7436);
or U8307 (N_8307,N_7525,N_7026);
xor U8308 (N_8308,N_7905,N_7369);
and U8309 (N_8309,N_7837,N_7459);
xnor U8310 (N_8310,N_7219,N_7774);
and U8311 (N_8311,N_7084,N_7357);
xor U8312 (N_8312,N_7025,N_7557);
or U8313 (N_8313,N_7391,N_7172);
or U8314 (N_8314,N_7584,N_7266);
and U8315 (N_8315,N_7290,N_7966);
or U8316 (N_8316,N_7330,N_7362);
and U8317 (N_8317,N_7614,N_7753);
or U8318 (N_8318,N_7102,N_7214);
or U8319 (N_8319,N_7739,N_7977);
nor U8320 (N_8320,N_7562,N_7293);
xor U8321 (N_8321,N_7902,N_7982);
or U8322 (N_8322,N_7942,N_7241);
or U8323 (N_8323,N_7721,N_7244);
nand U8324 (N_8324,N_7873,N_7284);
and U8325 (N_8325,N_7217,N_7978);
nor U8326 (N_8326,N_7930,N_7313);
or U8327 (N_8327,N_7316,N_7100);
nor U8328 (N_8328,N_7380,N_7496);
xor U8329 (N_8329,N_7072,N_7540);
xnor U8330 (N_8330,N_7716,N_7485);
and U8331 (N_8331,N_7594,N_7586);
xor U8332 (N_8332,N_7286,N_7486);
and U8333 (N_8333,N_7969,N_7489);
nand U8334 (N_8334,N_7127,N_7187);
nor U8335 (N_8335,N_7101,N_7780);
nand U8336 (N_8336,N_7817,N_7319);
xor U8337 (N_8337,N_7451,N_7384);
nand U8338 (N_8338,N_7583,N_7874);
xor U8339 (N_8339,N_7881,N_7519);
or U8340 (N_8340,N_7734,N_7639);
nand U8341 (N_8341,N_7796,N_7272);
nand U8342 (N_8342,N_7243,N_7468);
or U8343 (N_8343,N_7403,N_7816);
xor U8344 (N_8344,N_7689,N_7700);
and U8345 (N_8345,N_7999,N_7954);
nand U8346 (N_8346,N_7317,N_7422);
nor U8347 (N_8347,N_7755,N_7861);
nor U8348 (N_8348,N_7933,N_7103);
nor U8349 (N_8349,N_7707,N_7104);
nand U8350 (N_8350,N_7778,N_7824);
or U8351 (N_8351,N_7220,N_7094);
nand U8352 (N_8352,N_7042,N_7228);
or U8353 (N_8353,N_7488,N_7955);
nor U8354 (N_8354,N_7418,N_7344);
and U8355 (N_8355,N_7641,N_7213);
nor U8356 (N_8356,N_7517,N_7637);
or U8357 (N_8357,N_7771,N_7880);
and U8358 (N_8358,N_7770,N_7541);
or U8359 (N_8359,N_7439,N_7574);
or U8360 (N_8360,N_7417,N_7580);
xnor U8361 (N_8361,N_7715,N_7693);
nand U8362 (N_8362,N_7008,N_7173);
or U8363 (N_8363,N_7685,N_7212);
nand U8364 (N_8364,N_7859,N_7850);
xnor U8365 (N_8365,N_7587,N_7334);
and U8366 (N_8366,N_7150,N_7534);
nor U8367 (N_8367,N_7953,N_7535);
or U8368 (N_8368,N_7948,N_7687);
nand U8369 (N_8369,N_7226,N_7030);
or U8370 (N_8370,N_7560,N_7697);
nor U8371 (N_8371,N_7196,N_7386);
and U8372 (N_8372,N_7879,N_7301);
and U8373 (N_8373,N_7198,N_7124);
and U8374 (N_8374,N_7926,N_7416);
and U8375 (N_8375,N_7421,N_7827);
nand U8376 (N_8376,N_7189,N_7767);
xor U8377 (N_8377,N_7862,N_7068);
xnor U8378 (N_8378,N_7206,N_7190);
or U8379 (N_8379,N_7162,N_7667);
and U8380 (N_8380,N_7019,N_7834);
xor U8381 (N_8381,N_7504,N_7845);
and U8382 (N_8382,N_7397,N_7183);
or U8383 (N_8383,N_7203,N_7904);
or U8384 (N_8384,N_7852,N_7757);
nor U8385 (N_8385,N_7159,N_7702);
xor U8386 (N_8386,N_7811,N_7085);
or U8387 (N_8387,N_7256,N_7976);
nand U8388 (N_8388,N_7624,N_7961);
or U8389 (N_8389,N_7514,N_7413);
and U8390 (N_8390,N_7255,N_7646);
nand U8391 (N_8391,N_7177,N_7246);
nor U8392 (N_8392,N_7889,N_7133);
and U8393 (N_8393,N_7746,N_7623);
nor U8394 (N_8394,N_7106,N_7832);
nand U8395 (N_8395,N_7678,N_7288);
or U8396 (N_8396,N_7984,N_7368);
or U8397 (N_8397,N_7822,N_7636);
nor U8398 (N_8398,N_7523,N_7282);
xor U8399 (N_8399,N_7732,N_7526);
and U8400 (N_8400,N_7262,N_7654);
and U8401 (N_8401,N_7425,N_7216);
and U8402 (N_8402,N_7936,N_7178);
or U8403 (N_8403,N_7484,N_7745);
or U8404 (N_8404,N_7838,N_7882);
or U8405 (N_8405,N_7943,N_7993);
nor U8406 (N_8406,N_7900,N_7013);
xor U8407 (N_8407,N_7853,N_7151);
nor U8408 (N_8408,N_7532,N_7049);
nor U8409 (N_8409,N_7420,N_7511);
or U8410 (N_8410,N_7988,N_7409);
nand U8411 (N_8411,N_7432,N_7166);
or U8412 (N_8412,N_7750,N_7136);
and U8413 (N_8413,N_7012,N_7658);
nor U8414 (N_8414,N_7396,N_7393);
and U8415 (N_8415,N_7870,N_7690);
xnor U8416 (N_8416,N_7731,N_7260);
xor U8417 (N_8417,N_7625,N_7662);
nand U8418 (N_8418,N_7588,N_7363);
nand U8419 (N_8419,N_7752,N_7265);
or U8420 (N_8420,N_7776,N_7570);
and U8421 (N_8421,N_7782,N_7826);
and U8422 (N_8422,N_7867,N_7147);
nand U8423 (N_8423,N_7660,N_7278);
nand U8424 (N_8424,N_7398,N_7069);
nand U8425 (N_8425,N_7609,N_7318);
or U8426 (N_8426,N_7529,N_7729);
xnor U8427 (N_8427,N_7351,N_7543);
nor U8428 (N_8428,N_7082,N_7325);
and U8429 (N_8429,N_7435,N_7761);
nor U8430 (N_8430,N_7763,N_7634);
nor U8431 (N_8431,N_7184,N_7188);
or U8432 (N_8432,N_7937,N_7994);
nand U8433 (N_8433,N_7801,N_7231);
xor U8434 (N_8434,N_7596,N_7887);
and U8435 (N_8435,N_7825,N_7168);
xor U8436 (N_8436,N_7354,N_7508);
nor U8437 (N_8437,N_7321,N_7528);
nor U8438 (N_8438,N_7722,N_7098);
xnor U8439 (N_8439,N_7011,N_7615);
nor U8440 (N_8440,N_7239,N_7747);
and U8441 (N_8441,N_7968,N_7038);
or U8442 (N_8442,N_7192,N_7546);
nor U8443 (N_8443,N_7568,N_7161);
and U8444 (N_8444,N_7097,N_7302);
and U8445 (N_8445,N_7353,N_7740);
nand U8446 (N_8446,N_7201,N_7234);
or U8447 (N_8447,N_7176,N_7680);
and U8448 (N_8448,N_7164,N_7606);
and U8449 (N_8449,N_7604,N_7956);
and U8450 (N_8450,N_7350,N_7502);
xnor U8451 (N_8451,N_7908,N_7577);
or U8452 (N_8452,N_7871,N_7589);
xnor U8453 (N_8453,N_7230,N_7014);
and U8454 (N_8454,N_7495,N_7304);
or U8455 (N_8455,N_7208,N_7163);
and U8456 (N_8456,N_7470,N_7057);
xor U8457 (N_8457,N_7388,N_7647);
xor U8458 (N_8458,N_7411,N_7706);
or U8459 (N_8459,N_7345,N_7846);
xnor U8460 (N_8460,N_7128,N_7605);
and U8461 (N_8461,N_7248,N_7281);
xnor U8462 (N_8462,N_7000,N_7460);
nand U8463 (N_8463,N_7419,N_7622);
nand U8464 (N_8464,N_7267,N_7158);
xor U8465 (N_8465,N_7078,N_7045);
or U8466 (N_8466,N_7233,N_7631);
and U8467 (N_8467,N_7513,N_7927);
and U8468 (N_8468,N_7963,N_7372);
and U8469 (N_8469,N_7444,N_7527);
or U8470 (N_8470,N_7585,N_7480);
or U8471 (N_8471,N_7490,N_7314);
and U8472 (N_8472,N_7708,N_7399);
xnor U8473 (N_8473,N_7275,N_7733);
or U8474 (N_8474,N_7169,N_7911);
nand U8475 (N_8475,N_7113,N_7193);
xor U8476 (N_8476,N_7114,N_7857);
or U8477 (N_8477,N_7277,N_7611);
xnor U8478 (N_8478,N_7182,N_7521);
xnor U8479 (N_8479,N_7112,N_7651);
or U8480 (N_8480,N_7153,N_7765);
or U8481 (N_8481,N_7507,N_7790);
xor U8482 (N_8482,N_7053,N_7674);
or U8483 (N_8483,N_7131,N_7913);
xor U8484 (N_8484,N_7287,N_7194);
xor U8485 (N_8485,N_7020,N_7864);
xnor U8486 (N_8486,N_7914,N_7665);
or U8487 (N_8487,N_7257,N_7983);
or U8488 (N_8488,N_7896,N_7851);
xnor U8489 (N_8489,N_7342,N_7797);
or U8490 (N_8490,N_7115,N_7798);
or U8491 (N_8491,N_7554,N_7698);
nor U8492 (N_8492,N_7657,N_7352);
nor U8493 (N_8493,N_7620,N_7891);
nand U8494 (N_8494,N_7833,N_7174);
or U8495 (N_8495,N_7964,N_7628);
and U8496 (N_8496,N_7762,N_7627);
and U8497 (N_8497,N_7130,N_7555);
nor U8498 (N_8498,N_7222,N_7463);
nor U8499 (N_8499,N_7788,N_7454);
or U8500 (N_8500,N_7272,N_7328);
nand U8501 (N_8501,N_7996,N_7275);
nand U8502 (N_8502,N_7966,N_7433);
nor U8503 (N_8503,N_7844,N_7768);
or U8504 (N_8504,N_7116,N_7342);
and U8505 (N_8505,N_7488,N_7492);
and U8506 (N_8506,N_7445,N_7593);
nand U8507 (N_8507,N_7252,N_7230);
nor U8508 (N_8508,N_7180,N_7517);
nor U8509 (N_8509,N_7509,N_7282);
xor U8510 (N_8510,N_7212,N_7850);
or U8511 (N_8511,N_7868,N_7061);
and U8512 (N_8512,N_7049,N_7448);
nand U8513 (N_8513,N_7866,N_7847);
nor U8514 (N_8514,N_7902,N_7602);
nor U8515 (N_8515,N_7502,N_7927);
or U8516 (N_8516,N_7334,N_7817);
xnor U8517 (N_8517,N_7369,N_7400);
and U8518 (N_8518,N_7472,N_7142);
or U8519 (N_8519,N_7329,N_7531);
xnor U8520 (N_8520,N_7026,N_7492);
nand U8521 (N_8521,N_7051,N_7780);
xor U8522 (N_8522,N_7653,N_7336);
nand U8523 (N_8523,N_7891,N_7949);
and U8524 (N_8524,N_7144,N_7468);
and U8525 (N_8525,N_7960,N_7799);
xor U8526 (N_8526,N_7315,N_7318);
nand U8527 (N_8527,N_7880,N_7131);
and U8528 (N_8528,N_7607,N_7253);
nand U8529 (N_8529,N_7127,N_7565);
nand U8530 (N_8530,N_7030,N_7816);
nor U8531 (N_8531,N_7754,N_7323);
nor U8532 (N_8532,N_7917,N_7391);
nor U8533 (N_8533,N_7807,N_7226);
nor U8534 (N_8534,N_7588,N_7606);
xnor U8535 (N_8535,N_7973,N_7679);
and U8536 (N_8536,N_7129,N_7729);
nor U8537 (N_8537,N_7621,N_7814);
nand U8538 (N_8538,N_7803,N_7499);
xnor U8539 (N_8539,N_7639,N_7289);
and U8540 (N_8540,N_7359,N_7861);
or U8541 (N_8541,N_7534,N_7859);
nor U8542 (N_8542,N_7191,N_7173);
nand U8543 (N_8543,N_7823,N_7882);
and U8544 (N_8544,N_7510,N_7875);
nand U8545 (N_8545,N_7570,N_7375);
xnor U8546 (N_8546,N_7394,N_7281);
nor U8547 (N_8547,N_7405,N_7806);
nor U8548 (N_8548,N_7706,N_7626);
nor U8549 (N_8549,N_7003,N_7811);
or U8550 (N_8550,N_7401,N_7102);
nand U8551 (N_8551,N_7936,N_7442);
and U8552 (N_8552,N_7544,N_7272);
nand U8553 (N_8553,N_7892,N_7861);
or U8554 (N_8554,N_7211,N_7845);
nand U8555 (N_8555,N_7681,N_7096);
nor U8556 (N_8556,N_7578,N_7062);
and U8557 (N_8557,N_7837,N_7059);
or U8558 (N_8558,N_7449,N_7197);
or U8559 (N_8559,N_7305,N_7036);
nand U8560 (N_8560,N_7964,N_7707);
and U8561 (N_8561,N_7460,N_7061);
and U8562 (N_8562,N_7131,N_7860);
and U8563 (N_8563,N_7057,N_7949);
or U8564 (N_8564,N_7219,N_7731);
nor U8565 (N_8565,N_7790,N_7404);
nand U8566 (N_8566,N_7970,N_7287);
nand U8567 (N_8567,N_7099,N_7382);
or U8568 (N_8568,N_7334,N_7566);
or U8569 (N_8569,N_7394,N_7176);
or U8570 (N_8570,N_7947,N_7091);
xnor U8571 (N_8571,N_7576,N_7525);
nor U8572 (N_8572,N_7233,N_7881);
and U8573 (N_8573,N_7743,N_7599);
nand U8574 (N_8574,N_7641,N_7905);
xor U8575 (N_8575,N_7867,N_7594);
and U8576 (N_8576,N_7576,N_7643);
and U8577 (N_8577,N_7163,N_7515);
nor U8578 (N_8578,N_7950,N_7358);
nor U8579 (N_8579,N_7786,N_7649);
and U8580 (N_8580,N_7876,N_7794);
nand U8581 (N_8581,N_7925,N_7323);
and U8582 (N_8582,N_7034,N_7359);
xor U8583 (N_8583,N_7518,N_7396);
xor U8584 (N_8584,N_7884,N_7776);
or U8585 (N_8585,N_7490,N_7599);
nand U8586 (N_8586,N_7920,N_7487);
nand U8587 (N_8587,N_7410,N_7888);
nand U8588 (N_8588,N_7983,N_7855);
nand U8589 (N_8589,N_7939,N_7929);
xnor U8590 (N_8590,N_7753,N_7388);
or U8591 (N_8591,N_7919,N_7073);
xnor U8592 (N_8592,N_7974,N_7124);
nor U8593 (N_8593,N_7054,N_7877);
nand U8594 (N_8594,N_7444,N_7052);
xnor U8595 (N_8595,N_7145,N_7213);
or U8596 (N_8596,N_7576,N_7391);
xor U8597 (N_8597,N_7781,N_7471);
nand U8598 (N_8598,N_7233,N_7027);
nor U8599 (N_8599,N_7663,N_7023);
or U8600 (N_8600,N_7806,N_7090);
and U8601 (N_8601,N_7492,N_7720);
nand U8602 (N_8602,N_7243,N_7415);
nor U8603 (N_8603,N_7730,N_7909);
nor U8604 (N_8604,N_7243,N_7800);
and U8605 (N_8605,N_7800,N_7654);
nor U8606 (N_8606,N_7324,N_7863);
and U8607 (N_8607,N_7933,N_7940);
and U8608 (N_8608,N_7731,N_7099);
nand U8609 (N_8609,N_7499,N_7897);
or U8610 (N_8610,N_7476,N_7606);
xnor U8611 (N_8611,N_7809,N_7828);
xnor U8612 (N_8612,N_7514,N_7309);
xor U8613 (N_8613,N_7772,N_7970);
nand U8614 (N_8614,N_7388,N_7212);
or U8615 (N_8615,N_7735,N_7129);
nor U8616 (N_8616,N_7251,N_7944);
nor U8617 (N_8617,N_7784,N_7460);
xnor U8618 (N_8618,N_7537,N_7128);
nor U8619 (N_8619,N_7113,N_7933);
xnor U8620 (N_8620,N_7799,N_7769);
xnor U8621 (N_8621,N_7400,N_7515);
nor U8622 (N_8622,N_7829,N_7575);
and U8623 (N_8623,N_7950,N_7521);
nand U8624 (N_8624,N_7690,N_7740);
or U8625 (N_8625,N_7289,N_7353);
xor U8626 (N_8626,N_7871,N_7008);
nand U8627 (N_8627,N_7349,N_7366);
xor U8628 (N_8628,N_7196,N_7912);
nor U8629 (N_8629,N_7581,N_7181);
nor U8630 (N_8630,N_7487,N_7882);
xor U8631 (N_8631,N_7425,N_7102);
nor U8632 (N_8632,N_7998,N_7939);
xor U8633 (N_8633,N_7960,N_7366);
nand U8634 (N_8634,N_7526,N_7157);
nor U8635 (N_8635,N_7922,N_7709);
and U8636 (N_8636,N_7076,N_7996);
nor U8637 (N_8637,N_7906,N_7007);
or U8638 (N_8638,N_7476,N_7910);
and U8639 (N_8639,N_7223,N_7573);
or U8640 (N_8640,N_7557,N_7777);
and U8641 (N_8641,N_7743,N_7581);
xor U8642 (N_8642,N_7498,N_7868);
and U8643 (N_8643,N_7307,N_7648);
nor U8644 (N_8644,N_7146,N_7582);
xnor U8645 (N_8645,N_7736,N_7031);
and U8646 (N_8646,N_7801,N_7851);
or U8647 (N_8647,N_7149,N_7916);
nand U8648 (N_8648,N_7027,N_7246);
xnor U8649 (N_8649,N_7389,N_7390);
xor U8650 (N_8650,N_7300,N_7614);
nor U8651 (N_8651,N_7613,N_7067);
or U8652 (N_8652,N_7764,N_7674);
nor U8653 (N_8653,N_7234,N_7237);
and U8654 (N_8654,N_7226,N_7178);
nor U8655 (N_8655,N_7008,N_7077);
nor U8656 (N_8656,N_7323,N_7753);
xor U8657 (N_8657,N_7626,N_7641);
nor U8658 (N_8658,N_7663,N_7284);
and U8659 (N_8659,N_7695,N_7796);
nand U8660 (N_8660,N_7266,N_7423);
and U8661 (N_8661,N_7032,N_7396);
nand U8662 (N_8662,N_7101,N_7185);
and U8663 (N_8663,N_7360,N_7951);
nand U8664 (N_8664,N_7657,N_7110);
and U8665 (N_8665,N_7520,N_7740);
nand U8666 (N_8666,N_7328,N_7689);
and U8667 (N_8667,N_7177,N_7324);
and U8668 (N_8668,N_7990,N_7026);
and U8669 (N_8669,N_7989,N_7453);
nor U8670 (N_8670,N_7868,N_7658);
nand U8671 (N_8671,N_7547,N_7744);
or U8672 (N_8672,N_7398,N_7916);
nand U8673 (N_8673,N_7800,N_7756);
xnor U8674 (N_8674,N_7356,N_7387);
and U8675 (N_8675,N_7574,N_7450);
or U8676 (N_8676,N_7425,N_7678);
nor U8677 (N_8677,N_7958,N_7228);
nand U8678 (N_8678,N_7929,N_7746);
nand U8679 (N_8679,N_7533,N_7866);
nor U8680 (N_8680,N_7590,N_7544);
and U8681 (N_8681,N_7723,N_7745);
or U8682 (N_8682,N_7878,N_7948);
and U8683 (N_8683,N_7950,N_7502);
xor U8684 (N_8684,N_7340,N_7300);
or U8685 (N_8685,N_7704,N_7667);
nor U8686 (N_8686,N_7711,N_7453);
xor U8687 (N_8687,N_7473,N_7417);
xnor U8688 (N_8688,N_7758,N_7462);
xnor U8689 (N_8689,N_7063,N_7366);
xnor U8690 (N_8690,N_7541,N_7217);
nor U8691 (N_8691,N_7700,N_7321);
nand U8692 (N_8692,N_7142,N_7461);
nand U8693 (N_8693,N_7686,N_7883);
xnor U8694 (N_8694,N_7937,N_7070);
xor U8695 (N_8695,N_7201,N_7525);
xnor U8696 (N_8696,N_7833,N_7008);
or U8697 (N_8697,N_7035,N_7083);
and U8698 (N_8698,N_7550,N_7883);
and U8699 (N_8699,N_7557,N_7999);
and U8700 (N_8700,N_7128,N_7855);
and U8701 (N_8701,N_7658,N_7834);
and U8702 (N_8702,N_7925,N_7494);
and U8703 (N_8703,N_7031,N_7962);
or U8704 (N_8704,N_7176,N_7010);
or U8705 (N_8705,N_7098,N_7415);
nor U8706 (N_8706,N_7283,N_7666);
nand U8707 (N_8707,N_7147,N_7815);
nand U8708 (N_8708,N_7841,N_7317);
and U8709 (N_8709,N_7096,N_7952);
and U8710 (N_8710,N_7011,N_7658);
and U8711 (N_8711,N_7488,N_7917);
nand U8712 (N_8712,N_7975,N_7569);
or U8713 (N_8713,N_7072,N_7022);
xnor U8714 (N_8714,N_7619,N_7533);
and U8715 (N_8715,N_7012,N_7932);
or U8716 (N_8716,N_7465,N_7588);
xor U8717 (N_8717,N_7886,N_7676);
nor U8718 (N_8718,N_7425,N_7062);
or U8719 (N_8719,N_7415,N_7216);
nor U8720 (N_8720,N_7705,N_7749);
nor U8721 (N_8721,N_7609,N_7577);
nand U8722 (N_8722,N_7791,N_7944);
nor U8723 (N_8723,N_7458,N_7902);
nor U8724 (N_8724,N_7874,N_7956);
xnor U8725 (N_8725,N_7203,N_7962);
or U8726 (N_8726,N_7929,N_7080);
or U8727 (N_8727,N_7401,N_7855);
or U8728 (N_8728,N_7977,N_7366);
nand U8729 (N_8729,N_7094,N_7768);
nor U8730 (N_8730,N_7380,N_7563);
nand U8731 (N_8731,N_7083,N_7180);
and U8732 (N_8732,N_7491,N_7035);
xnor U8733 (N_8733,N_7186,N_7884);
or U8734 (N_8734,N_7317,N_7780);
or U8735 (N_8735,N_7052,N_7534);
or U8736 (N_8736,N_7452,N_7165);
and U8737 (N_8737,N_7701,N_7219);
xnor U8738 (N_8738,N_7284,N_7395);
or U8739 (N_8739,N_7388,N_7926);
nand U8740 (N_8740,N_7216,N_7135);
nand U8741 (N_8741,N_7846,N_7655);
or U8742 (N_8742,N_7305,N_7333);
and U8743 (N_8743,N_7145,N_7632);
or U8744 (N_8744,N_7755,N_7671);
xor U8745 (N_8745,N_7014,N_7401);
or U8746 (N_8746,N_7644,N_7106);
or U8747 (N_8747,N_7482,N_7052);
xor U8748 (N_8748,N_7513,N_7757);
nand U8749 (N_8749,N_7272,N_7300);
nand U8750 (N_8750,N_7020,N_7361);
nor U8751 (N_8751,N_7156,N_7262);
nand U8752 (N_8752,N_7171,N_7814);
xor U8753 (N_8753,N_7699,N_7424);
xor U8754 (N_8754,N_7722,N_7615);
nand U8755 (N_8755,N_7120,N_7911);
xnor U8756 (N_8756,N_7394,N_7947);
xnor U8757 (N_8757,N_7853,N_7828);
nand U8758 (N_8758,N_7140,N_7392);
and U8759 (N_8759,N_7179,N_7316);
xor U8760 (N_8760,N_7129,N_7607);
xor U8761 (N_8761,N_7608,N_7629);
nor U8762 (N_8762,N_7128,N_7293);
xnor U8763 (N_8763,N_7040,N_7167);
nor U8764 (N_8764,N_7640,N_7626);
nor U8765 (N_8765,N_7196,N_7174);
xor U8766 (N_8766,N_7520,N_7806);
and U8767 (N_8767,N_7454,N_7013);
nand U8768 (N_8768,N_7738,N_7558);
nor U8769 (N_8769,N_7406,N_7932);
or U8770 (N_8770,N_7047,N_7126);
or U8771 (N_8771,N_7886,N_7905);
and U8772 (N_8772,N_7471,N_7990);
xnor U8773 (N_8773,N_7947,N_7187);
nor U8774 (N_8774,N_7057,N_7430);
and U8775 (N_8775,N_7890,N_7388);
nor U8776 (N_8776,N_7786,N_7408);
xor U8777 (N_8777,N_7804,N_7943);
nand U8778 (N_8778,N_7049,N_7535);
or U8779 (N_8779,N_7938,N_7521);
nor U8780 (N_8780,N_7045,N_7607);
or U8781 (N_8781,N_7712,N_7911);
nand U8782 (N_8782,N_7614,N_7203);
nand U8783 (N_8783,N_7865,N_7904);
xor U8784 (N_8784,N_7345,N_7029);
and U8785 (N_8785,N_7392,N_7759);
and U8786 (N_8786,N_7035,N_7577);
or U8787 (N_8787,N_7938,N_7081);
xor U8788 (N_8788,N_7247,N_7564);
and U8789 (N_8789,N_7659,N_7312);
and U8790 (N_8790,N_7907,N_7746);
or U8791 (N_8791,N_7473,N_7440);
nand U8792 (N_8792,N_7864,N_7827);
or U8793 (N_8793,N_7908,N_7207);
nand U8794 (N_8794,N_7035,N_7967);
nand U8795 (N_8795,N_7989,N_7123);
xor U8796 (N_8796,N_7272,N_7627);
and U8797 (N_8797,N_7351,N_7577);
nand U8798 (N_8798,N_7224,N_7715);
nand U8799 (N_8799,N_7875,N_7377);
and U8800 (N_8800,N_7488,N_7541);
nor U8801 (N_8801,N_7939,N_7631);
nand U8802 (N_8802,N_7562,N_7179);
xnor U8803 (N_8803,N_7420,N_7956);
and U8804 (N_8804,N_7202,N_7837);
nand U8805 (N_8805,N_7066,N_7805);
and U8806 (N_8806,N_7975,N_7703);
and U8807 (N_8807,N_7410,N_7837);
nor U8808 (N_8808,N_7302,N_7382);
and U8809 (N_8809,N_7568,N_7442);
xor U8810 (N_8810,N_7466,N_7707);
nand U8811 (N_8811,N_7071,N_7528);
nand U8812 (N_8812,N_7483,N_7758);
or U8813 (N_8813,N_7741,N_7284);
and U8814 (N_8814,N_7767,N_7583);
and U8815 (N_8815,N_7933,N_7908);
nor U8816 (N_8816,N_7803,N_7965);
nand U8817 (N_8817,N_7094,N_7060);
and U8818 (N_8818,N_7671,N_7234);
nor U8819 (N_8819,N_7840,N_7077);
and U8820 (N_8820,N_7683,N_7534);
xnor U8821 (N_8821,N_7693,N_7497);
nand U8822 (N_8822,N_7164,N_7707);
xnor U8823 (N_8823,N_7069,N_7158);
or U8824 (N_8824,N_7112,N_7707);
or U8825 (N_8825,N_7573,N_7347);
and U8826 (N_8826,N_7375,N_7838);
xor U8827 (N_8827,N_7350,N_7258);
nand U8828 (N_8828,N_7164,N_7402);
nand U8829 (N_8829,N_7355,N_7716);
and U8830 (N_8830,N_7896,N_7592);
nand U8831 (N_8831,N_7621,N_7608);
and U8832 (N_8832,N_7273,N_7594);
xor U8833 (N_8833,N_7583,N_7315);
xor U8834 (N_8834,N_7930,N_7236);
and U8835 (N_8835,N_7935,N_7906);
nor U8836 (N_8836,N_7444,N_7645);
nand U8837 (N_8837,N_7743,N_7406);
nor U8838 (N_8838,N_7082,N_7111);
or U8839 (N_8839,N_7283,N_7765);
and U8840 (N_8840,N_7147,N_7355);
and U8841 (N_8841,N_7142,N_7606);
xor U8842 (N_8842,N_7895,N_7402);
nand U8843 (N_8843,N_7644,N_7002);
nand U8844 (N_8844,N_7706,N_7232);
xnor U8845 (N_8845,N_7074,N_7599);
xnor U8846 (N_8846,N_7199,N_7127);
or U8847 (N_8847,N_7704,N_7026);
or U8848 (N_8848,N_7053,N_7364);
or U8849 (N_8849,N_7960,N_7333);
nor U8850 (N_8850,N_7067,N_7458);
and U8851 (N_8851,N_7814,N_7081);
nor U8852 (N_8852,N_7160,N_7728);
and U8853 (N_8853,N_7436,N_7195);
and U8854 (N_8854,N_7087,N_7720);
or U8855 (N_8855,N_7584,N_7466);
xor U8856 (N_8856,N_7673,N_7395);
and U8857 (N_8857,N_7992,N_7593);
nor U8858 (N_8858,N_7664,N_7953);
or U8859 (N_8859,N_7162,N_7887);
or U8860 (N_8860,N_7131,N_7258);
nor U8861 (N_8861,N_7101,N_7754);
nor U8862 (N_8862,N_7746,N_7314);
or U8863 (N_8863,N_7300,N_7735);
nand U8864 (N_8864,N_7972,N_7524);
and U8865 (N_8865,N_7612,N_7361);
xnor U8866 (N_8866,N_7416,N_7336);
nor U8867 (N_8867,N_7447,N_7693);
or U8868 (N_8868,N_7155,N_7724);
or U8869 (N_8869,N_7501,N_7100);
nor U8870 (N_8870,N_7151,N_7307);
nor U8871 (N_8871,N_7631,N_7039);
xnor U8872 (N_8872,N_7472,N_7581);
and U8873 (N_8873,N_7267,N_7228);
xnor U8874 (N_8874,N_7191,N_7682);
nand U8875 (N_8875,N_7871,N_7633);
nand U8876 (N_8876,N_7556,N_7317);
nor U8877 (N_8877,N_7741,N_7509);
or U8878 (N_8878,N_7320,N_7638);
xnor U8879 (N_8879,N_7033,N_7301);
or U8880 (N_8880,N_7970,N_7410);
xor U8881 (N_8881,N_7097,N_7219);
or U8882 (N_8882,N_7166,N_7163);
and U8883 (N_8883,N_7086,N_7812);
nor U8884 (N_8884,N_7562,N_7928);
xor U8885 (N_8885,N_7990,N_7724);
or U8886 (N_8886,N_7276,N_7142);
nand U8887 (N_8887,N_7443,N_7412);
xnor U8888 (N_8888,N_7742,N_7074);
xor U8889 (N_8889,N_7286,N_7754);
or U8890 (N_8890,N_7555,N_7855);
or U8891 (N_8891,N_7417,N_7499);
nand U8892 (N_8892,N_7769,N_7831);
and U8893 (N_8893,N_7141,N_7697);
or U8894 (N_8894,N_7758,N_7684);
nor U8895 (N_8895,N_7998,N_7632);
nand U8896 (N_8896,N_7659,N_7825);
nor U8897 (N_8897,N_7482,N_7760);
xor U8898 (N_8898,N_7033,N_7981);
nand U8899 (N_8899,N_7252,N_7480);
and U8900 (N_8900,N_7473,N_7088);
nor U8901 (N_8901,N_7400,N_7656);
or U8902 (N_8902,N_7735,N_7965);
xor U8903 (N_8903,N_7475,N_7942);
nand U8904 (N_8904,N_7727,N_7796);
nor U8905 (N_8905,N_7614,N_7741);
xor U8906 (N_8906,N_7771,N_7411);
nand U8907 (N_8907,N_7802,N_7488);
and U8908 (N_8908,N_7544,N_7191);
xor U8909 (N_8909,N_7786,N_7431);
and U8910 (N_8910,N_7428,N_7164);
or U8911 (N_8911,N_7073,N_7177);
xor U8912 (N_8912,N_7101,N_7896);
or U8913 (N_8913,N_7522,N_7040);
or U8914 (N_8914,N_7733,N_7637);
nand U8915 (N_8915,N_7950,N_7568);
nand U8916 (N_8916,N_7333,N_7489);
or U8917 (N_8917,N_7414,N_7487);
nand U8918 (N_8918,N_7568,N_7588);
nand U8919 (N_8919,N_7912,N_7408);
and U8920 (N_8920,N_7833,N_7135);
nor U8921 (N_8921,N_7370,N_7318);
and U8922 (N_8922,N_7997,N_7943);
or U8923 (N_8923,N_7318,N_7092);
or U8924 (N_8924,N_7197,N_7117);
nand U8925 (N_8925,N_7223,N_7177);
xor U8926 (N_8926,N_7492,N_7990);
or U8927 (N_8927,N_7931,N_7254);
or U8928 (N_8928,N_7944,N_7542);
xnor U8929 (N_8929,N_7510,N_7929);
xor U8930 (N_8930,N_7440,N_7198);
nand U8931 (N_8931,N_7235,N_7422);
xnor U8932 (N_8932,N_7439,N_7472);
nand U8933 (N_8933,N_7082,N_7581);
or U8934 (N_8934,N_7258,N_7569);
xor U8935 (N_8935,N_7554,N_7751);
nor U8936 (N_8936,N_7983,N_7600);
or U8937 (N_8937,N_7915,N_7011);
nor U8938 (N_8938,N_7123,N_7779);
nor U8939 (N_8939,N_7524,N_7648);
nand U8940 (N_8940,N_7455,N_7835);
xnor U8941 (N_8941,N_7753,N_7688);
or U8942 (N_8942,N_7224,N_7770);
and U8943 (N_8943,N_7810,N_7564);
xnor U8944 (N_8944,N_7861,N_7214);
nand U8945 (N_8945,N_7681,N_7176);
xor U8946 (N_8946,N_7530,N_7078);
or U8947 (N_8947,N_7700,N_7415);
and U8948 (N_8948,N_7594,N_7070);
nand U8949 (N_8949,N_7523,N_7335);
xor U8950 (N_8950,N_7715,N_7461);
xor U8951 (N_8951,N_7544,N_7038);
or U8952 (N_8952,N_7294,N_7658);
nor U8953 (N_8953,N_7594,N_7882);
or U8954 (N_8954,N_7839,N_7532);
xor U8955 (N_8955,N_7012,N_7523);
nor U8956 (N_8956,N_7518,N_7596);
and U8957 (N_8957,N_7442,N_7903);
xnor U8958 (N_8958,N_7247,N_7194);
or U8959 (N_8959,N_7046,N_7325);
and U8960 (N_8960,N_7964,N_7740);
xnor U8961 (N_8961,N_7384,N_7670);
and U8962 (N_8962,N_7771,N_7988);
xor U8963 (N_8963,N_7793,N_7566);
xnor U8964 (N_8964,N_7496,N_7360);
xnor U8965 (N_8965,N_7884,N_7139);
xor U8966 (N_8966,N_7167,N_7456);
nor U8967 (N_8967,N_7013,N_7262);
xnor U8968 (N_8968,N_7279,N_7514);
nand U8969 (N_8969,N_7654,N_7557);
nor U8970 (N_8970,N_7288,N_7758);
nor U8971 (N_8971,N_7892,N_7547);
and U8972 (N_8972,N_7672,N_7090);
and U8973 (N_8973,N_7291,N_7742);
nor U8974 (N_8974,N_7016,N_7861);
nand U8975 (N_8975,N_7961,N_7685);
xnor U8976 (N_8976,N_7607,N_7651);
and U8977 (N_8977,N_7543,N_7383);
and U8978 (N_8978,N_7388,N_7818);
or U8979 (N_8979,N_7643,N_7120);
xnor U8980 (N_8980,N_7658,N_7515);
or U8981 (N_8981,N_7673,N_7108);
xnor U8982 (N_8982,N_7721,N_7038);
nand U8983 (N_8983,N_7152,N_7205);
and U8984 (N_8984,N_7723,N_7643);
and U8985 (N_8985,N_7335,N_7403);
nor U8986 (N_8986,N_7060,N_7966);
or U8987 (N_8987,N_7003,N_7573);
nor U8988 (N_8988,N_7277,N_7742);
and U8989 (N_8989,N_7495,N_7948);
or U8990 (N_8990,N_7092,N_7753);
xnor U8991 (N_8991,N_7476,N_7953);
xnor U8992 (N_8992,N_7534,N_7145);
nand U8993 (N_8993,N_7887,N_7827);
xnor U8994 (N_8994,N_7762,N_7193);
nor U8995 (N_8995,N_7406,N_7023);
nand U8996 (N_8996,N_7490,N_7638);
nor U8997 (N_8997,N_7872,N_7277);
nor U8998 (N_8998,N_7611,N_7390);
xor U8999 (N_8999,N_7294,N_7708);
and U9000 (N_9000,N_8802,N_8361);
xor U9001 (N_9001,N_8984,N_8735);
and U9002 (N_9002,N_8487,N_8759);
nand U9003 (N_9003,N_8946,N_8769);
nor U9004 (N_9004,N_8756,N_8336);
and U9005 (N_9005,N_8872,N_8883);
and U9006 (N_9006,N_8637,N_8874);
nand U9007 (N_9007,N_8933,N_8028);
or U9008 (N_9008,N_8180,N_8232);
nand U9009 (N_9009,N_8674,N_8750);
nand U9010 (N_9010,N_8424,N_8118);
nor U9011 (N_9011,N_8431,N_8638);
nor U9012 (N_9012,N_8112,N_8788);
or U9013 (N_9013,N_8468,N_8244);
xor U9014 (N_9014,N_8999,N_8319);
nor U9015 (N_9015,N_8557,N_8757);
and U9016 (N_9016,N_8950,N_8728);
and U9017 (N_9017,N_8850,N_8388);
or U9018 (N_9018,N_8768,N_8264);
xor U9019 (N_9019,N_8496,N_8177);
or U9020 (N_9020,N_8383,N_8574);
or U9021 (N_9021,N_8558,N_8868);
nor U9022 (N_9022,N_8831,N_8543);
or U9023 (N_9023,N_8240,N_8733);
xor U9024 (N_9024,N_8657,N_8707);
nor U9025 (N_9025,N_8708,N_8943);
and U9026 (N_9026,N_8207,N_8806);
nand U9027 (N_9027,N_8616,N_8605);
nand U9028 (N_9028,N_8562,N_8696);
xnor U9029 (N_9029,N_8408,N_8513);
or U9030 (N_9030,N_8398,N_8776);
or U9031 (N_9031,N_8393,N_8853);
and U9032 (N_9032,N_8667,N_8871);
nor U9033 (N_9033,N_8335,N_8681);
or U9034 (N_9034,N_8370,N_8991);
or U9035 (N_9035,N_8678,N_8745);
xor U9036 (N_9036,N_8985,N_8120);
nor U9037 (N_9037,N_8130,N_8194);
and U9038 (N_9038,N_8613,N_8066);
xor U9039 (N_9039,N_8978,N_8881);
or U9040 (N_9040,N_8820,N_8770);
and U9041 (N_9041,N_8552,N_8643);
xnor U9042 (N_9042,N_8173,N_8209);
nand U9043 (N_9043,N_8348,N_8719);
and U9044 (N_9044,N_8892,N_8094);
or U9045 (N_9045,N_8687,N_8111);
nor U9046 (N_9046,N_8146,N_8550);
nor U9047 (N_9047,N_8504,N_8332);
and U9048 (N_9048,N_8941,N_8294);
xnor U9049 (N_9049,N_8845,N_8299);
or U9050 (N_9050,N_8683,N_8144);
nor U9051 (N_9051,N_8127,N_8694);
or U9052 (N_9052,N_8572,N_8304);
or U9053 (N_9053,N_8726,N_8239);
or U9054 (N_9054,N_8055,N_8908);
nor U9055 (N_9055,N_8080,N_8163);
xor U9056 (N_9056,N_8639,N_8885);
or U9057 (N_9057,N_8379,N_8900);
nor U9058 (N_9058,N_8607,N_8901);
nand U9059 (N_9059,N_8053,N_8219);
nand U9060 (N_9060,N_8857,N_8436);
nor U9061 (N_9061,N_8193,N_8469);
and U9062 (N_9062,N_8480,N_8316);
or U9063 (N_9063,N_8349,N_8861);
and U9064 (N_9064,N_8352,N_8089);
and U9065 (N_9065,N_8916,N_8084);
nand U9066 (N_9066,N_8189,N_8256);
nand U9067 (N_9067,N_8277,N_8226);
or U9068 (N_9068,N_8037,N_8748);
nand U9069 (N_9069,N_8249,N_8477);
nand U9070 (N_9070,N_8346,N_8016);
or U9071 (N_9071,N_8470,N_8508);
nor U9072 (N_9072,N_8217,N_8679);
xnor U9073 (N_9073,N_8401,N_8576);
nand U9074 (N_9074,N_8526,N_8751);
xor U9075 (N_9075,N_8188,N_8444);
xnor U9076 (N_9076,N_8325,N_8419);
and U9077 (N_9077,N_8568,N_8823);
or U9078 (N_9078,N_8835,N_8108);
and U9079 (N_9079,N_8965,N_8204);
nand U9080 (N_9080,N_8791,N_8131);
and U9081 (N_9081,N_8921,N_8430);
nand U9082 (N_9082,N_8169,N_8721);
and U9083 (N_9083,N_8418,N_8877);
xnor U9084 (N_9084,N_8960,N_8390);
and U9085 (N_9085,N_8475,N_8454);
nand U9086 (N_9086,N_8251,N_8537);
or U9087 (N_9087,N_8712,N_8389);
nand U9088 (N_9088,N_8994,N_8830);
or U9089 (N_9089,N_8502,N_8732);
and U9090 (N_9090,N_8031,N_8579);
nor U9091 (N_9091,N_8865,N_8590);
and U9092 (N_9092,N_8715,N_8794);
or U9093 (N_9093,N_8971,N_8743);
nor U9094 (N_9094,N_8340,N_8573);
and U9095 (N_9095,N_8455,N_8292);
nand U9096 (N_9096,N_8754,N_8840);
or U9097 (N_9097,N_8822,N_8278);
nor U9098 (N_9098,N_8186,N_8979);
or U9099 (N_9099,N_8701,N_8964);
or U9100 (N_9100,N_8624,N_8859);
nand U9101 (N_9101,N_8191,N_8096);
nor U9102 (N_9102,N_8334,N_8364);
nor U9103 (N_9103,N_8143,N_8821);
nor U9104 (N_9104,N_8341,N_8261);
nor U9105 (N_9105,N_8847,N_8618);
and U9106 (N_9106,N_8106,N_8435);
and U9107 (N_9107,N_8365,N_8101);
xnor U9108 (N_9108,N_8631,N_8026);
nand U9109 (N_9109,N_8040,N_8529);
nand U9110 (N_9110,N_8531,N_8641);
or U9111 (N_9111,N_8786,N_8535);
and U9112 (N_9112,N_8539,N_8609);
xnor U9113 (N_9113,N_8784,N_8382);
nand U9114 (N_9114,N_8368,N_8825);
nor U9115 (N_9115,N_8816,N_8671);
or U9116 (N_9116,N_8875,N_8676);
and U9117 (N_9117,N_8035,N_8648);
or U9118 (N_9118,N_8595,N_8119);
and U9119 (N_9119,N_8934,N_8981);
and U9120 (N_9120,N_8048,N_8175);
nand U9121 (N_9121,N_8940,N_8915);
nor U9122 (N_9122,N_8109,N_8566);
nand U9123 (N_9123,N_8996,N_8328);
nand U9124 (N_9124,N_8499,N_8371);
and U9125 (N_9125,N_8922,N_8795);
and U9126 (N_9126,N_8744,N_8355);
nand U9127 (N_9127,N_8133,N_8484);
and U9128 (N_9128,N_8359,N_8377);
nor U9129 (N_9129,N_8503,N_8839);
nand U9130 (N_9130,N_8530,N_8547);
nor U9131 (N_9131,N_8524,N_8866);
or U9132 (N_9132,N_8034,N_8409);
or U9133 (N_9133,N_8826,N_8338);
or U9134 (N_9134,N_8212,N_8561);
xnor U9135 (N_9135,N_8760,N_8001);
nand U9136 (N_9136,N_8461,N_8152);
nand U9137 (N_9137,N_8944,N_8556);
or U9138 (N_9138,N_8620,N_8955);
xnor U9139 (N_9139,N_8017,N_8974);
nor U9140 (N_9140,N_8421,N_8310);
nor U9141 (N_9141,N_8460,N_8688);
nand U9142 (N_9142,N_8538,N_8913);
xnor U9143 (N_9143,N_8453,N_8402);
and U9144 (N_9144,N_8353,N_8227);
nand U9145 (N_9145,N_8771,N_8661);
or U9146 (N_9146,N_8646,N_8870);
and U9147 (N_9147,N_8911,N_8773);
xnor U9148 (N_9148,N_8014,N_8296);
xor U9149 (N_9149,N_8059,N_8774);
and U9150 (N_9150,N_8086,N_8967);
xnor U9151 (N_9151,N_8030,N_8029);
nor U9152 (N_9152,N_8002,N_8636);
nand U9153 (N_9153,N_8121,N_8909);
xor U9154 (N_9154,N_8819,N_8196);
and U9155 (N_9155,N_8890,N_8758);
or U9156 (N_9156,N_8652,N_8672);
nand U9157 (N_9157,N_8815,N_8238);
xnor U9158 (N_9158,N_8100,N_8019);
or U9159 (N_9159,N_8559,N_8314);
nor U9160 (N_9160,N_8237,N_8789);
or U9161 (N_9161,N_8333,N_8125);
xor U9162 (N_9162,N_8880,N_8507);
nand U9163 (N_9163,N_8357,N_8489);
xnor U9164 (N_9164,N_8128,N_8302);
xor U9165 (N_9165,N_8159,N_8710);
xnor U9166 (N_9166,N_8437,N_8044);
or U9167 (N_9167,N_8473,N_8841);
nor U9168 (N_9168,N_8665,N_8907);
nand U9169 (N_9169,N_8234,N_8536);
and U9170 (N_9170,N_8447,N_8288);
and U9171 (N_9171,N_8271,N_8324);
nand U9172 (N_9172,N_8814,N_8218);
and U9173 (N_9173,N_8367,N_8187);
nand U9174 (N_9174,N_8592,N_8117);
nor U9175 (N_9175,N_8472,N_8465);
nor U9176 (N_9176,N_8351,N_8702);
nand U9177 (N_9177,N_8575,N_8910);
or U9178 (N_9178,N_8033,N_8363);
xor U9179 (N_9179,N_8765,N_8762);
or U9180 (N_9180,N_8399,N_8129);
xnor U9181 (N_9181,N_8628,N_8013);
xnor U9182 (N_9182,N_8932,N_8553);
xnor U9183 (N_9183,N_8380,N_8356);
and U9184 (N_9184,N_8600,N_8659);
nor U9185 (N_9185,N_8809,N_8429);
and U9186 (N_9186,N_8801,N_8634);
nor U9187 (N_9187,N_8254,N_8483);
nor U9188 (N_9188,N_8474,N_8148);
and U9189 (N_9189,N_8606,N_8366);
nor U9190 (N_9190,N_8653,N_8602);
xnor U9191 (N_9191,N_8852,N_8441);
or U9192 (N_9192,N_8291,N_8884);
nand U9193 (N_9193,N_8904,N_8627);
nor U9194 (N_9194,N_8842,N_8279);
xnor U9195 (N_9195,N_8230,N_8918);
nand U9196 (N_9196,N_8591,N_8114);
nand U9197 (N_9197,N_8986,N_8467);
and U9198 (N_9198,N_8283,N_8988);
xor U9199 (N_9199,N_8838,N_8038);
nor U9200 (N_9200,N_8403,N_8738);
xor U9201 (N_9201,N_8775,N_8197);
nand U9202 (N_9202,N_8095,N_8581);
xnor U9203 (N_9203,N_8413,N_8949);
nor U9204 (N_9204,N_8376,N_8032);
nor U9205 (N_9205,N_8381,N_8587);
or U9206 (N_9206,N_8580,N_8521);
xor U9207 (N_9207,N_8200,N_8072);
and U9208 (N_9208,N_8995,N_8110);
nand U9209 (N_9209,N_8596,N_8983);
or U9210 (N_9210,N_8360,N_8003);
xor U9211 (N_9211,N_8577,N_8315);
nor U9212 (N_9212,N_8598,N_8860);
and U9213 (N_9213,N_8276,N_8534);
and U9214 (N_9214,N_8009,N_8584);
nor U9215 (N_9215,N_8190,N_8493);
xor U9216 (N_9216,N_8632,N_8384);
xnor U9217 (N_9217,N_8061,N_8451);
nand U9218 (N_9218,N_8166,N_8582);
and U9219 (N_9219,N_8064,N_8690);
or U9220 (N_9220,N_8843,N_8655);
or U9221 (N_9221,N_8548,N_8938);
nor U9222 (N_9222,N_8532,N_8666);
nand U9223 (N_9223,N_8057,N_8533);
xor U9224 (N_9224,N_8992,N_8067);
xnor U9225 (N_9225,N_8153,N_8394);
or U9226 (N_9226,N_8284,N_8780);
and U9227 (N_9227,N_8783,N_8720);
nor U9228 (N_9228,N_8697,N_8515);
nand U9229 (N_9229,N_8982,N_8873);
nor U9230 (N_9230,N_8422,N_8350);
nor U9231 (N_9231,N_8972,N_8115);
xor U9232 (N_9232,N_8252,N_8790);
or U9233 (N_9233,N_8851,N_8452);
xor U9234 (N_9234,N_8083,N_8043);
nand U9235 (N_9235,N_8746,N_8192);
and U9236 (N_9236,N_8862,N_8245);
and U9237 (N_9237,N_8198,N_8893);
nand U9238 (N_9238,N_8736,N_8387);
xnor U9239 (N_9239,N_8263,N_8203);
nor U9240 (N_9240,N_8936,N_8662);
or U9241 (N_9241,N_8416,N_8510);
nor U9242 (N_9242,N_8306,N_8076);
nand U9243 (N_9243,N_8682,N_8717);
nor U9244 (N_9244,N_8772,N_8796);
nand U9245 (N_9245,N_8425,N_8020);
nor U9246 (N_9246,N_8729,N_8063);
or U9247 (N_9247,N_8397,N_8528);
or U9248 (N_9248,N_8544,N_8924);
or U9249 (N_9249,N_8225,N_8597);
xor U9250 (N_9250,N_8275,N_8695);
nor U9251 (N_9251,N_8691,N_8085);
xor U9252 (N_9252,N_8763,N_8675);
nor U9253 (N_9253,N_8899,N_8301);
or U9254 (N_9254,N_8698,N_8411);
nor U9255 (N_9255,N_8412,N_8062);
nand U9256 (N_9256,N_8099,N_8311);
or U9257 (N_9257,N_8255,N_8185);
and U9258 (N_9258,N_8793,N_8650);
and U9259 (N_9259,N_8036,N_8052);
nand U9260 (N_9260,N_8817,N_8626);
nor U9261 (N_9261,N_8073,N_8214);
xnor U9262 (N_9262,N_8041,N_8642);
nand U9263 (N_9263,N_8813,N_8798);
and U9264 (N_9264,N_8405,N_8079);
nand U9265 (N_9265,N_8848,N_8199);
nor U9266 (N_9266,N_8093,N_8273);
xor U9267 (N_9267,N_8829,N_8959);
nor U9268 (N_9268,N_8337,N_8082);
nor U9269 (N_9269,N_8764,N_8268);
xnor U9270 (N_9270,N_8307,N_8170);
or U9271 (N_9271,N_8540,N_8007);
nor U9272 (N_9272,N_8787,N_8260);
nand U9273 (N_9273,N_8141,N_8242);
nand U9274 (N_9274,N_8722,N_8071);
xnor U9275 (N_9275,N_8375,N_8113);
nor U9276 (N_9276,N_8298,N_8223);
nand U9277 (N_9277,N_8329,N_8878);
nand U9278 (N_9278,N_8523,N_8545);
xor U9279 (N_9279,N_8272,N_8585);
nand U9280 (N_9280,N_8138,N_8280);
xnor U9281 (N_9281,N_8699,N_8948);
nor U9282 (N_9282,N_8505,N_8179);
xor U9283 (N_9283,N_8903,N_8888);
xor U9284 (N_9284,N_8541,N_8312);
xnor U9285 (N_9285,N_8195,N_8427);
or U9286 (N_9286,N_8737,N_8990);
nor U9287 (N_9287,N_8491,N_8520);
nand U9288 (N_9288,N_8182,N_8977);
and U9289 (N_9289,N_8202,N_8231);
nor U9290 (N_9290,N_8236,N_8420);
or U9291 (N_9291,N_8457,N_8395);
nand U9292 (N_9292,N_8181,N_8518);
or U9293 (N_9293,N_8511,N_8739);
and U9294 (N_9294,N_8134,N_8228);
or U9295 (N_9295,N_8810,N_8449);
nand U9296 (N_9296,N_8747,N_8807);
and U9297 (N_9297,N_8176,N_8406);
or U9298 (N_9298,N_8116,N_8285);
nor U9299 (N_9299,N_8047,N_8889);
and U9300 (N_9300,N_8253,N_8303);
nor U9301 (N_9301,N_8160,N_8614);
nand U9302 (N_9302,N_8439,N_8318);
or U9303 (N_9303,N_8132,N_8785);
nand U9304 (N_9304,N_8091,N_8976);
nor U9305 (N_9305,N_8258,N_8246);
nor U9306 (N_9306,N_8782,N_8863);
nor U9307 (N_9307,N_8858,N_8824);
nor U9308 (N_9308,N_8599,N_8068);
xnor U9309 (N_9309,N_8834,N_8867);
or U9310 (N_9310,N_8660,N_8725);
nand U9311 (N_9311,N_8570,N_8956);
nand U9312 (N_9312,N_8601,N_8257);
xor U9313 (N_9313,N_8897,N_8633);
or U9314 (N_9314,N_8827,N_8087);
and U9315 (N_9315,N_8400,N_8049);
and U9316 (N_9316,N_8206,N_8516);
and U9317 (N_9317,N_8459,N_8700);
or U9318 (N_9318,N_8321,N_8896);
xor U9319 (N_9319,N_8828,N_8248);
or U9320 (N_9320,N_8250,N_8446);
nand U9321 (N_9321,N_8649,N_8931);
nor U9322 (N_9322,N_8481,N_8781);
and U9323 (N_9323,N_8215,N_8339);
nor U9324 (N_9324,N_8313,N_8644);
nor U9325 (N_9325,N_8928,N_8706);
xor U9326 (N_9326,N_8869,N_8989);
and U9327 (N_9327,N_8973,N_8752);
nor U9328 (N_9328,N_8432,N_8755);
and U9329 (N_9329,N_8165,N_8058);
nor U9330 (N_9330,N_8617,N_8077);
nand U9331 (N_9331,N_8957,N_8282);
xor U9332 (N_9332,N_8372,N_8070);
nand U9333 (N_9333,N_8808,N_8391);
and U9334 (N_9334,N_8952,N_8517);
xnor U9335 (N_9335,N_8849,N_8963);
or U9336 (N_9336,N_8894,N_8069);
xor U9337 (N_9337,N_8433,N_8966);
nor U9338 (N_9338,N_8902,N_8525);
or U9339 (N_9339,N_8689,N_8056);
nand U9340 (N_9340,N_8104,N_8097);
xor U9341 (N_9341,N_8078,N_8274);
and U9342 (N_9342,N_8221,N_8293);
and U9343 (N_9343,N_8220,N_8494);
or U9344 (N_9344,N_8423,N_8000);
or U9345 (N_9345,N_8488,N_8320);
and U9346 (N_9346,N_8622,N_8135);
xnor U9347 (N_9347,N_8456,N_8050);
xnor U9348 (N_9348,N_8156,N_8373);
nand U9349 (N_9349,N_8927,N_8322);
nand U9350 (N_9350,N_8962,N_8448);
and U9351 (N_9351,N_8407,N_8554);
nor U9352 (N_9352,N_8442,N_8656);
nand U9353 (N_9353,N_8107,N_8286);
and U9354 (N_9354,N_8065,N_8331);
nor U9355 (N_9355,N_8330,N_8347);
xor U9356 (N_9356,N_8136,N_8327);
and U9357 (N_9357,N_8492,N_8137);
and U9358 (N_9358,N_8777,N_8567);
nand U9359 (N_9359,N_8914,N_8951);
xnor U9360 (N_9360,N_8919,N_8417);
nand U9361 (N_9361,N_8608,N_8023);
nand U9362 (N_9362,N_8478,N_8629);
and U9363 (N_9363,N_8718,N_8024);
nor U9364 (N_9364,N_8953,N_8445);
xor U9365 (N_9365,N_8742,N_8741);
nand U9366 (N_9366,N_8610,N_8415);
nand U9367 (N_9367,N_8895,N_8920);
xnor U9368 (N_9368,N_8876,N_8693);
or U9369 (N_9369,N_8571,N_8458);
and U9370 (N_9370,N_8929,N_8930);
or U9371 (N_9371,N_8386,N_8837);
xnor U9372 (N_9372,N_8168,N_8640);
xor U9373 (N_9373,N_8542,N_8619);
xor U9374 (N_9374,N_8027,N_8968);
nand U9375 (N_9375,N_8912,N_8476);
nor U9376 (N_9376,N_8854,N_8022);
nand U9377 (N_9377,N_8519,N_8612);
nor U9378 (N_9378,N_8647,N_8124);
nor U9379 (N_9379,N_8229,N_8378);
and U9380 (N_9380,N_8512,N_8692);
xnor U9381 (N_9381,N_8213,N_8224);
and U9382 (N_9382,N_8281,N_8266);
nor U9383 (N_9383,N_8404,N_8471);
xnor U9384 (N_9384,N_8727,N_8805);
or U9385 (N_9385,N_8522,N_8343);
or U9386 (N_9386,N_8551,N_8958);
nor U9387 (N_9387,N_8856,N_8147);
or U9388 (N_9388,N_8724,N_8184);
or U9389 (N_9389,N_8506,N_8150);
or U9390 (N_9390,N_8354,N_8882);
or U9391 (N_9391,N_8997,N_8440);
xnor U9392 (N_9392,N_8560,N_8730);
nand U9393 (N_9393,N_8317,N_8879);
and U9394 (N_9394,N_8906,N_8045);
or U9395 (N_9395,N_8300,N_8074);
and U9396 (N_9396,N_8886,N_8374);
nor U9397 (N_9397,N_8345,N_8438);
nand U9398 (N_9398,N_8797,N_8954);
nand U9399 (N_9399,N_8167,N_8549);
xor U9400 (N_9400,N_8993,N_8804);
and U9401 (N_9401,N_8164,N_8669);
xnor U9402 (N_9402,N_8490,N_8021);
xnor U9403 (N_9403,N_8767,N_8222);
nand U9404 (N_9404,N_8090,N_8015);
xor U9405 (N_9405,N_8102,N_8937);
and U9406 (N_9406,N_8723,N_8385);
and U9407 (N_9407,N_8625,N_8241);
xor U9408 (N_9408,N_8362,N_8259);
or U9409 (N_9409,N_8555,N_8235);
or U9410 (N_9410,N_8970,N_8426);
xnor U9411 (N_9411,N_8686,N_8621);
or U9412 (N_9412,N_8586,N_8799);
and U9413 (N_9413,N_8713,N_8514);
or U9414 (N_9414,N_8466,N_8939);
xnor U9415 (N_9415,N_8267,N_8887);
xor U9416 (N_9416,N_8800,N_8155);
nand U9417 (N_9417,N_8142,N_8092);
xnor U9418 (N_9418,N_8060,N_8703);
nand U9419 (N_9419,N_8042,N_8926);
xnor U9420 (N_9420,N_8326,N_8891);
xnor U9421 (N_9421,N_8500,N_8923);
or U9422 (N_9422,N_8677,N_8980);
or U9423 (N_9423,N_8172,N_8105);
nand U9424 (N_9424,N_8479,N_8969);
nor U9425 (N_9425,N_8846,N_8711);
xor U9426 (N_9426,N_8668,N_8342);
nor U9427 (N_9427,N_8247,N_8369);
nor U9428 (N_9428,N_8812,N_8075);
nand U9429 (N_9429,N_8987,N_8495);
nand U9430 (N_9430,N_8122,N_8464);
xnor U9431 (N_9431,N_8593,N_8947);
xor U9432 (N_9432,N_8008,N_8766);
nor U9433 (N_9433,N_8563,N_8265);
xor U9434 (N_9434,N_8588,N_8012);
or U9435 (N_9435,N_8216,N_8323);
nand U9436 (N_9436,N_8709,N_8836);
or U9437 (N_9437,N_8578,N_8233);
nand U9438 (N_9438,N_8546,N_8081);
xor U9439 (N_9439,N_8714,N_8208);
nand U9440 (N_9440,N_8039,N_8818);
and U9441 (N_9441,N_8149,N_8139);
and U9442 (N_9442,N_8615,N_8174);
nand U9443 (N_9443,N_8803,N_8779);
xor U9444 (N_9444,N_8685,N_8157);
or U9445 (N_9445,N_8344,N_8740);
nor U9446 (N_9446,N_8509,N_8054);
xor U9447 (N_9447,N_8396,N_8565);
or U9448 (N_9448,N_8716,N_8098);
nand U9449 (N_9449,N_8583,N_8654);
xnor U9450 (N_9450,N_8358,N_8410);
nor U9451 (N_9451,N_8010,N_8151);
and U9452 (N_9452,N_8486,N_8734);
or U9453 (N_9453,N_8428,N_8673);
nor U9454 (N_9454,N_8482,N_8603);
nand U9455 (N_9455,N_8501,N_8864);
or U9456 (N_9456,N_8898,N_8935);
xor U9457 (N_9457,N_8158,N_8705);
and U9458 (N_9458,N_8004,N_8414);
nand U9459 (N_9459,N_8145,N_8623);
nand U9460 (N_9460,N_8210,N_8018);
xor U9461 (N_9461,N_8704,N_8498);
nor U9462 (N_9462,N_8297,N_8998);
xnor U9463 (N_9463,N_8778,N_8961);
nand U9464 (N_9464,N_8611,N_8564);
and U9465 (N_9465,N_8604,N_8046);
nand U9466 (N_9466,N_8462,N_8211);
nor U9467 (N_9467,N_8243,N_8308);
nand U9468 (N_9468,N_8025,N_8450);
xnor U9469 (N_9469,N_8589,N_8855);
xnor U9470 (N_9470,N_8753,N_8645);
nand U9471 (N_9471,N_8975,N_8205);
nand U9472 (N_9472,N_8269,N_8103);
or U9473 (N_9473,N_8463,N_8663);
or U9474 (N_9474,N_8680,N_8792);
or U9475 (N_9475,N_8171,N_8749);
nor U9476 (N_9476,N_8183,N_8658);
nand U9477 (N_9477,N_8295,N_8917);
xor U9478 (N_9478,N_8811,N_8443);
or U9479 (N_9479,N_8392,N_8527);
nor U9480 (N_9480,N_8630,N_8844);
or U9481 (N_9481,N_8005,N_8178);
nand U9482 (N_9482,N_8497,N_8088);
xor U9483 (N_9483,N_8289,N_8434);
or U9484 (N_9484,N_8651,N_8011);
or U9485 (N_9485,N_8569,N_8201);
xnor U9486 (N_9486,N_8162,N_8161);
or U9487 (N_9487,N_8635,N_8664);
or U9488 (N_9488,N_8485,N_8126);
nor U9489 (N_9489,N_8670,N_8140);
nor U9490 (N_9490,N_8684,N_8262);
nor U9491 (N_9491,N_8942,N_8309);
nand U9492 (N_9492,N_8287,N_8270);
nand U9493 (N_9493,N_8154,N_8761);
xor U9494 (N_9494,N_8905,N_8051);
xnor U9495 (N_9495,N_8925,N_8832);
xnor U9496 (N_9496,N_8305,N_8123);
nor U9497 (N_9497,N_8290,N_8731);
nand U9498 (N_9498,N_8945,N_8006);
or U9499 (N_9499,N_8833,N_8594);
nand U9500 (N_9500,N_8674,N_8878);
nand U9501 (N_9501,N_8593,N_8986);
or U9502 (N_9502,N_8237,N_8140);
or U9503 (N_9503,N_8519,N_8116);
and U9504 (N_9504,N_8255,N_8248);
and U9505 (N_9505,N_8455,N_8261);
nor U9506 (N_9506,N_8795,N_8801);
and U9507 (N_9507,N_8257,N_8144);
and U9508 (N_9508,N_8142,N_8762);
nand U9509 (N_9509,N_8117,N_8624);
nor U9510 (N_9510,N_8838,N_8947);
xor U9511 (N_9511,N_8479,N_8553);
or U9512 (N_9512,N_8302,N_8787);
nor U9513 (N_9513,N_8656,N_8517);
nor U9514 (N_9514,N_8642,N_8313);
or U9515 (N_9515,N_8109,N_8295);
nor U9516 (N_9516,N_8749,N_8402);
or U9517 (N_9517,N_8847,N_8082);
or U9518 (N_9518,N_8732,N_8883);
nand U9519 (N_9519,N_8956,N_8919);
xnor U9520 (N_9520,N_8990,N_8604);
nand U9521 (N_9521,N_8785,N_8605);
or U9522 (N_9522,N_8091,N_8560);
and U9523 (N_9523,N_8281,N_8898);
and U9524 (N_9524,N_8410,N_8689);
nand U9525 (N_9525,N_8928,N_8023);
and U9526 (N_9526,N_8026,N_8938);
nor U9527 (N_9527,N_8746,N_8383);
nand U9528 (N_9528,N_8196,N_8795);
or U9529 (N_9529,N_8180,N_8957);
xor U9530 (N_9530,N_8372,N_8622);
or U9531 (N_9531,N_8692,N_8543);
or U9532 (N_9532,N_8217,N_8295);
nand U9533 (N_9533,N_8692,N_8523);
or U9534 (N_9534,N_8555,N_8424);
xnor U9535 (N_9535,N_8422,N_8667);
or U9536 (N_9536,N_8369,N_8584);
nand U9537 (N_9537,N_8295,N_8247);
nand U9538 (N_9538,N_8937,N_8096);
xnor U9539 (N_9539,N_8619,N_8635);
and U9540 (N_9540,N_8584,N_8908);
nor U9541 (N_9541,N_8862,N_8541);
or U9542 (N_9542,N_8424,N_8729);
nand U9543 (N_9543,N_8711,N_8635);
nor U9544 (N_9544,N_8499,N_8130);
xnor U9545 (N_9545,N_8160,N_8394);
or U9546 (N_9546,N_8043,N_8873);
and U9547 (N_9547,N_8430,N_8001);
nor U9548 (N_9548,N_8341,N_8840);
or U9549 (N_9549,N_8844,N_8239);
or U9550 (N_9550,N_8246,N_8278);
nand U9551 (N_9551,N_8148,N_8686);
nor U9552 (N_9552,N_8568,N_8701);
or U9553 (N_9553,N_8877,N_8133);
and U9554 (N_9554,N_8461,N_8405);
xnor U9555 (N_9555,N_8922,N_8248);
nand U9556 (N_9556,N_8309,N_8169);
xor U9557 (N_9557,N_8463,N_8276);
xor U9558 (N_9558,N_8707,N_8142);
nand U9559 (N_9559,N_8464,N_8838);
xnor U9560 (N_9560,N_8892,N_8775);
and U9561 (N_9561,N_8553,N_8485);
nand U9562 (N_9562,N_8473,N_8134);
nand U9563 (N_9563,N_8846,N_8785);
nand U9564 (N_9564,N_8548,N_8359);
or U9565 (N_9565,N_8298,N_8893);
or U9566 (N_9566,N_8295,N_8425);
nand U9567 (N_9567,N_8233,N_8291);
and U9568 (N_9568,N_8896,N_8962);
or U9569 (N_9569,N_8194,N_8695);
and U9570 (N_9570,N_8928,N_8916);
and U9571 (N_9571,N_8933,N_8032);
and U9572 (N_9572,N_8507,N_8764);
and U9573 (N_9573,N_8042,N_8992);
xnor U9574 (N_9574,N_8878,N_8915);
and U9575 (N_9575,N_8055,N_8108);
nand U9576 (N_9576,N_8300,N_8378);
xnor U9577 (N_9577,N_8055,N_8476);
xor U9578 (N_9578,N_8418,N_8321);
xnor U9579 (N_9579,N_8139,N_8677);
nand U9580 (N_9580,N_8162,N_8063);
nand U9581 (N_9581,N_8015,N_8757);
or U9582 (N_9582,N_8950,N_8577);
or U9583 (N_9583,N_8046,N_8523);
or U9584 (N_9584,N_8519,N_8385);
xnor U9585 (N_9585,N_8046,N_8433);
nand U9586 (N_9586,N_8487,N_8414);
and U9587 (N_9587,N_8963,N_8470);
or U9588 (N_9588,N_8280,N_8507);
or U9589 (N_9589,N_8914,N_8821);
nor U9590 (N_9590,N_8697,N_8630);
xnor U9591 (N_9591,N_8669,N_8134);
and U9592 (N_9592,N_8011,N_8337);
nand U9593 (N_9593,N_8010,N_8059);
nand U9594 (N_9594,N_8976,N_8930);
and U9595 (N_9595,N_8551,N_8475);
and U9596 (N_9596,N_8448,N_8869);
nand U9597 (N_9597,N_8458,N_8726);
and U9598 (N_9598,N_8979,N_8298);
and U9599 (N_9599,N_8214,N_8467);
and U9600 (N_9600,N_8138,N_8602);
and U9601 (N_9601,N_8668,N_8297);
nor U9602 (N_9602,N_8021,N_8682);
and U9603 (N_9603,N_8830,N_8200);
nand U9604 (N_9604,N_8378,N_8367);
or U9605 (N_9605,N_8145,N_8452);
xor U9606 (N_9606,N_8129,N_8423);
and U9607 (N_9607,N_8900,N_8166);
or U9608 (N_9608,N_8164,N_8920);
and U9609 (N_9609,N_8955,N_8990);
xor U9610 (N_9610,N_8486,N_8824);
xor U9611 (N_9611,N_8943,N_8268);
xor U9612 (N_9612,N_8632,N_8159);
nor U9613 (N_9613,N_8805,N_8588);
xnor U9614 (N_9614,N_8514,N_8066);
xnor U9615 (N_9615,N_8286,N_8124);
nor U9616 (N_9616,N_8190,N_8453);
or U9617 (N_9617,N_8657,N_8512);
nor U9618 (N_9618,N_8710,N_8579);
nand U9619 (N_9619,N_8423,N_8508);
and U9620 (N_9620,N_8715,N_8569);
nand U9621 (N_9621,N_8481,N_8096);
xnor U9622 (N_9622,N_8764,N_8008);
nor U9623 (N_9623,N_8933,N_8685);
and U9624 (N_9624,N_8082,N_8353);
xnor U9625 (N_9625,N_8432,N_8505);
or U9626 (N_9626,N_8172,N_8910);
or U9627 (N_9627,N_8939,N_8581);
nor U9628 (N_9628,N_8987,N_8582);
or U9629 (N_9629,N_8677,N_8608);
and U9630 (N_9630,N_8456,N_8650);
nor U9631 (N_9631,N_8231,N_8937);
xor U9632 (N_9632,N_8877,N_8254);
and U9633 (N_9633,N_8630,N_8498);
and U9634 (N_9634,N_8110,N_8081);
nor U9635 (N_9635,N_8228,N_8621);
or U9636 (N_9636,N_8408,N_8348);
nand U9637 (N_9637,N_8959,N_8260);
or U9638 (N_9638,N_8121,N_8427);
xnor U9639 (N_9639,N_8831,N_8791);
xnor U9640 (N_9640,N_8039,N_8273);
and U9641 (N_9641,N_8227,N_8175);
xnor U9642 (N_9642,N_8473,N_8611);
nand U9643 (N_9643,N_8674,N_8234);
and U9644 (N_9644,N_8457,N_8295);
nor U9645 (N_9645,N_8050,N_8960);
and U9646 (N_9646,N_8598,N_8639);
and U9647 (N_9647,N_8164,N_8560);
xnor U9648 (N_9648,N_8223,N_8326);
nor U9649 (N_9649,N_8527,N_8358);
or U9650 (N_9650,N_8565,N_8666);
nor U9651 (N_9651,N_8031,N_8126);
or U9652 (N_9652,N_8698,N_8868);
and U9653 (N_9653,N_8393,N_8168);
nand U9654 (N_9654,N_8494,N_8510);
xor U9655 (N_9655,N_8079,N_8077);
xor U9656 (N_9656,N_8371,N_8477);
nand U9657 (N_9657,N_8099,N_8758);
nand U9658 (N_9658,N_8771,N_8454);
xor U9659 (N_9659,N_8518,N_8276);
nand U9660 (N_9660,N_8568,N_8556);
nor U9661 (N_9661,N_8460,N_8830);
nand U9662 (N_9662,N_8836,N_8250);
nor U9663 (N_9663,N_8451,N_8913);
nand U9664 (N_9664,N_8763,N_8152);
or U9665 (N_9665,N_8415,N_8508);
xor U9666 (N_9666,N_8932,N_8244);
nor U9667 (N_9667,N_8969,N_8961);
nor U9668 (N_9668,N_8610,N_8663);
or U9669 (N_9669,N_8339,N_8569);
or U9670 (N_9670,N_8434,N_8821);
nand U9671 (N_9671,N_8415,N_8115);
and U9672 (N_9672,N_8100,N_8386);
nand U9673 (N_9673,N_8977,N_8564);
nor U9674 (N_9674,N_8113,N_8777);
and U9675 (N_9675,N_8665,N_8622);
or U9676 (N_9676,N_8552,N_8521);
nand U9677 (N_9677,N_8206,N_8514);
nor U9678 (N_9678,N_8167,N_8923);
nor U9679 (N_9679,N_8746,N_8368);
nand U9680 (N_9680,N_8454,N_8047);
xor U9681 (N_9681,N_8336,N_8865);
nand U9682 (N_9682,N_8223,N_8551);
xor U9683 (N_9683,N_8098,N_8502);
xnor U9684 (N_9684,N_8785,N_8022);
xnor U9685 (N_9685,N_8729,N_8317);
nor U9686 (N_9686,N_8548,N_8011);
nand U9687 (N_9687,N_8933,N_8308);
nor U9688 (N_9688,N_8862,N_8911);
xnor U9689 (N_9689,N_8636,N_8089);
xnor U9690 (N_9690,N_8282,N_8340);
xor U9691 (N_9691,N_8502,N_8158);
and U9692 (N_9692,N_8114,N_8624);
or U9693 (N_9693,N_8876,N_8677);
xor U9694 (N_9694,N_8873,N_8293);
nand U9695 (N_9695,N_8659,N_8850);
nor U9696 (N_9696,N_8619,N_8463);
or U9697 (N_9697,N_8951,N_8499);
or U9698 (N_9698,N_8385,N_8919);
nand U9699 (N_9699,N_8590,N_8438);
xor U9700 (N_9700,N_8290,N_8292);
or U9701 (N_9701,N_8723,N_8721);
xor U9702 (N_9702,N_8916,N_8797);
and U9703 (N_9703,N_8201,N_8982);
and U9704 (N_9704,N_8252,N_8335);
xnor U9705 (N_9705,N_8520,N_8398);
or U9706 (N_9706,N_8990,N_8483);
or U9707 (N_9707,N_8165,N_8940);
and U9708 (N_9708,N_8621,N_8144);
and U9709 (N_9709,N_8539,N_8765);
xnor U9710 (N_9710,N_8412,N_8943);
or U9711 (N_9711,N_8261,N_8391);
or U9712 (N_9712,N_8765,N_8655);
or U9713 (N_9713,N_8821,N_8299);
and U9714 (N_9714,N_8191,N_8577);
or U9715 (N_9715,N_8940,N_8614);
and U9716 (N_9716,N_8381,N_8365);
nor U9717 (N_9717,N_8335,N_8978);
or U9718 (N_9718,N_8352,N_8492);
or U9719 (N_9719,N_8095,N_8879);
nand U9720 (N_9720,N_8138,N_8530);
xor U9721 (N_9721,N_8508,N_8257);
xor U9722 (N_9722,N_8852,N_8178);
and U9723 (N_9723,N_8259,N_8178);
nor U9724 (N_9724,N_8444,N_8197);
nor U9725 (N_9725,N_8863,N_8839);
nor U9726 (N_9726,N_8278,N_8507);
nand U9727 (N_9727,N_8010,N_8171);
and U9728 (N_9728,N_8405,N_8726);
nand U9729 (N_9729,N_8950,N_8033);
nand U9730 (N_9730,N_8391,N_8436);
xor U9731 (N_9731,N_8666,N_8354);
nand U9732 (N_9732,N_8383,N_8117);
and U9733 (N_9733,N_8423,N_8590);
nand U9734 (N_9734,N_8382,N_8671);
and U9735 (N_9735,N_8907,N_8793);
or U9736 (N_9736,N_8673,N_8327);
and U9737 (N_9737,N_8986,N_8111);
nor U9738 (N_9738,N_8029,N_8054);
and U9739 (N_9739,N_8533,N_8621);
nand U9740 (N_9740,N_8587,N_8322);
or U9741 (N_9741,N_8909,N_8468);
or U9742 (N_9742,N_8462,N_8336);
xor U9743 (N_9743,N_8141,N_8824);
or U9744 (N_9744,N_8420,N_8889);
and U9745 (N_9745,N_8028,N_8926);
nor U9746 (N_9746,N_8890,N_8575);
nand U9747 (N_9747,N_8700,N_8185);
xnor U9748 (N_9748,N_8969,N_8512);
nand U9749 (N_9749,N_8799,N_8919);
xor U9750 (N_9750,N_8869,N_8111);
nand U9751 (N_9751,N_8472,N_8353);
xor U9752 (N_9752,N_8170,N_8926);
nor U9753 (N_9753,N_8864,N_8580);
xor U9754 (N_9754,N_8631,N_8633);
nor U9755 (N_9755,N_8621,N_8614);
nand U9756 (N_9756,N_8885,N_8381);
nand U9757 (N_9757,N_8830,N_8030);
nor U9758 (N_9758,N_8964,N_8089);
nand U9759 (N_9759,N_8843,N_8668);
or U9760 (N_9760,N_8921,N_8639);
nand U9761 (N_9761,N_8609,N_8654);
nor U9762 (N_9762,N_8639,N_8883);
xor U9763 (N_9763,N_8122,N_8021);
nor U9764 (N_9764,N_8964,N_8346);
nand U9765 (N_9765,N_8830,N_8974);
or U9766 (N_9766,N_8063,N_8898);
xnor U9767 (N_9767,N_8306,N_8996);
nor U9768 (N_9768,N_8609,N_8288);
and U9769 (N_9769,N_8049,N_8226);
nand U9770 (N_9770,N_8785,N_8160);
and U9771 (N_9771,N_8845,N_8725);
xnor U9772 (N_9772,N_8247,N_8914);
and U9773 (N_9773,N_8805,N_8615);
and U9774 (N_9774,N_8661,N_8597);
or U9775 (N_9775,N_8685,N_8035);
and U9776 (N_9776,N_8732,N_8897);
xor U9777 (N_9777,N_8522,N_8171);
and U9778 (N_9778,N_8623,N_8352);
or U9779 (N_9779,N_8817,N_8959);
or U9780 (N_9780,N_8144,N_8812);
and U9781 (N_9781,N_8519,N_8704);
nor U9782 (N_9782,N_8799,N_8866);
xnor U9783 (N_9783,N_8577,N_8607);
nor U9784 (N_9784,N_8418,N_8913);
nor U9785 (N_9785,N_8857,N_8599);
nand U9786 (N_9786,N_8993,N_8169);
nor U9787 (N_9787,N_8061,N_8259);
nor U9788 (N_9788,N_8656,N_8728);
nor U9789 (N_9789,N_8764,N_8716);
nor U9790 (N_9790,N_8645,N_8867);
nand U9791 (N_9791,N_8822,N_8841);
xor U9792 (N_9792,N_8601,N_8245);
xnor U9793 (N_9793,N_8225,N_8013);
and U9794 (N_9794,N_8072,N_8780);
nor U9795 (N_9795,N_8517,N_8578);
and U9796 (N_9796,N_8033,N_8630);
xor U9797 (N_9797,N_8499,N_8821);
nand U9798 (N_9798,N_8517,N_8277);
and U9799 (N_9799,N_8810,N_8119);
xor U9800 (N_9800,N_8194,N_8729);
nand U9801 (N_9801,N_8727,N_8520);
or U9802 (N_9802,N_8394,N_8971);
and U9803 (N_9803,N_8972,N_8881);
and U9804 (N_9804,N_8382,N_8636);
and U9805 (N_9805,N_8937,N_8040);
nand U9806 (N_9806,N_8313,N_8527);
nor U9807 (N_9807,N_8884,N_8387);
xor U9808 (N_9808,N_8107,N_8800);
xor U9809 (N_9809,N_8284,N_8909);
nor U9810 (N_9810,N_8710,N_8973);
xor U9811 (N_9811,N_8554,N_8874);
xor U9812 (N_9812,N_8422,N_8034);
nor U9813 (N_9813,N_8119,N_8162);
nor U9814 (N_9814,N_8831,N_8699);
nand U9815 (N_9815,N_8369,N_8861);
xor U9816 (N_9816,N_8456,N_8429);
nor U9817 (N_9817,N_8668,N_8622);
nand U9818 (N_9818,N_8873,N_8040);
nor U9819 (N_9819,N_8502,N_8010);
xor U9820 (N_9820,N_8462,N_8073);
or U9821 (N_9821,N_8459,N_8876);
or U9822 (N_9822,N_8123,N_8328);
and U9823 (N_9823,N_8010,N_8594);
xnor U9824 (N_9824,N_8953,N_8917);
xnor U9825 (N_9825,N_8836,N_8504);
nand U9826 (N_9826,N_8327,N_8641);
nor U9827 (N_9827,N_8499,N_8766);
and U9828 (N_9828,N_8743,N_8571);
xor U9829 (N_9829,N_8516,N_8517);
and U9830 (N_9830,N_8273,N_8554);
xor U9831 (N_9831,N_8287,N_8023);
or U9832 (N_9832,N_8603,N_8350);
nor U9833 (N_9833,N_8085,N_8053);
nand U9834 (N_9834,N_8376,N_8577);
or U9835 (N_9835,N_8638,N_8527);
xnor U9836 (N_9836,N_8475,N_8237);
nor U9837 (N_9837,N_8426,N_8977);
and U9838 (N_9838,N_8961,N_8303);
nor U9839 (N_9839,N_8306,N_8770);
nand U9840 (N_9840,N_8773,N_8917);
xnor U9841 (N_9841,N_8222,N_8950);
xnor U9842 (N_9842,N_8505,N_8446);
and U9843 (N_9843,N_8994,N_8620);
nor U9844 (N_9844,N_8762,N_8845);
and U9845 (N_9845,N_8555,N_8585);
or U9846 (N_9846,N_8181,N_8279);
xor U9847 (N_9847,N_8983,N_8968);
nand U9848 (N_9848,N_8694,N_8158);
and U9849 (N_9849,N_8693,N_8712);
nand U9850 (N_9850,N_8334,N_8227);
nand U9851 (N_9851,N_8676,N_8182);
and U9852 (N_9852,N_8898,N_8500);
xnor U9853 (N_9853,N_8113,N_8340);
or U9854 (N_9854,N_8238,N_8157);
or U9855 (N_9855,N_8708,N_8021);
or U9856 (N_9856,N_8477,N_8765);
and U9857 (N_9857,N_8642,N_8821);
and U9858 (N_9858,N_8112,N_8338);
nand U9859 (N_9859,N_8884,N_8612);
nor U9860 (N_9860,N_8902,N_8539);
or U9861 (N_9861,N_8568,N_8075);
or U9862 (N_9862,N_8080,N_8078);
nand U9863 (N_9863,N_8685,N_8857);
and U9864 (N_9864,N_8572,N_8458);
nor U9865 (N_9865,N_8470,N_8547);
xor U9866 (N_9866,N_8684,N_8484);
nor U9867 (N_9867,N_8796,N_8071);
or U9868 (N_9868,N_8457,N_8855);
and U9869 (N_9869,N_8195,N_8893);
nand U9870 (N_9870,N_8579,N_8906);
xor U9871 (N_9871,N_8926,N_8456);
and U9872 (N_9872,N_8100,N_8080);
nor U9873 (N_9873,N_8791,N_8051);
or U9874 (N_9874,N_8753,N_8828);
nand U9875 (N_9875,N_8926,N_8731);
and U9876 (N_9876,N_8720,N_8314);
nor U9877 (N_9877,N_8047,N_8409);
xor U9878 (N_9878,N_8282,N_8405);
or U9879 (N_9879,N_8930,N_8591);
nand U9880 (N_9880,N_8222,N_8617);
nand U9881 (N_9881,N_8302,N_8281);
xnor U9882 (N_9882,N_8051,N_8895);
or U9883 (N_9883,N_8635,N_8075);
or U9884 (N_9884,N_8733,N_8750);
or U9885 (N_9885,N_8727,N_8864);
nor U9886 (N_9886,N_8530,N_8141);
xnor U9887 (N_9887,N_8429,N_8988);
or U9888 (N_9888,N_8999,N_8328);
or U9889 (N_9889,N_8247,N_8441);
nand U9890 (N_9890,N_8463,N_8030);
xnor U9891 (N_9891,N_8745,N_8094);
or U9892 (N_9892,N_8356,N_8741);
or U9893 (N_9893,N_8367,N_8732);
nand U9894 (N_9894,N_8592,N_8598);
nand U9895 (N_9895,N_8657,N_8533);
nand U9896 (N_9896,N_8860,N_8935);
nand U9897 (N_9897,N_8122,N_8452);
nand U9898 (N_9898,N_8404,N_8663);
nor U9899 (N_9899,N_8266,N_8434);
nor U9900 (N_9900,N_8073,N_8429);
nor U9901 (N_9901,N_8173,N_8276);
nand U9902 (N_9902,N_8184,N_8150);
and U9903 (N_9903,N_8325,N_8715);
nand U9904 (N_9904,N_8781,N_8962);
nand U9905 (N_9905,N_8670,N_8795);
nor U9906 (N_9906,N_8202,N_8113);
and U9907 (N_9907,N_8670,N_8682);
nand U9908 (N_9908,N_8422,N_8360);
xor U9909 (N_9909,N_8520,N_8782);
xor U9910 (N_9910,N_8706,N_8468);
nand U9911 (N_9911,N_8018,N_8591);
and U9912 (N_9912,N_8752,N_8543);
nor U9913 (N_9913,N_8149,N_8473);
nor U9914 (N_9914,N_8115,N_8010);
nand U9915 (N_9915,N_8037,N_8699);
and U9916 (N_9916,N_8695,N_8766);
or U9917 (N_9917,N_8304,N_8746);
or U9918 (N_9918,N_8387,N_8399);
xnor U9919 (N_9919,N_8307,N_8439);
nor U9920 (N_9920,N_8273,N_8540);
nor U9921 (N_9921,N_8671,N_8486);
and U9922 (N_9922,N_8270,N_8096);
nor U9923 (N_9923,N_8678,N_8142);
nand U9924 (N_9924,N_8021,N_8467);
or U9925 (N_9925,N_8587,N_8162);
or U9926 (N_9926,N_8650,N_8490);
and U9927 (N_9927,N_8998,N_8863);
and U9928 (N_9928,N_8207,N_8599);
xnor U9929 (N_9929,N_8461,N_8126);
nor U9930 (N_9930,N_8010,N_8984);
nand U9931 (N_9931,N_8571,N_8872);
and U9932 (N_9932,N_8311,N_8091);
or U9933 (N_9933,N_8226,N_8741);
or U9934 (N_9934,N_8946,N_8936);
and U9935 (N_9935,N_8469,N_8876);
nand U9936 (N_9936,N_8817,N_8459);
nor U9937 (N_9937,N_8215,N_8487);
and U9938 (N_9938,N_8705,N_8546);
nor U9939 (N_9939,N_8472,N_8367);
xnor U9940 (N_9940,N_8300,N_8406);
nor U9941 (N_9941,N_8463,N_8494);
nor U9942 (N_9942,N_8181,N_8919);
xnor U9943 (N_9943,N_8388,N_8149);
nor U9944 (N_9944,N_8637,N_8599);
or U9945 (N_9945,N_8638,N_8607);
xnor U9946 (N_9946,N_8014,N_8152);
or U9947 (N_9947,N_8646,N_8296);
nor U9948 (N_9948,N_8074,N_8898);
nor U9949 (N_9949,N_8024,N_8816);
nand U9950 (N_9950,N_8487,N_8932);
or U9951 (N_9951,N_8448,N_8593);
xor U9952 (N_9952,N_8530,N_8639);
nand U9953 (N_9953,N_8817,N_8166);
or U9954 (N_9954,N_8342,N_8641);
xnor U9955 (N_9955,N_8949,N_8133);
nand U9956 (N_9956,N_8215,N_8315);
xnor U9957 (N_9957,N_8058,N_8780);
or U9958 (N_9958,N_8837,N_8787);
nand U9959 (N_9959,N_8916,N_8140);
or U9960 (N_9960,N_8303,N_8171);
nor U9961 (N_9961,N_8315,N_8115);
and U9962 (N_9962,N_8143,N_8937);
xnor U9963 (N_9963,N_8294,N_8990);
nor U9964 (N_9964,N_8165,N_8047);
nand U9965 (N_9965,N_8051,N_8445);
nor U9966 (N_9966,N_8204,N_8637);
and U9967 (N_9967,N_8418,N_8697);
nor U9968 (N_9968,N_8683,N_8466);
nor U9969 (N_9969,N_8141,N_8391);
nand U9970 (N_9970,N_8263,N_8348);
nand U9971 (N_9971,N_8152,N_8068);
and U9972 (N_9972,N_8907,N_8785);
xnor U9973 (N_9973,N_8389,N_8168);
nand U9974 (N_9974,N_8377,N_8374);
nand U9975 (N_9975,N_8013,N_8583);
xor U9976 (N_9976,N_8680,N_8890);
or U9977 (N_9977,N_8845,N_8682);
xnor U9978 (N_9978,N_8918,N_8059);
and U9979 (N_9979,N_8943,N_8077);
or U9980 (N_9980,N_8195,N_8121);
and U9981 (N_9981,N_8886,N_8558);
or U9982 (N_9982,N_8041,N_8174);
xnor U9983 (N_9983,N_8451,N_8177);
nor U9984 (N_9984,N_8707,N_8531);
nand U9985 (N_9985,N_8314,N_8854);
nand U9986 (N_9986,N_8647,N_8722);
or U9987 (N_9987,N_8403,N_8152);
or U9988 (N_9988,N_8910,N_8361);
or U9989 (N_9989,N_8199,N_8210);
and U9990 (N_9990,N_8746,N_8080);
nor U9991 (N_9991,N_8663,N_8001);
or U9992 (N_9992,N_8761,N_8299);
or U9993 (N_9993,N_8328,N_8551);
and U9994 (N_9994,N_8979,N_8604);
or U9995 (N_9995,N_8632,N_8032);
and U9996 (N_9996,N_8244,N_8272);
xor U9997 (N_9997,N_8642,N_8720);
and U9998 (N_9998,N_8687,N_8952);
xnor U9999 (N_9999,N_8871,N_8646);
nand U10000 (N_10000,N_9569,N_9315);
nand U10001 (N_10001,N_9802,N_9388);
or U10002 (N_10002,N_9651,N_9346);
nor U10003 (N_10003,N_9548,N_9086);
nor U10004 (N_10004,N_9520,N_9509);
xnor U10005 (N_10005,N_9056,N_9498);
nor U10006 (N_10006,N_9545,N_9752);
or U10007 (N_10007,N_9360,N_9298);
xor U10008 (N_10008,N_9739,N_9811);
nor U10009 (N_10009,N_9319,N_9849);
or U10010 (N_10010,N_9603,N_9282);
xnor U10011 (N_10011,N_9402,N_9986);
nand U10012 (N_10012,N_9429,N_9636);
or U10013 (N_10013,N_9890,N_9858);
and U10014 (N_10014,N_9547,N_9597);
and U10015 (N_10015,N_9445,N_9683);
or U10016 (N_10016,N_9249,N_9472);
and U10017 (N_10017,N_9118,N_9085);
nor U10018 (N_10018,N_9238,N_9945);
nand U10019 (N_10019,N_9613,N_9769);
nor U10020 (N_10020,N_9782,N_9399);
nand U10021 (N_10021,N_9253,N_9316);
nand U10022 (N_10022,N_9129,N_9908);
or U10023 (N_10023,N_9771,N_9966);
and U10024 (N_10024,N_9307,N_9648);
nand U10025 (N_10025,N_9047,N_9265);
or U10026 (N_10026,N_9022,N_9518);
xor U10027 (N_10027,N_9462,N_9492);
xnor U10028 (N_10028,N_9968,N_9278);
nand U10029 (N_10029,N_9630,N_9294);
xnor U10030 (N_10030,N_9337,N_9694);
or U10031 (N_10031,N_9586,N_9093);
and U10032 (N_10032,N_9293,N_9913);
or U10033 (N_10033,N_9091,N_9715);
nor U10034 (N_10034,N_9497,N_9286);
nand U10035 (N_10035,N_9731,N_9372);
xnor U10036 (N_10036,N_9026,N_9324);
or U10037 (N_10037,N_9042,N_9098);
nor U10038 (N_10038,N_9979,N_9289);
nand U10039 (N_10039,N_9927,N_9824);
xnor U10040 (N_10040,N_9842,N_9175);
nand U10041 (N_10041,N_9364,N_9117);
and U10042 (N_10042,N_9875,N_9181);
xor U10043 (N_10043,N_9521,N_9303);
xnor U10044 (N_10044,N_9736,N_9721);
nand U10045 (N_10045,N_9790,N_9809);
nor U10046 (N_10046,N_9246,N_9228);
and U10047 (N_10047,N_9274,N_9755);
or U10048 (N_10048,N_9850,N_9052);
or U10049 (N_10049,N_9335,N_9095);
nand U10050 (N_10050,N_9301,N_9976);
nor U10051 (N_10051,N_9990,N_9926);
nand U10052 (N_10052,N_9114,N_9427);
nor U10053 (N_10053,N_9594,N_9733);
nor U10054 (N_10054,N_9798,N_9442);
or U10055 (N_10055,N_9552,N_9124);
xor U10056 (N_10056,N_9835,N_9706);
and U10057 (N_10057,N_9078,N_9515);
nor U10058 (N_10058,N_9297,N_9856);
or U10059 (N_10059,N_9283,N_9717);
xor U10060 (N_10060,N_9024,N_9628);
and U10061 (N_10061,N_9876,N_9311);
nor U10062 (N_10062,N_9176,N_9368);
and U10063 (N_10063,N_9336,N_9256);
xor U10064 (N_10064,N_9896,N_9140);
xnor U10065 (N_10065,N_9861,N_9312);
or U10066 (N_10066,N_9952,N_9882);
nand U10067 (N_10067,N_9379,N_9351);
and U10068 (N_10068,N_9050,N_9574);
nor U10069 (N_10069,N_9138,N_9792);
nand U10070 (N_10070,N_9043,N_9419);
or U10071 (N_10071,N_9587,N_9076);
or U10072 (N_10072,N_9641,N_9729);
nand U10073 (N_10073,N_9322,N_9864);
nor U10074 (N_10074,N_9061,N_9620);
and U10075 (N_10075,N_9101,N_9167);
nor U10076 (N_10076,N_9543,N_9754);
nor U10077 (N_10077,N_9653,N_9542);
and U10078 (N_10078,N_9938,N_9075);
or U10079 (N_10079,N_9295,N_9252);
nand U10080 (N_10080,N_9227,N_9676);
nand U10081 (N_10081,N_9190,N_9268);
and U10082 (N_10082,N_9354,N_9994);
or U10083 (N_10083,N_9870,N_9204);
nand U10084 (N_10084,N_9777,N_9746);
xnor U10085 (N_10085,N_9776,N_9530);
nand U10086 (N_10086,N_9115,N_9753);
or U10087 (N_10087,N_9242,N_9598);
xnor U10088 (N_10088,N_9031,N_9436);
xnor U10089 (N_10089,N_9284,N_9959);
or U10090 (N_10090,N_9884,N_9046);
nor U10091 (N_10091,N_9206,N_9434);
or U10092 (N_10092,N_9059,N_9524);
nor U10093 (N_10093,N_9881,N_9655);
nor U10094 (N_10094,N_9055,N_9918);
or U10095 (N_10095,N_9121,N_9431);
nor U10096 (N_10096,N_9669,N_9173);
or U10097 (N_10097,N_9558,N_9860);
and U10098 (N_10098,N_9350,N_9762);
and U10099 (N_10099,N_9185,N_9488);
and U10100 (N_10100,N_9133,N_9212);
or U10101 (N_10101,N_9131,N_9536);
nor U10102 (N_10102,N_9557,N_9659);
xnor U10103 (N_10103,N_9421,N_9418);
xnor U10104 (N_10104,N_9723,N_9290);
nand U10105 (N_10105,N_9296,N_9533);
xor U10106 (N_10106,N_9203,N_9663);
xor U10107 (N_10107,N_9394,N_9012);
or U10108 (N_10108,N_9915,N_9631);
nor U10109 (N_10109,N_9711,N_9578);
nor U10110 (N_10110,N_9887,N_9825);
and U10111 (N_10111,N_9447,N_9826);
nand U10112 (N_10112,N_9189,N_9656);
and U10113 (N_10113,N_9590,N_9216);
nor U10114 (N_10114,N_9259,N_9963);
xor U10115 (N_10115,N_9099,N_9270);
or U10116 (N_10116,N_9044,N_9374);
xor U10117 (N_10117,N_9218,N_9983);
xnor U10118 (N_10118,N_9852,N_9068);
or U10119 (N_10119,N_9949,N_9995);
nor U10120 (N_10120,N_9458,N_9693);
and U10121 (N_10121,N_9673,N_9898);
nand U10122 (N_10122,N_9485,N_9271);
nor U10123 (N_10123,N_9378,N_9821);
and U10124 (N_10124,N_9725,N_9599);
or U10125 (N_10125,N_9160,N_9305);
xor U10126 (N_10126,N_9440,N_9505);
nand U10127 (N_10127,N_9540,N_9899);
and U10128 (N_10128,N_9658,N_9103);
or U10129 (N_10129,N_9347,N_9111);
and U10130 (N_10130,N_9255,N_9567);
xnor U10131 (N_10131,N_9832,N_9925);
nor U10132 (N_10132,N_9965,N_9865);
or U10133 (N_10133,N_9981,N_9154);
and U10134 (N_10134,N_9074,N_9261);
or U10135 (N_10135,N_9386,N_9199);
and U10136 (N_10136,N_9281,N_9116);
xor U10137 (N_10137,N_9555,N_9058);
nand U10138 (N_10138,N_9709,N_9734);
nor U10139 (N_10139,N_9622,N_9195);
and U10140 (N_10140,N_9584,N_9819);
and U10141 (N_10141,N_9407,N_9690);
or U10142 (N_10142,N_9843,N_9992);
nand U10143 (N_10143,N_9013,N_9499);
nor U10144 (N_10144,N_9110,N_9695);
or U10145 (N_10145,N_9495,N_9980);
xnor U10146 (N_10146,N_9147,N_9522);
or U10147 (N_10147,N_9900,N_9214);
or U10148 (N_10148,N_9778,N_9080);
and U10149 (N_10149,N_9200,N_9452);
or U10150 (N_10150,N_9537,N_9610);
nand U10151 (N_10151,N_9714,N_9756);
nor U10152 (N_10152,N_9396,N_9291);
xor U10153 (N_10153,N_9814,N_9930);
and U10154 (N_10154,N_9506,N_9716);
xor U10155 (N_10155,N_9519,N_9308);
and U10156 (N_10156,N_9743,N_9482);
xor U10157 (N_10157,N_9053,N_9634);
xnor U10158 (N_10158,N_9371,N_9340);
nor U10159 (N_10159,N_9551,N_9381);
and U10160 (N_10160,N_9119,N_9223);
nor U10161 (N_10161,N_9880,N_9765);
and U10162 (N_10162,N_9546,N_9389);
nor U10163 (N_10163,N_9331,N_9239);
and U10164 (N_10164,N_9132,N_9465);
and U10165 (N_10165,N_9840,N_9349);
or U10166 (N_10166,N_9642,N_9939);
or U10167 (N_10167,N_9572,N_9146);
and U10168 (N_10168,N_9457,N_9243);
and U10169 (N_10169,N_9623,N_9142);
nor U10170 (N_10170,N_9954,N_9991);
or U10171 (N_10171,N_9463,N_9940);
and U10172 (N_10172,N_9647,N_9127);
nor U10173 (N_10173,N_9392,N_9873);
nand U10174 (N_10174,N_9692,N_9484);
nand U10175 (N_10175,N_9184,N_9788);
xnor U10176 (N_10176,N_9928,N_9747);
nand U10177 (N_10177,N_9446,N_9207);
or U10178 (N_10178,N_9757,N_9014);
xor U10179 (N_10179,N_9164,N_9006);
or U10180 (N_10180,N_9352,N_9330);
or U10181 (N_10181,N_9191,N_9640);
nand U10182 (N_10182,N_9577,N_9269);
and U10183 (N_10183,N_9510,N_9363);
or U10184 (N_10184,N_9801,N_9919);
nand U10185 (N_10185,N_9914,N_9410);
nor U10186 (N_10186,N_9100,N_9438);
and U10187 (N_10187,N_9051,N_9070);
nor U10188 (N_10188,N_9707,N_9772);
and U10189 (N_10189,N_9508,N_9512);
xnor U10190 (N_10190,N_9745,N_9960);
xnor U10191 (N_10191,N_9135,N_9891);
nor U10192 (N_10192,N_9426,N_9561);
nor U10193 (N_10193,N_9784,N_9621);
or U10194 (N_10194,N_9468,N_9941);
or U10195 (N_10195,N_9358,N_9632);
or U10196 (N_10196,N_9748,N_9299);
or U10197 (N_10197,N_9432,N_9170);
nor U10198 (N_10198,N_9333,N_9174);
and U10199 (N_10199,N_9550,N_9500);
nor U10200 (N_10200,N_9652,N_9177);
nor U10201 (N_10201,N_9805,N_9329);
or U10202 (N_10202,N_9904,N_9219);
nand U10203 (N_10203,N_9607,N_9263);
and U10204 (N_10204,N_9531,N_9011);
nor U10205 (N_10205,N_9866,N_9837);
and U10206 (N_10206,N_9982,N_9084);
or U10207 (N_10207,N_9035,N_9917);
or U10208 (N_10208,N_9205,N_9403);
nand U10209 (N_10209,N_9341,N_9209);
and U10210 (N_10210,N_9325,N_9559);
xnor U10211 (N_10211,N_9041,N_9857);
or U10212 (N_10212,N_9049,N_9638);
nor U10213 (N_10213,N_9883,N_9439);
or U10214 (N_10214,N_9871,N_9906);
and U10215 (N_10215,N_9997,N_9751);
nand U10216 (N_10216,N_9128,N_9766);
nor U10217 (N_10217,N_9948,N_9886);
xnor U10218 (N_10218,N_9689,N_9724);
or U10219 (N_10219,N_9491,N_9496);
xnor U10220 (N_10220,N_9057,N_9064);
or U10221 (N_10221,N_9951,N_9781);
or U10222 (N_10222,N_9092,N_9812);
nand U10223 (N_10223,N_9564,N_9387);
nor U10224 (N_10224,N_9169,N_9661);
or U10225 (N_10225,N_9685,N_9194);
or U10226 (N_10226,N_9454,N_9107);
nor U10227 (N_10227,N_9909,N_9827);
and U10228 (N_10228,N_9596,N_9361);
nor U10229 (N_10229,N_9813,N_9637);
xor U10230 (N_10230,N_9310,N_9415);
and U10231 (N_10231,N_9338,N_9353);
or U10232 (N_10232,N_9159,N_9040);
and U10233 (N_10233,N_9863,N_9565);
and U10234 (N_10234,N_9595,N_9304);
nand U10235 (N_10235,N_9066,N_9513);
nor U10236 (N_10236,N_9339,N_9947);
xnor U10237 (N_10237,N_9503,N_9878);
or U10238 (N_10238,N_9730,N_9018);
or U10239 (N_10239,N_9845,N_9483);
nand U10240 (N_10240,N_9376,N_9470);
or U10241 (N_10241,N_9466,N_9580);
nor U10242 (N_10242,N_9460,N_9646);
or U10243 (N_10243,N_9675,N_9701);
nand U10244 (N_10244,N_9156,N_9601);
and U10245 (N_10245,N_9088,N_9532);
nand U10246 (N_10246,N_9507,N_9526);
xor U10247 (N_10247,N_9712,N_9773);
and U10248 (N_10248,N_9258,N_9625);
nor U10249 (N_10249,N_9624,N_9728);
or U10250 (N_10250,N_9538,N_9517);
xnor U10251 (N_10251,N_9967,N_9097);
nand U10252 (N_10252,N_9453,N_9065);
nor U10253 (N_10253,N_9060,N_9422);
or U10254 (N_10254,N_9617,N_9732);
or U10255 (N_10255,N_9034,N_9198);
nand U10256 (N_10256,N_9806,N_9950);
or U10257 (N_10257,N_9749,N_9944);
and U10258 (N_10258,N_9231,N_9414);
nand U10259 (N_10259,N_9592,N_9287);
xnor U10260 (N_10260,N_9375,N_9657);
and U10261 (N_10261,N_9089,N_9823);
and U10262 (N_10262,N_9145,N_9443);
nand U10263 (N_10263,N_9961,N_9187);
xnor U10264 (N_10264,N_9528,N_9467);
nand U10265 (N_10265,N_9393,N_9544);
and U10266 (N_10266,N_9910,N_9916);
xnor U10267 (N_10267,N_9831,N_9178);
xor U10268 (N_10268,N_9534,N_9390);
nor U10269 (N_10269,N_9942,N_9874);
xnor U10270 (N_10270,N_9527,N_9413);
xnor U10271 (N_10271,N_9273,N_9582);
xnor U10272 (N_10272,N_9702,N_9137);
xnor U10273 (N_10273,N_9213,N_9847);
nand U10274 (N_10274,N_9931,N_9365);
nand U10275 (N_10275,N_9869,N_9230);
and U10276 (N_10276,N_9989,N_9401);
nand U10277 (N_10277,N_9226,N_9962);
and U10278 (N_10278,N_9045,N_9314);
nor U10279 (N_10279,N_9614,N_9541);
nand U10280 (N_10280,N_9829,N_9568);
nand U10281 (N_10281,N_9015,N_9276);
nand U10282 (N_10282,N_9215,N_9416);
and U10283 (N_10283,N_9334,N_9957);
and U10284 (N_10284,N_9449,N_9744);
and U10285 (N_10285,N_9328,N_9794);
nand U10286 (N_10286,N_9775,N_9435);
xnor U10287 (N_10287,N_9188,N_9955);
or U10288 (N_10288,N_9722,N_9150);
xor U10289 (N_10289,N_9556,N_9566);
nor U10290 (N_10290,N_9490,N_9633);
and U10291 (N_10291,N_9946,N_9923);
or U10292 (N_10292,N_9583,N_9108);
nand U10293 (N_10293,N_9236,N_9936);
nor U10294 (N_10294,N_9077,N_9083);
xor U10295 (N_10295,N_9224,N_9313);
and U10296 (N_10296,N_9385,N_9677);
nand U10297 (N_10297,N_9841,N_9667);
nor U10298 (N_10298,N_9697,N_9851);
and U10299 (N_10299,N_9604,N_9999);
nor U10300 (N_10300,N_9241,N_9885);
nor U10301 (N_10301,N_9102,N_9958);
xor U10302 (N_10302,N_9395,N_9761);
nor U10303 (N_10303,N_9535,N_9616);
or U10304 (N_10304,N_9735,N_9588);
nand U10305 (N_10305,N_9810,N_9785);
and U10306 (N_10306,N_9019,N_9016);
and U10307 (N_10307,N_9643,N_9602);
and U10308 (N_10308,N_9033,N_9681);
nand U10309 (N_10309,N_9130,N_9705);
or U10310 (N_10310,N_9359,N_9245);
and U10311 (N_10311,N_9803,N_9589);
nand U10312 (N_10312,N_9032,N_9423);
or U10313 (N_10313,N_9366,N_9300);
and U10314 (N_10314,N_9929,N_9593);
and U10315 (N_10315,N_9023,N_9113);
or U10316 (N_10316,N_9902,N_9320);
and U10317 (N_10317,N_9171,N_9411);
nor U10318 (N_10318,N_9397,N_9839);
and U10319 (N_10319,N_9029,N_9501);
nor U10320 (N_10320,N_9877,N_9708);
nor U10321 (N_10321,N_9036,N_9005);
nand U10322 (N_10322,N_9853,N_9609);
nor U10323 (N_10323,N_9937,N_9678);
or U10324 (N_10324,N_9571,N_9816);
nand U10325 (N_10325,N_9525,N_9367);
xnor U10326 (N_10326,N_9451,N_9740);
xor U10327 (N_10327,N_9554,N_9345);
and U10328 (N_10328,N_9606,N_9973);
and U10329 (N_10329,N_9398,N_9815);
xnor U10330 (N_10330,N_9787,N_9846);
nor U10331 (N_10331,N_9644,N_9179);
and U10332 (N_10332,N_9838,N_9240);
and U10333 (N_10333,N_9348,N_9165);
nand U10334 (N_10334,N_9217,N_9808);
nand U10335 (N_10335,N_9072,N_9126);
xnor U10336 (N_10336,N_9428,N_9010);
and U10337 (N_10337,N_9618,N_9139);
and U10338 (N_10338,N_9844,N_9600);
xnor U10339 (N_10339,N_9894,N_9082);
xor U10340 (N_10340,N_9799,N_9575);
xnor U10341 (N_10341,N_9988,N_9459);
xnor U10342 (N_10342,N_9069,N_9087);
xnor U10343 (N_10343,N_9267,N_9612);
and U10344 (N_10344,N_9786,N_9017);
nor U10345 (N_10345,N_9232,N_9163);
nand U10346 (N_10346,N_9549,N_9514);
and U10347 (N_10347,N_9420,N_9235);
xor U10348 (N_10348,N_9605,N_9476);
xor U10349 (N_10349,N_9474,N_9125);
or U10350 (N_10350,N_9148,N_9934);
nor U10351 (N_10351,N_9244,N_9222);
or U10352 (N_10352,N_9713,N_9275);
or U10353 (N_10353,N_9079,N_9134);
and U10354 (N_10354,N_9668,N_9166);
and U10355 (N_10355,N_9738,N_9182);
nor U10356 (N_10356,N_9680,N_9956);
and U10357 (N_10357,N_9326,N_9473);
nand U10358 (N_10358,N_9817,N_9234);
and U10359 (N_10359,N_9048,N_9155);
or U10360 (N_10360,N_9037,N_9674);
nor U10361 (N_10361,N_9987,N_9479);
or U10362 (N_10362,N_9953,N_9264);
or U10363 (N_10363,N_9285,N_9562);
nor U10364 (N_10364,N_9964,N_9486);
or U10365 (N_10365,N_9000,N_9654);
nor U10366 (N_10366,N_9854,N_9943);
nand U10367 (N_10367,N_9789,N_9935);
and U10368 (N_10368,N_9292,N_9704);
xor U10369 (N_10369,N_9820,N_9237);
nor U10370 (N_10370,N_9073,N_9691);
or U10371 (N_10371,N_9020,N_9998);
and U10372 (N_10372,N_9469,N_9067);
or U10373 (N_10373,N_9323,N_9383);
nor U10374 (N_10374,N_9248,N_9581);
nor U10375 (N_10375,N_9382,N_9162);
nand U10376 (N_10376,N_9489,N_9855);
or U10377 (N_10377,N_9288,N_9409);
or U10378 (N_10378,N_9143,N_9627);
nor U10379 (N_10379,N_9280,N_9028);
xnor U10380 (N_10380,N_9985,N_9570);
and U10381 (N_10381,N_9027,N_9441);
xnor U10382 (N_10382,N_9975,N_9619);
nor U10383 (N_10383,N_9225,N_9591);
nor U10384 (N_10384,N_9796,N_9779);
and U10385 (N_10385,N_9974,N_9767);
or U10386 (N_10386,N_9272,N_9795);
xnor U10387 (N_10387,N_9406,N_9700);
xor U10388 (N_10388,N_9727,N_9480);
nand U10389 (N_10389,N_9062,N_9670);
nand U10390 (N_10390,N_9471,N_9626);
nand U10391 (N_10391,N_9141,N_9671);
and U10392 (N_10392,N_9201,N_9266);
and U10393 (N_10393,N_9412,N_9071);
and U10394 (N_10394,N_9400,N_9741);
nor U10395 (N_10395,N_9197,N_9684);
xor U10396 (N_10396,N_9151,N_9054);
and U10397 (N_10397,N_9122,N_9511);
xnor U10398 (N_10398,N_9905,N_9211);
nor U10399 (N_10399,N_9764,N_9493);
nand U10400 (N_10400,N_9615,N_9710);
xor U10401 (N_10401,N_9972,N_9193);
nand U10402 (N_10402,N_9149,N_9932);
xnor U10403 (N_10403,N_9897,N_9120);
and U10404 (N_10404,N_9144,N_9112);
or U10405 (N_10405,N_9196,N_9868);
xnor U10406 (N_10406,N_9257,N_9933);
or U10407 (N_10407,N_9828,N_9008);
or U10408 (N_10408,N_9742,N_9760);
and U10409 (N_10409,N_9660,N_9002);
xor U10410 (N_10410,N_9791,N_9220);
nor U10411 (N_10411,N_9699,N_9404);
xnor U10412 (N_10412,N_9090,N_9608);
nand U10413 (N_10413,N_9136,N_9993);
nor U10414 (N_10414,N_9001,N_9007);
and U10415 (N_10415,N_9254,N_9780);
nand U10416 (N_10416,N_9892,N_9461);
nor U10417 (N_10417,N_9202,N_9096);
xor U10418 (N_10418,N_9025,N_9342);
nand U10419 (N_10419,N_9377,N_9576);
xor U10420 (N_10420,N_9553,N_9487);
nand U10421 (N_10421,N_9081,N_9836);
nand U10422 (N_10422,N_9168,N_9317);
nand U10423 (N_10423,N_9343,N_9437);
and U10424 (N_10424,N_9094,N_9105);
nand U10425 (N_10425,N_9210,N_9158);
and U10426 (N_10426,N_9759,N_9830);
and U10427 (N_10427,N_9768,N_9356);
and U10428 (N_10428,N_9645,N_9318);
xor U10429 (N_10429,N_9448,N_9038);
xor U10430 (N_10430,N_9635,N_9425);
nor U10431 (N_10431,N_9970,N_9718);
or U10432 (N_10432,N_9260,N_9180);
nand U10433 (N_10433,N_9221,N_9424);
xnor U10434 (N_10434,N_9233,N_9106);
nor U10435 (N_10435,N_9996,N_9327);
nor U10436 (N_10436,N_9384,N_9560);
nor U10437 (N_10437,N_9879,N_9009);
nand U10438 (N_10438,N_9719,N_9464);
nor U10439 (N_10439,N_9478,N_9573);
or U10440 (N_10440,N_9247,N_9912);
or U10441 (N_10441,N_9822,N_9380);
and U10442 (N_10442,N_9893,N_9494);
or U10443 (N_10443,N_9003,N_9922);
or U10444 (N_10444,N_9611,N_9889);
nand U10445 (N_10445,N_9430,N_9834);
nor U10446 (N_10446,N_9585,N_9123);
or U10447 (N_10447,N_9357,N_9726);
nand U10448 (N_10448,N_9192,N_9502);
and U10449 (N_10449,N_9370,N_9978);
nand U10450 (N_10450,N_9679,N_9475);
or U10451 (N_10451,N_9797,N_9183);
or U10452 (N_10452,N_9186,N_9277);
and U10453 (N_10453,N_9455,N_9665);
and U10454 (N_10454,N_9369,N_9109);
and U10455 (N_10455,N_9504,N_9539);
or U10456 (N_10456,N_9172,N_9867);
nand U10457 (N_10457,N_9030,N_9672);
xor U10458 (N_10458,N_9862,N_9279);
or U10459 (N_10459,N_9523,N_9306);
or U10460 (N_10460,N_9450,N_9516);
or U10461 (N_10461,N_9859,N_9924);
xor U10462 (N_10462,N_9662,N_9444);
or U10463 (N_10463,N_9774,N_9686);
xor U10464 (N_10464,N_9639,N_9262);
nand U10465 (N_10465,N_9800,N_9650);
nand U10466 (N_10466,N_9833,N_9477);
xnor U10467 (N_10467,N_9698,N_9804);
nor U10468 (N_10468,N_9417,N_9344);
nand U10469 (N_10469,N_9250,N_9579);
nor U10470 (N_10470,N_9063,N_9903);
xor U10471 (N_10471,N_9004,N_9895);
nor U10472 (N_10472,N_9157,N_9362);
nand U10473 (N_10473,N_9309,N_9373);
nor U10474 (N_10474,N_9251,N_9161);
and U10475 (N_10475,N_9907,N_9971);
nor U10476 (N_10476,N_9302,N_9563);
nor U10477 (N_10477,N_9391,N_9984);
and U10478 (N_10478,N_9481,N_9104);
and U10479 (N_10479,N_9332,N_9229);
nand U10480 (N_10480,N_9408,N_9921);
nand U10481 (N_10481,N_9649,N_9793);
xnor U10482 (N_10482,N_9758,N_9529);
nor U10483 (N_10483,N_9770,N_9664);
or U10484 (N_10484,N_9763,N_9783);
nand U10485 (N_10485,N_9405,N_9687);
and U10486 (N_10486,N_9920,N_9969);
nand U10487 (N_10487,N_9208,N_9321);
nor U10488 (N_10488,N_9153,N_9872);
and U10489 (N_10489,N_9152,N_9901);
nor U10490 (N_10490,N_9696,N_9720);
and U10491 (N_10491,N_9911,N_9456);
or U10492 (N_10492,N_9888,N_9703);
or U10493 (N_10493,N_9355,N_9682);
nor U10494 (N_10494,N_9629,N_9666);
nor U10495 (N_10495,N_9750,N_9818);
nand U10496 (N_10496,N_9039,N_9433);
nor U10497 (N_10497,N_9977,N_9688);
nand U10498 (N_10498,N_9737,N_9807);
and U10499 (N_10499,N_9848,N_9021);
nand U10500 (N_10500,N_9692,N_9606);
nand U10501 (N_10501,N_9480,N_9134);
and U10502 (N_10502,N_9351,N_9100);
and U10503 (N_10503,N_9423,N_9140);
nor U10504 (N_10504,N_9893,N_9026);
or U10505 (N_10505,N_9449,N_9415);
or U10506 (N_10506,N_9182,N_9914);
or U10507 (N_10507,N_9909,N_9437);
or U10508 (N_10508,N_9910,N_9683);
or U10509 (N_10509,N_9370,N_9914);
xnor U10510 (N_10510,N_9671,N_9364);
or U10511 (N_10511,N_9931,N_9178);
nand U10512 (N_10512,N_9772,N_9139);
or U10513 (N_10513,N_9291,N_9883);
nand U10514 (N_10514,N_9052,N_9740);
nor U10515 (N_10515,N_9017,N_9527);
nand U10516 (N_10516,N_9614,N_9973);
xnor U10517 (N_10517,N_9923,N_9971);
and U10518 (N_10518,N_9052,N_9412);
and U10519 (N_10519,N_9319,N_9527);
nand U10520 (N_10520,N_9435,N_9793);
nand U10521 (N_10521,N_9558,N_9896);
xor U10522 (N_10522,N_9709,N_9111);
xor U10523 (N_10523,N_9615,N_9223);
and U10524 (N_10524,N_9102,N_9714);
and U10525 (N_10525,N_9948,N_9072);
nand U10526 (N_10526,N_9700,N_9525);
or U10527 (N_10527,N_9323,N_9622);
nor U10528 (N_10528,N_9835,N_9499);
xor U10529 (N_10529,N_9546,N_9604);
or U10530 (N_10530,N_9646,N_9270);
xnor U10531 (N_10531,N_9791,N_9225);
and U10532 (N_10532,N_9528,N_9240);
nand U10533 (N_10533,N_9777,N_9296);
and U10534 (N_10534,N_9185,N_9011);
or U10535 (N_10535,N_9452,N_9360);
nor U10536 (N_10536,N_9550,N_9319);
xnor U10537 (N_10537,N_9289,N_9943);
xnor U10538 (N_10538,N_9103,N_9134);
nand U10539 (N_10539,N_9360,N_9390);
and U10540 (N_10540,N_9782,N_9111);
or U10541 (N_10541,N_9948,N_9946);
and U10542 (N_10542,N_9760,N_9058);
nand U10543 (N_10543,N_9260,N_9961);
and U10544 (N_10544,N_9381,N_9602);
nand U10545 (N_10545,N_9011,N_9581);
or U10546 (N_10546,N_9015,N_9850);
nor U10547 (N_10547,N_9798,N_9852);
and U10548 (N_10548,N_9711,N_9957);
nand U10549 (N_10549,N_9004,N_9629);
and U10550 (N_10550,N_9024,N_9228);
nor U10551 (N_10551,N_9148,N_9981);
nand U10552 (N_10552,N_9386,N_9088);
xor U10553 (N_10553,N_9611,N_9459);
and U10554 (N_10554,N_9456,N_9258);
and U10555 (N_10555,N_9782,N_9883);
nor U10556 (N_10556,N_9482,N_9873);
nand U10557 (N_10557,N_9036,N_9932);
or U10558 (N_10558,N_9330,N_9009);
xnor U10559 (N_10559,N_9227,N_9060);
and U10560 (N_10560,N_9101,N_9230);
nor U10561 (N_10561,N_9345,N_9342);
nand U10562 (N_10562,N_9823,N_9684);
and U10563 (N_10563,N_9684,N_9104);
and U10564 (N_10564,N_9849,N_9962);
or U10565 (N_10565,N_9480,N_9312);
or U10566 (N_10566,N_9818,N_9379);
or U10567 (N_10567,N_9499,N_9303);
nor U10568 (N_10568,N_9025,N_9303);
nand U10569 (N_10569,N_9853,N_9215);
xnor U10570 (N_10570,N_9741,N_9525);
nand U10571 (N_10571,N_9234,N_9731);
nand U10572 (N_10572,N_9676,N_9830);
nand U10573 (N_10573,N_9229,N_9222);
and U10574 (N_10574,N_9139,N_9911);
xor U10575 (N_10575,N_9668,N_9545);
nor U10576 (N_10576,N_9494,N_9941);
nor U10577 (N_10577,N_9728,N_9855);
nor U10578 (N_10578,N_9562,N_9122);
and U10579 (N_10579,N_9216,N_9330);
nor U10580 (N_10580,N_9697,N_9469);
xnor U10581 (N_10581,N_9832,N_9186);
nor U10582 (N_10582,N_9322,N_9957);
and U10583 (N_10583,N_9499,N_9027);
or U10584 (N_10584,N_9411,N_9448);
and U10585 (N_10585,N_9276,N_9845);
xnor U10586 (N_10586,N_9002,N_9803);
nor U10587 (N_10587,N_9379,N_9782);
and U10588 (N_10588,N_9643,N_9323);
nand U10589 (N_10589,N_9391,N_9887);
nor U10590 (N_10590,N_9824,N_9232);
or U10591 (N_10591,N_9050,N_9729);
xor U10592 (N_10592,N_9271,N_9768);
and U10593 (N_10593,N_9383,N_9632);
nand U10594 (N_10594,N_9462,N_9675);
nor U10595 (N_10595,N_9019,N_9704);
xnor U10596 (N_10596,N_9054,N_9506);
and U10597 (N_10597,N_9568,N_9087);
nor U10598 (N_10598,N_9535,N_9548);
or U10599 (N_10599,N_9198,N_9592);
nand U10600 (N_10600,N_9900,N_9095);
xor U10601 (N_10601,N_9668,N_9407);
or U10602 (N_10602,N_9143,N_9497);
nor U10603 (N_10603,N_9700,N_9766);
nor U10604 (N_10604,N_9875,N_9449);
nand U10605 (N_10605,N_9481,N_9669);
or U10606 (N_10606,N_9388,N_9837);
nand U10607 (N_10607,N_9693,N_9047);
and U10608 (N_10608,N_9341,N_9519);
or U10609 (N_10609,N_9865,N_9743);
xnor U10610 (N_10610,N_9700,N_9622);
nand U10611 (N_10611,N_9640,N_9574);
and U10612 (N_10612,N_9894,N_9055);
nor U10613 (N_10613,N_9524,N_9683);
nand U10614 (N_10614,N_9956,N_9768);
nand U10615 (N_10615,N_9215,N_9545);
xnor U10616 (N_10616,N_9168,N_9095);
xor U10617 (N_10617,N_9728,N_9556);
or U10618 (N_10618,N_9914,N_9723);
or U10619 (N_10619,N_9721,N_9178);
nor U10620 (N_10620,N_9177,N_9674);
and U10621 (N_10621,N_9526,N_9824);
xor U10622 (N_10622,N_9895,N_9830);
nand U10623 (N_10623,N_9861,N_9976);
and U10624 (N_10624,N_9528,N_9811);
xor U10625 (N_10625,N_9599,N_9668);
nand U10626 (N_10626,N_9612,N_9746);
xor U10627 (N_10627,N_9539,N_9355);
and U10628 (N_10628,N_9594,N_9499);
xor U10629 (N_10629,N_9151,N_9915);
and U10630 (N_10630,N_9357,N_9599);
and U10631 (N_10631,N_9903,N_9074);
nand U10632 (N_10632,N_9899,N_9181);
nor U10633 (N_10633,N_9955,N_9644);
and U10634 (N_10634,N_9787,N_9222);
and U10635 (N_10635,N_9909,N_9071);
and U10636 (N_10636,N_9141,N_9754);
and U10637 (N_10637,N_9076,N_9849);
and U10638 (N_10638,N_9694,N_9320);
or U10639 (N_10639,N_9202,N_9180);
xor U10640 (N_10640,N_9126,N_9721);
xor U10641 (N_10641,N_9293,N_9397);
and U10642 (N_10642,N_9854,N_9433);
xnor U10643 (N_10643,N_9199,N_9736);
nor U10644 (N_10644,N_9826,N_9630);
nor U10645 (N_10645,N_9528,N_9819);
xor U10646 (N_10646,N_9083,N_9863);
nor U10647 (N_10647,N_9093,N_9067);
nand U10648 (N_10648,N_9763,N_9656);
nand U10649 (N_10649,N_9984,N_9865);
or U10650 (N_10650,N_9308,N_9816);
and U10651 (N_10651,N_9728,N_9382);
nand U10652 (N_10652,N_9824,N_9925);
nand U10653 (N_10653,N_9932,N_9500);
xor U10654 (N_10654,N_9356,N_9780);
or U10655 (N_10655,N_9258,N_9083);
and U10656 (N_10656,N_9701,N_9703);
xnor U10657 (N_10657,N_9931,N_9833);
and U10658 (N_10658,N_9223,N_9576);
and U10659 (N_10659,N_9599,N_9340);
and U10660 (N_10660,N_9019,N_9223);
nand U10661 (N_10661,N_9200,N_9965);
nand U10662 (N_10662,N_9290,N_9630);
or U10663 (N_10663,N_9637,N_9880);
xor U10664 (N_10664,N_9964,N_9454);
xnor U10665 (N_10665,N_9458,N_9609);
and U10666 (N_10666,N_9747,N_9121);
or U10667 (N_10667,N_9357,N_9399);
or U10668 (N_10668,N_9959,N_9485);
nor U10669 (N_10669,N_9953,N_9245);
and U10670 (N_10670,N_9347,N_9622);
and U10671 (N_10671,N_9158,N_9184);
and U10672 (N_10672,N_9468,N_9785);
and U10673 (N_10673,N_9506,N_9293);
xnor U10674 (N_10674,N_9778,N_9022);
nand U10675 (N_10675,N_9988,N_9569);
or U10676 (N_10676,N_9695,N_9609);
or U10677 (N_10677,N_9453,N_9612);
or U10678 (N_10678,N_9395,N_9810);
and U10679 (N_10679,N_9892,N_9476);
and U10680 (N_10680,N_9472,N_9246);
nor U10681 (N_10681,N_9502,N_9017);
xnor U10682 (N_10682,N_9261,N_9357);
nand U10683 (N_10683,N_9994,N_9834);
nand U10684 (N_10684,N_9695,N_9766);
and U10685 (N_10685,N_9013,N_9437);
xor U10686 (N_10686,N_9281,N_9783);
nor U10687 (N_10687,N_9692,N_9210);
or U10688 (N_10688,N_9414,N_9467);
nand U10689 (N_10689,N_9765,N_9216);
or U10690 (N_10690,N_9598,N_9460);
and U10691 (N_10691,N_9577,N_9592);
nand U10692 (N_10692,N_9113,N_9399);
and U10693 (N_10693,N_9401,N_9941);
or U10694 (N_10694,N_9772,N_9429);
nand U10695 (N_10695,N_9912,N_9921);
nor U10696 (N_10696,N_9981,N_9382);
and U10697 (N_10697,N_9250,N_9488);
and U10698 (N_10698,N_9371,N_9550);
nand U10699 (N_10699,N_9838,N_9316);
nor U10700 (N_10700,N_9315,N_9005);
nor U10701 (N_10701,N_9298,N_9392);
nand U10702 (N_10702,N_9487,N_9961);
and U10703 (N_10703,N_9879,N_9742);
nand U10704 (N_10704,N_9410,N_9998);
xor U10705 (N_10705,N_9228,N_9551);
or U10706 (N_10706,N_9252,N_9075);
xor U10707 (N_10707,N_9180,N_9607);
xnor U10708 (N_10708,N_9434,N_9431);
xor U10709 (N_10709,N_9196,N_9811);
nand U10710 (N_10710,N_9209,N_9190);
xor U10711 (N_10711,N_9856,N_9167);
or U10712 (N_10712,N_9380,N_9107);
nor U10713 (N_10713,N_9763,N_9928);
xnor U10714 (N_10714,N_9663,N_9900);
or U10715 (N_10715,N_9198,N_9284);
and U10716 (N_10716,N_9301,N_9535);
xor U10717 (N_10717,N_9360,N_9194);
nor U10718 (N_10718,N_9272,N_9444);
xor U10719 (N_10719,N_9642,N_9511);
nor U10720 (N_10720,N_9038,N_9856);
xor U10721 (N_10721,N_9607,N_9083);
xor U10722 (N_10722,N_9595,N_9779);
xor U10723 (N_10723,N_9362,N_9460);
xnor U10724 (N_10724,N_9017,N_9312);
nor U10725 (N_10725,N_9357,N_9816);
nand U10726 (N_10726,N_9956,N_9149);
and U10727 (N_10727,N_9453,N_9674);
or U10728 (N_10728,N_9506,N_9321);
xor U10729 (N_10729,N_9839,N_9374);
and U10730 (N_10730,N_9047,N_9175);
and U10731 (N_10731,N_9050,N_9323);
or U10732 (N_10732,N_9760,N_9134);
or U10733 (N_10733,N_9229,N_9154);
and U10734 (N_10734,N_9628,N_9268);
xor U10735 (N_10735,N_9895,N_9888);
or U10736 (N_10736,N_9560,N_9873);
xor U10737 (N_10737,N_9436,N_9205);
nand U10738 (N_10738,N_9588,N_9024);
nor U10739 (N_10739,N_9299,N_9019);
or U10740 (N_10740,N_9619,N_9977);
and U10741 (N_10741,N_9859,N_9404);
xor U10742 (N_10742,N_9698,N_9776);
or U10743 (N_10743,N_9437,N_9008);
nor U10744 (N_10744,N_9095,N_9741);
nor U10745 (N_10745,N_9578,N_9923);
nand U10746 (N_10746,N_9298,N_9075);
and U10747 (N_10747,N_9566,N_9494);
nand U10748 (N_10748,N_9619,N_9114);
or U10749 (N_10749,N_9283,N_9779);
nor U10750 (N_10750,N_9763,N_9478);
and U10751 (N_10751,N_9249,N_9555);
nand U10752 (N_10752,N_9385,N_9608);
or U10753 (N_10753,N_9542,N_9177);
and U10754 (N_10754,N_9622,N_9669);
and U10755 (N_10755,N_9384,N_9871);
or U10756 (N_10756,N_9759,N_9515);
nand U10757 (N_10757,N_9334,N_9043);
xnor U10758 (N_10758,N_9443,N_9853);
xor U10759 (N_10759,N_9531,N_9372);
nor U10760 (N_10760,N_9505,N_9027);
nand U10761 (N_10761,N_9724,N_9609);
nor U10762 (N_10762,N_9730,N_9055);
and U10763 (N_10763,N_9145,N_9118);
or U10764 (N_10764,N_9901,N_9206);
and U10765 (N_10765,N_9710,N_9010);
nor U10766 (N_10766,N_9524,N_9714);
and U10767 (N_10767,N_9375,N_9702);
nand U10768 (N_10768,N_9065,N_9362);
nand U10769 (N_10769,N_9355,N_9244);
xor U10770 (N_10770,N_9552,N_9912);
nor U10771 (N_10771,N_9470,N_9740);
or U10772 (N_10772,N_9669,N_9081);
xor U10773 (N_10773,N_9216,N_9333);
and U10774 (N_10774,N_9397,N_9530);
xor U10775 (N_10775,N_9801,N_9865);
nand U10776 (N_10776,N_9872,N_9951);
or U10777 (N_10777,N_9690,N_9858);
xor U10778 (N_10778,N_9916,N_9208);
nor U10779 (N_10779,N_9964,N_9140);
and U10780 (N_10780,N_9013,N_9290);
nand U10781 (N_10781,N_9328,N_9348);
nor U10782 (N_10782,N_9696,N_9652);
and U10783 (N_10783,N_9285,N_9880);
and U10784 (N_10784,N_9626,N_9692);
nor U10785 (N_10785,N_9510,N_9644);
xor U10786 (N_10786,N_9718,N_9205);
or U10787 (N_10787,N_9526,N_9903);
xor U10788 (N_10788,N_9532,N_9679);
or U10789 (N_10789,N_9534,N_9930);
nand U10790 (N_10790,N_9470,N_9007);
nor U10791 (N_10791,N_9819,N_9704);
nand U10792 (N_10792,N_9732,N_9354);
or U10793 (N_10793,N_9654,N_9796);
nor U10794 (N_10794,N_9470,N_9962);
nand U10795 (N_10795,N_9757,N_9583);
or U10796 (N_10796,N_9641,N_9054);
or U10797 (N_10797,N_9882,N_9555);
xnor U10798 (N_10798,N_9993,N_9595);
or U10799 (N_10799,N_9350,N_9292);
xnor U10800 (N_10800,N_9695,N_9182);
nor U10801 (N_10801,N_9439,N_9533);
nor U10802 (N_10802,N_9502,N_9135);
and U10803 (N_10803,N_9708,N_9667);
and U10804 (N_10804,N_9767,N_9766);
or U10805 (N_10805,N_9239,N_9696);
or U10806 (N_10806,N_9316,N_9804);
xor U10807 (N_10807,N_9004,N_9038);
nand U10808 (N_10808,N_9037,N_9266);
nor U10809 (N_10809,N_9937,N_9555);
or U10810 (N_10810,N_9587,N_9236);
and U10811 (N_10811,N_9502,N_9713);
nand U10812 (N_10812,N_9590,N_9474);
and U10813 (N_10813,N_9182,N_9034);
xor U10814 (N_10814,N_9873,N_9483);
nor U10815 (N_10815,N_9066,N_9229);
nand U10816 (N_10816,N_9458,N_9755);
nor U10817 (N_10817,N_9727,N_9160);
nor U10818 (N_10818,N_9196,N_9782);
nor U10819 (N_10819,N_9191,N_9394);
nand U10820 (N_10820,N_9521,N_9196);
and U10821 (N_10821,N_9179,N_9454);
and U10822 (N_10822,N_9949,N_9197);
or U10823 (N_10823,N_9174,N_9022);
nor U10824 (N_10824,N_9640,N_9987);
or U10825 (N_10825,N_9921,N_9373);
nor U10826 (N_10826,N_9225,N_9581);
nand U10827 (N_10827,N_9634,N_9306);
xnor U10828 (N_10828,N_9777,N_9705);
nand U10829 (N_10829,N_9767,N_9317);
nand U10830 (N_10830,N_9939,N_9766);
or U10831 (N_10831,N_9514,N_9239);
nor U10832 (N_10832,N_9393,N_9502);
nor U10833 (N_10833,N_9336,N_9190);
xnor U10834 (N_10834,N_9078,N_9247);
and U10835 (N_10835,N_9061,N_9698);
or U10836 (N_10836,N_9243,N_9366);
or U10837 (N_10837,N_9549,N_9618);
and U10838 (N_10838,N_9161,N_9748);
and U10839 (N_10839,N_9691,N_9872);
or U10840 (N_10840,N_9348,N_9613);
xor U10841 (N_10841,N_9754,N_9498);
or U10842 (N_10842,N_9894,N_9286);
and U10843 (N_10843,N_9061,N_9592);
and U10844 (N_10844,N_9570,N_9474);
nand U10845 (N_10845,N_9573,N_9928);
nor U10846 (N_10846,N_9641,N_9440);
and U10847 (N_10847,N_9285,N_9597);
nand U10848 (N_10848,N_9830,N_9367);
or U10849 (N_10849,N_9398,N_9152);
nand U10850 (N_10850,N_9835,N_9769);
nand U10851 (N_10851,N_9881,N_9845);
or U10852 (N_10852,N_9377,N_9977);
xnor U10853 (N_10853,N_9669,N_9734);
and U10854 (N_10854,N_9536,N_9238);
nand U10855 (N_10855,N_9975,N_9991);
and U10856 (N_10856,N_9749,N_9022);
nor U10857 (N_10857,N_9664,N_9731);
nand U10858 (N_10858,N_9252,N_9288);
nand U10859 (N_10859,N_9564,N_9212);
xor U10860 (N_10860,N_9584,N_9248);
xnor U10861 (N_10861,N_9481,N_9486);
and U10862 (N_10862,N_9522,N_9967);
nor U10863 (N_10863,N_9733,N_9477);
nor U10864 (N_10864,N_9950,N_9438);
xnor U10865 (N_10865,N_9108,N_9316);
and U10866 (N_10866,N_9457,N_9731);
nor U10867 (N_10867,N_9152,N_9543);
nand U10868 (N_10868,N_9968,N_9160);
or U10869 (N_10869,N_9241,N_9291);
nand U10870 (N_10870,N_9667,N_9545);
nor U10871 (N_10871,N_9440,N_9471);
nand U10872 (N_10872,N_9322,N_9626);
xor U10873 (N_10873,N_9434,N_9089);
or U10874 (N_10874,N_9552,N_9753);
nand U10875 (N_10875,N_9696,N_9599);
nor U10876 (N_10876,N_9236,N_9890);
xor U10877 (N_10877,N_9259,N_9022);
and U10878 (N_10878,N_9916,N_9959);
and U10879 (N_10879,N_9372,N_9760);
nand U10880 (N_10880,N_9430,N_9978);
xnor U10881 (N_10881,N_9886,N_9048);
nor U10882 (N_10882,N_9029,N_9900);
nand U10883 (N_10883,N_9769,N_9404);
xnor U10884 (N_10884,N_9179,N_9762);
or U10885 (N_10885,N_9230,N_9236);
nand U10886 (N_10886,N_9427,N_9498);
or U10887 (N_10887,N_9175,N_9098);
and U10888 (N_10888,N_9090,N_9468);
nor U10889 (N_10889,N_9226,N_9861);
xor U10890 (N_10890,N_9034,N_9639);
nor U10891 (N_10891,N_9184,N_9261);
nor U10892 (N_10892,N_9077,N_9842);
or U10893 (N_10893,N_9951,N_9932);
or U10894 (N_10894,N_9734,N_9352);
and U10895 (N_10895,N_9174,N_9445);
nor U10896 (N_10896,N_9549,N_9467);
nand U10897 (N_10897,N_9708,N_9007);
and U10898 (N_10898,N_9963,N_9155);
nand U10899 (N_10899,N_9785,N_9475);
nor U10900 (N_10900,N_9296,N_9994);
nor U10901 (N_10901,N_9666,N_9224);
and U10902 (N_10902,N_9553,N_9772);
nor U10903 (N_10903,N_9729,N_9442);
nand U10904 (N_10904,N_9525,N_9278);
or U10905 (N_10905,N_9920,N_9225);
nand U10906 (N_10906,N_9269,N_9645);
and U10907 (N_10907,N_9147,N_9279);
nor U10908 (N_10908,N_9705,N_9515);
nand U10909 (N_10909,N_9487,N_9822);
nor U10910 (N_10910,N_9483,N_9010);
nand U10911 (N_10911,N_9624,N_9400);
or U10912 (N_10912,N_9941,N_9044);
or U10913 (N_10913,N_9133,N_9462);
nor U10914 (N_10914,N_9419,N_9494);
nor U10915 (N_10915,N_9549,N_9196);
nor U10916 (N_10916,N_9806,N_9395);
and U10917 (N_10917,N_9173,N_9066);
or U10918 (N_10918,N_9152,N_9613);
and U10919 (N_10919,N_9095,N_9967);
nand U10920 (N_10920,N_9980,N_9933);
and U10921 (N_10921,N_9796,N_9167);
nor U10922 (N_10922,N_9308,N_9237);
xor U10923 (N_10923,N_9328,N_9027);
nand U10924 (N_10924,N_9094,N_9926);
and U10925 (N_10925,N_9069,N_9484);
xor U10926 (N_10926,N_9542,N_9737);
and U10927 (N_10927,N_9728,N_9898);
xnor U10928 (N_10928,N_9591,N_9873);
xnor U10929 (N_10929,N_9456,N_9971);
nand U10930 (N_10930,N_9291,N_9205);
or U10931 (N_10931,N_9526,N_9283);
nor U10932 (N_10932,N_9150,N_9000);
nor U10933 (N_10933,N_9181,N_9690);
nand U10934 (N_10934,N_9145,N_9685);
and U10935 (N_10935,N_9102,N_9018);
nand U10936 (N_10936,N_9575,N_9370);
and U10937 (N_10937,N_9981,N_9304);
nand U10938 (N_10938,N_9808,N_9908);
or U10939 (N_10939,N_9210,N_9877);
or U10940 (N_10940,N_9393,N_9423);
nand U10941 (N_10941,N_9925,N_9992);
and U10942 (N_10942,N_9545,N_9275);
and U10943 (N_10943,N_9660,N_9586);
xor U10944 (N_10944,N_9732,N_9231);
nor U10945 (N_10945,N_9567,N_9938);
xor U10946 (N_10946,N_9513,N_9497);
and U10947 (N_10947,N_9494,N_9541);
and U10948 (N_10948,N_9618,N_9960);
nor U10949 (N_10949,N_9402,N_9280);
or U10950 (N_10950,N_9578,N_9168);
nand U10951 (N_10951,N_9862,N_9173);
xnor U10952 (N_10952,N_9454,N_9880);
nor U10953 (N_10953,N_9453,N_9449);
nand U10954 (N_10954,N_9583,N_9707);
xor U10955 (N_10955,N_9757,N_9657);
xnor U10956 (N_10956,N_9186,N_9397);
nor U10957 (N_10957,N_9920,N_9145);
and U10958 (N_10958,N_9982,N_9079);
or U10959 (N_10959,N_9081,N_9314);
nor U10960 (N_10960,N_9509,N_9043);
or U10961 (N_10961,N_9156,N_9651);
and U10962 (N_10962,N_9403,N_9690);
nor U10963 (N_10963,N_9521,N_9416);
xnor U10964 (N_10964,N_9019,N_9849);
nand U10965 (N_10965,N_9967,N_9048);
and U10966 (N_10966,N_9748,N_9823);
nor U10967 (N_10967,N_9955,N_9947);
nor U10968 (N_10968,N_9173,N_9407);
nand U10969 (N_10969,N_9716,N_9167);
or U10970 (N_10970,N_9747,N_9799);
nor U10971 (N_10971,N_9723,N_9937);
nand U10972 (N_10972,N_9486,N_9049);
nand U10973 (N_10973,N_9885,N_9538);
xnor U10974 (N_10974,N_9752,N_9075);
and U10975 (N_10975,N_9658,N_9871);
xnor U10976 (N_10976,N_9345,N_9907);
or U10977 (N_10977,N_9436,N_9171);
xor U10978 (N_10978,N_9304,N_9023);
and U10979 (N_10979,N_9898,N_9278);
or U10980 (N_10980,N_9812,N_9206);
or U10981 (N_10981,N_9457,N_9585);
nand U10982 (N_10982,N_9060,N_9295);
xor U10983 (N_10983,N_9062,N_9784);
nor U10984 (N_10984,N_9904,N_9827);
nor U10985 (N_10985,N_9144,N_9558);
nand U10986 (N_10986,N_9913,N_9645);
xnor U10987 (N_10987,N_9566,N_9156);
nor U10988 (N_10988,N_9176,N_9220);
xor U10989 (N_10989,N_9811,N_9721);
and U10990 (N_10990,N_9035,N_9013);
nand U10991 (N_10991,N_9482,N_9208);
xnor U10992 (N_10992,N_9739,N_9141);
or U10993 (N_10993,N_9781,N_9913);
nor U10994 (N_10994,N_9005,N_9197);
nor U10995 (N_10995,N_9086,N_9337);
nand U10996 (N_10996,N_9605,N_9841);
or U10997 (N_10997,N_9480,N_9848);
xnor U10998 (N_10998,N_9179,N_9992);
and U10999 (N_10999,N_9289,N_9997);
or U11000 (N_11000,N_10764,N_10378);
nand U11001 (N_11001,N_10507,N_10663);
or U11002 (N_11002,N_10173,N_10226);
xnor U11003 (N_11003,N_10686,N_10315);
or U11004 (N_11004,N_10842,N_10558);
nor U11005 (N_11005,N_10871,N_10009);
xnor U11006 (N_11006,N_10598,N_10903);
or U11007 (N_11007,N_10697,N_10603);
and U11008 (N_11008,N_10153,N_10918);
xor U11009 (N_11009,N_10896,N_10347);
nand U11010 (N_11010,N_10829,N_10181);
and U11011 (N_11011,N_10374,N_10515);
xor U11012 (N_11012,N_10149,N_10152);
or U11013 (N_11013,N_10617,N_10502);
xnor U11014 (N_11014,N_10519,N_10214);
or U11015 (N_11015,N_10293,N_10339);
nor U11016 (N_11016,N_10823,N_10301);
and U11017 (N_11017,N_10593,N_10092);
nor U11018 (N_11018,N_10760,N_10360);
nand U11019 (N_11019,N_10338,N_10795);
nor U11020 (N_11020,N_10292,N_10522);
nor U11021 (N_11021,N_10583,N_10483);
and U11022 (N_11022,N_10727,N_10754);
or U11023 (N_11023,N_10341,N_10404);
xnor U11024 (N_11024,N_10366,N_10545);
xnor U11025 (N_11025,N_10131,N_10704);
or U11026 (N_11026,N_10731,N_10856);
or U11027 (N_11027,N_10385,N_10066);
nand U11028 (N_11028,N_10860,N_10208);
nor U11029 (N_11029,N_10223,N_10628);
or U11030 (N_11030,N_10201,N_10450);
or U11031 (N_11031,N_10845,N_10257);
or U11032 (N_11032,N_10677,N_10839);
nor U11033 (N_11033,N_10655,N_10342);
xnor U11034 (N_11034,N_10662,N_10915);
nor U11035 (N_11035,N_10249,N_10157);
or U11036 (N_11036,N_10565,N_10716);
nor U11037 (N_11037,N_10998,N_10863);
or U11038 (N_11038,N_10970,N_10984);
nand U11039 (N_11039,N_10571,N_10891);
nor U11040 (N_11040,N_10098,N_10321);
xnor U11041 (N_11041,N_10544,N_10075);
nand U11042 (N_11042,N_10311,N_10755);
or U11043 (N_11043,N_10403,N_10297);
nor U11044 (N_11044,N_10552,N_10804);
nand U11045 (N_11045,N_10095,N_10592);
xor U11046 (N_11046,N_10160,N_10955);
nand U11047 (N_11047,N_10254,N_10702);
nand U11048 (N_11048,N_10721,N_10904);
nand U11049 (N_11049,N_10947,N_10049);
nor U11050 (N_11050,N_10921,N_10635);
xor U11051 (N_11051,N_10966,N_10166);
nand U11052 (N_11052,N_10954,N_10642);
xor U11053 (N_11053,N_10849,N_10137);
or U11054 (N_11054,N_10022,N_10770);
or U11055 (N_11055,N_10456,N_10114);
nor U11056 (N_11056,N_10340,N_10855);
nor U11057 (N_11057,N_10211,N_10521);
and U11058 (N_11058,N_10975,N_10281);
nor U11059 (N_11059,N_10085,N_10619);
and U11060 (N_11060,N_10523,N_10818);
xnor U11061 (N_11061,N_10467,N_10768);
or U11062 (N_11062,N_10783,N_10636);
nor U11063 (N_11063,N_10255,N_10806);
and U11064 (N_11064,N_10553,N_10561);
nor U11065 (N_11065,N_10854,N_10132);
nor U11066 (N_11066,N_10123,N_10365);
xor U11067 (N_11067,N_10928,N_10825);
nor U11068 (N_11068,N_10604,N_10122);
xor U11069 (N_11069,N_10639,N_10399);
or U11070 (N_11070,N_10878,N_10511);
and U11071 (N_11071,N_10527,N_10786);
or U11072 (N_11072,N_10792,N_10684);
or U11073 (N_11073,N_10127,N_10685);
or U11074 (N_11074,N_10933,N_10911);
xnor U11075 (N_11075,N_10720,N_10660);
xnor U11076 (N_11076,N_10275,N_10950);
nand U11077 (N_11077,N_10186,N_10784);
or U11078 (N_11078,N_10352,N_10364);
or U11079 (N_11079,N_10269,N_10124);
xor U11080 (N_11080,N_10278,N_10081);
or U11081 (N_11081,N_10838,N_10291);
xnor U11082 (N_11082,N_10750,N_10045);
nand U11083 (N_11083,N_10048,N_10828);
nor U11084 (N_11084,N_10840,N_10566);
nand U11085 (N_11085,N_10105,N_10977);
or U11086 (N_11086,N_10451,N_10802);
or U11087 (N_11087,N_10890,N_10986);
nand U11088 (N_11088,N_10219,N_10960);
xnor U11089 (N_11089,N_10925,N_10886);
or U11090 (N_11090,N_10224,N_10433);
xnor U11091 (N_11091,N_10622,N_10021);
nand U11092 (N_11092,N_10674,N_10963);
xnor U11093 (N_11093,N_10446,N_10876);
xnor U11094 (N_11094,N_10514,N_10041);
nor U11095 (N_11095,N_10725,N_10334);
xnor U11096 (N_11096,N_10992,N_10455);
xnor U11097 (N_11097,N_10052,N_10314);
nor U11098 (N_11098,N_10099,N_10490);
nand U11099 (N_11099,N_10386,N_10030);
xor U11100 (N_11100,N_10423,N_10040);
and U11101 (N_11101,N_10333,N_10110);
nor U11102 (N_11102,N_10047,N_10262);
xor U11103 (N_11103,N_10466,N_10007);
and U11104 (N_11104,N_10656,N_10017);
and U11105 (N_11105,N_10962,N_10349);
nor U11106 (N_11106,N_10002,N_10665);
nor U11107 (N_11107,N_10145,N_10746);
and U11108 (N_11108,N_10393,N_10469);
or U11109 (N_11109,N_10621,N_10689);
nor U11110 (N_11110,N_10343,N_10348);
xnor U11111 (N_11111,N_10882,N_10695);
or U11112 (N_11112,N_10889,N_10816);
or U11113 (N_11113,N_10372,N_10381);
xnor U11114 (N_11114,N_10234,N_10189);
nor U11115 (N_11115,N_10406,N_10805);
and U11116 (N_11116,N_10948,N_10586);
xor U11117 (N_11117,N_10134,N_10946);
nor U11118 (N_11118,N_10533,N_10217);
nand U11119 (N_11119,N_10144,N_10481);
nor U11120 (N_11120,N_10879,N_10452);
xor U11121 (N_11121,N_10569,N_10215);
or U11122 (N_11122,N_10271,N_10958);
and U11123 (N_11123,N_10841,N_10135);
or U11124 (N_11124,N_10999,N_10243);
and U11125 (N_11125,N_10859,N_10119);
or U11126 (N_11126,N_10222,N_10492);
nor U11127 (N_11127,N_10159,N_10791);
nand U11128 (N_11128,N_10267,N_10408);
or U11129 (N_11129,N_10726,N_10705);
nor U11130 (N_11130,N_10298,N_10923);
nor U11131 (N_11131,N_10165,N_10638);
nor U11132 (N_11132,N_10542,N_10560);
or U11133 (N_11133,N_10733,N_10453);
and U11134 (N_11134,N_10847,N_10432);
nor U11135 (N_11135,N_10060,N_10988);
and U11136 (N_11136,N_10125,N_10761);
nand U11137 (N_11137,N_10648,N_10053);
or U11138 (N_11138,N_10897,N_10439);
nand U11139 (N_11139,N_10064,N_10086);
nor U11140 (N_11140,N_10182,N_10277);
xnor U11141 (N_11141,N_10901,N_10202);
and U11142 (N_11142,N_10163,N_10945);
and U11143 (N_11143,N_10518,N_10073);
xnor U11144 (N_11144,N_10104,N_10463);
or U11145 (N_11145,N_10100,N_10737);
nor U11146 (N_11146,N_10611,N_10525);
and U11147 (N_11147,N_10205,N_10212);
nor U11148 (N_11148,N_10517,N_10344);
and U11149 (N_11149,N_10461,N_10813);
xor U11150 (N_11150,N_10059,N_10142);
and U11151 (N_11151,N_10738,N_10943);
and U11152 (N_11152,N_10034,N_10155);
nand U11153 (N_11153,N_10116,N_10097);
or U11154 (N_11154,N_10907,N_10713);
nor U11155 (N_11155,N_10014,N_10076);
and U11156 (N_11156,N_10357,N_10494);
and U11157 (N_11157,N_10614,N_10834);
and U11158 (N_11158,N_10358,N_10150);
and U11159 (N_11159,N_10539,N_10169);
nand U11160 (N_11160,N_10646,N_10640);
nand U11161 (N_11161,N_10032,N_10887);
xnor U11162 (N_11162,N_10115,N_10995);
xor U11163 (N_11163,N_10884,N_10682);
or U11164 (N_11164,N_10661,N_10843);
nor U11165 (N_11165,N_10102,N_10071);
and U11166 (N_11166,N_10599,N_10734);
xor U11167 (N_11167,N_10745,N_10557);
or U11168 (N_11168,N_10128,N_10930);
xor U11169 (N_11169,N_10026,N_10996);
and U11170 (N_11170,N_10464,N_10039);
nor U11171 (N_11171,N_10801,N_10965);
or U11172 (N_11172,N_10307,N_10337);
nor U11173 (N_11173,N_10024,N_10562);
or U11174 (N_11174,N_10350,N_10934);
and U11175 (N_11175,N_10810,N_10020);
nand U11176 (N_11176,N_10659,N_10238);
and U11177 (N_11177,N_10289,N_10380);
nand U11178 (N_11178,N_10940,N_10579);
nor U11179 (N_11179,N_10596,N_10916);
nor U11180 (N_11180,N_10260,N_10192);
xnor U11181 (N_11181,N_10894,N_10367);
or U11182 (N_11182,N_10506,N_10536);
nor U11183 (N_11183,N_10303,N_10322);
or U11184 (N_11184,N_10430,N_10781);
nor U11185 (N_11185,N_10213,N_10793);
or U11186 (N_11186,N_10538,N_10417);
nand U11187 (N_11187,N_10835,N_10241);
or U11188 (N_11188,N_10748,N_10990);
nand U11189 (N_11189,N_10779,N_10209);
nand U11190 (N_11190,N_10531,N_10497);
and U11191 (N_11191,N_10005,N_10714);
xor U11192 (N_11192,N_10833,N_10447);
xnor U11193 (N_11193,N_10844,N_10265);
or U11194 (N_11194,N_10759,N_10831);
or U11195 (N_11195,N_10090,N_10185);
nor U11196 (N_11196,N_10459,N_10325);
xor U11197 (N_11197,N_10078,N_10851);
and U11198 (N_11198,N_10023,N_10126);
or U11199 (N_11199,N_10610,N_10753);
nand U11200 (N_11200,N_10836,N_10698);
nor U11201 (N_11201,N_10174,N_10796);
nand U11202 (N_11202,N_10729,N_10820);
nand U11203 (N_11203,N_10625,N_10161);
and U11204 (N_11204,N_10089,N_10535);
nand U11205 (N_11205,N_10711,N_10900);
nand U11206 (N_11206,N_10763,N_10093);
or U11207 (N_11207,N_10072,N_10111);
nand U11208 (N_11208,N_10549,N_10425);
nor U11209 (N_11209,N_10196,N_10935);
or U11210 (N_11210,N_10266,N_10862);
or U11211 (N_11211,N_10304,N_10667);
and U11212 (N_11212,N_10826,N_10058);
or U11213 (N_11213,N_10458,N_10248);
nand U11214 (N_11214,N_10246,N_10206);
nand U11215 (N_11215,N_10151,N_10789);
xnor U11216 (N_11216,N_10392,N_10120);
and U11217 (N_11217,N_10312,N_10285);
xnor U11218 (N_11218,N_10171,N_10487);
nand U11219 (N_11219,N_10382,N_10440);
nor U11220 (N_11220,N_10817,N_10268);
xor U11221 (N_11221,N_10431,N_10396);
nand U11222 (N_11222,N_10905,N_10832);
or U11223 (N_11223,N_10136,N_10567);
or U11224 (N_11224,N_10573,N_10630);
xnor U11225 (N_11225,N_10225,N_10585);
xor U11226 (N_11226,N_10387,N_10830);
xnor U11227 (N_11227,N_10680,N_10693);
and U11228 (N_11228,N_10936,N_10468);
nor U11229 (N_11229,N_10724,N_10790);
nand U11230 (N_11230,N_10143,N_10473);
nor U11231 (N_11231,N_10096,N_10669);
and U11232 (N_11232,N_10575,N_10769);
or U11233 (N_11233,N_10077,N_10233);
xor U11234 (N_11234,N_10274,N_10997);
nor U11235 (N_11235,N_10436,N_10356);
and U11236 (N_11236,N_10036,N_10867);
or U11237 (N_11237,N_10156,N_10013);
xor U11238 (N_11238,N_10426,N_10974);
nand U11239 (N_11239,N_10589,N_10778);
and U11240 (N_11240,N_10554,N_10270);
nand U11241 (N_11241,N_10637,N_10808);
nor U11242 (N_11242,N_10324,N_10400);
and U11243 (N_11243,N_10472,N_10551);
and U11244 (N_11244,N_10141,N_10158);
xnor U11245 (N_11245,N_10003,N_10164);
or U11246 (N_11246,N_10253,N_10133);
nand U11247 (N_11247,N_10079,N_10488);
or U11248 (N_11248,N_10602,N_10564);
and U11249 (N_11249,N_10620,N_10411);
and U11250 (N_11250,N_10687,N_10016);
and U11251 (N_11251,N_10728,N_10991);
or U11252 (N_11252,N_10025,N_10240);
or U11253 (N_11253,N_10751,N_10814);
and U11254 (N_11254,N_10658,N_10956);
and U11255 (N_11255,N_10187,N_10489);
or U11256 (N_11256,N_10994,N_10305);
nand U11257 (N_11257,N_10606,N_10063);
and U11258 (N_11258,N_10065,N_10074);
nand U11259 (N_11259,N_10649,N_10615);
nand U11260 (N_11260,N_10788,N_10474);
and U11261 (N_11261,N_10207,N_10528);
or U11262 (N_11262,N_10252,N_10730);
nand U11263 (N_11263,N_10942,N_10908);
nand U11264 (N_11264,N_10388,N_10037);
nor U11265 (N_11265,N_10979,N_10537);
xnor U11266 (N_11266,N_10824,N_10982);
xor U11267 (N_11267,N_10435,N_10971);
and U11268 (N_11268,N_10967,N_10251);
nand U11269 (N_11269,N_10676,N_10794);
or U11270 (N_11270,N_10410,N_10652);
or U11271 (N_11271,N_10087,N_10631);
nor U11272 (N_11272,N_10771,N_10609);
xnor U11273 (N_11273,N_10046,N_10191);
xnor U11274 (N_11274,N_10195,N_10235);
and U11275 (N_11275,N_10895,N_10595);
and U11276 (N_11276,N_10326,N_10300);
xor U11277 (N_11277,N_10499,N_10320);
nand U11278 (N_11278,N_10188,N_10370);
and U11279 (N_11279,N_10740,N_10263);
xnor U11280 (N_11280,N_10412,N_10616);
xnor U11281 (N_11281,N_10563,N_10503);
xor U11282 (N_11282,N_10148,N_10688);
nand U11283 (N_11283,N_10645,N_10922);
xor U11284 (N_11284,N_10938,N_10375);
and U11285 (N_11285,N_10837,N_10194);
xor U11286 (N_11286,N_10752,N_10772);
and U11287 (N_11287,N_10443,N_10397);
and U11288 (N_11288,N_10172,N_10944);
and U11289 (N_11289,N_10371,N_10821);
and U11290 (N_11290,N_10363,N_10739);
nand U11291 (N_11291,N_10556,N_10327);
or U11292 (N_11292,N_10989,N_10480);
nand U11293 (N_11293,N_10780,N_10866);
nand U11294 (N_11294,N_10401,N_10287);
or U11295 (N_11295,N_10785,N_10774);
and U11296 (N_11296,N_10283,N_10228);
and U11297 (N_11297,N_10787,N_10256);
nand U11298 (N_11298,N_10106,N_10766);
and U11299 (N_11299,N_10941,N_10437);
nand U11300 (N_11300,N_10310,N_10103);
or U11301 (N_11301,N_10546,N_10179);
and U11302 (N_11302,N_10203,N_10949);
xnor U11303 (N_11303,N_10968,N_10978);
nand U11304 (N_11304,N_10718,N_10330);
xor U11305 (N_11305,N_10284,N_10782);
or U11306 (N_11306,N_10345,N_10001);
nand U11307 (N_11307,N_10758,N_10743);
or U11308 (N_11308,N_10011,N_10861);
xor U11309 (N_11309,N_10885,N_10449);
or U11310 (N_11310,N_10694,N_10543);
xor U11311 (N_11311,N_10715,N_10247);
nor U11312 (N_11312,N_10245,N_10709);
and U11313 (N_11313,N_10657,N_10302);
nor U11314 (N_11314,N_10394,N_10541);
or U11315 (N_11315,N_10383,N_10741);
nor U11316 (N_11316,N_10259,N_10445);
xor U11317 (N_11317,N_10094,N_10218);
xor U11318 (N_11318,N_10038,N_10883);
and U11319 (N_11319,N_10578,N_10633);
xnor U11320 (N_11320,N_10776,N_10199);
and U11321 (N_11321,N_10762,N_10434);
or U11322 (N_11322,N_10624,N_10336);
nand U11323 (N_11323,N_10368,N_10476);
and U11324 (N_11324,N_10873,N_10594);
nor U11325 (N_11325,N_10416,N_10475);
nand U11326 (N_11326,N_10316,N_10204);
xnor U11327 (N_11327,N_10484,N_10675);
or U11328 (N_11328,N_10932,N_10902);
or U11329 (N_11329,N_10398,N_10373);
xnor U11330 (N_11330,N_10520,N_10613);
nand U11331 (N_11331,N_10717,N_10909);
nor U11332 (N_11332,N_10323,N_10872);
nand U11333 (N_11333,N_10898,N_10441);
and U11334 (N_11334,N_10061,N_10421);
or U11335 (N_11335,N_10130,N_10221);
xnor U11336 (N_11336,N_10912,N_10951);
nand U11337 (N_11337,N_10454,N_10299);
nand U11338 (N_11338,N_10550,N_10679);
or U11339 (N_11339,N_10588,N_10354);
and U11340 (N_11340,N_10193,N_10146);
nor U11341 (N_11341,N_10118,N_10177);
or U11342 (N_11342,N_10331,N_10953);
nand U11343 (N_11343,N_10290,N_10019);
nand U11344 (N_11344,N_10634,N_10462);
nand U11345 (N_11345,N_10570,N_10852);
and U11346 (N_11346,N_10369,N_10722);
or U11347 (N_11347,N_10815,N_10422);
and U11348 (N_11348,N_10083,N_10629);
nand U11349 (N_11349,N_10710,N_10236);
and U11350 (N_11350,N_10027,N_10627);
nor U11351 (N_11351,N_10910,N_10471);
or U11352 (N_11352,N_10532,N_10892);
xor U11353 (N_11353,N_10309,N_10757);
and U11354 (N_11354,N_10670,N_10961);
nor U11355 (N_11355,N_10590,N_10424);
nor U11356 (N_11356,N_10107,N_10210);
xor U11357 (N_11357,N_10505,N_10666);
nand U11358 (N_11358,N_10632,N_10395);
or U11359 (N_11359,N_10597,N_10198);
nand U11360 (N_11360,N_10881,N_10389);
nor U11361 (N_11361,N_10442,N_10308);
or U11362 (N_11362,N_10109,N_10332);
or U11363 (N_11363,N_10362,N_10485);
and U11364 (N_11364,N_10848,N_10390);
nand U11365 (N_11365,N_10313,N_10707);
nor U11366 (N_11366,N_10460,N_10244);
or U11367 (N_11367,N_10318,N_10591);
nor U11368 (N_11368,N_10568,N_10651);
and U11369 (N_11369,N_10601,N_10671);
xnor U11370 (N_11370,N_10138,N_10242);
nor U11371 (N_11371,N_10827,N_10800);
and U11372 (N_11372,N_10623,N_10108);
nand U11373 (N_11373,N_10712,N_10587);
or U11374 (N_11374,N_10976,N_10574);
xnor U11375 (N_11375,N_10858,N_10927);
nand U11376 (N_11376,N_10555,N_10919);
nand U11377 (N_11377,N_10029,N_10470);
or U11378 (N_11378,N_10015,N_10703);
nor U11379 (N_11379,N_10807,N_10673);
nand U11380 (N_11380,N_10981,N_10701);
nor U11381 (N_11381,N_10069,N_10280);
and U11382 (N_11382,N_10924,N_10050);
nand U11383 (N_11383,N_10735,N_10811);
and U11384 (N_11384,N_10668,N_10317);
and U11385 (N_11385,N_10272,N_10384);
xor U11386 (N_11386,N_10875,N_10584);
xnor U11387 (N_11387,N_10168,N_10121);
or U11388 (N_11388,N_10082,N_10361);
or U11389 (N_11389,N_10870,N_10690);
nand U11390 (N_11390,N_10319,N_10438);
and U11391 (N_11391,N_10865,N_10819);
xnor U11392 (N_11392,N_10864,N_10605);
or U11393 (N_11393,N_10524,N_10167);
xnor U11394 (N_11394,N_10732,N_10767);
nand U11395 (N_11395,N_10008,N_10959);
nor U11396 (N_11396,N_10427,N_10409);
or U11397 (N_11397,N_10929,N_10062);
xor U11398 (N_11398,N_10719,N_10190);
xor U11399 (N_11399,N_10985,N_10258);
nand U11400 (N_11400,N_10798,N_10035);
nand U11401 (N_11401,N_10056,N_10175);
xor U11402 (N_11402,N_10877,N_10006);
or U11403 (N_11403,N_10812,N_10391);
xor U11404 (N_11404,N_10282,N_10288);
and U11405 (N_11405,N_10154,N_10512);
and U11406 (N_11406,N_10612,N_10581);
xnor U11407 (N_11407,N_10033,N_10747);
nor U11408 (N_11408,N_10868,N_10180);
nand U11409 (N_11409,N_10799,N_10080);
nand U11410 (N_11410,N_10850,N_10526);
nand U11411 (N_11411,N_10377,N_10012);
nand U11412 (N_11412,N_10803,N_10893);
nor U11413 (N_11413,N_10482,N_10147);
or U11414 (N_11414,N_10335,N_10231);
xor U11415 (N_11415,N_10067,N_10448);
nor U11416 (N_11416,N_10286,N_10736);
nand U11417 (N_11417,N_10491,N_10140);
or U11418 (N_11418,N_10678,N_10742);
and U11419 (N_11419,N_10232,N_10580);
and U11420 (N_11420,N_10683,N_10402);
and U11421 (N_11421,N_10899,N_10869);
or U11422 (N_11422,N_10576,N_10913);
or U11423 (N_11423,N_10920,N_10846);
nand U11424 (N_11424,N_10917,N_10969);
xor U11425 (N_11425,N_10261,N_10444);
xnor U11426 (N_11426,N_10200,N_10641);
nand U11427 (N_11427,N_10723,N_10279);
or U11428 (N_11428,N_10972,N_10529);
nor U11429 (N_11429,N_10765,N_10486);
nand U11430 (N_11430,N_10376,N_10479);
nand U11431 (N_11431,N_10429,N_10239);
nor U11432 (N_11432,N_10043,N_10559);
and U11433 (N_11433,N_10773,N_10777);
nor U11434 (N_11434,N_10306,N_10647);
or U11435 (N_11435,N_10170,N_10407);
nor U11436 (N_11436,N_10744,N_10496);
and U11437 (N_11437,N_10184,N_10644);
nand U11438 (N_11438,N_10477,N_10548);
xor U11439 (N_11439,N_10057,N_10672);
and U11440 (N_11440,N_10084,N_10346);
nor U11441 (N_11441,N_10493,N_10540);
nor U11442 (N_11442,N_10295,N_10504);
nand U11443 (N_11443,N_10993,N_10508);
nor U11444 (N_11444,N_10822,N_10428);
nor U11445 (N_11445,N_10054,N_10415);
nand U11446 (N_11446,N_10607,N_10534);
or U11447 (N_11447,N_10572,N_10117);
nand U11448 (N_11448,N_10220,N_10857);
nand U11449 (N_11449,N_10957,N_10113);
or U11450 (N_11450,N_10414,N_10926);
and U11451 (N_11451,N_10987,N_10042);
xnor U11452 (N_11452,N_10413,N_10973);
nor U11453 (N_11453,N_10510,N_10355);
nor U11454 (N_11454,N_10706,N_10691);
nand U11455 (N_11455,N_10088,N_10010);
nand U11456 (N_11456,N_10353,N_10906);
nor U11457 (N_11457,N_10952,N_10276);
and U11458 (N_11458,N_10654,N_10178);
nor U11459 (N_11459,N_10931,N_10643);
xnor U11460 (N_11460,N_10070,N_10708);
xnor U11461 (N_11461,N_10500,N_10797);
nor U11462 (N_11462,N_10650,N_10880);
nand U11463 (N_11463,N_10964,N_10516);
nand U11464 (N_11464,N_10419,N_10914);
or U11465 (N_11465,N_10176,N_10101);
or U11466 (N_11466,N_10068,N_10756);
nand U11467 (N_11467,N_10618,N_10051);
or U11468 (N_11468,N_10749,N_10980);
and U11469 (N_11469,N_10229,N_10582);
nor U11470 (N_11470,N_10465,N_10939);
and U11471 (N_11471,N_10983,N_10264);
nor U11472 (N_11472,N_10055,N_10273);
or U11473 (N_11473,N_10328,N_10608);
xnor U11474 (N_11474,N_10457,N_10937);
nor U11475 (N_11475,N_10139,N_10162);
xor U11476 (N_11476,N_10031,N_10004);
xor U11477 (N_11477,N_10513,N_10018);
or U11478 (N_11478,N_10809,N_10028);
nand U11479 (N_11479,N_10044,N_10509);
xnor U11480 (N_11480,N_10183,N_10495);
or U11481 (N_11481,N_10501,N_10653);
and U11482 (N_11482,N_10418,N_10664);
and U11483 (N_11483,N_10091,N_10112);
nand U11484 (N_11484,N_10478,N_10250);
xor U11485 (N_11485,N_10874,N_10329);
xnor U11486 (N_11486,N_10700,N_10530);
nor U11487 (N_11487,N_10129,N_10237);
or U11488 (N_11488,N_10600,N_10577);
nor U11489 (N_11489,N_10230,N_10692);
nand U11490 (N_11490,N_10197,N_10216);
or U11491 (N_11491,N_10000,N_10359);
and U11492 (N_11492,N_10294,N_10626);
nor U11493 (N_11493,N_10775,N_10227);
nor U11494 (N_11494,N_10547,N_10888);
nor U11495 (N_11495,N_10681,N_10405);
nand U11496 (N_11496,N_10853,N_10379);
nor U11497 (N_11497,N_10699,N_10420);
nand U11498 (N_11498,N_10696,N_10498);
xnor U11499 (N_11499,N_10296,N_10351);
or U11500 (N_11500,N_10675,N_10370);
xor U11501 (N_11501,N_10827,N_10945);
nor U11502 (N_11502,N_10911,N_10236);
or U11503 (N_11503,N_10528,N_10667);
nand U11504 (N_11504,N_10220,N_10661);
xnor U11505 (N_11505,N_10391,N_10134);
nand U11506 (N_11506,N_10651,N_10968);
nor U11507 (N_11507,N_10807,N_10402);
nor U11508 (N_11508,N_10015,N_10402);
nand U11509 (N_11509,N_10303,N_10310);
xnor U11510 (N_11510,N_10535,N_10326);
nor U11511 (N_11511,N_10289,N_10660);
and U11512 (N_11512,N_10623,N_10700);
and U11513 (N_11513,N_10337,N_10364);
and U11514 (N_11514,N_10477,N_10581);
xor U11515 (N_11515,N_10713,N_10383);
nand U11516 (N_11516,N_10713,N_10965);
nor U11517 (N_11517,N_10330,N_10115);
and U11518 (N_11518,N_10614,N_10021);
or U11519 (N_11519,N_10307,N_10474);
nand U11520 (N_11520,N_10930,N_10786);
nand U11521 (N_11521,N_10018,N_10264);
and U11522 (N_11522,N_10949,N_10657);
or U11523 (N_11523,N_10567,N_10353);
nand U11524 (N_11524,N_10820,N_10619);
xor U11525 (N_11525,N_10583,N_10611);
nand U11526 (N_11526,N_10778,N_10848);
nand U11527 (N_11527,N_10403,N_10220);
xor U11528 (N_11528,N_10783,N_10477);
xor U11529 (N_11529,N_10233,N_10934);
xor U11530 (N_11530,N_10112,N_10572);
nor U11531 (N_11531,N_10167,N_10518);
nand U11532 (N_11532,N_10098,N_10797);
nand U11533 (N_11533,N_10718,N_10884);
or U11534 (N_11534,N_10974,N_10236);
and U11535 (N_11535,N_10921,N_10374);
nand U11536 (N_11536,N_10686,N_10303);
nand U11537 (N_11537,N_10754,N_10732);
or U11538 (N_11538,N_10549,N_10516);
nor U11539 (N_11539,N_10249,N_10446);
nand U11540 (N_11540,N_10445,N_10239);
nor U11541 (N_11541,N_10627,N_10117);
xnor U11542 (N_11542,N_10609,N_10817);
or U11543 (N_11543,N_10580,N_10382);
nand U11544 (N_11544,N_10723,N_10106);
or U11545 (N_11545,N_10951,N_10200);
or U11546 (N_11546,N_10526,N_10418);
xor U11547 (N_11547,N_10364,N_10186);
nor U11548 (N_11548,N_10644,N_10099);
or U11549 (N_11549,N_10312,N_10479);
nand U11550 (N_11550,N_10510,N_10531);
nand U11551 (N_11551,N_10244,N_10645);
and U11552 (N_11552,N_10292,N_10990);
and U11553 (N_11553,N_10751,N_10244);
xnor U11554 (N_11554,N_10275,N_10116);
xnor U11555 (N_11555,N_10439,N_10450);
nor U11556 (N_11556,N_10083,N_10353);
nand U11557 (N_11557,N_10532,N_10082);
and U11558 (N_11558,N_10126,N_10029);
and U11559 (N_11559,N_10371,N_10670);
and U11560 (N_11560,N_10481,N_10764);
and U11561 (N_11561,N_10903,N_10546);
nand U11562 (N_11562,N_10267,N_10843);
nor U11563 (N_11563,N_10645,N_10841);
and U11564 (N_11564,N_10646,N_10756);
or U11565 (N_11565,N_10947,N_10304);
xnor U11566 (N_11566,N_10849,N_10194);
or U11567 (N_11567,N_10243,N_10573);
nor U11568 (N_11568,N_10658,N_10415);
or U11569 (N_11569,N_10621,N_10878);
or U11570 (N_11570,N_10070,N_10397);
and U11571 (N_11571,N_10277,N_10477);
nor U11572 (N_11572,N_10702,N_10884);
nand U11573 (N_11573,N_10283,N_10652);
and U11574 (N_11574,N_10839,N_10808);
and U11575 (N_11575,N_10221,N_10362);
and U11576 (N_11576,N_10033,N_10102);
nor U11577 (N_11577,N_10138,N_10264);
and U11578 (N_11578,N_10679,N_10886);
xor U11579 (N_11579,N_10450,N_10217);
nor U11580 (N_11580,N_10721,N_10092);
nand U11581 (N_11581,N_10535,N_10532);
nor U11582 (N_11582,N_10024,N_10512);
and U11583 (N_11583,N_10739,N_10072);
nand U11584 (N_11584,N_10402,N_10625);
nor U11585 (N_11585,N_10800,N_10619);
or U11586 (N_11586,N_10304,N_10518);
nor U11587 (N_11587,N_10233,N_10569);
or U11588 (N_11588,N_10266,N_10768);
or U11589 (N_11589,N_10483,N_10884);
nor U11590 (N_11590,N_10978,N_10515);
or U11591 (N_11591,N_10145,N_10797);
xor U11592 (N_11592,N_10500,N_10331);
nand U11593 (N_11593,N_10605,N_10485);
nand U11594 (N_11594,N_10572,N_10828);
nor U11595 (N_11595,N_10402,N_10783);
or U11596 (N_11596,N_10227,N_10838);
and U11597 (N_11597,N_10019,N_10863);
nand U11598 (N_11598,N_10816,N_10153);
or U11599 (N_11599,N_10373,N_10979);
nor U11600 (N_11600,N_10725,N_10391);
nand U11601 (N_11601,N_10557,N_10281);
or U11602 (N_11602,N_10399,N_10976);
nand U11603 (N_11603,N_10071,N_10760);
nor U11604 (N_11604,N_10109,N_10162);
xnor U11605 (N_11605,N_10609,N_10168);
or U11606 (N_11606,N_10641,N_10381);
or U11607 (N_11607,N_10321,N_10211);
or U11608 (N_11608,N_10586,N_10833);
xor U11609 (N_11609,N_10771,N_10192);
or U11610 (N_11610,N_10367,N_10856);
xor U11611 (N_11611,N_10899,N_10941);
or U11612 (N_11612,N_10169,N_10325);
or U11613 (N_11613,N_10025,N_10573);
nand U11614 (N_11614,N_10606,N_10167);
nand U11615 (N_11615,N_10124,N_10450);
nand U11616 (N_11616,N_10421,N_10336);
xor U11617 (N_11617,N_10942,N_10018);
or U11618 (N_11618,N_10423,N_10918);
and U11619 (N_11619,N_10264,N_10012);
nor U11620 (N_11620,N_10668,N_10482);
nor U11621 (N_11621,N_10479,N_10346);
or U11622 (N_11622,N_10230,N_10999);
nand U11623 (N_11623,N_10364,N_10733);
and U11624 (N_11624,N_10095,N_10661);
xor U11625 (N_11625,N_10858,N_10172);
or U11626 (N_11626,N_10954,N_10660);
nand U11627 (N_11627,N_10976,N_10317);
nor U11628 (N_11628,N_10101,N_10074);
nand U11629 (N_11629,N_10985,N_10995);
xor U11630 (N_11630,N_10945,N_10624);
nor U11631 (N_11631,N_10827,N_10048);
nor U11632 (N_11632,N_10306,N_10794);
and U11633 (N_11633,N_10544,N_10401);
xor U11634 (N_11634,N_10787,N_10719);
xnor U11635 (N_11635,N_10895,N_10890);
and U11636 (N_11636,N_10627,N_10098);
nand U11637 (N_11637,N_10235,N_10524);
nor U11638 (N_11638,N_10899,N_10856);
nand U11639 (N_11639,N_10328,N_10484);
nand U11640 (N_11640,N_10573,N_10203);
xnor U11641 (N_11641,N_10554,N_10663);
nor U11642 (N_11642,N_10053,N_10867);
xor U11643 (N_11643,N_10086,N_10386);
nor U11644 (N_11644,N_10639,N_10884);
xor U11645 (N_11645,N_10679,N_10149);
nor U11646 (N_11646,N_10031,N_10502);
nor U11647 (N_11647,N_10469,N_10559);
and U11648 (N_11648,N_10803,N_10990);
nand U11649 (N_11649,N_10259,N_10989);
nand U11650 (N_11650,N_10933,N_10884);
nor U11651 (N_11651,N_10482,N_10942);
xor U11652 (N_11652,N_10858,N_10313);
nand U11653 (N_11653,N_10448,N_10830);
nor U11654 (N_11654,N_10185,N_10360);
xnor U11655 (N_11655,N_10751,N_10510);
nand U11656 (N_11656,N_10634,N_10307);
nor U11657 (N_11657,N_10500,N_10537);
nor U11658 (N_11658,N_10953,N_10001);
nand U11659 (N_11659,N_10218,N_10283);
or U11660 (N_11660,N_10214,N_10275);
nor U11661 (N_11661,N_10094,N_10061);
nor U11662 (N_11662,N_10493,N_10863);
nor U11663 (N_11663,N_10731,N_10444);
or U11664 (N_11664,N_10790,N_10016);
xor U11665 (N_11665,N_10699,N_10300);
or U11666 (N_11666,N_10127,N_10876);
xnor U11667 (N_11667,N_10634,N_10212);
or U11668 (N_11668,N_10305,N_10306);
and U11669 (N_11669,N_10097,N_10431);
nand U11670 (N_11670,N_10787,N_10064);
xnor U11671 (N_11671,N_10896,N_10008);
nand U11672 (N_11672,N_10233,N_10470);
nand U11673 (N_11673,N_10946,N_10760);
or U11674 (N_11674,N_10149,N_10830);
or U11675 (N_11675,N_10305,N_10071);
and U11676 (N_11676,N_10516,N_10735);
and U11677 (N_11677,N_10823,N_10930);
nor U11678 (N_11678,N_10859,N_10178);
nor U11679 (N_11679,N_10763,N_10344);
and U11680 (N_11680,N_10862,N_10729);
or U11681 (N_11681,N_10859,N_10705);
and U11682 (N_11682,N_10538,N_10683);
nand U11683 (N_11683,N_10043,N_10731);
or U11684 (N_11684,N_10082,N_10996);
and U11685 (N_11685,N_10552,N_10360);
or U11686 (N_11686,N_10369,N_10125);
and U11687 (N_11687,N_10121,N_10868);
or U11688 (N_11688,N_10153,N_10876);
xor U11689 (N_11689,N_10048,N_10191);
and U11690 (N_11690,N_10110,N_10446);
and U11691 (N_11691,N_10396,N_10475);
xor U11692 (N_11692,N_10510,N_10819);
and U11693 (N_11693,N_10916,N_10372);
or U11694 (N_11694,N_10285,N_10495);
or U11695 (N_11695,N_10475,N_10641);
xnor U11696 (N_11696,N_10314,N_10568);
and U11697 (N_11697,N_10005,N_10656);
and U11698 (N_11698,N_10993,N_10589);
nor U11699 (N_11699,N_10656,N_10504);
or U11700 (N_11700,N_10231,N_10552);
and U11701 (N_11701,N_10064,N_10648);
or U11702 (N_11702,N_10424,N_10331);
xnor U11703 (N_11703,N_10831,N_10558);
nand U11704 (N_11704,N_10332,N_10486);
and U11705 (N_11705,N_10115,N_10672);
nand U11706 (N_11706,N_10978,N_10554);
and U11707 (N_11707,N_10019,N_10259);
or U11708 (N_11708,N_10743,N_10974);
nor U11709 (N_11709,N_10880,N_10241);
and U11710 (N_11710,N_10498,N_10877);
nand U11711 (N_11711,N_10228,N_10625);
and U11712 (N_11712,N_10520,N_10667);
nand U11713 (N_11713,N_10780,N_10528);
nor U11714 (N_11714,N_10360,N_10909);
or U11715 (N_11715,N_10278,N_10969);
and U11716 (N_11716,N_10595,N_10038);
nor U11717 (N_11717,N_10276,N_10121);
xor U11718 (N_11718,N_10897,N_10403);
nor U11719 (N_11719,N_10383,N_10707);
or U11720 (N_11720,N_10547,N_10471);
xor U11721 (N_11721,N_10655,N_10081);
nor U11722 (N_11722,N_10214,N_10358);
and U11723 (N_11723,N_10047,N_10504);
nor U11724 (N_11724,N_10127,N_10525);
or U11725 (N_11725,N_10411,N_10657);
xor U11726 (N_11726,N_10839,N_10444);
and U11727 (N_11727,N_10582,N_10704);
and U11728 (N_11728,N_10231,N_10461);
nand U11729 (N_11729,N_10819,N_10945);
and U11730 (N_11730,N_10118,N_10259);
nor U11731 (N_11731,N_10326,N_10546);
and U11732 (N_11732,N_10086,N_10801);
and U11733 (N_11733,N_10462,N_10996);
xor U11734 (N_11734,N_10533,N_10916);
nor U11735 (N_11735,N_10500,N_10695);
nand U11736 (N_11736,N_10241,N_10309);
or U11737 (N_11737,N_10296,N_10643);
xnor U11738 (N_11738,N_10793,N_10931);
nand U11739 (N_11739,N_10391,N_10865);
xor U11740 (N_11740,N_10884,N_10616);
nand U11741 (N_11741,N_10989,N_10938);
nand U11742 (N_11742,N_10349,N_10074);
and U11743 (N_11743,N_10889,N_10083);
and U11744 (N_11744,N_10888,N_10445);
and U11745 (N_11745,N_10838,N_10766);
nor U11746 (N_11746,N_10051,N_10946);
nand U11747 (N_11747,N_10112,N_10849);
and U11748 (N_11748,N_10832,N_10605);
and U11749 (N_11749,N_10443,N_10565);
nand U11750 (N_11750,N_10891,N_10787);
nand U11751 (N_11751,N_10957,N_10680);
nand U11752 (N_11752,N_10342,N_10281);
and U11753 (N_11753,N_10282,N_10927);
xor U11754 (N_11754,N_10421,N_10004);
xor U11755 (N_11755,N_10971,N_10197);
or U11756 (N_11756,N_10614,N_10376);
nor U11757 (N_11757,N_10978,N_10864);
and U11758 (N_11758,N_10144,N_10264);
nand U11759 (N_11759,N_10646,N_10399);
nor U11760 (N_11760,N_10686,N_10856);
nor U11761 (N_11761,N_10768,N_10530);
nor U11762 (N_11762,N_10558,N_10884);
nand U11763 (N_11763,N_10086,N_10575);
and U11764 (N_11764,N_10527,N_10248);
or U11765 (N_11765,N_10551,N_10733);
and U11766 (N_11766,N_10296,N_10563);
and U11767 (N_11767,N_10122,N_10819);
nor U11768 (N_11768,N_10833,N_10489);
or U11769 (N_11769,N_10571,N_10018);
nand U11770 (N_11770,N_10261,N_10611);
nand U11771 (N_11771,N_10170,N_10256);
and U11772 (N_11772,N_10124,N_10034);
nor U11773 (N_11773,N_10847,N_10309);
and U11774 (N_11774,N_10980,N_10794);
nand U11775 (N_11775,N_10510,N_10598);
or U11776 (N_11776,N_10556,N_10189);
nor U11777 (N_11777,N_10449,N_10833);
and U11778 (N_11778,N_10944,N_10798);
nand U11779 (N_11779,N_10040,N_10762);
xor U11780 (N_11780,N_10624,N_10845);
and U11781 (N_11781,N_10351,N_10912);
nor U11782 (N_11782,N_10541,N_10279);
or U11783 (N_11783,N_10673,N_10175);
and U11784 (N_11784,N_10856,N_10152);
xor U11785 (N_11785,N_10779,N_10049);
nand U11786 (N_11786,N_10195,N_10675);
nand U11787 (N_11787,N_10169,N_10971);
or U11788 (N_11788,N_10588,N_10138);
and U11789 (N_11789,N_10558,N_10013);
nand U11790 (N_11790,N_10263,N_10882);
nor U11791 (N_11791,N_10550,N_10659);
and U11792 (N_11792,N_10231,N_10544);
nor U11793 (N_11793,N_10602,N_10332);
nor U11794 (N_11794,N_10793,N_10365);
and U11795 (N_11795,N_10239,N_10318);
or U11796 (N_11796,N_10366,N_10948);
nand U11797 (N_11797,N_10393,N_10378);
nand U11798 (N_11798,N_10954,N_10793);
or U11799 (N_11799,N_10064,N_10894);
xor U11800 (N_11800,N_10441,N_10439);
or U11801 (N_11801,N_10257,N_10603);
or U11802 (N_11802,N_10664,N_10310);
nor U11803 (N_11803,N_10713,N_10135);
nor U11804 (N_11804,N_10689,N_10289);
and U11805 (N_11805,N_10343,N_10609);
nand U11806 (N_11806,N_10943,N_10328);
and U11807 (N_11807,N_10742,N_10588);
and U11808 (N_11808,N_10858,N_10444);
or U11809 (N_11809,N_10170,N_10446);
and U11810 (N_11810,N_10882,N_10405);
and U11811 (N_11811,N_10633,N_10331);
and U11812 (N_11812,N_10501,N_10479);
nand U11813 (N_11813,N_10866,N_10439);
or U11814 (N_11814,N_10047,N_10442);
xor U11815 (N_11815,N_10754,N_10929);
nor U11816 (N_11816,N_10879,N_10599);
nor U11817 (N_11817,N_10887,N_10244);
and U11818 (N_11818,N_10863,N_10974);
nor U11819 (N_11819,N_10907,N_10085);
nand U11820 (N_11820,N_10690,N_10121);
nand U11821 (N_11821,N_10167,N_10580);
or U11822 (N_11822,N_10253,N_10926);
xnor U11823 (N_11823,N_10184,N_10065);
or U11824 (N_11824,N_10642,N_10344);
nand U11825 (N_11825,N_10459,N_10405);
xor U11826 (N_11826,N_10501,N_10822);
xnor U11827 (N_11827,N_10005,N_10208);
nor U11828 (N_11828,N_10361,N_10970);
and U11829 (N_11829,N_10140,N_10899);
nand U11830 (N_11830,N_10089,N_10406);
xor U11831 (N_11831,N_10296,N_10857);
or U11832 (N_11832,N_10938,N_10216);
and U11833 (N_11833,N_10711,N_10218);
and U11834 (N_11834,N_10602,N_10732);
nor U11835 (N_11835,N_10232,N_10692);
or U11836 (N_11836,N_10353,N_10909);
and U11837 (N_11837,N_10853,N_10382);
and U11838 (N_11838,N_10064,N_10748);
and U11839 (N_11839,N_10279,N_10269);
nand U11840 (N_11840,N_10444,N_10283);
xor U11841 (N_11841,N_10707,N_10294);
xnor U11842 (N_11842,N_10053,N_10817);
or U11843 (N_11843,N_10178,N_10500);
nand U11844 (N_11844,N_10086,N_10441);
nand U11845 (N_11845,N_10527,N_10368);
and U11846 (N_11846,N_10820,N_10470);
nor U11847 (N_11847,N_10224,N_10739);
xor U11848 (N_11848,N_10377,N_10026);
nor U11849 (N_11849,N_10105,N_10671);
nor U11850 (N_11850,N_10064,N_10060);
nand U11851 (N_11851,N_10543,N_10383);
or U11852 (N_11852,N_10110,N_10274);
or U11853 (N_11853,N_10668,N_10644);
and U11854 (N_11854,N_10840,N_10591);
and U11855 (N_11855,N_10347,N_10719);
xnor U11856 (N_11856,N_10919,N_10558);
nand U11857 (N_11857,N_10682,N_10547);
and U11858 (N_11858,N_10697,N_10118);
nand U11859 (N_11859,N_10857,N_10485);
and U11860 (N_11860,N_10344,N_10237);
or U11861 (N_11861,N_10311,N_10262);
xor U11862 (N_11862,N_10998,N_10391);
or U11863 (N_11863,N_10939,N_10867);
or U11864 (N_11864,N_10862,N_10182);
nand U11865 (N_11865,N_10394,N_10524);
nor U11866 (N_11866,N_10923,N_10760);
nand U11867 (N_11867,N_10656,N_10391);
xor U11868 (N_11868,N_10172,N_10713);
xnor U11869 (N_11869,N_10143,N_10717);
or U11870 (N_11870,N_10711,N_10858);
nor U11871 (N_11871,N_10074,N_10889);
xor U11872 (N_11872,N_10468,N_10362);
xor U11873 (N_11873,N_10887,N_10563);
and U11874 (N_11874,N_10135,N_10565);
nand U11875 (N_11875,N_10144,N_10744);
nor U11876 (N_11876,N_10296,N_10720);
or U11877 (N_11877,N_10750,N_10460);
and U11878 (N_11878,N_10128,N_10556);
and U11879 (N_11879,N_10809,N_10067);
nand U11880 (N_11880,N_10850,N_10100);
nor U11881 (N_11881,N_10209,N_10543);
or U11882 (N_11882,N_10665,N_10765);
xor U11883 (N_11883,N_10369,N_10796);
and U11884 (N_11884,N_10693,N_10082);
or U11885 (N_11885,N_10709,N_10290);
or U11886 (N_11886,N_10204,N_10349);
nand U11887 (N_11887,N_10900,N_10270);
nand U11888 (N_11888,N_10872,N_10607);
xor U11889 (N_11889,N_10540,N_10665);
xor U11890 (N_11890,N_10741,N_10090);
nand U11891 (N_11891,N_10369,N_10329);
nand U11892 (N_11892,N_10520,N_10335);
nand U11893 (N_11893,N_10333,N_10991);
nand U11894 (N_11894,N_10617,N_10706);
xnor U11895 (N_11895,N_10724,N_10376);
nor U11896 (N_11896,N_10120,N_10207);
or U11897 (N_11897,N_10546,N_10404);
nor U11898 (N_11898,N_10473,N_10939);
and U11899 (N_11899,N_10565,N_10803);
xor U11900 (N_11900,N_10953,N_10624);
or U11901 (N_11901,N_10785,N_10620);
nand U11902 (N_11902,N_10028,N_10005);
xor U11903 (N_11903,N_10112,N_10560);
nand U11904 (N_11904,N_10144,N_10142);
nand U11905 (N_11905,N_10674,N_10418);
or U11906 (N_11906,N_10235,N_10588);
or U11907 (N_11907,N_10190,N_10784);
xor U11908 (N_11908,N_10601,N_10672);
nand U11909 (N_11909,N_10652,N_10791);
nand U11910 (N_11910,N_10628,N_10334);
nor U11911 (N_11911,N_10923,N_10231);
nor U11912 (N_11912,N_10899,N_10435);
and U11913 (N_11913,N_10798,N_10360);
xor U11914 (N_11914,N_10342,N_10536);
and U11915 (N_11915,N_10209,N_10384);
or U11916 (N_11916,N_10663,N_10721);
and U11917 (N_11917,N_10930,N_10524);
nor U11918 (N_11918,N_10638,N_10206);
xnor U11919 (N_11919,N_10609,N_10847);
nor U11920 (N_11920,N_10493,N_10018);
nor U11921 (N_11921,N_10865,N_10130);
nand U11922 (N_11922,N_10219,N_10506);
or U11923 (N_11923,N_10675,N_10288);
and U11924 (N_11924,N_10086,N_10456);
and U11925 (N_11925,N_10512,N_10683);
nand U11926 (N_11926,N_10086,N_10378);
nor U11927 (N_11927,N_10146,N_10789);
xnor U11928 (N_11928,N_10847,N_10046);
and U11929 (N_11929,N_10755,N_10332);
and U11930 (N_11930,N_10506,N_10385);
and U11931 (N_11931,N_10919,N_10733);
nand U11932 (N_11932,N_10838,N_10190);
xnor U11933 (N_11933,N_10261,N_10034);
nand U11934 (N_11934,N_10556,N_10546);
nand U11935 (N_11935,N_10276,N_10594);
nand U11936 (N_11936,N_10610,N_10287);
and U11937 (N_11937,N_10449,N_10270);
nand U11938 (N_11938,N_10064,N_10469);
xor U11939 (N_11939,N_10706,N_10657);
or U11940 (N_11940,N_10897,N_10057);
and U11941 (N_11941,N_10219,N_10844);
and U11942 (N_11942,N_10709,N_10226);
nand U11943 (N_11943,N_10754,N_10347);
or U11944 (N_11944,N_10776,N_10070);
or U11945 (N_11945,N_10326,N_10183);
nor U11946 (N_11946,N_10996,N_10586);
and U11947 (N_11947,N_10133,N_10627);
xnor U11948 (N_11948,N_10423,N_10244);
nor U11949 (N_11949,N_10280,N_10634);
nor U11950 (N_11950,N_10943,N_10594);
xor U11951 (N_11951,N_10169,N_10807);
nor U11952 (N_11952,N_10145,N_10254);
or U11953 (N_11953,N_10572,N_10813);
xor U11954 (N_11954,N_10947,N_10372);
nand U11955 (N_11955,N_10732,N_10457);
xnor U11956 (N_11956,N_10460,N_10444);
or U11957 (N_11957,N_10281,N_10148);
or U11958 (N_11958,N_10233,N_10047);
xor U11959 (N_11959,N_10348,N_10392);
and U11960 (N_11960,N_10065,N_10260);
nor U11961 (N_11961,N_10633,N_10045);
and U11962 (N_11962,N_10523,N_10435);
or U11963 (N_11963,N_10641,N_10419);
nand U11964 (N_11964,N_10625,N_10711);
or U11965 (N_11965,N_10869,N_10044);
or U11966 (N_11966,N_10049,N_10927);
or U11967 (N_11967,N_10401,N_10294);
xnor U11968 (N_11968,N_10511,N_10334);
and U11969 (N_11969,N_10757,N_10837);
or U11970 (N_11970,N_10181,N_10370);
nand U11971 (N_11971,N_10956,N_10829);
and U11972 (N_11972,N_10754,N_10657);
and U11973 (N_11973,N_10615,N_10042);
xor U11974 (N_11974,N_10371,N_10540);
xor U11975 (N_11975,N_10964,N_10451);
nand U11976 (N_11976,N_10872,N_10551);
and U11977 (N_11977,N_10857,N_10554);
xor U11978 (N_11978,N_10654,N_10532);
and U11979 (N_11979,N_10906,N_10263);
nand U11980 (N_11980,N_10270,N_10736);
or U11981 (N_11981,N_10286,N_10069);
nor U11982 (N_11982,N_10467,N_10301);
and U11983 (N_11983,N_10908,N_10391);
and U11984 (N_11984,N_10047,N_10494);
nor U11985 (N_11985,N_10849,N_10046);
or U11986 (N_11986,N_10398,N_10019);
and U11987 (N_11987,N_10825,N_10057);
nand U11988 (N_11988,N_10075,N_10849);
nand U11989 (N_11989,N_10456,N_10937);
or U11990 (N_11990,N_10801,N_10762);
nand U11991 (N_11991,N_10012,N_10817);
nand U11992 (N_11992,N_10094,N_10132);
nand U11993 (N_11993,N_10826,N_10232);
nand U11994 (N_11994,N_10106,N_10707);
nand U11995 (N_11995,N_10413,N_10362);
xor U11996 (N_11996,N_10324,N_10087);
and U11997 (N_11997,N_10343,N_10380);
xor U11998 (N_11998,N_10553,N_10249);
nand U11999 (N_11999,N_10103,N_10869);
or U12000 (N_12000,N_11363,N_11718);
and U12001 (N_12001,N_11944,N_11369);
nor U12002 (N_12002,N_11243,N_11744);
nor U12003 (N_12003,N_11602,N_11372);
and U12004 (N_12004,N_11194,N_11448);
nor U12005 (N_12005,N_11925,N_11181);
or U12006 (N_12006,N_11604,N_11464);
and U12007 (N_12007,N_11964,N_11748);
or U12008 (N_12008,N_11077,N_11493);
nor U12009 (N_12009,N_11467,N_11587);
nor U12010 (N_12010,N_11578,N_11528);
xnor U12011 (N_12011,N_11025,N_11230);
and U12012 (N_12012,N_11118,N_11348);
or U12013 (N_12013,N_11111,N_11033);
nor U12014 (N_12014,N_11569,N_11091);
nand U12015 (N_12015,N_11553,N_11839);
and U12016 (N_12016,N_11040,N_11392);
or U12017 (N_12017,N_11263,N_11438);
and U12018 (N_12018,N_11217,N_11252);
and U12019 (N_12019,N_11843,N_11772);
nor U12020 (N_12020,N_11982,N_11024);
nor U12021 (N_12021,N_11271,N_11761);
xnor U12022 (N_12022,N_11513,N_11399);
or U12023 (N_12023,N_11196,N_11690);
and U12024 (N_12024,N_11164,N_11981);
nor U12025 (N_12025,N_11110,N_11965);
nor U12026 (N_12026,N_11841,N_11276);
xor U12027 (N_12027,N_11031,N_11305);
and U12028 (N_12028,N_11650,N_11092);
or U12029 (N_12029,N_11142,N_11222);
nand U12030 (N_12030,N_11300,N_11155);
or U12031 (N_12031,N_11818,N_11732);
and U12032 (N_12032,N_11525,N_11901);
and U12033 (N_12033,N_11488,N_11970);
and U12034 (N_12034,N_11803,N_11016);
and U12035 (N_12035,N_11617,N_11371);
nor U12036 (N_12036,N_11038,N_11910);
nand U12037 (N_12037,N_11461,N_11408);
or U12038 (N_12038,N_11572,N_11504);
xor U12039 (N_12039,N_11104,N_11869);
nand U12040 (N_12040,N_11746,N_11559);
or U12041 (N_12041,N_11888,N_11254);
and U12042 (N_12042,N_11045,N_11470);
or U12043 (N_12043,N_11855,N_11814);
nand U12044 (N_12044,N_11103,N_11229);
nor U12045 (N_12045,N_11793,N_11264);
nor U12046 (N_12046,N_11825,N_11460);
nor U12047 (N_12047,N_11941,N_11066);
or U12048 (N_12048,N_11342,N_11220);
nand U12049 (N_12049,N_11757,N_11483);
nand U12050 (N_12050,N_11861,N_11562);
nand U12051 (N_12051,N_11863,N_11554);
xor U12052 (N_12052,N_11389,N_11688);
and U12053 (N_12053,N_11773,N_11445);
xnor U12054 (N_12054,N_11902,N_11245);
nand U12055 (N_12055,N_11734,N_11093);
and U12056 (N_12056,N_11157,N_11939);
and U12057 (N_12057,N_11132,N_11019);
xnor U12058 (N_12058,N_11766,N_11433);
xnor U12059 (N_12059,N_11440,N_11236);
and U12060 (N_12060,N_11691,N_11089);
nor U12061 (N_12061,N_11210,N_11121);
nand U12062 (N_12062,N_11439,N_11899);
nand U12063 (N_12063,N_11619,N_11410);
nand U12064 (N_12064,N_11361,N_11611);
or U12065 (N_12065,N_11677,N_11852);
nand U12066 (N_12066,N_11849,N_11332);
and U12067 (N_12067,N_11740,N_11655);
nand U12068 (N_12068,N_11983,N_11726);
or U12069 (N_12069,N_11540,N_11208);
or U12070 (N_12070,N_11323,N_11224);
nand U12071 (N_12071,N_11897,N_11756);
xor U12072 (N_12072,N_11890,N_11596);
xor U12073 (N_12073,N_11645,N_11681);
nor U12074 (N_12074,N_11898,N_11268);
and U12075 (N_12075,N_11937,N_11857);
nor U12076 (N_12076,N_11518,N_11895);
xnor U12077 (N_12077,N_11636,N_11162);
nand U12078 (N_12078,N_11146,N_11749);
or U12079 (N_12079,N_11286,N_11736);
or U12080 (N_12080,N_11283,N_11973);
or U12081 (N_12081,N_11752,N_11651);
nand U12082 (N_12082,N_11737,N_11123);
and U12083 (N_12083,N_11282,N_11912);
and U12084 (N_12084,N_11495,N_11931);
nand U12085 (N_12085,N_11711,N_11062);
xor U12086 (N_12086,N_11624,N_11694);
nor U12087 (N_12087,N_11152,N_11786);
or U12088 (N_12088,N_11696,N_11850);
nand U12089 (N_12089,N_11076,N_11835);
or U12090 (N_12090,N_11991,N_11679);
or U12091 (N_12091,N_11247,N_11889);
xnor U12092 (N_12092,N_11451,N_11797);
xnor U12093 (N_12093,N_11138,N_11635);
nor U12094 (N_12094,N_11792,N_11992);
or U12095 (N_12095,N_11277,N_11427);
nand U12096 (N_12096,N_11980,N_11350);
nor U12097 (N_12097,N_11447,N_11833);
and U12098 (N_12098,N_11259,N_11086);
xnor U12099 (N_12099,N_11358,N_11179);
and U12100 (N_12100,N_11919,N_11543);
xnor U12101 (N_12101,N_11585,N_11794);
or U12102 (N_12102,N_11057,N_11760);
nand U12103 (N_12103,N_11722,N_11891);
xor U12104 (N_12104,N_11446,N_11697);
nand U12105 (N_12105,N_11203,N_11771);
nand U12106 (N_12106,N_11892,N_11715);
and U12107 (N_12107,N_11612,N_11933);
nand U12108 (N_12108,N_11468,N_11339);
or U12109 (N_12109,N_11729,N_11163);
or U12110 (N_12110,N_11848,N_11584);
or U12111 (N_12111,N_11812,N_11436);
nor U12112 (N_12112,N_11261,N_11506);
nor U12113 (N_12113,N_11357,N_11634);
or U12114 (N_12114,N_11564,N_11683);
and U12115 (N_12115,N_11047,N_11692);
nor U12116 (N_12116,N_11943,N_11637);
or U12117 (N_12117,N_11918,N_11876);
or U12118 (N_12118,N_11213,N_11327);
and U12119 (N_12119,N_11158,N_11237);
and U12120 (N_12120,N_11599,N_11826);
nor U12121 (N_12121,N_11595,N_11494);
nor U12122 (N_12122,N_11514,N_11275);
or U12123 (N_12123,N_11087,N_11065);
and U12124 (N_12124,N_11806,N_11633);
or U12125 (N_12125,N_11838,N_11127);
nor U12126 (N_12126,N_11886,N_11364);
nor U12127 (N_12127,N_11844,N_11106);
xor U12128 (N_12128,N_11720,N_11731);
or U12129 (N_12129,N_11824,N_11529);
or U12130 (N_12130,N_11547,N_11882);
nand U12131 (N_12131,N_11625,N_11568);
nor U12132 (N_12132,N_11708,N_11523);
and U12133 (N_12133,N_11510,N_11974);
xor U12134 (N_12134,N_11490,N_11192);
and U12135 (N_12135,N_11821,N_11597);
nand U12136 (N_12136,N_11977,N_11039);
and U12137 (N_12137,N_11796,N_11022);
nand U12138 (N_12138,N_11951,N_11102);
xnor U12139 (N_12139,N_11374,N_11541);
xor U12140 (N_12140,N_11462,N_11030);
nor U12141 (N_12141,N_11647,N_11990);
xor U12142 (N_12142,N_11575,N_11840);
nand U12143 (N_12143,N_11054,N_11714);
and U12144 (N_12144,N_11505,N_11516);
and U12145 (N_12145,N_11425,N_11444);
nor U12146 (N_12146,N_11519,N_11166);
nand U12147 (N_12147,N_11485,N_11005);
xnor U12148 (N_12148,N_11487,N_11116);
and U12149 (N_12149,N_11649,N_11082);
or U12150 (N_12150,N_11207,N_11453);
or U12151 (N_12151,N_11417,N_11463);
xnor U12152 (N_12152,N_11884,N_11627);
xor U12153 (N_12153,N_11682,N_11819);
xnor U12154 (N_12154,N_11570,N_11067);
and U12155 (N_12155,N_11362,N_11209);
nand U12156 (N_12156,N_11542,N_11950);
nand U12157 (N_12157,N_11548,N_11112);
xor U12158 (N_12158,N_11319,N_11287);
and U12159 (N_12159,N_11430,N_11903);
or U12160 (N_12160,N_11469,N_11338);
and U12161 (N_12161,N_11044,N_11450);
nand U12162 (N_12162,N_11945,N_11013);
nor U12163 (N_12163,N_11134,N_11255);
nand U12164 (N_12164,N_11957,N_11791);
and U12165 (N_12165,N_11193,N_11537);
and U12166 (N_12166,N_11457,N_11337);
and U12167 (N_12167,N_11307,N_11795);
xnor U12168 (N_12168,N_11001,N_11706);
or U12169 (N_12169,N_11741,N_11807);
nor U12170 (N_12170,N_11285,N_11909);
nand U12171 (N_12171,N_11588,N_11280);
xnor U12172 (N_12172,N_11947,N_11404);
nand U12173 (N_12173,N_11508,N_11401);
and U12174 (N_12174,N_11815,N_11403);
xnor U12175 (N_12175,N_11967,N_11769);
nor U12176 (N_12176,N_11799,N_11422);
and U12177 (N_12177,N_11418,N_11698);
xnor U12178 (N_12178,N_11297,N_11143);
xor U12179 (N_12179,N_11336,N_11183);
and U12180 (N_12180,N_11662,N_11386);
nand U12181 (N_12181,N_11221,N_11334);
nor U12182 (N_12182,N_11871,N_11566);
xnor U12183 (N_12183,N_11060,N_11703);
or U12184 (N_12184,N_11994,N_11189);
or U12185 (N_12185,N_11070,N_11191);
or U12186 (N_12186,N_11292,N_11184);
nor U12187 (N_12187,N_11136,N_11658);
and U12188 (N_12188,N_11712,N_11501);
and U12189 (N_12189,N_11244,N_11032);
nand U12190 (N_12190,N_11673,N_11622);
or U12191 (N_12191,N_11932,N_11411);
and U12192 (N_12192,N_11789,N_11449);
xor U12193 (N_12193,N_11721,N_11675);
and U12194 (N_12194,N_11028,N_11180);
and U12195 (N_12195,N_11281,N_11552);
or U12196 (N_12196,N_11754,N_11412);
or U12197 (N_12197,N_11787,N_11249);
xnor U12198 (N_12198,N_11859,N_11988);
nand U12199 (N_12199,N_11303,N_11666);
or U12200 (N_12200,N_11148,N_11441);
or U12201 (N_12201,N_11428,N_11081);
xnor U12202 (N_12202,N_11742,N_11896);
and U12203 (N_12203,N_11115,N_11571);
xnor U12204 (N_12204,N_11836,N_11242);
and U12205 (N_12205,N_11996,N_11214);
nand U12206 (N_12206,N_11317,N_11156);
and U12207 (N_12207,N_11478,N_11080);
and U12208 (N_12208,N_11266,N_11785);
nor U12209 (N_12209,N_11665,N_11423);
nor U12210 (N_12210,N_11075,N_11656);
nand U12211 (N_12211,N_11379,N_11809);
or U12212 (N_12212,N_11751,N_11653);
nand U12213 (N_12213,N_11608,N_11420);
and U12214 (N_12214,N_11432,N_11544);
nor U12215 (N_12215,N_11875,N_11798);
and U12216 (N_12216,N_11832,N_11680);
nand U12217 (N_12217,N_11830,N_11927);
or U12218 (N_12218,N_11375,N_11880);
nand U12219 (N_12219,N_11185,N_11195);
or U12220 (N_12220,N_11705,N_11328);
nand U12221 (N_12221,N_11670,N_11003);
xor U12222 (N_12222,N_11605,N_11701);
nor U12223 (N_12223,N_11130,N_11421);
or U12224 (N_12224,N_11002,N_11971);
nand U12225 (N_12225,N_11061,N_11709);
xnor U12226 (N_12226,N_11739,N_11397);
xnor U12227 (N_12227,N_11802,N_11015);
nand U12228 (N_12228,N_11878,N_11784);
or U12229 (N_12229,N_11862,N_11538);
and U12230 (N_12230,N_11790,N_11966);
nand U12231 (N_12231,N_11476,N_11567);
nor U12232 (N_12232,N_11924,N_11856);
and U12233 (N_12233,N_11465,N_11241);
nor U12234 (N_12234,N_11099,N_11190);
or U12235 (N_12235,N_11043,N_11172);
or U12236 (N_12236,N_11131,N_11642);
or U12237 (N_12237,N_11452,N_11068);
nor U12238 (N_12238,N_11010,N_11592);
and U12239 (N_12239,N_11046,N_11955);
nor U12240 (N_12240,N_11177,N_11288);
nor U12241 (N_12241,N_11206,N_11913);
and U12242 (N_12242,N_11048,N_11289);
xor U12243 (N_12243,N_11735,N_11550);
nor U12244 (N_12244,N_11351,N_11188);
or U12245 (N_12245,N_11512,N_11484);
and U12246 (N_12246,N_11186,N_11227);
or U12247 (N_12247,N_11382,N_11151);
nand U12248 (N_12248,N_11233,N_11916);
or U12249 (N_12249,N_11942,N_11956);
or U12250 (N_12250,N_11041,N_11128);
and U12251 (N_12251,N_11866,N_11346);
nor U12252 (N_12252,N_11962,N_11728);
and U12253 (N_12253,N_11969,N_11434);
or U12254 (N_12254,N_11834,N_11667);
and U12255 (N_12255,N_11109,N_11272);
xor U12256 (N_12256,N_11187,N_11384);
nor U12257 (N_12257,N_11580,N_11455);
xor U12258 (N_12258,N_11816,N_11893);
nand U12259 (N_12259,N_11657,N_11074);
nor U12260 (N_12260,N_11777,N_11579);
xor U12261 (N_12261,N_11788,N_11979);
or U12262 (N_12262,N_11313,N_11489);
nand U12263 (N_12263,N_11299,N_11879);
nand U12264 (N_12264,N_11270,N_11576);
nor U12265 (N_12265,N_11049,N_11398);
or U12266 (N_12266,N_11098,N_11854);
xnor U12267 (N_12267,N_11034,N_11551);
xor U12268 (N_12268,N_11354,N_11725);
or U12269 (N_12269,N_11402,N_11008);
or U12270 (N_12270,N_11717,N_11563);
or U12271 (N_12271,N_11377,N_11928);
nand U12272 (N_12272,N_11699,N_11783);
nor U12273 (N_12273,N_11908,N_11150);
xor U12274 (N_12274,N_11904,N_11822);
xnor U12275 (N_12275,N_11072,N_11558);
and U12276 (N_12276,N_11056,N_11700);
and U12277 (N_12277,N_11561,N_11312);
and U12278 (N_12278,N_11119,N_11765);
and U12279 (N_12279,N_11205,N_11395);
nand U12280 (N_12280,N_11331,N_11120);
nand U12281 (N_12281,N_11154,N_11808);
nor U12282 (N_12282,N_11366,N_11987);
nor U12283 (N_12283,N_11733,N_11324);
xor U12284 (N_12284,N_11409,N_11231);
nand U12285 (N_12285,N_11767,N_11607);
or U12286 (N_12286,N_11406,N_11674);
nand U12287 (N_12287,N_11020,N_11574);
and U12288 (N_12288,N_11845,N_11429);
xor U12289 (N_12289,N_11995,N_11606);
nand U12290 (N_12290,N_11173,N_11321);
nand U12291 (N_12291,N_11594,N_11929);
nor U12292 (N_12292,N_11546,N_11911);
xnor U12293 (N_12293,N_11813,N_11456);
and U12294 (N_12294,N_11480,N_11027);
or U12295 (N_12295,N_11641,N_11290);
xnor U12296 (N_12296,N_11129,N_11923);
nor U12297 (N_12297,N_11710,N_11745);
or U12298 (N_12298,N_11341,N_11472);
or U12299 (N_12299,N_11664,N_11435);
and U12300 (N_12300,N_11105,N_11774);
nor U12301 (N_12301,N_11628,N_11431);
or U12302 (N_12302,N_11326,N_11630);
nor U12303 (N_12303,N_11723,N_11847);
xor U12304 (N_12304,N_11122,N_11517);
or U12305 (N_12305,N_11764,N_11085);
nand U12306 (N_12306,N_11829,N_11269);
or U12307 (N_12307,N_11952,N_11058);
xnor U12308 (N_12308,N_11414,N_11521);
and U12309 (N_12309,N_11646,N_11695);
xor U12310 (N_12310,N_11780,N_11114);
nand U12311 (N_12311,N_11643,N_11533);
nand U12312 (N_12312,N_11426,N_11250);
nor U12313 (N_12313,N_11278,N_11021);
nand U12314 (N_12314,N_11330,N_11376);
or U12315 (N_12315,N_11496,N_11870);
xnor U12316 (N_12316,N_11026,N_11831);
nor U12317 (N_12317,N_11094,N_11652);
nand U12318 (N_12318,N_11492,N_11084);
and U12319 (N_12319,N_11820,N_11877);
or U12320 (N_12320,N_11997,N_11858);
nand U12321 (N_12321,N_11800,N_11125);
nand U12322 (N_12322,N_11212,N_11581);
xor U12323 (N_12323,N_11894,N_11640);
or U12324 (N_12324,N_11873,N_11394);
nor U12325 (N_12325,N_11126,N_11088);
and U12326 (N_12326,N_11353,N_11023);
and U12327 (N_12327,N_11144,N_11459);
or U12328 (N_12328,N_11175,N_11917);
or U12329 (N_12329,N_11586,N_11295);
nor U12330 (N_12330,N_11135,N_11293);
nor U12331 (N_12331,N_11770,N_11405);
nand U12332 (N_12332,N_11169,N_11671);
or U12333 (N_12333,N_11614,N_11344);
nand U12334 (N_12334,N_11416,N_11265);
xor U12335 (N_12335,N_11133,N_11491);
or U12336 (N_12336,N_11101,N_11390);
and U12337 (N_12337,N_11811,N_11267);
nand U12338 (N_12338,N_11583,N_11368);
xor U12339 (N_12339,N_11284,N_11343);
or U12340 (N_12340,N_11827,N_11975);
nor U12341 (N_12341,N_11753,N_11437);
or U12342 (N_12342,N_11724,N_11096);
nand U12343 (N_12343,N_11147,N_11885);
xor U12344 (N_12344,N_11978,N_11298);
and U12345 (N_12345,N_11644,N_11631);
nand U12346 (N_12346,N_11618,N_11176);
nand U12347 (N_12347,N_11872,N_11986);
or U12348 (N_12348,N_11659,N_11515);
and U12349 (N_12349,N_11958,N_11663);
nor U12350 (N_12350,N_11383,N_11549);
nand U12351 (N_12351,N_11590,N_11388);
or U12352 (N_12352,N_11380,N_11454);
nor U12353 (N_12353,N_11949,N_11874);
and U12354 (N_12354,N_11522,N_11145);
or U12355 (N_12355,N_11704,N_11443);
nor U12356 (N_12356,N_11935,N_11329);
xor U12357 (N_12357,N_11968,N_11356);
nand U12358 (N_12358,N_11253,N_11593);
nor U12359 (N_12359,N_11322,N_11851);
nand U12360 (N_12360,N_11926,N_11998);
or U12361 (N_12361,N_11349,N_11707);
or U12362 (N_12362,N_11486,N_11174);
nand U12363 (N_12363,N_11499,N_11415);
or U12364 (N_12364,N_11778,N_11000);
and U12365 (N_12365,N_11017,N_11301);
or U12366 (N_12366,N_11310,N_11340);
nand U12367 (N_12367,N_11258,N_11325);
or U12368 (N_12368,N_11846,N_11900);
or U12369 (N_12369,N_11532,N_11226);
and U12370 (N_12370,N_11475,N_11768);
nand U12371 (N_12371,N_11279,N_11314);
xor U12372 (N_12372,N_11407,N_11167);
or U12373 (N_12373,N_11396,N_11984);
xnor U12374 (N_12374,N_11672,N_11613);
and U12375 (N_12375,N_11867,N_11837);
nand U12376 (N_12376,N_11097,N_11661);
nand U12377 (N_12377,N_11479,N_11573);
xnor U12378 (N_12378,N_11993,N_11530);
nand U12379 (N_12379,N_11201,N_11477);
nand U12380 (N_12380,N_11365,N_11234);
xnor U12381 (N_12381,N_11320,N_11758);
nand U12382 (N_12382,N_11042,N_11137);
or U12383 (N_12383,N_11083,N_11507);
xor U12384 (N_12384,N_11498,N_11999);
or U12385 (N_12385,N_11064,N_11959);
xnor U12386 (N_12386,N_11881,N_11055);
nand U12387 (N_12387,N_11198,N_11079);
and U12388 (N_12388,N_11256,N_11117);
nand U12389 (N_12389,N_11161,N_11200);
or U12390 (N_12390,N_11260,N_11577);
nor U12391 (N_12391,N_11621,N_11306);
nor U12392 (N_12392,N_11311,N_11355);
or U12393 (N_12393,N_11702,N_11828);
or U12394 (N_12394,N_11948,N_11051);
xnor U12395 (N_12395,N_11853,N_11620);
nor U12396 (N_12396,N_11626,N_11527);
xor U12397 (N_12397,N_11381,N_11302);
and U12398 (N_12398,N_11639,N_11373);
xnor U12399 (N_12399,N_11385,N_11865);
and U12400 (N_12400,N_11262,N_11050);
nor U12401 (N_12401,N_11014,N_11615);
xnor U12402 (N_12402,N_11616,N_11333);
nand U12403 (N_12403,N_11170,N_11335);
xnor U12404 (N_12404,N_11603,N_11171);
nor U12405 (N_12405,N_11378,N_11178);
nor U12406 (N_12406,N_11304,N_11442);
and U12407 (N_12407,N_11199,N_11922);
and U12408 (N_12408,N_11387,N_11141);
nor U12409 (N_12409,N_11946,N_11750);
nand U12410 (N_12410,N_11458,N_11011);
or U12411 (N_12411,N_11810,N_11248);
nor U12412 (N_12412,N_11907,N_11842);
nand U12413 (N_12413,N_11960,N_11560);
xor U12414 (N_12414,N_11108,N_11914);
nor U12415 (N_12415,N_11763,N_11318);
or U12416 (N_12416,N_11029,N_11609);
nand U12417 (N_12417,N_11693,N_11887);
nor U12418 (N_12418,N_11052,N_11526);
nand U12419 (N_12419,N_11685,N_11823);
nor U12420 (N_12420,N_11905,N_11360);
nand U12421 (N_12421,N_11938,N_11782);
nor U12422 (N_12422,N_11009,N_11296);
and U12423 (N_12423,N_11601,N_11555);
xor U12424 (N_12424,N_11954,N_11713);
and U12425 (N_12425,N_11976,N_11308);
nor U12426 (N_12426,N_11535,N_11759);
xnor U12427 (N_12427,N_11294,N_11113);
xnor U12428 (N_12428,N_11915,N_11095);
or U12429 (N_12429,N_11497,N_11520);
xor U12430 (N_12430,N_11149,N_11124);
xor U12431 (N_12431,N_11805,N_11315);
nand U12432 (N_12432,N_11921,N_11972);
and U12433 (N_12433,N_11291,N_11139);
xnor U12434 (N_12434,N_11738,N_11069);
and U12435 (N_12435,N_11687,N_11218);
nor U12436 (N_12436,N_11063,N_11598);
and U12437 (N_12437,N_11035,N_11012);
and U12438 (N_12438,N_11182,N_11159);
nor U12439 (N_12439,N_11400,N_11235);
or U12440 (N_12440,N_11153,N_11686);
nand U12441 (N_12441,N_11589,N_11503);
xnor U12442 (N_12442,N_11053,N_11669);
and U12443 (N_12443,N_11565,N_11036);
xnor U12444 (N_12444,N_11660,N_11775);
or U12445 (N_12445,N_11007,N_11239);
xor U12446 (N_12446,N_11274,N_11864);
xnor U12447 (N_12447,N_11018,N_11367);
xor U12448 (N_12448,N_11719,N_11545);
xnor U12449 (N_12449,N_11934,N_11524);
xor U12450 (N_12450,N_11240,N_11689);
or U12451 (N_12451,N_11059,N_11920);
nor U12452 (N_12452,N_11779,N_11107);
or U12453 (N_12453,N_11370,N_11246);
xor U12454 (N_12454,N_11225,N_11073);
nor U12455 (N_12455,N_11502,N_11776);
nor U12456 (N_12456,N_11953,N_11100);
or U12457 (N_12457,N_11743,N_11638);
nor U12458 (N_12458,N_11654,N_11202);
xnor U12459 (N_12459,N_11359,N_11391);
nor U12460 (N_12460,N_11762,N_11716);
or U12461 (N_12461,N_11471,N_11801);
and U12462 (N_12462,N_11215,N_11090);
and U12463 (N_12463,N_11668,N_11232);
and U12464 (N_12464,N_11610,N_11004);
or U12465 (N_12465,N_11509,N_11273);
and U12466 (N_12466,N_11860,N_11557);
nand U12467 (N_12467,N_11868,N_11781);
or U12468 (N_12468,N_11419,N_11309);
nor U12469 (N_12469,N_11071,N_11219);
nor U12470 (N_12470,N_11536,N_11989);
xor U12471 (N_12471,N_11676,N_11204);
nand U12472 (N_12472,N_11473,N_11684);
and U12473 (N_12473,N_11481,N_11936);
nor U12474 (N_12474,N_11474,N_11591);
xnor U12475 (N_12475,N_11500,N_11539);
or U12476 (N_12476,N_11165,N_11632);
and U12477 (N_12477,N_11006,N_11582);
and U12478 (N_12478,N_11393,N_11648);
nor U12479 (N_12479,N_11963,N_11347);
nand U12480 (N_12480,N_11730,N_11037);
or U12481 (N_12481,N_11316,N_11160);
nor U12482 (N_12482,N_11251,N_11078);
nand U12483 (N_12483,N_11985,N_11747);
xnor U12484 (N_12484,N_11140,N_11556);
xnor U12485 (N_12485,N_11623,N_11238);
nand U12486 (N_12486,N_11817,N_11961);
nor U12487 (N_12487,N_11466,N_11940);
nor U12488 (N_12488,N_11511,N_11883);
nand U12489 (N_12489,N_11930,N_11534);
xnor U12490 (N_12490,N_11216,N_11211);
xor U12491 (N_12491,N_11531,N_11482);
nor U12492 (N_12492,N_11600,N_11413);
nand U12493 (N_12493,N_11223,N_11804);
and U12494 (N_12494,N_11755,N_11228);
or U12495 (N_12495,N_11424,N_11352);
nor U12496 (N_12496,N_11345,N_11906);
and U12497 (N_12497,N_11678,N_11197);
nand U12498 (N_12498,N_11257,N_11168);
or U12499 (N_12499,N_11629,N_11727);
xnor U12500 (N_12500,N_11922,N_11658);
nand U12501 (N_12501,N_11946,N_11766);
nor U12502 (N_12502,N_11993,N_11884);
nor U12503 (N_12503,N_11999,N_11977);
and U12504 (N_12504,N_11815,N_11741);
nand U12505 (N_12505,N_11144,N_11484);
nand U12506 (N_12506,N_11083,N_11451);
xnor U12507 (N_12507,N_11970,N_11391);
xor U12508 (N_12508,N_11332,N_11736);
nor U12509 (N_12509,N_11237,N_11950);
and U12510 (N_12510,N_11397,N_11869);
and U12511 (N_12511,N_11991,N_11370);
or U12512 (N_12512,N_11859,N_11990);
nand U12513 (N_12513,N_11560,N_11605);
or U12514 (N_12514,N_11282,N_11449);
nand U12515 (N_12515,N_11839,N_11722);
nor U12516 (N_12516,N_11530,N_11514);
and U12517 (N_12517,N_11072,N_11682);
nor U12518 (N_12518,N_11256,N_11920);
nor U12519 (N_12519,N_11318,N_11256);
nand U12520 (N_12520,N_11466,N_11858);
and U12521 (N_12521,N_11933,N_11359);
or U12522 (N_12522,N_11871,N_11129);
xor U12523 (N_12523,N_11380,N_11780);
nor U12524 (N_12524,N_11386,N_11413);
xnor U12525 (N_12525,N_11454,N_11690);
or U12526 (N_12526,N_11749,N_11200);
nor U12527 (N_12527,N_11404,N_11242);
and U12528 (N_12528,N_11483,N_11695);
nand U12529 (N_12529,N_11721,N_11289);
xor U12530 (N_12530,N_11845,N_11156);
nand U12531 (N_12531,N_11499,N_11649);
nor U12532 (N_12532,N_11685,N_11821);
or U12533 (N_12533,N_11705,N_11751);
or U12534 (N_12534,N_11344,N_11556);
nor U12535 (N_12535,N_11226,N_11941);
nor U12536 (N_12536,N_11938,N_11431);
and U12537 (N_12537,N_11936,N_11965);
nand U12538 (N_12538,N_11751,N_11825);
xor U12539 (N_12539,N_11802,N_11906);
nand U12540 (N_12540,N_11603,N_11473);
xor U12541 (N_12541,N_11831,N_11549);
nor U12542 (N_12542,N_11997,N_11795);
or U12543 (N_12543,N_11710,N_11078);
xor U12544 (N_12544,N_11345,N_11788);
xnor U12545 (N_12545,N_11140,N_11801);
xnor U12546 (N_12546,N_11253,N_11999);
xnor U12547 (N_12547,N_11472,N_11487);
and U12548 (N_12548,N_11839,N_11283);
nor U12549 (N_12549,N_11062,N_11761);
nand U12550 (N_12550,N_11572,N_11262);
xnor U12551 (N_12551,N_11351,N_11293);
or U12552 (N_12552,N_11550,N_11148);
and U12553 (N_12553,N_11049,N_11099);
or U12554 (N_12554,N_11787,N_11378);
or U12555 (N_12555,N_11933,N_11925);
or U12556 (N_12556,N_11048,N_11336);
nand U12557 (N_12557,N_11939,N_11980);
xor U12558 (N_12558,N_11625,N_11573);
or U12559 (N_12559,N_11753,N_11176);
and U12560 (N_12560,N_11224,N_11796);
nand U12561 (N_12561,N_11461,N_11591);
nor U12562 (N_12562,N_11340,N_11476);
xnor U12563 (N_12563,N_11398,N_11616);
nor U12564 (N_12564,N_11528,N_11647);
nand U12565 (N_12565,N_11782,N_11709);
or U12566 (N_12566,N_11004,N_11388);
and U12567 (N_12567,N_11460,N_11562);
nand U12568 (N_12568,N_11327,N_11871);
nor U12569 (N_12569,N_11514,N_11697);
or U12570 (N_12570,N_11443,N_11385);
or U12571 (N_12571,N_11822,N_11019);
and U12572 (N_12572,N_11059,N_11802);
xnor U12573 (N_12573,N_11321,N_11648);
or U12574 (N_12574,N_11108,N_11208);
xnor U12575 (N_12575,N_11286,N_11285);
nor U12576 (N_12576,N_11273,N_11002);
nor U12577 (N_12577,N_11472,N_11456);
and U12578 (N_12578,N_11031,N_11638);
nand U12579 (N_12579,N_11124,N_11946);
and U12580 (N_12580,N_11082,N_11087);
xnor U12581 (N_12581,N_11597,N_11160);
nand U12582 (N_12582,N_11225,N_11984);
nor U12583 (N_12583,N_11458,N_11177);
and U12584 (N_12584,N_11068,N_11430);
nand U12585 (N_12585,N_11476,N_11806);
and U12586 (N_12586,N_11018,N_11142);
or U12587 (N_12587,N_11082,N_11287);
nor U12588 (N_12588,N_11891,N_11565);
nor U12589 (N_12589,N_11961,N_11354);
and U12590 (N_12590,N_11000,N_11937);
or U12591 (N_12591,N_11630,N_11168);
and U12592 (N_12592,N_11182,N_11469);
or U12593 (N_12593,N_11848,N_11686);
nand U12594 (N_12594,N_11076,N_11356);
nand U12595 (N_12595,N_11890,N_11747);
and U12596 (N_12596,N_11061,N_11581);
or U12597 (N_12597,N_11929,N_11487);
nand U12598 (N_12598,N_11432,N_11915);
or U12599 (N_12599,N_11953,N_11845);
xnor U12600 (N_12600,N_11483,N_11069);
xnor U12601 (N_12601,N_11915,N_11006);
nand U12602 (N_12602,N_11271,N_11964);
or U12603 (N_12603,N_11786,N_11927);
nor U12604 (N_12604,N_11985,N_11024);
or U12605 (N_12605,N_11632,N_11447);
nor U12606 (N_12606,N_11862,N_11260);
xor U12607 (N_12607,N_11544,N_11547);
xnor U12608 (N_12608,N_11797,N_11341);
xor U12609 (N_12609,N_11254,N_11297);
nand U12610 (N_12610,N_11969,N_11773);
nand U12611 (N_12611,N_11124,N_11856);
and U12612 (N_12612,N_11712,N_11927);
xnor U12613 (N_12613,N_11069,N_11114);
xnor U12614 (N_12614,N_11250,N_11683);
nand U12615 (N_12615,N_11889,N_11972);
nand U12616 (N_12616,N_11762,N_11043);
or U12617 (N_12617,N_11400,N_11332);
or U12618 (N_12618,N_11212,N_11514);
nand U12619 (N_12619,N_11580,N_11216);
nor U12620 (N_12620,N_11438,N_11373);
xnor U12621 (N_12621,N_11359,N_11911);
nor U12622 (N_12622,N_11569,N_11878);
or U12623 (N_12623,N_11765,N_11079);
nor U12624 (N_12624,N_11591,N_11984);
or U12625 (N_12625,N_11247,N_11430);
or U12626 (N_12626,N_11519,N_11522);
xnor U12627 (N_12627,N_11534,N_11376);
xor U12628 (N_12628,N_11459,N_11728);
nor U12629 (N_12629,N_11832,N_11333);
xnor U12630 (N_12630,N_11822,N_11699);
xor U12631 (N_12631,N_11067,N_11782);
or U12632 (N_12632,N_11171,N_11092);
nor U12633 (N_12633,N_11789,N_11203);
or U12634 (N_12634,N_11525,N_11180);
and U12635 (N_12635,N_11142,N_11801);
or U12636 (N_12636,N_11875,N_11878);
nor U12637 (N_12637,N_11396,N_11824);
nand U12638 (N_12638,N_11762,N_11244);
nand U12639 (N_12639,N_11530,N_11105);
and U12640 (N_12640,N_11931,N_11860);
nor U12641 (N_12641,N_11186,N_11759);
nor U12642 (N_12642,N_11313,N_11671);
and U12643 (N_12643,N_11470,N_11107);
nor U12644 (N_12644,N_11365,N_11359);
or U12645 (N_12645,N_11841,N_11217);
nor U12646 (N_12646,N_11946,N_11825);
nor U12647 (N_12647,N_11588,N_11284);
nand U12648 (N_12648,N_11196,N_11010);
xnor U12649 (N_12649,N_11871,N_11916);
nand U12650 (N_12650,N_11882,N_11564);
xor U12651 (N_12651,N_11693,N_11788);
or U12652 (N_12652,N_11380,N_11428);
xnor U12653 (N_12653,N_11927,N_11708);
xnor U12654 (N_12654,N_11446,N_11942);
nor U12655 (N_12655,N_11182,N_11885);
or U12656 (N_12656,N_11386,N_11564);
nor U12657 (N_12657,N_11635,N_11270);
xor U12658 (N_12658,N_11120,N_11069);
nor U12659 (N_12659,N_11662,N_11320);
nor U12660 (N_12660,N_11802,N_11503);
nand U12661 (N_12661,N_11976,N_11954);
and U12662 (N_12662,N_11956,N_11226);
xor U12663 (N_12663,N_11490,N_11292);
or U12664 (N_12664,N_11525,N_11724);
and U12665 (N_12665,N_11225,N_11303);
and U12666 (N_12666,N_11847,N_11272);
and U12667 (N_12667,N_11405,N_11129);
or U12668 (N_12668,N_11866,N_11423);
xnor U12669 (N_12669,N_11418,N_11358);
nor U12670 (N_12670,N_11826,N_11401);
and U12671 (N_12671,N_11198,N_11346);
xor U12672 (N_12672,N_11054,N_11323);
and U12673 (N_12673,N_11962,N_11781);
xor U12674 (N_12674,N_11199,N_11859);
nor U12675 (N_12675,N_11462,N_11392);
or U12676 (N_12676,N_11121,N_11773);
nand U12677 (N_12677,N_11650,N_11148);
nand U12678 (N_12678,N_11169,N_11908);
nor U12679 (N_12679,N_11993,N_11807);
xor U12680 (N_12680,N_11714,N_11443);
or U12681 (N_12681,N_11891,N_11280);
nor U12682 (N_12682,N_11378,N_11441);
and U12683 (N_12683,N_11858,N_11159);
nor U12684 (N_12684,N_11739,N_11151);
nand U12685 (N_12685,N_11799,N_11408);
and U12686 (N_12686,N_11327,N_11188);
or U12687 (N_12687,N_11681,N_11598);
xnor U12688 (N_12688,N_11136,N_11642);
xnor U12689 (N_12689,N_11869,N_11796);
or U12690 (N_12690,N_11099,N_11420);
and U12691 (N_12691,N_11772,N_11335);
nor U12692 (N_12692,N_11971,N_11836);
or U12693 (N_12693,N_11503,N_11140);
or U12694 (N_12694,N_11313,N_11084);
nand U12695 (N_12695,N_11457,N_11787);
and U12696 (N_12696,N_11994,N_11473);
and U12697 (N_12697,N_11243,N_11335);
xor U12698 (N_12698,N_11250,N_11542);
or U12699 (N_12699,N_11559,N_11452);
nor U12700 (N_12700,N_11306,N_11361);
or U12701 (N_12701,N_11967,N_11548);
nor U12702 (N_12702,N_11314,N_11863);
nand U12703 (N_12703,N_11800,N_11912);
nor U12704 (N_12704,N_11921,N_11370);
nand U12705 (N_12705,N_11644,N_11419);
or U12706 (N_12706,N_11602,N_11191);
or U12707 (N_12707,N_11083,N_11248);
nand U12708 (N_12708,N_11484,N_11754);
xnor U12709 (N_12709,N_11440,N_11530);
or U12710 (N_12710,N_11873,N_11731);
and U12711 (N_12711,N_11403,N_11190);
and U12712 (N_12712,N_11404,N_11915);
nor U12713 (N_12713,N_11005,N_11629);
and U12714 (N_12714,N_11770,N_11189);
and U12715 (N_12715,N_11098,N_11972);
nor U12716 (N_12716,N_11854,N_11568);
or U12717 (N_12717,N_11829,N_11221);
nand U12718 (N_12718,N_11980,N_11780);
nand U12719 (N_12719,N_11101,N_11439);
nor U12720 (N_12720,N_11800,N_11000);
nand U12721 (N_12721,N_11666,N_11634);
xnor U12722 (N_12722,N_11367,N_11683);
nand U12723 (N_12723,N_11290,N_11418);
nor U12724 (N_12724,N_11341,N_11948);
or U12725 (N_12725,N_11009,N_11928);
and U12726 (N_12726,N_11987,N_11152);
nor U12727 (N_12727,N_11585,N_11508);
or U12728 (N_12728,N_11360,N_11787);
or U12729 (N_12729,N_11627,N_11436);
xnor U12730 (N_12730,N_11594,N_11549);
and U12731 (N_12731,N_11858,N_11374);
nor U12732 (N_12732,N_11860,N_11781);
and U12733 (N_12733,N_11871,N_11467);
nand U12734 (N_12734,N_11472,N_11477);
xor U12735 (N_12735,N_11101,N_11614);
xor U12736 (N_12736,N_11309,N_11466);
or U12737 (N_12737,N_11828,N_11376);
nor U12738 (N_12738,N_11877,N_11084);
nand U12739 (N_12739,N_11912,N_11410);
or U12740 (N_12740,N_11738,N_11491);
nand U12741 (N_12741,N_11847,N_11452);
or U12742 (N_12742,N_11758,N_11391);
nor U12743 (N_12743,N_11161,N_11418);
and U12744 (N_12744,N_11559,N_11822);
nor U12745 (N_12745,N_11895,N_11279);
nand U12746 (N_12746,N_11280,N_11965);
nor U12747 (N_12747,N_11122,N_11932);
and U12748 (N_12748,N_11894,N_11511);
nand U12749 (N_12749,N_11631,N_11905);
or U12750 (N_12750,N_11223,N_11413);
or U12751 (N_12751,N_11333,N_11759);
or U12752 (N_12752,N_11364,N_11540);
nor U12753 (N_12753,N_11901,N_11550);
xor U12754 (N_12754,N_11543,N_11418);
nand U12755 (N_12755,N_11713,N_11097);
nand U12756 (N_12756,N_11598,N_11118);
and U12757 (N_12757,N_11001,N_11986);
nor U12758 (N_12758,N_11671,N_11632);
and U12759 (N_12759,N_11429,N_11163);
and U12760 (N_12760,N_11463,N_11233);
and U12761 (N_12761,N_11002,N_11180);
or U12762 (N_12762,N_11941,N_11560);
and U12763 (N_12763,N_11320,N_11517);
and U12764 (N_12764,N_11064,N_11352);
or U12765 (N_12765,N_11347,N_11061);
xor U12766 (N_12766,N_11986,N_11623);
xor U12767 (N_12767,N_11881,N_11392);
and U12768 (N_12768,N_11354,N_11478);
xnor U12769 (N_12769,N_11196,N_11318);
nand U12770 (N_12770,N_11683,N_11262);
xnor U12771 (N_12771,N_11933,N_11517);
nand U12772 (N_12772,N_11683,N_11289);
xor U12773 (N_12773,N_11452,N_11851);
and U12774 (N_12774,N_11423,N_11724);
or U12775 (N_12775,N_11469,N_11450);
nand U12776 (N_12776,N_11444,N_11175);
nor U12777 (N_12777,N_11967,N_11005);
and U12778 (N_12778,N_11201,N_11953);
or U12779 (N_12779,N_11418,N_11813);
and U12780 (N_12780,N_11664,N_11032);
nor U12781 (N_12781,N_11314,N_11132);
and U12782 (N_12782,N_11320,N_11376);
xor U12783 (N_12783,N_11930,N_11541);
nand U12784 (N_12784,N_11805,N_11896);
and U12785 (N_12785,N_11306,N_11877);
xor U12786 (N_12786,N_11752,N_11522);
nor U12787 (N_12787,N_11726,N_11280);
or U12788 (N_12788,N_11293,N_11211);
or U12789 (N_12789,N_11969,N_11329);
xnor U12790 (N_12790,N_11644,N_11327);
and U12791 (N_12791,N_11933,N_11467);
nor U12792 (N_12792,N_11897,N_11721);
nand U12793 (N_12793,N_11129,N_11173);
and U12794 (N_12794,N_11570,N_11118);
and U12795 (N_12795,N_11897,N_11916);
or U12796 (N_12796,N_11635,N_11215);
xnor U12797 (N_12797,N_11554,N_11875);
xnor U12798 (N_12798,N_11523,N_11001);
nand U12799 (N_12799,N_11799,N_11867);
xnor U12800 (N_12800,N_11006,N_11021);
nor U12801 (N_12801,N_11113,N_11420);
or U12802 (N_12802,N_11465,N_11606);
and U12803 (N_12803,N_11373,N_11364);
nor U12804 (N_12804,N_11711,N_11995);
or U12805 (N_12805,N_11445,N_11885);
and U12806 (N_12806,N_11320,N_11597);
nand U12807 (N_12807,N_11351,N_11149);
xnor U12808 (N_12808,N_11156,N_11353);
and U12809 (N_12809,N_11164,N_11277);
nand U12810 (N_12810,N_11134,N_11328);
nand U12811 (N_12811,N_11638,N_11983);
nor U12812 (N_12812,N_11991,N_11776);
xnor U12813 (N_12813,N_11112,N_11773);
xnor U12814 (N_12814,N_11250,N_11306);
xnor U12815 (N_12815,N_11429,N_11139);
or U12816 (N_12816,N_11707,N_11393);
and U12817 (N_12817,N_11401,N_11038);
nand U12818 (N_12818,N_11552,N_11025);
and U12819 (N_12819,N_11835,N_11135);
nand U12820 (N_12820,N_11828,N_11469);
nand U12821 (N_12821,N_11025,N_11794);
nor U12822 (N_12822,N_11959,N_11504);
xnor U12823 (N_12823,N_11986,N_11899);
and U12824 (N_12824,N_11375,N_11543);
or U12825 (N_12825,N_11789,N_11139);
and U12826 (N_12826,N_11812,N_11226);
nor U12827 (N_12827,N_11401,N_11477);
xnor U12828 (N_12828,N_11786,N_11097);
and U12829 (N_12829,N_11756,N_11983);
or U12830 (N_12830,N_11526,N_11600);
and U12831 (N_12831,N_11701,N_11848);
nor U12832 (N_12832,N_11911,N_11091);
or U12833 (N_12833,N_11078,N_11883);
nor U12834 (N_12834,N_11449,N_11804);
nand U12835 (N_12835,N_11855,N_11491);
xnor U12836 (N_12836,N_11133,N_11321);
xnor U12837 (N_12837,N_11183,N_11837);
and U12838 (N_12838,N_11235,N_11293);
and U12839 (N_12839,N_11129,N_11994);
nor U12840 (N_12840,N_11412,N_11205);
nor U12841 (N_12841,N_11847,N_11888);
or U12842 (N_12842,N_11185,N_11434);
nand U12843 (N_12843,N_11685,N_11014);
nand U12844 (N_12844,N_11038,N_11725);
or U12845 (N_12845,N_11248,N_11933);
nor U12846 (N_12846,N_11132,N_11331);
xnor U12847 (N_12847,N_11284,N_11406);
nor U12848 (N_12848,N_11496,N_11458);
or U12849 (N_12849,N_11380,N_11086);
nand U12850 (N_12850,N_11435,N_11675);
or U12851 (N_12851,N_11860,N_11043);
xnor U12852 (N_12852,N_11186,N_11174);
xor U12853 (N_12853,N_11331,N_11579);
and U12854 (N_12854,N_11052,N_11313);
xor U12855 (N_12855,N_11869,N_11228);
or U12856 (N_12856,N_11925,N_11247);
nand U12857 (N_12857,N_11657,N_11150);
xnor U12858 (N_12858,N_11676,N_11856);
nor U12859 (N_12859,N_11757,N_11511);
nand U12860 (N_12860,N_11813,N_11171);
xnor U12861 (N_12861,N_11756,N_11913);
xnor U12862 (N_12862,N_11936,N_11530);
nand U12863 (N_12863,N_11277,N_11987);
nor U12864 (N_12864,N_11465,N_11170);
and U12865 (N_12865,N_11799,N_11510);
or U12866 (N_12866,N_11794,N_11590);
or U12867 (N_12867,N_11279,N_11582);
nand U12868 (N_12868,N_11082,N_11378);
and U12869 (N_12869,N_11179,N_11260);
xor U12870 (N_12870,N_11357,N_11236);
nand U12871 (N_12871,N_11823,N_11035);
and U12872 (N_12872,N_11710,N_11992);
and U12873 (N_12873,N_11622,N_11456);
xnor U12874 (N_12874,N_11052,N_11748);
and U12875 (N_12875,N_11517,N_11909);
or U12876 (N_12876,N_11838,N_11473);
xnor U12877 (N_12877,N_11108,N_11241);
nor U12878 (N_12878,N_11609,N_11237);
nand U12879 (N_12879,N_11156,N_11143);
xor U12880 (N_12880,N_11643,N_11206);
nand U12881 (N_12881,N_11175,N_11257);
nor U12882 (N_12882,N_11543,N_11502);
xnor U12883 (N_12883,N_11986,N_11365);
nor U12884 (N_12884,N_11440,N_11508);
or U12885 (N_12885,N_11889,N_11684);
or U12886 (N_12886,N_11997,N_11655);
or U12887 (N_12887,N_11449,N_11630);
or U12888 (N_12888,N_11422,N_11471);
or U12889 (N_12889,N_11140,N_11641);
nor U12890 (N_12890,N_11987,N_11113);
or U12891 (N_12891,N_11015,N_11152);
and U12892 (N_12892,N_11791,N_11998);
or U12893 (N_12893,N_11386,N_11586);
or U12894 (N_12894,N_11867,N_11286);
and U12895 (N_12895,N_11667,N_11185);
or U12896 (N_12896,N_11708,N_11984);
xnor U12897 (N_12897,N_11659,N_11191);
nand U12898 (N_12898,N_11957,N_11538);
nand U12899 (N_12899,N_11762,N_11292);
and U12900 (N_12900,N_11680,N_11704);
nand U12901 (N_12901,N_11700,N_11902);
or U12902 (N_12902,N_11049,N_11255);
or U12903 (N_12903,N_11937,N_11746);
nor U12904 (N_12904,N_11566,N_11288);
nand U12905 (N_12905,N_11157,N_11300);
or U12906 (N_12906,N_11195,N_11100);
xnor U12907 (N_12907,N_11520,N_11394);
nor U12908 (N_12908,N_11810,N_11715);
and U12909 (N_12909,N_11786,N_11175);
xnor U12910 (N_12910,N_11296,N_11941);
xor U12911 (N_12911,N_11484,N_11775);
nand U12912 (N_12912,N_11594,N_11099);
or U12913 (N_12913,N_11540,N_11548);
and U12914 (N_12914,N_11928,N_11243);
and U12915 (N_12915,N_11546,N_11542);
and U12916 (N_12916,N_11730,N_11782);
nor U12917 (N_12917,N_11654,N_11602);
xnor U12918 (N_12918,N_11781,N_11557);
xor U12919 (N_12919,N_11745,N_11098);
nand U12920 (N_12920,N_11435,N_11964);
or U12921 (N_12921,N_11729,N_11402);
nand U12922 (N_12922,N_11925,N_11419);
nor U12923 (N_12923,N_11230,N_11474);
nor U12924 (N_12924,N_11229,N_11727);
xor U12925 (N_12925,N_11214,N_11306);
and U12926 (N_12926,N_11565,N_11154);
nand U12927 (N_12927,N_11456,N_11579);
and U12928 (N_12928,N_11337,N_11436);
nand U12929 (N_12929,N_11821,N_11456);
or U12930 (N_12930,N_11304,N_11154);
or U12931 (N_12931,N_11410,N_11789);
nor U12932 (N_12932,N_11108,N_11462);
and U12933 (N_12933,N_11177,N_11425);
nand U12934 (N_12934,N_11597,N_11569);
and U12935 (N_12935,N_11663,N_11434);
xnor U12936 (N_12936,N_11033,N_11018);
nand U12937 (N_12937,N_11322,N_11919);
nand U12938 (N_12938,N_11747,N_11745);
nand U12939 (N_12939,N_11378,N_11642);
nand U12940 (N_12940,N_11407,N_11951);
nand U12941 (N_12941,N_11205,N_11889);
nand U12942 (N_12942,N_11508,N_11971);
nand U12943 (N_12943,N_11875,N_11594);
nor U12944 (N_12944,N_11391,N_11826);
and U12945 (N_12945,N_11228,N_11962);
xnor U12946 (N_12946,N_11308,N_11726);
xor U12947 (N_12947,N_11449,N_11323);
xor U12948 (N_12948,N_11423,N_11801);
or U12949 (N_12949,N_11255,N_11448);
nand U12950 (N_12950,N_11213,N_11564);
or U12951 (N_12951,N_11023,N_11895);
nand U12952 (N_12952,N_11735,N_11058);
nor U12953 (N_12953,N_11044,N_11022);
and U12954 (N_12954,N_11664,N_11549);
and U12955 (N_12955,N_11972,N_11127);
xor U12956 (N_12956,N_11148,N_11938);
nand U12957 (N_12957,N_11542,N_11716);
or U12958 (N_12958,N_11368,N_11886);
xor U12959 (N_12959,N_11283,N_11274);
xnor U12960 (N_12960,N_11043,N_11237);
and U12961 (N_12961,N_11861,N_11180);
nor U12962 (N_12962,N_11999,N_11948);
or U12963 (N_12963,N_11966,N_11951);
or U12964 (N_12964,N_11914,N_11438);
or U12965 (N_12965,N_11295,N_11294);
or U12966 (N_12966,N_11874,N_11537);
nor U12967 (N_12967,N_11522,N_11115);
nor U12968 (N_12968,N_11372,N_11378);
or U12969 (N_12969,N_11197,N_11552);
and U12970 (N_12970,N_11710,N_11152);
and U12971 (N_12971,N_11576,N_11086);
nand U12972 (N_12972,N_11471,N_11213);
and U12973 (N_12973,N_11395,N_11583);
xor U12974 (N_12974,N_11752,N_11887);
xor U12975 (N_12975,N_11966,N_11101);
and U12976 (N_12976,N_11029,N_11821);
xnor U12977 (N_12977,N_11884,N_11068);
xnor U12978 (N_12978,N_11654,N_11488);
and U12979 (N_12979,N_11199,N_11910);
nor U12980 (N_12980,N_11808,N_11072);
and U12981 (N_12981,N_11517,N_11862);
or U12982 (N_12982,N_11715,N_11545);
nor U12983 (N_12983,N_11218,N_11791);
nand U12984 (N_12984,N_11763,N_11907);
nor U12985 (N_12985,N_11364,N_11704);
nor U12986 (N_12986,N_11591,N_11278);
nor U12987 (N_12987,N_11404,N_11936);
nand U12988 (N_12988,N_11231,N_11204);
nand U12989 (N_12989,N_11601,N_11321);
and U12990 (N_12990,N_11571,N_11444);
or U12991 (N_12991,N_11205,N_11692);
xnor U12992 (N_12992,N_11955,N_11793);
and U12993 (N_12993,N_11563,N_11047);
and U12994 (N_12994,N_11241,N_11920);
or U12995 (N_12995,N_11401,N_11464);
nor U12996 (N_12996,N_11295,N_11298);
and U12997 (N_12997,N_11378,N_11360);
or U12998 (N_12998,N_11237,N_11945);
and U12999 (N_12999,N_11965,N_11086);
nor U13000 (N_13000,N_12987,N_12514);
or U13001 (N_13001,N_12474,N_12612);
xnor U13002 (N_13002,N_12685,N_12969);
or U13003 (N_13003,N_12870,N_12505);
or U13004 (N_13004,N_12980,N_12196);
nor U13005 (N_13005,N_12486,N_12169);
xnor U13006 (N_13006,N_12047,N_12974);
nand U13007 (N_13007,N_12268,N_12271);
and U13008 (N_13008,N_12761,N_12684);
nand U13009 (N_13009,N_12831,N_12602);
nand U13010 (N_13010,N_12719,N_12640);
and U13011 (N_13011,N_12305,N_12093);
and U13012 (N_13012,N_12767,N_12226);
and U13013 (N_13013,N_12130,N_12478);
or U13014 (N_13014,N_12187,N_12195);
xor U13015 (N_13015,N_12119,N_12067);
nor U13016 (N_13016,N_12725,N_12429);
xor U13017 (N_13017,N_12989,N_12132);
and U13018 (N_13018,N_12356,N_12006);
or U13019 (N_13019,N_12787,N_12515);
or U13020 (N_13020,N_12216,N_12586);
xor U13021 (N_13021,N_12708,N_12524);
nor U13022 (N_13022,N_12701,N_12774);
xnor U13023 (N_13023,N_12802,N_12583);
and U13024 (N_13024,N_12202,N_12975);
nor U13025 (N_13025,N_12882,N_12318);
xnor U13026 (N_13026,N_12888,N_12168);
xnor U13027 (N_13027,N_12872,N_12957);
nand U13028 (N_13028,N_12278,N_12698);
and U13029 (N_13029,N_12813,N_12471);
nor U13030 (N_13030,N_12864,N_12080);
nor U13031 (N_13031,N_12150,N_12186);
nand U13032 (N_13032,N_12741,N_12308);
xor U13033 (N_13033,N_12376,N_12727);
or U13034 (N_13034,N_12798,N_12823);
or U13035 (N_13035,N_12898,N_12479);
nor U13036 (N_13036,N_12952,N_12419);
xor U13037 (N_13037,N_12559,N_12424);
xnor U13038 (N_13038,N_12073,N_12133);
and U13039 (N_13039,N_12814,N_12796);
and U13040 (N_13040,N_12282,N_12921);
nand U13041 (N_13041,N_12103,N_12311);
nor U13042 (N_13042,N_12615,N_12136);
or U13043 (N_13043,N_12634,N_12074);
nand U13044 (N_13044,N_12241,N_12214);
nand U13045 (N_13045,N_12225,N_12248);
nor U13046 (N_13046,N_12060,N_12812);
xor U13047 (N_13047,N_12387,N_12222);
nand U13048 (N_13048,N_12807,N_12569);
nand U13049 (N_13049,N_12404,N_12631);
xnor U13050 (N_13050,N_12999,N_12686);
or U13051 (N_13051,N_12399,N_12899);
and U13052 (N_13052,N_12673,N_12843);
nand U13053 (N_13053,N_12726,N_12373);
nor U13054 (N_13054,N_12537,N_12525);
or U13055 (N_13055,N_12317,N_12238);
or U13056 (N_13056,N_12852,N_12639);
xor U13057 (N_13057,N_12721,N_12031);
nor U13058 (N_13058,N_12897,N_12599);
nand U13059 (N_13059,N_12914,N_12100);
nor U13060 (N_13060,N_12942,N_12454);
nand U13061 (N_13061,N_12094,N_12160);
and U13062 (N_13062,N_12797,N_12502);
and U13063 (N_13063,N_12344,N_12688);
nand U13064 (N_13064,N_12061,N_12265);
nand U13065 (N_13065,N_12492,N_12617);
or U13066 (N_13066,N_12346,N_12841);
nand U13067 (N_13067,N_12664,N_12995);
or U13068 (N_13068,N_12567,N_12484);
xnor U13069 (N_13069,N_12778,N_12626);
xor U13070 (N_13070,N_12013,N_12303);
or U13071 (N_13071,N_12333,N_12704);
xnor U13072 (N_13072,N_12397,N_12585);
or U13073 (N_13073,N_12923,N_12218);
nor U13074 (N_13074,N_12712,N_12827);
and U13075 (N_13075,N_12293,N_12577);
or U13076 (N_13076,N_12945,N_12543);
xor U13077 (N_13077,N_12352,N_12944);
or U13078 (N_13078,N_12855,N_12190);
nand U13079 (N_13079,N_12723,N_12326);
nor U13080 (N_13080,N_12476,N_12710);
nor U13081 (N_13081,N_12157,N_12242);
nor U13082 (N_13082,N_12371,N_12752);
nand U13083 (N_13083,N_12233,N_12811);
and U13084 (N_13084,N_12635,N_12620);
nor U13085 (N_13085,N_12739,N_12402);
nor U13086 (N_13086,N_12354,N_12596);
and U13087 (N_13087,N_12724,N_12536);
and U13088 (N_13088,N_12732,N_12267);
and U13089 (N_13089,N_12637,N_12744);
nor U13090 (N_13090,N_12877,N_12571);
xor U13091 (N_13091,N_12264,N_12188);
xnor U13092 (N_13092,N_12319,N_12603);
nand U13093 (N_13093,N_12057,N_12258);
nand U13094 (N_13094,N_12205,N_12842);
nor U13095 (N_13095,N_12137,N_12667);
and U13096 (N_13096,N_12269,N_12309);
nand U13097 (N_13097,N_12895,N_12192);
nor U13098 (N_13098,N_12351,N_12947);
or U13099 (N_13099,N_12290,N_12117);
and U13100 (N_13100,N_12489,N_12754);
xnor U13101 (N_13101,N_12693,N_12388);
or U13102 (N_13102,N_12528,N_12716);
nor U13103 (N_13103,N_12553,N_12848);
nor U13104 (N_13104,N_12825,N_12237);
nor U13105 (N_13105,N_12772,N_12678);
and U13106 (N_13106,N_12223,N_12917);
nor U13107 (N_13107,N_12343,N_12535);
nand U13108 (N_13108,N_12792,N_12621);
nor U13109 (N_13109,N_12874,N_12102);
and U13110 (N_13110,N_12370,N_12682);
nand U13111 (N_13111,N_12036,N_12353);
xor U13112 (N_13112,N_12003,N_12277);
nand U13113 (N_13113,N_12506,N_12081);
xnor U13114 (N_13114,N_12367,N_12624);
nand U13115 (N_13115,N_12784,N_12089);
xnor U13116 (N_13116,N_12283,N_12949);
and U13117 (N_13117,N_12126,N_12611);
xor U13118 (N_13118,N_12208,N_12955);
xnor U13119 (N_13119,N_12885,N_12022);
and U13120 (N_13120,N_12614,N_12856);
nor U13121 (N_13121,N_12289,N_12322);
or U13122 (N_13122,N_12288,N_12138);
and U13123 (N_13123,N_12206,N_12307);
xor U13124 (N_13124,N_12412,N_12876);
nor U13125 (N_13125,N_12950,N_12445);
or U13126 (N_13126,N_12581,N_12135);
nor U13127 (N_13127,N_12517,N_12433);
nor U13128 (N_13128,N_12737,N_12016);
nand U13129 (N_13129,N_12951,N_12927);
nor U13130 (N_13130,N_12526,N_12253);
nor U13131 (N_13131,N_12240,N_12275);
nor U13132 (N_13132,N_12751,N_12560);
nor U13133 (N_13133,N_12015,N_12211);
or U13134 (N_13134,N_12722,N_12042);
and U13135 (N_13135,N_12155,N_12665);
and U13136 (N_13136,N_12879,N_12762);
nand U13137 (N_13137,N_12257,N_12279);
nand U13138 (N_13138,N_12391,N_12312);
xnor U13139 (N_13139,N_12436,N_12558);
and U13140 (N_13140,N_12795,N_12996);
or U13141 (N_13141,N_12111,N_12799);
and U13142 (N_13142,N_12636,N_12608);
xnor U13143 (N_13143,N_12859,N_12830);
or U13144 (N_13144,N_12504,N_12591);
nor U13145 (N_13145,N_12134,N_12541);
nand U13146 (N_13146,N_12368,N_12301);
and U13147 (N_13147,N_12758,N_12338);
or U13148 (N_13148,N_12193,N_12925);
and U13149 (N_13149,N_12260,N_12456);
xor U13150 (N_13150,N_12007,N_12284);
nor U13151 (N_13151,N_12437,N_12400);
nor U13152 (N_13152,N_12200,N_12452);
and U13153 (N_13153,N_12262,N_12418);
or U13154 (N_13154,N_12972,N_12958);
nor U13155 (N_13155,N_12121,N_12129);
and U13156 (N_13156,N_12125,N_12442);
or U13157 (N_13157,N_12025,N_12116);
or U13158 (N_13158,N_12033,N_12491);
nand U13159 (N_13159,N_12444,N_12713);
and U13160 (N_13160,N_12450,N_12998);
and U13161 (N_13161,N_12887,N_12295);
or U13162 (N_13162,N_12315,N_12058);
nor U13163 (N_13163,N_12820,N_12853);
nor U13164 (N_13164,N_12669,N_12959);
and U13165 (N_13165,N_12858,N_12764);
nand U13166 (N_13166,N_12847,N_12824);
and U13167 (N_13167,N_12236,N_12689);
and U13168 (N_13168,N_12646,N_12156);
nor U13169 (N_13169,N_12970,N_12203);
nand U13170 (N_13170,N_12838,N_12546);
or U13171 (N_13171,N_12728,N_12485);
xnor U13172 (N_13172,N_12234,N_12177);
xor U13173 (N_13173,N_12300,N_12781);
nor U13174 (N_13174,N_12334,N_12670);
xor U13175 (N_13175,N_12935,N_12922);
nor U13176 (N_13176,N_12041,N_12556);
nor U13177 (N_13177,N_12549,N_12964);
nand U13178 (N_13178,N_12413,N_12576);
and U13179 (N_13179,N_12176,N_12050);
xnor U13180 (N_13180,N_12566,N_12868);
and U13181 (N_13181,N_12372,N_12747);
and U13182 (N_13182,N_12361,N_12916);
nor U13183 (N_13183,N_12377,N_12512);
nand U13184 (N_13184,N_12034,N_12336);
nor U13185 (N_13185,N_12630,N_12229);
nor U13186 (N_13186,N_12490,N_12776);
nand U13187 (N_13187,N_12940,N_12750);
nand U13188 (N_13188,N_12092,N_12616);
or U13189 (N_13189,N_12956,N_12893);
nand U13190 (N_13190,N_12963,N_12421);
and U13191 (N_13191,N_12742,N_12829);
or U13192 (N_13192,N_12846,N_12481);
xnor U13193 (N_13193,N_12840,N_12244);
nor U13194 (N_13194,N_12984,N_12349);
nor U13195 (N_13195,N_12816,N_12106);
or U13196 (N_13196,N_12965,N_12869);
and U13197 (N_13197,N_12551,N_12532);
and U13198 (N_13198,N_12018,N_12627);
or U13199 (N_13199,N_12906,N_12901);
and U13200 (N_13200,N_12523,N_12008);
nand U13201 (N_13201,N_12801,N_12185);
and U13202 (N_13202,N_12574,N_12066);
nand U13203 (N_13203,N_12329,N_12657);
nor U13204 (N_13204,N_12065,N_12118);
nor U13205 (N_13205,N_12903,N_12409);
xnor U13206 (N_13206,N_12280,N_12194);
nand U13207 (N_13207,N_12494,N_12509);
xnor U13208 (N_13208,N_12335,N_12513);
xor U13209 (N_13209,N_12120,N_12276);
and U13210 (N_13210,N_12930,N_12651);
xor U13211 (N_13211,N_12932,N_12172);
xor U13212 (N_13212,N_12518,N_12470);
and U13213 (N_13213,N_12755,N_12393);
and U13214 (N_13214,N_12162,N_12228);
or U13215 (N_13215,N_12466,N_12961);
or U13216 (N_13216,N_12681,N_12939);
xnor U13217 (N_13217,N_12976,N_12141);
or U13218 (N_13218,N_12604,N_12497);
and U13219 (N_13219,N_12587,N_12522);
or U13220 (N_13220,N_12866,N_12675);
and U13221 (N_13221,N_12913,N_12625);
or U13222 (N_13222,N_12565,N_12731);
nor U13223 (N_13223,N_12662,N_12108);
or U13224 (N_13224,N_12337,N_12407);
nor U13225 (N_13225,N_12316,N_12966);
or U13226 (N_13226,N_12428,N_12451);
xnor U13227 (N_13227,N_12147,N_12729);
or U13228 (N_13228,N_12836,N_12467);
nand U13229 (N_13229,N_12482,N_12423);
nor U13230 (N_13230,N_12589,N_12339);
xnor U13231 (N_13231,N_12032,N_12871);
nor U13232 (N_13232,N_12676,N_12562);
and U13233 (N_13233,N_12235,N_12706);
and U13234 (N_13234,N_12915,N_12642);
xnor U13235 (N_13235,N_12937,N_12068);
nand U13236 (N_13236,N_12496,N_12993);
nand U13237 (N_13237,N_12886,N_12910);
xor U13238 (N_13238,N_12692,N_12691);
nand U13239 (N_13239,N_12516,N_12374);
nor U13240 (N_13240,N_12891,N_12212);
or U13241 (N_13241,N_12540,N_12900);
or U13242 (N_13242,N_12904,N_12341);
xnor U13243 (N_13243,N_12826,N_12062);
or U13244 (N_13244,N_12143,N_12833);
xnor U13245 (N_13245,N_12148,N_12573);
or U13246 (N_13246,N_12191,N_12325);
or U13247 (N_13247,N_12817,N_12076);
nor U13248 (N_13248,N_12063,N_12656);
nor U13249 (N_13249,N_12189,N_12793);
and U13250 (N_13250,N_12382,N_12358);
and U13251 (N_13251,N_12531,N_12593);
nand U13252 (N_13252,N_12668,N_12170);
nand U13253 (N_13253,N_12046,N_12239);
xnor U13254 (N_13254,N_12294,N_12839);
nor U13255 (N_13255,N_12821,N_12345);
nand U13256 (N_13256,N_12366,N_12035);
and U13257 (N_13257,N_12458,N_12340);
nand U13258 (N_13258,N_12746,N_12079);
xor U13259 (N_13259,N_12991,N_12666);
or U13260 (N_13260,N_12590,N_12714);
and U13261 (N_13261,N_12968,N_12483);
nand U13262 (N_13262,N_12861,N_12173);
or U13263 (N_13263,N_12461,N_12112);
nor U13264 (N_13264,N_12123,N_12997);
nand U13265 (N_13265,N_12263,N_12849);
xor U13266 (N_13266,N_12931,N_12430);
or U13267 (N_13267,N_12435,N_12809);
xor U13268 (N_13268,N_12398,N_12889);
xnor U13269 (N_13269,N_12113,N_12149);
and U13270 (N_13270,N_12447,N_12197);
nor U13271 (N_13271,N_12250,N_12417);
nand U13272 (N_13272,N_12142,N_12232);
and U13273 (N_13273,N_12605,N_12053);
nor U13274 (N_13274,N_12440,N_12894);
xor U13275 (N_13275,N_12702,N_12002);
nor U13276 (N_13276,N_12028,N_12270);
nor U13277 (N_13277,N_12380,N_12570);
or U13278 (N_13278,N_12672,N_12777);
or U13279 (N_13279,N_12355,N_12564);
or U13280 (N_13280,N_12677,N_12324);
and U13281 (N_13281,N_12039,N_12427);
nor U13282 (N_13282,N_12804,N_12198);
or U13283 (N_13283,N_12055,N_12365);
nand U13284 (N_13284,N_12740,N_12563);
xor U13285 (N_13285,N_12694,N_12510);
or U13286 (N_13286,N_12711,N_12643);
and U13287 (N_13287,N_12633,N_12071);
or U13288 (N_13288,N_12507,N_12070);
and U13289 (N_13289,N_12806,N_12401);
nor U13290 (N_13290,N_12568,N_12153);
or U13291 (N_13291,N_12863,N_12629);
nand U13292 (N_13292,N_12166,N_12215);
nor U13293 (N_13293,N_12994,N_12773);
and U13294 (N_13294,N_12285,N_12896);
nand U13295 (N_13295,N_12539,N_12680);
and U13296 (N_13296,N_12674,N_12363);
or U13297 (N_13297,N_12822,N_12151);
or U13298 (N_13298,N_12499,N_12273);
or U13299 (N_13299,N_12431,N_12707);
nor U13300 (N_13300,N_12908,N_12828);
nor U13301 (N_13301,N_12310,N_12037);
nand U13302 (N_13302,N_12131,N_12029);
nor U13303 (N_13303,N_12010,N_12128);
xor U13304 (N_13304,N_12385,N_12231);
nand U13305 (N_13305,N_12146,N_12099);
nand U13306 (N_13306,N_12054,N_12395);
xor U13307 (N_13307,N_12544,N_12109);
nand U13308 (N_13308,N_12928,N_12052);
nand U13309 (N_13309,N_12648,N_12019);
and U13310 (N_13310,N_12655,N_12511);
or U13311 (N_13311,N_12297,N_12924);
nor U13312 (N_13312,N_12632,N_12983);
or U13313 (N_13313,N_12455,N_12808);
and U13314 (N_13314,N_12127,N_12375);
nor U13315 (N_13315,N_12299,N_12446);
and U13316 (N_13316,N_12075,N_12249);
xor U13317 (N_13317,N_12703,N_12800);
xor U13318 (N_13318,N_12919,N_12459);
and U13319 (N_13319,N_12520,N_12790);
nand U13320 (N_13320,N_12867,N_12059);
nor U13321 (N_13321,N_12696,N_12503);
and U13322 (N_13322,N_12292,N_12005);
xnor U13323 (N_13323,N_12152,N_12579);
nand U13324 (N_13324,N_12323,N_12521);
nand U13325 (N_13325,N_12770,N_12815);
or U13326 (N_13326,N_12415,N_12938);
nand U13327 (N_13327,N_12224,N_12392);
nand U13328 (N_13328,N_12905,N_12769);
and U13329 (N_13329,N_12735,N_12654);
and U13330 (N_13330,N_12488,N_12911);
nor U13331 (N_13331,N_12001,N_12749);
nor U13332 (N_13332,N_12139,N_12012);
nand U13333 (N_13333,N_12199,N_12743);
or U13334 (N_13334,N_12881,N_12548);
or U13335 (N_13335,N_12406,N_12165);
or U13336 (N_13336,N_12783,N_12227);
nand U13337 (N_13337,N_12962,N_12663);
xor U13338 (N_13338,N_12441,N_12607);
or U13339 (N_13339,N_12687,N_12545);
nor U13340 (N_13340,N_12718,N_12953);
and U13341 (N_13341,N_12943,N_12408);
nand U13342 (N_13342,N_12394,N_12246);
and U13343 (N_13343,N_12933,N_12048);
and U13344 (N_13344,N_12088,N_12462);
or U13345 (N_13345,N_12175,N_12348);
xor U13346 (N_13346,N_12990,N_12878);
or U13347 (N_13347,N_12946,N_12086);
nand U13348 (N_13348,N_12845,N_12085);
xnor U13349 (N_13349,N_12658,N_12645);
or U13350 (N_13350,N_12973,N_12313);
nand U13351 (N_13351,N_12087,N_12369);
nand U13352 (N_13352,N_12217,N_12107);
nand U13353 (N_13353,N_12463,N_12328);
and U13354 (N_13354,N_12929,N_12552);
and U13355 (N_13355,N_12542,N_12439);
nor U13356 (N_13356,N_12298,N_12768);
or U13357 (N_13357,N_12164,N_12835);
or U13358 (N_13358,N_12738,N_12347);
and U13359 (N_13359,N_12056,N_12763);
nor U13360 (N_13360,N_12644,N_12434);
and U13361 (N_13361,N_12892,N_12251);
or U13362 (N_13362,N_12803,N_12850);
nor U13363 (N_13363,N_12396,N_12272);
or U13364 (N_13364,N_12095,N_12122);
and U13365 (N_13365,N_12557,N_12017);
and U13366 (N_13366,N_12660,N_12912);
nand U13367 (N_13367,N_12104,N_12572);
nand U13368 (N_13368,N_12247,N_12971);
xnor U13369 (N_13369,N_12844,N_12043);
nand U13370 (N_13370,N_12771,N_12389);
or U13371 (N_13371,N_12049,N_12259);
xor U13372 (N_13372,N_12105,N_12159);
nor U13373 (N_13373,N_12554,N_12954);
or U13374 (N_13374,N_12533,N_12291);
and U13375 (N_13375,N_12880,N_12204);
xor U13376 (N_13376,N_12873,N_12145);
or U13377 (N_13377,N_12473,N_12810);
nand U13378 (N_13378,N_12985,N_12083);
xor U13379 (N_13379,N_12530,N_12302);
and U13380 (N_13380,N_12000,N_12628);
and U13381 (N_13381,N_12851,N_12760);
nor U13382 (N_13382,N_12487,N_12734);
nor U13383 (N_13383,N_12786,N_12219);
or U13384 (N_13384,N_12287,N_12582);
nor U13385 (N_13385,N_12026,N_12992);
xor U13386 (N_13386,N_12171,N_12306);
or U13387 (N_13387,N_12834,N_12432);
xnor U13388 (N_13388,N_12449,N_12154);
or U13389 (N_13389,N_12296,N_12243);
or U13390 (N_13390,N_12378,N_12027);
nor U13391 (N_13391,N_12183,N_12819);
nand U13392 (N_13392,N_12865,N_12805);
nand U13393 (N_13393,N_12756,N_12044);
xnor U13394 (N_13394,N_12715,N_12321);
and U13395 (N_13395,N_12020,N_12788);
nand U13396 (N_13396,N_12619,N_12332);
or U13397 (N_13397,N_12926,N_12578);
xor U13398 (N_13398,N_12304,N_12084);
xnor U13399 (N_13399,N_12004,N_12469);
xnor U13400 (N_13400,N_12534,N_12350);
and U13401 (N_13401,N_12832,N_12671);
nor U13402 (N_13402,N_12457,N_12072);
nand U13403 (N_13403,N_12979,N_12230);
xor U13404 (N_13404,N_12178,N_12717);
nor U13405 (N_13405,N_12606,N_12884);
nand U13406 (N_13406,N_12386,N_12420);
nor U13407 (N_13407,N_12918,N_12038);
and U13408 (N_13408,N_12699,N_12405);
nor U13409 (N_13409,N_12857,N_12320);
nor U13410 (N_13410,N_12330,N_12045);
xor U13411 (N_13411,N_12281,N_12220);
nand U13412 (N_13412,N_12201,N_12213);
and U13413 (N_13413,N_12410,N_12261);
or U13414 (N_13414,N_12091,N_12221);
and U13415 (N_13415,N_12623,N_12064);
nand U13416 (N_13416,N_12609,N_12818);
nor U13417 (N_13417,N_12077,N_12453);
xor U13418 (N_13418,N_12697,N_12357);
xnor U13419 (N_13419,N_12286,N_12659);
and U13420 (N_13420,N_12519,N_12854);
and U13421 (N_13421,N_12791,N_12759);
or U13422 (N_13422,N_12598,N_12575);
nor U13423 (N_13423,N_12101,N_12595);
or U13424 (N_13424,N_12948,N_12592);
xor U13425 (N_13425,N_12981,N_12890);
or U13426 (N_13426,N_12647,N_12601);
nor U13427 (N_13427,N_12733,N_12529);
xnor U13428 (N_13428,N_12547,N_12096);
and U13429 (N_13429,N_12179,N_12837);
xor U13430 (N_13430,N_12014,N_12360);
and U13431 (N_13431,N_12023,N_12690);
nand U13432 (N_13432,N_12789,N_12794);
xnor U13433 (N_13433,N_12051,N_12140);
xor U13434 (N_13434,N_12766,N_12584);
or U13435 (N_13435,N_12757,N_12683);
nor U13436 (N_13436,N_12941,N_12909);
nand U13437 (N_13437,N_12425,N_12438);
and U13438 (N_13438,N_12465,N_12069);
nor U13439 (N_13439,N_12362,N_12254);
and U13440 (N_13440,N_12021,N_12753);
and U13441 (N_13441,N_12650,N_12098);
or U13442 (N_13442,N_12936,N_12460);
nor U13443 (N_13443,N_12765,N_12695);
and U13444 (N_13444,N_12009,N_12390);
xor U13445 (N_13445,N_12314,N_12653);
xor U13446 (N_13446,N_12477,N_12468);
xor U13447 (N_13447,N_12161,N_12167);
nand U13448 (N_13448,N_12090,N_12907);
or U13449 (N_13449,N_12610,N_12082);
xnor U13450 (N_13450,N_12383,N_12252);
nor U13451 (N_13451,N_12780,N_12245);
or U13452 (N_13452,N_12745,N_12414);
and U13453 (N_13453,N_12207,N_12158);
nor U13454 (N_13454,N_12498,N_12030);
xnor U13455 (N_13455,N_12403,N_12527);
nand U13456 (N_13456,N_12594,N_12988);
nor U13457 (N_13457,N_12555,N_12274);
nand U13458 (N_13458,N_12184,N_12124);
nor U13459 (N_13459,N_12011,N_12618);
and U13460 (N_13460,N_12097,N_12779);
and U13461 (N_13461,N_12209,N_12597);
or U13462 (N_13462,N_12256,N_12652);
nor U13463 (N_13463,N_12480,N_12883);
xor U13464 (N_13464,N_12649,N_12210);
nand U13465 (N_13465,N_12641,N_12359);
and U13466 (N_13466,N_12182,N_12679);
nand U13467 (N_13467,N_12720,N_12342);
or U13468 (N_13468,N_12416,N_12934);
xor U13469 (N_13469,N_12475,N_12902);
or U13470 (N_13470,N_12782,N_12588);
and U13471 (N_13471,N_12144,N_12967);
nor U13472 (N_13472,N_12730,N_12364);
xor U13473 (N_13473,N_12977,N_12550);
nor U13474 (N_13474,N_12613,N_12862);
or U13475 (N_13475,N_12174,N_12709);
and U13476 (N_13476,N_12181,N_12622);
or U13477 (N_13477,N_12561,N_12700);
and U13478 (N_13478,N_12114,N_12785);
xor U13479 (N_13479,N_12327,N_12493);
and U13480 (N_13480,N_12448,N_12384);
and U13481 (N_13481,N_12040,N_12422);
nand U13482 (N_13482,N_12464,N_12860);
nor U13483 (N_13483,N_12501,N_12600);
and U13484 (N_13484,N_12508,N_12411);
nand U13485 (N_13485,N_12331,N_12426);
or U13486 (N_13486,N_12538,N_12638);
and U13487 (N_13487,N_12748,N_12255);
nand U13488 (N_13488,N_12110,N_12705);
nand U13489 (N_13489,N_12379,N_12163);
xor U13490 (N_13490,N_12661,N_12472);
nor U13491 (N_13491,N_12500,N_12495);
and U13492 (N_13492,N_12982,N_12443);
and U13493 (N_13493,N_12875,N_12180);
xor U13494 (N_13494,N_12978,N_12266);
nor U13495 (N_13495,N_12775,N_12078);
and U13496 (N_13496,N_12580,N_12920);
nand U13497 (N_13497,N_12960,N_12115);
and U13498 (N_13498,N_12986,N_12736);
xor U13499 (N_13499,N_12381,N_12024);
or U13500 (N_13500,N_12013,N_12944);
nand U13501 (N_13501,N_12116,N_12418);
xnor U13502 (N_13502,N_12934,N_12779);
xor U13503 (N_13503,N_12805,N_12736);
nor U13504 (N_13504,N_12536,N_12579);
xor U13505 (N_13505,N_12632,N_12880);
and U13506 (N_13506,N_12711,N_12835);
nand U13507 (N_13507,N_12694,N_12337);
and U13508 (N_13508,N_12429,N_12351);
nor U13509 (N_13509,N_12399,N_12815);
nor U13510 (N_13510,N_12978,N_12317);
or U13511 (N_13511,N_12576,N_12286);
nor U13512 (N_13512,N_12139,N_12930);
nor U13513 (N_13513,N_12890,N_12169);
xor U13514 (N_13514,N_12670,N_12492);
or U13515 (N_13515,N_12000,N_12853);
nor U13516 (N_13516,N_12746,N_12810);
xor U13517 (N_13517,N_12275,N_12793);
nor U13518 (N_13518,N_12847,N_12543);
xnor U13519 (N_13519,N_12879,N_12962);
and U13520 (N_13520,N_12060,N_12802);
nor U13521 (N_13521,N_12105,N_12366);
and U13522 (N_13522,N_12454,N_12024);
nand U13523 (N_13523,N_12859,N_12553);
xnor U13524 (N_13524,N_12806,N_12709);
xor U13525 (N_13525,N_12255,N_12647);
and U13526 (N_13526,N_12823,N_12757);
nor U13527 (N_13527,N_12430,N_12992);
and U13528 (N_13528,N_12713,N_12787);
xor U13529 (N_13529,N_12046,N_12428);
or U13530 (N_13530,N_12476,N_12328);
and U13531 (N_13531,N_12828,N_12555);
nor U13532 (N_13532,N_12908,N_12753);
xor U13533 (N_13533,N_12938,N_12476);
or U13534 (N_13534,N_12108,N_12680);
nand U13535 (N_13535,N_12084,N_12905);
nand U13536 (N_13536,N_12417,N_12194);
or U13537 (N_13537,N_12095,N_12480);
or U13538 (N_13538,N_12993,N_12002);
nor U13539 (N_13539,N_12770,N_12097);
nand U13540 (N_13540,N_12001,N_12460);
nand U13541 (N_13541,N_12033,N_12159);
and U13542 (N_13542,N_12848,N_12063);
nand U13543 (N_13543,N_12101,N_12062);
or U13544 (N_13544,N_12556,N_12501);
and U13545 (N_13545,N_12646,N_12817);
xnor U13546 (N_13546,N_12341,N_12852);
nor U13547 (N_13547,N_12705,N_12836);
or U13548 (N_13548,N_12749,N_12764);
xor U13549 (N_13549,N_12650,N_12778);
nand U13550 (N_13550,N_12584,N_12943);
or U13551 (N_13551,N_12189,N_12344);
nand U13552 (N_13552,N_12206,N_12176);
xnor U13553 (N_13553,N_12010,N_12692);
nor U13554 (N_13554,N_12616,N_12182);
xnor U13555 (N_13555,N_12519,N_12626);
and U13556 (N_13556,N_12381,N_12568);
xor U13557 (N_13557,N_12816,N_12183);
and U13558 (N_13558,N_12065,N_12896);
and U13559 (N_13559,N_12089,N_12399);
nand U13560 (N_13560,N_12047,N_12004);
and U13561 (N_13561,N_12195,N_12183);
xnor U13562 (N_13562,N_12948,N_12658);
nor U13563 (N_13563,N_12908,N_12257);
nor U13564 (N_13564,N_12698,N_12957);
or U13565 (N_13565,N_12601,N_12807);
nand U13566 (N_13566,N_12248,N_12153);
and U13567 (N_13567,N_12710,N_12754);
and U13568 (N_13568,N_12946,N_12512);
and U13569 (N_13569,N_12409,N_12621);
xnor U13570 (N_13570,N_12669,N_12819);
xor U13571 (N_13571,N_12523,N_12227);
nor U13572 (N_13572,N_12861,N_12096);
nand U13573 (N_13573,N_12247,N_12852);
and U13574 (N_13574,N_12231,N_12505);
xor U13575 (N_13575,N_12911,N_12733);
nor U13576 (N_13576,N_12407,N_12162);
and U13577 (N_13577,N_12099,N_12119);
xnor U13578 (N_13578,N_12852,N_12724);
nor U13579 (N_13579,N_12597,N_12837);
nand U13580 (N_13580,N_12586,N_12870);
xor U13581 (N_13581,N_12797,N_12501);
and U13582 (N_13582,N_12000,N_12346);
or U13583 (N_13583,N_12790,N_12013);
xnor U13584 (N_13584,N_12421,N_12306);
xnor U13585 (N_13585,N_12803,N_12704);
nor U13586 (N_13586,N_12847,N_12249);
nand U13587 (N_13587,N_12749,N_12614);
or U13588 (N_13588,N_12901,N_12300);
and U13589 (N_13589,N_12329,N_12103);
and U13590 (N_13590,N_12070,N_12281);
xor U13591 (N_13591,N_12425,N_12744);
nor U13592 (N_13592,N_12996,N_12219);
nor U13593 (N_13593,N_12422,N_12365);
nand U13594 (N_13594,N_12078,N_12095);
nand U13595 (N_13595,N_12108,N_12126);
nor U13596 (N_13596,N_12973,N_12702);
and U13597 (N_13597,N_12898,N_12419);
or U13598 (N_13598,N_12115,N_12599);
or U13599 (N_13599,N_12332,N_12539);
nand U13600 (N_13600,N_12199,N_12228);
and U13601 (N_13601,N_12436,N_12104);
nor U13602 (N_13602,N_12699,N_12955);
nor U13603 (N_13603,N_12845,N_12065);
xnor U13604 (N_13604,N_12721,N_12379);
nand U13605 (N_13605,N_12808,N_12918);
nand U13606 (N_13606,N_12515,N_12194);
or U13607 (N_13607,N_12392,N_12248);
xnor U13608 (N_13608,N_12444,N_12706);
and U13609 (N_13609,N_12107,N_12517);
nand U13610 (N_13610,N_12744,N_12029);
nor U13611 (N_13611,N_12108,N_12356);
nand U13612 (N_13612,N_12539,N_12372);
nor U13613 (N_13613,N_12482,N_12396);
xnor U13614 (N_13614,N_12779,N_12440);
or U13615 (N_13615,N_12082,N_12268);
or U13616 (N_13616,N_12154,N_12554);
nor U13617 (N_13617,N_12908,N_12361);
nor U13618 (N_13618,N_12666,N_12777);
nand U13619 (N_13619,N_12492,N_12678);
or U13620 (N_13620,N_12348,N_12801);
nand U13621 (N_13621,N_12804,N_12520);
or U13622 (N_13622,N_12048,N_12770);
and U13623 (N_13623,N_12365,N_12190);
and U13624 (N_13624,N_12495,N_12836);
nor U13625 (N_13625,N_12153,N_12074);
xor U13626 (N_13626,N_12692,N_12993);
xnor U13627 (N_13627,N_12384,N_12909);
or U13628 (N_13628,N_12548,N_12927);
and U13629 (N_13629,N_12445,N_12209);
or U13630 (N_13630,N_12962,N_12087);
and U13631 (N_13631,N_12237,N_12929);
nor U13632 (N_13632,N_12349,N_12646);
nand U13633 (N_13633,N_12706,N_12662);
nand U13634 (N_13634,N_12110,N_12483);
or U13635 (N_13635,N_12849,N_12455);
and U13636 (N_13636,N_12850,N_12669);
and U13637 (N_13637,N_12535,N_12332);
nor U13638 (N_13638,N_12648,N_12201);
and U13639 (N_13639,N_12801,N_12601);
or U13640 (N_13640,N_12881,N_12357);
and U13641 (N_13641,N_12620,N_12962);
nor U13642 (N_13642,N_12133,N_12344);
nor U13643 (N_13643,N_12038,N_12011);
nor U13644 (N_13644,N_12832,N_12804);
nor U13645 (N_13645,N_12330,N_12518);
xor U13646 (N_13646,N_12077,N_12791);
nor U13647 (N_13647,N_12981,N_12201);
xnor U13648 (N_13648,N_12085,N_12335);
and U13649 (N_13649,N_12152,N_12893);
xor U13650 (N_13650,N_12194,N_12939);
or U13651 (N_13651,N_12867,N_12868);
and U13652 (N_13652,N_12675,N_12871);
nor U13653 (N_13653,N_12148,N_12701);
xnor U13654 (N_13654,N_12584,N_12154);
or U13655 (N_13655,N_12548,N_12270);
nand U13656 (N_13656,N_12462,N_12327);
nor U13657 (N_13657,N_12839,N_12045);
xor U13658 (N_13658,N_12431,N_12566);
nor U13659 (N_13659,N_12928,N_12000);
nor U13660 (N_13660,N_12078,N_12829);
xnor U13661 (N_13661,N_12946,N_12185);
xnor U13662 (N_13662,N_12292,N_12586);
nand U13663 (N_13663,N_12232,N_12174);
or U13664 (N_13664,N_12250,N_12297);
nor U13665 (N_13665,N_12259,N_12352);
nand U13666 (N_13666,N_12089,N_12527);
nor U13667 (N_13667,N_12843,N_12870);
xor U13668 (N_13668,N_12749,N_12428);
or U13669 (N_13669,N_12339,N_12604);
and U13670 (N_13670,N_12575,N_12639);
xnor U13671 (N_13671,N_12475,N_12092);
or U13672 (N_13672,N_12455,N_12049);
or U13673 (N_13673,N_12684,N_12178);
or U13674 (N_13674,N_12357,N_12565);
and U13675 (N_13675,N_12580,N_12751);
nand U13676 (N_13676,N_12882,N_12071);
or U13677 (N_13677,N_12868,N_12749);
xor U13678 (N_13678,N_12125,N_12708);
xnor U13679 (N_13679,N_12854,N_12223);
xnor U13680 (N_13680,N_12815,N_12173);
xor U13681 (N_13681,N_12049,N_12423);
or U13682 (N_13682,N_12745,N_12041);
and U13683 (N_13683,N_12742,N_12974);
nand U13684 (N_13684,N_12380,N_12164);
nand U13685 (N_13685,N_12485,N_12016);
xnor U13686 (N_13686,N_12936,N_12430);
xor U13687 (N_13687,N_12818,N_12108);
or U13688 (N_13688,N_12904,N_12813);
or U13689 (N_13689,N_12555,N_12844);
or U13690 (N_13690,N_12967,N_12363);
nand U13691 (N_13691,N_12353,N_12482);
xnor U13692 (N_13692,N_12351,N_12344);
nor U13693 (N_13693,N_12693,N_12814);
nor U13694 (N_13694,N_12735,N_12877);
xor U13695 (N_13695,N_12628,N_12878);
nor U13696 (N_13696,N_12892,N_12692);
xnor U13697 (N_13697,N_12704,N_12940);
nand U13698 (N_13698,N_12610,N_12904);
nor U13699 (N_13699,N_12111,N_12295);
and U13700 (N_13700,N_12445,N_12321);
xnor U13701 (N_13701,N_12376,N_12373);
and U13702 (N_13702,N_12616,N_12374);
and U13703 (N_13703,N_12398,N_12511);
and U13704 (N_13704,N_12896,N_12403);
or U13705 (N_13705,N_12372,N_12634);
nor U13706 (N_13706,N_12881,N_12840);
nor U13707 (N_13707,N_12337,N_12283);
or U13708 (N_13708,N_12368,N_12491);
xnor U13709 (N_13709,N_12013,N_12083);
xor U13710 (N_13710,N_12407,N_12755);
xor U13711 (N_13711,N_12344,N_12987);
xor U13712 (N_13712,N_12617,N_12395);
xor U13713 (N_13713,N_12356,N_12793);
or U13714 (N_13714,N_12460,N_12234);
and U13715 (N_13715,N_12164,N_12226);
nor U13716 (N_13716,N_12840,N_12356);
nor U13717 (N_13717,N_12121,N_12172);
nand U13718 (N_13718,N_12606,N_12611);
and U13719 (N_13719,N_12513,N_12347);
xor U13720 (N_13720,N_12772,N_12729);
nor U13721 (N_13721,N_12248,N_12422);
or U13722 (N_13722,N_12698,N_12530);
xnor U13723 (N_13723,N_12355,N_12246);
nand U13724 (N_13724,N_12116,N_12682);
and U13725 (N_13725,N_12858,N_12160);
or U13726 (N_13726,N_12802,N_12077);
xnor U13727 (N_13727,N_12676,N_12345);
and U13728 (N_13728,N_12347,N_12397);
and U13729 (N_13729,N_12904,N_12861);
xnor U13730 (N_13730,N_12879,N_12185);
xnor U13731 (N_13731,N_12137,N_12057);
nand U13732 (N_13732,N_12787,N_12081);
and U13733 (N_13733,N_12271,N_12931);
xnor U13734 (N_13734,N_12659,N_12233);
xor U13735 (N_13735,N_12774,N_12073);
or U13736 (N_13736,N_12295,N_12734);
or U13737 (N_13737,N_12360,N_12477);
or U13738 (N_13738,N_12848,N_12229);
and U13739 (N_13739,N_12437,N_12498);
or U13740 (N_13740,N_12055,N_12153);
xnor U13741 (N_13741,N_12603,N_12966);
xor U13742 (N_13742,N_12843,N_12329);
and U13743 (N_13743,N_12630,N_12669);
xor U13744 (N_13744,N_12588,N_12058);
or U13745 (N_13745,N_12454,N_12131);
xor U13746 (N_13746,N_12530,N_12642);
nor U13747 (N_13747,N_12251,N_12633);
nor U13748 (N_13748,N_12041,N_12861);
nand U13749 (N_13749,N_12265,N_12597);
and U13750 (N_13750,N_12801,N_12201);
xnor U13751 (N_13751,N_12940,N_12847);
nor U13752 (N_13752,N_12211,N_12337);
xnor U13753 (N_13753,N_12595,N_12963);
or U13754 (N_13754,N_12192,N_12547);
or U13755 (N_13755,N_12195,N_12780);
nor U13756 (N_13756,N_12730,N_12715);
nand U13757 (N_13757,N_12956,N_12394);
and U13758 (N_13758,N_12288,N_12987);
or U13759 (N_13759,N_12840,N_12337);
nor U13760 (N_13760,N_12348,N_12257);
xor U13761 (N_13761,N_12884,N_12396);
nor U13762 (N_13762,N_12702,N_12202);
xnor U13763 (N_13763,N_12203,N_12982);
nor U13764 (N_13764,N_12835,N_12443);
or U13765 (N_13765,N_12356,N_12190);
nand U13766 (N_13766,N_12439,N_12844);
or U13767 (N_13767,N_12034,N_12994);
xnor U13768 (N_13768,N_12954,N_12515);
or U13769 (N_13769,N_12068,N_12314);
nor U13770 (N_13770,N_12804,N_12377);
nor U13771 (N_13771,N_12172,N_12195);
xor U13772 (N_13772,N_12399,N_12945);
and U13773 (N_13773,N_12076,N_12689);
nand U13774 (N_13774,N_12168,N_12541);
xnor U13775 (N_13775,N_12540,N_12506);
or U13776 (N_13776,N_12503,N_12289);
and U13777 (N_13777,N_12948,N_12502);
or U13778 (N_13778,N_12027,N_12073);
xor U13779 (N_13779,N_12745,N_12647);
nor U13780 (N_13780,N_12746,N_12495);
or U13781 (N_13781,N_12636,N_12313);
and U13782 (N_13782,N_12972,N_12040);
nand U13783 (N_13783,N_12721,N_12972);
nor U13784 (N_13784,N_12415,N_12851);
or U13785 (N_13785,N_12681,N_12062);
xnor U13786 (N_13786,N_12284,N_12522);
or U13787 (N_13787,N_12263,N_12982);
nand U13788 (N_13788,N_12371,N_12684);
nor U13789 (N_13789,N_12677,N_12636);
nand U13790 (N_13790,N_12306,N_12214);
nand U13791 (N_13791,N_12135,N_12050);
nor U13792 (N_13792,N_12370,N_12103);
or U13793 (N_13793,N_12703,N_12962);
nor U13794 (N_13794,N_12776,N_12209);
and U13795 (N_13795,N_12794,N_12635);
nand U13796 (N_13796,N_12912,N_12934);
nor U13797 (N_13797,N_12378,N_12209);
or U13798 (N_13798,N_12259,N_12131);
or U13799 (N_13799,N_12655,N_12697);
xor U13800 (N_13800,N_12065,N_12984);
and U13801 (N_13801,N_12523,N_12530);
or U13802 (N_13802,N_12945,N_12849);
xor U13803 (N_13803,N_12522,N_12365);
nand U13804 (N_13804,N_12238,N_12320);
nand U13805 (N_13805,N_12515,N_12729);
xnor U13806 (N_13806,N_12049,N_12066);
xor U13807 (N_13807,N_12253,N_12236);
nor U13808 (N_13808,N_12595,N_12407);
xor U13809 (N_13809,N_12666,N_12576);
xor U13810 (N_13810,N_12370,N_12572);
nor U13811 (N_13811,N_12762,N_12342);
or U13812 (N_13812,N_12932,N_12303);
xor U13813 (N_13813,N_12168,N_12293);
and U13814 (N_13814,N_12262,N_12356);
nor U13815 (N_13815,N_12587,N_12586);
nor U13816 (N_13816,N_12774,N_12228);
or U13817 (N_13817,N_12752,N_12030);
and U13818 (N_13818,N_12701,N_12494);
or U13819 (N_13819,N_12641,N_12100);
or U13820 (N_13820,N_12244,N_12336);
or U13821 (N_13821,N_12783,N_12419);
xor U13822 (N_13822,N_12307,N_12336);
or U13823 (N_13823,N_12759,N_12474);
nor U13824 (N_13824,N_12956,N_12774);
or U13825 (N_13825,N_12067,N_12606);
and U13826 (N_13826,N_12905,N_12229);
or U13827 (N_13827,N_12219,N_12047);
and U13828 (N_13828,N_12393,N_12240);
nor U13829 (N_13829,N_12281,N_12240);
nand U13830 (N_13830,N_12569,N_12609);
nor U13831 (N_13831,N_12697,N_12702);
and U13832 (N_13832,N_12465,N_12447);
nor U13833 (N_13833,N_12730,N_12249);
nand U13834 (N_13834,N_12048,N_12784);
nand U13835 (N_13835,N_12289,N_12658);
and U13836 (N_13836,N_12687,N_12044);
nand U13837 (N_13837,N_12599,N_12737);
or U13838 (N_13838,N_12971,N_12439);
xnor U13839 (N_13839,N_12671,N_12411);
and U13840 (N_13840,N_12755,N_12195);
and U13841 (N_13841,N_12291,N_12396);
nor U13842 (N_13842,N_12938,N_12470);
xor U13843 (N_13843,N_12247,N_12909);
nor U13844 (N_13844,N_12060,N_12285);
xnor U13845 (N_13845,N_12959,N_12664);
xor U13846 (N_13846,N_12261,N_12795);
nor U13847 (N_13847,N_12567,N_12089);
xnor U13848 (N_13848,N_12627,N_12485);
nor U13849 (N_13849,N_12633,N_12300);
nor U13850 (N_13850,N_12192,N_12089);
and U13851 (N_13851,N_12542,N_12734);
and U13852 (N_13852,N_12276,N_12937);
xor U13853 (N_13853,N_12858,N_12236);
xor U13854 (N_13854,N_12246,N_12106);
or U13855 (N_13855,N_12263,N_12520);
nand U13856 (N_13856,N_12330,N_12183);
nor U13857 (N_13857,N_12018,N_12897);
and U13858 (N_13858,N_12963,N_12192);
or U13859 (N_13859,N_12297,N_12091);
or U13860 (N_13860,N_12877,N_12573);
or U13861 (N_13861,N_12455,N_12522);
nand U13862 (N_13862,N_12438,N_12228);
nand U13863 (N_13863,N_12489,N_12003);
nor U13864 (N_13864,N_12901,N_12290);
xnor U13865 (N_13865,N_12333,N_12377);
or U13866 (N_13866,N_12268,N_12262);
nand U13867 (N_13867,N_12063,N_12058);
nor U13868 (N_13868,N_12695,N_12032);
nor U13869 (N_13869,N_12459,N_12183);
xnor U13870 (N_13870,N_12181,N_12008);
nand U13871 (N_13871,N_12278,N_12723);
and U13872 (N_13872,N_12830,N_12227);
or U13873 (N_13873,N_12698,N_12796);
or U13874 (N_13874,N_12792,N_12701);
nand U13875 (N_13875,N_12842,N_12295);
xnor U13876 (N_13876,N_12300,N_12367);
or U13877 (N_13877,N_12716,N_12997);
and U13878 (N_13878,N_12873,N_12725);
or U13879 (N_13879,N_12455,N_12859);
and U13880 (N_13880,N_12344,N_12428);
or U13881 (N_13881,N_12737,N_12237);
nand U13882 (N_13882,N_12361,N_12061);
or U13883 (N_13883,N_12676,N_12187);
xor U13884 (N_13884,N_12851,N_12256);
nand U13885 (N_13885,N_12465,N_12748);
nor U13886 (N_13886,N_12237,N_12478);
or U13887 (N_13887,N_12005,N_12693);
or U13888 (N_13888,N_12689,N_12860);
nor U13889 (N_13889,N_12811,N_12334);
and U13890 (N_13890,N_12434,N_12218);
or U13891 (N_13891,N_12916,N_12021);
or U13892 (N_13892,N_12077,N_12422);
and U13893 (N_13893,N_12156,N_12285);
nand U13894 (N_13894,N_12777,N_12523);
nor U13895 (N_13895,N_12145,N_12177);
or U13896 (N_13896,N_12987,N_12508);
and U13897 (N_13897,N_12500,N_12651);
or U13898 (N_13898,N_12755,N_12490);
xor U13899 (N_13899,N_12684,N_12516);
nor U13900 (N_13900,N_12124,N_12508);
xor U13901 (N_13901,N_12301,N_12683);
nor U13902 (N_13902,N_12813,N_12831);
and U13903 (N_13903,N_12667,N_12261);
and U13904 (N_13904,N_12216,N_12186);
and U13905 (N_13905,N_12811,N_12852);
xor U13906 (N_13906,N_12883,N_12063);
xnor U13907 (N_13907,N_12174,N_12412);
and U13908 (N_13908,N_12874,N_12508);
nand U13909 (N_13909,N_12745,N_12614);
or U13910 (N_13910,N_12783,N_12679);
nand U13911 (N_13911,N_12514,N_12988);
or U13912 (N_13912,N_12879,N_12587);
nand U13913 (N_13913,N_12815,N_12228);
xnor U13914 (N_13914,N_12146,N_12366);
or U13915 (N_13915,N_12953,N_12176);
nand U13916 (N_13916,N_12067,N_12676);
or U13917 (N_13917,N_12850,N_12189);
nand U13918 (N_13918,N_12417,N_12631);
nor U13919 (N_13919,N_12492,N_12683);
nor U13920 (N_13920,N_12788,N_12630);
nand U13921 (N_13921,N_12255,N_12151);
xor U13922 (N_13922,N_12541,N_12045);
or U13923 (N_13923,N_12132,N_12913);
and U13924 (N_13924,N_12418,N_12360);
nor U13925 (N_13925,N_12913,N_12523);
nor U13926 (N_13926,N_12469,N_12266);
nor U13927 (N_13927,N_12768,N_12376);
or U13928 (N_13928,N_12332,N_12360);
nor U13929 (N_13929,N_12352,N_12859);
xnor U13930 (N_13930,N_12107,N_12944);
and U13931 (N_13931,N_12016,N_12574);
nand U13932 (N_13932,N_12374,N_12517);
or U13933 (N_13933,N_12938,N_12620);
xnor U13934 (N_13934,N_12958,N_12389);
or U13935 (N_13935,N_12540,N_12784);
and U13936 (N_13936,N_12877,N_12594);
nand U13937 (N_13937,N_12139,N_12450);
xnor U13938 (N_13938,N_12010,N_12694);
or U13939 (N_13939,N_12494,N_12091);
and U13940 (N_13940,N_12268,N_12488);
or U13941 (N_13941,N_12718,N_12693);
and U13942 (N_13942,N_12539,N_12163);
or U13943 (N_13943,N_12312,N_12193);
or U13944 (N_13944,N_12453,N_12315);
xor U13945 (N_13945,N_12063,N_12263);
nand U13946 (N_13946,N_12790,N_12323);
xor U13947 (N_13947,N_12264,N_12289);
xor U13948 (N_13948,N_12929,N_12028);
nand U13949 (N_13949,N_12667,N_12447);
nand U13950 (N_13950,N_12757,N_12570);
xnor U13951 (N_13951,N_12456,N_12742);
xnor U13952 (N_13952,N_12396,N_12013);
and U13953 (N_13953,N_12106,N_12682);
nand U13954 (N_13954,N_12256,N_12340);
nand U13955 (N_13955,N_12346,N_12873);
nand U13956 (N_13956,N_12644,N_12112);
xor U13957 (N_13957,N_12624,N_12915);
nor U13958 (N_13958,N_12021,N_12301);
xor U13959 (N_13959,N_12251,N_12442);
nand U13960 (N_13960,N_12499,N_12182);
and U13961 (N_13961,N_12722,N_12543);
or U13962 (N_13962,N_12260,N_12441);
and U13963 (N_13963,N_12649,N_12056);
and U13964 (N_13964,N_12459,N_12102);
or U13965 (N_13965,N_12489,N_12136);
nand U13966 (N_13966,N_12993,N_12201);
xnor U13967 (N_13967,N_12274,N_12515);
xnor U13968 (N_13968,N_12112,N_12146);
and U13969 (N_13969,N_12901,N_12931);
and U13970 (N_13970,N_12010,N_12059);
nor U13971 (N_13971,N_12819,N_12682);
xor U13972 (N_13972,N_12334,N_12141);
nor U13973 (N_13973,N_12269,N_12137);
and U13974 (N_13974,N_12211,N_12341);
nor U13975 (N_13975,N_12084,N_12083);
nor U13976 (N_13976,N_12244,N_12129);
nand U13977 (N_13977,N_12056,N_12569);
nand U13978 (N_13978,N_12654,N_12190);
or U13979 (N_13979,N_12940,N_12627);
or U13980 (N_13980,N_12727,N_12572);
or U13981 (N_13981,N_12909,N_12638);
xor U13982 (N_13982,N_12418,N_12485);
xnor U13983 (N_13983,N_12763,N_12418);
xnor U13984 (N_13984,N_12954,N_12522);
and U13985 (N_13985,N_12795,N_12550);
and U13986 (N_13986,N_12338,N_12542);
xor U13987 (N_13987,N_12998,N_12551);
nand U13988 (N_13988,N_12790,N_12627);
xnor U13989 (N_13989,N_12835,N_12957);
nor U13990 (N_13990,N_12350,N_12442);
or U13991 (N_13991,N_12845,N_12887);
nor U13992 (N_13992,N_12184,N_12327);
or U13993 (N_13993,N_12943,N_12576);
or U13994 (N_13994,N_12911,N_12840);
or U13995 (N_13995,N_12659,N_12750);
xor U13996 (N_13996,N_12982,N_12423);
or U13997 (N_13997,N_12401,N_12706);
or U13998 (N_13998,N_12457,N_12181);
nand U13999 (N_13999,N_12867,N_12222);
xor U14000 (N_14000,N_13581,N_13056);
or U14001 (N_14001,N_13548,N_13628);
nand U14002 (N_14002,N_13843,N_13546);
xor U14003 (N_14003,N_13924,N_13239);
and U14004 (N_14004,N_13313,N_13600);
or U14005 (N_14005,N_13820,N_13137);
or U14006 (N_14006,N_13980,N_13587);
or U14007 (N_14007,N_13810,N_13723);
or U14008 (N_14008,N_13374,N_13627);
xnor U14009 (N_14009,N_13123,N_13113);
xnor U14010 (N_14010,N_13541,N_13172);
nand U14011 (N_14011,N_13630,N_13444);
xor U14012 (N_14012,N_13453,N_13883);
and U14013 (N_14013,N_13108,N_13086);
nor U14014 (N_14014,N_13064,N_13827);
and U14015 (N_14015,N_13614,N_13162);
nand U14016 (N_14016,N_13101,N_13046);
nand U14017 (N_14017,N_13584,N_13325);
or U14018 (N_14018,N_13375,N_13503);
or U14019 (N_14019,N_13177,N_13315);
nand U14020 (N_14020,N_13700,N_13021);
and U14021 (N_14021,N_13276,N_13815);
xor U14022 (N_14022,N_13864,N_13801);
nand U14023 (N_14023,N_13765,N_13710);
nor U14024 (N_14024,N_13590,N_13649);
nand U14025 (N_14025,N_13194,N_13040);
or U14026 (N_14026,N_13533,N_13154);
and U14027 (N_14027,N_13084,N_13519);
and U14028 (N_14028,N_13944,N_13898);
nand U14029 (N_14029,N_13271,N_13348);
xnor U14030 (N_14030,N_13957,N_13770);
or U14031 (N_14031,N_13520,N_13821);
and U14032 (N_14032,N_13126,N_13211);
nor U14033 (N_14033,N_13911,N_13975);
nand U14034 (N_14034,N_13814,N_13925);
nand U14035 (N_14035,N_13009,N_13940);
nor U14036 (N_14036,N_13717,N_13709);
xor U14037 (N_14037,N_13999,N_13228);
or U14038 (N_14038,N_13718,N_13391);
or U14039 (N_14039,N_13722,N_13007);
or U14040 (N_14040,N_13256,N_13532);
and U14041 (N_14041,N_13462,N_13085);
xor U14042 (N_14042,N_13932,N_13159);
nand U14043 (N_14043,N_13759,N_13849);
and U14044 (N_14044,N_13903,N_13212);
nor U14045 (N_14045,N_13218,N_13362);
and U14046 (N_14046,N_13730,N_13262);
or U14047 (N_14047,N_13433,N_13384);
nor U14048 (N_14048,N_13324,N_13420);
and U14049 (N_14049,N_13869,N_13110);
nor U14050 (N_14050,N_13750,N_13835);
or U14051 (N_14051,N_13876,N_13415);
nor U14052 (N_14052,N_13209,N_13141);
xor U14053 (N_14053,N_13233,N_13363);
xor U14054 (N_14054,N_13557,N_13594);
nand U14055 (N_14055,N_13592,N_13024);
nor U14056 (N_14056,N_13173,N_13307);
nor U14057 (N_14057,N_13298,N_13715);
nand U14058 (N_14058,N_13776,N_13634);
nor U14059 (N_14059,N_13997,N_13254);
nor U14060 (N_14060,N_13422,N_13398);
or U14061 (N_14061,N_13777,N_13358);
nand U14062 (N_14062,N_13045,N_13439);
nand U14063 (N_14063,N_13906,N_13329);
xnor U14064 (N_14064,N_13031,N_13409);
nand U14065 (N_14065,N_13939,N_13185);
nor U14066 (N_14066,N_13583,N_13392);
and U14067 (N_14067,N_13961,N_13977);
nand U14068 (N_14068,N_13204,N_13521);
nand U14069 (N_14069,N_13000,N_13248);
xor U14070 (N_14070,N_13234,N_13602);
nor U14071 (N_14071,N_13861,N_13522);
and U14072 (N_14072,N_13757,N_13564);
or U14073 (N_14073,N_13314,N_13673);
and U14074 (N_14074,N_13549,N_13896);
xnor U14075 (N_14075,N_13741,N_13011);
and U14076 (N_14076,N_13933,N_13247);
nand U14077 (N_14077,N_13454,N_13958);
xnor U14078 (N_14078,N_13342,N_13487);
nor U14079 (N_14079,N_13726,N_13902);
or U14080 (N_14080,N_13037,N_13518);
and U14081 (N_14081,N_13962,N_13819);
nor U14082 (N_14082,N_13465,N_13260);
nor U14083 (N_14083,N_13451,N_13643);
xnor U14084 (N_14084,N_13704,N_13073);
xnor U14085 (N_14085,N_13699,N_13484);
or U14086 (N_14086,N_13778,N_13702);
xnor U14087 (N_14087,N_13766,N_13216);
nand U14088 (N_14088,N_13095,N_13339);
nor U14089 (N_14089,N_13432,N_13582);
or U14090 (N_14090,N_13251,N_13580);
or U14091 (N_14091,N_13772,N_13201);
or U14092 (N_14092,N_13192,N_13371);
xnor U14093 (N_14093,N_13812,N_13620);
nor U14094 (N_14094,N_13554,N_13938);
nor U14095 (N_14095,N_13461,N_13565);
and U14096 (N_14096,N_13823,N_13662);
nand U14097 (N_14097,N_13394,N_13966);
nor U14098 (N_14098,N_13603,N_13979);
nand U14099 (N_14099,N_13929,N_13756);
and U14100 (N_14100,N_13403,N_13197);
nor U14101 (N_14101,N_13107,N_13641);
nand U14102 (N_14102,N_13800,N_13555);
nand U14103 (N_14103,N_13285,N_13663);
or U14104 (N_14104,N_13142,N_13449);
and U14105 (N_14105,N_13585,N_13118);
nand U14106 (N_14106,N_13379,N_13891);
and U14107 (N_14107,N_13186,N_13199);
and U14108 (N_14108,N_13690,N_13091);
nand U14109 (N_14109,N_13479,N_13556);
nand U14110 (N_14110,N_13301,N_13727);
nand U14111 (N_14111,N_13593,N_13292);
nand U14112 (N_14112,N_13624,N_13317);
and U14113 (N_14113,N_13544,N_13402);
nor U14114 (N_14114,N_13005,N_13751);
nand U14115 (N_14115,N_13240,N_13296);
and U14116 (N_14116,N_13951,N_13346);
or U14117 (N_14117,N_13908,N_13825);
nor U14118 (N_14118,N_13245,N_13724);
and U14119 (N_14119,N_13882,N_13886);
nand U14120 (N_14120,N_13563,N_13026);
nor U14121 (N_14121,N_13542,N_13488);
nor U14122 (N_14122,N_13236,N_13865);
or U14123 (N_14123,N_13716,N_13436);
and U14124 (N_14124,N_13050,N_13680);
nand U14125 (N_14125,N_13794,N_13918);
and U14126 (N_14126,N_13619,N_13033);
xnor U14127 (N_14127,N_13832,N_13761);
nor U14128 (N_14128,N_13134,N_13809);
nor U14129 (N_14129,N_13611,N_13983);
nand U14130 (N_14130,N_13745,N_13993);
or U14131 (N_14131,N_13639,N_13573);
and U14132 (N_14132,N_13399,N_13203);
nand U14133 (N_14133,N_13854,N_13839);
and U14134 (N_14134,N_13121,N_13534);
or U14135 (N_14135,N_13472,N_13791);
xnor U14136 (N_14136,N_13691,N_13104);
nand U14137 (N_14137,N_13106,N_13874);
or U14138 (N_14138,N_13482,N_13987);
nor U14139 (N_14139,N_13613,N_13257);
nor U14140 (N_14140,N_13102,N_13842);
or U14141 (N_14141,N_13622,N_13176);
nor U14142 (N_14142,N_13266,N_13885);
nor U14143 (N_14143,N_13020,N_13509);
and U14144 (N_14144,N_13366,N_13596);
xor U14145 (N_14145,N_13469,N_13848);
and U14146 (N_14146,N_13122,N_13658);
and U14147 (N_14147,N_13261,N_13151);
nand U14148 (N_14148,N_13226,N_13599);
nor U14149 (N_14149,N_13408,N_13686);
nand U14150 (N_14150,N_13166,N_13308);
or U14151 (N_14151,N_13115,N_13650);
xor U14152 (N_14152,N_13517,N_13023);
xor U14153 (N_14153,N_13536,N_13438);
or U14154 (N_14154,N_13274,N_13179);
nand U14155 (N_14155,N_13167,N_13735);
nand U14156 (N_14156,N_13258,N_13213);
or U14157 (N_14157,N_13719,N_13783);
nor U14158 (N_14158,N_13205,N_13077);
nand U14159 (N_14159,N_13497,N_13025);
and U14160 (N_14160,N_13284,N_13075);
or U14161 (N_14161,N_13644,N_13286);
nand U14162 (N_14162,N_13250,N_13341);
and U14163 (N_14163,N_13889,N_13065);
or U14164 (N_14164,N_13019,N_13076);
nand U14165 (N_14165,N_13180,N_13605);
or U14166 (N_14166,N_13930,N_13830);
xnor U14167 (N_14167,N_13922,N_13935);
and U14168 (N_14168,N_13041,N_13516);
xor U14169 (N_14169,N_13335,N_13551);
and U14170 (N_14170,N_13665,N_13305);
nor U14171 (N_14171,N_13505,N_13540);
and U14172 (N_14172,N_13858,N_13004);
or U14173 (N_14173,N_13066,N_13867);
nand U14174 (N_14174,N_13357,N_13460);
nor U14175 (N_14175,N_13851,N_13749);
and U14176 (N_14176,N_13871,N_13214);
or U14177 (N_14177,N_13664,N_13053);
xor U14178 (N_14178,N_13318,N_13788);
nand U14179 (N_14179,N_13155,N_13395);
nand U14180 (N_14180,N_13822,N_13733);
xor U14181 (N_14181,N_13049,N_13913);
nor U14182 (N_14182,N_13178,N_13941);
nand U14183 (N_14183,N_13208,N_13368);
nor U14184 (N_14184,N_13547,N_13720);
nor U14185 (N_14185,N_13734,N_13758);
nand U14186 (N_14186,N_13143,N_13901);
nand U14187 (N_14187,N_13838,N_13976);
xor U14188 (N_14188,N_13014,N_13070);
nor U14189 (N_14189,N_13967,N_13900);
xnor U14190 (N_14190,N_13390,N_13708);
nand U14191 (N_14191,N_13824,N_13012);
and U14192 (N_14192,N_13942,N_13195);
xnor U14193 (N_14193,N_13857,N_13743);
and U14194 (N_14194,N_13184,N_13606);
nor U14195 (N_14195,N_13738,N_13418);
xnor U14196 (N_14196,N_13237,N_13294);
and U14197 (N_14197,N_13361,N_13968);
or U14198 (N_14198,N_13131,N_13464);
nor U14199 (N_14199,N_13381,N_13198);
or U14200 (N_14200,N_13696,N_13456);
nor U14201 (N_14201,N_13471,N_13895);
nor U14202 (N_14202,N_13931,N_13295);
or U14203 (N_14203,N_13607,N_13183);
nor U14204 (N_14204,N_13333,N_13369);
nor U14205 (N_14205,N_13279,N_13642);
nand U14206 (N_14206,N_13986,N_13003);
or U14207 (N_14207,N_13786,N_13133);
or U14208 (N_14208,N_13921,N_13561);
and U14209 (N_14209,N_13376,N_13356);
nor U14210 (N_14210,N_13175,N_13515);
or U14211 (N_14211,N_13648,N_13388);
nor U14212 (N_14212,N_13656,N_13351);
nor U14213 (N_14213,N_13631,N_13744);
or U14214 (N_14214,N_13588,N_13928);
nor U14215 (N_14215,N_13904,N_13287);
or U14216 (N_14216,N_13330,N_13117);
or U14217 (N_14217,N_13569,N_13425);
and U14218 (N_14218,N_13069,N_13319);
or U14219 (N_14219,N_13907,N_13470);
nand U14220 (N_14220,N_13872,N_13586);
and U14221 (N_14221,N_13998,N_13316);
nand U14222 (N_14222,N_13164,N_13281);
xor U14223 (N_14223,N_13343,N_13253);
or U14224 (N_14224,N_13112,N_13496);
xnor U14225 (N_14225,N_13481,N_13171);
nor U14226 (N_14226,N_13909,N_13452);
and U14227 (N_14227,N_13217,N_13808);
and U14228 (N_14228,N_13514,N_13467);
xor U14229 (N_14229,N_13063,N_13174);
xor U14230 (N_14230,N_13447,N_13372);
nor U14231 (N_14231,N_13651,N_13135);
nand U14232 (N_14232,N_13675,N_13666);
nand U14233 (N_14233,N_13670,N_13168);
or U14234 (N_14234,N_13074,N_13767);
and U14235 (N_14235,N_13996,N_13032);
and U14236 (N_14236,N_13833,N_13491);
or U14237 (N_14237,N_13311,N_13132);
xor U14238 (N_14238,N_13780,N_13919);
or U14239 (N_14239,N_13952,N_13992);
or U14240 (N_14240,N_13990,N_13147);
or U14241 (N_14241,N_13016,N_13897);
xnor U14242 (N_14242,N_13309,N_13015);
nand U14243 (N_14243,N_13235,N_13169);
nand U14244 (N_14244,N_13047,N_13430);
or U14245 (N_14245,N_13672,N_13082);
or U14246 (N_14246,N_13625,N_13637);
or U14247 (N_14247,N_13712,N_13834);
nand U14248 (N_14248,N_13303,N_13249);
nand U14249 (N_14249,N_13633,N_13576);
or U14250 (N_14250,N_13412,N_13753);
or U14251 (N_14251,N_13655,N_13423);
nor U14252 (N_14252,N_13746,N_13732);
nor U14253 (N_14253,N_13579,N_13378);
or U14254 (N_14254,N_13873,N_13448);
nand U14255 (N_14255,N_13721,N_13994);
nand U14256 (N_14256,N_13511,N_13893);
nor U14257 (N_14257,N_13689,N_13530);
and U14258 (N_14258,N_13034,N_13693);
xor U14259 (N_14259,N_13779,N_13936);
or U14260 (N_14260,N_13042,N_13193);
nand U14261 (N_14261,N_13528,N_13754);
nand U14262 (N_14262,N_13773,N_13948);
xor U14263 (N_14263,N_13653,N_13784);
or U14264 (N_14264,N_13685,N_13232);
nor U14265 (N_14265,N_13729,N_13125);
or U14266 (N_14266,N_13382,N_13140);
or U14267 (N_14267,N_13310,N_13377);
and U14268 (N_14268,N_13828,N_13798);
xor U14269 (N_14269,N_13181,N_13450);
or U14270 (N_14270,N_13538,N_13934);
nor U14271 (N_14271,N_13806,N_13280);
nand U14272 (N_14272,N_13960,N_13275);
nand U14273 (N_14273,N_13574,N_13100);
and U14274 (N_14274,N_13081,N_13492);
nor U14275 (N_14275,N_13289,N_13411);
or U14276 (N_14276,N_13269,N_13618);
xnor U14277 (N_14277,N_13706,N_13238);
nand U14278 (N_14278,N_13446,N_13923);
or U14279 (N_14279,N_13553,N_13668);
and U14280 (N_14280,N_13971,N_13406);
or U14281 (N_14281,N_13762,N_13424);
nand U14282 (N_14282,N_13048,N_13974);
or U14283 (N_14283,N_13455,N_13972);
nand U14284 (N_14284,N_13850,N_13252);
nand U14285 (N_14285,N_13494,N_13389);
nand U14286 (N_14286,N_13457,N_13621);
nand U14287 (N_14287,N_13768,N_13959);
xor U14288 (N_14288,N_13344,N_13230);
nand U14289 (N_14289,N_13984,N_13413);
or U14290 (N_14290,N_13635,N_13079);
xor U14291 (N_14291,N_13558,N_13352);
and U14292 (N_14292,N_13202,N_13512);
xor U14293 (N_14293,N_13359,N_13035);
nor U14294 (N_14294,N_13092,N_13499);
xor U14295 (N_14295,N_13905,N_13504);
xnor U14296 (N_14296,N_13157,N_13419);
and U14297 (N_14297,N_13323,N_13291);
xor U14298 (N_14298,N_13793,N_13054);
and U14299 (N_14299,N_13831,N_13725);
xor U14300 (N_14300,N_13697,N_13350);
and U14301 (N_14301,N_13604,N_13340);
nand U14302 (N_14302,N_13953,N_13892);
nand U14303 (N_14303,N_13401,N_13659);
nand U14304 (N_14304,N_13881,N_13227);
xnor U14305 (N_14305,N_13062,N_13529);
or U14306 (N_14306,N_13705,N_13364);
xnor U14307 (N_14307,N_13888,N_13608);
xor U14308 (N_14308,N_13242,N_13473);
or U14309 (N_14309,N_13191,N_13052);
xnor U14310 (N_14310,N_13807,N_13890);
and U14311 (N_14311,N_13416,N_13950);
nor U14312 (N_14312,N_13853,N_13410);
or U14313 (N_14313,N_13739,N_13139);
xnor U14314 (N_14314,N_13914,N_13552);
and U14315 (N_14315,N_13638,N_13083);
xor U14316 (N_14316,N_13636,N_13617);
xnor U14317 (N_14317,N_13243,N_13225);
nor U14318 (N_14318,N_13103,N_13674);
nor U14319 (N_14319,N_13769,N_13785);
xnor U14320 (N_14320,N_13545,N_13485);
or U14321 (N_14321,N_13844,N_13337);
and U14322 (N_14322,N_13626,N_13327);
nand U14323 (N_14323,N_13578,N_13567);
nor U14324 (N_14324,N_13837,N_13127);
nand U14325 (N_14325,N_13099,N_13714);
and U14326 (N_14326,N_13144,N_13523);
nor U14327 (N_14327,N_13796,N_13027);
xor U14328 (N_14328,N_13428,N_13787);
nor U14329 (N_14329,N_13632,N_13029);
nor U14330 (N_14330,N_13441,N_13331);
nand U14331 (N_14331,N_13852,N_13591);
and U14332 (N_14332,N_13043,N_13894);
and U14333 (N_14333,N_13474,N_13840);
or U14334 (N_14334,N_13707,N_13096);
nor U14335 (N_14335,N_13222,N_13055);
nor U14336 (N_14336,N_13506,N_13160);
xor U14337 (N_14337,N_13263,N_13334);
xor U14338 (N_14338,N_13550,N_13661);
nand U14339 (N_14339,N_13332,N_13845);
or U14340 (N_14340,N_13434,N_13568);
nand U14341 (N_14341,N_13797,N_13476);
and U14342 (N_14342,N_13669,N_13763);
and U14343 (N_14343,N_13060,N_13915);
nor U14344 (N_14344,N_13038,N_13061);
or U14345 (N_14345,N_13970,N_13559);
xnor U14346 (N_14346,N_13677,N_13513);
or U14347 (N_14347,N_13483,N_13443);
or U14348 (N_14348,N_13124,N_13165);
or U14349 (N_14349,N_13946,N_13152);
or U14350 (N_14350,N_13955,N_13775);
nand U14351 (N_14351,N_13836,N_13989);
or U14352 (N_14352,N_13737,N_13829);
nand U14353 (N_14353,N_13109,N_13302);
nand U14354 (N_14354,N_13846,N_13463);
and U14355 (N_14355,N_13044,N_13790);
nand U14356 (N_14356,N_13866,N_13995);
xor U14357 (N_14357,N_13304,N_13681);
xor U14358 (N_14358,N_13200,N_13071);
and U14359 (N_14359,N_13093,N_13490);
xnor U14360 (N_14360,N_13030,N_13145);
nand U14361 (N_14361,N_13880,N_13577);
or U14362 (N_14362,N_13264,N_13560);
nor U14363 (N_14363,N_13426,N_13421);
or U14364 (N_14364,N_13347,N_13068);
or U14365 (N_14365,N_13489,N_13445);
and U14366 (N_14366,N_13130,N_13698);
nor U14367 (N_14367,N_13945,N_13396);
xor U14368 (N_14368,N_13789,N_13713);
nor U14369 (N_14369,N_13480,N_13982);
or U14370 (N_14370,N_13207,N_13969);
nor U14371 (N_14371,N_13146,N_13010);
nand U14372 (N_14372,N_13244,N_13562);
and U14373 (N_14373,N_13535,N_13414);
nand U14374 (N_14374,N_13017,N_13189);
and U14375 (N_14375,N_13774,N_13616);
xor U14376 (N_14376,N_13170,N_13646);
or U14377 (N_14377,N_13855,N_13507);
nor U14378 (N_14378,N_13912,N_13153);
xor U14379 (N_14379,N_13190,N_13863);
or U14380 (N_14380,N_13059,N_13028);
and U14381 (N_14381,N_13684,N_13956);
or U14382 (N_14382,N_13826,N_13373);
or U14383 (N_14383,N_13657,N_13387);
nor U14384 (N_14384,N_13740,N_13654);
and U14385 (N_14385,N_13259,N_13802);
and U14386 (N_14386,N_13206,N_13543);
or U14387 (N_14387,N_13385,N_13268);
nor U14388 (N_14388,N_13129,N_13752);
xor U14389 (N_14389,N_13601,N_13078);
nor U14390 (N_14390,N_13405,N_13210);
xor U14391 (N_14391,N_13682,N_13196);
or U14392 (N_14392,N_13229,N_13355);
xor U14393 (N_14393,N_13293,N_13612);
or U14394 (N_14394,N_13524,N_13215);
and U14395 (N_14395,N_13300,N_13008);
nor U14396 (N_14396,N_13879,N_13088);
xor U14397 (N_14397,N_13917,N_13610);
nor U14398 (N_14398,N_13531,N_13417);
nand U14399 (N_14399,N_13188,N_13321);
and U14400 (N_14400,N_13435,N_13246);
xnor U14401 (N_14401,N_13477,N_13964);
and U14402 (N_14402,N_13652,N_13006);
or U14403 (N_14403,N_13671,N_13380);
and U14404 (N_14404,N_13629,N_13051);
nand U14405 (N_14405,N_13817,N_13943);
xor U14406 (N_14406,N_13527,N_13120);
and U14407 (N_14407,N_13711,N_13597);
nor U14408 (N_14408,N_13098,N_13887);
or U14409 (N_14409,N_13978,N_13731);
nand U14410 (N_14410,N_13057,N_13067);
or U14411 (N_14411,N_13036,N_13781);
nand U14412 (N_14412,N_13223,N_13322);
and U14413 (N_14413,N_13973,N_13615);
or U14414 (N_14414,N_13265,N_13220);
xnor U14415 (N_14415,N_13755,N_13805);
or U14416 (N_14416,N_13001,N_13018);
xor U14417 (N_14417,N_13841,N_13161);
nor U14418 (N_14418,N_13429,N_13742);
nand U14419 (N_14419,N_13272,N_13221);
nor U14420 (N_14420,N_13393,N_13988);
and U14421 (N_14421,N_13799,N_13566);
nand U14422 (N_14422,N_13878,N_13383);
and U14423 (N_14423,N_13926,N_13920);
nor U14424 (N_14424,N_13150,N_13813);
and U14425 (N_14425,N_13495,N_13136);
nand U14426 (N_14426,N_13116,N_13965);
xor U14427 (N_14427,N_13623,N_13128);
xor U14428 (N_14428,N_13510,N_13187);
or U14429 (N_14429,N_13508,N_13458);
xnor U14430 (N_14430,N_13609,N_13645);
xnor U14431 (N_14431,N_13400,N_13667);
nor U14432 (N_14432,N_13090,N_13692);
nand U14433 (N_14433,N_13089,N_13985);
and U14434 (N_14434,N_13360,N_13148);
or U14435 (N_14435,N_13255,N_13440);
nand U14436 (N_14436,N_13267,N_13916);
xor U14437 (N_14437,N_13320,N_13764);
or U14438 (N_14438,N_13937,N_13437);
nor U14439 (N_14439,N_13899,N_13367);
and U14440 (N_14440,N_13875,N_13336);
nand U14441 (N_14441,N_13312,N_13688);
nor U14442 (N_14442,N_13299,N_13349);
or U14443 (N_14443,N_13442,N_13502);
xor U14444 (N_14444,N_13338,N_13386);
or U14445 (N_14445,N_13679,N_13114);
or U14446 (N_14446,N_13306,N_13991);
and U14447 (N_14447,N_13877,N_13910);
xor U14448 (N_14448,N_13094,N_13326);
xnor U14449 (N_14449,N_13282,N_13747);
nand U14450 (N_14450,N_13283,N_13478);
xnor U14451 (N_14451,N_13678,N_13748);
or U14452 (N_14452,N_13771,N_13466);
or U14453 (N_14453,N_13703,N_13105);
nand U14454 (N_14454,N_13486,N_13728);
nand U14455 (N_14455,N_13370,N_13694);
and U14456 (N_14456,N_13353,N_13241);
or U14457 (N_14457,N_13818,N_13097);
or U14458 (N_14458,N_13468,N_13475);
nand U14459 (N_14459,N_13589,N_13493);
xor U14460 (N_14460,N_13288,N_13647);
or U14461 (N_14461,N_13111,N_13277);
xor U14462 (N_14462,N_13816,N_13149);
xor U14463 (N_14463,N_13427,N_13660);
nor U14464 (N_14464,N_13002,N_13595);
or U14465 (N_14465,N_13598,N_13022);
and U14466 (N_14466,N_13795,N_13884);
and U14467 (N_14467,N_13860,N_13119);
nor U14468 (N_14468,N_13687,N_13862);
nand U14469 (N_14469,N_13270,N_13290);
xor U14470 (N_14470,N_13297,N_13570);
nor U14471 (N_14471,N_13571,N_13803);
nand U14472 (N_14472,N_13963,N_13575);
xnor U14473 (N_14473,N_13501,N_13736);
and U14474 (N_14474,N_13328,N_13397);
and U14475 (N_14475,N_13695,N_13182);
xor U14476 (N_14476,N_13572,N_13231);
nor U14477 (N_14477,N_13954,N_13947);
or U14478 (N_14478,N_13949,N_13273);
and U14479 (N_14479,N_13219,N_13498);
nand U14480 (N_14480,N_13859,N_13701);
or U14481 (N_14481,N_13683,N_13526);
and U14482 (N_14482,N_13804,N_13365);
xnor U14483 (N_14483,N_13525,N_13345);
xor U14484 (N_14484,N_13640,N_13856);
xnor U14485 (N_14485,N_13224,N_13072);
xnor U14486 (N_14486,N_13868,N_13080);
xnor U14487 (N_14487,N_13676,N_13158);
nor U14488 (N_14488,N_13847,N_13163);
xor U14489 (N_14489,N_13039,N_13760);
xor U14490 (N_14490,N_13431,N_13058);
and U14491 (N_14491,N_13354,N_13156);
nor U14492 (N_14492,N_13981,N_13404);
nor U14493 (N_14493,N_13537,N_13811);
nor U14494 (N_14494,N_13792,N_13278);
and U14495 (N_14495,N_13459,N_13500);
nor U14496 (N_14496,N_13927,N_13013);
and U14497 (N_14497,N_13138,N_13087);
nor U14498 (N_14498,N_13407,N_13782);
and U14499 (N_14499,N_13870,N_13539);
and U14500 (N_14500,N_13286,N_13473);
nor U14501 (N_14501,N_13186,N_13386);
or U14502 (N_14502,N_13820,N_13899);
and U14503 (N_14503,N_13002,N_13991);
nor U14504 (N_14504,N_13978,N_13252);
nor U14505 (N_14505,N_13860,N_13846);
or U14506 (N_14506,N_13710,N_13864);
xor U14507 (N_14507,N_13846,N_13130);
and U14508 (N_14508,N_13194,N_13870);
xnor U14509 (N_14509,N_13700,N_13611);
nor U14510 (N_14510,N_13676,N_13381);
nor U14511 (N_14511,N_13874,N_13974);
and U14512 (N_14512,N_13532,N_13530);
and U14513 (N_14513,N_13225,N_13500);
xnor U14514 (N_14514,N_13647,N_13453);
and U14515 (N_14515,N_13820,N_13083);
or U14516 (N_14516,N_13994,N_13448);
xor U14517 (N_14517,N_13901,N_13751);
nand U14518 (N_14518,N_13042,N_13176);
nor U14519 (N_14519,N_13119,N_13730);
xor U14520 (N_14520,N_13088,N_13717);
nand U14521 (N_14521,N_13903,N_13079);
or U14522 (N_14522,N_13171,N_13259);
nand U14523 (N_14523,N_13129,N_13355);
xnor U14524 (N_14524,N_13274,N_13908);
nor U14525 (N_14525,N_13750,N_13484);
nand U14526 (N_14526,N_13146,N_13990);
nand U14527 (N_14527,N_13425,N_13175);
nor U14528 (N_14528,N_13433,N_13818);
or U14529 (N_14529,N_13095,N_13818);
nand U14530 (N_14530,N_13962,N_13870);
nand U14531 (N_14531,N_13916,N_13437);
nor U14532 (N_14532,N_13906,N_13627);
nor U14533 (N_14533,N_13086,N_13673);
nor U14534 (N_14534,N_13462,N_13761);
xor U14535 (N_14535,N_13255,N_13827);
or U14536 (N_14536,N_13706,N_13675);
or U14537 (N_14537,N_13290,N_13858);
or U14538 (N_14538,N_13121,N_13080);
nor U14539 (N_14539,N_13194,N_13107);
xnor U14540 (N_14540,N_13183,N_13425);
nor U14541 (N_14541,N_13483,N_13438);
nand U14542 (N_14542,N_13407,N_13553);
and U14543 (N_14543,N_13025,N_13810);
nand U14544 (N_14544,N_13094,N_13497);
nor U14545 (N_14545,N_13883,N_13306);
or U14546 (N_14546,N_13409,N_13299);
nor U14547 (N_14547,N_13003,N_13448);
and U14548 (N_14548,N_13496,N_13311);
nor U14549 (N_14549,N_13640,N_13674);
and U14550 (N_14550,N_13858,N_13582);
xnor U14551 (N_14551,N_13351,N_13248);
or U14552 (N_14552,N_13551,N_13731);
nand U14553 (N_14553,N_13299,N_13557);
nor U14554 (N_14554,N_13960,N_13189);
xnor U14555 (N_14555,N_13682,N_13614);
or U14556 (N_14556,N_13792,N_13779);
nor U14557 (N_14557,N_13938,N_13818);
nand U14558 (N_14558,N_13454,N_13502);
nor U14559 (N_14559,N_13537,N_13674);
and U14560 (N_14560,N_13858,N_13036);
xnor U14561 (N_14561,N_13403,N_13690);
xnor U14562 (N_14562,N_13869,N_13501);
nor U14563 (N_14563,N_13905,N_13230);
or U14564 (N_14564,N_13537,N_13187);
nor U14565 (N_14565,N_13756,N_13329);
and U14566 (N_14566,N_13181,N_13978);
or U14567 (N_14567,N_13542,N_13050);
and U14568 (N_14568,N_13934,N_13885);
xor U14569 (N_14569,N_13486,N_13996);
or U14570 (N_14570,N_13930,N_13389);
xor U14571 (N_14571,N_13251,N_13067);
xnor U14572 (N_14572,N_13739,N_13587);
nor U14573 (N_14573,N_13576,N_13358);
xnor U14574 (N_14574,N_13112,N_13323);
and U14575 (N_14575,N_13111,N_13779);
nand U14576 (N_14576,N_13468,N_13966);
nand U14577 (N_14577,N_13375,N_13762);
or U14578 (N_14578,N_13170,N_13174);
or U14579 (N_14579,N_13708,N_13750);
nand U14580 (N_14580,N_13612,N_13197);
nand U14581 (N_14581,N_13204,N_13815);
and U14582 (N_14582,N_13138,N_13342);
nor U14583 (N_14583,N_13850,N_13483);
nor U14584 (N_14584,N_13124,N_13258);
nor U14585 (N_14585,N_13369,N_13086);
xnor U14586 (N_14586,N_13647,N_13883);
xnor U14587 (N_14587,N_13842,N_13511);
xor U14588 (N_14588,N_13312,N_13347);
and U14589 (N_14589,N_13837,N_13031);
xnor U14590 (N_14590,N_13658,N_13615);
xnor U14591 (N_14591,N_13688,N_13870);
xor U14592 (N_14592,N_13619,N_13244);
or U14593 (N_14593,N_13782,N_13528);
xnor U14594 (N_14594,N_13713,N_13000);
and U14595 (N_14595,N_13085,N_13548);
or U14596 (N_14596,N_13685,N_13913);
xnor U14597 (N_14597,N_13682,N_13072);
and U14598 (N_14598,N_13086,N_13902);
nand U14599 (N_14599,N_13212,N_13288);
nor U14600 (N_14600,N_13153,N_13763);
nor U14601 (N_14601,N_13210,N_13073);
xor U14602 (N_14602,N_13321,N_13246);
and U14603 (N_14603,N_13415,N_13177);
xnor U14604 (N_14604,N_13150,N_13582);
nand U14605 (N_14605,N_13159,N_13620);
nor U14606 (N_14606,N_13141,N_13481);
xor U14607 (N_14607,N_13120,N_13210);
nor U14608 (N_14608,N_13001,N_13801);
xor U14609 (N_14609,N_13406,N_13884);
and U14610 (N_14610,N_13397,N_13544);
or U14611 (N_14611,N_13368,N_13869);
xnor U14612 (N_14612,N_13856,N_13009);
and U14613 (N_14613,N_13711,N_13287);
xor U14614 (N_14614,N_13271,N_13155);
nor U14615 (N_14615,N_13928,N_13733);
nor U14616 (N_14616,N_13182,N_13135);
or U14617 (N_14617,N_13938,N_13099);
or U14618 (N_14618,N_13048,N_13841);
nor U14619 (N_14619,N_13947,N_13727);
or U14620 (N_14620,N_13386,N_13937);
and U14621 (N_14621,N_13897,N_13458);
and U14622 (N_14622,N_13804,N_13218);
nand U14623 (N_14623,N_13323,N_13757);
or U14624 (N_14624,N_13207,N_13646);
xnor U14625 (N_14625,N_13101,N_13630);
nor U14626 (N_14626,N_13997,N_13402);
and U14627 (N_14627,N_13539,N_13096);
nand U14628 (N_14628,N_13764,N_13258);
nor U14629 (N_14629,N_13955,N_13816);
or U14630 (N_14630,N_13756,N_13706);
or U14631 (N_14631,N_13647,N_13355);
nand U14632 (N_14632,N_13332,N_13949);
or U14633 (N_14633,N_13009,N_13140);
and U14634 (N_14634,N_13320,N_13745);
nor U14635 (N_14635,N_13545,N_13352);
nand U14636 (N_14636,N_13475,N_13356);
nand U14637 (N_14637,N_13760,N_13614);
and U14638 (N_14638,N_13382,N_13487);
or U14639 (N_14639,N_13688,N_13894);
xor U14640 (N_14640,N_13139,N_13467);
xor U14641 (N_14641,N_13468,N_13576);
or U14642 (N_14642,N_13918,N_13743);
xnor U14643 (N_14643,N_13918,N_13531);
or U14644 (N_14644,N_13319,N_13961);
or U14645 (N_14645,N_13915,N_13450);
and U14646 (N_14646,N_13083,N_13941);
and U14647 (N_14647,N_13126,N_13401);
nand U14648 (N_14648,N_13771,N_13082);
and U14649 (N_14649,N_13432,N_13562);
nand U14650 (N_14650,N_13176,N_13106);
nor U14651 (N_14651,N_13652,N_13418);
or U14652 (N_14652,N_13285,N_13492);
nor U14653 (N_14653,N_13259,N_13150);
or U14654 (N_14654,N_13844,N_13950);
nor U14655 (N_14655,N_13859,N_13954);
xnor U14656 (N_14656,N_13828,N_13178);
nor U14657 (N_14657,N_13032,N_13122);
or U14658 (N_14658,N_13368,N_13633);
nand U14659 (N_14659,N_13891,N_13666);
xor U14660 (N_14660,N_13109,N_13018);
and U14661 (N_14661,N_13588,N_13704);
nand U14662 (N_14662,N_13588,N_13597);
xor U14663 (N_14663,N_13562,N_13416);
nand U14664 (N_14664,N_13337,N_13887);
or U14665 (N_14665,N_13891,N_13385);
or U14666 (N_14666,N_13832,N_13983);
xor U14667 (N_14667,N_13566,N_13540);
or U14668 (N_14668,N_13970,N_13928);
or U14669 (N_14669,N_13472,N_13114);
and U14670 (N_14670,N_13371,N_13586);
nor U14671 (N_14671,N_13355,N_13920);
nand U14672 (N_14672,N_13625,N_13609);
and U14673 (N_14673,N_13822,N_13287);
nor U14674 (N_14674,N_13907,N_13475);
nor U14675 (N_14675,N_13401,N_13245);
xnor U14676 (N_14676,N_13349,N_13946);
and U14677 (N_14677,N_13148,N_13223);
xor U14678 (N_14678,N_13607,N_13885);
nand U14679 (N_14679,N_13459,N_13202);
and U14680 (N_14680,N_13368,N_13636);
nand U14681 (N_14681,N_13885,N_13442);
xnor U14682 (N_14682,N_13594,N_13797);
nor U14683 (N_14683,N_13532,N_13475);
xor U14684 (N_14684,N_13832,N_13098);
nor U14685 (N_14685,N_13005,N_13918);
nand U14686 (N_14686,N_13924,N_13572);
nand U14687 (N_14687,N_13830,N_13974);
or U14688 (N_14688,N_13743,N_13800);
and U14689 (N_14689,N_13094,N_13793);
nand U14690 (N_14690,N_13311,N_13440);
or U14691 (N_14691,N_13439,N_13704);
and U14692 (N_14692,N_13283,N_13534);
xor U14693 (N_14693,N_13743,N_13792);
xor U14694 (N_14694,N_13833,N_13394);
nand U14695 (N_14695,N_13523,N_13189);
nand U14696 (N_14696,N_13588,N_13955);
nand U14697 (N_14697,N_13208,N_13659);
or U14698 (N_14698,N_13493,N_13602);
and U14699 (N_14699,N_13013,N_13221);
xor U14700 (N_14700,N_13731,N_13382);
or U14701 (N_14701,N_13135,N_13761);
and U14702 (N_14702,N_13449,N_13865);
nor U14703 (N_14703,N_13015,N_13174);
and U14704 (N_14704,N_13697,N_13756);
nand U14705 (N_14705,N_13955,N_13872);
nand U14706 (N_14706,N_13523,N_13237);
nor U14707 (N_14707,N_13685,N_13063);
and U14708 (N_14708,N_13545,N_13595);
or U14709 (N_14709,N_13398,N_13778);
nor U14710 (N_14710,N_13058,N_13109);
nand U14711 (N_14711,N_13840,N_13207);
nor U14712 (N_14712,N_13772,N_13713);
or U14713 (N_14713,N_13815,N_13641);
nor U14714 (N_14714,N_13999,N_13424);
nand U14715 (N_14715,N_13564,N_13766);
and U14716 (N_14716,N_13862,N_13556);
nand U14717 (N_14717,N_13784,N_13869);
nand U14718 (N_14718,N_13169,N_13449);
xnor U14719 (N_14719,N_13667,N_13014);
nor U14720 (N_14720,N_13425,N_13812);
and U14721 (N_14721,N_13849,N_13351);
or U14722 (N_14722,N_13960,N_13669);
nor U14723 (N_14723,N_13950,N_13817);
nand U14724 (N_14724,N_13506,N_13189);
and U14725 (N_14725,N_13256,N_13686);
nand U14726 (N_14726,N_13713,N_13414);
nor U14727 (N_14727,N_13140,N_13535);
nand U14728 (N_14728,N_13136,N_13985);
nand U14729 (N_14729,N_13402,N_13882);
and U14730 (N_14730,N_13630,N_13901);
nor U14731 (N_14731,N_13636,N_13737);
and U14732 (N_14732,N_13305,N_13282);
or U14733 (N_14733,N_13170,N_13915);
xor U14734 (N_14734,N_13212,N_13284);
xnor U14735 (N_14735,N_13421,N_13433);
and U14736 (N_14736,N_13914,N_13348);
or U14737 (N_14737,N_13960,N_13070);
or U14738 (N_14738,N_13414,N_13445);
or U14739 (N_14739,N_13453,N_13881);
nand U14740 (N_14740,N_13864,N_13570);
nand U14741 (N_14741,N_13285,N_13175);
xor U14742 (N_14742,N_13751,N_13596);
and U14743 (N_14743,N_13600,N_13238);
nor U14744 (N_14744,N_13844,N_13663);
and U14745 (N_14745,N_13714,N_13456);
xor U14746 (N_14746,N_13172,N_13406);
xor U14747 (N_14747,N_13172,N_13627);
and U14748 (N_14748,N_13248,N_13657);
or U14749 (N_14749,N_13034,N_13368);
nand U14750 (N_14750,N_13330,N_13020);
or U14751 (N_14751,N_13123,N_13914);
xor U14752 (N_14752,N_13632,N_13426);
nand U14753 (N_14753,N_13741,N_13808);
and U14754 (N_14754,N_13061,N_13430);
xnor U14755 (N_14755,N_13337,N_13081);
or U14756 (N_14756,N_13152,N_13798);
xor U14757 (N_14757,N_13349,N_13875);
nand U14758 (N_14758,N_13742,N_13733);
nand U14759 (N_14759,N_13770,N_13693);
and U14760 (N_14760,N_13420,N_13925);
and U14761 (N_14761,N_13717,N_13049);
nor U14762 (N_14762,N_13365,N_13247);
nor U14763 (N_14763,N_13402,N_13787);
nand U14764 (N_14764,N_13569,N_13233);
nor U14765 (N_14765,N_13047,N_13169);
nor U14766 (N_14766,N_13094,N_13182);
nor U14767 (N_14767,N_13165,N_13152);
nor U14768 (N_14768,N_13269,N_13036);
nand U14769 (N_14769,N_13324,N_13156);
xnor U14770 (N_14770,N_13903,N_13067);
or U14771 (N_14771,N_13451,N_13587);
or U14772 (N_14772,N_13627,N_13958);
and U14773 (N_14773,N_13670,N_13500);
nand U14774 (N_14774,N_13963,N_13704);
nor U14775 (N_14775,N_13328,N_13150);
xor U14776 (N_14776,N_13753,N_13876);
or U14777 (N_14777,N_13472,N_13673);
and U14778 (N_14778,N_13445,N_13693);
xor U14779 (N_14779,N_13644,N_13988);
and U14780 (N_14780,N_13422,N_13711);
nand U14781 (N_14781,N_13730,N_13112);
nand U14782 (N_14782,N_13990,N_13004);
nor U14783 (N_14783,N_13485,N_13807);
xnor U14784 (N_14784,N_13371,N_13760);
or U14785 (N_14785,N_13914,N_13028);
nor U14786 (N_14786,N_13337,N_13692);
nand U14787 (N_14787,N_13481,N_13755);
and U14788 (N_14788,N_13711,N_13306);
nand U14789 (N_14789,N_13921,N_13447);
and U14790 (N_14790,N_13291,N_13286);
or U14791 (N_14791,N_13231,N_13643);
nand U14792 (N_14792,N_13222,N_13708);
and U14793 (N_14793,N_13951,N_13826);
and U14794 (N_14794,N_13073,N_13384);
or U14795 (N_14795,N_13103,N_13804);
and U14796 (N_14796,N_13223,N_13533);
and U14797 (N_14797,N_13753,N_13180);
or U14798 (N_14798,N_13220,N_13014);
nand U14799 (N_14799,N_13904,N_13485);
and U14800 (N_14800,N_13253,N_13296);
and U14801 (N_14801,N_13980,N_13331);
xor U14802 (N_14802,N_13137,N_13810);
xor U14803 (N_14803,N_13136,N_13583);
nand U14804 (N_14804,N_13568,N_13457);
or U14805 (N_14805,N_13471,N_13922);
or U14806 (N_14806,N_13440,N_13370);
xnor U14807 (N_14807,N_13785,N_13407);
nand U14808 (N_14808,N_13236,N_13198);
nor U14809 (N_14809,N_13491,N_13943);
nand U14810 (N_14810,N_13770,N_13502);
xnor U14811 (N_14811,N_13635,N_13005);
or U14812 (N_14812,N_13108,N_13512);
xor U14813 (N_14813,N_13436,N_13617);
nor U14814 (N_14814,N_13331,N_13699);
nor U14815 (N_14815,N_13965,N_13440);
nor U14816 (N_14816,N_13653,N_13314);
nand U14817 (N_14817,N_13313,N_13459);
and U14818 (N_14818,N_13736,N_13649);
nor U14819 (N_14819,N_13872,N_13376);
and U14820 (N_14820,N_13389,N_13236);
or U14821 (N_14821,N_13140,N_13402);
nand U14822 (N_14822,N_13295,N_13753);
nand U14823 (N_14823,N_13858,N_13987);
or U14824 (N_14824,N_13747,N_13695);
nand U14825 (N_14825,N_13473,N_13200);
or U14826 (N_14826,N_13428,N_13215);
xor U14827 (N_14827,N_13797,N_13104);
nand U14828 (N_14828,N_13389,N_13223);
and U14829 (N_14829,N_13078,N_13099);
xnor U14830 (N_14830,N_13778,N_13327);
nor U14831 (N_14831,N_13555,N_13775);
nor U14832 (N_14832,N_13902,N_13673);
xor U14833 (N_14833,N_13416,N_13432);
xnor U14834 (N_14834,N_13095,N_13140);
nand U14835 (N_14835,N_13488,N_13938);
and U14836 (N_14836,N_13048,N_13836);
nor U14837 (N_14837,N_13263,N_13488);
and U14838 (N_14838,N_13961,N_13860);
nor U14839 (N_14839,N_13345,N_13011);
nor U14840 (N_14840,N_13645,N_13454);
or U14841 (N_14841,N_13709,N_13254);
nor U14842 (N_14842,N_13103,N_13838);
nand U14843 (N_14843,N_13946,N_13228);
or U14844 (N_14844,N_13551,N_13176);
nor U14845 (N_14845,N_13506,N_13515);
xnor U14846 (N_14846,N_13973,N_13667);
nand U14847 (N_14847,N_13983,N_13120);
nor U14848 (N_14848,N_13184,N_13455);
nand U14849 (N_14849,N_13602,N_13529);
nand U14850 (N_14850,N_13801,N_13630);
nand U14851 (N_14851,N_13754,N_13287);
or U14852 (N_14852,N_13386,N_13968);
or U14853 (N_14853,N_13338,N_13783);
xor U14854 (N_14854,N_13766,N_13182);
nand U14855 (N_14855,N_13042,N_13297);
or U14856 (N_14856,N_13700,N_13467);
nor U14857 (N_14857,N_13791,N_13431);
and U14858 (N_14858,N_13061,N_13324);
xnor U14859 (N_14859,N_13208,N_13566);
xnor U14860 (N_14860,N_13408,N_13872);
nand U14861 (N_14861,N_13984,N_13354);
and U14862 (N_14862,N_13796,N_13492);
nand U14863 (N_14863,N_13212,N_13923);
or U14864 (N_14864,N_13971,N_13237);
and U14865 (N_14865,N_13944,N_13401);
nor U14866 (N_14866,N_13179,N_13237);
nand U14867 (N_14867,N_13279,N_13388);
nand U14868 (N_14868,N_13976,N_13003);
and U14869 (N_14869,N_13899,N_13585);
xnor U14870 (N_14870,N_13250,N_13270);
or U14871 (N_14871,N_13378,N_13568);
xor U14872 (N_14872,N_13895,N_13317);
xnor U14873 (N_14873,N_13289,N_13357);
nor U14874 (N_14874,N_13185,N_13659);
nand U14875 (N_14875,N_13166,N_13649);
nand U14876 (N_14876,N_13964,N_13097);
or U14877 (N_14877,N_13385,N_13570);
nor U14878 (N_14878,N_13755,N_13435);
xnor U14879 (N_14879,N_13409,N_13310);
xor U14880 (N_14880,N_13079,N_13597);
xor U14881 (N_14881,N_13706,N_13198);
xor U14882 (N_14882,N_13922,N_13596);
nand U14883 (N_14883,N_13046,N_13174);
and U14884 (N_14884,N_13229,N_13302);
nor U14885 (N_14885,N_13172,N_13826);
xor U14886 (N_14886,N_13302,N_13663);
nand U14887 (N_14887,N_13541,N_13943);
nor U14888 (N_14888,N_13950,N_13858);
or U14889 (N_14889,N_13887,N_13744);
nor U14890 (N_14890,N_13869,N_13878);
or U14891 (N_14891,N_13826,N_13037);
nor U14892 (N_14892,N_13620,N_13958);
and U14893 (N_14893,N_13577,N_13725);
nor U14894 (N_14894,N_13981,N_13704);
or U14895 (N_14895,N_13191,N_13303);
nand U14896 (N_14896,N_13265,N_13611);
xnor U14897 (N_14897,N_13978,N_13910);
xor U14898 (N_14898,N_13546,N_13954);
and U14899 (N_14899,N_13211,N_13007);
or U14900 (N_14900,N_13850,N_13165);
xnor U14901 (N_14901,N_13681,N_13485);
and U14902 (N_14902,N_13832,N_13965);
or U14903 (N_14903,N_13335,N_13374);
nor U14904 (N_14904,N_13561,N_13172);
and U14905 (N_14905,N_13076,N_13426);
xnor U14906 (N_14906,N_13274,N_13264);
xor U14907 (N_14907,N_13628,N_13695);
xor U14908 (N_14908,N_13327,N_13605);
nor U14909 (N_14909,N_13458,N_13975);
xor U14910 (N_14910,N_13686,N_13693);
or U14911 (N_14911,N_13669,N_13658);
and U14912 (N_14912,N_13576,N_13773);
nand U14913 (N_14913,N_13850,N_13266);
xnor U14914 (N_14914,N_13896,N_13491);
and U14915 (N_14915,N_13444,N_13584);
xor U14916 (N_14916,N_13451,N_13734);
nand U14917 (N_14917,N_13499,N_13020);
and U14918 (N_14918,N_13632,N_13950);
and U14919 (N_14919,N_13345,N_13654);
or U14920 (N_14920,N_13353,N_13708);
or U14921 (N_14921,N_13835,N_13338);
xnor U14922 (N_14922,N_13761,N_13747);
nand U14923 (N_14923,N_13634,N_13447);
or U14924 (N_14924,N_13050,N_13668);
nor U14925 (N_14925,N_13282,N_13738);
or U14926 (N_14926,N_13248,N_13470);
nor U14927 (N_14927,N_13844,N_13693);
nand U14928 (N_14928,N_13343,N_13594);
nor U14929 (N_14929,N_13914,N_13405);
nand U14930 (N_14930,N_13355,N_13197);
nor U14931 (N_14931,N_13919,N_13895);
xor U14932 (N_14932,N_13949,N_13315);
or U14933 (N_14933,N_13277,N_13614);
or U14934 (N_14934,N_13179,N_13871);
nand U14935 (N_14935,N_13234,N_13348);
xor U14936 (N_14936,N_13459,N_13870);
or U14937 (N_14937,N_13734,N_13971);
or U14938 (N_14938,N_13842,N_13664);
and U14939 (N_14939,N_13706,N_13883);
and U14940 (N_14940,N_13191,N_13651);
xor U14941 (N_14941,N_13468,N_13116);
nand U14942 (N_14942,N_13332,N_13037);
and U14943 (N_14943,N_13205,N_13446);
nor U14944 (N_14944,N_13227,N_13641);
and U14945 (N_14945,N_13750,N_13499);
or U14946 (N_14946,N_13235,N_13541);
xor U14947 (N_14947,N_13247,N_13858);
xor U14948 (N_14948,N_13336,N_13293);
and U14949 (N_14949,N_13727,N_13996);
xor U14950 (N_14950,N_13562,N_13564);
or U14951 (N_14951,N_13453,N_13000);
and U14952 (N_14952,N_13615,N_13389);
and U14953 (N_14953,N_13517,N_13898);
nand U14954 (N_14954,N_13256,N_13105);
nand U14955 (N_14955,N_13644,N_13536);
or U14956 (N_14956,N_13806,N_13587);
nand U14957 (N_14957,N_13985,N_13798);
and U14958 (N_14958,N_13069,N_13306);
or U14959 (N_14959,N_13349,N_13213);
nand U14960 (N_14960,N_13312,N_13879);
nor U14961 (N_14961,N_13340,N_13513);
nor U14962 (N_14962,N_13279,N_13968);
xor U14963 (N_14963,N_13656,N_13908);
and U14964 (N_14964,N_13141,N_13626);
and U14965 (N_14965,N_13672,N_13433);
nand U14966 (N_14966,N_13347,N_13712);
or U14967 (N_14967,N_13389,N_13316);
and U14968 (N_14968,N_13225,N_13132);
xnor U14969 (N_14969,N_13972,N_13799);
or U14970 (N_14970,N_13878,N_13436);
and U14971 (N_14971,N_13249,N_13739);
nand U14972 (N_14972,N_13236,N_13912);
nand U14973 (N_14973,N_13967,N_13892);
xor U14974 (N_14974,N_13050,N_13090);
and U14975 (N_14975,N_13393,N_13958);
or U14976 (N_14976,N_13318,N_13018);
nor U14977 (N_14977,N_13439,N_13662);
or U14978 (N_14978,N_13116,N_13290);
nand U14979 (N_14979,N_13955,N_13480);
nor U14980 (N_14980,N_13204,N_13936);
nor U14981 (N_14981,N_13322,N_13956);
xor U14982 (N_14982,N_13821,N_13162);
and U14983 (N_14983,N_13805,N_13044);
xnor U14984 (N_14984,N_13234,N_13815);
nand U14985 (N_14985,N_13776,N_13887);
nor U14986 (N_14986,N_13252,N_13439);
and U14987 (N_14987,N_13504,N_13356);
nand U14988 (N_14988,N_13752,N_13705);
and U14989 (N_14989,N_13100,N_13037);
xnor U14990 (N_14990,N_13827,N_13238);
and U14991 (N_14991,N_13544,N_13647);
nor U14992 (N_14992,N_13329,N_13894);
nand U14993 (N_14993,N_13325,N_13680);
nand U14994 (N_14994,N_13524,N_13649);
nand U14995 (N_14995,N_13376,N_13903);
and U14996 (N_14996,N_13218,N_13489);
xnor U14997 (N_14997,N_13094,N_13285);
nor U14998 (N_14998,N_13468,N_13785);
nor U14999 (N_14999,N_13354,N_13549);
xnor U15000 (N_15000,N_14089,N_14747);
or U15001 (N_15001,N_14495,N_14347);
xor U15002 (N_15002,N_14986,N_14081);
and U15003 (N_15003,N_14267,N_14927);
and U15004 (N_15004,N_14360,N_14162);
nor U15005 (N_15005,N_14981,N_14186);
and U15006 (N_15006,N_14296,N_14865);
xor U15007 (N_15007,N_14717,N_14300);
and U15008 (N_15008,N_14657,N_14402);
nand U15009 (N_15009,N_14197,N_14555);
nand U15010 (N_15010,N_14893,N_14411);
nor U15011 (N_15011,N_14547,N_14899);
nand U15012 (N_15012,N_14769,N_14345);
xor U15013 (N_15013,N_14012,N_14118);
or U15014 (N_15014,N_14781,N_14131);
and U15015 (N_15015,N_14768,N_14970);
or U15016 (N_15016,N_14286,N_14892);
nand U15017 (N_15017,N_14461,N_14193);
or U15018 (N_15018,N_14835,N_14082);
xor U15019 (N_15019,N_14706,N_14280);
xor U15020 (N_15020,N_14651,N_14303);
xnor U15021 (N_15021,N_14984,N_14056);
xnor U15022 (N_15022,N_14189,N_14240);
nor U15023 (N_15023,N_14227,N_14766);
xor U15024 (N_15024,N_14611,N_14932);
nor U15025 (N_15025,N_14423,N_14649);
and U15026 (N_15026,N_14204,N_14053);
nor U15027 (N_15027,N_14359,N_14900);
nand U15028 (N_15028,N_14704,N_14966);
xnor U15029 (N_15029,N_14285,N_14687);
or U15030 (N_15030,N_14061,N_14613);
and U15031 (N_15031,N_14075,N_14940);
or U15032 (N_15032,N_14665,N_14109);
xnor U15033 (N_15033,N_14178,N_14748);
and U15034 (N_15034,N_14920,N_14770);
or U15035 (N_15035,N_14701,N_14369);
or U15036 (N_15036,N_14339,N_14074);
or U15037 (N_15037,N_14046,N_14225);
nor U15038 (N_15038,N_14678,N_14585);
xnor U15039 (N_15039,N_14034,N_14011);
nand U15040 (N_15040,N_14365,N_14887);
or U15041 (N_15041,N_14564,N_14808);
xor U15042 (N_15042,N_14840,N_14960);
xnor U15043 (N_15043,N_14543,N_14854);
xor U15044 (N_15044,N_14179,N_14834);
and U15045 (N_15045,N_14608,N_14630);
nand U15046 (N_15046,N_14432,N_14507);
nand U15047 (N_15047,N_14526,N_14381);
nor U15048 (N_15048,N_14083,N_14644);
or U15049 (N_15049,N_14888,N_14048);
and U15050 (N_15050,N_14326,N_14418);
and U15051 (N_15051,N_14260,N_14828);
nor U15052 (N_15052,N_14950,N_14801);
and U15053 (N_15053,N_14764,N_14372);
nand U15054 (N_15054,N_14815,N_14894);
nand U15055 (N_15055,N_14389,N_14831);
and U15056 (N_15056,N_14362,N_14095);
nor U15057 (N_15057,N_14698,N_14667);
nand U15058 (N_15058,N_14187,N_14292);
and U15059 (N_15059,N_14924,N_14107);
xnor U15060 (N_15060,N_14587,N_14420);
and U15061 (N_15061,N_14895,N_14858);
or U15062 (N_15062,N_14168,N_14029);
nor U15063 (N_15063,N_14444,N_14383);
nor U15064 (N_15064,N_14914,N_14897);
and U15065 (N_15065,N_14597,N_14263);
nand U15066 (N_15066,N_14164,N_14876);
and U15067 (N_15067,N_14404,N_14689);
nor U15068 (N_15068,N_14491,N_14958);
nor U15069 (N_15069,N_14196,N_14645);
and U15070 (N_15070,N_14295,N_14283);
nor U15071 (N_15071,N_14250,N_14980);
or U15072 (N_15072,N_14321,N_14972);
and U15073 (N_15073,N_14489,N_14836);
nand U15074 (N_15074,N_14134,N_14494);
nand U15075 (N_15075,N_14675,N_14505);
nand U15076 (N_15076,N_14155,N_14376);
nor U15077 (N_15077,N_14301,N_14676);
xor U15078 (N_15078,N_14382,N_14013);
xnor U15079 (N_15079,N_14143,N_14680);
or U15080 (N_15080,N_14414,N_14968);
and U15081 (N_15081,N_14396,N_14331);
nor U15082 (N_15082,N_14860,N_14621);
xor U15083 (N_15083,N_14985,N_14614);
nand U15084 (N_15084,N_14310,N_14610);
and U15085 (N_15085,N_14846,N_14291);
xnor U15086 (N_15086,N_14503,N_14567);
nand U15087 (N_15087,N_14866,N_14115);
xor U15088 (N_15088,N_14631,N_14108);
nand U15089 (N_15089,N_14424,N_14007);
nand U15090 (N_15090,N_14111,N_14745);
and U15091 (N_15091,N_14758,N_14742);
xor U15092 (N_15092,N_14504,N_14125);
or U15093 (N_15093,N_14902,N_14415);
and U15094 (N_15094,N_14379,N_14183);
nand U15095 (N_15095,N_14563,N_14009);
or U15096 (N_15096,N_14730,N_14150);
nor U15097 (N_15097,N_14071,N_14599);
and U15098 (N_15098,N_14190,N_14992);
and U15099 (N_15099,N_14248,N_14732);
xnor U15100 (N_15100,N_14774,N_14441);
nand U15101 (N_15101,N_14579,N_14949);
and U15102 (N_15102,N_14664,N_14670);
or U15103 (N_15103,N_14219,N_14609);
xor U15104 (N_15104,N_14635,N_14752);
and U15105 (N_15105,N_14884,N_14064);
xnor U15106 (N_15106,N_14384,N_14492);
nand U15107 (N_15107,N_14575,N_14161);
xnor U15108 (N_15108,N_14625,N_14158);
nor U15109 (N_15109,N_14642,N_14775);
and U15110 (N_15110,N_14661,N_14788);
or U15111 (N_15111,N_14440,N_14400);
nor U15112 (N_15112,N_14998,N_14978);
and U15113 (N_15113,N_14031,N_14983);
and U15114 (N_15114,N_14697,N_14232);
xor U15115 (N_15115,N_14032,N_14080);
nand U15116 (N_15116,N_14088,N_14103);
or U15117 (N_15117,N_14800,N_14353);
xor U15118 (N_15118,N_14911,N_14184);
nor U15119 (N_15119,N_14206,N_14238);
xor U15120 (N_15120,N_14929,N_14794);
nor U15121 (N_15121,N_14050,N_14915);
nand U15122 (N_15122,N_14205,N_14332);
and U15123 (N_15123,N_14553,N_14349);
and U15124 (N_15124,N_14044,N_14956);
xor U15125 (N_15125,N_14410,N_14090);
xnor U15126 (N_15126,N_14133,N_14746);
nand U15127 (N_15127,N_14693,N_14191);
xnor U15128 (N_15128,N_14449,N_14485);
xor U15129 (N_15129,N_14991,N_14925);
nor U15130 (N_15130,N_14595,N_14091);
and U15131 (N_15131,N_14037,N_14928);
nor U15132 (N_15132,N_14772,N_14535);
nand U15133 (N_15133,N_14576,N_14761);
and U15134 (N_15134,N_14959,N_14817);
nor U15135 (N_15135,N_14167,N_14848);
nand U15136 (N_15136,N_14935,N_14026);
and U15137 (N_15137,N_14798,N_14122);
nand U15138 (N_15138,N_14076,N_14603);
and U15139 (N_15139,N_14216,N_14106);
xor U15140 (N_15140,N_14662,N_14528);
nand U15141 (N_15141,N_14307,N_14853);
nor U15142 (N_15142,N_14316,N_14674);
nor U15143 (N_15143,N_14428,N_14964);
or U15144 (N_15144,N_14215,N_14207);
nor U15145 (N_15145,N_14456,N_14348);
xnor U15146 (N_15146,N_14738,N_14004);
or U15147 (N_15147,N_14923,N_14171);
nand U15148 (N_15148,N_14508,N_14509);
xnor U15149 (N_15149,N_14040,N_14878);
nor U15150 (N_15150,N_14357,N_14656);
or U15151 (N_15151,N_14198,N_14045);
or U15152 (N_15152,N_14500,N_14862);
nor U15153 (N_15153,N_14429,N_14018);
nor U15154 (N_15154,N_14014,N_14921);
xnor U15155 (N_15155,N_14453,N_14713);
nand U15156 (N_15156,N_14773,N_14129);
nand U15157 (N_15157,N_14350,N_14487);
nor U15158 (N_15158,N_14600,N_14623);
or U15159 (N_15159,N_14844,N_14533);
or U15160 (N_15160,N_14364,N_14582);
and U15161 (N_15161,N_14025,N_14245);
nand U15162 (N_15162,N_14833,N_14476);
nand U15163 (N_15163,N_14974,N_14138);
or U15164 (N_15164,N_14692,N_14266);
nand U15165 (N_15165,N_14536,N_14633);
nand U15166 (N_15166,N_14521,N_14721);
or U15167 (N_15167,N_14757,N_14142);
and U15168 (N_15168,N_14629,N_14513);
nand U15169 (N_15169,N_14087,N_14430);
and U15170 (N_15170,N_14110,N_14446);
or U15171 (N_15171,N_14017,N_14518);
and U15172 (N_15172,N_14628,N_14636);
or U15173 (N_15173,N_14727,N_14851);
and U15174 (N_15174,N_14308,N_14724);
or U15175 (N_15175,N_14023,N_14767);
xor U15176 (N_15176,N_14220,N_14673);
and U15177 (N_15177,N_14361,N_14395);
xnor U15178 (N_15178,N_14159,N_14417);
and U15179 (N_15179,N_14523,N_14367);
and U15180 (N_15180,N_14455,N_14457);
or U15181 (N_15181,N_14021,N_14254);
or U15182 (N_15182,N_14471,N_14392);
nor U15183 (N_15183,N_14030,N_14114);
nand U15184 (N_15184,N_14473,N_14284);
or U15185 (N_15185,N_14722,N_14314);
nand U15186 (N_15186,N_14771,N_14099);
or U15187 (N_15187,N_14463,N_14971);
nor U15188 (N_15188,N_14059,N_14522);
and U15189 (N_15189,N_14409,N_14313);
xor U15190 (N_15190,N_14156,N_14538);
and U15191 (N_15191,N_14826,N_14136);
or U15192 (N_15192,N_14468,N_14304);
or U15193 (N_15193,N_14639,N_14231);
nand U15194 (N_15194,N_14646,N_14258);
nand U15195 (N_15195,N_14945,N_14439);
and U15196 (N_15196,N_14907,N_14256);
xor U15197 (N_15197,N_14065,N_14351);
nor U15198 (N_15198,N_14333,N_14824);
nor U15199 (N_15199,N_14627,N_14632);
nor U15200 (N_15200,N_14062,N_14294);
and U15201 (N_15201,N_14228,N_14847);
nand U15202 (N_15202,N_14224,N_14965);
or U15203 (N_15203,N_14917,N_14281);
nand U15204 (N_15204,N_14754,N_14490);
nor U15205 (N_15205,N_14837,N_14330);
and U15206 (N_15206,N_14253,N_14696);
xnor U15207 (N_15207,N_14527,N_14789);
and U15208 (N_15208,N_14434,N_14967);
nand U15209 (N_15209,N_14070,N_14211);
and U15210 (N_15210,N_14055,N_14270);
and U15211 (N_15211,N_14883,N_14908);
or U15212 (N_15212,N_14856,N_14782);
xnor U15213 (N_15213,N_14058,N_14822);
xor U15214 (N_15214,N_14290,N_14530);
nand U15215 (N_15215,N_14277,N_14130);
nand U15216 (N_15216,N_14711,N_14057);
and U15217 (N_15217,N_14319,N_14702);
xor U15218 (N_15218,N_14885,N_14811);
xnor U15219 (N_15219,N_14556,N_14501);
nand U15220 (N_15220,N_14024,N_14243);
xnor U15221 (N_15221,N_14804,N_14723);
xnor U15222 (N_15222,N_14868,N_14830);
and U15223 (N_15223,N_14352,N_14340);
or U15224 (N_15224,N_14433,N_14545);
or U15225 (N_15225,N_14199,N_14092);
and U15226 (N_15226,N_14787,N_14244);
nand U15227 (N_15227,N_14705,N_14712);
and U15228 (N_15228,N_14760,N_14126);
or U15229 (N_15229,N_14317,N_14117);
or U15230 (N_15230,N_14222,N_14707);
or U15231 (N_15231,N_14470,N_14719);
nand U15232 (N_15232,N_14279,N_14241);
and U15233 (N_15233,N_14309,N_14650);
xor U15234 (N_15234,N_14944,N_14480);
nand U15235 (N_15235,N_14035,N_14478);
and U15236 (N_15236,N_14979,N_14010);
or U15237 (N_15237,N_14648,N_14094);
nor U15238 (N_15238,N_14934,N_14042);
or U15239 (N_15239,N_14652,N_14618);
and U15240 (N_15240,N_14413,N_14584);
nand U15241 (N_15241,N_14861,N_14436);
xnor U15242 (N_15242,N_14085,N_14829);
or U15243 (N_15243,N_14688,N_14268);
or U15244 (N_15244,N_14412,N_14969);
nor U15245 (N_15245,N_14852,N_14939);
nand U15246 (N_15246,N_14904,N_14212);
and U15247 (N_15247,N_14666,N_14322);
nor U15248 (N_15248,N_14873,N_14496);
nor U15249 (N_15249,N_14259,N_14141);
nor U15250 (N_15250,N_14278,N_14020);
nor U15251 (N_15251,N_14948,N_14566);
or U15252 (N_15252,N_14481,N_14843);
xnor U15253 (N_15253,N_14452,N_14443);
nand U15254 (N_15254,N_14229,N_14954);
nor U15255 (N_15255,N_14957,N_14398);
xnor U15256 (N_15256,N_14683,N_14931);
xnor U15257 (N_15257,N_14063,N_14663);
nand U15258 (N_15258,N_14438,N_14731);
xor U15259 (N_15259,N_14825,N_14990);
and U15260 (N_15260,N_14377,N_14881);
or U15261 (N_15261,N_14407,N_14919);
xnor U15262 (N_15262,N_14421,N_14202);
nor U15263 (N_15263,N_14519,N_14262);
nand U15264 (N_15264,N_14778,N_14640);
or U15265 (N_15265,N_14735,N_14235);
and U15266 (N_15266,N_14725,N_14736);
or U15267 (N_15267,N_14341,N_14586);
nor U15268 (N_15268,N_14849,N_14975);
nand U15269 (N_15269,N_14247,N_14390);
or U15270 (N_15270,N_14298,N_14318);
or U15271 (N_15271,N_14820,N_14716);
nand U15272 (N_15272,N_14976,N_14550);
and U15273 (N_15273,N_14234,N_14226);
nor U15274 (N_15274,N_14174,N_14388);
and U15275 (N_15275,N_14137,N_14249);
and U15276 (N_15276,N_14022,N_14839);
and U15277 (N_15277,N_14203,N_14751);
nor U15278 (N_15278,N_14146,N_14066);
or U15279 (N_15279,N_14669,N_14151);
nand U15280 (N_15280,N_14874,N_14261);
nor U15281 (N_15281,N_14139,N_14739);
and U15282 (N_15282,N_14242,N_14072);
and U15283 (N_15283,N_14544,N_14889);
xor U15284 (N_15284,N_14938,N_14877);
and U15285 (N_15285,N_14378,N_14510);
xor U15286 (N_15286,N_14287,N_14546);
or U15287 (N_15287,N_14880,N_14098);
nor U15288 (N_15288,N_14016,N_14548);
nor U15289 (N_15289,N_14431,N_14568);
or U15290 (N_15290,N_14387,N_14454);
nand U15291 (N_15291,N_14185,N_14819);
nor U15292 (N_15292,N_14329,N_14426);
and U15293 (N_15293,N_14459,N_14619);
or U15294 (N_15294,N_14274,N_14482);
nand U15295 (N_15295,N_14905,N_14565);
nor U15296 (N_15296,N_14160,N_14132);
xnor U15297 (N_15297,N_14346,N_14105);
and U15298 (N_15298,N_14246,N_14344);
nand U15299 (N_15299,N_14394,N_14943);
and U15300 (N_15300,N_14909,N_14622);
nor U15301 (N_15301,N_14593,N_14660);
xnor U15302 (N_15302,N_14451,N_14315);
nand U15303 (N_15303,N_14408,N_14176);
or U15304 (N_15304,N_14233,N_14078);
nand U15305 (N_15305,N_14996,N_14741);
nor U15306 (N_15306,N_14542,N_14524);
xor U15307 (N_15307,N_14729,N_14684);
or U15308 (N_15308,N_14192,N_14520);
and U15309 (N_15309,N_14583,N_14734);
nor U15310 (N_15310,N_14560,N_14264);
nor U15311 (N_15311,N_14571,N_14539);
xnor U15312 (N_15312,N_14681,N_14120);
xnor U15313 (N_15313,N_14867,N_14901);
xor U15314 (N_15314,N_14643,N_14615);
and U15315 (N_15315,N_14994,N_14784);
nor U15316 (N_15316,N_14805,N_14323);
nor U15317 (N_15317,N_14437,N_14755);
xor U15318 (N_15318,N_14799,N_14872);
nor U15319 (N_15319,N_14276,N_14282);
nor U15320 (N_15320,N_14015,N_14488);
and U15321 (N_15321,N_14785,N_14373);
xor U15322 (N_15322,N_14855,N_14606);
nor U15323 (N_15323,N_14325,N_14910);
nor U15324 (N_15324,N_14149,N_14366);
and U15325 (N_15325,N_14715,N_14355);
nor U15326 (N_15326,N_14416,N_14561);
xor U15327 (N_15327,N_14779,N_14783);
nor U15328 (N_15328,N_14517,N_14653);
nand U15329 (N_15329,N_14821,N_14690);
or U15330 (N_15330,N_14493,N_14685);
xnor U15331 (N_15331,N_14882,N_14385);
nand U15332 (N_15332,N_14208,N_14067);
nor U15333 (N_15333,N_14695,N_14620);
or U15334 (N_15334,N_14054,N_14272);
nor U15335 (N_15335,N_14857,N_14525);
and U15336 (N_15336,N_14218,N_14896);
or U15337 (N_15337,N_14006,N_14638);
xnor U15338 (N_15338,N_14484,N_14273);
and U15339 (N_15339,N_14327,N_14918);
nand U15340 (N_15340,N_14467,N_14955);
nand U15341 (N_15341,N_14047,N_14708);
or U15342 (N_15342,N_14947,N_14079);
or U15343 (N_15343,N_14589,N_14569);
xor U15344 (N_15344,N_14818,N_14864);
nor U15345 (N_15345,N_14210,N_14119);
and U15346 (N_15346,N_14093,N_14588);
or U15347 (N_15347,N_14374,N_14338);
and U15348 (N_15348,N_14827,N_14195);
nor U15349 (N_15349,N_14871,N_14356);
xor U15350 (N_15350,N_14617,N_14406);
nor U15351 (N_15351,N_14127,N_14534);
and U15352 (N_15352,N_14634,N_14182);
or U15353 (N_15353,N_14709,N_14759);
xor U15354 (N_15354,N_14305,N_14405);
xnor U15355 (N_15355,N_14573,N_14570);
or U15356 (N_15356,N_14624,N_14435);
or U15357 (N_15357,N_14288,N_14401);
nor U15358 (N_15358,N_14989,N_14194);
nor U15359 (N_15359,N_14097,N_14562);
nor U15360 (N_15360,N_14933,N_14714);
and U15361 (N_15361,N_14086,N_14033);
nand U15362 (N_15362,N_14841,N_14863);
nand U15363 (N_15363,N_14879,N_14733);
and U15364 (N_15364,N_14397,N_14393);
nor U15365 (N_15365,N_14213,N_14039);
or U15366 (N_15366,N_14886,N_14486);
or U15367 (N_15367,N_14180,N_14152);
or U15368 (N_15368,N_14124,N_14311);
nand U15369 (N_15369,N_14594,N_14299);
nor U15370 (N_15370,N_14541,N_14458);
xor U15371 (N_15371,N_14572,N_14946);
or U15372 (N_15372,N_14647,N_14049);
nor U15373 (N_15373,N_14237,N_14641);
nand U15374 (N_15374,N_14654,N_14121);
and U15375 (N_15375,N_14465,N_14000);
and U15376 (N_15376,N_14590,N_14051);
nor U15377 (N_15377,N_14368,N_14462);
xor U15378 (N_15378,N_14659,N_14442);
xnor U15379 (N_15379,N_14027,N_14516);
xor U15380 (N_15380,N_14380,N_14812);
or U15381 (N_15381,N_14765,N_14993);
nand U15382 (N_15382,N_14201,N_14140);
xnor U15383 (N_15383,N_14147,N_14483);
and U15384 (N_15384,N_14941,N_14041);
and U15385 (N_15385,N_14558,N_14069);
nor U15386 (N_15386,N_14354,N_14474);
nand U15387 (N_15387,N_14112,N_14912);
or U15388 (N_15388,N_14810,N_14786);
or U15389 (N_15389,N_14616,N_14809);
or U15390 (N_15390,N_14977,N_14221);
or U15391 (N_15391,N_14806,N_14251);
nor U15392 (N_15392,N_14655,N_14559);
and U15393 (N_15393,N_14200,N_14170);
xnor U15394 (N_15394,N_14128,N_14425);
nand U15395 (N_15395,N_14607,N_14293);
xnor U15396 (N_15396,N_14100,N_14792);
or U15397 (N_15397,N_14497,N_14743);
xor U15398 (N_15398,N_14334,N_14916);
nor U15399 (N_15399,N_14028,N_14999);
and U15400 (N_15400,N_14953,N_14371);
nor U15401 (N_15401,N_14472,N_14145);
xor U15402 (N_15402,N_14165,N_14869);
and U15403 (N_15403,N_14358,N_14002);
nand U15404 (N_15404,N_14814,N_14591);
or U15405 (N_15405,N_14942,N_14596);
or U15406 (N_15406,N_14703,N_14464);
or U15407 (N_15407,N_14602,N_14859);
xnor U15408 (N_15408,N_14823,N_14604);
xor U15409 (N_15409,N_14343,N_14995);
nand U15410 (N_15410,N_14803,N_14554);
xor U15411 (N_15411,N_14008,N_14302);
or U15412 (N_15412,N_14551,N_14797);
and U15413 (N_15413,N_14891,N_14658);
xor U15414 (N_15414,N_14740,N_14531);
xor U15415 (N_15415,N_14154,N_14898);
xnor U15416 (N_15416,N_14549,N_14239);
nand U15417 (N_15417,N_14096,N_14399);
xnor U15418 (N_15418,N_14001,N_14123);
nand U15419 (N_15419,N_14577,N_14906);
and U15420 (N_15420,N_14963,N_14601);
xnor U15421 (N_15421,N_14297,N_14104);
nand U15422 (N_15422,N_14951,N_14166);
nand U15423 (N_15423,N_14529,N_14447);
or U15424 (N_15424,N_14791,N_14790);
or U15425 (N_15425,N_14903,N_14700);
or U15426 (N_15426,N_14997,N_14557);
nor U15427 (N_15427,N_14626,N_14961);
or U15428 (N_15428,N_14515,N_14209);
and U15429 (N_15429,N_14838,N_14574);
or U15430 (N_15430,N_14077,N_14101);
nor U15431 (N_15431,N_14328,N_14973);
nor U15432 (N_15432,N_14188,N_14612);
and U15433 (N_15433,N_14477,N_14342);
nand U15434 (N_15434,N_14499,N_14875);
or U15435 (N_15435,N_14845,N_14175);
xor U15436 (N_15436,N_14217,N_14637);
xnor U15437 (N_15437,N_14445,N_14450);
nor U15438 (N_15438,N_14460,N_14922);
or U15439 (N_15439,N_14255,N_14363);
nor U15440 (N_15440,N_14498,N_14753);
xor U15441 (N_15441,N_14084,N_14236);
xnor U15442 (N_15442,N_14306,N_14335);
nor U15443 (N_15443,N_14479,N_14511);
nand U15444 (N_15444,N_14370,N_14005);
nor U15445 (N_15445,N_14552,N_14982);
nor U15446 (N_15446,N_14832,N_14312);
nor U15447 (N_15447,N_14116,N_14506);
and U15448 (N_15448,N_14391,N_14936);
nand U15449 (N_15449,N_14148,N_14173);
or U15450 (N_15450,N_14271,N_14038);
xor U15451 (N_15451,N_14793,N_14726);
nor U15452 (N_15452,N_14605,N_14718);
nand U15453 (N_15453,N_14060,N_14157);
xnor U15454 (N_15454,N_14469,N_14036);
or U15455 (N_15455,N_14802,N_14850);
and U15456 (N_15456,N_14913,N_14169);
or U15457 (N_15457,N_14749,N_14578);
nand U15458 (N_15458,N_14762,N_14403);
nand U15459 (N_15459,N_14987,N_14214);
nand U15460 (N_15460,N_14842,N_14750);
nand U15461 (N_15461,N_14937,N_14807);
nor U15462 (N_15462,N_14672,N_14813);
and U15463 (N_15463,N_14686,N_14890);
nand U15464 (N_15464,N_14275,N_14581);
nor U15465 (N_15465,N_14537,N_14475);
xor U15466 (N_15466,N_14073,N_14512);
nand U15467 (N_15467,N_14052,N_14336);
nand U15468 (N_15468,N_14003,N_14699);
xnor U15469 (N_15469,N_14223,N_14710);
nand U15470 (N_15470,N_14375,N_14795);
or U15471 (N_15471,N_14952,N_14043);
nand U15472 (N_15472,N_14514,N_14153);
and U15473 (N_15473,N_14962,N_14427);
nand U15474 (N_15474,N_14466,N_14756);
or U15475 (N_15475,N_14257,N_14682);
and U15476 (N_15476,N_14320,N_14252);
nand U15477 (N_15477,N_14068,N_14776);
nand U15478 (N_15478,N_14102,N_14598);
nand U15479 (N_15479,N_14540,N_14163);
or U15480 (N_15480,N_14419,N_14728);
nand U15481 (N_15481,N_14930,N_14532);
and U15482 (N_15482,N_14679,N_14386);
nand U15483 (N_15483,N_14448,N_14796);
and U15484 (N_15484,N_14737,N_14926);
or U15485 (N_15485,N_14988,N_14422);
nor U15486 (N_15486,N_14019,N_14870);
nor U15487 (N_15487,N_14677,N_14289);
or U15488 (N_15488,N_14671,N_14720);
and U15489 (N_15489,N_14172,N_14230);
nand U15490 (N_15490,N_14592,N_14777);
xor U15491 (N_15491,N_14265,N_14694);
xnor U15492 (N_15492,N_14816,N_14135);
or U15493 (N_15493,N_14744,N_14691);
nor U15494 (N_15494,N_14324,N_14144);
nand U15495 (N_15495,N_14177,N_14181);
xnor U15496 (N_15496,N_14580,N_14763);
and U15497 (N_15497,N_14113,N_14269);
xor U15498 (N_15498,N_14780,N_14502);
xor U15499 (N_15499,N_14337,N_14668);
nor U15500 (N_15500,N_14865,N_14493);
nand U15501 (N_15501,N_14136,N_14421);
and U15502 (N_15502,N_14317,N_14786);
and U15503 (N_15503,N_14144,N_14189);
or U15504 (N_15504,N_14842,N_14608);
nor U15505 (N_15505,N_14306,N_14766);
and U15506 (N_15506,N_14575,N_14432);
and U15507 (N_15507,N_14477,N_14617);
nor U15508 (N_15508,N_14022,N_14600);
xnor U15509 (N_15509,N_14401,N_14532);
or U15510 (N_15510,N_14541,N_14123);
or U15511 (N_15511,N_14000,N_14061);
and U15512 (N_15512,N_14094,N_14500);
nor U15513 (N_15513,N_14494,N_14432);
or U15514 (N_15514,N_14773,N_14511);
or U15515 (N_15515,N_14996,N_14915);
xor U15516 (N_15516,N_14783,N_14713);
xor U15517 (N_15517,N_14362,N_14067);
or U15518 (N_15518,N_14967,N_14056);
xor U15519 (N_15519,N_14193,N_14900);
or U15520 (N_15520,N_14293,N_14355);
or U15521 (N_15521,N_14898,N_14454);
nand U15522 (N_15522,N_14225,N_14135);
nand U15523 (N_15523,N_14887,N_14172);
nor U15524 (N_15524,N_14440,N_14613);
nor U15525 (N_15525,N_14045,N_14300);
and U15526 (N_15526,N_14788,N_14240);
xor U15527 (N_15527,N_14734,N_14022);
and U15528 (N_15528,N_14873,N_14497);
nand U15529 (N_15529,N_14110,N_14838);
xor U15530 (N_15530,N_14808,N_14412);
and U15531 (N_15531,N_14701,N_14554);
and U15532 (N_15532,N_14265,N_14448);
or U15533 (N_15533,N_14147,N_14839);
or U15534 (N_15534,N_14446,N_14684);
nor U15535 (N_15535,N_14894,N_14812);
and U15536 (N_15536,N_14730,N_14403);
or U15537 (N_15537,N_14088,N_14713);
or U15538 (N_15538,N_14969,N_14698);
or U15539 (N_15539,N_14755,N_14186);
nand U15540 (N_15540,N_14672,N_14278);
nor U15541 (N_15541,N_14565,N_14699);
xor U15542 (N_15542,N_14593,N_14667);
and U15543 (N_15543,N_14023,N_14984);
or U15544 (N_15544,N_14144,N_14227);
and U15545 (N_15545,N_14529,N_14389);
and U15546 (N_15546,N_14041,N_14734);
xnor U15547 (N_15547,N_14937,N_14825);
or U15548 (N_15548,N_14988,N_14341);
or U15549 (N_15549,N_14162,N_14443);
and U15550 (N_15550,N_14720,N_14475);
or U15551 (N_15551,N_14422,N_14935);
or U15552 (N_15552,N_14991,N_14267);
nand U15553 (N_15553,N_14953,N_14470);
nor U15554 (N_15554,N_14692,N_14533);
or U15555 (N_15555,N_14710,N_14381);
or U15556 (N_15556,N_14855,N_14349);
and U15557 (N_15557,N_14821,N_14086);
or U15558 (N_15558,N_14903,N_14062);
nand U15559 (N_15559,N_14732,N_14304);
or U15560 (N_15560,N_14547,N_14908);
nor U15561 (N_15561,N_14575,N_14095);
xnor U15562 (N_15562,N_14015,N_14695);
xor U15563 (N_15563,N_14805,N_14199);
nand U15564 (N_15564,N_14184,N_14480);
and U15565 (N_15565,N_14827,N_14274);
nand U15566 (N_15566,N_14219,N_14737);
nor U15567 (N_15567,N_14694,N_14564);
or U15568 (N_15568,N_14318,N_14509);
nand U15569 (N_15569,N_14889,N_14585);
and U15570 (N_15570,N_14279,N_14886);
xor U15571 (N_15571,N_14348,N_14297);
or U15572 (N_15572,N_14701,N_14533);
xnor U15573 (N_15573,N_14094,N_14590);
nor U15574 (N_15574,N_14662,N_14563);
nand U15575 (N_15575,N_14963,N_14533);
or U15576 (N_15576,N_14366,N_14689);
or U15577 (N_15577,N_14926,N_14388);
nor U15578 (N_15578,N_14416,N_14803);
nor U15579 (N_15579,N_14418,N_14151);
nor U15580 (N_15580,N_14521,N_14458);
xor U15581 (N_15581,N_14083,N_14393);
xnor U15582 (N_15582,N_14208,N_14989);
nand U15583 (N_15583,N_14398,N_14137);
and U15584 (N_15584,N_14301,N_14437);
or U15585 (N_15585,N_14605,N_14210);
nor U15586 (N_15586,N_14681,N_14460);
xnor U15587 (N_15587,N_14592,N_14486);
and U15588 (N_15588,N_14656,N_14680);
nand U15589 (N_15589,N_14906,N_14161);
nand U15590 (N_15590,N_14362,N_14883);
nor U15591 (N_15591,N_14614,N_14732);
xnor U15592 (N_15592,N_14997,N_14765);
and U15593 (N_15593,N_14311,N_14848);
and U15594 (N_15594,N_14129,N_14716);
nor U15595 (N_15595,N_14010,N_14461);
and U15596 (N_15596,N_14308,N_14516);
xor U15597 (N_15597,N_14952,N_14411);
and U15598 (N_15598,N_14548,N_14783);
xnor U15599 (N_15599,N_14816,N_14275);
nand U15600 (N_15600,N_14131,N_14763);
nor U15601 (N_15601,N_14408,N_14333);
nor U15602 (N_15602,N_14652,N_14857);
xor U15603 (N_15603,N_14725,N_14433);
nand U15604 (N_15604,N_14806,N_14156);
xnor U15605 (N_15605,N_14265,N_14732);
xnor U15606 (N_15606,N_14260,N_14696);
nor U15607 (N_15607,N_14354,N_14546);
nand U15608 (N_15608,N_14027,N_14802);
or U15609 (N_15609,N_14817,N_14147);
xor U15610 (N_15610,N_14325,N_14738);
and U15611 (N_15611,N_14522,N_14193);
xnor U15612 (N_15612,N_14049,N_14752);
nand U15613 (N_15613,N_14944,N_14306);
xor U15614 (N_15614,N_14291,N_14430);
nand U15615 (N_15615,N_14013,N_14296);
nand U15616 (N_15616,N_14065,N_14721);
nand U15617 (N_15617,N_14874,N_14421);
or U15618 (N_15618,N_14680,N_14544);
nand U15619 (N_15619,N_14643,N_14734);
and U15620 (N_15620,N_14350,N_14815);
or U15621 (N_15621,N_14856,N_14750);
and U15622 (N_15622,N_14276,N_14178);
xnor U15623 (N_15623,N_14889,N_14336);
xor U15624 (N_15624,N_14830,N_14183);
or U15625 (N_15625,N_14287,N_14908);
nand U15626 (N_15626,N_14279,N_14636);
xor U15627 (N_15627,N_14185,N_14117);
or U15628 (N_15628,N_14182,N_14464);
and U15629 (N_15629,N_14531,N_14010);
or U15630 (N_15630,N_14625,N_14545);
nor U15631 (N_15631,N_14135,N_14859);
nor U15632 (N_15632,N_14592,N_14643);
nor U15633 (N_15633,N_14777,N_14047);
nand U15634 (N_15634,N_14854,N_14163);
nand U15635 (N_15635,N_14617,N_14221);
xor U15636 (N_15636,N_14936,N_14698);
nor U15637 (N_15637,N_14146,N_14217);
nor U15638 (N_15638,N_14753,N_14078);
nor U15639 (N_15639,N_14634,N_14880);
nand U15640 (N_15640,N_14711,N_14415);
nor U15641 (N_15641,N_14119,N_14003);
nand U15642 (N_15642,N_14416,N_14895);
and U15643 (N_15643,N_14650,N_14533);
and U15644 (N_15644,N_14701,N_14328);
xor U15645 (N_15645,N_14716,N_14873);
or U15646 (N_15646,N_14410,N_14598);
xor U15647 (N_15647,N_14581,N_14267);
nand U15648 (N_15648,N_14494,N_14230);
xnor U15649 (N_15649,N_14177,N_14391);
xnor U15650 (N_15650,N_14990,N_14583);
xnor U15651 (N_15651,N_14274,N_14070);
and U15652 (N_15652,N_14277,N_14756);
xor U15653 (N_15653,N_14101,N_14045);
nand U15654 (N_15654,N_14152,N_14319);
nor U15655 (N_15655,N_14187,N_14439);
nor U15656 (N_15656,N_14763,N_14628);
or U15657 (N_15657,N_14538,N_14371);
and U15658 (N_15658,N_14839,N_14044);
and U15659 (N_15659,N_14037,N_14939);
xor U15660 (N_15660,N_14198,N_14699);
and U15661 (N_15661,N_14053,N_14542);
or U15662 (N_15662,N_14583,N_14958);
nand U15663 (N_15663,N_14561,N_14814);
and U15664 (N_15664,N_14676,N_14176);
nand U15665 (N_15665,N_14402,N_14971);
xor U15666 (N_15666,N_14006,N_14002);
and U15667 (N_15667,N_14418,N_14282);
nor U15668 (N_15668,N_14935,N_14086);
or U15669 (N_15669,N_14901,N_14710);
xor U15670 (N_15670,N_14589,N_14580);
nand U15671 (N_15671,N_14837,N_14285);
and U15672 (N_15672,N_14822,N_14739);
or U15673 (N_15673,N_14085,N_14902);
nor U15674 (N_15674,N_14340,N_14119);
nor U15675 (N_15675,N_14144,N_14558);
xnor U15676 (N_15676,N_14192,N_14793);
or U15677 (N_15677,N_14678,N_14196);
nand U15678 (N_15678,N_14688,N_14087);
nand U15679 (N_15679,N_14004,N_14507);
nand U15680 (N_15680,N_14788,N_14277);
and U15681 (N_15681,N_14011,N_14493);
nor U15682 (N_15682,N_14843,N_14188);
and U15683 (N_15683,N_14873,N_14485);
nand U15684 (N_15684,N_14978,N_14697);
or U15685 (N_15685,N_14732,N_14030);
xnor U15686 (N_15686,N_14747,N_14830);
and U15687 (N_15687,N_14264,N_14585);
nor U15688 (N_15688,N_14963,N_14423);
and U15689 (N_15689,N_14449,N_14036);
and U15690 (N_15690,N_14109,N_14296);
or U15691 (N_15691,N_14470,N_14619);
or U15692 (N_15692,N_14085,N_14417);
nand U15693 (N_15693,N_14451,N_14678);
nand U15694 (N_15694,N_14361,N_14291);
nand U15695 (N_15695,N_14460,N_14002);
nand U15696 (N_15696,N_14472,N_14877);
xor U15697 (N_15697,N_14347,N_14175);
xor U15698 (N_15698,N_14418,N_14504);
nand U15699 (N_15699,N_14128,N_14846);
and U15700 (N_15700,N_14130,N_14418);
nor U15701 (N_15701,N_14309,N_14640);
nand U15702 (N_15702,N_14528,N_14958);
and U15703 (N_15703,N_14997,N_14333);
nor U15704 (N_15704,N_14674,N_14418);
and U15705 (N_15705,N_14436,N_14662);
or U15706 (N_15706,N_14121,N_14186);
nand U15707 (N_15707,N_14890,N_14043);
xnor U15708 (N_15708,N_14650,N_14112);
nand U15709 (N_15709,N_14751,N_14148);
or U15710 (N_15710,N_14896,N_14529);
or U15711 (N_15711,N_14800,N_14008);
xnor U15712 (N_15712,N_14580,N_14460);
nor U15713 (N_15713,N_14933,N_14902);
nand U15714 (N_15714,N_14239,N_14413);
nor U15715 (N_15715,N_14915,N_14016);
or U15716 (N_15716,N_14563,N_14719);
nor U15717 (N_15717,N_14567,N_14408);
or U15718 (N_15718,N_14898,N_14726);
nand U15719 (N_15719,N_14359,N_14124);
or U15720 (N_15720,N_14165,N_14769);
or U15721 (N_15721,N_14788,N_14251);
nand U15722 (N_15722,N_14057,N_14274);
xnor U15723 (N_15723,N_14740,N_14092);
nand U15724 (N_15724,N_14672,N_14340);
and U15725 (N_15725,N_14716,N_14742);
nor U15726 (N_15726,N_14214,N_14061);
nand U15727 (N_15727,N_14373,N_14554);
or U15728 (N_15728,N_14310,N_14182);
nand U15729 (N_15729,N_14655,N_14671);
xnor U15730 (N_15730,N_14745,N_14982);
or U15731 (N_15731,N_14728,N_14624);
or U15732 (N_15732,N_14137,N_14958);
and U15733 (N_15733,N_14365,N_14385);
nand U15734 (N_15734,N_14165,N_14172);
nand U15735 (N_15735,N_14673,N_14077);
nor U15736 (N_15736,N_14177,N_14293);
and U15737 (N_15737,N_14759,N_14312);
xor U15738 (N_15738,N_14675,N_14545);
nor U15739 (N_15739,N_14153,N_14201);
nor U15740 (N_15740,N_14323,N_14166);
and U15741 (N_15741,N_14998,N_14408);
nor U15742 (N_15742,N_14052,N_14647);
nand U15743 (N_15743,N_14433,N_14564);
xnor U15744 (N_15744,N_14104,N_14453);
xnor U15745 (N_15745,N_14789,N_14772);
and U15746 (N_15746,N_14340,N_14966);
nand U15747 (N_15747,N_14752,N_14711);
or U15748 (N_15748,N_14721,N_14062);
or U15749 (N_15749,N_14712,N_14761);
nand U15750 (N_15750,N_14170,N_14411);
nor U15751 (N_15751,N_14443,N_14247);
xnor U15752 (N_15752,N_14583,N_14722);
or U15753 (N_15753,N_14491,N_14089);
and U15754 (N_15754,N_14247,N_14128);
or U15755 (N_15755,N_14485,N_14998);
xor U15756 (N_15756,N_14838,N_14964);
and U15757 (N_15757,N_14487,N_14081);
nor U15758 (N_15758,N_14077,N_14300);
and U15759 (N_15759,N_14805,N_14367);
xor U15760 (N_15760,N_14812,N_14743);
and U15761 (N_15761,N_14967,N_14196);
and U15762 (N_15762,N_14485,N_14770);
nand U15763 (N_15763,N_14748,N_14560);
or U15764 (N_15764,N_14362,N_14438);
or U15765 (N_15765,N_14802,N_14693);
or U15766 (N_15766,N_14121,N_14015);
xor U15767 (N_15767,N_14227,N_14624);
nor U15768 (N_15768,N_14743,N_14031);
nor U15769 (N_15769,N_14455,N_14787);
or U15770 (N_15770,N_14552,N_14535);
nand U15771 (N_15771,N_14404,N_14534);
xor U15772 (N_15772,N_14657,N_14019);
xor U15773 (N_15773,N_14375,N_14431);
nand U15774 (N_15774,N_14003,N_14260);
and U15775 (N_15775,N_14047,N_14483);
nor U15776 (N_15776,N_14043,N_14963);
nand U15777 (N_15777,N_14948,N_14536);
nor U15778 (N_15778,N_14847,N_14082);
xor U15779 (N_15779,N_14826,N_14919);
and U15780 (N_15780,N_14953,N_14860);
nand U15781 (N_15781,N_14900,N_14930);
and U15782 (N_15782,N_14765,N_14688);
xor U15783 (N_15783,N_14769,N_14887);
nand U15784 (N_15784,N_14546,N_14846);
or U15785 (N_15785,N_14437,N_14093);
nor U15786 (N_15786,N_14180,N_14996);
and U15787 (N_15787,N_14781,N_14247);
and U15788 (N_15788,N_14822,N_14977);
nor U15789 (N_15789,N_14689,N_14164);
and U15790 (N_15790,N_14544,N_14397);
xor U15791 (N_15791,N_14634,N_14078);
or U15792 (N_15792,N_14914,N_14169);
and U15793 (N_15793,N_14476,N_14044);
nor U15794 (N_15794,N_14031,N_14322);
and U15795 (N_15795,N_14513,N_14667);
xor U15796 (N_15796,N_14307,N_14141);
or U15797 (N_15797,N_14104,N_14671);
nand U15798 (N_15798,N_14089,N_14516);
nand U15799 (N_15799,N_14562,N_14960);
and U15800 (N_15800,N_14382,N_14049);
or U15801 (N_15801,N_14517,N_14535);
xnor U15802 (N_15802,N_14544,N_14101);
nand U15803 (N_15803,N_14604,N_14927);
nor U15804 (N_15804,N_14634,N_14330);
xor U15805 (N_15805,N_14619,N_14453);
xnor U15806 (N_15806,N_14139,N_14274);
and U15807 (N_15807,N_14396,N_14020);
nand U15808 (N_15808,N_14240,N_14821);
and U15809 (N_15809,N_14467,N_14522);
xor U15810 (N_15810,N_14672,N_14257);
or U15811 (N_15811,N_14386,N_14450);
xor U15812 (N_15812,N_14006,N_14926);
nand U15813 (N_15813,N_14280,N_14780);
nand U15814 (N_15814,N_14996,N_14463);
or U15815 (N_15815,N_14827,N_14263);
and U15816 (N_15816,N_14315,N_14147);
nand U15817 (N_15817,N_14216,N_14528);
and U15818 (N_15818,N_14660,N_14970);
xor U15819 (N_15819,N_14365,N_14474);
nor U15820 (N_15820,N_14890,N_14433);
nor U15821 (N_15821,N_14189,N_14486);
or U15822 (N_15822,N_14501,N_14667);
nand U15823 (N_15823,N_14695,N_14574);
xor U15824 (N_15824,N_14402,N_14227);
xor U15825 (N_15825,N_14455,N_14424);
or U15826 (N_15826,N_14753,N_14760);
xor U15827 (N_15827,N_14168,N_14505);
xnor U15828 (N_15828,N_14683,N_14754);
or U15829 (N_15829,N_14024,N_14379);
and U15830 (N_15830,N_14869,N_14660);
and U15831 (N_15831,N_14269,N_14080);
xor U15832 (N_15832,N_14082,N_14372);
and U15833 (N_15833,N_14528,N_14646);
or U15834 (N_15834,N_14030,N_14343);
xor U15835 (N_15835,N_14882,N_14859);
nand U15836 (N_15836,N_14602,N_14352);
nand U15837 (N_15837,N_14759,N_14175);
nand U15838 (N_15838,N_14641,N_14291);
nand U15839 (N_15839,N_14601,N_14418);
nand U15840 (N_15840,N_14409,N_14731);
or U15841 (N_15841,N_14469,N_14638);
and U15842 (N_15842,N_14932,N_14592);
and U15843 (N_15843,N_14885,N_14175);
nor U15844 (N_15844,N_14617,N_14062);
nand U15845 (N_15845,N_14656,N_14920);
or U15846 (N_15846,N_14970,N_14275);
or U15847 (N_15847,N_14740,N_14640);
xnor U15848 (N_15848,N_14547,N_14340);
or U15849 (N_15849,N_14999,N_14830);
nand U15850 (N_15850,N_14153,N_14801);
xor U15851 (N_15851,N_14048,N_14139);
xnor U15852 (N_15852,N_14222,N_14295);
xnor U15853 (N_15853,N_14254,N_14584);
xor U15854 (N_15854,N_14713,N_14920);
xnor U15855 (N_15855,N_14670,N_14240);
xnor U15856 (N_15856,N_14917,N_14592);
or U15857 (N_15857,N_14243,N_14008);
nand U15858 (N_15858,N_14729,N_14404);
and U15859 (N_15859,N_14037,N_14259);
nand U15860 (N_15860,N_14329,N_14164);
nor U15861 (N_15861,N_14235,N_14611);
and U15862 (N_15862,N_14543,N_14010);
xnor U15863 (N_15863,N_14700,N_14103);
and U15864 (N_15864,N_14259,N_14385);
nor U15865 (N_15865,N_14213,N_14284);
xor U15866 (N_15866,N_14610,N_14186);
nor U15867 (N_15867,N_14934,N_14369);
or U15868 (N_15868,N_14549,N_14427);
or U15869 (N_15869,N_14421,N_14891);
and U15870 (N_15870,N_14156,N_14787);
and U15871 (N_15871,N_14919,N_14219);
nor U15872 (N_15872,N_14327,N_14464);
nand U15873 (N_15873,N_14283,N_14770);
nor U15874 (N_15874,N_14372,N_14527);
xor U15875 (N_15875,N_14510,N_14560);
and U15876 (N_15876,N_14138,N_14096);
or U15877 (N_15877,N_14946,N_14154);
and U15878 (N_15878,N_14766,N_14554);
or U15879 (N_15879,N_14201,N_14749);
nor U15880 (N_15880,N_14862,N_14282);
xor U15881 (N_15881,N_14161,N_14037);
and U15882 (N_15882,N_14510,N_14024);
nor U15883 (N_15883,N_14890,N_14839);
nor U15884 (N_15884,N_14815,N_14582);
xnor U15885 (N_15885,N_14539,N_14573);
nor U15886 (N_15886,N_14518,N_14576);
or U15887 (N_15887,N_14980,N_14795);
nor U15888 (N_15888,N_14930,N_14444);
or U15889 (N_15889,N_14903,N_14570);
nand U15890 (N_15890,N_14078,N_14858);
xor U15891 (N_15891,N_14218,N_14908);
or U15892 (N_15892,N_14477,N_14167);
nor U15893 (N_15893,N_14720,N_14140);
or U15894 (N_15894,N_14219,N_14521);
and U15895 (N_15895,N_14465,N_14827);
xnor U15896 (N_15896,N_14272,N_14881);
nor U15897 (N_15897,N_14878,N_14260);
nand U15898 (N_15898,N_14762,N_14624);
or U15899 (N_15899,N_14191,N_14637);
or U15900 (N_15900,N_14874,N_14541);
and U15901 (N_15901,N_14366,N_14977);
nor U15902 (N_15902,N_14374,N_14089);
xor U15903 (N_15903,N_14007,N_14590);
or U15904 (N_15904,N_14847,N_14130);
or U15905 (N_15905,N_14678,N_14181);
xnor U15906 (N_15906,N_14486,N_14029);
and U15907 (N_15907,N_14048,N_14229);
or U15908 (N_15908,N_14557,N_14625);
and U15909 (N_15909,N_14265,N_14045);
nand U15910 (N_15910,N_14626,N_14342);
or U15911 (N_15911,N_14581,N_14098);
and U15912 (N_15912,N_14488,N_14212);
nor U15913 (N_15913,N_14128,N_14111);
or U15914 (N_15914,N_14766,N_14365);
or U15915 (N_15915,N_14117,N_14340);
and U15916 (N_15916,N_14558,N_14445);
or U15917 (N_15917,N_14196,N_14549);
nand U15918 (N_15918,N_14136,N_14652);
or U15919 (N_15919,N_14716,N_14195);
or U15920 (N_15920,N_14267,N_14910);
and U15921 (N_15921,N_14273,N_14630);
xnor U15922 (N_15922,N_14461,N_14650);
nor U15923 (N_15923,N_14538,N_14030);
nand U15924 (N_15924,N_14616,N_14512);
nor U15925 (N_15925,N_14495,N_14538);
and U15926 (N_15926,N_14185,N_14112);
nor U15927 (N_15927,N_14963,N_14119);
or U15928 (N_15928,N_14100,N_14074);
and U15929 (N_15929,N_14394,N_14097);
or U15930 (N_15930,N_14932,N_14322);
nand U15931 (N_15931,N_14198,N_14271);
or U15932 (N_15932,N_14836,N_14069);
and U15933 (N_15933,N_14560,N_14283);
and U15934 (N_15934,N_14412,N_14536);
and U15935 (N_15935,N_14116,N_14524);
nand U15936 (N_15936,N_14233,N_14869);
nand U15937 (N_15937,N_14165,N_14545);
or U15938 (N_15938,N_14672,N_14784);
xnor U15939 (N_15939,N_14065,N_14470);
nor U15940 (N_15940,N_14203,N_14973);
xnor U15941 (N_15941,N_14082,N_14040);
or U15942 (N_15942,N_14348,N_14868);
nand U15943 (N_15943,N_14594,N_14679);
nand U15944 (N_15944,N_14448,N_14318);
or U15945 (N_15945,N_14654,N_14013);
xor U15946 (N_15946,N_14691,N_14137);
and U15947 (N_15947,N_14106,N_14929);
nor U15948 (N_15948,N_14310,N_14200);
xor U15949 (N_15949,N_14486,N_14259);
and U15950 (N_15950,N_14557,N_14363);
nor U15951 (N_15951,N_14948,N_14865);
or U15952 (N_15952,N_14740,N_14938);
nor U15953 (N_15953,N_14278,N_14087);
xnor U15954 (N_15954,N_14511,N_14695);
nor U15955 (N_15955,N_14385,N_14419);
xnor U15956 (N_15956,N_14587,N_14244);
xor U15957 (N_15957,N_14040,N_14341);
or U15958 (N_15958,N_14343,N_14582);
nand U15959 (N_15959,N_14367,N_14868);
nand U15960 (N_15960,N_14739,N_14512);
xor U15961 (N_15961,N_14784,N_14065);
xnor U15962 (N_15962,N_14561,N_14205);
nor U15963 (N_15963,N_14659,N_14931);
and U15964 (N_15964,N_14706,N_14810);
nor U15965 (N_15965,N_14717,N_14699);
nand U15966 (N_15966,N_14569,N_14742);
xor U15967 (N_15967,N_14436,N_14265);
nand U15968 (N_15968,N_14054,N_14631);
nand U15969 (N_15969,N_14641,N_14487);
and U15970 (N_15970,N_14824,N_14151);
nand U15971 (N_15971,N_14704,N_14084);
nand U15972 (N_15972,N_14248,N_14352);
xor U15973 (N_15973,N_14157,N_14993);
nor U15974 (N_15974,N_14234,N_14119);
xor U15975 (N_15975,N_14522,N_14254);
or U15976 (N_15976,N_14830,N_14323);
nor U15977 (N_15977,N_14463,N_14263);
or U15978 (N_15978,N_14790,N_14280);
xor U15979 (N_15979,N_14182,N_14846);
or U15980 (N_15980,N_14110,N_14142);
or U15981 (N_15981,N_14645,N_14824);
or U15982 (N_15982,N_14294,N_14095);
nor U15983 (N_15983,N_14556,N_14827);
nand U15984 (N_15984,N_14991,N_14904);
or U15985 (N_15985,N_14783,N_14810);
or U15986 (N_15986,N_14851,N_14020);
nand U15987 (N_15987,N_14008,N_14664);
nand U15988 (N_15988,N_14050,N_14788);
xnor U15989 (N_15989,N_14463,N_14737);
and U15990 (N_15990,N_14332,N_14213);
nand U15991 (N_15991,N_14794,N_14150);
or U15992 (N_15992,N_14244,N_14187);
nor U15993 (N_15993,N_14123,N_14749);
xnor U15994 (N_15994,N_14673,N_14021);
and U15995 (N_15995,N_14048,N_14266);
and U15996 (N_15996,N_14543,N_14604);
and U15997 (N_15997,N_14990,N_14955);
nor U15998 (N_15998,N_14532,N_14250);
and U15999 (N_15999,N_14691,N_14347);
nand U16000 (N_16000,N_15151,N_15577);
xor U16001 (N_16001,N_15351,N_15024);
and U16002 (N_16002,N_15877,N_15342);
or U16003 (N_16003,N_15242,N_15600);
xnor U16004 (N_16004,N_15887,N_15703);
or U16005 (N_16005,N_15038,N_15779);
and U16006 (N_16006,N_15130,N_15996);
or U16007 (N_16007,N_15604,N_15840);
nand U16008 (N_16008,N_15168,N_15911);
nor U16009 (N_16009,N_15700,N_15311);
and U16010 (N_16010,N_15166,N_15689);
and U16011 (N_16011,N_15948,N_15743);
nand U16012 (N_16012,N_15012,N_15320);
and U16013 (N_16013,N_15581,N_15451);
or U16014 (N_16014,N_15216,N_15832);
xor U16015 (N_16015,N_15898,N_15464);
nor U16016 (N_16016,N_15715,N_15650);
nand U16017 (N_16017,N_15393,N_15000);
nor U16018 (N_16018,N_15082,N_15558);
xor U16019 (N_16019,N_15058,N_15034);
or U16020 (N_16020,N_15666,N_15125);
xnor U16021 (N_16021,N_15248,N_15892);
xor U16022 (N_16022,N_15052,N_15008);
xnor U16023 (N_16023,N_15372,N_15035);
xnor U16024 (N_16024,N_15375,N_15423);
xnor U16025 (N_16025,N_15701,N_15730);
nand U16026 (N_16026,N_15014,N_15200);
nand U16027 (N_16027,N_15308,N_15591);
xor U16028 (N_16028,N_15925,N_15993);
xnor U16029 (N_16029,N_15210,N_15835);
nor U16030 (N_16030,N_15607,N_15603);
nor U16031 (N_16031,N_15405,N_15146);
nor U16032 (N_16032,N_15473,N_15940);
xnor U16033 (N_16033,N_15520,N_15163);
xnor U16034 (N_16034,N_15127,N_15916);
and U16035 (N_16035,N_15465,N_15447);
and U16036 (N_16036,N_15837,N_15851);
nor U16037 (N_16037,N_15425,N_15212);
nand U16038 (N_16038,N_15893,N_15376);
xor U16039 (N_16039,N_15852,N_15463);
xor U16040 (N_16040,N_15139,N_15866);
nor U16041 (N_16041,N_15816,N_15858);
nand U16042 (N_16042,N_15628,N_15224);
nand U16043 (N_16043,N_15665,N_15062);
nor U16044 (N_16044,N_15512,N_15098);
nor U16045 (N_16045,N_15566,N_15957);
xor U16046 (N_16046,N_15740,N_15292);
or U16047 (N_16047,N_15551,N_15099);
nand U16048 (N_16048,N_15506,N_15507);
or U16049 (N_16049,N_15361,N_15050);
or U16050 (N_16050,N_15266,N_15394);
xnor U16051 (N_16051,N_15992,N_15455);
or U16052 (N_16052,N_15335,N_15379);
nand U16053 (N_16053,N_15717,N_15928);
or U16054 (N_16054,N_15259,N_15720);
or U16055 (N_16055,N_15129,N_15088);
or U16056 (N_16056,N_15980,N_15849);
nor U16057 (N_16057,N_15587,N_15675);
or U16058 (N_16058,N_15913,N_15883);
nor U16059 (N_16059,N_15422,N_15286);
nand U16060 (N_16060,N_15638,N_15491);
or U16061 (N_16061,N_15757,N_15805);
nor U16062 (N_16062,N_15854,N_15170);
nand U16063 (N_16063,N_15390,N_15873);
or U16064 (N_16064,N_15252,N_15289);
and U16065 (N_16065,N_15702,N_15956);
xor U16066 (N_16066,N_15640,N_15258);
xnor U16067 (N_16067,N_15695,N_15358);
or U16068 (N_16068,N_15201,N_15440);
xor U16069 (N_16069,N_15119,N_15309);
or U16070 (N_16070,N_15525,N_15148);
nor U16071 (N_16071,N_15729,N_15909);
and U16072 (N_16072,N_15821,N_15579);
nor U16073 (N_16073,N_15350,N_15775);
xnor U16074 (N_16074,N_15841,N_15986);
and U16075 (N_16075,N_15514,N_15827);
and U16076 (N_16076,N_15784,N_15486);
and U16077 (N_16077,N_15232,N_15408);
nand U16078 (N_16078,N_15677,N_15172);
or U16079 (N_16079,N_15636,N_15132);
nor U16080 (N_16080,N_15633,N_15070);
nand U16081 (N_16081,N_15795,N_15274);
xnor U16082 (N_16082,N_15040,N_15739);
or U16083 (N_16083,N_15882,N_15509);
and U16084 (N_16084,N_15179,N_15078);
xnor U16085 (N_16085,N_15086,N_15183);
xnor U16086 (N_16086,N_15443,N_15524);
nor U16087 (N_16087,N_15287,N_15659);
and U16088 (N_16088,N_15339,N_15671);
or U16089 (N_16089,N_15206,N_15921);
nor U16090 (N_16090,N_15781,N_15806);
nor U16091 (N_16091,N_15269,N_15303);
and U16092 (N_16092,N_15084,N_15648);
and U16093 (N_16093,N_15064,N_15871);
and U16094 (N_16094,N_15714,N_15111);
and U16095 (N_16095,N_15178,N_15780);
or U16096 (N_16096,N_15977,N_15467);
xor U16097 (N_16097,N_15502,N_15409);
xnor U16098 (N_16098,N_15760,N_15985);
or U16099 (N_16099,N_15748,N_15523);
nand U16100 (N_16100,N_15769,N_15978);
and U16101 (N_16101,N_15371,N_15057);
and U16102 (N_16102,N_15173,N_15613);
xor U16103 (N_16103,N_15114,N_15138);
nor U16104 (N_16104,N_15679,N_15391);
or U16105 (N_16105,N_15112,N_15763);
or U16106 (N_16106,N_15068,N_15243);
xnor U16107 (N_16107,N_15645,N_15856);
nor U16108 (N_16108,N_15688,N_15401);
xor U16109 (N_16109,N_15534,N_15255);
or U16110 (N_16110,N_15060,N_15018);
and U16111 (N_16111,N_15133,N_15678);
or U16112 (N_16112,N_15517,N_15131);
xor U16113 (N_16113,N_15949,N_15233);
xnor U16114 (N_16114,N_15270,N_15260);
nor U16115 (N_16115,N_15942,N_15972);
nor U16116 (N_16116,N_15338,N_15975);
nand U16117 (N_16117,N_15313,N_15356);
and U16118 (N_16118,N_15554,N_15189);
nand U16119 (N_16119,N_15021,N_15096);
and U16120 (N_16120,N_15322,N_15522);
and U16121 (N_16121,N_15500,N_15295);
and U16122 (N_16122,N_15941,N_15343);
nand U16123 (N_16123,N_15113,N_15503);
or U16124 (N_16124,N_15623,N_15249);
and U16125 (N_16125,N_15672,N_15753);
xor U16126 (N_16126,N_15987,N_15478);
xor U16127 (N_16127,N_15360,N_15354);
and U16128 (N_16128,N_15939,N_15412);
or U16129 (N_16129,N_15960,N_15533);
or U16130 (N_16130,N_15271,N_15218);
nor U16131 (N_16131,N_15262,N_15175);
and U16132 (N_16132,N_15722,N_15934);
nor U16133 (N_16133,N_15818,N_15876);
xor U16134 (N_16134,N_15758,N_15999);
nand U16135 (N_16135,N_15728,N_15263);
or U16136 (N_16136,N_15707,N_15685);
xnor U16137 (N_16137,N_15899,N_15799);
or U16138 (N_16138,N_15970,N_15718);
or U16139 (N_16139,N_15469,N_15560);
and U16140 (N_16140,N_15627,N_15143);
and U16141 (N_16141,N_15006,N_15699);
nand U16142 (N_16142,N_15845,N_15615);
and U16143 (N_16143,N_15219,N_15997);
nand U16144 (N_16144,N_15823,N_15240);
xnor U16145 (N_16145,N_15275,N_15066);
and U16146 (N_16146,N_15791,N_15167);
xor U16147 (N_16147,N_15452,N_15013);
nand U16148 (N_16148,N_15919,N_15348);
xor U16149 (N_16149,N_15253,N_15680);
and U16150 (N_16150,N_15855,N_15374);
xor U16151 (N_16151,N_15436,N_15141);
and U16152 (N_16152,N_15437,N_15237);
nand U16153 (N_16153,N_15485,N_15541);
or U16154 (N_16154,N_15332,N_15302);
nor U16155 (N_16155,N_15570,N_15466);
or U16156 (N_16156,N_15184,N_15569);
nand U16157 (N_16157,N_15563,N_15345);
and U16158 (N_16158,N_15053,N_15482);
and U16159 (N_16159,N_15930,N_15629);
xnor U16160 (N_16160,N_15809,N_15367);
or U16161 (N_16161,N_15198,N_15380);
nand U16162 (N_16162,N_15429,N_15819);
or U16163 (N_16163,N_15528,N_15527);
and U16164 (N_16164,N_15634,N_15480);
or U16165 (N_16165,N_15829,N_15220);
or U16166 (N_16166,N_15272,N_15931);
or U16167 (N_16167,N_15268,N_15540);
and U16168 (N_16168,N_15370,N_15914);
nor U16169 (N_16169,N_15642,N_15384);
and U16170 (N_16170,N_15626,N_15785);
nand U16171 (N_16171,N_15697,N_15284);
nor U16172 (N_16172,N_15349,N_15029);
xnor U16173 (N_16173,N_15918,N_15649);
nand U16174 (N_16174,N_15885,N_15056);
nand U16175 (N_16175,N_15054,N_15585);
xnor U16176 (N_16176,N_15108,N_15085);
nand U16177 (N_16177,N_15160,N_15831);
nand U16178 (N_16178,N_15814,N_15202);
or U16179 (N_16179,N_15011,N_15592);
and U16180 (N_16180,N_15750,N_15860);
and U16181 (N_16181,N_15494,N_15770);
and U16182 (N_16182,N_15565,N_15761);
or U16183 (N_16183,N_15059,N_15398);
nand U16184 (N_16184,N_15105,N_15618);
nand U16185 (N_16185,N_15214,N_15142);
xnor U16186 (N_16186,N_15647,N_15044);
or U16187 (N_16187,N_15306,N_15476);
nor U16188 (N_16188,N_15435,N_15438);
and U16189 (N_16189,N_15811,N_15294);
and U16190 (N_16190,N_15842,N_15706);
nor U16191 (N_16191,N_15330,N_15955);
xor U16192 (N_16192,N_15813,N_15646);
nor U16193 (N_16193,N_15479,N_15869);
xor U16194 (N_16194,N_15225,N_15929);
nor U16195 (N_16195,N_15530,N_15602);
nand U16196 (N_16196,N_15550,N_15895);
nor U16197 (N_16197,N_15428,N_15974);
or U16198 (N_16198,N_15555,N_15280);
nor U16199 (N_16199,N_15181,N_15802);
xnor U16200 (N_16200,N_15395,N_15872);
nand U16201 (N_16201,N_15884,N_15386);
nor U16202 (N_16202,N_15709,N_15116);
nand U16203 (N_16203,N_15747,N_15484);
xor U16204 (N_16204,N_15962,N_15406);
or U16205 (N_16205,N_15559,N_15952);
and U16206 (N_16206,N_15288,N_15850);
and U16207 (N_16207,N_15036,N_15341);
nor U16208 (N_16208,N_15246,N_15783);
or U16209 (N_16209,N_15598,N_15497);
xor U16210 (N_16210,N_15643,N_15276);
and U16211 (N_16211,N_15357,N_15118);
nand U16212 (N_16212,N_15725,N_15724);
and U16213 (N_16213,N_15669,N_15595);
xnor U16214 (N_16214,N_15828,N_15065);
nor U16215 (N_16215,N_15211,N_15298);
and U16216 (N_16216,N_15947,N_15848);
xnor U16217 (N_16217,N_15089,N_15325);
nand U16218 (N_16218,N_15093,N_15710);
xnor U16219 (N_16219,N_15542,N_15983);
xnor U16220 (N_16220,N_15316,N_15387);
and U16221 (N_16221,N_15472,N_15180);
nand U16222 (N_16222,N_15005,N_15622);
and U16223 (N_16223,N_15267,N_15578);
xnor U16224 (N_16224,N_15159,N_15461);
or U16225 (N_16225,N_15215,N_15277);
nand U16226 (N_16226,N_15807,N_15122);
nand U16227 (N_16227,N_15857,N_15247);
nand U16228 (N_16228,N_15989,N_15990);
xnor U16229 (N_16229,N_15967,N_15241);
xor U16230 (N_16230,N_15896,N_15102);
or U16231 (N_16231,N_15862,N_15556);
or U16232 (N_16232,N_15880,N_15961);
nor U16233 (N_16233,N_15025,N_15333);
or U16234 (N_16234,N_15954,N_15373);
and U16235 (N_16235,N_15879,N_15191);
xor U16236 (N_16236,N_15593,N_15644);
nand U16237 (N_16237,N_15107,N_15123);
or U16238 (N_16238,N_15654,N_15421);
or U16239 (N_16239,N_15926,N_15511);
or U16240 (N_16240,N_15994,N_15771);
xor U16241 (N_16241,N_15881,N_15489);
or U16242 (N_16242,N_15442,N_15457);
nand U16243 (N_16243,N_15727,N_15496);
and U16244 (N_16244,N_15766,N_15953);
or U16245 (N_16245,N_15825,N_15532);
and U16246 (N_16246,N_15261,N_15334);
nor U16247 (N_16247,N_15217,N_15731);
nor U16248 (N_16248,N_15844,N_15007);
nor U16249 (N_16249,N_15768,N_15834);
or U16250 (N_16250,N_15608,N_15794);
xnor U16251 (N_16251,N_15145,N_15583);
xor U16252 (N_16252,N_15299,N_15477);
or U16253 (N_16253,N_15304,N_15419);
nor U16254 (N_16254,N_15772,N_15120);
nor U16255 (N_16255,N_15072,N_15833);
nor U16256 (N_16256,N_15943,N_15870);
nor U16257 (N_16257,N_15529,N_15935);
and U16258 (N_16258,N_15045,N_15291);
or U16259 (N_16259,N_15028,N_15501);
nand U16260 (N_16260,N_15382,N_15667);
xor U16261 (N_16261,N_15450,N_15264);
xor U16262 (N_16262,N_15446,N_15104);
and U16263 (N_16263,N_15016,N_15988);
nor U16264 (N_16264,N_15966,N_15097);
nor U16265 (N_16265,N_15314,N_15543);
nor U16266 (N_16266,N_15580,N_15301);
and U16267 (N_16267,N_15745,N_15756);
and U16268 (N_16268,N_15030,N_15199);
xor U16269 (N_16269,N_15483,N_15182);
or U16270 (N_16270,N_15973,N_15470);
or U16271 (N_16271,N_15959,N_15459);
and U16272 (N_16272,N_15213,N_15346);
or U16273 (N_16273,N_15300,N_15708);
xnor U16274 (N_16274,N_15468,N_15231);
xor U16275 (N_16275,N_15998,N_15188);
or U16276 (N_16276,N_15019,N_15150);
nand U16277 (N_16277,N_15658,N_15655);
nor U16278 (N_16278,N_15273,N_15900);
nand U16279 (N_16279,N_15568,N_15734);
or U16280 (N_16280,N_15510,N_15936);
nand U16281 (N_16281,N_15787,N_15203);
or U16282 (N_16282,N_15599,N_15927);
and U16283 (N_16283,N_15683,N_15377);
nor U16284 (N_16284,N_15773,N_15846);
nor U16285 (N_16285,N_15817,N_15504);
nand U16286 (N_16286,N_15951,N_15684);
and U16287 (N_16287,N_15586,N_15063);
or U16288 (N_16288,N_15596,N_15741);
nor U16289 (N_16289,N_15245,N_15023);
and U16290 (N_16290,N_15995,N_15265);
nor U16291 (N_16291,N_15414,N_15474);
xor U16292 (N_16292,N_15337,N_15315);
or U16293 (N_16293,N_15562,N_15329);
nand U16294 (N_16294,N_15144,N_15719);
nand U16295 (N_16295,N_15984,N_15445);
and U16296 (N_16296,N_15307,N_15194);
and U16297 (N_16297,N_15022,N_15427);
xor U16298 (N_16298,N_15531,N_15415);
xnor U16299 (N_16299,N_15456,N_15095);
nand U16300 (N_16300,N_15069,N_15020);
nor U16301 (N_16301,N_15938,N_15789);
xnor U16302 (N_16302,N_15824,N_15733);
xnor U16303 (N_16303,N_15889,N_15723);
xor U16304 (N_16304,N_15347,N_15193);
and U16305 (N_16305,N_15251,N_15051);
or U16306 (N_16306,N_15544,N_15229);
nor U16307 (N_16307,N_15597,N_15278);
xnor U16308 (N_16308,N_15905,N_15515);
nand U16309 (N_16309,N_15110,N_15207);
or U16310 (N_16310,N_15673,N_15396);
xor U16311 (N_16311,N_15134,N_15381);
xor U16312 (N_16312,N_15692,N_15864);
xor U16313 (N_16313,N_15431,N_15553);
nor U16314 (N_16314,N_15801,N_15336);
and U16315 (N_16315,N_15576,N_15475);
nand U16316 (N_16316,N_15061,N_15664);
nand U16317 (N_16317,N_15037,N_15681);
or U16318 (N_16318,N_15352,N_15043);
or U16319 (N_16319,N_15526,N_15810);
nor U16320 (N_16320,N_15958,N_15176);
nor U16321 (N_16321,N_15670,N_15594);
nand U16322 (N_16322,N_15950,N_15621);
xor U16323 (N_16323,N_15564,N_15624);
and U16324 (N_16324,N_15762,N_15076);
nor U16325 (N_16325,N_15606,N_15487);
and U16326 (N_16326,N_15331,N_15124);
xnor U16327 (N_16327,N_15290,N_15651);
and U16328 (N_16328,N_15344,N_15742);
nand U16329 (N_16329,N_15676,N_15536);
nor U16330 (N_16330,N_15094,N_15392);
nand U16331 (N_16331,N_15792,N_15878);
nand U16332 (N_16332,N_15886,N_15490);
and U16333 (N_16333,N_15726,N_15937);
and U16334 (N_16334,N_15661,N_15296);
and U16335 (N_16335,N_15326,N_15567);
nor U16336 (N_16336,N_15800,N_15901);
nand U16337 (N_16337,N_15652,N_15327);
xnor U16338 (N_16338,N_15946,N_15822);
and U16339 (N_16339,N_15385,N_15238);
nor U16340 (N_16340,N_15046,N_15031);
xor U16341 (N_16341,N_15162,N_15355);
nor U16342 (N_16342,N_15735,N_15538);
or U16343 (N_16343,N_15788,N_15388);
nor U16344 (N_16344,N_15874,N_15574);
nand U16345 (N_16345,N_15424,N_15808);
nand U16346 (N_16346,N_15945,N_15744);
nor U16347 (N_16347,N_15430,N_15859);
nand U16348 (N_16348,N_15906,N_15932);
xor U16349 (N_16349,N_15010,N_15782);
and U16350 (N_16350,N_15917,N_15413);
and U16351 (N_16351,N_15009,N_15281);
xnor U16352 (N_16352,N_15410,N_15048);
and U16353 (N_16353,N_15631,N_15796);
nor U16354 (N_16354,N_15910,N_15674);
or U16355 (N_16355,N_15236,N_15204);
nor U16356 (N_16356,N_15904,N_15765);
and U16357 (N_16357,N_15039,N_15407);
xor U16358 (N_16358,N_15197,N_15963);
nor U16359 (N_16359,N_15508,N_15169);
and U16360 (N_16360,N_15032,N_15836);
or U16361 (N_16361,N_15924,N_15310);
nand U16362 (N_16362,N_15493,N_15297);
and U16363 (N_16363,N_15353,N_15912);
nand U16364 (N_16364,N_15793,N_15619);
xnor U16365 (N_16365,N_15363,N_15979);
nand U16366 (N_16366,N_15227,N_15915);
nor U16367 (N_16367,N_15418,N_15081);
nand U16368 (N_16368,N_15965,N_15324);
nor U16369 (N_16369,N_15049,N_15365);
nor U16370 (N_16370,N_15693,N_15090);
nand U16371 (N_16371,N_15609,N_15091);
nand U16372 (N_16372,N_15283,N_15891);
xor U16373 (N_16373,N_15516,N_15389);
or U16374 (N_16374,N_15933,N_15863);
and U16375 (N_16375,N_15402,N_15981);
nor U16376 (N_16376,N_15017,N_15230);
or U16377 (N_16377,N_15420,N_15187);
xor U16378 (N_16378,N_15902,N_15653);
and U16379 (N_16379,N_15630,N_15115);
xor U16380 (N_16380,N_15976,N_15546);
or U16381 (N_16381,N_15448,N_15026);
and U16382 (N_16382,N_15121,N_15908);
nand U16383 (N_16383,N_15545,N_15471);
nand U16384 (N_16384,N_15635,N_15055);
or U16385 (N_16385,N_15293,N_15033);
nor U16386 (N_16386,N_15752,N_15694);
nand U16387 (N_16387,N_15969,N_15399);
nand U16388 (N_16388,N_15738,N_15537);
nand U16389 (N_16389,N_15226,N_15152);
xnor U16390 (N_16390,N_15364,N_15454);
xnor U16391 (N_16391,N_15704,N_15186);
and U16392 (N_16392,N_15746,N_15366);
and U16393 (N_16393,N_15092,N_15136);
or U16394 (N_16394,N_15157,N_15584);
xnor U16395 (N_16395,N_15798,N_15109);
xor U16396 (N_16396,N_15620,N_15103);
nor U16397 (N_16397,N_15126,N_15767);
and U16398 (N_16398,N_15164,N_15632);
nand U16399 (N_16399,N_15128,N_15433);
or U16400 (N_16400,N_15080,N_15149);
nor U16401 (N_16401,N_15764,N_15610);
or U16402 (N_16402,N_15481,N_15209);
or U16403 (N_16403,N_15922,N_15755);
nor U16404 (N_16404,N_15074,N_15495);
nand U16405 (N_16405,N_15790,N_15894);
or U16406 (N_16406,N_15696,N_15171);
or U16407 (N_16407,N_15462,N_15751);
and U16408 (N_16408,N_15982,N_15687);
nand U16409 (N_16409,N_15663,N_15359);
or U16410 (N_16410,N_15439,N_15441);
or U16411 (N_16411,N_15397,N_15101);
and U16412 (N_16412,N_15888,N_15154);
xor U16413 (N_16413,N_15549,N_15140);
and U16414 (N_16414,N_15657,N_15498);
xor U16415 (N_16415,N_15668,N_15601);
and U16416 (N_16416,N_15254,N_15572);
nor U16417 (N_16417,N_15458,N_15234);
or U16418 (N_16418,N_15721,N_15165);
and U16419 (N_16419,N_15228,N_15737);
xor U16420 (N_16420,N_15812,N_15190);
nor U16421 (N_16421,N_15573,N_15041);
and U16422 (N_16422,N_15285,N_15611);
or U16423 (N_16423,N_15426,N_15605);
or U16424 (N_16424,N_15417,N_15161);
or U16425 (N_16425,N_15196,N_15614);
and U16426 (N_16426,N_15944,N_15535);
or U16427 (N_16427,N_15843,N_15073);
nand U16428 (N_16428,N_15340,N_15319);
or U16429 (N_16429,N_15552,N_15083);
and U16430 (N_16430,N_15691,N_15158);
nor U16431 (N_16431,N_15590,N_15153);
or U16432 (N_16432,N_15867,N_15732);
or U16433 (N_16433,N_15075,N_15778);
and U16434 (N_16434,N_15042,N_15815);
nor U16435 (N_16435,N_15003,N_15561);
nand U16436 (N_16436,N_15575,N_15612);
nor U16437 (N_16437,N_15416,N_15369);
and U16438 (N_16438,N_15279,N_15077);
xor U16439 (N_16439,N_15192,N_15004);
nand U16440 (N_16440,N_15513,N_15015);
and U16441 (N_16441,N_15505,N_15705);
nor U16442 (N_16442,N_15305,N_15449);
nor U16443 (N_16443,N_15047,N_15890);
nand U16444 (N_16444,N_15135,N_15521);
nor U16445 (N_16445,N_15321,N_15839);
nor U16446 (N_16446,N_15362,N_15754);
nor U16447 (N_16447,N_15662,N_15641);
nor U16448 (N_16448,N_15971,N_15001);
and U16449 (N_16449,N_15155,N_15830);
or U16450 (N_16450,N_15195,N_15712);
or U16451 (N_16451,N_15239,N_15071);
and U16452 (N_16452,N_15400,N_15847);
xor U16453 (N_16453,N_15323,N_15403);
or U16454 (N_16454,N_15312,N_15444);
or U16455 (N_16455,N_15432,N_15100);
or U16456 (N_16456,N_15838,N_15222);
xor U16457 (N_16457,N_15964,N_15625);
xnor U16458 (N_16458,N_15776,N_15759);
or U16459 (N_16459,N_15453,N_15660);
nand U16460 (N_16460,N_15589,N_15548);
and U16461 (N_16461,N_15786,N_15804);
nand U16462 (N_16462,N_15434,N_15920);
and U16463 (N_16463,N_15318,N_15582);
xnor U16464 (N_16464,N_15698,N_15539);
xor U16465 (N_16465,N_15690,N_15282);
nand U16466 (N_16466,N_15682,N_15002);
nand U16467 (N_16467,N_15244,N_15117);
nor U16468 (N_16468,N_15820,N_15923);
or U16469 (N_16469,N_15777,N_15250);
and U16470 (N_16470,N_15713,N_15803);
or U16471 (N_16471,N_15156,N_15404);
nor U16472 (N_16472,N_15588,N_15547);
or U16473 (N_16473,N_15235,N_15383);
and U16474 (N_16474,N_15571,N_15185);
nand U16475 (N_16475,N_15865,N_15079);
nor U16476 (N_16476,N_15617,N_15991);
nand U16477 (N_16477,N_15106,N_15907);
nor U16478 (N_16478,N_15177,N_15087);
xnor U16479 (N_16479,N_15749,N_15639);
nor U16480 (N_16480,N_15774,N_15897);
and U16481 (N_16481,N_15328,N_15317);
nand U16482 (N_16482,N_15616,N_15903);
nor U16483 (N_16483,N_15257,N_15711);
nand U16484 (N_16484,N_15736,N_15368);
nand U16485 (N_16485,N_15518,N_15174);
nand U16486 (N_16486,N_15499,N_15716);
nor U16487 (N_16487,N_15488,N_15861);
or U16488 (N_16488,N_15460,N_15147);
nor U16489 (N_16489,N_15637,N_15205);
nor U16490 (N_16490,N_15137,N_15853);
nor U16491 (N_16491,N_15027,N_15797);
or U16492 (N_16492,N_15223,N_15519);
nor U16493 (N_16493,N_15826,N_15221);
and U16494 (N_16494,N_15656,N_15256);
xnor U16495 (N_16495,N_15492,N_15557);
or U16496 (N_16496,N_15968,N_15868);
xor U16497 (N_16497,N_15411,N_15875);
nand U16498 (N_16498,N_15208,N_15686);
and U16499 (N_16499,N_15378,N_15067);
nand U16500 (N_16500,N_15335,N_15916);
and U16501 (N_16501,N_15174,N_15682);
nand U16502 (N_16502,N_15281,N_15363);
nand U16503 (N_16503,N_15977,N_15364);
nand U16504 (N_16504,N_15294,N_15970);
and U16505 (N_16505,N_15242,N_15257);
xnor U16506 (N_16506,N_15079,N_15049);
nand U16507 (N_16507,N_15083,N_15652);
nand U16508 (N_16508,N_15727,N_15211);
and U16509 (N_16509,N_15494,N_15417);
xor U16510 (N_16510,N_15023,N_15951);
or U16511 (N_16511,N_15848,N_15355);
and U16512 (N_16512,N_15349,N_15291);
and U16513 (N_16513,N_15147,N_15689);
nand U16514 (N_16514,N_15628,N_15218);
or U16515 (N_16515,N_15737,N_15222);
and U16516 (N_16516,N_15752,N_15225);
and U16517 (N_16517,N_15325,N_15397);
xnor U16518 (N_16518,N_15343,N_15047);
nor U16519 (N_16519,N_15571,N_15246);
xnor U16520 (N_16520,N_15282,N_15797);
and U16521 (N_16521,N_15752,N_15771);
or U16522 (N_16522,N_15246,N_15688);
or U16523 (N_16523,N_15405,N_15116);
and U16524 (N_16524,N_15144,N_15635);
xnor U16525 (N_16525,N_15836,N_15252);
xor U16526 (N_16526,N_15943,N_15538);
and U16527 (N_16527,N_15291,N_15883);
and U16528 (N_16528,N_15667,N_15040);
nor U16529 (N_16529,N_15703,N_15251);
or U16530 (N_16530,N_15844,N_15860);
or U16531 (N_16531,N_15329,N_15309);
nand U16532 (N_16532,N_15014,N_15436);
and U16533 (N_16533,N_15015,N_15160);
nor U16534 (N_16534,N_15541,N_15926);
and U16535 (N_16535,N_15102,N_15680);
nand U16536 (N_16536,N_15284,N_15375);
or U16537 (N_16537,N_15038,N_15543);
and U16538 (N_16538,N_15723,N_15967);
xor U16539 (N_16539,N_15584,N_15828);
nor U16540 (N_16540,N_15791,N_15306);
nor U16541 (N_16541,N_15046,N_15565);
nor U16542 (N_16542,N_15219,N_15855);
xor U16543 (N_16543,N_15251,N_15634);
nor U16544 (N_16544,N_15567,N_15325);
nand U16545 (N_16545,N_15054,N_15253);
and U16546 (N_16546,N_15987,N_15670);
and U16547 (N_16547,N_15309,N_15914);
nor U16548 (N_16548,N_15437,N_15838);
and U16549 (N_16549,N_15186,N_15629);
nand U16550 (N_16550,N_15850,N_15703);
xor U16551 (N_16551,N_15656,N_15726);
or U16552 (N_16552,N_15546,N_15326);
nor U16553 (N_16553,N_15351,N_15838);
or U16554 (N_16554,N_15230,N_15980);
nand U16555 (N_16555,N_15283,N_15513);
nand U16556 (N_16556,N_15045,N_15267);
or U16557 (N_16557,N_15796,N_15743);
xnor U16558 (N_16558,N_15862,N_15375);
nand U16559 (N_16559,N_15450,N_15899);
or U16560 (N_16560,N_15153,N_15796);
and U16561 (N_16561,N_15774,N_15772);
nor U16562 (N_16562,N_15811,N_15349);
nor U16563 (N_16563,N_15229,N_15943);
or U16564 (N_16564,N_15824,N_15261);
and U16565 (N_16565,N_15741,N_15705);
nand U16566 (N_16566,N_15204,N_15875);
and U16567 (N_16567,N_15764,N_15668);
and U16568 (N_16568,N_15836,N_15446);
nand U16569 (N_16569,N_15576,N_15314);
nor U16570 (N_16570,N_15900,N_15978);
xor U16571 (N_16571,N_15084,N_15104);
nor U16572 (N_16572,N_15502,N_15204);
and U16573 (N_16573,N_15661,N_15136);
and U16574 (N_16574,N_15171,N_15729);
xor U16575 (N_16575,N_15755,N_15563);
xnor U16576 (N_16576,N_15227,N_15972);
or U16577 (N_16577,N_15632,N_15189);
xor U16578 (N_16578,N_15813,N_15474);
nor U16579 (N_16579,N_15062,N_15650);
nand U16580 (N_16580,N_15189,N_15680);
or U16581 (N_16581,N_15833,N_15767);
nand U16582 (N_16582,N_15409,N_15959);
nor U16583 (N_16583,N_15336,N_15388);
xnor U16584 (N_16584,N_15526,N_15196);
or U16585 (N_16585,N_15160,N_15593);
nand U16586 (N_16586,N_15169,N_15124);
and U16587 (N_16587,N_15795,N_15668);
and U16588 (N_16588,N_15380,N_15500);
xor U16589 (N_16589,N_15589,N_15016);
nor U16590 (N_16590,N_15921,N_15401);
nor U16591 (N_16591,N_15026,N_15282);
nor U16592 (N_16592,N_15286,N_15172);
and U16593 (N_16593,N_15588,N_15363);
nor U16594 (N_16594,N_15273,N_15413);
nand U16595 (N_16595,N_15263,N_15486);
or U16596 (N_16596,N_15106,N_15975);
and U16597 (N_16597,N_15442,N_15073);
nor U16598 (N_16598,N_15508,N_15577);
and U16599 (N_16599,N_15959,N_15348);
xor U16600 (N_16600,N_15483,N_15410);
and U16601 (N_16601,N_15435,N_15945);
nor U16602 (N_16602,N_15456,N_15826);
or U16603 (N_16603,N_15472,N_15436);
xor U16604 (N_16604,N_15167,N_15363);
and U16605 (N_16605,N_15927,N_15150);
nor U16606 (N_16606,N_15184,N_15208);
and U16607 (N_16607,N_15685,N_15832);
nand U16608 (N_16608,N_15153,N_15621);
nor U16609 (N_16609,N_15349,N_15817);
or U16610 (N_16610,N_15821,N_15358);
xnor U16611 (N_16611,N_15072,N_15672);
or U16612 (N_16612,N_15633,N_15108);
nand U16613 (N_16613,N_15491,N_15346);
or U16614 (N_16614,N_15504,N_15484);
and U16615 (N_16615,N_15860,N_15525);
and U16616 (N_16616,N_15421,N_15620);
and U16617 (N_16617,N_15081,N_15058);
nor U16618 (N_16618,N_15810,N_15274);
or U16619 (N_16619,N_15951,N_15823);
xor U16620 (N_16620,N_15544,N_15671);
nor U16621 (N_16621,N_15491,N_15226);
xor U16622 (N_16622,N_15301,N_15418);
or U16623 (N_16623,N_15199,N_15749);
xnor U16624 (N_16624,N_15963,N_15621);
xor U16625 (N_16625,N_15779,N_15087);
nor U16626 (N_16626,N_15397,N_15886);
or U16627 (N_16627,N_15726,N_15685);
nand U16628 (N_16628,N_15174,N_15722);
xor U16629 (N_16629,N_15023,N_15852);
nor U16630 (N_16630,N_15272,N_15846);
and U16631 (N_16631,N_15172,N_15105);
or U16632 (N_16632,N_15676,N_15019);
and U16633 (N_16633,N_15253,N_15506);
and U16634 (N_16634,N_15663,N_15226);
and U16635 (N_16635,N_15374,N_15831);
and U16636 (N_16636,N_15214,N_15400);
and U16637 (N_16637,N_15290,N_15501);
xor U16638 (N_16638,N_15963,N_15945);
or U16639 (N_16639,N_15738,N_15655);
xor U16640 (N_16640,N_15742,N_15667);
nand U16641 (N_16641,N_15301,N_15505);
and U16642 (N_16642,N_15147,N_15838);
and U16643 (N_16643,N_15950,N_15151);
nand U16644 (N_16644,N_15355,N_15467);
and U16645 (N_16645,N_15389,N_15515);
and U16646 (N_16646,N_15347,N_15944);
nand U16647 (N_16647,N_15922,N_15966);
nand U16648 (N_16648,N_15753,N_15780);
nor U16649 (N_16649,N_15696,N_15397);
or U16650 (N_16650,N_15422,N_15039);
or U16651 (N_16651,N_15253,N_15724);
and U16652 (N_16652,N_15151,N_15615);
or U16653 (N_16653,N_15194,N_15467);
nand U16654 (N_16654,N_15585,N_15856);
nand U16655 (N_16655,N_15845,N_15644);
nor U16656 (N_16656,N_15471,N_15197);
nand U16657 (N_16657,N_15769,N_15008);
xnor U16658 (N_16658,N_15490,N_15091);
xnor U16659 (N_16659,N_15877,N_15869);
nand U16660 (N_16660,N_15881,N_15570);
nor U16661 (N_16661,N_15807,N_15126);
and U16662 (N_16662,N_15221,N_15497);
nand U16663 (N_16663,N_15374,N_15143);
nor U16664 (N_16664,N_15833,N_15094);
and U16665 (N_16665,N_15625,N_15749);
nand U16666 (N_16666,N_15114,N_15326);
xor U16667 (N_16667,N_15708,N_15231);
nor U16668 (N_16668,N_15786,N_15020);
nand U16669 (N_16669,N_15280,N_15737);
xnor U16670 (N_16670,N_15461,N_15479);
nor U16671 (N_16671,N_15356,N_15943);
xnor U16672 (N_16672,N_15635,N_15902);
or U16673 (N_16673,N_15457,N_15657);
nand U16674 (N_16674,N_15420,N_15903);
nor U16675 (N_16675,N_15683,N_15031);
nor U16676 (N_16676,N_15271,N_15018);
nor U16677 (N_16677,N_15694,N_15736);
and U16678 (N_16678,N_15796,N_15283);
and U16679 (N_16679,N_15078,N_15537);
xnor U16680 (N_16680,N_15998,N_15075);
or U16681 (N_16681,N_15061,N_15779);
nand U16682 (N_16682,N_15604,N_15131);
and U16683 (N_16683,N_15141,N_15199);
and U16684 (N_16684,N_15573,N_15263);
or U16685 (N_16685,N_15288,N_15745);
or U16686 (N_16686,N_15572,N_15562);
and U16687 (N_16687,N_15080,N_15977);
nor U16688 (N_16688,N_15873,N_15389);
or U16689 (N_16689,N_15886,N_15361);
or U16690 (N_16690,N_15907,N_15042);
or U16691 (N_16691,N_15840,N_15136);
and U16692 (N_16692,N_15005,N_15313);
or U16693 (N_16693,N_15835,N_15742);
or U16694 (N_16694,N_15654,N_15054);
or U16695 (N_16695,N_15441,N_15567);
or U16696 (N_16696,N_15118,N_15794);
and U16697 (N_16697,N_15814,N_15816);
and U16698 (N_16698,N_15766,N_15049);
nor U16699 (N_16699,N_15821,N_15750);
nor U16700 (N_16700,N_15013,N_15311);
xor U16701 (N_16701,N_15965,N_15242);
and U16702 (N_16702,N_15138,N_15305);
or U16703 (N_16703,N_15337,N_15041);
xnor U16704 (N_16704,N_15212,N_15672);
nand U16705 (N_16705,N_15307,N_15706);
xnor U16706 (N_16706,N_15592,N_15851);
and U16707 (N_16707,N_15761,N_15896);
nor U16708 (N_16708,N_15238,N_15837);
or U16709 (N_16709,N_15189,N_15078);
xnor U16710 (N_16710,N_15382,N_15562);
nand U16711 (N_16711,N_15907,N_15311);
or U16712 (N_16712,N_15771,N_15988);
nand U16713 (N_16713,N_15835,N_15967);
and U16714 (N_16714,N_15501,N_15275);
nand U16715 (N_16715,N_15439,N_15909);
or U16716 (N_16716,N_15610,N_15801);
or U16717 (N_16717,N_15866,N_15230);
xor U16718 (N_16718,N_15407,N_15030);
or U16719 (N_16719,N_15357,N_15067);
nand U16720 (N_16720,N_15568,N_15467);
or U16721 (N_16721,N_15118,N_15915);
nor U16722 (N_16722,N_15273,N_15645);
and U16723 (N_16723,N_15423,N_15726);
nand U16724 (N_16724,N_15438,N_15889);
nand U16725 (N_16725,N_15911,N_15685);
or U16726 (N_16726,N_15512,N_15445);
and U16727 (N_16727,N_15285,N_15347);
or U16728 (N_16728,N_15635,N_15121);
nand U16729 (N_16729,N_15331,N_15363);
and U16730 (N_16730,N_15789,N_15437);
nand U16731 (N_16731,N_15990,N_15160);
or U16732 (N_16732,N_15795,N_15395);
nor U16733 (N_16733,N_15456,N_15117);
xor U16734 (N_16734,N_15701,N_15479);
and U16735 (N_16735,N_15378,N_15294);
and U16736 (N_16736,N_15595,N_15408);
nor U16737 (N_16737,N_15246,N_15359);
xor U16738 (N_16738,N_15458,N_15516);
xor U16739 (N_16739,N_15990,N_15042);
xnor U16740 (N_16740,N_15268,N_15469);
nand U16741 (N_16741,N_15038,N_15465);
nand U16742 (N_16742,N_15305,N_15018);
nand U16743 (N_16743,N_15466,N_15649);
nand U16744 (N_16744,N_15867,N_15459);
nand U16745 (N_16745,N_15300,N_15443);
and U16746 (N_16746,N_15314,N_15275);
xnor U16747 (N_16747,N_15263,N_15256);
or U16748 (N_16748,N_15882,N_15401);
and U16749 (N_16749,N_15121,N_15356);
or U16750 (N_16750,N_15678,N_15267);
nor U16751 (N_16751,N_15847,N_15372);
xor U16752 (N_16752,N_15268,N_15608);
or U16753 (N_16753,N_15231,N_15738);
nand U16754 (N_16754,N_15183,N_15288);
nor U16755 (N_16755,N_15178,N_15648);
nor U16756 (N_16756,N_15476,N_15852);
nor U16757 (N_16757,N_15781,N_15208);
nor U16758 (N_16758,N_15535,N_15223);
nor U16759 (N_16759,N_15818,N_15983);
and U16760 (N_16760,N_15904,N_15342);
nand U16761 (N_16761,N_15059,N_15687);
and U16762 (N_16762,N_15495,N_15114);
nor U16763 (N_16763,N_15127,N_15991);
or U16764 (N_16764,N_15847,N_15190);
xor U16765 (N_16765,N_15982,N_15324);
and U16766 (N_16766,N_15890,N_15300);
and U16767 (N_16767,N_15233,N_15914);
and U16768 (N_16768,N_15108,N_15014);
nand U16769 (N_16769,N_15484,N_15805);
nand U16770 (N_16770,N_15390,N_15740);
or U16771 (N_16771,N_15074,N_15168);
nor U16772 (N_16772,N_15515,N_15795);
or U16773 (N_16773,N_15569,N_15791);
or U16774 (N_16774,N_15385,N_15091);
nor U16775 (N_16775,N_15457,N_15979);
xnor U16776 (N_16776,N_15891,N_15848);
and U16777 (N_16777,N_15017,N_15902);
and U16778 (N_16778,N_15781,N_15620);
and U16779 (N_16779,N_15706,N_15262);
xor U16780 (N_16780,N_15380,N_15743);
nor U16781 (N_16781,N_15224,N_15641);
and U16782 (N_16782,N_15484,N_15904);
xor U16783 (N_16783,N_15827,N_15014);
or U16784 (N_16784,N_15204,N_15443);
and U16785 (N_16785,N_15804,N_15398);
or U16786 (N_16786,N_15299,N_15378);
xor U16787 (N_16787,N_15677,N_15072);
nor U16788 (N_16788,N_15442,N_15739);
or U16789 (N_16789,N_15647,N_15287);
or U16790 (N_16790,N_15191,N_15930);
xnor U16791 (N_16791,N_15400,N_15668);
or U16792 (N_16792,N_15950,N_15443);
and U16793 (N_16793,N_15304,N_15659);
nand U16794 (N_16794,N_15248,N_15007);
nor U16795 (N_16795,N_15876,N_15526);
xnor U16796 (N_16796,N_15438,N_15564);
and U16797 (N_16797,N_15267,N_15065);
or U16798 (N_16798,N_15750,N_15308);
nand U16799 (N_16799,N_15363,N_15770);
nand U16800 (N_16800,N_15515,N_15559);
nor U16801 (N_16801,N_15064,N_15973);
and U16802 (N_16802,N_15746,N_15204);
nor U16803 (N_16803,N_15280,N_15349);
and U16804 (N_16804,N_15693,N_15263);
or U16805 (N_16805,N_15563,N_15836);
xnor U16806 (N_16806,N_15643,N_15321);
and U16807 (N_16807,N_15982,N_15186);
or U16808 (N_16808,N_15134,N_15418);
xor U16809 (N_16809,N_15492,N_15112);
and U16810 (N_16810,N_15526,N_15646);
nand U16811 (N_16811,N_15297,N_15694);
nand U16812 (N_16812,N_15566,N_15397);
xnor U16813 (N_16813,N_15918,N_15768);
nor U16814 (N_16814,N_15026,N_15354);
xor U16815 (N_16815,N_15215,N_15366);
nor U16816 (N_16816,N_15398,N_15378);
and U16817 (N_16817,N_15968,N_15624);
nor U16818 (N_16818,N_15251,N_15970);
xnor U16819 (N_16819,N_15012,N_15816);
nand U16820 (N_16820,N_15603,N_15646);
xnor U16821 (N_16821,N_15524,N_15632);
or U16822 (N_16822,N_15797,N_15198);
or U16823 (N_16823,N_15640,N_15539);
xnor U16824 (N_16824,N_15640,N_15530);
nor U16825 (N_16825,N_15949,N_15928);
nand U16826 (N_16826,N_15588,N_15665);
and U16827 (N_16827,N_15706,N_15976);
nand U16828 (N_16828,N_15448,N_15127);
and U16829 (N_16829,N_15130,N_15912);
xor U16830 (N_16830,N_15441,N_15977);
or U16831 (N_16831,N_15301,N_15189);
and U16832 (N_16832,N_15196,N_15446);
and U16833 (N_16833,N_15036,N_15309);
and U16834 (N_16834,N_15767,N_15846);
or U16835 (N_16835,N_15383,N_15549);
nor U16836 (N_16836,N_15167,N_15411);
or U16837 (N_16837,N_15624,N_15927);
nor U16838 (N_16838,N_15238,N_15844);
xor U16839 (N_16839,N_15118,N_15912);
and U16840 (N_16840,N_15276,N_15230);
xor U16841 (N_16841,N_15577,N_15197);
or U16842 (N_16842,N_15077,N_15500);
or U16843 (N_16843,N_15272,N_15507);
xnor U16844 (N_16844,N_15948,N_15844);
or U16845 (N_16845,N_15543,N_15205);
nand U16846 (N_16846,N_15760,N_15633);
nor U16847 (N_16847,N_15215,N_15367);
nand U16848 (N_16848,N_15593,N_15996);
xnor U16849 (N_16849,N_15833,N_15013);
xor U16850 (N_16850,N_15668,N_15893);
and U16851 (N_16851,N_15126,N_15304);
nor U16852 (N_16852,N_15226,N_15652);
or U16853 (N_16853,N_15651,N_15624);
nor U16854 (N_16854,N_15530,N_15332);
nor U16855 (N_16855,N_15756,N_15819);
nor U16856 (N_16856,N_15926,N_15849);
nand U16857 (N_16857,N_15813,N_15557);
xnor U16858 (N_16858,N_15601,N_15560);
and U16859 (N_16859,N_15871,N_15860);
and U16860 (N_16860,N_15608,N_15066);
and U16861 (N_16861,N_15844,N_15618);
nor U16862 (N_16862,N_15659,N_15487);
nor U16863 (N_16863,N_15912,N_15287);
or U16864 (N_16864,N_15466,N_15513);
xor U16865 (N_16865,N_15724,N_15352);
nor U16866 (N_16866,N_15513,N_15920);
nor U16867 (N_16867,N_15357,N_15103);
xnor U16868 (N_16868,N_15406,N_15941);
nor U16869 (N_16869,N_15570,N_15033);
xor U16870 (N_16870,N_15046,N_15624);
and U16871 (N_16871,N_15752,N_15539);
nor U16872 (N_16872,N_15083,N_15883);
nand U16873 (N_16873,N_15327,N_15236);
or U16874 (N_16874,N_15117,N_15452);
and U16875 (N_16875,N_15063,N_15642);
and U16876 (N_16876,N_15774,N_15863);
nor U16877 (N_16877,N_15811,N_15014);
nor U16878 (N_16878,N_15114,N_15657);
nor U16879 (N_16879,N_15873,N_15664);
and U16880 (N_16880,N_15769,N_15322);
nand U16881 (N_16881,N_15024,N_15879);
and U16882 (N_16882,N_15114,N_15533);
xnor U16883 (N_16883,N_15748,N_15349);
xor U16884 (N_16884,N_15344,N_15399);
or U16885 (N_16885,N_15661,N_15305);
and U16886 (N_16886,N_15549,N_15330);
nor U16887 (N_16887,N_15405,N_15003);
xor U16888 (N_16888,N_15098,N_15024);
and U16889 (N_16889,N_15239,N_15047);
nand U16890 (N_16890,N_15031,N_15816);
or U16891 (N_16891,N_15851,N_15567);
and U16892 (N_16892,N_15050,N_15418);
or U16893 (N_16893,N_15938,N_15456);
and U16894 (N_16894,N_15996,N_15928);
xor U16895 (N_16895,N_15871,N_15290);
and U16896 (N_16896,N_15891,N_15844);
nor U16897 (N_16897,N_15637,N_15683);
nand U16898 (N_16898,N_15004,N_15840);
or U16899 (N_16899,N_15758,N_15814);
nor U16900 (N_16900,N_15904,N_15766);
or U16901 (N_16901,N_15392,N_15437);
or U16902 (N_16902,N_15333,N_15480);
nand U16903 (N_16903,N_15341,N_15193);
xor U16904 (N_16904,N_15557,N_15645);
and U16905 (N_16905,N_15414,N_15506);
nand U16906 (N_16906,N_15856,N_15263);
nand U16907 (N_16907,N_15690,N_15659);
or U16908 (N_16908,N_15375,N_15859);
nand U16909 (N_16909,N_15940,N_15323);
nand U16910 (N_16910,N_15931,N_15351);
nor U16911 (N_16911,N_15274,N_15270);
xnor U16912 (N_16912,N_15276,N_15575);
or U16913 (N_16913,N_15217,N_15070);
nor U16914 (N_16914,N_15393,N_15222);
and U16915 (N_16915,N_15121,N_15443);
or U16916 (N_16916,N_15527,N_15863);
nand U16917 (N_16917,N_15236,N_15669);
and U16918 (N_16918,N_15456,N_15401);
nor U16919 (N_16919,N_15431,N_15045);
nor U16920 (N_16920,N_15054,N_15594);
nor U16921 (N_16921,N_15717,N_15427);
nor U16922 (N_16922,N_15823,N_15629);
nor U16923 (N_16923,N_15786,N_15864);
and U16924 (N_16924,N_15175,N_15034);
xnor U16925 (N_16925,N_15873,N_15071);
nor U16926 (N_16926,N_15324,N_15685);
nand U16927 (N_16927,N_15188,N_15565);
or U16928 (N_16928,N_15390,N_15310);
nor U16929 (N_16929,N_15253,N_15232);
nand U16930 (N_16930,N_15994,N_15821);
xnor U16931 (N_16931,N_15874,N_15774);
or U16932 (N_16932,N_15645,N_15998);
and U16933 (N_16933,N_15442,N_15393);
or U16934 (N_16934,N_15757,N_15431);
and U16935 (N_16935,N_15007,N_15416);
xor U16936 (N_16936,N_15800,N_15705);
nor U16937 (N_16937,N_15644,N_15776);
nor U16938 (N_16938,N_15749,N_15703);
and U16939 (N_16939,N_15124,N_15858);
or U16940 (N_16940,N_15860,N_15280);
nand U16941 (N_16941,N_15145,N_15976);
or U16942 (N_16942,N_15018,N_15379);
or U16943 (N_16943,N_15054,N_15945);
xor U16944 (N_16944,N_15589,N_15512);
and U16945 (N_16945,N_15036,N_15576);
and U16946 (N_16946,N_15465,N_15156);
xor U16947 (N_16947,N_15913,N_15566);
and U16948 (N_16948,N_15699,N_15848);
nor U16949 (N_16949,N_15872,N_15710);
or U16950 (N_16950,N_15934,N_15051);
xnor U16951 (N_16951,N_15159,N_15812);
nand U16952 (N_16952,N_15882,N_15052);
nand U16953 (N_16953,N_15699,N_15800);
or U16954 (N_16954,N_15136,N_15588);
xor U16955 (N_16955,N_15013,N_15890);
or U16956 (N_16956,N_15506,N_15264);
nor U16957 (N_16957,N_15157,N_15786);
or U16958 (N_16958,N_15518,N_15461);
nand U16959 (N_16959,N_15683,N_15711);
and U16960 (N_16960,N_15961,N_15174);
or U16961 (N_16961,N_15803,N_15461);
nand U16962 (N_16962,N_15407,N_15058);
nor U16963 (N_16963,N_15740,N_15844);
and U16964 (N_16964,N_15378,N_15613);
nand U16965 (N_16965,N_15575,N_15091);
xnor U16966 (N_16966,N_15583,N_15134);
nand U16967 (N_16967,N_15181,N_15818);
and U16968 (N_16968,N_15651,N_15387);
nand U16969 (N_16969,N_15460,N_15330);
xnor U16970 (N_16970,N_15438,N_15751);
or U16971 (N_16971,N_15761,N_15921);
and U16972 (N_16972,N_15209,N_15819);
xnor U16973 (N_16973,N_15667,N_15839);
or U16974 (N_16974,N_15407,N_15552);
and U16975 (N_16975,N_15647,N_15164);
and U16976 (N_16976,N_15711,N_15141);
nor U16977 (N_16977,N_15288,N_15197);
nor U16978 (N_16978,N_15397,N_15077);
nand U16979 (N_16979,N_15901,N_15545);
xor U16980 (N_16980,N_15826,N_15404);
nand U16981 (N_16981,N_15871,N_15564);
and U16982 (N_16982,N_15806,N_15225);
and U16983 (N_16983,N_15425,N_15507);
nor U16984 (N_16984,N_15170,N_15094);
nor U16985 (N_16985,N_15534,N_15951);
and U16986 (N_16986,N_15938,N_15247);
and U16987 (N_16987,N_15867,N_15454);
nor U16988 (N_16988,N_15552,N_15116);
or U16989 (N_16989,N_15349,N_15483);
xnor U16990 (N_16990,N_15435,N_15697);
xnor U16991 (N_16991,N_15784,N_15063);
nand U16992 (N_16992,N_15966,N_15316);
nand U16993 (N_16993,N_15280,N_15000);
xnor U16994 (N_16994,N_15750,N_15651);
nand U16995 (N_16995,N_15711,N_15724);
xor U16996 (N_16996,N_15586,N_15075);
and U16997 (N_16997,N_15663,N_15856);
nand U16998 (N_16998,N_15080,N_15746);
nor U16999 (N_16999,N_15900,N_15475);
or U17000 (N_17000,N_16845,N_16737);
xnor U17001 (N_17001,N_16374,N_16042);
or U17002 (N_17002,N_16565,N_16660);
or U17003 (N_17003,N_16753,N_16038);
and U17004 (N_17004,N_16609,N_16037);
nand U17005 (N_17005,N_16978,N_16671);
and U17006 (N_17006,N_16085,N_16640);
xnor U17007 (N_17007,N_16125,N_16452);
nor U17008 (N_17008,N_16213,N_16227);
nor U17009 (N_17009,N_16303,N_16943);
xnor U17010 (N_17010,N_16929,N_16380);
nor U17011 (N_17011,N_16349,N_16500);
and U17012 (N_17012,N_16655,N_16796);
xnor U17013 (N_17013,N_16546,N_16164);
xnor U17014 (N_17014,N_16048,N_16391);
xnor U17015 (N_17015,N_16249,N_16439);
or U17016 (N_17016,N_16714,N_16051);
nor U17017 (N_17017,N_16952,N_16430);
nor U17018 (N_17018,N_16973,N_16091);
nor U17019 (N_17019,N_16088,N_16657);
or U17020 (N_17020,N_16922,N_16661);
nand U17021 (N_17021,N_16616,N_16646);
nor U17022 (N_17022,N_16955,N_16353);
xnor U17023 (N_17023,N_16842,N_16719);
nand U17024 (N_17024,N_16941,N_16309);
nor U17025 (N_17025,N_16871,N_16912);
or U17026 (N_17026,N_16862,N_16369);
and U17027 (N_17027,N_16462,N_16907);
nor U17028 (N_17028,N_16998,N_16666);
and U17029 (N_17029,N_16731,N_16139);
nor U17030 (N_17030,N_16972,N_16035);
xnor U17031 (N_17031,N_16276,N_16734);
nand U17032 (N_17032,N_16224,N_16788);
nor U17033 (N_17033,N_16549,N_16957);
xnor U17034 (N_17034,N_16300,N_16808);
or U17035 (N_17035,N_16449,N_16581);
and U17036 (N_17036,N_16223,N_16852);
and U17037 (N_17037,N_16096,N_16415);
or U17038 (N_17038,N_16521,N_16823);
nand U17039 (N_17039,N_16687,N_16909);
xor U17040 (N_17040,N_16207,N_16018);
nand U17041 (N_17041,N_16115,N_16744);
or U17042 (N_17042,N_16028,N_16116);
nand U17043 (N_17043,N_16890,N_16780);
xor U17044 (N_17044,N_16846,N_16335);
and U17045 (N_17045,N_16323,N_16005);
nor U17046 (N_17046,N_16228,N_16481);
nor U17047 (N_17047,N_16056,N_16601);
nand U17048 (N_17048,N_16149,N_16385);
or U17049 (N_17049,N_16694,N_16988);
or U17050 (N_17050,N_16059,N_16459);
and U17051 (N_17051,N_16670,N_16641);
nor U17052 (N_17052,N_16338,N_16285);
xnor U17053 (N_17053,N_16494,N_16302);
xnor U17054 (N_17054,N_16121,N_16937);
nand U17055 (N_17055,N_16327,N_16861);
nor U17056 (N_17056,N_16069,N_16282);
nor U17057 (N_17057,N_16133,N_16058);
and U17058 (N_17058,N_16013,N_16156);
or U17059 (N_17059,N_16326,N_16736);
nand U17060 (N_17060,N_16638,N_16238);
nand U17061 (N_17061,N_16777,N_16667);
or U17062 (N_17062,N_16821,N_16294);
xor U17063 (N_17063,N_16509,N_16100);
xnor U17064 (N_17064,N_16931,N_16488);
nor U17065 (N_17065,N_16954,N_16273);
xnor U17066 (N_17066,N_16991,N_16816);
or U17067 (N_17067,N_16087,N_16109);
xor U17068 (N_17068,N_16183,N_16317);
or U17069 (N_17069,N_16935,N_16754);
xor U17070 (N_17070,N_16315,N_16726);
nor U17071 (N_17071,N_16226,N_16547);
nor U17072 (N_17072,N_16767,N_16659);
xnor U17073 (N_17073,N_16310,N_16897);
and U17074 (N_17074,N_16468,N_16131);
and U17075 (N_17075,N_16932,N_16411);
nand U17076 (N_17076,N_16432,N_16102);
nor U17077 (N_17077,N_16355,N_16266);
xnor U17078 (N_17078,N_16901,N_16197);
nor U17079 (N_17079,N_16812,N_16877);
and U17080 (N_17080,N_16105,N_16400);
xnor U17081 (N_17081,N_16648,N_16498);
nor U17082 (N_17082,N_16985,N_16225);
nor U17083 (N_17083,N_16321,N_16518);
nand U17084 (N_17084,N_16829,N_16728);
nand U17085 (N_17085,N_16429,N_16182);
nor U17086 (N_17086,N_16160,N_16709);
and U17087 (N_17087,N_16596,N_16017);
and U17088 (N_17088,N_16206,N_16210);
and U17089 (N_17089,N_16624,N_16367);
nor U17090 (N_17090,N_16128,N_16372);
nand U17091 (N_17091,N_16471,N_16440);
nand U17092 (N_17092,N_16524,N_16567);
nor U17093 (N_17093,N_16376,N_16097);
xnor U17094 (N_17094,N_16178,N_16482);
or U17095 (N_17095,N_16365,N_16428);
nor U17096 (N_17096,N_16497,N_16373);
nor U17097 (N_17097,N_16994,N_16838);
and U17098 (N_17098,N_16913,N_16112);
xor U17099 (N_17099,N_16268,N_16553);
or U17100 (N_17100,N_16775,N_16061);
nand U17101 (N_17101,N_16403,N_16964);
nor U17102 (N_17102,N_16702,N_16122);
or U17103 (N_17103,N_16850,N_16426);
and U17104 (N_17104,N_16378,N_16774);
or U17105 (N_17105,N_16712,N_16538);
nor U17106 (N_17106,N_16129,N_16078);
nand U17107 (N_17107,N_16577,N_16730);
nand U17108 (N_17108,N_16633,N_16067);
or U17109 (N_17109,N_16405,N_16643);
nor U17110 (N_17110,N_16689,N_16718);
and U17111 (N_17111,N_16408,N_16404);
nand U17112 (N_17112,N_16570,N_16504);
nand U17113 (N_17113,N_16847,N_16407);
nand U17114 (N_17114,N_16412,N_16642);
nand U17115 (N_17115,N_16352,N_16729);
nor U17116 (N_17116,N_16990,N_16022);
xor U17117 (N_17117,N_16493,N_16906);
nand U17118 (N_17118,N_16047,N_16746);
nand U17119 (N_17119,N_16260,N_16107);
and U17120 (N_17120,N_16123,N_16084);
nand U17121 (N_17121,N_16849,N_16592);
nand U17122 (N_17122,N_16540,N_16695);
and U17123 (N_17123,N_16126,N_16575);
and U17124 (N_17124,N_16668,N_16065);
and U17125 (N_17125,N_16235,N_16794);
xnor U17126 (N_17126,N_16366,N_16942);
xor U17127 (N_17127,N_16340,N_16159);
xor U17128 (N_17128,N_16627,N_16764);
xnor U17129 (N_17129,N_16992,N_16090);
nor U17130 (N_17130,N_16915,N_16157);
and U17131 (N_17131,N_16066,N_16933);
or U17132 (N_17132,N_16830,N_16008);
or U17133 (N_17133,N_16717,N_16630);
or U17134 (N_17134,N_16401,N_16771);
or U17135 (N_17135,N_16211,N_16834);
nand U17136 (N_17136,N_16793,N_16168);
nand U17137 (N_17137,N_16072,N_16926);
nor U17138 (N_17138,N_16899,N_16370);
nand U17139 (N_17139,N_16124,N_16948);
nor U17140 (N_17140,N_16598,N_16856);
or U17141 (N_17141,N_16765,N_16590);
xor U17142 (N_17142,N_16778,N_16247);
nor U17143 (N_17143,N_16284,N_16800);
nor U17144 (N_17144,N_16137,N_16305);
nor U17145 (N_17145,N_16288,N_16086);
nand U17146 (N_17146,N_16081,N_16036);
and U17147 (N_17147,N_16987,N_16701);
xnor U17148 (N_17148,N_16986,N_16316);
nor U17149 (N_17149,N_16611,N_16219);
nor U17150 (N_17150,N_16620,N_16818);
nor U17151 (N_17151,N_16200,N_16446);
and U17152 (N_17152,N_16614,N_16076);
nand U17153 (N_17153,N_16347,N_16716);
and U17154 (N_17154,N_16189,N_16073);
and U17155 (N_17155,N_16381,N_16757);
and U17156 (N_17156,N_16445,N_16786);
and U17157 (N_17157,N_16256,N_16231);
and U17158 (N_17158,N_16761,N_16117);
nor U17159 (N_17159,N_16878,N_16466);
nand U17160 (N_17160,N_16398,N_16708);
nand U17161 (N_17161,N_16433,N_16650);
nor U17162 (N_17162,N_16594,N_16113);
nor U17163 (N_17163,N_16704,N_16141);
and U17164 (N_17164,N_16891,N_16479);
and U17165 (N_17165,N_16216,N_16186);
or U17166 (N_17166,N_16417,N_16951);
or U17167 (N_17167,N_16055,N_16612);
or U17168 (N_17168,N_16114,N_16148);
nor U17169 (N_17169,N_16568,N_16617);
nand U17170 (N_17170,N_16892,N_16527);
and U17171 (N_17171,N_16184,N_16212);
and U17172 (N_17172,N_16817,N_16306);
or U17173 (N_17173,N_16959,N_16467);
and U17174 (N_17174,N_16499,N_16437);
nand U17175 (N_17175,N_16679,N_16104);
xnor U17176 (N_17176,N_16928,N_16738);
and U17177 (N_17177,N_16257,N_16561);
xor U17178 (N_17178,N_16587,N_16755);
nor U17179 (N_17179,N_16881,N_16111);
xor U17180 (N_17180,N_16192,N_16523);
nand U17181 (N_17181,N_16593,N_16873);
xor U17182 (N_17182,N_16875,N_16208);
or U17183 (N_17183,N_16656,N_16278);
nor U17184 (N_17184,N_16060,N_16040);
nand U17185 (N_17185,N_16876,N_16155);
or U17186 (N_17186,N_16784,N_16236);
nand U17187 (N_17187,N_16889,N_16879);
and U17188 (N_17188,N_16371,N_16574);
nor U17189 (N_17189,N_16664,N_16763);
nand U17190 (N_17190,N_16304,N_16244);
nand U17191 (N_17191,N_16531,N_16644);
nor U17192 (N_17192,N_16919,N_16027);
nor U17193 (N_17193,N_16799,N_16825);
or U17194 (N_17194,N_16677,N_16075);
nand U17195 (N_17195,N_16629,N_16248);
nand U17196 (N_17196,N_16914,N_16054);
nand U17197 (N_17197,N_16921,N_16484);
xor U17198 (N_17198,N_16550,N_16153);
and U17199 (N_17199,N_16501,N_16181);
nand U17200 (N_17200,N_16451,N_16289);
xnor U17201 (N_17201,N_16770,N_16680);
xor U17202 (N_17202,N_16406,N_16585);
or U17203 (N_17203,N_16956,N_16064);
and U17204 (N_17204,N_16140,N_16621);
nor U17205 (N_17205,N_16029,N_16607);
and U17206 (N_17206,N_16345,N_16789);
or U17207 (N_17207,N_16217,N_16025);
and U17208 (N_17208,N_16474,N_16456);
xnor U17209 (N_17209,N_16662,N_16743);
or U17210 (N_17210,N_16893,N_16350);
nand U17211 (N_17211,N_16110,N_16286);
xnor U17212 (N_17212,N_16421,N_16868);
xor U17213 (N_17213,N_16172,N_16924);
xnor U17214 (N_17214,N_16724,N_16198);
nand U17215 (N_17215,N_16602,N_16797);
xor U17216 (N_17216,N_16416,N_16293);
and U17217 (N_17217,N_16245,N_16342);
nand U17218 (N_17218,N_16950,N_16635);
nand U17219 (N_17219,N_16977,N_16166);
nand U17220 (N_17220,N_16740,N_16050);
xor U17221 (N_17221,N_16552,N_16475);
or U17222 (N_17222,N_16608,N_16274);
or U17223 (N_17223,N_16544,N_16525);
xor U17224 (N_17224,N_16308,N_16205);
and U17225 (N_17225,N_16558,N_16958);
nand U17226 (N_17226,N_16402,N_16424);
nand U17227 (N_17227,N_16209,N_16887);
nor U17228 (N_17228,N_16572,N_16835);
xnor U17229 (N_17229,N_16083,N_16867);
nor U17230 (N_17230,N_16858,N_16554);
xnor U17231 (N_17231,N_16751,N_16969);
nor U17232 (N_17232,N_16344,N_16324);
nor U17233 (N_17233,N_16357,N_16898);
nor U17234 (N_17234,N_16280,N_16760);
xnor U17235 (N_17235,N_16966,N_16171);
nor U17236 (N_17236,N_16420,N_16291);
and U17237 (N_17237,N_16311,N_16983);
nor U17238 (N_17238,N_16619,N_16343);
and U17239 (N_17239,N_16710,N_16307);
and U17240 (N_17240,N_16979,N_16865);
nor U17241 (N_17241,N_16707,N_16043);
nor U17242 (N_17242,N_16545,N_16672);
or U17243 (N_17243,N_16487,N_16092);
nor U17244 (N_17244,N_16146,N_16174);
or U17245 (N_17245,N_16806,N_16804);
or U17246 (N_17246,N_16927,N_16222);
and U17247 (N_17247,N_16706,N_16422);
xor U17248 (N_17248,N_16827,N_16506);
and U17249 (N_17249,N_16375,N_16283);
or U17250 (N_17250,N_16354,N_16682);
nor U17251 (N_17251,N_16610,N_16271);
nand U17252 (N_17252,N_16551,N_16281);
nand U17253 (N_17253,N_16089,N_16472);
or U17254 (N_17254,N_16194,N_16191);
or U17255 (N_17255,N_16534,N_16588);
xor U17256 (N_17256,N_16505,N_16175);
nand U17257 (N_17257,N_16857,N_16215);
or U17258 (N_17258,N_16169,N_16173);
nand U17259 (N_17259,N_16934,N_16508);
nand U17260 (N_17260,N_16015,N_16193);
and U17261 (N_17261,N_16364,N_16678);
nand U17262 (N_17262,N_16782,N_16787);
and U17263 (N_17263,N_16947,N_16318);
nor U17264 (N_17264,N_16469,N_16815);
or U17265 (N_17265,N_16254,N_16241);
or U17266 (N_17266,N_16233,N_16458);
or U17267 (N_17267,N_16143,N_16563);
nor U17268 (N_17268,N_16536,N_16802);
and U17269 (N_17269,N_16399,N_16533);
xnor U17270 (N_17270,N_16295,N_16997);
or U17271 (N_17271,N_16436,N_16414);
and U17272 (N_17272,N_16049,N_16332);
nor U17273 (N_17273,N_16134,N_16615);
or U17274 (N_17274,N_16605,N_16328);
or U17275 (N_17275,N_16578,N_16267);
nor U17276 (N_17276,N_16622,N_16438);
and U17277 (N_17277,N_16519,N_16095);
or U17278 (N_17278,N_16068,N_16180);
and U17279 (N_17279,N_16296,N_16014);
nand U17280 (N_17280,N_16251,N_16108);
nand U17281 (N_17281,N_16938,N_16801);
xor U17282 (N_17282,N_16388,N_16106);
nand U17283 (N_17283,N_16455,N_16976);
or U17284 (N_17284,N_16700,N_16348);
nand U17285 (N_17285,N_16790,N_16496);
xor U17286 (N_17286,N_16480,N_16094);
nand U17287 (N_17287,N_16855,N_16221);
and U17288 (N_17288,N_16099,N_16541);
or U17289 (N_17289,N_16749,N_16098);
nor U17290 (N_17290,N_16888,N_16167);
or U17291 (N_17291,N_16711,N_16024);
or U17292 (N_17292,N_16831,N_16297);
or U17293 (N_17293,N_16637,N_16674);
and U17294 (N_17294,N_16434,N_16566);
nor U17295 (N_17295,N_16016,N_16591);
or U17296 (N_17296,N_16910,N_16669);
nor U17297 (N_17297,N_16517,N_16154);
xor U17298 (N_17298,N_16880,N_16242);
or U17299 (N_17299,N_16649,N_16093);
and U17300 (N_17300,N_16361,N_16557);
or U17301 (N_17301,N_16623,N_16395);
xnor U17302 (N_17302,N_16511,N_16239);
and U17303 (N_17303,N_16936,N_16034);
or U17304 (N_17304,N_16632,N_16562);
and U17305 (N_17305,N_16826,N_16331);
nor U17306 (N_17306,N_16625,N_16522);
nor U17307 (N_17307,N_16190,N_16177);
and U17308 (N_17308,N_16044,N_16903);
or U17309 (N_17309,N_16651,N_16392);
or U17310 (N_17310,N_16261,N_16170);
xor U17311 (N_17311,N_16776,N_16975);
nand U17312 (N_17312,N_16690,N_16447);
nand U17313 (N_17313,N_16158,N_16514);
or U17314 (N_17314,N_16485,N_16745);
nor U17315 (N_17315,N_16844,N_16337);
xnor U17316 (N_17316,N_16923,N_16009);
nor U17317 (N_17317,N_16971,N_16940);
xnor U17318 (N_17318,N_16684,N_16580);
xor U17319 (N_17319,N_16454,N_16379);
and U17320 (N_17320,N_16489,N_16863);
nand U17321 (N_17321,N_16299,N_16516);
nand U17322 (N_17322,N_16866,N_16628);
nand U17323 (N_17323,N_16441,N_16031);
nor U17324 (N_17324,N_16735,N_16502);
or U17325 (N_17325,N_16739,N_16811);
nor U17326 (N_17326,N_16444,N_16460);
nand U17327 (N_17327,N_16162,N_16033);
nand U17328 (N_17328,N_16232,N_16962);
xor U17329 (N_17329,N_16002,N_16384);
or U17330 (N_17330,N_16859,N_16152);
or U17331 (N_17331,N_16742,N_16699);
nand U17332 (N_17332,N_16253,N_16358);
nand U17333 (N_17333,N_16409,N_16077);
xnor U17334 (N_17334,N_16030,N_16179);
xor U17335 (N_17335,N_16012,N_16006);
xnor U17336 (N_17336,N_16675,N_16272);
or U17337 (N_17337,N_16658,N_16949);
xnor U17338 (N_17338,N_16758,N_16393);
xor U17339 (N_17339,N_16798,N_16756);
xor U17340 (N_17340,N_16532,N_16082);
or U17341 (N_17341,N_16886,N_16410);
nor U17342 (N_17342,N_16457,N_16813);
xor U17343 (N_17343,N_16853,N_16925);
and U17344 (N_17344,N_16431,N_16663);
xor U17345 (N_17345,N_16769,N_16138);
nand U17346 (N_17346,N_16766,N_16142);
nor U17347 (N_17347,N_16387,N_16229);
and U17348 (N_17348,N_16723,N_16750);
nor U17349 (N_17349,N_16240,N_16698);
and U17350 (N_17350,N_16683,N_16301);
nor U17351 (N_17351,N_16872,N_16636);
nor U17352 (N_17352,N_16968,N_16526);
or U17353 (N_17353,N_16673,N_16559);
nor U17354 (N_17354,N_16870,N_16995);
or U17355 (N_17355,N_16443,N_16389);
nor U17356 (N_17356,N_16470,N_16250);
nor U17357 (N_17357,N_16188,N_16270);
nand U17358 (N_17358,N_16974,N_16528);
or U17359 (N_17359,N_16262,N_16537);
nand U17360 (N_17360,N_16483,N_16539);
nand U17361 (N_17361,N_16900,N_16555);
nor U17362 (N_17362,N_16127,N_16599);
nor U17363 (N_17363,N_16394,N_16356);
nor U17364 (N_17364,N_16639,N_16895);
nand U17365 (N_17365,N_16752,N_16686);
and U17366 (N_17366,N_16287,N_16839);
and U17367 (N_17367,N_16851,N_16841);
and U17368 (N_17368,N_16258,N_16052);
and U17369 (N_17369,N_16762,N_16564);
nand U17370 (N_17370,N_16368,N_16916);
and U17371 (N_17371,N_16011,N_16201);
or U17372 (N_17372,N_16960,N_16981);
and U17373 (N_17373,N_16589,N_16860);
xor U17374 (N_17374,N_16713,N_16453);
nor U17375 (N_17375,N_16885,N_16320);
or U17376 (N_17376,N_16722,N_16584);
xor U17377 (N_17377,N_16070,N_16118);
nand U17378 (N_17378,N_16945,N_16010);
or U17379 (N_17379,N_16150,N_16720);
or U17380 (N_17380,N_16917,N_16199);
and U17381 (N_17381,N_16832,N_16634);
or U17382 (N_17382,N_16814,N_16325);
and U17383 (N_17383,N_16843,N_16848);
nor U17384 (N_17384,N_16996,N_16195);
xor U17385 (N_17385,N_16779,N_16147);
nand U17386 (N_17386,N_16882,N_16019);
nor U17387 (N_17387,N_16967,N_16529);
nor U17388 (N_17388,N_16290,N_16999);
and U17389 (N_17389,N_16606,N_16363);
and U17390 (N_17390,N_16869,N_16252);
nor U17391 (N_17391,N_16715,N_16319);
and U17392 (N_17392,N_16822,N_16151);
and U17393 (N_17393,N_16419,N_16904);
nor U17394 (N_17394,N_16103,N_16548);
xnor U17395 (N_17395,N_16597,N_16645);
nor U17396 (N_17396,N_16676,N_16530);
nor U17397 (N_17397,N_16259,N_16136);
or U17398 (N_17398,N_16057,N_16603);
or U17399 (N_17399,N_16542,N_16980);
xor U17400 (N_17400,N_16101,N_16697);
nand U17401 (N_17401,N_16579,N_16275);
xnor U17402 (N_17402,N_16383,N_16161);
nand U17403 (N_17403,N_16185,N_16360);
nand U17404 (N_17404,N_16573,N_16571);
nor U17405 (N_17405,N_16423,N_16390);
and U17406 (N_17406,N_16512,N_16359);
xnor U17407 (N_17407,N_16586,N_16336);
and U17408 (N_17408,N_16450,N_16946);
xnor U17409 (N_17409,N_16833,N_16448);
or U17410 (N_17410,N_16004,N_16944);
xor U17411 (N_17411,N_16733,N_16809);
and U17412 (N_17412,N_16080,N_16618);
and U17413 (N_17413,N_16039,N_16418);
nand U17414 (N_17414,N_16196,N_16569);
or U17415 (N_17415,N_16237,N_16230);
nand U17416 (N_17416,N_16819,N_16377);
xnor U17417 (N_17417,N_16074,N_16836);
nand U17418 (N_17418,N_16220,N_16595);
and U17419 (N_17419,N_16135,N_16071);
or U17420 (N_17420,N_16486,N_16810);
xor U17421 (N_17421,N_16351,N_16894);
nand U17422 (N_17422,N_16463,N_16464);
nand U17423 (N_17423,N_16785,N_16792);
xnor U17424 (N_17424,N_16854,N_16298);
nand U17425 (N_17425,N_16747,N_16490);
xor U17426 (N_17426,N_16727,N_16970);
and U17427 (N_17427,N_16246,N_16492);
nor U17428 (N_17428,N_16626,N_16692);
or U17429 (N_17429,N_16465,N_16911);
nand U17430 (N_17430,N_16007,N_16313);
nor U17431 (N_17431,N_16119,N_16243);
nand U17432 (N_17432,N_16582,N_16427);
or U17433 (N_17433,N_16053,N_16510);
nor U17434 (N_17434,N_16314,N_16652);
nor U17435 (N_17435,N_16515,N_16218);
or U17436 (N_17436,N_16144,N_16312);
nand U17437 (N_17437,N_16828,N_16908);
nor U17438 (N_17438,N_16026,N_16725);
xor U17439 (N_17439,N_16003,N_16883);
or U17440 (N_17440,N_16329,N_16681);
and U17441 (N_17441,N_16292,N_16993);
nand U17442 (N_17442,N_16902,N_16791);
or U17443 (N_17443,N_16984,N_16214);
or U17444 (N_17444,N_16965,N_16543);
or U17445 (N_17445,N_16896,N_16203);
xnor U17446 (N_17446,N_16269,N_16783);
nor U17447 (N_17447,N_16583,N_16560);
nor U17448 (N_17448,N_16795,N_16333);
nand U17449 (N_17449,N_16535,N_16079);
nor U17450 (N_17450,N_16120,N_16691);
or U17451 (N_17451,N_16062,N_16930);
or U17452 (N_17452,N_16130,N_16461);
or U17453 (N_17453,N_16920,N_16693);
or U17454 (N_17454,N_16768,N_16647);
and U17455 (N_17455,N_16413,N_16021);
or U17456 (N_17456,N_16513,N_16478);
nand U17457 (N_17457,N_16032,N_16665);
xor U17458 (N_17458,N_16145,N_16346);
nor U17459 (N_17459,N_16264,N_16781);
nand U17460 (N_17460,N_16442,N_16397);
xor U17461 (N_17461,N_16654,N_16600);
or U17462 (N_17462,N_16685,N_16772);
nand U17463 (N_17463,N_16631,N_16386);
xnor U17464 (N_17464,N_16653,N_16202);
or U17465 (N_17465,N_16805,N_16382);
xnor U17466 (N_17466,N_16803,N_16020);
and U17467 (N_17467,N_16473,N_16023);
nor U17468 (N_17468,N_16163,N_16263);
nand U17469 (N_17469,N_16187,N_16435);
and U17470 (N_17470,N_16759,N_16884);
nor U17471 (N_17471,N_16425,N_16696);
xnor U17472 (N_17472,N_16063,N_16864);
nand U17473 (N_17473,N_16824,N_16476);
nor U17474 (N_17474,N_16322,N_16046);
nand U17475 (N_17475,N_16576,N_16905);
or U17476 (N_17476,N_16001,N_16982);
or U17477 (N_17477,N_16953,N_16807);
or U17478 (N_17478,N_16165,N_16989);
xor U17479 (N_17479,N_16495,N_16613);
nor U17480 (N_17480,N_16277,N_16334);
and U17481 (N_17481,N_16477,N_16732);
and U17482 (N_17482,N_16918,N_16703);
and U17483 (N_17483,N_16265,N_16963);
and U17484 (N_17484,N_16396,N_16279);
or U17485 (N_17485,N_16341,N_16939);
and U17486 (N_17486,N_16748,N_16362);
or U17487 (N_17487,N_16132,N_16705);
nor U17488 (N_17488,N_16204,N_16491);
nand U17489 (N_17489,N_16520,N_16041);
xor U17490 (N_17490,N_16255,N_16339);
nand U17491 (N_17491,N_16045,N_16556);
nor U17492 (N_17492,N_16741,N_16507);
or U17493 (N_17493,N_16503,N_16820);
xnor U17494 (N_17494,N_16840,N_16330);
xnor U17495 (N_17495,N_16000,N_16721);
and U17496 (N_17496,N_16773,N_16176);
or U17497 (N_17497,N_16874,N_16234);
and U17498 (N_17498,N_16688,N_16837);
nand U17499 (N_17499,N_16961,N_16604);
nor U17500 (N_17500,N_16011,N_16366);
and U17501 (N_17501,N_16589,N_16379);
nor U17502 (N_17502,N_16858,N_16518);
nand U17503 (N_17503,N_16315,N_16539);
or U17504 (N_17504,N_16060,N_16030);
nor U17505 (N_17505,N_16568,N_16135);
nor U17506 (N_17506,N_16379,N_16638);
nand U17507 (N_17507,N_16134,N_16438);
xor U17508 (N_17508,N_16743,N_16251);
xor U17509 (N_17509,N_16659,N_16992);
xor U17510 (N_17510,N_16741,N_16857);
xnor U17511 (N_17511,N_16419,N_16060);
or U17512 (N_17512,N_16320,N_16642);
and U17513 (N_17513,N_16880,N_16434);
or U17514 (N_17514,N_16939,N_16167);
xnor U17515 (N_17515,N_16771,N_16324);
xor U17516 (N_17516,N_16165,N_16595);
nand U17517 (N_17517,N_16028,N_16249);
nor U17518 (N_17518,N_16861,N_16683);
nor U17519 (N_17519,N_16836,N_16577);
nor U17520 (N_17520,N_16299,N_16205);
or U17521 (N_17521,N_16091,N_16075);
xnor U17522 (N_17522,N_16275,N_16743);
and U17523 (N_17523,N_16794,N_16834);
and U17524 (N_17524,N_16410,N_16198);
nor U17525 (N_17525,N_16884,N_16921);
or U17526 (N_17526,N_16334,N_16550);
xnor U17527 (N_17527,N_16675,N_16200);
nor U17528 (N_17528,N_16499,N_16751);
and U17529 (N_17529,N_16786,N_16061);
or U17530 (N_17530,N_16948,N_16113);
xnor U17531 (N_17531,N_16601,N_16394);
nor U17532 (N_17532,N_16001,N_16996);
xor U17533 (N_17533,N_16983,N_16003);
nand U17534 (N_17534,N_16597,N_16005);
nand U17535 (N_17535,N_16055,N_16682);
and U17536 (N_17536,N_16513,N_16149);
xnor U17537 (N_17537,N_16343,N_16770);
nand U17538 (N_17538,N_16834,N_16697);
nand U17539 (N_17539,N_16903,N_16900);
xnor U17540 (N_17540,N_16067,N_16949);
and U17541 (N_17541,N_16376,N_16028);
nor U17542 (N_17542,N_16341,N_16138);
nand U17543 (N_17543,N_16380,N_16629);
nand U17544 (N_17544,N_16381,N_16882);
and U17545 (N_17545,N_16899,N_16321);
xor U17546 (N_17546,N_16416,N_16302);
nand U17547 (N_17547,N_16941,N_16088);
or U17548 (N_17548,N_16194,N_16069);
and U17549 (N_17549,N_16359,N_16187);
nor U17550 (N_17550,N_16230,N_16551);
nor U17551 (N_17551,N_16229,N_16123);
nor U17552 (N_17552,N_16184,N_16436);
and U17553 (N_17553,N_16671,N_16856);
and U17554 (N_17554,N_16907,N_16150);
or U17555 (N_17555,N_16358,N_16456);
xor U17556 (N_17556,N_16368,N_16456);
xnor U17557 (N_17557,N_16344,N_16526);
nor U17558 (N_17558,N_16404,N_16674);
nor U17559 (N_17559,N_16098,N_16946);
nor U17560 (N_17560,N_16505,N_16248);
nand U17561 (N_17561,N_16633,N_16997);
nand U17562 (N_17562,N_16487,N_16790);
nand U17563 (N_17563,N_16112,N_16979);
or U17564 (N_17564,N_16342,N_16897);
and U17565 (N_17565,N_16325,N_16782);
and U17566 (N_17566,N_16618,N_16394);
and U17567 (N_17567,N_16673,N_16021);
nand U17568 (N_17568,N_16295,N_16881);
nor U17569 (N_17569,N_16814,N_16961);
nand U17570 (N_17570,N_16607,N_16944);
xor U17571 (N_17571,N_16155,N_16127);
nand U17572 (N_17572,N_16983,N_16985);
nand U17573 (N_17573,N_16006,N_16168);
nand U17574 (N_17574,N_16796,N_16388);
nor U17575 (N_17575,N_16564,N_16023);
xor U17576 (N_17576,N_16279,N_16649);
and U17577 (N_17577,N_16890,N_16759);
and U17578 (N_17578,N_16836,N_16236);
nand U17579 (N_17579,N_16087,N_16920);
xnor U17580 (N_17580,N_16928,N_16836);
xor U17581 (N_17581,N_16975,N_16747);
xnor U17582 (N_17582,N_16370,N_16765);
nor U17583 (N_17583,N_16388,N_16752);
nor U17584 (N_17584,N_16574,N_16226);
xor U17585 (N_17585,N_16033,N_16774);
nor U17586 (N_17586,N_16655,N_16884);
or U17587 (N_17587,N_16571,N_16395);
xnor U17588 (N_17588,N_16623,N_16742);
and U17589 (N_17589,N_16460,N_16456);
nor U17590 (N_17590,N_16466,N_16169);
and U17591 (N_17591,N_16759,N_16963);
nand U17592 (N_17592,N_16691,N_16541);
or U17593 (N_17593,N_16902,N_16961);
nand U17594 (N_17594,N_16101,N_16950);
nand U17595 (N_17595,N_16239,N_16097);
nand U17596 (N_17596,N_16279,N_16218);
xnor U17597 (N_17597,N_16657,N_16662);
and U17598 (N_17598,N_16719,N_16651);
or U17599 (N_17599,N_16981,N_16869);
or U17600 (N_17600,N_16870,N_16767);
and U17601 (N_17601,N_16357,N_16756);
and U17602 (N_17602,N_16774,N_16272);
xor U17603 (N_17603,N_16910,N_16215);
nand U17604 (N_17604,N_16862,N_16512);
nor U17605 (N_17605,N_16469,N_16942);
xnor U17606 (N_17606,N_16966,N_16056);
nor U17607 (N_17607,N_16112,N_16536);
or U17608 (N_17608,N_16078,N_16147);
and U17609 (N_17609,N_16098,N_16103);
or U17610 (N_17610,N_16973,N_16413);
nor U17611 (N_17611,N_16867,N_16787);
nor U17612 (N_17612,N_16434,N_16476);
nand U17613 (N_17613,N_16679,N_16972);
nand U17614 (N_17614,N_16044,N_16323);
nor U17615 (N_17615,N_16495,N_16612);
and U17616 (N_17616,N_16770,N_16431);
xnor U17617 (N_17617,N_16274,N_16178);
xor U17618 (N_17618,N_16163,N_16336);
xor U17619 (N_17619,N_16355,N_16879);
nor U17620 (N_17620,N_16442,N_16171);
nor U17621 (N_17621,N_16532,N_16475);
nor U17622 (N_17622,N_16247,N_16438);
nor U17623 (N_17623,N_16621,N_16310);
and U17624 (N_17624,N_16242,N_16238);
nand U17625 (N_17625,N_16043,N_16023);
xnor U17626 (N_17626,N_16020,N_16325);
nor U17627 (N_17627,N_16708,N_16782);
xor U17628 (N_17628,N_16270,N_16240);
nand U17629 (N_17629,N_16535,N_16347);
nor U17630 (N_17630,N_16508,N_16447);
nand U17631 (N_17631,N_16414,N_16160);
or U17632 (N_17632,N_16063,N_16355);
or U17633 (N_17633,N_16615,N_16801);
nand U17634 (N_17634,N_16178,N_16342);
xnor U17635 (N_17635,N_16613,N_16910);
xnor U17636 (N_17636,N_16106,N_16513);
nand U17637 (N_17637,N_16963,N_16877);
and U17638 (N_17638,N_16445,N_16994);
nand U17639 (N_17639,N_16810,N_16546);
nor U17640 (N_17640,N_16905,N_16756);
or U17641 (N_17641,N_16053,N_16266);
nor U17642 (N_17642,N_16604,N_16757);
and U17643 (N_17643,N_16350,N_16072);
xnor U17644 (N_17644,N_16750,N_16174);
or U17645 (N_17645,N_16000,N_16746);
and U17646 (N_17646,N_16395,N_16307);
and U17647 (N_17647,N_16018,N_16445);
nor U17648 (N_17648,N_16130,N_16691);
xor U17649 (N_17649,N_16528,N_16557);
and U17650 (N_17650,N_16670,N_16406);
and U17651 (N_17651,N_16472,N_16027);
or U17652 (N_17652,N_16045,N_16759);
xor U17653 (N_17653,N_16072,N_16098);
nand U17654 (N_17654,N_16559,N_16726);
and U17655 (N_17655,N_16018,N_16679);
xor U17656 (N_17656,N_16343,N_16673);
nor U17657 (N_17657,N_16943,N_16889);
and U17658 (N_17658,N_16834,N_16670);
nand U17659 (N_17659,N_16138,N_16218);
or U17660 (N_17660,N_16507,N_16032);
nor U17661 (N_17661,N_16599,N_16005);
or U17662 (N_17662,N_16121,N_16620);
nor U17663 (N_17663,N_16164,N_16319);
xnor U17664 (N_17664,N_16203,N_16804);
nand U17665 (N_17665,N_16969,N_16175);
xor U17666 (N_17666,N_16677,N_16901);
or U17667 (N_17667,N_16807,N_16310);
nand U17668 (N_17668,N_16486,N_16649);
and U17669 (N_17669,N_16426,N_16729);
or U17670 (N_17670,N_16339,N_16977);
or U17671 (N_17671,N_16141,N_16594);
or U17672 (N_17672,N_16339,N_16731);
and U17673 (N_17673,N_16523,N_16411);
and U17674 (N_17674,N_16661,N_16715);
xnor U17675 (N_17675,N_16212,N_16384);
and U17676 (N_17676,N_16033,N_16871);
nor U17677 (N_17677,N_16058,N_16575);
and U17678 (N_17678,N_16288,N_16123);
nand U17679 (N_17679,N_16252,N_16191);
nor U17680 (N_17680,N_16818,N_16800);
nor U17681 (N_17681,N_16059,N_16914);
and U17682 (N_17682,N_16658,N_16511);
and U17683 (N_17683,N_16681,N_16394);
nor U17684 (N_17684,N_16590,N_16540);
nand U17685 (N_17685,N_16432,N_16591);
nand U17686 (N_17686,N_16014,N_16645);
and U17687 (N_17687,N_16990,N_16408);
and U17688 (N_17688,N_16587,N_16365);
xnor U17689 (N_17689,N_16249,N_16819);
nand U17690 (N_17690,N_16732,N_16170);
and U17691 (N_17691,N_16417,N_16569);
nor U17692 (N_17692,N_16470,N_16128);
nor U17693 (N_17693,N_16290,N_16300);
nor U17694 (N_17694,N_16672,N_16719);
xnor U17695 (N_17695,N_16188,N_16844);
nand U17696 (N_17696,N_16162,N_16110);
or U17697 (N_17697,N_16378,N_16535);
xor U17698 (N_17698,N_16320,N_16072);
xnor U17699 (N_17699,N_16447,N_16140);
xor U17700 (N_17700,N_16452,N_16805);
or U17701 (N_17701,N_16261,N_16202);
and U17702 (N_17702,N_16729,N_16681);
or U17703 (N_17703,N_16872,N_16282);
nor U17704 (N_17704,N_16849,N_16449);
xnor U17705 (N_17705,N_16634,N_16728);
xor U17706 (N_17706,N_16534,N_16418);
and U17707 (N_17707,N_16690,N_16862);
xor U17708 (N_17708,N_16376,N_16114);
nand U17709 (N_17709,N_16757,N_16107);
xor U17710 (N_17710,N_16959,N_16092);
or U17711 (N_17711,N_16856,N_16946);
nor U17712 (N_17712,N_16649,N_16769);
and U17713 (N_17713,N_16701,N_16800);
and U17714 (N_17714,N_16834,N_16413);
or U17715 (N_17715,N_16965,N_16706);
nand U17716 (N_17716,N_16607,N_16895);
and U17717 (N_17717,N_16672,N_16065);
and U17718 (N_17718,N_16797,N_16468);
xnor U17719 (N_17719,N_16576,N_16111);
xor U17720 (N_17720,N_16152,N_16213);
and U17721 (N_17721,N_16566,N_16820);
nor U17722 (N_17722,N_16205,N_16714);
and U17723 (N_17723,N_16404,N_16735);
and U17724 (N_17724,N_16277,N_16117);
nand U17725 (N_17725,N_16361,N_16772);
nor U17726 (N_17726,N_16396,N_16850);
and U17727 (N_17727,N_16036,N_16693);
or U17728 (N_17728,N_16290,N_16911);
and U17729 (N_17729,N_16163,N_16446);
nand U17730 (N_17730,N_16238,N_16821);
and U17731 (N_17731,N_16609,N_16925);
nand U17732 (N_17732,N_16050,N_16542);
nand U17733 (N_17733,N_16982,N_16008);
nor U17734 (N_17734,N_16603,N_16926);
nand U17735 (N_17735,N_16864,N_16327);
xnor U17736 (N_17736,N_16328,N_16388);
xnor U17737 (N_17737,N_16101,N_16549);
nor U17738 (N_17738,N_16124,N_16872);
xnor U17739 (N_17739,N_16321,N_16046);
nand U17740 (N_17740,N_16641,N_16967);
nand U17741 (N_17741,N_16293,N_16887);
and U17742 (N_17742,N_16719,N_16529);
nand U17743 (N_17743,N_16280,N_16550);
or U17744 (N_17744,N_16477,N_16046);
and U17745 (N_17745,N_16355,N_16255);
nor U17746 (N_17746,N_16416,N_16086);
and U17747 (N_17747,N_16753,N_16968);
xor U17748 (N_17748,N_16781,N_16951);
nor U17749 (N_17749,N_16577,N_16284);
nor U17750 (N_17750,N_16171,N_16016);
xor U17751 (N_17751,N_16961,N_16466);
nand U17752 (N_17752,N_16805,N_16258);
and U17753 (N_17753,N_16188,N_16291);
nor U17754 (N_17754,N_16235,N_16501);
or U17755 (N_17755,N_16438,N_16352);
nand U17756 (N_17756,N_16341,N_16566);
and U17757 (N_17757,N_16866,N_16837);
xor U17758 (N_17758,N_16919,N_16269);
nor U17759 (N_17759,N_16755,N_16763);
nor U17760 (N_17760,N_16080,N_16157);
nand U17761 (N_17761,N_16712,N_16958);
nor U17762 (N_17762,N_16980,N_16040);
or U17763 (N_17763,N_16787,N_16965);
nor U17764 (N_17764,N_16536,N_16843);
xnor U17765 (N_17765,N_16228,N_16234);
nor U17766 (N_17766,N_16568,N_16828);
xnor U17767 (N_17767,N_16769,N_16202);
and U17768 (N_17768,N_16476,N_16944);
xor U17769 (N_17769,N_16275,N_16472);
xnor U17770 (N_17770,N_16753,N_16983);
and U17771 (N_17771,N_16686,N_16851);
and U17772 (N_17772,N_16078,N_16449);
or U17773 (N_17773,N_16693,N_16718);
or U17774 (N_17774,N_16633,N_16933);
nor U17775 (N_17775,N_16045,N_16749);
and U17776 (N_17776,N_16330,N_16355);
nor U17777 (N_17777,N_16318,N_16796);
and U17778 (N_17778,N_16635,N_16795);
or U17779 (N_17779,N_16349,N_16868);
or U17780 (N_17780,N_16456,N_16942);
nor U17781 (N_17781,N_16565,N_16386);
nor U17782 (N_17782,N_16591,N_16126);
nand U17783 (N_17783,N_16624,N_16491);
or U17784 (N_17784,N_16024,N_16330);
and U17785 (N_17785,N_16949,N_16679);
nand U17786 (N_17786,N_16709,N_16536);
xnor U17787 (N_17787,N_16526,N_16337);
and U17788 (N_17788,N_16893,N_16357);
and U17789 (N_17789,N_16198,N_16555);
and U17790 (N_17790,N_16023,N_16951);
and U17791 (N_17791,N_16924,N_16137);
and U17792 (N_17792,N_16555,N_16573);
and U17793 (N_17793,N_16923,N_16278);
nand U17794 (N_17794,N_16339,N_16476);
nor U17795 (N_17795,N_16963,N_16352);
and U17796 (N_17796,N_16284,N_16346);
nand U17797 (N_17797,N_16241,N_16448);
and U17798 (N_17798,N_16238,N_16491);
xnor U17799 (N_17799,N_16058,N_16096);
or U17800 (N_17800,N_16345,N_16044);
nand U17801 (N_17801,N_16249,N_16205);
nand U17802 (N_17802,N_16145,N_16322);
nor U17803 (N_17803,N_16739,N_16149);
xor U17804 (N_17804,N_16153,N_16577);
and U17805 (N_17805,N_16189,N_16219);
or U17806 (N_17806,N_16059,N_16157);
or U17807 (N_17807,N_16382,N_16550);
nand U17808 (N_17808,N_16173,N_16388);
and U17809 (N_17809,N_16362,N_16325);
or U17810 (N_17810,N_16086,N_16474);
or U17811 (N_17811,N_16520,N_16122);
nand U17812 (N_17812,N_16077,N_16679);
xor U17813 (N_17813,N_16068,N_16941);
nand U17814 (N_17814,N_16008,N_16239);
or U17815 (N_17815,N_16920,N_16317);
nor U17816 (N_17816,N_16553,N_16305);
nor U17817 (N_17817,N_16287,N_16168);
nand U17818 (N_17818,N_16528,N_16370);
or U17819 (N_17819,N_16174,N_16498);
nor U17820 (N_17820,N_16344,N_16851);
nand U17821 (N_17821,N_16736,N_16052);
nand U17822 (N_17822,N_16831,N_16000);
nand U17823 (N_17823,N_16777,N_16519);
or U17824 (N_17824,N_16746,N_16298);
nand U17825 (N_17825,N_16007,N_16747);
and U17826 (N_17826,N_16033,N_16611);
nand U17827 (N_17827,N_16035,N_16851);
or U17828 (N_17828,N_16790,N_16159);
or U17829 (N_17829,N_16591,N_16095);
xnor U17830 (N_17830,N_16223,N_16056);
nor U17831 (N_17831,N_16425,N_16831);
and U17832 (N_17832,N_16537,N_16221);
nand U17833 (N_17833,N_16453,N_16173);
xnor U17834 (N_17834,N_16607,N_16691);
nor U17835 (N_17835,N_16671,N_16487);
and U17836 (N_17836,N_16464,N_16425);
or U17837 (N_17837,N_16618,N_16999);
and U17838 (N_17838,N_16716,N_16084);
nor U17839 (N_17839,N_16456,N_16312);
or U17840 (N_17840,N_16395,N_16779);
and U17841 (N_17841,N_16122,N_16938);
nand U17842 (N_17842,N_16500,N_16003);
and U17843 (N_17843,N_16650,N_16781);
xor U17844 (N_17844,N_16128,N_16102);
and U17845 (N_17845,N_16885,N_16809);
nand U17846 (N_17846,N_16836,N_16393);
xor U17847 (N_17847,N_16423,N_16379);
and U17848 (N_17848,N_16079,N_16620);
nand U17849 (N_17849,N_16416,N_16978);
xnor U17850 (N_17850,N_16307,N_16384);
and U17851 (N_17851,N_16031,N_16454);
xor U17852 (N_17852,N_16905,N_16659);
nor U17853 (N_17853,N_16003,N_16409);
and U17854 (N_17854,N_16629,N_16635);
nand U17855 (N_17855,N_16103,N_16924);
nand U17856 (N_17856,N_16060,N_16352);
nand U17857 (N_17857,N_16588,N_16300);
or U17858 (N_17858,N_16104,N_16376);
nor U17859 (N_17859,N_16153,N_16879);
and U17860 (N_17860,N_16672,N_16098);
or U17861 (N_17861,N_16322,N_16981);
and U17862 (N_17862,N_16919,N_16642);
and U17863 (N_17863,N_16344,N_16437);
or U17864 (N_17864,N_16456,N_16101);
or U17865 (N_17865,N_16613,N_16899);
or U17866 (N_17866,N_16087,N_16495);
and U17867 (N_17867,N_16657,N_16310);
xor U17868 (N_17868,N_16319,N_16300);
nor U17869 (N_17869,N_16617,N_16277);
and U17870 (N_17870,N_16248,N_16369);
nor U17871 (N_17871,N_16398,N_16872);
nor U17872 (N_17872,N_16223,N_16963);
or U17873 (N_17873,N_16362,N_16521);
xor U17874 (N_17874,N_16789,N_16288);
nand U17875 (N_17875,N_16240,N_16258);
nor U17876 (N_17876,N_16435,N_16423);
nor U17877 (N_17877,N_16772,N_16878);
nand U17878 (N_17878,N_16336,N_16526);
nor U17879 (N_17879,N_16535,N_16503);
nor U17880 (N_17880,N_16213,N_16518);
or U17881 (N_17881,N_16181,N_16510);
nand U17882 (N_17882,N_16571,N_16157);
nand U17883 (N_17883,N_16675,N_16038);
xor U17884 (N_17884,N_16636,N_16097);
xor U17885 (N_17885,N_16164,N_16040);
and U17886 (N_17886,N_16056,N_16797);
or U17887 (N_17887,N_16054,N_16460);
or U17888 (N_17888,N_16387,N_16223);
or U17889 (N_17889,N_16407,N_16276);
or U17890 (N_17890,N_16927,N_16236);
and U17891 (N_17891,N_16770,N_16283);
nand U17892 (N_17892,N_16504,N_16402);
and U17893 (N_17893,N_16486,N_16062);
nand U17894 (N_17894,N_16414,N_16876);
nor U17895 (N_17895,N_16329,N_16370);
or U17896 (N_17896,N_16218,N_16582);
and U17897 (N_17897,N_16140,N_16258);
nor U17898 (N_17898,N_16459,N_16494);
or U17899 (N_17899,N_16987,N_16456);
nor U17900 (N_17900,N_16538,N_16161);
and U17901 (N_17901,N_16556,N_16287);
nor U17902 (N_17902,N_16365,N_16597);
xor U17903 (N_17903,N_16663,N_16683);
xnor U17904 (N_17904,N_16028,N_16944);
nor U17905 (N_17905,N_16818,N_16610);
xor U17906 (N_17906,N_16571,N_16661);
xnor U17907 (N_17907,N_16948,N_16676);
and U17908 (N_17908,N_16043,N_16027);
nor U17909 (N_17909,N_16338,N_16700);
xor U17910 (N_17910,N_16388,N_16141);
or U17911 (N_17911,N_16875,N_16758);
nor U17912 (N_17912,N_16535,N_16815);
xor U17913 (N_17913,N_16243,N_16947);
nand U17914 (N_17914,N_16718,N_16686);
nand U17915 (N_17915,N_16009,N_16249);
and U17916 (N_17916,N_16301,N_16366);
nand U17917 (N_17917,N_16550,N_16074);
or U17918 (N_17918,N_16802,N_16320);
xnor U17919 (N_17919,N_16866,N_16934);
or U17920 (N_17920,N_16278,N_16240);
or U17921 (N_17921,N_16641,N_16159);
nand U17922 (N_17922,N_16967,N_16181);
nor U17923 (N_17923,N_16417,N_16058);
and U17924 (N_17924,N_16106,N_16597);
nor U17925 (N_17925,N_16997,N_16078);
xor U17926 (N_17926,N_16469,N_16707);
nor U17927 (N_17927,N_16561,N_16737);
or U17928 (N_17928,N_16847,N_16405);
or U17929 (N_17929,N_16884,N_16905);
nor U17930 (N_17930,N_16013,N_16080);
xnor U17931 (N_17931,N_16090,N_16144);
nor U17932 (N_17932,N_16064,N_16505);
nand U17933 (N_17933,N_16008,N_16558);
or U17934 (N_17934,N_16279,N_16784);
nor U17935 (N_17935,N_16341,N_16745);
nand U17936 (N_17936,N_16311,N_16064);
nor U17937 (N_17937,N_16492,N_16017);
or U17938 (N_17938,N_16338,N_16632);
or U17939 (N_17939,N_16457,N_16814);
xnor U17940 (N_17940,N_16557,N_16017);
or U17941 (N_17941,N_16611,N_16695);
or U17942 (N_17942,N_16445,N_16197);
nor U17943 (N_17943,N_16046,N_16292);
nor U17944 (N_17944,N_16288,N_16836);
and U17945 (N_17945,N_16197,N_16832);
nand U17946 (N_17946,N_16166,N_16665);
nor U17947 (N_17947,N_16092,N_16402);
nor U17948 (N_17948,N_16113,N_16472);
or U17949 (N_17949,N_16223,N_16206);
and U17950 (N_17950,N_16986,N_16344);
and U17951 (N_17951,N_16665,N_16375);
nand U17952 (N_17952,N_16643,N_16169);
nand U17953 (N_17953,N_16914,N_16061);
or U17954 (N_17954,N_16657,N_16960);
nor U17955 (N_17955,N_16743,N_16868);
xor U17956 (N_17956,N_16669,N_16403);
nor U17957 (N_17957,N_16591,N_16101);
nand U17958 (N_17958,N_16282,N_16415);
nand U17959 (N_17959,N_16633,N_16349);
nor U17960 (N_17960,N_16725,N_16014);
and U17961 (N_17961,N_16229,N_16146);
nand U17962 (N_17962,N_16564,N_16011);
and U17963 (N_17963,N_16079,N_16189);
and U17964 (N_17964,N_16179,N_16031);
nand U17965 (N_17965,N_16285,N_16393);
or U17966 (N_17966,N_16833,N_16988);
nand U17967 (N_17967,N_16167,N_16975);
nand U17968 (N_17968,N_16056,N_16410);
nor U17969 (N_17969,N_16175,N_16771);
or U17970 (N_17970,N_16342,N_16136);
nor U17971 (N_17971,N_16869,N_16056);
nand U17972 (N_17972,N_16968,N_16862);
or U17973 (N_17973,N_16164,N_16157);
nor U17974 (N_17974,N_16284,N_16265);
or U17975 (N_17975,N_16709,N_16650);
nor U17976 (N_17976,N_16350,N_16533);
xnor U17977 (N_17977,N_16847,N_16033);
or U17978 (N_17978,N_16617,N_16395);
and U17979 (N_17979,N_16111,N_16952);
or U17980 (N_17980,N_16577,N_16645);
nor U17981 (N_17981,N_16564,N_16285);
and U17982 (N_17982,N_16127,N_16439);
xnor U17983 (N_17983,N_16931,N_16668);
nor U17984 (N_17984,N_16522,N_16403);
or U17985 (N_17985,N_16051,N_16816);
xor U17986 (N_17986,N_16446,N_16945);
xnor U17987 (N_17987,N_16184,N_16094);
nor U17988 (N_17988,N_16533,N_16027);
nor U17989 (N_17989,N_16346,N_16000);
and U17990 (N_17990,N_16095,N_16367);
nand U17991 (N_17991,N_16724,N_16220);
and U17992 (N_17992,N_16767,N_16867);
and U17993 (N_17993,N_16163,N_16824);
and U17994 (N_17994,N_16650,N_16044);
xor U17995 (N_17995,N_16522,N_16831);
nor U17996 (N_17996,N_16055,N_16148);
nor U17997 (N_17997,N_16595,N_16786);
and U17998 (N_17998,N_16266,N_16894);
nor U17999 (N_17999,N_16341,N_16216);
xnor U18000 (N_18000,N_17085,N_17851);
nor U18001 (N_18001,N_17253,N_17523);
and U18002 (N_18002,N_17105,N_17667);
and U18003 (N_18003,N_17129,N_17058);
or U18004 (N_18004,N_17005,N_17010);
or U18005 (N_18005,N_17850,N_17399);
nor U18006 (N_18006,N_17741,N_17266);
nand U18007 (N_18007,N_17090,N_17421);
xnor U18008 (N_18008,N_17844,N_17080);
and U18009 (N_18009,N_17219,N_17494);
nand U18010 (N_18010,N_17541,N_17201);
nor U18011 (N_18011,N_17736,N_17830);
or U18012 (N_18012,N_17789,N_17819);
and U18013 (N_18013,N_17134,N_17318);
and U18014 (N_18014,N_17576,N_17986);
xor U18015 (N_18015,N_17743,N_17021);
and U18016 (N_18016,N_17904,N_17867);
or U18017 (N_18017,N_17978,N_17972);
or U18018 (N_18018,N_17766,N_17346);
and U18019 (N_18019,N_17653,N_17485);
xor U18020 (N_18020,N_17094,N_17498);
and U18021 (N_18021,N_17968,N_17301);
and U18022 (N_18022,N_17983,N_17344);
nor U18023 (N_18023,N_17567,N_17024);
or U18024 (N_18024,N_17483,N_17896);
and U18025 (N_18025,N_17918,N_17173);
and U18026 (N_18026,N_17232,N_17803);
xnor U18027 (N_18027,N_17098,N_17869);
and U18028 (N_18028,N_17103,N_17153);
nand U18029 (N_18029,N_17744,N_17397);
xnor U18030 (N_18030,N_17988,N_17964);
xor U18031 (N_18031,N_17514,N_17855);
nand U18032 (N_18032,N_17303,N_17176);
xor U18033 (N_18033,N_17734,N_17965);
nor U18034 (N_18034,N_17463,N_17490);
nand U18035 (N_18035,N_17990,N_17525);
or U18036 (N_18036,N_17345,N_17834);
xnor U18037 (N_18037,N_17617,N_17782);
nand U18038 (N_18038,N_17499,N_17033);
or U18039 (N_18039,N_17070,N_17293);
xor U18040 (N_18040,N_17280,N_17190);
or U18041 (N_18041,N_17724,N_17439);
nor U18042 (N_18042,N_17754,N_17276);
nand U18043 (N_18043,N_17012,N_17601);
nand U18044 (N_18044,N_17703,N_17756);
or U18045 (N_18045,N_17057,N_17360);
or U18046 (N_18046,N_17967,N_17611);
nand U18047 (N_18047,N_17702,N_17627);
or U18048 (N_18048,N_17875,N_17832);
or U18049 (N_18049,N_17079,N_17258);
nand U18050 (N_18050,N_17477,N_17681);
nand U18051 (N_18051,N_17763,N_17113);
xnor U18052 (N_18052,N_17150,N_17952);
xnor U18053 (N_18053,N_17308,N_17051);
xor U18054 (N_18054,N_17448,N_17372);
nor U18055 (N_18055,N_17535,N_17287);
and U18056 (N_18056,N_17456,N_17050);
or U18057 (N_18057,N_17092,N_17846);
xnor U18058 (N_18058,N_17487,N_17445);
or U18059 (N_18059,N_17532,N_17404);
nand U18060 (N_18060,N_17479,N_17778);
and U18061 (N_18061,N_17809,N_17274);
xnor U18062 (N_18062,N_17250,N_17154);
xnor U18063 (N_18063,N_17292,N_17779);
xor U18064 (N_18064,N_17504,N_17859);
nand U18065 (N_18065,N_17704,N_17164);
or U18066 (N_18066,N_17424,N_17314);
nor U18067 (N_18067,N_17296,N_17429);
or U18068 (N_18068,N_17670,N_17542);
xnor U18069 (N_18069,N_17249,N_17116);
nand U18070 (N_18070,N_17179,N_17997);
or U18071 (N_18071,N_17014,N_17174);
nor U18072 (N_18072,N_17631,N_17822);
nor U18073 (N_18073,N_17947,N_17999);
or U18074 (N_18074,N_17570,N_17242);
and U18075 (N_18075,N_17141,N_17267);
nand U18076 (N_18076,N_17353,N_17003);
or U18077 (N_18077,N_17261,N_17211);
xnor U18078 (N_18078,N_17086,N_17534);
or U18079 (N_18079,N_17957,N_17886);
nor U18080 (N_18080,N_17874,N_17520);
nand U18081 (N_18081,N_17112,N_17143);
xnor U18082 (N_18082,N_17884,N_17686);
nand U18083 (N_18083,N_17671,N_17157);
and U18084 (N_18084,N_17528,N_17434);
xor U18085 (N_18085,N_17979,N_17698);
or U18086 (N_18086,N_17807,N_17139);
xor U18087 (N_18087,N_17664,N_17548);
and U18088 (N_18088,N_17889,N_17996);
xnor U18089 (N_18089,N_17794,N_17450);
or U18090 (N_18090,N_17742,N_17688);
nand U18091 (N_18091,N_17843,N_17797);
nand U18092 (N_18092,N_17127,N_17642);
nor U18093 (N_18093,N_17501,N_17609);
and U18094 (N_18094,N_17371,N_17598);
nand U18095 (N_18095,N_17604,N_17186);
nor U18096 (N_18096,N_17387,N_17449);
nand U18097 (N_18097,N_17426,N_17633);
nand U18098 (N_18098,N_17800,N_17695);
or U18099 (N_18099,N_17619,N_17084);
xor U18100 (N_18100,N_17599,N_17035);
and U18101 (N_18101,N_17749,N_17100);
xor U18102 (N_18102,N_17827,N_17217);
and U18103 (N_18103,N_17002,N_17218);
nand U18104 (N_18104,N_17311,N_17823);
xor U18105 (N_18105,N_17299,N_17748);
or U18106 (N_18106,N_17189,N_17578);
xor U18107 (N_18107,N_17561,N_17717);
or U18108 (N_18108,N_17286,N_17409);
nor U18109 (N_18109,N_17746,N_17795);
nand U18110 (N_18110,N_17270,N_17753);
xor U18111 (N_18111,N_17418,N_17281);
or U18112 (N_18112,N_17412,N_17970);
and U18113 (N_18113,N_17569,N_17814);
xnor U18114 (N_18114,N_17715,N_17919);
nand U18115 (N_18115,N_17665,N_17783);
or U18116 (N_18116,N_17771,N_17503);
nor U18117 (N_18117,N_17185,N_17691);
nor U18118 (N_18118,N_17597,N_17928);
nor U18119 (N_18119,N_17446,N_17768);
xnor U18120 (N_18120,N_17197,N_17980);
xnor U18121 (N_18121,N_17687,N_17130);
nand U18122 (N_18122,N_17038,N_17312);
or U18123 (N_18123,N_17354,N_17204);
xnor U18124 (N_18124,N_17815,N_17854);
nand U18125 (N_18125,N_17984,N_17405);
xnor U18126 (N_18126,N_17781,N_17659);
nand U18127 (N_18127,N_17240,N_17628);
xnor U18128 (N_18128,N_17958,N_17581);
nand U18129 (N_18129,N_17168,N_17882);
nand U18130 (N_18130,N_17828,N_17626);
or U18131 (N_18131,N_17401,N_17364);
nand U18132 (N_18132,N_17425,N_17481);
and U18133 (N_18133,N_17899,N_17095);
nand U18134 (N_18134,N_17145,N_17706);
or U18135 (N_18135,N_17773,N_17478);
and U18136 (N_18136,N_17662,N_17272);
and U18137 (N_18137,N_17923,N_17011);
or U18138 (N_18138,N_17638,N_17006);
xnor U18139 (N_18139,N_17661,N_17977);
and U18140 (N_18140,N_17676,N_17927);
nand U18141 (N_18141,N_17911,N_17871);
nand U18142 (N_18142,N_17786,N_17547);
or U18143 (N_18143,N_17063,N_17909);
xor U18144 (N_18144,N_17133,N_17410);
nor U18145 (N_18145,N_17269,N_17386);
and U18146 (N_18146,N_17720,N_17298);
nand U18147 (N_18147,N_17256,N_17976);
nand U18148 (N_18148,N_17654,N_17842);
nor U18149 (N_18149,N_17602,N_17398);
nand U18150 (N_18150,N_17319,N_17252);
nand U18151 (N_18151,N_17075,N_17735);
nand U18152 (N_18152,N_17845,N_17333);
nand U18153 (N_18153,N_17488,N_17457);
xor U18154 (N_18154,N_17621,N_17673);
nand U18155 (N_18155,N_17072,N_17942);
and U18156 (N_18156,N_17572,N_17689);
nand U18157 (N_18157,N_17852,N_17194);
nand U18158 (N_18158,N_17235,N_17166);
and U18159 (N_18159,N_17169,N_17683);
xor U18160 (N_18160,N_17739,N_17998);
or U18161 (N_18161,N_17632,N_17374);
nand U18162 (N_18162,N_17920,N_17061);
nor U18163 (N_18163,N_17044,N_17873);
xnor U18164 (N_18164,N_17881,N_17437);
nor U18165 (N_18165,N_17275,N_17564);
nand U18166 (N_18166,N_17556,N_17036);
xor U18167 (N_18167,N_17496,N_17907);
nor U18168 (N_18168,N_17708,N_17473);
xor U18169 (N_18169,N_17304,N_17975);
nand U18170 (N_18170,N_17951,N_17530);
nand U18171 (N_18171,N_17625,N_17028);
nand U18172 (N_18172,N_17898,N_17295);
nand U18173 (N_18173,N_17337,N_17073);
or U18174 (N_18174,N_17885,N_17509);
and U18175 (N_18175,N_17559,N_17901);
nand U18176 (N_18176,N_17963,N_17959);
and U18177 (N_18177,N_17914,N_17955);
nand U18178 (N_18178,N_17305,N_17801);
and U18179 (N_18179,N_17289,N_17165);
or U18180 (N_18180,N_17402,N_17593);
nand U18181 (N_18181,N_17519,N_17861);
xor U18182 (N_18182,N_17384,N_17931);
nand U18183 (N_18183,N_17191,N_17224);
nand U18184 (N_18184,N_17956,N_17042);
and U18185 (N_18185,N_17788,N_17394);
nor U18186 (N_18186,N_17151,N_17725);
nand U18187 (N_18187,N_17257,N_17356);
nand U18188 (N_18188,N_17202,N_17738);
nor U18189 (N_18189,N_17336,N_17316);
nand U18190 (N_18190,N_17974,N_17682);
or U18191 (N_18191,N_17325,N_17486);
and U18192 (N_18192,N_17641,N_17728);
or U18193 (N_18193,N_17290,N_17362);
or U18194 (N_18194,N_17156,N_17447);
xor U18195 (N_18195,N_17536,N_17701);
or U18196 (N_18196,N_17428,N_17056);
and U18197 (N_18197,N_17315,N_17962);
and U18198 (N_18198,N_17306,N_17125);
or U18199 (N_18199,N_17833,N_17769);
nand U18200 (N_18200,N_17147,N_17294);
nand U18201 (N_18201,N_17518,N_17656);
or U18202 (N_18202,N_17214,N_17106);
nand U18203 (N_18203,N_17560,N_17533);
nand U18204 (N_18204,N_17666,N_17181);
or U18205 (N_18205,N_17903,N_17973);
nand U18206 (N_18206,N_17892,N_17030);
nand U18207 (N_18207,N_17444,N_17966);
nor U18208 (N_18208,N_17588,N_17894);
xnor U18209 (N_18209,N_17663,N_17243);
nand U18210 (N_18210,N_17751,N_17328);
nor U18211 (N_18211,N_17089,N_17639);
nand U18212 (N_18212,N_17538,N_17069);
and U18213 (N_18213,N_17423,N_17373);
xnor U18214 (N_18214,N_17029,N_17101);
or U18215 (N_18215,N_17992,N_17378);
xnor U18216 (N_18216,N_17205,N_17195);
nor U18217 (N_18217,N_17022,N_17432);
and U18218 (N_18218,N_17025,N_17714);
and U18219 (N_18219,N_17945,N_17610);
nand U18220 (N_18220,N_17913,N_17711);
nor U18221 (N_18221,N_17731,N_17438);
nor U18222 (N_18222,N_17452,N_17055);
nand U18223 (N_18223,N_17821,N_17453);
or U18224 (N_18224,N_17138,N_17805);
and U18225 (N_18225,N_17902,N_17497);
or U18226 (N_18226,N_17136,N_17732);
or U18227 (N_18227,N_17210,N_17228);
nor U18228 (N_18228,N_17120,N_17613);
and U18229 (N_18229,N_17227,N_17464);
and U18230 (N_18230,N_17829,N_17471);
and U18231 (N_18231,N_17196,N_17239);
and U18232 (N_18232,N_17590,N_17826);
and U18233 (N_18233,N_17745,N_17868);
nand U18234 (N_18234,N_17981,N_17225);
nand U18235 (N_18235,N_17142,N_17989);
xnor U18236 (N_18236,N_17417,N_17046);
nor U18237 (N_18237,N_17813,N_17411);
and U18238 (N_18238,N_17772,N_17922);
and U18239 (N_18239,N_17877,N_17937);
or U18240 (N_18240,N_17515,N_17148);
and U18241 (N_18241,N_17987,N_17493);
nand U18242 (N_18242,N_17921,N_17361);
nor U18243 (N_18243,N_17104,N_17660);
or U18244 (N_18244,N_17511,N_17692);
nor U18245 (N_18245,N_17128,N_17229);
xnor U18246 (N_18246,N_17340,N_17607);
nand U18247 (N_18247,N_17934,N_17929);
xnor U18248 (N_18248,N_17505,N_17161);
xor U18249 (N_18249,N_17347,N_17825);
nand U18250 (N_18250,N_17775,N_17469);
xor U18251 (N_18251,N_17900,N_17693);
xnor U18252 (N_18252,N_17279,N_17009);
and U18253 (N_18253,N_17370,N_17117);
and U18254 (N_18254,N_17119,N_17953);
and U18255 (N_18255,N_17575,N_17777);
xor U18256 (N_18256,N_17152,N_17074);
nor U18257 (N_18257,N_17137,N_17936);
and U18258 (N_18258,N_17237,N_17650);
nor U18259 (N_18259,N_17329,N_17122);
nand U18260 (N_18260,N_17076,N_17589);
and U18261 (N_18261,N_17222,N_17375);
nor U18262 (N_18262,N_17032,N_17792);
or U18263 (N_18263,N_17517,N_17950);
and U18264 (N_18264,N_17259,N_17635);
and U18265 (N_18265,N_17524,N_17470);
xor U18266 (N_18266,N_17537,N_17472);
and U18267 (N_18267,N_17355,N_17727);
and U18268 (N_18268,N_17461,N_17040);
nand U18269 (N_18269,N_17502,N_17574);
nor U18270 (N_18270,N_17184,N_17455);
nand U18271 (N_18271,N_17352,N_17880);
and U18272 (N_18272,N_17835,N_17573);
and U18273 (N_18273,N_17761,N_17182);
xor U18274 (N_18274,N_17458,N_17059);
or U18275 (N_18275,N_17297,N_17349);
and U18276 (N_18276,N_17313,N_17162);
and U18277 (N_18277,N_17837,N_17710);
xor U18278 (N_18278,N_17467,N_17132);
and U18279 (N_18279,N_17924,N_17144);
and U18280 (N_18280,N_17796,N_17812);
nand U18281 (N_18281,N_17677,N_17415);
nand U18282 (N_18282,N_17484,N_17413);
and U18283 (N_18283,N_17954,N_17649);
nor U18284 (N_18284,N_17912,N_17740);
or U18285 (N_18285,N_17065,N_17555);
xor U18286 (N_18286,N_17764,N_17480);
xor U18287 (N_18287,N_17915,N_17752);
nor U18288 (N_18288,N_17414,N_17798);
nor U18289 (N_18289,N_17465,N_17348);
or U18290 (N_18290,N_17696,N_17188);
xnor U18291 (N_18291,N_17856,N_17192);
and U18292 (N_18292,N_17993,N_17407);
xor U18293 (N_18293,N_17960,N_17668);
nand U18294 (N_18294,N_17849,N_17278);
xor U18295 (N_18295,N_17321,N_17858);
and U18296 (N_18296,N_17791,N_17508);
nand U18297 (N_18297,N_17571,N_17140);
xnor U18298 (N_18298,N_17608,N_17804);
nor U18299 (N_18299,N_17718,N_17540);
nor U18300 (N_18300,N_17200,N_17969);
and U18301 (N_18301,N_17004,N_17291);
and U18302 (N_18302,N_17338,N_17645);
xor U18303 (N_18303,N_17332,N_17707);
nand U18304 (N_18304,N_17674,N_17087);
nand U18305 (N_18305,N_17723,N_17624);
or U18306 (N_18306,N_17603,N_17383);
or U18307 (N_18307,N_17857,N_17614);
xor U18308 (N_18308,N_17254,N_17251);
nor U18309 (N_18309,N_17341,N_17392);
xnor U18310 (N_18310,N_17379,N_17238);
xor U18311 (N_18311,N_17932,N_17351);
nand U18312 (N_18312,N_17118,N_17226);
nor U18313 (N_18313,N_17700,N_17212);
or U18314 (N_18314,N_17187,N_17039);
or U18315 (N_18315,N_17015,N_17554);
nor U18316 (N_18316,N_17521,N_17784);
nor U18317 (N_18317,N_17043,N_17543);
and U18318 (N_18318,N_17760,N_17462);
and U18319 (N_18319,N_17774,N_17108);
nor U18320 (N_18320,N_17612,N_17234);
xnor U18321 (N_18321,N_17099,N_17531);
nand U18322 (N_18322,N_17460,N_17780);
nand U18323 (N_18323,N_17283,N_17553);
and U18324 (N_18324,N_17793,N_17331);
nand U18325 (N_18325,N_17435,N_17762);
nand U18326 (N_18326,N_17091,N_17557);
xnor U18327 (N_18327,N_17083,N_17390);
or U18328 (N_18328,N_17114,N_17178);
nor U18329 (N_18329,N_17180,N_17672);
or U18330 (N_18330,N_17408,N_17595);
and U18331 (N_18331,N_17811,N_17680);
nor U18332 (N_18332,N_17600,N_17926);
and U18333 (N_18333,N_17019,N_17018);
nor U18334 (N_18334,N_17558,N_17391);
nor U18335 (N_18335,N_17618,N_17655);
and U18336 (N_18336,N_17657,N_17388);
nor U18337 (N_18337,N_17241,N_17121);
and U18338 (N_18338,N_17324,N_17658);
nand U18339 (N_18339,N_17053,N_17562);
nor U18340 (N_18340,N_17406,N_17077);
and U18341 (N_18341,N_17622,N_17605);
xnor U18342 (N_18342,N_17897,N_17171);
xnor U18343 (N_18343,N_17433,N_17806);
or U18344 (N_18344,N_17248,N_17381);
nand U18345 (N_18345,N_17123,N_17264);
nor U18346 (N_18346,N_17770,N_17062);
and U18347 (N_18347,N_17277,N_17369);
nand U18348 (N_18348,N_17377,N_17307);
nor U18349 (N_18349,N_17081,N_17334);
nand U18350 (N_18350,N_17047,N_17995);
xor U18351 (N_18351,N_17818,N_17982);
and U18352 (N_18352,N_17093,N_17579);
or U18353 (N_18353,N_17459,N_17016);
nor U18354 (N_18354,N_17096,N_17840);
and U18355 (N_18355,N_17159,N_17716);
and U18356 (N_18356,N_17203,N_17694);
xnor U18357 (N_18357,N_17640,N_17879);
or U18358 (N_18358,N_17454,N_17906);
nand U18359 (N_18359,N_17422,N_17726);
and U18360 (N_18360,N_17317,N_17757);
nand U18361 (N_18361,N_17568,N_17637);
xnor U18362 (N_18362,N_17506,N_17644);
nor U18363 (N_18363,N_17719,N_17207);
xnor U18364 (N_18364,N_17949,N_17870);
nor U18365 (N_18365,N_17935,N_17078);
and U18366 (N_18366,N_17385,N_17917);
xnor U18367 (N_18367,N_17847,N_17623);
nand U18368 (N_18368,N_17585,N_17669);
nor U18369 (N_18369,N_17071,N_17045);
and U18370 (N_18370,N_17747,N_17468);
xor U18371 (N_18371,N_17546,N_17482);
nand U18372 (N_18372,N_17451,N_17023);
or U18373 (N_18373,N_17008,N_17048);
or U18374 (N_18374,N_17862,N_17697);
and U18375 (N_18375,N_17905,N_17309);
or U18376 (N_18376,N_17634,N_17865);
xor U18377 (N_18377,N_17580,N_17785);
and U18378 (N_18378,N_17516,N_17991);
nand U18379 (N_18379,N_17343,N_17592);
or U18380 (N_18380,N_17759,N_17790);
or U18381 (N_18381,N_17209,N_17787);
nor U18382 (N_18382,N_17323,N_17442);
nor U18383 (N_18383,N_17041,N_17111);
and U18384 (N_18384,N_17170,N_17288);
or U18385 (N_18385,N_17419,N_17594);
nand U18386 (N_18386,N_17326,N_17591);
nor U18387 (N_18387,N_17737,N_17596);
nand U18388 (N_18388,N_17420,N_17647);
and U18389 (N_18389,N_17236,N_17273);
or U18390 (N_18390,N_17587,N_17427);
nand U18391 (N_18391,N_17436,N_17491);
or U18392 (N_18392,N_17730,N_17544);
or U18393 (N_18393,N_17526,N_17577);
nand U18394 (N_18394,N_17925,N_17330);
and U18395 (N_18395,N_17146,N_17322);
xnor U18396 (N_18396,N_17878,N_17939);
nand U18397 (N_18397,N_17755,N_17365);
nor U18398 (N_18398,N_17495,N_17513);
and U18399 (N_18399,N_17001,N_17284);
xnor U18400 (N_18400,N_17810,N_17615);
nor U18401 (N_18401,N_17853,N_17750);
or U18402 (N_18402,N_17193,N_17102);
nor U18403 (N_18403,N_17895,N_17838);
nor U18404 (N_18404,N_17910,N_17097);
or U18405 (N_18405,N_17223,N_17916);
nand U18406 (N_18406,N_17522,N_17946);
and U18407 (N_18407,N_17690,N_17155);
or U18408 (N_18408,N_17864,N_17158);
nor U18409 (N_18409,N_17262,N_17215);
nor U18410 (N_18410,N_17586,N_17068);
or U18411 (N_18411,N_17883,N_17020);
and U18412 (N_18412,N_17049,N_17646);
nor U18413 (N_18413,N_17216,N_17876);
or U18414 (N_18414,N_17507,N_17848);
or U18415 (N_18415,N_17510,N_17767);
xnor U18416 (N_18416,N_17206,N_17891);
and U18417 (N_18417,N_17163,N_17994);
xnor U18418 (N_18418,N_17860,N_17160);
nand U18419 (N_18419,N_17088,N_17636);
xor U18420 (N_18420,N_17395,N_17124);
or U18421 (N_18421,N_17231,N_17255);
xor U18422 (N_18422,N_17335,N_17802);
nand U18423 (N_18423,N_17389,N_17443);
xor U18424 (N_18424,N_17031,N_17866);
and U18425 (N_18425,N_17363,N_17474);
nand U18426 (N_18426,N_17552,N_17943);
nand U18427 (N_18427,N_17948,N_17026);
xnor U18428 (N_18428,N_17713,N_17198);
nor U18429 (N_18429,N_17282,N_17149);
nand U18430 (N_18430,N_17380,N_17551);
or U18431 (N_18431,N_17441,N_17930);
nand U18432 (N_18432,N_17475,N_17064);
xor U18433 (N_18433,N_17177,N_17172);
nor U18434 (N_18434,N_17893,N_17416);
and U18435 (N_18435,N_17110,N_17841);
or U18436 (N_18436,N_17135,N_17400);
or U18437 (N_18437,N_17115,N_17246);
xnor U18438 (N_18438,N_17403,N_17652);
or U18439 (N_18439,N_17839,N_17629);
or U18440 (N_18440,N_17971,N_17382);
nor U18441 (N_18441,N_17027,N_17000);
and U18442 (N_18442,N_17630,N_17220);
nor U18443 (N_18443,N_17836,N_17271);
or U18444 (N_18444,N_17244,N_17938);
xor U18445 (N_18445,N_17933,N_17489);
or U18446 (N_18446,N_17643,N_17476);
and U18447 (N_18447,N_17678,N_17366);
nor U18448 (N_18448,N_17583,N_17648);
or U18449 (N_18449,N_17620,N_17733);
xor U18450 (N_18450,N_17017,N_17007);
nor U18451 (N_18451,N_17940,N_17888);
or U18452 (N_18452,N_17808,N_17961);
or U18453 (N_18453,N_17500,N_17230);
or U18454 (N_18454,N_17765,N_17052);
nor U18455 (N_18455,N_17545,N_17529);
or U18456 (N_18456,N_17985,N_17431);
and U18457 (N_18457,N_17872,N_17221);
and U18458 (N_18458,N_17721,N_17034);
nand U18459 (N_18459,N_17167,N_17310);
or U18460 (N_18460,N_17941,N_17816);
xnor U18461 (N_18461,N_17359,N_17566);
and U18462 (N_18462,N_17263,N_17890);
nor U18463 (N_18463,N_17067,N_17245);
or U18464 (N_18464,N_17679,N_17208);
nor U18465 (N_18465,N_17887,N_17539);
nor U18466 (N_18466,N_17054,N_17320);
nor U18467 (N_18467,N_17820,N_17651);
or U18468 (N_18468,N_17863,N_17302);
nor U18469 (N_18469,N_17675,N_17831);
nand U18470 (N_18470,N_17183,N_17376);
nand U18471 (N_18471,N_17350,N_17699);
nand U18472 (N_18472,N_17709,N_17233);
nand U18473 (N_18473,N_17393,N_17265);
nor U18474 (N_18474,N_17908,N_17527);
nor U18475 (N_18475,N_17729,N_17082);
and U18476 (N_18476,N_17512,N_17013);
nand U18477 (N_18477,N_17824,N_17606);
and U18478 (N_18478,N_17466,N_17260);
nand U18479 (N_18479,N_17944,N_17107);
and U18480 (N_18480,N_17712,N_17430);
nand U18481 (N_18481,N_17357,N_17758);
nor U18482 (N_18482,N_17126,N_17367);
and U18483 (N_18483,N_17339,N_17799);
and U18484 (N_18484,N_17285,N_17817);
or U18485 (N_18485,N_17685,N_17213);
xor U18486 (N_18486,N_17616,N_17582);
xor U18487 (N_18487,N_17247,N_17066);
or U18488 (N_18488,N_17300,N_17565);
xnor U18489 (N_18489,N_17131,N_17549);
or U18490 (N_18490,N_17776,N_17175);
or U18491 (N_18491,N_17060,N_17396);
and U18492 (N_18492,N_17037,N_17705);
nor U18493 (N_18493,N_17199,N_17440);
or U18494 (N_18494,N_17342,N_17358);
and U18495 (N_18495,N_17563,N_17368);
nor U18496 (N_18496,N_17492,N_17268);
and U18497 (N_18497,N_17550,N_17109);
nor U18498 (N_18498,N_17684,N_17327);
nand U18499 (N_18499,N_17722,N_17584);
xnor U18500 (N_18500,N_17367,N_17062);
nand U18501 (N_18501,N_17567,N_17970);
or U18502 (N_18502,N_17594,N_17951);
and U18503 (N_18503,N_17129,N_17687);
nand U18504 (N_18504,N_17650,N_17477);
or U18505 (N_18505,N_17285,N_17101);
nor U18506 (N_18506,N_17475,N_17827);
and U18507 (N_18507,N_17790,N_17055);
nand U18508 (N_18508,N_17922,N_17176);
xnor U18509 (N_18509,N_17841,N_17566);
or U18510 (N_18510,N_17256,N_17449);
nand U18511 (N_18511,N_17904,N_17561);
nor U18512 (N_18512,N_17895,N_17059);
or U18513 (N_18513,N_17187,N_17631);
and U18514 (N_18514,N_17867,N_17123);
nor U18515 (N_18515,N_17529,N_17947);
or U18516 (N_18516,N_17845,N_17081);
xnor U18517 (N_18517,N_17473,N_17535);
or U18518 (N_18518,N_17319,N_17663);
nor U18519 (N_18519,N_17762,N_17699);
nor U18520 (N_18520,N_17760,N_17334);
xor U18521 (N_18521,N_17340,N_17202);
and U18522 (N_18522,N_17843,N_17492);
xnor U18523 (N_18523,N_17478,N_17954);
nand U18524 (N_18524,N_17096,N_17508);
xor U18525 (N_18525,N_17909,N_17551);
xor U18526 (N_18526,N_17039,N_17767);
xnor U18527 (N_18527,N_17858,N_17788);
xnor U18528 (N_18528,N_17628,N_17001);
xnor U18529 (N_18529,N_17050,N_17602);
nand U18530 (N_18530,N_17805,N_17479);
nand U18531 (N_18531,N_17406,N_17316);
nand U18532 (N_18532,N_17262,N_17323);
nand U18533 (N_18533,N_17104,N_17670);
or U18534 (N_18534,N_17905,N_17178);
xor U18535 (N_18535,N_17851,N_17449);
nand U18536 (N_18536,N_17704,N_17412);
or U18537 (N_18537,N_17660,N_17251);
nor U18538 (N_18538,N_17826,N_17064);
and U18539 (N_18539,N_17461,N_17762);
and U18540 (N_18540,N_17322,N_17046);
nor U18541 (N_18541,N_17080,N_17429);
nor U18542 (N_18542,N_17320,N_17072);
nor U18543 (N_18543,N_17866,N_17375);
or U18544 (N_18544,N_17685,N_17922);
xor U18545 (N_18545,N_17813,N_17041);
nand U18546 (N_18546,N_17155,N_17689);
or U18547 (N_18547,N_17267,N_17066);
and U18548 (N_18548,N_17910,N_17872);
and U18549 (N_18549,N_17287,N_17563);
xor U18550 (N_18550,N_17118,N_17817);
nor U18551 (N_18551,N_17969,N_17889);
xor U18552 (N_18552,N_17505,N_17654);
xor U18553 (N_18553,N_17919,N_17942);
xor U18554 (N_18554,N_17145,N_17754);
or U18555 (N_18555,N_17004,N_17997);
nand U18556 (N_18556,N_17947,N_17003);
or U18557 (N_18557,N_17197,N_17728);
and U18558 (N_18558,N_17144,N_17680);
nor U18559 (N_18559,N_17239,N_17366);
and U18560 (N_18560,N_17384,N_17395);
or U18561 (N_18561,N_17121,N_17609);
and U18562 (N_18562,N_17751,N_17423);
xor U18563 (N_18563,N_17652,N_17492);
nand U18564 (N_18564,N_17803,N_17473);
and U18565 (N_18565,N_17315,N_17560);
or U18566 (N_18566,N_17765,N_17413);
nor U18567 (N_18567,N_17255,N_17658);
and U18568 (N_18568,N_17761,N_17766);
or U18569 (N_18569,N_17742,N_17815);
and U18570 (N_18570,N_17535,N_17560);
nand U18571 (N_18571,N_17432,N_17510);
and U18572 (N_18572,N_17375,N_17374);
xnor U18573 (N_18573,N_17253,N_17322);
nor U18574 (N_18574,N_17531,N_17007);
or U18575 (N_18575,N_17199,N_17354);
nand U18576 (N_18576,N_17332,N_17593);
nor U18577 (N_18577,N_17369,N_17872);
nor U18578 (N_18578,N_17185,N_17733);
and U18579 (N_18579,N_17195,N_17042);
nand U18580 (N_18580,N_17241,N_17332);
nor U18581 (N_18581,N_17631,N_17455);
nor U18582 (N_18582,N_17817,N_17166);
or U18583 (N_18583,N_17997,N_17443);
nor U18584 (N_18584,N_17858,N_17099);
nand U18585 (N_18585,N_17561,N_17311);
nor U18586 (N_18586,N_17917,N_17288);
or U18587 (N_18587,N_17178,N_17642);
xnor U18588 (N_18588,N_17290,N_17191);
and U18589 (N_18589,N_17834,N_17395);
nand U18590 (N_18590,N_17253,N_17517);
xor U18591 (N_18591,N_17578,N_17210);
or U18592 (N_18592,N_17079,N_17814);
nor U18593 (N_18593,N_17863,N_17604);
nand U18594 (N_18594,N_17122,N_17579);
xnor U18595 (N_18595,N_17791,N_17064);
nor U18596 (N_18596,N_17329,N_17012);
and U18597 (N_18597,N_17557,N_17499);
nor U18598 (N_18598,N_17376,N_17795);
or U18599 (N_18599,N_17387,N_17637);
and U18600 (N_18600,N_17506,N_17576);
nand U18601 (N_18601,N_17041,N_17628);
and U18602 (N_18602,N_17167,N_17654);
or U18603 (N_18603,N_17063,N_17430);
or U18604 (N_18604,N_17749,N_17579);
or U18605 (N_18605,N_17974,N_17732);
xor U18606 (N_18606,N_17421,N_17451);
nand U18607 (N_18607,N_17485,N_17114);
nor U18608 (N_18608,N_17521,N_17006);
xnor U18609 (N_18609,N_17778,N_17972);
or U18610 (N_18610,N_17244,N_17942);
or U18611 (N_18611,N_17185,N_17135);
xor U18612 (N_18612,N_17949,N_17892);
and U18613 (N_18613,N_17455,N_17813);
or U18614 (N_18614,N_17278,N_17966);
nor U18615 (N_18615,N_17673,N_17777);
xor U18616 (N_18616,N_17073,N_17254);
or U18617 (N_18617,N_17512,N_17718);
and U18618 (N_18618,N_17446,N_17620);
or U18619 (N_18619,N_17738,N_17238);
nor U18620 (N_18620,N_17766,N_17914);
nand U18621 (N_18621,N_17595,N_17910);
or U18622 (N_18622,N_17603,N_17578);
xnor U18623 (N_18623,N_17967,N_17201);
xor U18624 (N_18624,N_17299,N_17908);
nand U18625 (N_18625,N_17250,N_17104);
and U18626 (N_18626,N_17608,N_17769);
nor U18627 (N_18627,N_17616,N_17654);
nor U18628 (N_18628,N_17519,N_17089);
nor U18629 (N_18629,N_17902,N_17250);
or U18630 (N_18630,N_17740,N_17261);
or U18631 (N_18631,N_17496,N_17992);
xnor U18632 (N_18632,N_17794,N_17906);
and U18633 (N_18633,N_17850,N_17290);
xnor U18634 (N_18634,N_17544,N_17336);
xor U18635 (N_18635,N_17197,N_17554);
nor U18636 (N_18636,N_17434,N_17922);
or U18637 (N_18637,N_17325,N_17561);
or U18638 (N_18638,N_17129,N_17390);
and U18639 (N_18639,N_17795,N_17720);
nor U18640 (N_18640,N_17512,N_17270);
nor U18641 (N_18641,N_17060,N_17649);
nor U18642 (N_18642,N_17625,N_17262);
or U18643 (N_18643,N_17425,N_17050);
and U18644 (N_18644,N_17327,N_17899);
xnor U18645 (N_18645,N_17092,N_17901);
and U18646 (N_18646,N_17227,N_17248);
and U18647 (N_18647,N_17357,N_17417);
and U18648 (N_18648,N_17875,N_17945);
xor U18649 (N_18649,N_17956,N_17878);
or U18650 (N_18650,N_17936,N_17410);
xnor U18651 (N_18651,N_17150,N_17607);
nand U18652 (N_18652,N_17585,N_17664);
xor U18653 (N_18653,N_17663,N_17958);
and U18654 (N_18654,N_17662,N_17781);
and U18655 (N_18655,N_17101,N_17038);
nand U18656 (N_18656,N_17148,N_17465);
xnor U18657 (N_18657,N_17799,N_17326);
xor U18658 (N_18658,N_17739,N_17064);
nor U18659 (N_18659,N_17768,N_17856);
nand U18660 (N_18660,N_17963,N_17742);
nand U18661 (N_18661,N_17334,N_17452);
and U18662 (N_18662,N_17108,N_17601);
and U18663 (N_18663,N_17946,N_17202);
nand U18664 (N_18664,N_17666,N_17922);
nor U18665 (N_18665,N_17741,N_17949);
nand U18666 (N_18666,N_17536,N_17417);
xnor U18667 (N_18667,N_17021,N_17127);
xnor U18668 (N_18668,N_17639,N_17027);
nand U18669 (N_18669,N_17582,N_17990);
or U18670 (N_18670,N_17466,N_17918);
and U18671 (N_18671,N_17370,N_17615);
nor U18672 (N_18672,N_17283,N_17748);
and U18673 (N_18673,N_17243,N_17251);
nor U18674 (N_18674,N_17398,N_17744);
and U18675 (N_18675,N_17521,N_17165);
and U18676 (N_18676,N_17674,N_17585);
xnor U18677 (N_18677,N_17683,N_17498);
nor U18678 (N_18678,N_17699,N_17169);
nand U18679 (N_18679,N_17288,N_17776);
and U18680 (N_18680,N_17354,N_17069);
and U18681 (N_18681,N_17074,N_17466);
nand U18682 (N_18682,N_17550,N_17612);
and U18683 (N_18683,N_17967,N_17327);
nor U18684 (N_18684,N_17127,N_17631);
nand U18685 (N_18685,N_17399,N_17160);
and U18686 (N_18686,N_17712,N_17530);
xnor U18687 (N_18687,N_17878,N_17760);
or U18688 (N_18688,N_17338,N_17066);
and U18689 (N_18689,N_17864,N_17148);
and U18690 (N_18690,N_17765,N_17823);
or U18691 (N_18691,N_17358,N_17181);
and U18692 (N_18692,N_17194,N_17373);
or U18693 (N_18693,N_17320,N_17548);
xnor U18694 (N_18694,N_17077,N_17565);
xnor U18695 (N_18695,N_17888,N_17229);
and U18696 (N_18696,N_17005,N_17873);
xor U18697 (N_18697,N_17360,N_17897);
and U18698 (N_18698,N_17684,N_17200);
and U18699 (N_18699,N_17174,N_17501);
nand U18700 (N_18700,N_17905,N_17429);
xnor U18701 (N_18701,N_17482,N_17342);
nand U18702 (N_18702,N_17355,N_17053);
nor U18703 (N_18703,N_17681,N_17499);
nor U18704 (N_18704,N_17207,N_17078);
xnor U18705 (N_18705,N_17518,N_17793);
xor U18706 (N_18706,N_17620,N_17626);
nand U18707 (N_18707,N_17479,N_17503);
or U18708 (N_18708,N_17039,N_17399);
and U18709 (N_18709,N_17186,N_17029);
xor U18710 (N_18710,N_17435,N_17939);
or U18711 (N_18711,N_17259,N_17720);
or U18712 (N_18712,N_17276,N_17729);
nand U18713 (N_18713,N_17221,N_17737);
nand U18714 (N_18714,N_17165,N_17648);
and U18715 (N_18715,N_17958,N_17939);
nor U18716 (N_18716,N_17397,N_17359);
xnor U18717 (N_18717,N_17195,N_17561);
nand U18718 (N_18718,N_17984,N_17941);
nand U18719 (N_18719,N_17769,N_17345);
nor U18720 (N_18720,N_17838,N_17271);
or U18721 (N_18721,N_17244,N_17211);
and U18722 (N_18722,N_17209,N_17329);
nor U18723 (N_18723,N_17767,N_17165);
nor U18724 (N_18724,N_17114,N_17788);
nor U18725 (N_18725,N_17732,N_17400);
nand U18726 (N_18726,N_17527,N_17064);
and U18727 (N_18727,N_17380,N_17401);
nor U18728 (N_18728,N_17795,N_17305);
or U18729 (N_18729,N_17071,N_17453);
and U18730 (N_18730,N_17643,N_17291);
nand U18731 (N_18731,N_17863,N_17193);
nand U18732 (N_18732,N_17199,N_17788);
or U18733 (N_18733,N_17695,N_17685);
xnor U18734 (N_18734,N_17586,N_17090);
and U18735 (N_18735,N_17742,N_17263);
nand U18736 (N_18736,N_17644,N_17397);
nand U18737 (N_18737,N_17676,N_17524);
and U18738 (N_18738,N_17183,N_17192);
nand U18739 (N_18739,N_17942,N_17022);
or U18740 (N_18740,N_17254,N_17371);
nor U18741 (N_18741,N_17950,N_17253);
and U18742 (N_18742,N_17969,N_17931);
nor U18743 (N_18743,N_17691,N_17600);
nor U18744 (N_18744,N_17780,N_17164);
or U18745 (N_18745,N_17771,N_17219);
nand U18746 (N_18746,N_17524,N_17901);
xor U18747 (N_18747,N_17145,N_17892);
and U18748 (N_18748,N_17398,N_17919);
and U18749 (N_18749,N_17146,N_17982);
or U18750 (N_18750,N_17661,N_17140);
and U18751 (N_18751,N_17380,N_17211);
xor U18752 (N_18752,N_17572,N_17987);
and U18753 (N_18753,N_17192,N_17607);
or U18754 (N_18754,N_17001,N_17320);
nor U18755 (N_18755,N_17261,N_17983);
nor U18756 (N_18756,N_17910,N_17339);
xnor U18757 (N_18757,N_17649,N_17582);
nand U18758 (N_18758,N_17961,N_17119);
and U18759 (N_18759,N_17787,N_17025);
xor U18760 (N_18760,N_17356,N_17443);
xor U18761 (N_18761,N_17250,N_17571);
nor U18762 (N_18762,N_17292,N_17065);
nor U18763 (N_18763,N_17679,N_17647);
and U18764 (N_18764,N_17899,N_17049);
nor U18765 (N_18765,N_17539,N_17477);
or U18766 (N_18766,N_17082,N_17848);
nor U18767 (N_18767,N_17088,N_17262);
nor U18768 (N_18768,N_17455,N_17689);
or U18769 (N_18769,N_17683,N_17752);
nand U18770 (N_18770,N_17766,N_17306);
nor U18771 (N_18771,N_17918,N_17894);
or U18772 (N_18772,N_17281,N_17884);
or U18773 (N_18773,N_17847,N_17705);
xor U18774 (N_18774,N_17189,N_17020);
nand U18775 (N_18775,N_17614,N_17191);
nand U18776 (N_18776,N_17473,N_17415);
nand U18777 (N_18777,N_17107,N_17952);
and U18778 (N_18778,N_17360,N_17446);
and U18779 (N_18779,N_17068,N_17183);
or U18780 (N_18780,N_17108,N_17161);
nor U18781 (N_18781,N_17777,N_17795);
or U18782 (N_18782,N_17717,N_17627);
or U18783 (N_18783,N_17732,N_17833);
and U18784 (N_18784,N_17183,N_17542);
or U18785 (N_18785,N_17750,N_17084);
xor U18786 (N_18786,N_17885,N_17014);
nor U18787 (N_18787,N_17809,N_17183);
nor U18788 (N_18788,N_17210,N_17850);
nor U18789 (N_18789,N_17184,N_17604);
nand U18790 (N_18790,N_17719,N_17530);
xnor U18791 (N_18791,N_17129,N_17957);
nor U18792 (N_18792,N_17166,N_17500);
nand U18793 (N_18793,N_17425,N_17981);
xnor U18794 (N_18794,N_17700,N_17131);
nand U18795 (N_18795,N_17082,N_17777);
nand U18796 (N_18796,N_17845,N_17485);
and U18797 (N_18797,N_17786,N_17834);
nand U18798 (N_18798,N_17109,N_17529);
nand U18799 (N_18799,N_17066,N_17243);
xnor U18800 (N_18800,N_17203,N_17480);
nor U18801 (N_18801,N_17685,N_17599);
nand U18802 (N_18802,N_17470,N_17260);
xor U18803 (N_18803,N_17499,N_17309);
or U18804 (N_18804,N_17795,N_17157);
nand U18805 (N_18805,N_17561,N_17401);
and U18806 (N_18806,N_17657,N_17062);
xnor U18807 (N_18807,N_17336,N_17153);
nor U18808 (N_18808,N_17186,N_17540);
nor U18809 (N_18809,N_17065,N_17423);
xor U18810 (N_18810,N_17775,N_17766);
or U18811 (N_18811,N_17853,N_17890);
and U18812 (N_18812,N_17149,N_17057);
and U18813 (N_18813,N_17511,N_17891);
xor U18814 (N_18814,N_17144,N_17341);
nor U18815 (N_18815,N_17081,N_17898);
nand U18816 (N_18816,N_17065,N_17950);
nand U18817 (N_18817,N_17023,N_17520);
nor U18818 (N_18818,N_17719,N_17700);
nand U18819 (N_18819,N_17187,N_17706);
nand U18820 (N_18820,N_17826,N_17495);
or U18821 (N_18821,N_17844,N_17120);
nand U18822 (N_18822,N_17461,N_17979);
nand U18823 (N_18823,N_17133,N_17613);
nor U18824 (N_18824,N_17937,N_17215);
nor U18825 (N_18825,N_17867,N_17869);
nand U18826 (N_18826,N_17590,N_17721);
nor U18827 (N_18827,N_17866,N_17935);
xnor U18828 (N_18828,N_17960,N_17904);
or U18829 (N_18829,N_17860,N_17690);
or U18830 (N_18830,N_17828,N_17383);
nor U18831 (N_18831,N_17245,N_17394);
and U18832 (N_18832,N_17597,N_17250);
nand U18833 (N_18833,N_17898,N_17902);
or U18834 (N_18834,N_17239,N_17120);
nand U18835 (N_18835,N_17067,N_17395);
xnor U18836 (N_18836,N_17110,N_17028);
nor U18837 (N_18837,N_17137,N_17276);
and U18838 (N_18838,N_17322,N_17873);
nor U18839 (N_18839,N_17713,N_17138);
and U18840 (N_18840,N_17726,N_17361);
xor U18841 (N_18841,N_17818,N_17573);
or U18842 (N_18842,N_17834,N_17459);
and U18843 (N_18843,N_17406,N_17510);
nor U18844 (N_18844,N_17580,N_17684);
xor U18845 (N_18845,N_17658,N_17712);
and U18846 (N_18846,N_17957,N_17214);
nand U18847 (N_18847,N_17169,N_17434);
nand U18848 (N_18848,N_17702,N_17840);
xor U18849 (N_18849,N_17679,N_17126);
xnor U18850 (N_18850,N_17365,N_17936);
and U18851 (N_18851,N_17942,N_17269);
xnor U18852 (N_18852,N_17562,N_17541);
nor U18853 (N_18853,N_17697,N_17578);
or U18854 (N_18854,N_17369,N_17362);
nand U18855 (N_18855,N_17307,N_17684);
nand U18856 (N_18856,N_17898,N_17649);
or U18857 (N_18857,N_17001,N_17851);
or U18858 (N_18858,N_17194,N_17127);
and U18859 (N_18859,N_17587,N_17964);
and U18860 (N_18860,N_17371,N_17728);
xnor U18861 (N_18861,N_17760,N_17893);
nor U18862 (N_18862,N_17870,N_17449);
and U18863 (N_18863,N_17112,N_17811);
xnor U18864 (N_18864,N_17126,N_17055);
or U18865 (N_18865,N_17134,N_17475);
or U18866 (N_18866,N_17258,N_17340);
or U18867 (N_18867,N_17497,N_17528);
xnor U18868 (N_18868,N_17709,N_17528);
xnor U18869 (N_18869,N_17443,N_17780);
nor U18870 (N_18870,N_17807,N_17207);
nor U18871 (N_18871,N_17404,N_17277);
and U18872 (N_18872,N_17858,N_17228);
xnor U18873 (N_18873,N_17379,N_17140);
nand U18874 (N_18874,N_17682,N_17533);
xor U18875 (N_18875,N_17780,N_17338);
xnor U18876 (N_18876,N_17383,N_17752);
xor U18877 (N_18877,N_17051,N_17856);
or U18878 (N_18878,N_17109,N_17049);
and U18879 (N_18879,N_17899,N_17484);
and U18880 (N_18880,N_17937,N_17956);
nor U18881 (N_18881,N_17343,N_17384);
nor U18882 (N_18882,N_17104,N_17705);
and U18883 (N_18883,N_17353,N_17112);
nor U18884 (N_18884,N_17194,N_17714);
xor U18885 (N_18885,N_17140,N_17209);
and U18886 (N_18886,N_17106,N_17048);
nand U18887 (N_18887,N_17064,N_17568);
xnor U18888 (N_18888,N_17536,N_17740);
nor U18889 (N_18889,N_17519,N_17937);
nor U18890 (N_18890,N_17085,N_17274);
nor U18891 (N_18891,N_17801,N_17595);
nand U18892 (N_18892,N_17335,N_17029);
or U18893 (N_18893,N_17037,N_17762);
or U18894 (N_18894,N_17101,N_17363);
xnor U18895 (N_18895,N_17282,N_17878);
and U18896 (N_18896,N_17890,N_17375);
or U18897 (N_18897,N_17718,N_17701);
and U18898 (N_18898,N_17162,N_17020);
and U18899 (N_18899,N_17350,N_17599);
xor U18900 (N_18900,N_17943,N_17984);
or U18901 (N_18901,N_17917,N_17384);
or U18902 (N_18902,N_17025,N_17199);
xor U18903 (N_18903,N_17970,N_17816);
nand U18904 (N_18904,N_17043,N_17269);
xnor U18905 (N_18905,N_17089,N_17484);
and U18906 (N_18906,N_17922,N_17770);
nor U18907 (N_18907,N_17621,N_17763);
xnor U18908 (N_18908,N_17987,N_17510);
and U18909 (N_18909,N_17924,N_17415);
and U18910 (N_18910,N_17791,N_17746);
or U18911 (N_18911,N_17406,N_17632);
and U18912 (N_18912,N_17573,N_17209);
nand U18913 (N_18913,N_17766,N_17121);
xnor U18914 (N_18914,N_17595,N_17774);
nor U18915 (N_18915,N_17298,N_17524);
xor U18916 (N_18916,N_17603,N_17309);
or U18917 (N_18917,N_17165,N_17494);
and U18918 (N_18918,N_17024,N_17972);
nand U18919 (N_18919,N_17725,N_17076);
xor U18920 (N_18920,N_17290,N_17997);
and U18921 (N_18921,N_17177,N_17575);
xnor U18922 (N_18922,N_17529,N_17133);
or U18923 (N_18923,N_17694,N_17678);
nor U18924 (N_18924,N_17507,N_17675);
nor U18925 (N_18925,N_17122,N_17747);
and U18926 (N_18926,N_17262,N_17806);
xnor U18927 (N_18927,N_17343,N_17174);
xor U18928 (N_18928,N_17415,N_17664);
nor U18929 (N_18929,N_17091,N_17661);
xor U18930 (N_18930,N_17516,N_17877);
xor U18931 (N_18931,N_17204,N_17971);
xor U18932 (N_18932,N_17319,N_17321);
and U18933 (N_18933,N_17826,N_17308);
xnor U18934 (N_18934,N_17790,N_17842);
xor U18935 (N_18935,N_17141,N_17278);
or U18936 (N_18936,N_17920,N_17172);
nand U18937 (N_18937,N_17602,N_17191);
nand U18938 (N_18938,N_17992,N_17422);
nand U18939 (N_18939,N_17964,N_17981);
xnor U18940 (N_18940,N_17999,N_17763);
and U18941 (N_18941,N_17493,N_17475);
nor U18942 (N_18942,N_17113,N_17501);
nor U18943 (N_18943,N_17140,N_17282);
xnor U18944 (N_18944,N_17313,N_17697);
or U18945 (N_18945,N_17224,N_17479);
and U18946 (N_18946,N_17889,N_17314);
xor U18947 (N_18947,N_17236,N_17003);
xor U18948 (N_18948,N_17540,N_17319);
nand U18949 (N_18949,N_17805,N_17276);
nand U18950 (N_18950,N_17323,N_17740);
xnor U18951 (N_18951,N_17517,N_17257);
nand U18952 (N_18952,N_17804,N_17698);
and U18953 (N_18953,N_17136,N_17860);
xor U18954 (N_18954,N_17284,N_17536);
or U18955 (N_18955,N_17593,N_17976);
or U18956 (N_18956,N_17989,N_17194);
xnor U18957 (N_18957,N_17793,N_17379);
and U18958 (N_18958,N_17859,N_17283);
or U18959 (N_18959,N_17894,N_17718);
or U18960 (N_18960,N_17351,N_17713);
xnor U18961 (N_18961,N_17230,N_17446);
nor U18962 (N_18962,N_17128,N_17606);
xnor U18963 (N_18963,N_17330,N_17474);
xor U18964 (N_18964,N_17989,N_17274);
nor U18965 (N_18965,N_17881,N_17698);
nand U18966 (N_18966,N_17937,N_17601);
xnor U18967 (N_18967,N_17022,N_17351);
or U18968 (N_18968,N_17417,N_17116);
or U18969 (N_18969,N_17918,N_17374);
or U18970 (N_18970,N_17255,N_17396);
nand U18971 (N_18971,N_17932,N_17512);
or U18972 (N_18972,N_17129,N_17197);
nand U18973 (N_18973,N_17000,N_17429);
xnor U18974 (N_18974,N_17632,N_17675);
xor U18975 (N_18975,N_17351,N_17437);
nand U18976 (N_18976,N_17746,N_17368);
and U18977 (N_18977,N_17786,N_17650);
and U18978 (N_18978,N_17083,N_17002);
nor U18979 (N_18979,N_17278,N_17438);
nand U18980 (N_18980,N_17064,N_17134);
or U18981 (N_18981,N_17910,N_17565);
and U18982 (N_18982,N_17117,N_17085);
xnor U18983 (N_18983,N_17153,N_17834);
nand U18984 (N_18984,N_17573,N_17412);
or U18985 (N_18985,N_17024,N_17676);
and U18986 (N_18986,N_17968,N_17750);
and U18987 (N_18987,N_17272,N_17294);
nor U18988 (N_18988,N_17220,N_17517);
or U18989 (N_18989,N_17967,N_17552);
nand U18990 (N_18990,N_17463,N_17108);
or U18991 (N_18991,N_17331,N_17734);
or U18992 (N_18992,N_17410,N_17983);
and U18993 (N_18993,N_17641,N_17407);
nand U18994 (N_18994,N_17114,N_17935);
or U18995 (N_18995,N_17573,N_17612);
and U18996 (N_18996,N_17315,N_17343);
and U18997 (N_18997,N_17559,N_17627);
nand U18998 (N_18998,N_17174,N_17280);
nor U18999 (N_18999,N_17202,N_17891);
and U19000 (N_19000,N_18550,N_18283);
or U19001 (N_19001,N_18538,N_18435);
xor U19002 (N_19002,N_18328,N_18988);
or U19003 (N_19003,N_18629,N_18131);
nand U19004 (N_19004,N_18309,N_18513);
nor U19005 (N_19005,N_18395,N_18167);
and U19006 (N_19006,N_18020,N_18113);
nor U19007 (N_19007,N_18368,N_18168);
nor U19008 (N_19008,N_18519,N_18372);
or U19009 (N_19009,N_18024,N_18798);
nand U19010 (N_19010,N_18149,N_18455);
or U19011 (N_19011,N_18312,N_18674);
nand U19012 (N_19012,N_18363,N_18892);
or U19013 (N_19013,N_18802,N_18948);
nor U19014 (N_19014,N_18890,N_18402);
nand U19015 (N_19015,N_18597,N_18018);
and U19016 (N_19016,N_18457,N_18545);
or U19017 (N_19017,N_18710,N_18831);
and U19018 (N_19018,N_18045,N_18794);
xor U19019 (N_19019,N_18590,N_18684);
nor U19020 (N_19020,N_18301,N_18554);
nand U19021 (N_19021,N_18872,N_18733);
nand U19022 (N_19022,N_18007,N_18456);
or U19023 (N_19023,N_18420,N_18050);
xor U19024 (N_19024,N_18716,N_18370);
xnor U19025 (N_19025,N_18291,N_18496);
xnor U19026 (N_19026,N_18767,N_18622);
xnor U19027 (N_19027,N_18446,N_18177);
nor U19028 (N_19028,N_18134,N_18670);
nand U19029 (N_19029,N_18005,N_18919);
xor U19030 (N_19030,N_18627,N_18524);
xnor U19031 (N_19031,N_18347,N_18305);
nand U19032 (N_19032,N_18595,N_18964);
nor U19033 (N_19033,N_18717,N_18781);
or U19034 (N_19034,N_18043,N_18815);
xnor U19035 (N_19035,N_18607,N_18863);
xnor U19036 (N_19036,N_18965,N_18047);
nand U19037 (N_19037,N_18317,N_18832);
nor U19038 (N_19038,N_18388,N_18540);
xor U19039 (N_19039,N_18745,N_18313);
xor U19040 (N_19040,N_18405,N_18861);
nor U19041 (N_19041,N_18940,N_18011);
and U19042 (N_19042,N_18763,N_18895);
nand U19043 (N_19043,N_18805,N_18827);
xnor U19044 (N_19044,N_18661,N_18858);
nand U19045 (N_19045,N_18515,N_18101);
nand U19046 (N_19046,N_18025,N_18421);
or U19047 (N_19047,N_18508,N_18450);
and U19048 (N_19048,N_18578,N_18908);
nor U19049 (N_19049,N_18937,N_18991);
xnor U19050 (N_19050,N_18956,N_18636);
and U19051 (N_19051,N_18231,N_18913);
nor U19052 (N_19052,N_18083,N_18926);
nor U19053 (N_19053,N_18423,N_18377);
nand U19054 (N_19054,N_18434,N_18306);
nor U19055 (N_19055,N_18136,N_18860);
and U19056 (N_19056,N_18768,N_18072);
xnor U19057 (N_19057,N_18776,N_18202);
nand U19058 (N_19058,N_18944,N_18995);
nand U19059 (N_19059,N_18806,N_18062);
and U19060 (N_19060,N_18633,N_18383);
and U19061 (N_19061,N_18785,N_18775);
xnor U19062 (N_19062,N_18734,N_18037);
nand U19063 (N_19063,N_18138,N_18464);
or U19064 (N_19064,N_18625,N_18004);
and U19065 (N_19065,N_18255,N_18330);
nand U19066 (N_19066,N_18962,N_18443);
xor U19067 (N_19067,N_18546,N_18753);
or U19068 (N_19068,N_18250,N_18928);
nor U19069 (N_19069,N_18563,N_18335);
or U19070 (N_19070,N_18295,N_18010);
nor U19071 (N_19071,N_18950,N_18534);
nand U19072 (N_19072,N_18410,N_18536);
or U19073 (N_19073,N_18205,N_18182);
xnor U19074 (N_19074,N_18938,N_18756);
nor U19075 (N_19075,N_18981,N_18204);
nor U19076 (N_19076,N_18656,N_18602);
nor U19077 (N_19077,N_18677,N_18373);
nor U19078 (N_19078,N_18079,N_18638);
or U19079 (N_19079,N_18253,N_18853);
nor U19080 (N_19080,N_18234,N_18259);
nand U19081 (N_19081,N_18752,N_18146);
and U19082 (N_19082,N_18277,N_18478);
xnor U19083 (N_19083,N_18833,N_18996);
nand U19084 (N_19084,N_18128,N_18348);
and U19085 (N_19085,N_18647,N_18145);
or U19086 (N_19086,N_18132,N_18310);
nor U19087 (N_19087,N_18196,N_18361);
nor U19088 (N_19088,N_18346,N_18034);
or U19089 (N_19089,N_18970,N_18787);
nor U19090 (N_19090,N_18172,N_18409);
nor U19091 (N_19091,N_18932,N_18960);
and U19092 (N_19092,N_18572,N_18403);
nor U19093 (N_19093,N_18855,N_18162);
xor U19094 (N_19094,N_18015,N_18151);
xnor U19095 (N_19095,N_18800,N_18213);
xor U19096 (N_19096,N_18654,N_18605);
and U19097 (N_19097,N_18352,N_18706);
or U19098 (N_19098,N_18275,N_18525);
nor U19099 (N_19099,N_18364,N_18958);
xnor U19100 (N_19100,N_18491,N_18046);
nor U19101 (N_19101,N_18618,N_18567);
and U19102 (N_19102,N_18116,N_18603);
xor U19103 (N_19103,N_18163,N_18576);
and U19104 (N_19104,N_18642,N_18056);
nor U19105 (N_19105,N_18099,N_18085);
nand U19106 (N_19106,N_18570,N_18235);
nor U19107 (N_19107,N_18561,N_18127);
nand U19108 (N_19108,N_18093,N_18594);
nand U19109 (N_19109,N_18342,N_18048);
and U19110 (N_19110,N_18529,N_18125);
or U19111 (N_19111,N_18621,N_18510);
or U19112 (N_19112,N_18440,N_18771);
nand U19113 (N_19113,N_18564,N_18917);
nand U19114 (N_19114,N_18140,N_18987);
and U19115 (N_19115,N_18122,N_18176);
nand U19116 (N_19116,N_18119,N_18783);
and U19117 (N_19117,N_18817,N_18747);
nand U19118 (N_19118,N_18862,N_18886);
or U19119 (N_19119,N_18533,N_18465);
and U19120 (N_19120,N_18918,N_18233);
nor U19121 (N_19121,N_18822,N_18497);
or U19122 (N_19122,N_18930,N_18267);
xnor U19123 (N_19123,N_18030,N_18573);
and U19124 (N_19124,N_18194,N_18644);
nor U19125 (N_19125,N_18723,N_18754);
nor U19126 (N_19126,N_18111,N_18531);
nand U19127 (N_19127,N_18216,N_18103);
nand U19128 (N_19128,N_18387,N_18362);
or U19129 (N_19129,N_18582,N_18485);
nor U19130 (N_19130,N_18596,N_18198);
or U19131 (N_19131,N_18121,N_18825);
and U19132 (N_19132,N_18552,N_18057);
and U19133 (N_19133,N_18294,N_18019);
nor U19134 (N_19134,N_18542,N_18566);
nand U19135 (N_19135,N_18087,N_18321);
and U19136 (N_19136,N_18844,N_18489);
or U19137 (N_19137,N_18547,N_18726);
nand U19138 (N_19138,N_18589,N_18027);
nand U19139 (N_19139,N_18732,N_18555);
nand U19140 (N_19140,N_18049,N_18110);
and U19141 (N_19141,N_18158,N_18943);
nor U19142 (N_19142,N_18114,N_18159);
or U19143 (N_19143,N_18139,N_18588);
or U19144 (N_19144,N_18014,N_18413);
xnor U19145 (N_19145,N_18419,N_18657);
or U19146 (N_19146,N_18678,N_18171);
or U19147 (N_19147,N_18495,N_18467);
nand U19148 (N_19148,N_18444,N_18070);
nor U19149 (N_19149,N_18179,N_18984);
and U19150 (N_19150,N_18432,N_18929);
or U19151 (N_19151,N_18215,N_18088);
or U19152 (N_19152,N_18487,N_18469);
nor U19153 (N_19153,N_18986,N_18226);
xnor U19154 (N_19154,N_18008,N_18797);
nor U19155 (N_19155,N_18484,N_18773);
xor U19156 (N_19156,N_18738,N_18838);
or U19157 (N_19157,N_18760,N_18166);
xor U19158 (N_19158,N_18120,N_18278);
nand U19159 (N_19159,N_18795,N_18634);
and U19160 (N_19160,N_18297,N_18448);
or U19161 (N_19161,N_18548,N_18889);
nor U19162 (N_19162,N_18620,N_18708);
or U19163 (N_19163,N_18315,N_18923);
nand U19164 (N_19164,N_18914,N_18282);
nor U19165 (N_19165,N_18189,N_18000);
and U19166 (N_19166,N_18568,N_18668);
xor U19167 (N_19167,N_18195,N_18839);
nor U19168 (N_19168,N_18461,N_18532);
nor U19169 (N_19169,N_18682,N_18556);
nand U19170 (N_19170,N_18915,N_18022);
nor U19171 (N_19171,N_18156,N_18302);
and U19172 (N_19172,N_18199,N_18724);
or U19173 (N_19173,N_18906,N_18583);
xnor U19174 (N_19174,N_18812,N_18701);
xor U19175 (N_19175,N_18982,N_18316);
nor U19176 (N_19176,N_18424,N_18666);
xnor U19177 (N_19177,N_18868,N_18408);
and U19178 (N_19178,N_18418,N_18428);
or U19179 (N_19179,N_18907,N_18396);
and U19180 (N_19180,N_18813,N_18990);
nor U19181 (N_19181,N_18837,N_18933);
nand U19182 (N_19182,N_18126,N_18371);
or U19183 (N_19183,N_18675,N_18615);
nor U19184 (N_19184,N_18791,N_18878);
or U19185 (N_19185,N_18221,N_18051);
or U19186 (N_19186,N_18530,N_18242);
xnor U19187 (N_19187,N_18694,N_18504);
or U19188 (N_19188,N_18341,N_18599);
or U19189 (N_19189,N_18207,N_18269);
and U19190 (N_19190,N_18332,N_18528);
or U19191 (N_19191,N_18150,N_18068);
nand U19192 (N_19192,N_18322,N_18730);
nor U19193 (N_19193,N_18503,N_18522);
xnor U19194 (N_19194,N_18911,N_18271);
xor U19195 (N_19195,N_18327,N_18350);
and U19196 (N_19196,N_18857,N_18512);
nand U19197 (N_19197,N_18592,N_18075);
nand U19198 (N_19198,N_18288,N_18107);
xnor U19199 (N_19199,N_18035,N_18690);
nand U19200 (N_19200,N_18343,N_18673);
or U19201 (N_19201,N_18197,N_18850);
nor U19202 (N_19202,N_18811,N_18641);
xnor U19203 (N_19203,N_18575,N_18792);
nand U19204 (N_19204,N_18663,N_18466);
or U19205 (N_19205,N_18721,N_18819);
nor U19206 (N_19206,N_18091,N_18270);
xor U19207 (N_19207,N_18285,N_18142);
and U19208 (N_19208,N_18842,N_18584);
and U19209 (N_19209,N_18579,N_18585);
nand U19210 (N_19210,N_18076,N_18474);
nand U19211 (N_19211,N_18009,N_18662);
nand U19212 (N_19212,N_18696,N_18251);
or U19213 (N_19213,N_18400,N_18203);
xor U19214 (N_19214,N_18214,N_18574);
and U19215 (N_19215,N_18971,N_18386);
and U19216 (N_19216,N_18698,N_18651);
nor U19217 (N_19217,N_18337,N_18472);
or U19218 (N_19218,N_18784,N_18617);
xnor U19219 (N_19219,N_18246,N_18966);
or U19220 (N_19220,N_18208,N_18947);
or U19221 (N_19221,N_18591,N_18994);
or U19222 (N_19222,N_18002,N_18660);
and U19223 (N_19223,N_18909,N_18081);
nand U19224 (N_19224,N_18632,N_18961);
nand U19225 (N_19225,N_18065,N_18845);
xnor U19226 (N_19226,N_18631,N_18129);
or U19227 (N_19227,N_18431,N_18897);
or U19228 (N_19228,N_18206,N_18693);
xor U19229 (N_19229,N_18260,N_18899);
xnor U19230 (N_19230,N_18643,N_18218);
and U19231 (N_19231,N_18351,N_18358);
nor U19232 (N_19232,N_18628,N_18479);
xor U19233 (N_19233,N_18058,N_18846);
or U19234 (N_19234,N_18509,N_18967);
nor U19235 (N_19235,N_18580,N_18953);
nor U19236 (N_19236,N_18714,N_18980);
nand U19237 (N_19237,N_18016,N_18764);
nor U19238 (N_19238,N_18707,N_18921);
and U19239 (N_19239,N_18757,N_18157);
and U19240 (N_19240,N_18376,N_18963);
nand U19241 (N_19241,N_18679,N_18265);
and U19242 (N_19242,N_18229,N_18108);
nor U19243 (N_19243,N_18407,N_18720);
or U19244 (N_19244,N_18080,N_18818);
xor U19245 (N_19245,N_18289,N_18669);
or U19246 (N_19246,N_18830,N_18069);
or U19247 (N_19247,N_18659,N_18160);
or U19248 (N_19248,N_18033,N_18880);
nand U19249 (N_19249,N_18284,N_18728);
and U19250 (N_19250,N_18606,N_18779);
or U19251 (N_19251,N_18598,N_18587);
or U19252 (N_19252,N_18191,N_18325);
nor U19253 (N_19253,N_18211,N_18712);
or U19254 (N_19254,N_18877,N_18061);
or U19255 (N_19255,N_18280,N_18185);
and U19256 (N_19256,N_18492,N_18823);
or U19257 (N_19257,N_18686,N_18239);
and U19258 (N_19258,N_18268,N_18230);
or U19259 (N_19259,N_18241,N_18169);
nand U19260 (N_19260,N_18648,N_18417);
nand U19261 (N_19261,N_18249,N_18066);
or U19262 (N_19262,N_18137,N_18793);
nand U19263 (N_19263,N_18298,N_18148);
and U19264 (N_19264,N_18406,N_18307);
or U19265 (N_19265,N_18646,N_18702);
xor U19266 (N_19266,N_18073,N_18053);
or U19267 (N_19267,N_18840,N_18097);
or U19268 (N_19268,N_18200,N_18700);
and U19269 (N_19269,N_18856,N_18729);
nand U19270 (N_19270,N_18436,N_18742);
and U19271 (N_19271,N_18799,N_18021);
nand U19272 (N_19272,N_18972,N_18261);
or U19273 (N_19273,N_18074,N_18577);
xnor U19274 (N_19274,N_18296,N_18292);
nor U19275 (N_19275,N_18586,N_18224);
nand U19276 (N_19276,N_18334,N_18885);
and U19277 (N_19277,N_18055,N_18626);
or U19278 (N_19278,N_18257,N_18985);
and U19279 (N_19279,N_18433,N_18319);
nand U19280 (N_19280,N_18256,N_18476);
nor U19281 (N_19281,N_18975,N_18506);
and U19282 (N_19282,N_18244,N_18925);
nand U19283 (N_19283,N_18539,N_18109);
nand U19284 (N_19284,N_18095,N_18124);
and U19285 (N_19285,N_18003,N_18320);
and U19286 (N_19286,N_18652,N_18789);
nand U19287 (N_19287,N_18883,N_18637);
xnor U19288 (N_19288,N_18697,N_18187);
or U19289 (N_19289,N_18834,N_18905);
nand U19290 (N_19290,N_18875,N_18100);
or U19291 (N_19291,N_18471,N_18378);
nand U19292 (N_19292,N_18006,N_18748);
nor U19293 (N_19293,N_18184,N_18248);
xor U19294 (N_19294,N_18425,N_18106);
xnor U19295 (N_19295,N_18688,N_18954);
nand U19296 (N_19296,N_18365,N_18841);
or U19297 (N_19297,N_18640,N_18604);
nand U19298 (N_19298,N_18765,N_18314);
or U19299 (N_19299,N_18152,N_18969);
or U19300 (N_19300,N_18102,N_18777);
nor U19301 (N_19301,N_18992,N_18153);
nand U19302 (N_19302,N_18380,N_18355);
nor U19303 (N_19303,N_18593,N_18366);
nand U19304 (N_19304,N_18397,N_18393);
xor U19305 (N_19305,N_18836,N_18404);
nor U19306 (N_19306,N_18477,N_18681);
or U19307 (N_19307,N_18821,N_18181);
or U19308 (N_19308,N_18064,N_18826);
or U19309 (N_19309,N_18141,N_18609);
nor U19310 (N_19310,N_18349,N_18357);
nand U19311 (N_19311,N_18384,N_18769);
xnor U19312 (N_19312,N_18155,N_18537);
xnor U19313 (N_19313,N_18683,N_18354);
or U19314 (N_19314,N_18903,N_18161);
nand U19315 (N_19315,N_18154,N_18252);
nor U19316 (N_19316,N_18635,N_18067);
nor U19317 (N_19317,N_18382,N_18511);
nand U19318 (N_19318,N_18664,N_18243);
or U19319 (N_19319,N_18237,N_18725);
or U19320 (N_19320,N_18401,N_18900);
nor U19321 (N_19321,N_18927,N_18997);
nand U19322 (N_19322,N_18655,N_18272);
and U19323 (N_19323,N_18311,N_18262);
and U19324 (N_19324,N_18778,N_18608);
or U19325 (N_19325,N_18521,N_18543);
nor U19326 (N_19326,N_18135,N_18326);
xnor U19327 (N_19327,N_18345,N_18475);
or U19328 (N_19328,N_18569,N_18115);
and U19329 (N_19329,N_18807,N_18869);
nor U19330 (N_19330,N_18032,N_18117);
or U19331 (N_19331,N_18758,N_18737);
and U19332 (N_19332,N_18864,N_18870);
nor U19333 (N_19333,N_18974,N_18026);
and U19334 (N_19334,N_18422,N_18174);
xor U19335 (N_19335,N_18118,N_18227);
nor U19336 (N_19336,N_18993,N_18581);
and U19337 (N_19337,N_18353,N_18887);
or U19338 (N_19338,N_18619,N_18462);
xnor U19339 (N_19339,N_18225,N_18374);
nand U19340 (N_19340,N_18505,N_18977);
nand U19341 (N_19341,N_18323,N_18193);
nor U19342 (N_19342,N_18945,N_18920);
and U19343 (N_19343,N_18412,N_18415);
xnor U19344 (N_19344,N_18959,N_18293);
nor U19345 (N_19345,N_18715,N_18916);
and U19346 (N_19346,N_18254,N_18849);
or U19347 (N_19347,N_18931,N_18266);
nor U19348 (N_19348,N_18544,N_18013);
xor U19349 (N_19349,N_18437,N_18976);
and U19350 (N_19350,N_18759,N_18517);
nand U19351 (N_19351,N_18133,N_18803);
xor U19352 (N_19352,N_18442,N_18687);
nand U19353 (N_19353,N_18790,N_18391);
and U19354 (N_19354,N_18222,N_18553);
nand U19355 (N_19355,N_18866,N_18499);
or U19356 (N_19356,N_18814,N_18264);
xnor U19357 (N_19357,N_18052,N_18653);
xor U19358 (N_19358,N_18468,N_18894);
nor U19359 (N_19359,N_18077,N_18175);
xor U19360 (N_19360,N_18094,N_18600);
or U19361 (N_19361,N_18247,N_18143);
xnor U19362 (N_19362,N_18957,N_18209);
and U19363 (N_19363,N_18500,N_18924);
nor U19364 (N_19364,N_18516,N_18676);
nor U19365 (N_19365,N_18601,N_18761);
xnor U19366 (N_19366,N_18876,N_18939);
or U19367 (N_19367,N_18245,N_18274);
nor U19368 (N_19368,N_18501,N_18782);
nor U19369 (N_19369,N_18874,N_18824);
and U19370 (N_19370,N_18744,N_18999);
and U19371 (N_19371,N_18611,N_18390);
nor U19372 (N_19372,N_18898,N_18884);
nand U19373 (N_19373,N_18685,N_18623);
xor U19374 (N_19374,N_18859,N_18144);
xor U19375 (N_19375,N_18852,N_18796);
nand U19376 (N_19376,N_18190,N_18183);
and U19377 (N_19377,N_18340,N_18178);
nor U19378 (N_19378,N_18040,N_18089);
xnor U19379 (N_19379,N_18801,N_18851);
and U19380 (N_19380,N_18041,N_18236);
nor U19381 (N_19381,N_18273,N_18854);
and U19382 (N_19382,N_18983,N_18452);
and U19383 (N_19383,N_18459,N_18755);
or U19384 (N_19384,N_18470,N_18494);
nand U19385 (N_19385,N_18458,N_18809);
nand U19386 (N_19386,N_18695,N_18689);
and U19387 (N_19387,N_18650,N_18810);
nand U19388 (N_19388,N_18188,N_18012);
nand U19389 (N_19389,N_18735,N_18054);
xnor U19390 (N_19390,N_18219,N_18078);
or U19391 (N_19391,N_18303,N_18170);
and U19392 (N_19392,N_18228,N_18445);
nor U19393 (N_19393,N_18902,N_18722);
or U19394 (N_19394,N_18463,N_18086);
nand U19395 (N_19395,N_18258,N_18367);
nor U19396 (N_19396,N_18028,N_18718);
nand U19397 (N_19397,N_18952,N_18571);
xor U19398 (N_19398,N_18473,N_18816);
nand U19399 (N_19399,N_18711,N_18427);
or U19400 (N_19400,N_18780,N_18082);
nor U19401 (N_19401,N_18829,N_18092);
nor U19402 (N_19402,N_18879,N_18039);
nand U19403 (N_19403,N_18667,N_18704);
nand U19404 (N_19404,N_18526,N_18217);
nor U19405 (N_19405,N_18451,N_18703);
nand U19406 (N_19406,N_18324,N_18551);
xnor U19407 (N_19407,N_18562,N_18535);
or U19408 (N_19408,N_18416,N_18979);
and U19409 (N_19409,N_18336,N_18483);
and U19410 (N_19410,N_18286,N_18518);
xor U19411 (N_19411,N_18105,N_18389);
xnor U19412 (N_19412,N_18750,N_18029);
xor U19413 (N_19413,N_18867,N_18071);
nand U19414 (N_19414,N_18036,N_18290);
xor U19415 (N_19415,N_18762,N_18498);
and U19416 (N_19416,N_18523,N_18480);
and U19417 (N_19417,N_18287,N_18359);
or U19418 (N_19418,N_18882,N_18808);
and U19419 (N_19419,N_18951,N_18130);
and U19420 (N_19420,N_18719,N_18490);
nand U19421 (N_19421,N_18090,N_18507);
nand U19422 (N_19422,N_18514,N_18098);
and U19423 (N_19423,N_18743,N_18038);
nor U19424 (N_19424,N_18460,N_18912);
or U19425 (N_19425,N_18624,N_18186);
xor U19426 (N_19426,N_18904,N_18220);
nand U19427 (N_19427,N_18240,N_18835);
xnor U19428 (N_19428,N_18385,N_18429);
or U19429 (N_19429,N_18936,N_18671);
or U19430 (N_19430,N_18164,N_18447);
nand U19431 (N_19431,N_18740,N_18665);
nand U19432 (N_19432,N_18430,N_18847);
or U19433 (N_19433,N_18888,N_18398);
xnor U19434 (N_19434,N_18173,N_18104);
nor U19435 (N_19435,N_18770,N_18672);
xor U19436 (N_19436,N_18713,N_18059);
or U19437 (N_19437,N_18998,N_18788);
nor U19438 (N_19438,N_18658,N_18333);
nor U19439 (N_19439,N_18379,N_18941);
xnor U19440 (N_19440,N_18699,N_18680);
xor U19441 (N_19441,N_18973,N_18749);
xor U19442 (N_19442,N_18772,N_18614);
xor U19443 (N_19443,N_18238,N_18165);
and U19444 (N_19444,N_18192,N_18339);
and U19445 (N_19445,N_18084,N_18527);
nand U19446 (N_19446,N_18786,N_18843);
xor U19447 (N_19447,N_18630,N_18881);
nor U19448 (N_19448,N_18493,N_18147);
nor U19449 (N_19449,N_18549,N_18329);
xor U19450 (N_19450,N_18731,N_18934);
nand U19451 (N_19451,N_18439,N_18044);
nand U19452 (N_19452,N_18318,N_18441);
nand U19453 (N_19453,N_18559,N_18210);
and U19454 (N_19454,N_18481,N_18482);
or U19455 (N_19455,N_18645,N_18922);
xor U19456 (N_19456,N_18560,N_18502);
or U19457 (N_19457,N_18123,N_18893);
or U19458 (N_19458,N_18063,N_18201);
nand U19459 (N_19459,N_18612,N_18017);
nand U19460 (N_19460,N_18774,N_18453);
and U19461 (N_19461,N_18610,N_18968);
or U19462 (N_19462,N_18649,N_18276);
xor U19463 (N_19463,N_18375,N_18212);
or U19464 (N_19464,N_18989,N_18001);
nor U19465 (N_19465,N_18873,N_18031);
nor U19466 (N_19466,N_18828,N_18223);
and U19467 (N_19467,N_18331,N_18394);
nor U19468 (N_19468,N_18613,N_18486);
nand U19469 (N_19469,N_18449,N_18739);
and U19470 (N_19470,N_18709,N_18871);
nand U19471 (N_19471,N_18565,N_18414);
or U19472 (N_19472,N_18978,N_18096);
and U19473 (N_19473,N_18541,N_18955);
nor U19474 (N_19474,N_18691,N_18896);
xnor U19475 (N_19475,N_18232,N_18804);
xor U19476 (N_19476,N_18891,N_18304);
and U19477 (N_19477,N_18338,N_18727);
xnor U19478 (N_19478,N_18705,N_18023);
nor U19479 (N_19479,N_18308,N_18392);
nand U19480 (N_19480,N_18300,N_18399);
nand U19481 (N_19481,N_18281,N_18360);
or U19482 (N_19482,N_18942,N_18766);
and U19483 (N_19483,N_18848,N_18746);
nand U19484 (N_19484,N_18557,N_18381);
xnor U19485 (N_19485,N_18411,N_18263);
xor U19486 (N_19486,N_18558,N_18356);
and U19487 (N_19487,N_18910,N_18692);
nand U19488 (N_19488,N_18279,N_18946);
and U19489 (N_19489,N_18751,N_18741);
or U19490 (N_19490,N_18949,N_18865);
nor U19491 (N_19491,N_18180,N_18935);
and U19492 (N_19492,N_18369,N_18438);
or U19493 (N_19493,N_18060,N_18520);
and U19494 (N_19494,N_18736,N_18639);
or U19495 (N_19495,N_18426,N_18112);
or U19496 (N_19496,N_18488,N_18042);
xor U19497 (N_19497,N_18901,N_18820);
nor U19498 (N_19498,N_18454,N_18344);
xnor U19499 (N_19499,N_18616,N_18299);
or U19500 (N_19500,N_18632,N_18330);
or U19501 (N_19501,N_18263,N_18573);
or U19502 (N_19502,N_18019,N_18331);
xnor U19503 (N_19503,N_18773,N_18956);
and U19504 (N_19504,N_18348,N_18787);
nand U19505 (N_19505,N_18220,N_18673);
and U19506 (N_19506,N_18279,N_18619);
nand U19507 (N_19507,N_18429,N_18236);
and U19508 (N_19508,N_18758,N_18952);
nor U19509 (N_19509,N_18516,N_18809);
xnor U19510 (N_19510,N_18005,N_18383);
and U19511 (N_19511,N_18484,N_18600);
xor U19512 (N_19512,N_18934,N_18580);
or U19513 (N_19513,N_18525,N_18695);
xnor U19514 (N_19514,N_18526,N_18139);
xor U19515 (N_19515,N_18723,N_18706);
and U19516 (N_19516,N_18705,N_18272);
nand U19517 (N_19517,N_18594,N_18401);
nor U19518 (N_19518,N_18949,N_18080);
xnor U19519 (N_19519,N_18922,N_18346);
nand U19520 (N_19520,N_18919,N_18831);
and U19521 (N_19521,N_18220,N_18252);
or U19522 (N_19522,N_18322,N_18547);
nand U19523 (N_19523,N_18551,N_18612);
xor U19524 (N_19524,N_18718,N_18277);
and U19525 (N_19525,N_18402,N_18471);
or U19526 (N_19526,N_18444,N_18255);
or U19527 (N_19527,N_18254,N_18762);
xnor U19528 (N_19528,N_18751,N_18112);
or U19529 (N_19529,N_18380,N_18267);
nor U19530 (N_19530,N_18357,N_18735);
and U19531 (N_19531,N_18702,N_18188);
nor U19532 (N_19532,N_18418,N_18201);
or U19533 (N_19533,N_18159,N_18378);
or U19534 (N_19534,N_18443,N_18832);
nand U19535 (N_19535,N_18022,N_18671);
xor U19536 (N_19536,N_18907,N_18100);
or U19537 (N_19537,N_18395,N_18868);
nand U19538 (N_19538,N_18268,N_18255);
nand U19539 (N_19539,N_18848,N_18745);
nor U19540 (N_19540,N_18286,N_18687);
or U19541 (N_19541,N_18568,N_18575);
xor U19542 (N_19542,N_18167,N_18589);
and U19543 (N_19543,N_18841,N_18271);
or U19544 (N_19544,N_18014,N_18706);
xor U19545 (N_19545,N_18497,N_18306);
xor U19546 (N_19546,N_18210,N_18799);
nand U19547 (N_19547,N_18585,N_18157);
and U19548 (N_19548,N_18254,N_18396);
nand U19549 (N_19549,N_18324,N_18244);
xnor U19550 (N_19550,N_18901,N_18246);
or U19551 (N_19551,N_18249,N_18145);
and U19552 (N_19552,N_18549,N_18928);
nor U19553 (N_19553,N_18060,N_18077);
and U19554 (N_19554,N_18870,N_18621);
or U19555 (N_19555,N_18441,N_18756);
nor U19556 (N_19556,N_18787,N_18400);
nand U19557 (N_19557,N_18324,N_18163);
xnor U19558 (N_19558,N_18636,N_18678);
and U19559 (N_19559,N_18291,N_18442);
xnor U19560 (N_19560,N_18432,N_18662);
xnor U19561 (N_19561,N_18993,N_18927);
and U19562 (N_19562,N_18272,N_18005);
nor U19563 (N_19563,N_18857,N_18547);
xnor U19564 (N_19564,N_18437,N_18939);
and U19565 (N_19565,N_18238,N_18530);
nor U19566 (N_19566,N_18223,N_18603);
nor U19567 (N_19567,N_18844,N_18554);
and U19568 (N_19568,N_18067,N_18867);
nor U19569 (N_19569,N_18929,N_18280);
and U19570 (N_19570,N_18996,N_18924);
and U19571 (N_19571,N_18560,N_18682);
or U19572 (N_19572,N_18788,N_18414);
or U19573 (N_19573,N_18376,N_18697);
nand U19574 (N_19574,N_18051,N_18066);
xnor U19575 (N_19575,N_18112,N_18261);
nand U19576 (N_19576,N_18619,N_18159);
or U19577 (N_19577,N_18649,N_18949);
or U19578 (N_19578,N_18788,N_18140);
and U19579 (N_19579,N_18222,N_18725);
and U19580 (N_19580,N_18824,N_18676);
xor U19581 (N_19581,N_18438,N_18107);
or U19582 (N_19582,N_18919,N_18868);
and U19583 (N_19583,N_18969,N_18685);
nand U19584 (N_19584,N_18507,N_18086);
nor U19585 (N_19585,N_18701,N_18488);
nor U19586 (N_19586,N_18492,N_18685);
or U19587 (N_19587,N_18192,N_18545);
or U19588 (N_19588,N_18286,N_18447);
and U19589 (N_19589,N_18523,N_18910);
xor U19590 (N_19590,N_18642,N_18916);
or U19591 (N_19591,N_18669,N_18804);
and U19592 (N_19592,N_18709,N_18214);
nand U19593 (N_19593,N_18523,N_18665);
nor U19594 (N_19594,N_18233,N_18718);
and U19595 (N_19595,N_18398,N_18149);
xnor U19596 (N_19596,N_18602,N_18122);
or U19597 (N_19597,N_18069,N_18437);
and U19598 (N_19598,N_18611,N_18986);
xnor U19599 (N_19599,N_18391,N_18263);
nand U19600 (N_19600,N_18574,N_18629);
xnor U19601 (N_19601,N_18479,N_18494);
nor U19602 (N_19602,N_18650,N_18306);
nand U19603 (N_19603,N_18469,N_18733);
xnor U19604 (N_19604,N_18387,N_18315);
or U19605 (N_19605,N_18413,N_18785);
nand U19606 (N_19606,N_18538,N_18655);
nor U19607 (N_19607,N_18998,N_18847);
xnor U19608 (N_19608,N_18534,N_18122);
and U19609 (N_19609,N_18125,N_18978);
nor U19610 (N_19610,N_18772,N_18638);
and U19611 (N_19611,N_18429,N_18203);
nor U19612 (N_19612,N_18142,N_18565);
nand U19613 (N_19613,N_18409,N_18569);
nand U19614 (N_19614,N_18476,N_18120);
and U19615 (N_19615,N_18148,N_18638);
xor U19616 (N_19616,N_18572,N_18675);
xor U19617 (N_19617,N_18671,N_18622);
and U19618 (N_19618,N_18345,N_18418);
or U19619 (N_19619,N_18140,N_18238);
xnor U19620 (N_19620,N_18231,N_18899);
or U19621 (N_19621,N_18300,N_18764);
nor U19622 (N_19622,N_18933,N_18203);
and U19623 (N_19623,N_18798,N_18669);
or U19624 (N_19624,N_18477,N_18002);
nor U19625 (N_19625,N_18171,N_18905);
xnor U19626 (N_19626,N_18529,N_18922);
nor U19627 (N_19627,N_18244,N_18868);
nand U19628 (N_19628,N_18204,N_18177);
and U19629 (N_19629,N_18000,N_18202);
xor U19630 (N_19630,N_18112,N_18021);
or U19631 (N_19631,N_18446,N_18304);
or U19632 (N_19632,N_18836,N_18069);
and U19633 (N_19633,N_18066,N_18417);
and U19634 (N_19634,N_18612,N_18651);
nor U19635 (N_19635,N_18159,N_18919);
and U19636 (N_19636,N_18865,N_18265);
and U19637 (N_19637,N_18655,N_18290);
or U19638 (N_19638,N_18075,N_18635);
or U19639 (N_19639,N_18899,N_18672);
nor U19640 (N_19640,N_18070,N_18156);
nor U19641 (N_19641,N_18959,N_18456);
xnor U19642 (N_19642,N_18650,N_18967);
nand U19643 (N_19643,N_18101,N_18825);
xnor U19644 (N_19644,N_18055,N_18953);
nand U19645 (N_19645,N_18142,N_18298);
nand U19646 (N_19646,N_18171,N_18389);
nand U19647 (N_19647,N_18150,N_18136);
nand U19648 (N_19648,N_18886,N_18993);
nand U19649 (N_19649,N_18780,N_18939);
nor U19650 (N_19650,N_18499,N_18894);
and U19651 (N_19651,N_18280,N_18839);
or U19652 (N_19652,N_18821,N_18088);
xnor U19653 (N_19653,N_18070,N_18910);
nand U19654 (N_19654,N_18762,N_18830);
and U19655 (N_19655,N_18008,N_18489);
and U19656 (N_19656,N_18150,N_18229);
nor U19657 (N_19657,N_18446,N_18323);
xor U19658 (N_19658,N_18422,N_18503);
or U19659 (N_19659,N_18340,N_18626);
nor U19660 (N_19660,N_18494,N_18905);
xnor U19661 (N_19661,N_18692,N_18144);
xnor U19662 (N_19662,N_18485,N_18111);
nand U19663 (N_19663,N_18988,N_18258);
and U19664 (N_19664,N_18052,N_18854);
xnor U19665 (N_19665,N_18792,N_18496);
nor U19666 (N_19666,N_18896,N_18931);
xnor U19667 (N_19667,N_18170,N_18017);
nor U19668 (N_19668,N_18860,N_18851);
and U19669 (N_19669,N_18805,N_18962);
nor U19670 (N_19670,N_18471,N_18197);
or U19671 (N_19671,N_18509,N_18059);
nor U19672 (N_19672,N_18840,N_18976);
nand U19673 (N_19673,N_18557,N_18875);
xor U19674 (N_19674,N_18714,N_18685);
or U19675 (N_19675,N_18829,N_18996);
nand U19676 (N_19676,N_18397,N_18191);
or U19677 (N_19677,N_18395,N_18397);
or U19678 (N_19678,N_18435,N_18363);
or U19679 (N_19679,N_18488,N_18706);
xor U19680 (N_19680,N_18546,N_18704);
xor U19681 (N_19681,N_18712,N_18398);
and U19682 (N_19682,N_18636,N_18028);
and U19683 (N_19683,N_18047,N_18170);
xor U19684 (N_19684,N_18480,N_18931);
nor U19685 (N_19685,N_18235,N_18764);
xor U19686 (N_19686,N_18298,N_18093);
nand U19687 (N_19687,N_18957,N_18631);
nor U19688 (N_19688,N_18494,N_18391);
or U19689 (N_19689,N_18904,N_18375);
nor U19690 (N_19690,N_18526,N_18726);
and U19691 (N_19691,N_18094,N_18339);
xor U19692 (N_19692,N_18097,N_18609);
and U19693 (N_19693,N_18421,N_18852);
xor U19694 (N_19694,N_18219,N_18692);
nor U19695 (N_19695,N_18649,N_18064);
nor U19696 (N_19696,N_18622,N_18984);
nor U19697 (N_19697,N_18209,N_18886);
and U19698 (N_19698,N_18270,N_18046);
nand U19699 (N_19699,N_18709,N_18485);
and U19700 (N_19700,N_18221,N_18075);
and U19701 (N_19701,N_18494,N_18401);
xor U19702 (N_19702,N_18304,N_18315);
xnor U19703 (N_19703,N_18548,N_18910);
xor U19704 (N_19704,N_18113,N_18829);
xnor U19705 (N_19705,N_18976,N_18455);
nor U19706 (N_19706,N_18571,N_18194);
nand U19707 (N_19707,N_18531,N_18808);
and U19708 (N_19708,N_18879,N_18910);
xor U19709 (N_19709,N_18243,N_18261);
xor U19710 (N_19710,N_18614,N_18211);
and U19711 (N_19711,N_18723,N_18214);
or U19712 (N_19712,N_18281,N_18524);
xor U19713 (N_19713,N_18726,N_18946);
and U19714 (N_19714,N_18425,N_18663);
nor U19715 (N_19715,N_18013,N_18236);
nand U19716 (N_19716,N_18541,N_18684);
nand U19717 (N_19717,N_18186,N_18482);
xnor U19718 (N_19718,N_18094,N_18643);
nand U19719 (N_19719,N_18195,N_18406);
nand U19720 (N_19720,N_18669,N_18796);
and U19721 (N_19721,N_18987,N_18519);
xnor U19722 (N_19722,N_18333,N_18575);
nand U19723 (N_19723,N_18628,N_18313);
nand U19724 (N_19724,N_18619,N_18120);
or U19725 (N_19725,N_18391,N_18797);
and U19726 (N_19726,N_18266,N_18966);
and U19727 (N_19727,N_18017,N_18258);
or U19728 (N_19728,N_18256,N_18105);
and U19729 (N_19729,N_18966,N_18646);
and U19730 (N_19730,N_18566,N_18087);
and U19731 (N_19731,N_18932,N_18319);
xor U19732 (N_19732,N_18279,N_18836);
nor U19733 (N_19733,N_18565,N_18563);
xor U19734 (N_19734,N_18690,N_18968);
nand U19735 (N_19735,N_18329,N_18078);
or U19736 (N_19736,N_18111,N_18224);
nand U19737 (N_19737,N_18612,N_18902);
or U19738 (N_19738,N_18944,N_18828);
nand U19739 (N_19739,N_18772,N_18767);
or U19740 (N_19740,N_18826,N_18459);
or U19741 (N_19741,N_18225,N_18759);
nor U19742 (N_19742,N_18855,N_18781);
nor U19743 (N_19743,N_18399,N_18409);
nand U19744 (N_19744,N_18155,N_18154);
nand U19745 (N_19745,N_18766,N_18536);
xor U19746 (N_19746,N_18313,N_18327);
nand U19747 (N_19747,N_18999,N_18264);
nor U19748 (N_19748,N_18752,N_18268);
or U19749 (N_19749,N_18533,N_18873);
nand U19750 (N_19750,N_18574,N_18450);
or U19751 (N_19751,N_18067,N_18697);
xnor U19752 (N_19752,N_18689,N_18083);
or U19753 (N_19753,N_18224,N_18157);
and U19754 (N_19754,N_18122,N_18166);
xor U19755 (N_19755,N_18138,N_18995);
xor U19756 (N_19756,N_18805,N_18612);
or U19757 (N_19757,N_18945,N_18055);
nor U19758 (N_19758,N_18092,N_18100);
or U19759 (N_19759,N_18675,N_18476);
and U19760 (N_19760,N_18645,N_18234);
nand U19761 (N_19761,N_18923,N_18598);
nor U19762 (N_19762,N_18307,N_18305);
nand U19763 (N_19763,N_18914,N_18009);
and U19764 (N_19764,N_18519,N_18165);
nor U19765 (N_19765,N_18412,N_18483);
or U19766 (N_19766,N_18859,N_18140);
or U19767 (N_19767,N_18505,N_18213);
nor U19768 (N_19768,N_18941,N_18914);
xor U19769 (N_19769,N_18548,N_18171);
xor U19770 (N_19770,N_18826,N_18668);
nor U19771 (N_19771,N_18169,N_18257);
xor U19772 (N_19772,N_18530,N_18463);
or U19773 (N_19773,N_18509,N_18274);
nor U19774 (N_19774,N_18979,N_18167);
nand U19775 (N_19775,N_18674,N_18194);
nand U19776 (N_19776,N_18172,N_18846);
nor U19777 (N_19777,N_18477,N_18439);
nand U19778 (N_19778,N_18296,N_18824);
and U19779 (N_19779,N_18408,N_18483);
or U19780 (N_19780,N_18743,N_18622);
or U19781 (N_19781,N_18811,N_18187);
and U19782 (N_19782,N_18095,N_18376);
nand U19783 (N_19783,N_18818,N_18575);
or U19784 (N_19784,N_18015,N_18963);
nand U19785 (N_19785,N_18447,N_18515);
or U19786 (N_19786,N_18573,N_18555);
nand U19787 (N_19787,N_18649,N_18641);
nand U19788 (N_19788,N_18576,N_18259);
xnor U19789 (N_19789,N_18572,N_18699);
or U19790 (N_19790,N_18162,N_18421);
nor U19791 (N_19791,N_18381,N_18465);
nor U19792 (N_19792,N_18210,N_18809);
and U19793 (N_19793,N_18604,N_18554);
nand U19794 (N_19794,N_18998,N_18826);
nand U19795 (N_19795,N_18499,N_18153);
or U19796 (N_19796,N_18497,N_18434);
xnor U19797 (N_19797,N_18427,N_18584);
and U19798 (N_19798,N_18080,N_18936);
xnor U19799 (N_19799,N_18115,N_18523);
nand U19800 (N_19800,N_18956,N_18157);
and U19801 (N_19801,N_18882,N_18212);
or U19802 (N_19802,N_18367,N_18006);
nor U19803 (N_19803,N_18955,N_18905);
and U19804 (N_19804,N_18226,N_18479);
or U19805 (N_19805,N_18324,N_18296);
xnor U19806 (N_19806,N_18969,N_18437);
nand U19807 (N_19807,N_18027,N_18379);
or U19808 (N_19808,N_18216,N_18000);
xnor U19809 (N_19809,N_18301,N_18870);
or U19810 (N_19810,N_18993,N_18789);
xor U19811 (N_19811,N_18524,N_18143);
xor U19812 (N_19812,N_18868,N_18366);
and U19813 (N_19813,N_18129,N_18109);
and U19814 (N_19814,N_18902,N_18431);
xnor U19815 (N_19815,N_18017,N_18617);
and U19816 (N_19816,N_18499,N_18668);
nor U19817 (N_19817,N_18752,N_18407);
or U19818 (N_19818,N_18759,N_18346);
nor U19819 (N_19819,N_18288,N_18825);
nor U19820 (N_19820,N_18216,N_18799);
nand U19821 (N_19821,N_18106,N_18188);
nand U19822 (N_19822,N_18152,N_18621);
nor U19823 (N_19823,N_18119,N_18513);
or U19824 (N_19824,N_18811,N_18079);
xor U19825 (N_19825,N_18776,N_18387);
xor U19826 (N_19826,N_18559,N_18724);
nand U19827 (N_19827,N_18504,N_18625);
xor U19828 (N_19828,N_18284,N_18975);
nor U19829 (N_19829,N_18614,N_18314);
nand U19830 (N_19830,N_18944,N_18256);
xnor U19831 (N_19831,N_18865,N_18199);
nor U19832 (N_19832,N_18877,N_18139);
and U19833 (N_19833,N_18345,N_18218);
and U19834 (N_19834,N_18446,N_18569);
xor U19835 (N_19835,N_18336,N_18743);
and U19836 (N_19836,N_18479,N_18758);
nand U19837 (N_19837,N_18840,N_18121);
xnor U19838 (N_19838,N_18786,N_18998);
and U19839 (N_19839,N_18993,N_18958);
xnor U19840 (N_19840,N_18132,N_18693);
and U19841 (N_19841,N_18158,N_18216);
nor U19842 (N_19842,N_18289,N_18071);
nor U19843 (N_19843,N_18148,N_18716);
nor U19844 (N_19844,N_18147,N_18817);
xor U19845 (N_19845,N_18662,N_18664);
nor U19846 (N_19846,N_18368,N_18222);
or U19847 (N_19847,N_18494,N_18879);
xor U19848 (N_19848,N_18241,N_18735);
or U19849 (N_19849,N_18614,N_18490);
and U19850 (N_19850,N_18781,N_18883);
xor U19851 (N_19851,N_18938,N_18490);
xnor U19852 (N_19852,N_18118,N_18919);
or U19853 (N_19853,N_18384,N_18876);
nor U19854 (N_19854,N_18015,N_18179);
and U19855 (N_19855,N_18372,N_18259);
nor U19856 (N_19856,N_18313,N_18037);
nand U19857 (N_19857,N_18293,N_18704);
xor U19858 (N_19858,N_18110,N_18810);
nand U19859 (N_19859,N_18726,N_18484);
nand U19860 (N_19860,N_18117,N_18075);
and U19861 (N_19861,N_18368,N_18770);
or U19862 (N_19862,N_18570,N_18192);
or U19863 (N_19863,N_18109,N_18546);
or U19864 (N_19864,N_18719,N_18849);
nand U19865 (N_19865,N_18981,N_18215);
xor U19866 (N_19866,N_18897,N_18702);
or U19867 (N_19867,N_18952,N_18948);
and U19868 (N_19868,N_18707,N_18684);
and U19869 (N_19869,N_18606,N_18594);
xnor U19870 (N_19870,N_18676,N_18249);
nor U19871 (N_19871,N_18380,N_18394);
xnor U19872 (N_19872,N_18189,N_18900);
and U19873 (N_19873,N_18749,N_18459);
nand U19874 (N_19874,N_18296,N_18237);
and U19875 (N_19875,N_18614,N_18083);
nor U19876 (N_19876,N_18901,N_18831);
xor U19877 (N_19877,N_18144,N_18568);
or U19878 (N_19878,N_18274,N_18978);
and U19879 (N_19879,N_18289,N_18728);
or U19880 (N_19880,N_18927,N_18211);
nor U19881 (N_19881,N_18259,N_18450);
and U19882 (N_19882,N_18567,N_18655);
or U19883 (N_19883,N_18899,N_18631);
xor U19884 (N_19884,N_18739,N_18754);
or U19885 (N_19885,N_18600,N_18217);
nor U19886 (N_19886,N_18854,N_18919);
nand U19887 (N_19887,N_18881,N_18986);
nor U19888 (N_19888,N_18954,N_18222);
or U19889 (N_19889,N_18870,N_18622);
and U19890 (N_19890,N_18915,N_18945);
or U19891 (N_19891,N_18298,N_18761);
and U19892 (N_19892,N_18747,N_18553);
or U19893 (N_19893,N_18720,N_18132);
nand U19894 (N_19894,N_18101,N_18901);
xor U19895 (N_19895,N_18569,N_18918);
and U19896 (N_19896,N_18494,N_18282);
and U19897 (N_19897,N_18776,N_18888);
nor U19898 (N_19898,N_18973,N_18245);
nand U19899 (N_19899,N_18810,N_18624);
or U19900 (N_19900,N_18009,N_18708);
nand U19901 (N_19901,N_18992,N_18717);
nand U19902 (N_19902,N_18734,N_18466);
or U19903 (N_19903,N_18972,N_18385);
or U19904 (N_19904,N_18402,N_18312);
nor U19905 (N_19905,N_18336,N_18278);
nor U19906 (N_19906,N_18592,N_18421);
nor U19907 (N_19907,N_18527,N_18012);
or U19908 (N_19908,N_18157,N_18191);
nor U19909 (N_19909,N_18217,N_18132);
or U19910 (N_19910,N_18218,N_18704);
nor U19911 (N_19911,N_18519,N_18099);
nand U19912 (N_19912,N_18551,N_18344);
xor U19913 (N_19913,N_18163,N_18540);
and U19914 (N_19914,N_18176,N_18732);
nor U19915 (N_19915,N_18598,N_18770);
xor U19916 (N_19916,N_18026,N_18828);
nand U19917 (N_19917,N_18709,N_18212);
nor U19918 (N_19918,N_18699,N_18245);
or U19919 (N_19919,N_18410,N_18880);
nor U19920 (N_19920,N_18336,N_18332);
xor U19921 (N_19921,N_18361,N_18671);
or U19922 (N_19922,N_18432,N_18033);
or U19923 (N_19923,N_18942,N_18949);
xnor U19924 (N_19924,N_18647,N_18238);
or U19925 (N_19925,N_18204,N_18150);
nand U19926 (N_19926,N_18396,N_18457);
or U19927 (N_19927,N_18539,N_18127);
nand U19928 (N_19928,N_18826,N_18655);
xnor U19929 (N_19929,N_18541,N_18474);
nand U19930 (N_19930,N_18592,N_18363);
xnor U19931 (N_19931,N_18259,N_18226);
and U19932 (N_19932,N_18245,N_18713);
xor U19933 (N_19933,N_18323,N_18654);
and U19934 (N_19934,N_18067,N_18784);
or U19935 (N_19935,N_18015,N_18667);
or U19936 (N_19936,N_18466,N_18748);
xnor U19937 (N_19937,N_18579,N_18594);
nor U19938 (N_19938,N_18605,N_18634);
or U19939 (N_19939,N_18312,N_18557);
and U19940 (N_19940,N_18661,N_18428);
nor U19941 (N_19941,N_18489,N_18224);
and U19942 (N_19942,N_18126,N_18394);
and U19943 (N_19943,N_18988,N_18197);
and U19944 (N_19944,N_18511,N_18281);
nand U19945 (N_19945,N_18268,N_18331);
and U19946 (N_19946,N_18095,N_18659);
and U19947 (N_19947,N_18611,N_18883);
or U19948 (N_19948,N_18123,N_18479);
and U19949 (N_19949,N_18393,N_18572);
xor U19950 (N_19950,N_18865,N_18197);
xor U19951 (N_19951,N_18469,N_18738);
nor U19952 (N_19952,N_18911,N_18138);
xnor U19953 (N_19953,N_18812,N_18759);
nand U19954 (N_19954,N_18651,N_18761);
or U19955 (N_19955,N_18491,N_18672);
and U19956 (N_19956,N_18650,N_18968);
nand U19957 (N_19957,N_18962,N_18170);
and U19958 (N_19958,N_18374,N_18665);
xor U19959 (N_19959,N_18873,N_18760);
nor U19960 (N_19960,N_18207,N_18510);
or U19961 (N_19961,N_18642,N_18265);
xnor U19962 (N_19962,N_18351,N_18685);
and U19963 (N_19963,N_18743,N_18809);
and U19964 (N_19964,N_18993,N_18282);
nor U19965 (N_19965,N_18925,N_18515);
or U19966 (N_19966,N_18343,N_18988);
nand U19967 (N_19967,N_18661,N_18276);
or U19968 (N_19968,N_18755,N_18806);
nand U19969 (N_19969,N_18834,N_18605);
and U19970 (N_19970,N_18194,N_18788);
and U19971 (N_19971,N_18601,N_18347);
and U19972 (N_19972,N_18815,N_18831);
xor U19973 (N_19973,N_18420,N_18606);
and U19974 (N_19974,N_18570,N_18150);
and U19975 (N_19975,N_18060,N_18818);
nand U19976 (N_19976,N_18384,N_18271);
and U19977 (N_19977,N_18428,N_18861);
nand U19978 (N_19978,N_18514,N_18729);
xor U19979 (N_19979,N_18698,N_18764);
or U19980 (N_19980,N_18361,N_18084);
and U19981 (N_19981,N_18018,N_18407);
and U19982 (N_19982,N_18740,N_18116);
nand U19983 (N_19983,N_18796,N_18625);
or U19984 (N_19984,N_18359,N_18091);
xnor U19985 (N_19985,N_18995,N_18561);
nor U19986 (N_19986,N_18765,N_18972);
or U19987 (N_19987,N_18179,N_18945);
nor U19988 (N_19988,N_18285,N_18216);
and U19989 (N_19989,N_18616,N_18314);
nand U19990 (N_19990,N_18087,N_18358);
xor U19991 (N_19991,N_18750,N_18636);
nor U19992 (N_19992,N_18278,N_18558);
or U19993 (N_19993,N_18776,N_18014);
and U19994 (N_19994,N_18744,N_18769);
or U19995 (N_19995,N_18611,N_18460);
or U19996 (N_19996,N_18595,N_18312);
nor U19997 (N_19997,N_18958,N_18833);
or U19998 (N_19998,N_18208,N_18929);
xor U19999 (N_19999,N_18131,N_18563);
nand UO_0 (O_0,N_19756,N_19686);
or UO_1 (O_1,N_19357,N_19378);
or UO_2 (O_2,N_19234,N_19184);
nor UO_3 (O_3,N_19645,N_19029);
or UO_4 (O_4,N_19914,N_19680);
or UO_5 (O_5,N_19219,N_19589);
or UO_6 (O_6,N_19274,N_19804);
nor UO_7 (O_7,N_19245,N_19170);
and UO_8 (O_8,N_19660,N_19685);
and UO_9 (O_9,N_19407,N_19421);
or UO_10 (O_10,N_19146,N_19555);
and UO_11 (O_11,N_19494,N_19635);
xnor UO_12 (O_12,N_19431,N_19710);
or UO_13 (O_13,N_19725,N_19567);
nand UO_14 (O_14,N_19639,N_19846);
xor UO_15 (O_15,N_19736,N_19876);
xor UO_16 (O_16,N_19483,N_19998);
nor UO_17 (O_17,N_19770,N_19180);
nor UO_18 (O_18,N_19528,N_19491);
nand UO_19 (O_19,N_19350,N_19132);
or UO_20 (O_20,N_19993,N_19949);
or UO_21 (O_21,N_19349,N_19739);
or UO_22 (O_22,N_19664,N_19301);
or UO_23 (O_23,N_19189,N_19723);
or UO_24 (O_24,N_19936,N_19800);
xor UO_25 (O_25,N_19294,N_19355);
nand UO_26 (O_26,N_19403,N_19977);
nand UO_27 (O_27,N_19580,N_19394);
and UO_28 (O_28,N_19133,N_19161);
nor UO_29 (O_29,N_19741,N_19776);
nor UO_30 (O_30,N_19514,N_19588);
and UO_31 (O_31,N_19925,N_19707);
and UO_32 (O_32,N_19320,N_19693);
xor UO_33 (O_33,N_19651,N_19466);
nand UO_34 (O_34,N_19190,N_19401);
nand UO_35 (O_35,N_19318,N_19726);
nor UO_36 (O_36,N_19969,N_19308);
xor UO_37 (O_37,N_19072,N_19338);
or UO_38 (O_38,N_19211,N_19802);
nand UO_39 (O_39,N_19337,N_19326);
nand UO_40 (O_40,N_19005,N_19542);
or UO_41 (O_41,N_19445,N_19507);
or UO_42 (O_42,N_19862,N_19478);
xor UO_43 (O_43,N_19922,N_19851);
nor UO_44 (O_44,N_19314,N_19109);
nand UO_45 (O_45,N_19408,N_19263);
xnor UO_46 (O_46,N_19480,N_19481);
and UO_47 (O_47,N_19857,N_19637);
nor UO_48 (O_48,N_19044,N_19402);
nand UO_49 (O_49,N_19997,N_19387);
and UO_50 (O_50,N_19533,N_19961);
nor UO_51 (O_51,N_19046,N_19575);
xor UO_52 (O_52,N_19400,N_19142);
or UO_53 (O_53,N_19617,N_19957);
xor UO_54 (O_54,N_19796,N_19539);
or UO_55 (O_55,N_19573,N_19614);
nor UO_56 (O_56,N_19469,N_19447);
nand UO_57 (O_57,N_19593,N_19935);
or UO_58 (O_58,N_19926,N_19098);
or UO_59 (O_59,N_19782,N_19248);
xnor UO_60 (O_60,N_19310,N_19819);
and UO_61 (O_61,N_19893,N_19476);
xor UO_62 (O_62,N_19939,N_19856);
or UO_63 (O_63,N_19655,N_19284);
and UO_64 (O_64,N_19689,N_19388);
nor UO_65 (O_65,N_19092,N_19143);
or UO_66 (O_66,N_19041,N_19026);
and UO_67 (O_67,N_19502,N_19743);
and UO_68 (O_68,N_19891,N_19004);
xnor UO_69 (O_69,N_19526,N_19759);
or UO_70 (O_70,N_19049,N_19264);
nor UO_71 (O_71,N_19232,N_19195);
xnor UO_72 (O_72,N_19106,N_19391);
nand UO_73 (O_73,N_19968,N_19485);
nor UO_74 (O_74,N_19442,N_19894);
xnor UO_75 (O_75,N_19592,N_19799);
xor UO_76 (O_76,N_19951,N_19569);
xnor UO_77 (O_77,N_19608,N_19147);
nor UO_78 (O_78,N_19169,N_19873);
xnor UO_79 (O_79,N_19410,N_19538);
and UO_80 (O_80,N_19972,N_19917);
nor UO_81 (O_81,N_19241,N_19631);
or UO_82 (O_82,N_19424,N_19684);
nand UO_83 (O_83,N_19229,N_19192);
nor UO_84 (O_84,N_19446,N_19050);
or UO_85 (O_85,N_19059,N_19701);
xor UO_86 (O_86,N_19669,N_19080);
nand UO_87 (O_87,N_19420,N_19121);
and UO_88 (O_88,N_19602,N_19215);
or UO_89 (O_89,N_19768,N_19316);
and UO_90 (O_90,N_19305,N_19227);
or UO_91 (O_91,N_19534,N_19766);
nand UO_92 (O_92,N_19489,N_19027);
nor UO_93 (O_93,N_19508,N_19166);
nor UO_94 (O_94,N_19913,N_19299);
or UO_95 (O_95,N_19666,N_19762);
nor UO_96 (O_96,N_19596,N_19735);
and UO_97 (O_97,N_19647,N_19490);
nand UO_98 (O_98,N_19619,N_19641);
xnor UO_99 (O_99,N_19482,N_19249);
nor UO_100 (O_100,N_19709,N_19942);
and UO_101 (O_101,N_19681,N_19979);
or UO_102 (O_102,N_19501,N_19373);
xor UO_103 (O_103,N_19174,N_19985);
nor UO_104 (O_104,N_19927,N_19761);
nor UO_105 (O_105,N_19820,N_19676);
nor UO_106 (O_106,N_19493,N_19946);
xor UO_107 (O_107,N_19611,N_19730);
xnor UO_108 (O_108,N_19235,N_19495);
xnor UO_109 (O_109,N_19467,N_19858);
and UO_110 (O_110,N_19734,N_19148);
and UO_111 (O_111,N_19019,N_19042);
nor UO_112 (O_112,N_19065,N_19714);
nor UO_113 (O_113,N_19784,N_19070);
and UO_114 (O_114,N_19456,N_19071);
and UO_115 (O_115,N_19090,N_19982);
nor UO_116 (O_116,N_19869,N_19053);
or UO_117 (O_117,N_19329,N_19035);
or UO_118 (O_118,N_19771,N_19716);
nor UO_119 (O_119,N_19398,N_19022);
nor UO_120 (O_120,N_19656,N_19540);
and UO_121 (O_121,N_19559,N_19433);
or UO_122 (O_122,N_19545,N_19976);
nand UO_123 (O_123,N_19034,N_19111);
or UO_124 (O_124,N_19001,N_19067);
and UO_125 (O_125,N_19124,N_19187);
or UO_126 (O_126,N_19191,N_19535);
and UO_127 (O_127,N_19809,N_19564);
xnor UO_128 (O_128,N_19943,N_19156);
or UO_129 (O_129,N_19811,N_19667);
xnor UO_130 (O_130,N_19956,N_19341);
xnor UO_131 (O_131,N_19319,N_19607);
xor UO_132 (O_132,N_19342,N_19921);
xnor UO_133 (O_133,N_19082,N_19722);
or UO_134 (O_134,N_19585,N_19074);
xor UO_135 (O_135,N_19638,N_19966);
xnor UO_136 (O_136,N_19986,N_19778);
nand UO_137 (O_137,N_19268,N_19687);
nand UO_138 (O_138,N_19878,N_19874);
xnor UO_139 (O_139,N_19464,N_19554);
and UO_140 (O_140,N_19854,N_19868);
or UO_141 (O_141,N_19813,N_19753);
and UO_142 (O_142,N_19713,N_19162);
xor UO_143 (O_143,N_19983,N_19783);
xor UO_144 (O_144,N_19282,N_19313);
or UO_145 (O_145,N_19965,N_19068);
nor UO_146 (O_146,N_19863,N_19231);
or UO_147 (O_147,N_19824,N_19731);
and UO_148 (O_148,N_19193,N_19210);
or UO_149 (O_149,N_19995,N_19934);
nor UO_150 (O_150,N_19706,N_19733);
nor UO_151 (O_151,N_19742,N_19422);
or UO_152 (O_152,N_19060,N_19024);
nor UO_153 (O_153,N_19774,N_19910);
nand UO_154 (O_154,N_19586,N_19529);
nand UO_155 (O_155,N_19441,N_19176);
nor UO_156 (O_156,N_19242,N_19119);
and UO_157 (O_157,N_19902,N_19702);
nand UO_158 (O_158,N_19703,N_19890);
nand UO_159 (O_159,N_19786,N_19428);
and UO_160 (O_160,N_19964,N_19099);
or UO_161 (O_161,N_19157,N_19978);
nand UO_162 (O_162,N_19247,N_19275);
xor UO_163 (O_163,N_19371,N_19785);
or UO_164 (O_164,N_19841,N_19419);
nand UO_165 (O_165,N_19389,N_19039);
nor UO_166 (O_166,N_19165,N_19945);
and UO_167 (O_167,N_19801,N_19110);
nor UO_168 (O_168,N_19947,N_19405);
and UO_169 (O_169,N_19918,N_19375);
and UO_170 (O_170,N_19788,N_19272);
or UO_171 (O_171,N_19845,N_19999);
nand UO_172 (O_172,N_19128,N_19454);
nand UO_173 (O_173,N_19045,N_19828);
or UO_174 (O_174,N_19852,N_19652);
and UO_175 (O_175,N_19087,N_19201);
xnor UO_176 (O_176,N_19425,N_19740);
xnor UO_177 (O_177,N_19105,N_19458);
or UO_178 (O_178,N_19861,N_19412);
nand UO_179 (O_179,N_19830,N_19167);
or UO_180 (O_180,N_19043,N_19246);
nand UO_181 (O_181,N_19054,N_19295);
and UO_182 (O_182,N_19817,N_19769);
or UO_183 (O_183,N_19336,N_19806);
nand UO_184 (O_184,N_19537,N_19896);
nor UO_185 (O_185,N_19088,N_19640);
xnor UO_186 (O_186,N_19720,N_19780);
and UO_187 (O_187,N_19552,N_19395);
nand UO_188 (O_188,N_19291,N_19217);
nor UO_189 (O_189,N_19240,N_19807);
xnor UO_190 (O_190,N_19136,N_19056);
nand UO_191 (O_191,N_19279,N_19306);
or UO_192 (O_192,N_19871,N_19882);
nand UO_193 (O_193,N_19598,N_19565);
or UO_194 (O_194,N_19516,N_19627);
nor UO_195 (O_195,N_19816,N_19787);
nand UO_196 (O_196,N_19037,N_19673);
nand UO_197 (O_197,N_19557,N_19522);
nand UO_198 (O_198,N_19351,N_19909);
or UO_199 (O_199,N_19453,N_19629);
nand UO_200 (O_200,N_19950,N_19153);
xnor UO_201 (O_201,N_19257,N_19175);
and UO_202 (O_202,N_19171,N_19550);
and UO_203 (O_203,N_19737,N_19524);
nand UO_204 (O_204,N_19948,N_19113);
and UO_205 (O_205,N_19286,N_19228);
xnor UO_206 (O_206,N_19302,N_19324);
or UO_207 (O_207,N_19665,N_19962);
or UO_208 (O_208,N_19623,N_19886);
or UO_209 (O_209,N_19475,N_19530);
nand UO_210 (O_210,N_19512,N_19287);
nor UO_211 (O_211,N_19527,N_19462);
xnor UO_212 (O_212,N_19277,N_19758);
nand UO_213 (O_213,N_19877,N_19061);
nor UO_214 (O_214,N_19487,N_19825);
xor UO_215 (O_215,N_19590,N_19497);
and UO_216 (O_216,N_19202,N_19595);
xor UO_217 (O_217,N_19085,N_19578);
nand UO_218 (O_218,N_19293,N_19864);
or UO_219 (O_219,N_19510,N_19657);
or UO_220 (O_220,N_19653,N_19505);
nand UO_221 (O_221,N_19831,N_19610);
nor UO_222 (O_222,N_19691,N_19859);
xor UO_223 (O_223,N_19380,N_19298);
nand UO_224 (O_224,N_19304,N_19131);
nor UO_225 (O_225,N_19973,N_19003);
nor UO_226 (O_226,N_19523,N_19810);
nand UO_227 (O_227,N_19411,N_19536);
nand UO_228 (O_228,N_19519,N_19836);
nand UO_229 (O_229,N_19152,N_19429);
or UO_230 (O_230,N_19755,N_19233);
xor UO_231 (O_231,N_19750,N_19362);
nor UO_232 (O_232,N_19430,N_19568);
nor UO_233 (O_233,N_19712,N_19690);
xor UO_234 (O_234,N_19057,N_19205);
xnor UO_235 (O_235,N_19333,N_19853);
and UO_236 (O_236,N_19449,N_19815);
xor UO_237 (O_237,N_19718,N_19963);
nor UO_238 (O_238,N_19584,N_19339);
or UO_239 (O_239,N_19239,N_19721);
and UO_240 (O_240,N_19376,N_19630);
or UO_241 (O_241,N_19311,N_19079);
or UO_242 (O_242,N_19423,N_19102);
xnor UO_243 (O_243,N_19374,N_19347);
nand UO_244 (O_244,N_19181,N_19149);
and UO_245 (O_245,N_19895,N_19618);
xnor UO_246 (O_246,N_19020,N_19500);
nand UO_247 (O_247,N_19254,N_19805);
xor UO_248 (O_248,N_19765,N_19354);
nor UO_249 (O_249,N_19236,N_19560);
and UO_250 (O_250,N_19426,N_19448);
and UO_251 (O_251,N_19107,N_19620);
and UO_252 (O_252,N_19566,N_19151);
nor UO_253 (O_253,N_19207,N_19484);
and UO_254 (O_254,N_19016,N_19437);
and UO_255 (O_255,N_19808,N_19708);
xnor UO_256 (O_256,N_19971,N_19238);
nand UO_257 (O_257,N_19541,N_19358);
or UO_258 (O_258,N_19463,N_19159);
and UO_259 (O_259,N_19897,N_19138);
and UO_260 (O_260,N_19221,N_19276);
nor UO_261 (O_261,N_19738,N_19717);
and UO_262 (O_262,N_19797,N_19790);
nor UO_263 (O_263,N_19571,N_19970);
or UO_264 (O_264,N_19069,N_19084);
nor UO_265 (O_265,N_19129,N_19518);
nand UO_266 (O_266,N_19827,N_19532);
and UO_267 (O_267,N_19317,N_19609);
and UO_268 (O_268,N_19014,N_19081);
or UO_269 (O_269,N_19255,N_19220);
nor UO_270 (O_270,N_19066,N_19646);
xor UO_271 (O_271,N_19370,N_19021);
nor UO_272 (O_272,N_19872,N_19118);
and UO_273 (O_273,N_19729,N_19688);
nor UO_274 (O_274,N_19504,N_19929);
and UO_275 (O_275,N_19867,N_19615);
xnor UO_276 (O_276,N_19551,N_19889);
or UO_277 (O_277,N_19616,N_19297);
and UO_278 (O_278,N_19002,N_19125);
or UO_279 (O_279,N_19103,N_19377);
nand UO_280 (O_280,N_19732,N_19984);
and UO_281 (O_281,N_19506,N_19763);
nor UO_282 (O_282,N_19661,N_19218);
and UO_283 (O_283,N_19775,N_19648);
and UO_284 (O_284,N_19335,N_19840);
nor UO_285 (O_285,N_19887,N_19940);
nand UO_286 (O_286,N_19100,N_19793);
nand UO_287 (O_287,N_19679,N_19990);
and UO_288 (O_288,N_19383,N_19040);
nand UO_289 (O_289,N_19260,N_19622);
and UO_290 (O_290,N_19671,N_19017);
xnor UO_291 (O_291,N_19850,N_19328);
or UO_292 (O_292,N_19916,N_19579);
xor UO_293 (O_293,N_19322,N_19773);
xor UO_294 (O_294,N_19803,N_19757);
nand UO_295 (O_295,N_19572,N_19015);
or UO_296 (O_296,N_19699,N_19209);
nor UO_297 (O_297,N_19285,N_19381);
or UO_298 (O_298,N_19674,N_19860);
or UO_299 (O_299,N_19694,N_19188);
nand UO_300 (O_300,N_19791,N_19839);
xor UO_301 (O_301,N_19468,N_19222);
nand UO_302 (O_302,N_19473,N_19032);
nor UO_303 (O_303,N_19006,N_19499);
nand UO_304 (O_304,N_19392,N_19382);
nor UO_305 (O_305,N_19327,N_19944);
nor UO_306 (O_306,N_19583,N_19443);
xnor UO_307 (O_307,N_19980,N_19632);
xnor UO_308 (O_308,N_19789,N_19278);
nand UO_309 (O_309,N_19140,N_19288);
nor UO_310 (O_310,N_19633,N_19751);
nor UO_311 (O_311,N_19814,N_19884);
xnor UO_312 (O_312,N_19312,N_19353);
nor UO_313 (O_313,N_19108,N_19393);
and UO_314 (O_314,N_19521,N_19465);
nand UO_315 (O_315,N_19052,N_19745);
or UO_316 (O_316,N_19030,N_19139);
xor UO_317 (O_317,N_19928,N_19352);
nor UO_318 (O_318,N_19332,N_19628);
and UO_319 (O_319,N_19346,N_19991);
and UO_320 (O_320,N_19436,N_19435);
or UO_321 (O_321,N_19920,N_19952);
xnor UO_322 (O_322,N_19933,N_19517);
xor UO_323 (O_323,N_19083,N_19182);
or UO_324 (O_324,N_19855,N_19603);
nand UO_325 (O_325,N_19062,N_19256);
or UO_326 (O_326,N_19273,N_19958);
nor UO_327 (O_327,N_19649,N_19197);
nor UO_328 (O_328,N_19698,N_19835);
nor UO_329 (O_329,N_19230,N_19204);
and UO_330 (O_330,N_19163,N_19636);
and UO_331 (O_331,N_19697,N_19911);
xnor UO_332 (O_332,N_19267,N_19621);
xor UO_333 (O_333,N_19912,N_19091);
xnor UO_334 (O_334,N_19104,N_19659);
or UO_335 (O_335,N_19258,N_19460);
nand UO_336 (O_336,N_19179,N_19472);
nand UO_337 (O_337,N_19283,N_19144);
or UO_338 (O_338,N_19549,N_19413);
nor UO_339 (O_339,N_19826,N_19018);
xnor UO_340 (O_340,N_19658,N_19344);
nor UO_341 (O_341,N_19281,N_19767);
nand UO_342 (O_342,N_19094,N_19558);
and UO_343 (O_343,N_19941,N_19073);
xor UO_344 (O_344,N_19172,N_19821);
nand UO_345 (O_345,N_19634,N_19838);
nor UO_346 (O_346,N_19866,N_19543);
and UO_347 (O_347,N_19334,N_19503);
xor UO_348 (O_348,N_19955,N_19309);
or UO_349 (O_349,N_19194,N_19642);
or UO_350 (O_350,N_19892,N_19682);
or UO_351 (O_351,N_19781,N_19544);
or UO_352 (O_352,N_19954,N_19183);
xor UO_353 (O_353,N_19988,N_19792);
nor UO_354 (O_354,N_19009,N_19368);
nand UO_355 (O_355,N_19012,N_19663);
xor UO_356 (O_356,N_19471,N_19064);
nor UO_357 (O_357,N_19315,N_19123);
nand UO_358 (O_358,N_19626,N_19498);
xor UO_359 (O_359,N_19325,N_19719);
nor UO_360 (O_360,N_19879,N_19923);
and UO_361 (O_361,N_19601,N_19974);
xnor UO_362 (O_362,N_19843,N_19457);
xor UO_363 (O_363,N_19168,N_19396);
nand UO_364 (O_364,N_19496,N_19265);
and UO_365 (O_365,N_19086,N_19127);
and UO_366 (O_366,N_19880,N_19900);
nor UO_367 (O_367,N_19416,N_19677);
and UO_368 (O_368,N_19023,N_19063);
and UO_369 (O_369,N_19008,N_19292);
and UO_370 (O_370,N_19606,N_19137);
xor UO_371 (O_371,N_19114,N_19372);
xnor UO_372 (O_372,N_19672,N_19531);
xor UO_373 (O_373,N_19678,N_19348);
nand UO_374 (O_374,N_19754,N_19477);
and UO_375 (O_375,N_19130,N_19078);
nor UO_376 (O_376,N_19613,N_19440);
nor UO_377 (O_377,N_19705,N_19812);
and UO_378 (O_378,N_19777,N_19844);
nor UO_379 (O_379,N_19270,N_19899);
or UO_380 (O_380,N_19290,N_19390);
nor UO_381 (O_381,N_19199,N_19562);
and UO_382 (O_382,N_19888,N_19818);
nand UO_383 (O_383,N_19520,N_19384);
or UO_384 (O_384,N_19379,N_19055);
and UO_385 (O_385,N_19244,N_19361);
nand UO_386 (O_386,N_19794,N_19903);
nand UO_387 (O_387,N_19459,N_19591);
nor UO_388 (O_388,N_19904,N_19206);
nand UO_389 (O_389,N_19415,N_19600);
xor UO_390 (O_390,N_19832,N_19605);
nand UO_391 (O_391,N_19488,N_19077);
xor UO_392 (O_392,N_19451,N_19574);
xnor UO_393 (O_393,N_19967,N_19266);
xor UO_394 (O_394,N_19216,N_19919);
nor UO_395 (O_395,N_19749,N_19007);
nand UO_396 (O_396,N_19515,N_19668);
nand UO_397 (O_397,N_19624,N_19747);
nor UO_398 (O_398,N_19905,N_19164);
nor UO_399 (O_399,N_19764,N_19200);
or UO_400 (O_400,N_19849,N_19363);
xor UO_401 (O_401,N_19924,N_19289);
xor UO_402 (O_402,N_19570,N_19406);
nand UO_403 (O_403,N_19875,N_19427);
xnor UO_404 (O_404,N_19261,N_19937);
or UO_405 (O_405,N_19321,N_19259);
or UO_406 (O_406,N_19696,N_19834);
nor UO_407 (O_407,N_19173,N_19604);
xnor UO_408 (O_408,N_19576,N_19213);
nor UO_409 (O_409,N_19076,N_19025);
or UO_410 (O_410,N_19033,N_19096);
or UO_411 (O_411,N_19262,N_19695);
nor UO_412 (O_412,N_19135,N_19196);
xnor UO_413 (O_413,N_19343,N_19010);
and UO_414 (O_414,N_19367,N_19582);
and UO_415 (O_415,N_19746,N_19058);
xnor UO_416 (O_416,N_19748,N_19345);
nor UO_417 (O_417,N_19744,N_19612);
nand UO_418 (O_418,N_19439,N_19901);
nor UO_419 (O_419,N_19994,N_19975);
nor UO_420 (O_420,N_19728,N_19364);
nand UO_421 (O_421,N_19145,N_19870);
or UO_422 (O_422,N_19548,N_19865);
xnor UO_423 (O_423,N_19906,N_19455);
xnor UO_424 (O_424,N_19959,N_19048);
or UO_425 (O_425,N_19883,N_19644);
xnor UO_426 (O_426,N_19546,N_19432);
or UO_427 (O_427,N_19158,N_19450);
xnor UO_428 (O_428,N_19331,N_19154);
xnor UO_429 (O_429,N_19960,N_19126);
xnor UO_430 (O_430,N_19177,N_19307);
nand UO_431 (O_431,N_19452,N_19386);
xor UO_432 (O_432,N_19438,N_19915);
and UO_433 (O_433,N_19134,N_19587);
xor UO_434 (O_434,N_19795,N_19237);
or UO_435 (O_435,N_19989,N_19296);
xor UO_436 (O_436,N_19417,N_19185);
nor UO_437 (O_437,N_19093,N_19662);
nor UO_438 (O_438,N_19198,N_19178);
nand UO_439 (O_439,N_19155,N_19101);
xor UO_440 (O_440,N_19837,N_19252);
nand UO_441 (O_441,N_19898,N_19885);
and UO_442 (O_442,N_19075,N_19366);
xor UO_443 (O_443,N_19938,N_19654);
nor UO_444 (O_444,N_19116,N_19577);
or UO_445 (O_445,N_19594,N_19479);
or UO_446 (O_446,N_19444,N_19829);
nor UO_447 (O_447,N_19397,N_19798);
xnor UO_448 (O_448,N_19385,N_19409);
nor UO_449 (O_449,N_19226,N_19280);
nand UO_450 (O_450,N_19330,N_19115);
nand UO_451 (O_451,N_19847,N_19160);
nor UO_452 (O_452,N_19097,N_19842);
or UO_453 (O_453,N_19996,N_19563);
and UO_454 (O_454,N_19556,N_19112);
xnor UO_455 (O_455,N_19643,N_19931);
nand UO_456 (O_456,N_19881,N_19987);
xor UO_457 (O_457,N_19122,N_19365);
and UO_458 (O_458,N_19513,N_19547);
and UO_459 (O_459,N_19907,N_19760);
or UO_460 (O_460,N_19704,N_19223);
nand UO_461 (O_461,N_19038,N_19414);
or UO_462 (O_462,N_19461,N_19700);
xor UO_463 (O_463,N_19492,N_19028);
nor UO_464 (O_464,N_19597,N_19300);
nand UO_465 (O_465,N_19243,N_19212);
xnor UO_466 (O_466,N_19599,N_19225);
and UO_467 (O_467,N_19908,N_19253);
nand UO_468 (O_468,N_19117,N_19359);
nand UO_469 (O_469,N_19715,N_19675);
nand UO_470 (O_470,N_19992,N_19525);
and UO_471 (O_471,N_19470,N_19271);
nor UO_472 (O_472,N_19981,N_19724);
nor UO_473 (O_473,N_19932,N_19224);
nand UO_474 (O_474,N_19051,N_19186);
nor UO_475 (O_475,N_19848,N_19303);
xnor UO_476 (O_476,N_19474,N_19683);
and UO_477 (O_477,N_19727,N_19095);
or UO_478 (O_478,N_19772,N_19692);
nand UO_479 (O_479,N_19779,N_19150);
and UO_480 (O_480,N_19930,N_19434);
xnor UO_481 (O_481,N_19000,N_19141);
or UO_482 (O_482,N_19120,N_19833);
nor UO_483 (O_483,N_19013,N_19250);
nand UO_484 (O_484,N_19625,N_19214);
xor UO_485 (O_485,N_19031,N_19269);
and UO_486 (O_486,N_19752,N_19208);
nor UO_487 (O_487,N_19251,N_19511);
nor UO_488 (O_488,N_19340,N_19418);
and UO_489 (O_489,N_19360,N_19036);
or UO_490 (O_490,N_19356,N_19399);
and UO_491 (O_491,N_19670,N_19404);
xnor UO_492 (O_492,N_19581,N_19650);
or UO_493 (O_493,N_19822,N_19553);
xor UO_494 (O_494,N_19323,N_19823);
and UO_495 (O_495,N_19047,N_19011);
or UO_496 (O_496,N_19486,N_19089);
nand UO_497 (O_497,N_19953,N_19203);
xor UO_498 (O_498,N_19509,N_19561);
nor UO_499 (O_499,N_19711,N_19369);
and UO_500 (O_500,N_19422,N_19259);
nor UO_501 (O_501,N_19376,N_19643);
xnor UO_502 (O_502,N_19620,N_19100);
or UO_503 (O_503,N_19786,N_19733);
and UO_504 (O_504,N_19796,N_19697);
xor UO_505 (O_505,N_19178,N_19998);
and UO_506 (O_506,N_19287,N_19173);
nor UO_507 (O_507,N_19625,N_19518);
xnor UO_508 (O_508,N_19826,N_19072);
nor UO_509 (O_509,N_19014,N_19401);
xor UO_510 (O_510,N_19585,N_19730);
nand UO_511 (O_511,N_19736,N_19254);
nor UO_512 (O_512,N_19958,N_19628);
or UO_513 (O_513,N_19360,N_19272);
or UO_514 (O_514,N_19087,N_19795);
or UO_515 (O_515,N_19295,N_19091);
xnor UO_516 (O_516,N_19287,N_19446);
nand UO_517 (O_517,N_19369,N_19882);
or UO_518 (O_518,N_19973,N_19563);
xnor UO_519 (O_519,N_19007,N_19728);
nand UO_520 (O_520,N_19722,N_19075);
nor UO_521 (O_521,N_19000,N_19280);
or UO_522 (O_522,N_19021,N_19777);
xnor UO_523 (O_523,N_19437,N_19367);
or UO_524 (O_524,N_19669,N_19633);
nand UO_525 (O_525,N_19967,N_19903);
or UO_526 (O_526,N_19809,N_19953);
nand UO_527 (O_527,N_19165,N_19680);
and UO_528 (O_528,N_19320,N_19316);
or UO_529 (O_529,N_19521,N_19610);
xnor UO_530 (O_530,N_19643,N_19519);
nor UO_531 (O_531,N_19329,N_19851);
nand UO_532 (O_532,N_19219,N_19047);
nor UO_533 (O_533,N_19313,N_19465);
and UO_534 (O_534,N_19957,N_19778);
nor UO_535 (O_535,N_19995,N_19556);
nor UO_536 (O_536,N_19057,N_19680);
nor UO_537 (O_537,N_19993,N_19400);
nand UO_538 (O_538,N_19998,N_19822);
nand UO_539 (O_539,N_19295,N_19221);
or UO_540 (O_540,N_19708,N_19806);
nor UO_541 (O_541,N_19828,N_19784);
and UO_542 (O_542,N_19950,N_19676);
and UO_543 (O_543,N_19318,N_19841);
or UO_544 (O_544,N_19858,N_19093);
nand UO_545 (O_545,N_19085,N_19546);
nand UO_546 (O_546,N_19557,N_19409);
nand UO_547 (O_547,N_19064,N_19612);
or UO_548 (O_548,N_19592,N_19562);
and UO_549 (O_549,N_19483,N_19605);
nand UO_550 (O_550,N_19300,N_19303);
nand UO_551 (O_551,N_19424,N_19067);
and UO_552 (O_552,N_19015,N_19261);
and UO_553 (O_553,N_19961,N_19875);
nand UO_554 (O_554,N_19076,N_19938);
or UO_555 (O_555,N_19713,N_19957);
nand UO_556 (O_556,N_19640,N_19193);
nor UO_557 (O_557,N_19639,N_19565);
nor UO_558 (O_558,N_19724,N_19551);
nand UO_559 (O_559,N_19533,N_19145);
or UO_560 (O_560,N_19646,N_19510);
nor UO_561 (O_561,N_19010,N_19566);
xnor UO_562 (O_562,N_19261,N_19003);
nand UO_563 (O_563,N_19132,N_19503);
nand UO_564 (O_564,N_19622,N_19270);
and UO_565 (O_565,N_19174,N_19690);
nand UO_566 (O_566,N_19358,N_19620);
xnor UO_567 (O_567,N_19509,N_19130);
or UO_568 (O_568,N_19793,N_19456);
xnor UO_569 (O_569,N_19208,N_19019);
and UO_570 (O_570,N_19817,N_19614);
or UO_571 (O_571,N_19881,N_19519);
or UO_572 (O_572,N_19071,N_19213);
nor UO_573 (O_573,N_19049,N_19429);
nor UO_574 (O_574,N_19701,N_19791);
and UO_575 (O_575,N_19184,N_19090);
and UO_576 (O_576,N_19018,N_19751);
nand UO_577 (O_577,N_19059,N_19036);
nand UO_578 (O_578,N_19913,N_19688);
nor UO_579 (O_579,N_19893,N_19220);
nor UO_580 (O_580,N_19525,N_19829);
nand UO_581 (O_581,N_19224,N_19319);
or UO_582 (O_582,N_19222,N_19654);
and UO_583 (O_583,N_19189,N_19955);
nor UO_584 (O_584,N_19959,N_19783);
or UO_585 (O_585,N_19341,N_19612);
and UO_586 (O_586,N_19368,N_19717);
xor UO_587 (O_587,N_19164,N_19503);
nor UO_588 (O_588,N_19429,N_19680);
and UO_589 (O_589,N_19469,N_19424);
or UO_590 (O_590,N_19578,N_19777);
or UO_591 (O_591,N_19955,N_19027);
or UO_592 (O_592,N_19015,N_19001);
or UO_593 (O_593,N_19214,N_19133);
and UO_594 (O_594,N_19113,N_19592);
or UO_595 (O_595,N_19378,N_19263);
nand UO_596 (O_596,N_19510,N_19157);
xor UO_597 (O_597,N_19584,N_19503);
and UO_598 (O_598,N_19672,N_19681);
nand UO_599 (O_599,N_19994,N_19774);
nand UO_600 (O_600,N_19550,N_19090);
xor UO_601 (O_601,N_19064,N_19734);
nand UO_602 (O_602,N_19299,N_19635);
xor UO_603 (O_603,N_19210,N_19435);
nand UO_604 (O_604,N_19705,N_19219);
xor UO_605 (O_605,N_19625,N_19767);
nor UO_606 (O_606,N_19912,N_19079);
xor UO_607 (O_607,N_19819,N_19632);
or UO_608 (O_608,N_19755,N_19425);
or UO_609 (O_609,N_19644,N_19042);
xor UO_610 (O_610,N_19246,N_19536);
and UO_611 (O_611,N_19432,N_19246);
xnor UO_612 (O_612,N_19828,N_19430);
or UO_613 (O_613,N_19479,N_19860);
or UO_614 (O_614,N_19790,N_19111);
and UO_615 (O_615,N_19303,N_19881);
or UO_616 (O_616,N_19397,N_19555);
and UO_617 (O_617,N_19434,N_19509);
nand UO_618 (O_618,N_19918,N_19294);
and UO_619 (O_619,N_19620,N_19059);
xor UO_620 (O_620,N_19464,N_19503);
or UO_621 (O_621,N_19842,N_19643);
xnor UO_622 (O_622,N_19730,N_19064);
nand UO_623 (O_623,N_19883,N_19684);
or UO_624 (O_624,N_19236,N_19207);
xor UO_625 (O_625,N_19190,N_19743);
or UO_626 (O_626,N_19551,N_19522);
nand UO_627 (O_627,N_19789,N_19157);
and UO_628 (O_628,N_19964,N_19942);
or UO_629 (O_629,N_19444,N_19174);
xor UO_630 (O_630,N_19916,N_19208);
xnor UO_631 (O_631,N_19923,N_19402);
nor UO_632 (O_632,N_19803,N_19907);
nor UO_633 (O_633,N_19787,N_19614);
or UO_634 (O_634,N_19899,N_19828);
nand UO_635 (O_635,N_19832,N_19812);
nand UO_636 (O_636,N_19196,N_19537);
xor UO_637 (O_637,N_19438,N_19920);
or UO_638 (O_638,N_19964,N_19687);
nor UO_639 (O_639,N_19891,N_19111);
nor UO_640 (O_640,N_19002,N_19267);
nand UO_641 (O_641,N_19735,N_19327);
nand UO_642 (O_642,N_19072,N_19444);
nand UO_643 (O_643,N_19338,N_19220);
xor UO_644 (O_644,N_19985,N_19352);
and UO_645 (O_645,N_19897,N_19539);
nor UO_646 (O_646,N_19193,N_19055);
and UO_647 (O_647,N_19142,N_19551);
or UO_648 (O_648,N_19786,N_19783);
and UO_649 (O_649,N_19917,N_19596);
nor UO_650 (O_650,N_19608,N_19165);
and UO_651 (O_651,N_19349,N_19237);
xnor UO_652 (O_652,N_19937,N_19547);
or UO_653 (O_653,N_19362,N_19075);
nor UO_654 (O_654,N_19909,N_19605);
xnor UO_655 (O_655,N_19011,N_19999);
or UO_656 (O_656,N_19590,N_19937);
or UO_657 (O_657,N_19297,N_19174);
nor UO_658 (O_658,N_19770,N_19545);
nor UO_659 (O_659,N_19883,N_19392);
or UO_660 (O_660,N_19427,N_19785);
or UO_661 (O_661,N_19746,N_19155);
nor UO_662 (O_662,N_19897,N_19506);
xor UO_663 (O_663,N_19122,N_19795);
nand UO_664 (O_664,N_19361,N_19060);
or UO_665 (O_665,N_19154,N_19094);
and UO_666 (O_666,N_19775,N_19779);
xnor UO_667 (O_667,N_19575,N_19803);
xnor UO_668 (O_668,N_19679,N_19781);
or UO_669 (O_669,N_19405,N_19064);
and UO_670 (O_670,N_19016,N_19512);
xnor UO_671 (O_671,N_19955,N_19292);
nor UO_672 (O_672,N_19944,N_19684);
nor UO_673 (O_673,N_19479,N_19721);
xor UO_674 (O_674,N_19530,N_19608);
or UO_675 (O_675,N_19450,N_19406);
and UO_676 (O_676,N_19782,N_19585);
or UO_677 (O_677,N_19750,N_19458);
nand UO_678 (O_678,N_19858,N_19376);
nand UO_679 (O_679,N_19577,N_19222);
nor UO_680 (O_680,N_19974,N_19462);
nand UO_681 (O_681,N_19515,N_19695);
or UO_682 (O_682,N_19813,N_19510);
xnor UO_683 (O_683,N_19029,N_19446);
and UO_684 (O_684,N_19129,N_19063);
and UO_685 (O_685,N_19701,N_19391);
nand UO_686 (O_686,N_19140,N_19146);
and UO_687 (O_687,N_19592,N_19432);
xor UO_688 (O_688,N_19340,N_19590);
nand UO_689 (O_689,N_19852,N_19730);
xnor UO_690 (O_690,N_19945,N_19245);
xor UO_691 (O_691,N_19170,N_19246);
or UO_692 (O_692,N_19354,N_19867);
nor UO_693 (O_693,N_19282,N_19193);
or UO_694 (O_694,N_19376,N_19863);
and UO_695 (O_695,N_19280,N_19166);
and UO_696 (O_696,N_19497,N_19958);
or UO_697 (O_697,N_19820,N_19273);
xor UO_698 (O_698,N_19534,N_19457);
or UO_699 (O_699,N_19574,N_19703);
or UO_700 (O_700,N_19373,N_19114);
and UO_701 (O_701,N_19570,N_19481);
nor UO_702 (O_702,N_19201,N_19945);
nor UO_703 (O_703,N_19433,N_19753);
or UO_704 (O_704,N_19165,N_19161);
xor UO_705 (O_705,N_19698,N_19450);
nor UO_706 (O_706,N_19475,N_19179);
and UO_707 (O_707,N_19054,N_19099);
nor UO_708 (O_708,N_19188,N_19693);
nor UO_709 (O_709,N_19635,N_19450);
nand UO_710 (O_710,N_19175,N_19085);
xnor UO_711 (O_711,N_19322,N_19856);
nor UO_712 (O_712,N_19997,N_19543);
and UO_713 (O_713,N_19352,N_19647);
and UO_714 (O_714,N_19192,N_19878);
and UO_715 (O_715,N_19755,N_19601);
nand UO_716 (O_716,N_19926,N_19703);
or UO_717 (O_717,N_19649,N_19057);
and UO_718 (O_718,N_19892,N_19129);
xor UO_719 (O_719,N_19347,N_19647);
nand UO_720 (O_720,N_19929,N_19054);
or UO_721 (O_721,N_19456,N_19902);
nand UO_722 (O_722,N_19990,N_19085);
nand UO_723 (O_723,N_19472,N_19595);
and UO_724 (O_724,N_19638,N_19904);
nand UO_725 (O_725,N_19916,N_19848);
xor UO_726 (O_726,N_19614,N_19798);
nor UO_727 (O_727,N_19078,N_19382);
or UO_728 (O_728,N_19274,N_19276);
nor UO_729 (O_729,N_19951,N_19332);
or UO_730 (O_730,N_19730,N_19754);
nor UO_731 (O_731,N_19261,N_19296);
nand UO_732 (O_732,N_19211,N_19809);
and UO_733 (O_733,N_19181,N_19165);
nor UO_734 (O_734,N_19908,N_19269);
and UO_735 (O_735,N_19053,N_19818);
xnor UO_736 (O_736,N_19263,N_19787);
nand UO_737 (O_737,N_19270,N_19883);
nor UO_738 (O_738,N_19205,N_19353);
and UO_739 (O_739,N_19819,N_19488);
xnor UO_740 (O_740,N_19711,N_19587);
nand UO_741 (O_741,N_19340,N_19112);
or UO_742 (O_742,N_19195,N_19426);
nor UO_743 (O_743,N_19505,N_19992);
nand UO_744 (O_744,N_19689,N_19764);
nand UO_745 (O_745,N_19922,N_19051);
nand UO_746 (O_746,N_19008,N_19956);
xnor UO_747 (O_747,N_19944,N_19374);
nand UO_748 (O_748,N_19432,N_19193);
or UO_749 (O_749,N_19371,N_19278);
nor UO_750 (O_750,N_19761,N_19573);
nand UO_751 (O_751,N_19831,N_19809);
or UO_752 (O_752,N_19050,N_19009);
and UO_753 (O_753,N_19772,N_19960);
nand UO_754 (O_754,N_19621,N_19958);
or UO_755 (O_755,N_19716,N_19739);
xnor UO_756 (O_756,N_19779,N_19704);
or UO_757 (O_757,N_19455,N_19482);
or UO_758 (O_758,N_19649,N_19074);
nand UO_759 (O_759,N_19474,N_19478);
xor UO_760 (O_760,N_19811,N_19535);
or UO_761 (O_761,N_19317,N_19047);
nor UO_762 (O_762,N_19807,N_19792);
or UO_763 (O_763,N_19443,N_19718);
or UO_764 (O_764,N_19682,N_19903);
or UO_765 (O_765,N_19218,N_19871);
xor UO_766 (O_766,N_19320,N_19694);
xor UO_767 (O_767,N_19524,N_19652);
and UO_768 (O_768,N_19643,N_19422);
and UO_769 (O_769,N_19284,N_19315);
or UO_770 (O_770,N_19634,N_19519);
nor UO_771 (O_771,N_19085,N_19984);
nor UO_772 (O_772,N_19222,N_19413);
nand UO_773 (O_773,N_19280,N_19131);
and UO_774 (O_774,N_19872,N_19210);
and UO_775 (O_775,N_19767,N_19448);
xor UO_776 (O_776,N_19549,N_19819);
or UO_777 (O_777,N_19247,N_19793);
and UO_778 (O_778,N_19569,N_19564);
nand UO_779 (O_779,N_19542,N_19443);
and UO_780 (O_780,N_19056,N_19460);
and UO_781 (O_781,N_19429,N_19110);
and UO_782 (O_782,N_19674,N_19673);
or UO_783 (O_783,N_19640,N_19222);
xor UO_784 (O_784,N_19971,N_19530);
nand UO_785 (O_785,N_19452,N_19664);
nand UO_786 (O_786,N_19444,N_19573);
xnor UO_787 (O_787,N_19349,N_19148);
or UO_788 (O_788,N_19321,N_19930);
or UO_789 (O_789,N_19879,N_19927);
or UO_790 (O_790,N_19556,N_19990);
nor UO_791 (O_791,N_19073,N_19923);
or UO_792 (O_792,N_19756,N_19385);
nand UO_793 (O_793,N_19764,N_19815);
and UO_794 (O_794,N_19352,N_19053);
xor UO_795 (O_795,N_19957,N_19044);
xnor UO_796 (O_796,N_19913,N_19759);
and UO_797 (O_797,N_19774,N_19298);
nor UO_798 (O_798,N_19055,N_19221);
or UO_799 (O_799,N_19577,N_19140);
or UO_800 (O_800,N_19582,N_19906);
xnor UO_801 (O_801,N_19395,N_19861);
or UO_802 (O_802,N_19601,N_19862);
nor UO_803 (O_803,N_19721,N_19991);
or UO_804 (O_804,N_19603,N_19917);
xor UO_805 (O_805,N_19078,N_19557);
and UO_806 (O_806,N_19331,N_19491);
or UO_807 (O_807,N_19131,N_19297);
or UO_808 (O_808,N_19603,N_19862);
or UO_809 (O_809,N_19492,N_19869);
nand UO_810 (O_810,N_19202,N_19999);
nor UO_811 (O_811,N_19094,N_19396);
or UO_812 (O_812,N_19246,N_19277);
xnor UO_813 (O_813,N_19378,N_19359);
xor UO_814 (O_814,N_19019,N_19854);
nand UO_815 (O_815,N_19889,N_19682);
xor UO_816 (O_816,N_19958,N_19922);
nand UO_817 (O_817,N_19605,N_19221);
nor UO_818 (O_818,N_19698,N_19378);
and UO_819 (O_819,N_19267,N_19234);
or UO_820 (O_820,N_19301,N_19005);
nand UO_821 (O_821,N_19756,N_19616);
or UO_822 (O_822,N_19916,N_19279);
nand UO_823 (O_823,N_19572,N_19105);
nor UO_824 (O_824,N_19273,N_19457);
nand UO_825 (O_825,N_19018,N_19127);
nor UO_826 (O_826,N_19924,N_19420);
nand UO_827 (O_827,N_19437,N_19572);
nor UO_828 (O_828,N_19611,N_19939);
nand UO_829 (O_829,N_19015,N_19536);
xor UO_830 (O_830,N_19365,N_19137);
or UO_831 (O_831,N_19988,N_19470);
nor UO_832 (O_832,N_19752,N_19480);
nor UO_833 (O_833,N_19744,N_19900);
and UO_834 (O_834,N_19668,N_19945);
or UO_835 (O_835,N_19974,N_19854);
xnor UO_836 (O_836,N_19057,N_19848);
or UO_837 (O_837,N_19996,N_19078);
nor UO_838 (O_838,N_19832,N_19200);
xnor UO_839 (O_839,N_19668,N_19265);
xnor UO_840 (O_840,N_19456,N_19080);
nand UO_841 (O_841,N_19304,N_19372);
nor UO_842 (O_842,N_19007,N_19745);
nand UO_843 (O_843,N_19244,N_19060);
nor UO_844 (O_844,N_19997,N_19228);
xor UO_845 (O_845,N_19798,N_19227);
nor UO_846 (O_846,N_19994,N_19745);
and UO_847 (O_847,N_19035,N_19927);
and UO_848 (O_848,N_19754,N_19273);
or UO_849 (O_849,N_19445,N_19412);
nor UO_850 (O_850,N_19260,N_19665);
xor UO_851 (O_851,N_19255,N_19324);
nand UO_852 (O_852,N_19975,N_19347);
nand UO_853 (O_853,N_19028,N_19729);
or UO_854 (O_854,N_19830,N_19519);
nor UO_855 (O_855,N_19439,N_19557);
xnor UO_856 (O_856,N_19801,N_19569);
nand UO_857 (O_857,N_19744,N_19561);
and UO_858 (O_858,N_19353,N_19081);
nand UO_859 (O_859,N_19874,N_19387);
nor UO_860 (O_860,N_19910,N_19551);
nor UO_861 (O_861,N_19694,N_19850);
nand UO_862 (O_862,N_19141,N_19425);
and UO_863 (O_863,N_19374,N_19613);
nand UO_864 (O_864,N_19444,N_19112);
or UO_865 (O_865,N_19955,N_19538);
and UO_866 (O_866,N_19955,N_19256);
nand UO_867 (O_867,N_19493,N_19257);
xnor UO_868 (O_868,N_19938,N_19712);
nor UO_869 (O_869,N_19944,N_19109);
nor UO_870 (O_870,N_19010,N_19885);
xor UO_871 (O_871,N_19753,N_19574);
or UO_872 (O_872,N_19641,N_19628);
or UO_873 (O_873,N_19209,N_19264);
xnor UO_874 (O_874,N_19881,N_19274);
and UO_875 (O_875,N_19030,N_19202);
and UO_876 (O_876,N_19174,N_19735);
nor UO_877 (O_877,N_19451,N_19703);
or UO_878 (O_878,N_19950,N_19027);
or UO_879 (O_879,N_19983,N_19176);
and UO_880 (O_880,N_19986,N_19616);
and UO_881 (O_881,N_19474,N_19367);
or UO_882 (O_882,N_19857,N_19389);
xnor UO_883 (O_883,N_19496,N_19639);
xor UO_884 (O_884,N_19084,N_19011);
or UO_885 (O_885,N_19875,N_19483);
and UO_886 (O_886,N_19867,N_19714);
or UO_887 (O_887,N_19384,N_19725);
xnor UO_888 (O_888,N_19912,N_19777);
nor UO_889 (O_889,N_19508,N_19773);
xor UO_890 (O_890,N_19582,N_19174);
nand UO_891 (O_891,N_19938,N_19695);
nor UO_892 (O_892,N_19786,N_19678);
nand UO_893 (O_893,N_19518,N_19121);
or UO_894 (O_894,N_19170,N_19819);
nor UO_895 (O_895,N_19314,N_19025);
and UO_896 (O_896,N_19340,N_19425);
or UO_897 (O_897,N_19129,N_19314);
xnor UO_898 (O_898,N_19141,N_19937);
nor UO_899 (O_899,N_19158,N_19582);
and UO_900 (O_900,N_19143,N_19864);
nand UO_901 (O_901,N_19287,N_19520);
and UO_902 (O_902,N_19044,N_19151);
nand UO_903 (O_903,N_19041,N_19096);
nor UO_904 (O_904,N_19453,N_19300);
nand UO_905 (O_905,N_19320,N_19205);
nand UO_906 (O_906,N_19901,N_19284);
and UO_907 (O_907,N_19757,N_19637);
and UO_908 (O_908,N_19573,N_19008);
xor UO_909 (O_909,N_19019,N_19305);
or UO_910 (O_910,N_19819,N_19491);
or UO_911 (O_911,N_19267,N_19524);
nand UO_912 (O_912,N_19521,N_19254);
and UO_913 (O_913,N_19533,N_19546);
and UO_914 (O_914,N_19894,N_19688);
or UO_915 (O_915,N_19087,N_19682);
nand UO_916 (O_916,N_19845,N_19754);
or UO_917 (O_917,N_19573,N_19409);
xnor UO_918 (O_918,N_19262,N_19113);
nor UO_919 (O_919,N_19675,N_19280);
or UO_920 (O_920,N_19739,N_19298);
nand UO_921 (O_921,N_19684,N_19190);
xnor UO_922 (O_922,N_19277,N_19572);
nor UO_923 (O_923,N_19527,N_19694);
nand UO_924 (O_924,N_19301,N_19966);
nand UO_925 (O_925,N_19177,N_19484);
nand UO_926 (O_926,N_19554,N_19866);
or UO_927 (O_927,N_19797,N_19309);
xor UO_928 (O_928,N_19501,N_19439);
or UO_929 (O_929,N_19172,N_19040);
and UO_930 (O_930,N_19540,N_19403);
nand UO_931 (O_931,N_19124,N_19595);
nor UO_932 (O_932,N_19458,N_19355);
nor UO_933 (O_933,N_19101,N_19780);
and UO_934 (O_934,N_19014,N_19246);
nand UO_935 (O_935,N_19136,N_19821);
xor UO_936 (O_936,N_19021,N_19264);
or UO_937 (O_937,N_19337,N_19146);
nand UO_938 (O_938,N_19812,N_19434);
nand UO_939 (O_939,N_19611,N_19119);
and UO_940 (O_940,N_19769,N_19716);
and UO_941 (O_941,N_19422,N_19433);
xor UO_942 (O_942,N_19510,N_19598);
xnor UO_943 (O_943,N_19052,N_19119);
nand UO_944 (O_944,N_19793,N_19480);
xor UO_945 (O_945,N_19029,N_19672);
nand UO_946 (O_946,N_19863,N_19355);
and UO_947 (O_947,N_19941,N_19323);
or UO_948 (O_948,N_19911,N_19167);
nor UO_949 (O_949,N_19297,N_19053);
or UO_950 (O_950,N_19026,N_19201);
nor UO_951 (O_951,N_19205,N_19265);
nor UO_952 (O_952,N_19029,N_19678);
and UO_953 (O_953,N_19498,N_19922);
nand UO_954 (O_954,N_19608,N_19223);
and UO_955 (O_955,N_19555,N_19618);
or UO_956 (O_956,N_19481,N_19643);
xor UO_957 (O_957,N_19466,N_19461);
nor UO_958 (O_958,N_19060,N_19658);
and UO_959 (O_959,N_19205,N_19981);
xor UO_960 (O_960,N_19789,N_19411);
and UO_961 (O_961,N_19385,N_19447);
nor UO_962 (O_962,N_19967,N_19348);
and UO_963 (O_963,N_19957,N_19396);
nand UO_964 (O_964,N_19519,N_19343);
nor UO_965 (O_965,N_19971,N_19067);
xor UO_966 (O_966,N_19444,N_19366);
nor UO_967 (O_967,N_19598,N_19034);
or UO_968 (O_968,N_19021,N_19303);
xor UO_969 (O_969,N_19105,N_19720);
nand UO_970 (O_970,N_19010,N_19653);
nand UO_971 (O_971,N_19027,N_19313);
xor UO_972 (O_972,N_19600,N_19845);
nand UO_973 (O_973,N_19415,N_19629);
or UO_974 (O_974,N_19558,N_19963);
nand UO_975 (O_975,N_19077,N_19143);
or UO_976 (O_976,N_19819,N_19577);
and UO_977 (O_977,N_19476,N_19488);
and UO_978 (O_978,N_19822,N_19481);
or UO_979 (O_979,N_19935,N_19718);
and UO_980 (O_980,N_19063,N_19505);
and UO_981 (O_981,N_19063,N_19555);
nor UO_982 (O_982,N_19031,N_19170);
or UO_983 (O_983,N_19155,N_19869);
and UO_984 (O_984,N_19844,N_19662);
nor UO_985 (O_985,N_19570,N_19405);
nor UO_986 (O_986,N_19316,N_19100);
nor UO_987 (O_987,N_19246,N_19769);
xnor UO_988 (O_988,N_19671,N_19175);
xnor UO_989 (O_989,N_19951,N_19379);
nand UO_990 (O_990,N_19154,N_19627);
nand UO_991 (O_991,N_19182,N_19731);
and UO_992 (O_992,N_19795,N_19742);
and UO_993 (O_993,N_19957,N_19405);
nand UO_994 (O_994,N_19806,N_19544);
xnor UO_995 (O_995,N_19484,N_19494);
nand UO_996 (O_996,N_19830,N_19643);
nor UO_997 (O_997,N_19026,N_19487);
and UO_998 (O_998,N_19465,N_19058);
or UO_999 (O_999,N_19771,N_19730);
and UO_1000 (O_1000,N_19454,N_19841);
and UO_1001 (O_1001,N_19440,N_19827);
or UO_1002 (O_1002,N_19698,N_19971);
xnor UO_1003 (O_1003,N_19642,N_19059);
xor UO_1004 (O_1004,N_19556,N_19678);
or UO_1005 (O_1005,N_19338,N_19555);
or UO_1006 (O_1006,N_19526,N_19656);
and UO_1007 (O_1007,N_19448,N_19999);
xnor UO_1008 (O_1008,N_19146,N_19091);
nor UO_1009 (O_1009,N_19020,N_19405);
and UO_1010 (O_1010,N_19826,N_19853);
nor UO_1011 (O_1011,N_19083,N_19299);
and UO_1012 (O_1012,N_19924,N_19026);
and UO_1013 (O_1013,N_19723,N_19502);
and UO_1014 (O_1014,N_19135,N_19485);
xnor UO_1015 (O_1015,N_19789,N_19871);
and UO_1016 (O_1016,N_19824,N_19459);
or UO_1017 (O_1017,N_19851,N_19368);
xnor UO_1018 (O_1018,N_19654,N_19856);
nand UO_1019 (O_1019,N_19574,N_19803);
or UO_1020 (O_1020,N_19817,N_19603);
and UO_1021 (O_1021,N_19793,N_19253);
and UO_1022 (O_1022,N_19559,N_19443);
or UO_1023 (O_1023,N_19034,N_19576);
and UO_1024 (O_1024,N_19866,N_19440);
nor UO_1025 (O_1025,N_19029,N_19221);
and UO_1026 (O_1026,N_19333,N_19748);
or UO_1027 (O_1027,N_19392,N_19451);
nand UO_1028 (O_1028,N_19287,N_19068);
xor UO_1029 (O_1029,N_19642,N_19133);
nand UO_1030 (O_1030,N_19421,N_19402);
or UO_1031 (O_1031,N_19794,N_19924);
xnor UO_1032 (O_1032,N_19242,N_19769);
nor UO_1033 (O_1033,N_19275,N_19680);
and UO_1034 (O_1034,N_19629,N_19284);
xor UO_1035 (O_1035,N_19606,N_19627);
or UO_1036 (O_1036,N_19692,N_19136);
xnor UO_1037 (O_1037,N_19296,N_19816);
nand UO_1038 (O_1038,N_19239,N_19020);
nand UO_1039 (O_1039,N_19029,N_19480);
nand UO_1040 (O_1040,N_19440,N_19185);
nor UO_1041 (O_1041,N_19257,N_19352);
xnor UO_1042 (O_1042,N_19515,N_19993);
or UO_1043 (O_1043,N_19586,N_19000);
xnor UO_1044 (O_1044,N_19513,N_19658);
xnor UO_1045 (O_1045,N_19954,N_19586);
nor UO_1046 (O_1046,N_19950,N_19086);
and UO_1047 (O_1047,N_19135,N_19360);
nor UO_1048 (O_1048,N_19099,N_19703);
nor UO_1049 (O_1049,N_19615,N_19845);
or UO_1050 (O_1050,N_19696,N_19952);
xor UO_1051 (O_1051,N_19078,N_19533);
nor UO_1052 (O_1052,N_19367,N_19613);
nor UO_1053 (O_1053,N_19483,N_19184);
nand UO_1054 (O_1054,N_19513,N_19476);
or UO_1055 (O_1055,N_19503,N_19508);
xor UO_1056 (O_1056,N_19287,N_19800);
nor UO_1057 (O_1057,N_19314,N_19617);
nand UO_1058 (O_1058,N_19248,N_19908);
nand UO_1059 (O_1059,N_19027,N_19555);
and UO_1060 (O_1060,N_19050,N_19381);
xor UO_1061 (O_1061,N_19696,N_19494);
and UO_1062 (O_1062,N_19746,N_19597);
and UO_1063 (O_1063,N_19269,N_19439);
nor UO_1064 (O_1064,N_19848,N_19799);
and UO_1065 (O_1065,N_19500,N_19669);
and UO_1066 (O_1066,N_19515,N_19594);
nor UO_1067 (O_1067,N_19471,N_19515);
or UO_1068 (O_1068,N_19876,N_19295);
nor UO_1069 (O_1069,N_19688,N_19594);
xor UO_1070 (O_1070,N_19087,N_19864);
nor UO_1071 (O_1071,N_19488,N_19132);
or UO_1072 (O_1072,N_19794,N_19825);
nand UO_1073 (O_1073,N_19855,N_19962);
nand UO_1074 (O_1074,N_19117,N_19288);
and UO_1075 (O_1075,N_19884,N_19969);
xor UO_1076 (O_1076,N_19695,N_19414);
nor UO_1077 (O_1077,N_19149,N_19702);
nand UO_1078 (O_1078,N_19675,N_19897);
nand UO_1079 (O_1079,N_19057,N_19557);
nand UO_1080 (O_1080,N_19774,N_19882);
or UO_1081 (O_1081,N_19227,N_19483);
xor UO_1082 (O_1082,N_19636,N_19505);
nor UO_1083 (O_1083,N_19573,N_19207);
nand UO_1084 (O_1084,N_19465,N_19356);
nor UO_1085 (O_1085,N_19585,N_19632);
nand UO_1086 (O_1086,N_19612,N_19580);
or UO_1087 (O_1087,N_19509,N_19303);
or UO_1088 (O_1088,N_19553,N_19583);
xnor UO_1089 (O_1089,N_19813,N_19778);
xor UO_1090 (O_1090,N_19994,N_19859);
nor UO_1091 (O_1091,N_19299,N_19215);
nand UO_1092 (O_1092,N_19701,N_19338);
nand UO_1093 (O_1093,N_19720,N_19219);
nand UO_1094 (O_1094,N_19745,N_19675);
nor UO_1095 (O_1095,N_19006,N_19105);
and UO_1096 (O_1096,N_19569,N_19154);
or UO_1097 (O_1097,N_19067,N_19997);
or UO_1098 (O_1098,N_19108,N_19030);
or UO_1099 (O_1099,N_19753,N_19650);
nand UO_1100 (O_1100,N_19882,N_19200);
and UO_1101 (O_1101,N_19427,N_19242);
nor UO_1102 (O_1102,N_19790,N_19308);
nor UO_1103 (O_1103,N_19250,N_19760);
or UO_1104 (O_1104,N_19372,N_19992);
xnor UO_1105 (O_1105,N_19829,N_19046);
xor UO_1106 (O_1106,N_19831,N_19600);
nand UO_1107 (O_1107,N_19405,N_19106);
xnor UO_1108 (O_1108,N_19551,N_19178);
nor UO_1109 (O_1109,N_19185,N_19523);
or UO_1110 (O_1110,N_19692,N_19317);
nor UO_1111 (O_1111,N_19781,N_19419);
and UO_1112 (O_1112,N_19952,N_19678);
or UO_1113 (O_1113,N_19924,N_19171);
nor UO_1114 (O_1114,N_19552,N_19053);
nand UO_1115 (O_1115,N_19999,N_19793);
and UO_1116 (O_1116,N_19762,N_19348);
or UO_1117 (O_1117,N_19009,N_19222);
and UO_1118 (O_1118,N_19898,N_19409);
and UO_1119 (O_1119,N_19144,N_19793);
and UO_1120 (O_1120,N_19576,N_19988);
and UO_1121 (O_1121,N_19729,N_19550);
nand UO_1122 (O_1122,N_19879,N_19991);
nand UO_1123 (O_1123,N_19951,N_19981);
xnor UO_1124 (O_1124,N_19046,N_19420);
nand UO_1125 (O_1125,N_19432,N_19900);
nor UO_1126 (O_1126,N_19860,N_19398);
or UO_1127 (O_1127,N_19196,N_19719);
xor UO_1128 (O_1128,N_19311,N_19775);
xor UO_1129 (O_1129,N_19784,N_19823);
nand UO_1130 (O_1130,N_19513,N_19766);
nor UO_1131 (O_1131,N_19044,N_19355);
nand UO_1132 (O_1132,N_19389,N_19802);
nor UO_1133 (O_1133,N_19470,N_19445);
nor UO_1134 (O_1134,N_19326,N_19598);
nor UO_1135 (O_1135,N_19339,N_19979);
and UO_1136 (O_1136,N_19571,N_19388);
nand UO_1137 (O_1137,N_19824,N_19190);
or UO_1138 (O_1138,N_19150,N_19423);
or UO_1139 (O_1139,N_19626,N_19072);
xnor UO_1140 (O_1140,N_19591,N_19322);
nor UO_1141 (O_1141,N_19739,N_19358);
and UO_1142 (O_1142,N_19898,N_19907);
nand UO_1143 (O_1143,N_19808,N_19254);
xnor UO_1144 (O_1144,N_19539,N_19258);
and UO_1145 (O_1145,N_19171,N_19178);
and UO_1146 (O_1146,N_19047,N_19016);
nor UO_1147 (O_1147,N_19247,N_19471);
xnor UO_1148 (O_1148,N_19511,N_19529);
nor UO_1149 (O_1149,N_19339,N_19211);
or UO_1150 (O_1150,N_19115,N_19208);
or UO_1151 (O_1151,N_19557,N_19988);
or UO_1152 (O_1152,N_19594,N_19501);
nand UO_1153 (O_1153,N_19757,N_19267);
and UO_1154 (O_1154,N_19092,N_19916);
nand UO_1155 (O_1155,N_19657,N_19788);
xnor UO_1156 (O_1156,N_19045,N_19495);
or UO_1157 (O_1157,N_19835,N_19905);
and UO_1158 (O_1158,N_19856,N_19582);
xnor UO_1159 (O_1159,N_19544,N_19496);
or UO_1160 (O_1160,N_19279,N_19577);
and UO_1161 (O_1161,N_19027,N_19194);
xor UO_1162 (O_1162,N_19098,N_19019);
and UO_1163 (O_1163,N_19189,N_19298);
xor UO_1164 (O_1164,N_19416,N_19259);
and UO_1165 (O_1165,N_19359,N_19973);
or UO_1166 (O_1166,N_19008,N_19756);
nor UO_1167 (O_1167,N_19440,N_19256);
or UO_1168 (O_1168,N_19457,N_19555);
nor UO_1169 (O_1169,N_19940,N_19190);
nor UO_1170 (O_1170,N_19709,N_19400);
nand UO_1171 (O_1171,N_19228,N_19447);
and UO_1172 (O_1172,N_19387,N_19408);
and UO_1173 (O_1173,N_19827,N_19736);
xnor UO_1174 (O_1174,N_19612,N_19151);
and UO_1175 (O_1175,N_19445,N_19942);
nor UO_1176 (O_1176,N_19470,N_19736);
nor UO_1177 (O_1177,N_19012,N_19100);
nor UO_1178 (O_1178,N_19010,N_19180);
xor UO_1179 (O_1179,N_19255,N_19980);
nand UO_1180 (O_1180,N_19904,N_19011);
and UO_1181 (O_1181,N_19598,N_19747);
nor UO_1182 (O_1182,N_19162,N_19566);
or UO_1183 (O_1183,N_19342,N_19139);
xnor UO_1184 (O_1184,N_19110,N_19474);
and UO_1185 (O_1185,N_19982,N_19197);
and UO_1186 (O_1186,N_19094,N_19210);
nand UO_1187 (O_1187,N_19807,N_19725);
nand UO_1188 (O_1188,N_19952,N_19329);
or UO_1189 (O_1189,N_19955,N_19719);
nor UO_1190 (O_1190,N_19039,N_19064);
xor UO_1191 (O_1191,N_19857,N_19414);
nor UO_1192 (O_1192,N_19839,N_19024);
nor UO_1193 (O_1193,N_19531,N_19958);
and UO_1194 (O_1194,N_19322,N_19561);
or UO_1195 (O_1195,N_19755,N_19327);
and UO_1196 (O_1196,N_19987,N_19769);
and UO_1197 (O_1197,N_19036,N_19117);
nor UO_1198 (O_1198,N_19149,N_19224);
xnor UO_1199 (O_1199,N_19063,N_19029);
nor UO_1200 (O_1200,N_19699,N_19510);
xor UO_1201 (O_1201,N_19091,N_19463);
nor UO_1202 (O_1202,N_19659,N_19752);
nor UO_1203 (O_1203,N_19838,N_19640);
xor UO_1204 (O_1204,N_19257,N_19169);
and UO_1205 (O_1205,N_19134,N_19945);
or UO_1206 (O_1206,N_19583,N_19020);
xor UO_1207 (O_1207,N_19904,N_19602);
nand UO_1208 (O_1208,N_19904,N_19221);
and UO_1209 (O_1209,N_19425,N_19711);
nor UO_1210 (O_1210,N_19529,N_19920);
xnor UO_1211 (O_1211,N_19024,N_19446);
or UO_1212 (O_1212,N_19134,N_19220);
xor UO_1213 (O_1213,N_19972,N_19718);
nor UO_1214 (O_1214,N_19825,N_19357);
and UO_1215 (O_1215,N_19426,N_19978);
nand UO_1216 (O_1216,N_19151,N_19025);
nand UO_1217 (O_1217,N_19686,N_19629);
and UO_1218 (O_1218,N_19756,N_19709);
xnor UO_1219 (O_1219,N_19805,N_19801);
nor UO_1220 (O_1220,N_19473,N_19706);
nand UO_1221 (O_1221,N_19098,N_19344);
xnor UO_1222 (O_1222,N_19142,N_19199);
nor UO_1223 (O_1223,N_19871,N_19466);
or UO_1224 (O_1224,N_19607,N_19059);
xor UO_1225 (O_1225,N_19797,N_19180);
nor UO_1226 (O_1226,N_19924,N_19244);
nor UO_1227 (O_1227,N_19559,N_19951);
and UO_1228 (O_1228,N_19423,N_19347);
nor UO_1229 (O_1229,N_19720,N_19233);
and UO_1230 (O_1230,N_19741,N_19159);
xnor UO_1231 (O_1231,N_19186,N_19978);
and UO_1232 (O_1232,N_19709,N_19421);
or UO_1233 (O_1233,N_19081,N_19507);
xnor UO_1234 (O_1234,N_19834,N_19484);
nand UO_1235 (O_1235,N_19342,N_19482);
nand UO_1236 (O_1236,N_19544,N_19871);
nand UO_1237 (O_1237,N_19534,N_19439);
xor UO_1238 (O_1238,N_19814,N_19653);
and UO_1239 (O_1239,N_19756,N_19748);
nor UO_1240 (O_1240,N_19162,N_19291);
nor UO_1241 (O_1241,N_19100,N_19901);
nand UO_1242 (O_1242,N_19445,N_19807);
nor UO_1243 (O_1243,N_19072,N_19497);
nand UO_1244 (O_1244,N_19127,N_19973);
nor UO_1245 (O_1245,N_19711,N_19438);
nor UO_1246 (O_1246,N_19416,N_19581);
xor UO_1247 (O_1247,N_19634,N_19620);
or UO_1248 (O_1248,N_19599,N_19459);
or UO_1249 (O_1249,N_19032,N_19094);
nor UO_1250 (O_1250,N_19499,N_19158);
xor UO_1251 (O_1251,N_19336,N_19777);
xnor UO_1252 (O_1252,N_19810,N_19038);
xnor UO_1253 (O_1253,N_19718,N_19771);
and UO_1254 (O_1254,N_19462,N_19563);
nand UO_1255 (O_1255,N_19970,N_19236);
nand UO_1256 (O_1256,N_19231,N_19030);
nand UO_1257 (O_1257,N_19402,N_19014);
nor UO_1258 (O_1258,N_19307,N_19446);
or UO_1259 (O_1259,N_19387,N_19045);
nand UO_1260 (O_1260,N_19563,N_19484);
or UO_1261 (O_1261,N_19596,N_19898);
nor UO_1262 (O_1262,N_19318,N_19736);
nand UO_1263 (O_1263,N_19546,N_19573);
xor UO_1264 (O_1264,N_19795,N_19861);
and UO_1265 (O_1265,N_19049,N_19572);
nor UO_1266 (O_1266,N_19323,N_19108);
or UO_1267 (O_1267,N_19486,N_19695);
nand UO_1268 (O_1268,N_19690,N_19473);
or UO_1269 (O_1269,N_19897,N_19356);
nor UO_1270 (O_1270,N_19078,N_19748);
or UO_1271 (O_1271,N_19681,N_19248);
xnor UO_1272 (O_1272,N_19381,N_19254);
xnor UO_1273 (O_1273,N_19237,N_19063);
nand UO_1274 (O_1274,N_19351,N_19525);
nor UO_1275 (O_1275,N_19796,N_19037);
nor UO_1276 (O_1276,N_19905,N_19960);
nor UO_1277 (O_1277,N_19338,N_19068);
xor UO_1278 (O_1278,N_19847,N_19319);
xnor UO_1279 (O_1279,N_19370,N_19744);
nor UO_1280 (O_1280,N_19242,N_19044);
xnor UO_1281 (O_1281,N_19381,N_19630);
nand UO_1282 (O_1282,N_19778,N_19332);
and UO_1283 (O_1283,N_19748,N_19031);
nor UO_1284 (O_1284,N_19679,N_19342);
and UO_1285 (O_1285,N_19614,N_19759);
xnor UO_1286 (O_1286,N_19128,N_19955);
nand UO_1287 (O_1287,N_19483,N_19377);
or UO_1288 (O_1288,N_19838,N_19060);
or UO_1289 (O_1289,N_19533,N_19920);
nand UO_1290 (O_1290,N_19693,N_19319);
or UO_1291 (O_1291,N_19414,N_19307);
xnor UO_1292 (O_1292,N_19417,N_19073);
or UO_1293 (O_1293,N_19940,N_19977);
xnor UO_1294 (O_1294,N_19457,N_19104);
nand UO_1295 (O_1295,N_19451,N_19730);
nor UO_1296 (O_1296,N_19230,N_19428);
nand UO_1297 (O_1297,N_19765,N_19658);
xnor UO_1298 (O_1298,N_19943,N_19015);
nor UO_1299 (O_1299,N_19899,N_19863);
or UO_1300 (O_1300,N_19939,N_19380);
nor UO_1301 (O_1301,N_19750,N_19286);
nor UO_1302 (O_1302,N_19855,N_19544);
nand UO_1303 (O_1303,N_19313,N_19883);
nand UO_1304 (O_1304,N_19370,N_19265);
xor UO_1305 (O_1305,N_19590,N_19259);
nand UO_1306 (O_1306,N_19592,N_19497);
nor UO_1307 (O_1307,N_19092,N_19710);
and UO_1308 (O_1308,N_19477,N_19809);
nor UO_1309 (O_1309,N_19676,N_19965);
or UO_1310 (O_1310,N_19279,N_19951);
and UO_1311 (O_1311,N_19235,N_19641);
nor UO_1312 (O_1312,N_19793,N_19191);
xor UO_1313 (O_1313,N_19839,N_19729);
xnor UO_1314 (O_1314,N_19315,N_19063);
and UO_1315 (O_1315,N_19812,N_19540);
xnor UO_1316 (O_1316,N_19729,N_19353);
nand UO_1317 (O_1317,N_19267,N_19967);
nand UO_1318 (O_1318,N_19581,N_19030);
or UO_1319 (O_1319,N_19741,N_19410);
or UO_1320 (O_1320,N_19274,N_19729);
nand UO_1321 (O_1321,N_19384,N_19890);
or UO_1322 (O_1322,N_19835,N_19701);
or UO_1323 (O_1323,N_19090,N_19265);
xnor UO_1324 (O_1324,N_19477,N_19191);
nor UO_1325 (O_1325,N_19473,N_19917);
or UO_1326 (O_1326,N_19150,N_19172);
or UO_1327 (O_1327,N_19616,N_19207);
nand UO_1328 (O_1328,N_19415,N_19708);
nand UO_1329 (O_1329,N_19881,N_19606);
xor UO_1330 (O_1330,N_19268,N_19037);
xor UO_1331 (O_1331,N_19249,N_19359);
and UO_1332 (O_1332,N_19135,N_19463);
xor UO_1333 (O_1333,N_19148,N_19015);
nand UO_1334 (O_1334,N_19073,N_19717);
and UO_1335 (O_1335,N_19194,N_19314);
or UO_1336 (O_1336,N_19831,N_19160);
and UO_1337 (O_1337,N_19653,N_19911);
nor UO_1338 (O_1338,N_19279,N_19991);
or UO_1339 (O_1339,N_19460,N_19621);
nand UO_1340 (O_1340,N_19098,N_19105);
nand UO_1341 (O_1341,N_19663,N_19706);
or UO_1342 (O_1342,N_19796,N_19352);
xnor UO_1343 (O_1343,N_19892,N_19070);
and UO_1344 (O_1344,N_19599,N_19151);
or UO_1345 (O_1345,N_19263,N_19039);
nand UO_1346 (O_1346,N_19855,N_19814);
or UO_1347 (O_1347,N_19421,N_19785);
xnor UO_1348 (O_1348,N_19075,N_19364);
xor UO_1349 (O_1349,N_19999,N_19491);
or UO_1350 (O_1350,N_19319,N_19950);
nor UO_1351 (O_1351,N_19349,N_19451);
and UO_1352 (O_1352,N_19565,N_19065);
xnor UO_1353 (O_1353,N_19789,N_19451);
xor UO_1354 (O_1354,N_19352,N_19657);
nor UO_1355 (O_1355,N_19422,N_19658);
nor UO_1356 (O_1356,N_19657,N_19366);
nor UO_1357 (O_1357,N_19775,N_19700);
and UO_1358 (O_1358,N_19280,N_19476);
and UO_1359 (O_1359,N_19234,N_19875);
nand UO_1360 (O_1360,N_19705,N_19322);
xor UO_1361 (O_1361,N_19077,N_19328);
nor UO_1362 (O_1362,N_19659,N_19908);
nand UO_1363 (O_1363,N_19023,N_19567);
and UO_1364 (O_1364,N_19831,N_19824);
xnor UO_1365 (O_1365,N_19691,N_19160);
and UO_1366 (O_1366,N_19052,N_19802);
nor UO_1367 (O_1367,N_19376,N_19060);
or UO_1368 (O_1368,N_19032,N_19249);
nand UO_1369 (O_1369,N_19528,N_19130);
xnor UO_1370 (O_1370,N_19004,N_19913);
and UO_1371 (O_1371,N_19287,N_19297);
nor UO_1372 (O_1372,N_19524,N_19206);
and UO_1373 (O_1373,N_19550,N_19765);
or UO_1374 (O_1374,N_19292,N_19456);
xor UO_1375 (O_1375,N_19148,N_19341);
or UO_1376 (O_1376,N_19818,N_19151);
nor UO_1377 (O_1377,N_19380,N_19128);
and UO_1378 (O_1378,N_19204,N_19880);
xor UO_1379 (O_1379,N_19513,N_19136);
or UO_1380 (O_1380,N_19596,N_19502);
nand UO_1381 (O_1381,N_19840,N_19852);
and UO_1382 (O_1382,N_19076,N_19611);
and UO_1383 (O_1383,N_19433,N_19136);
nand UO_1384 (O_1384,N_19436,N_19654);
or UO_1385 (O_1385,N_19143,N_19505);
nand UO_1386 (O_1386,N_19552,N_19195);
nand UO_1387 (O_1387,N_19991,N_19913);
xnor UO_1388 (O_1388,N_19665,N_19146);
and UO_1389 (O_1389,N_19398,N_19403);
xnor UO_1390 (O_1390,N_19650,N_19959);
and UO_1391 (O_1391,N_19016,N_19426);
xnor UO_1392 (O_1392,N_19229,N_19885);
nor UO_1393 (O_1393,N_19900,N_19741);
and UO_1394 (O_1394,N_19130,N_19406);
nand UO_1395 (O_1395,N_19973,N_19697);
nand UO_1396 (O_1396,N_19502,N_19746);
or UO_1397 (O_1397,N_19664,N_19012);
xnor UO_1398 (O_1398,N_19639,N_19943);
nor UO_1399 (O_1399,N_19676,N_19053);
xor UO_1400 (O_1400,N_19197,N_19915);
and UO_1401 (O_1401,N_19923,N_19077);
nand UO_1402 (O_1402,N_19355,N_19734);
xor UO_1403 (O_1403,N_19708,N_19265);
and UO_1404 (O_1404,N_19110,N_19482);
nor UO_1405 (O_1405,N_19546,N_19348);
nor UO_1406 (O_1406,N_19352,N_19542);
or UO_1407 (O_1407,N_19381,N_19428);
nand UO_1408 (O_1408,N_19623,N_19980);
nor UO_1409 (O_1409,N_19754,N_19621);
xor UO_1410 (O_1410,N_19652,N_19074);
and UO_1411 (O_1411,N_19973,N_19799);
nand UO_1412 (O_1412,N_19195,N_19771);
xnor UO_1413 (O_1413,N_19706,N_19118);
and UO_1414 (O_1414,N_19468,N_19217);
and UO_1415 (O_1415,N_19387,N_19063);
xnor UO_1416 (O_1416,N_19481,N_19083);
xor UO_1417 (O_1417,N_19709,N_19845);
or UO_1418 (O_1418,N_19376,N_19401);
nand UO_1419 (O_1419,N_19327,N_19282);
or UO_1420 (O_1420,N_19534,N_19236);
nor UO_1421 (O_1421,N_19910,N_19926);
nor UO_1422 (O_1422,N_19975,N_19714);
or UO_1423 (O_1423,N_19843,N_19838);
nand UO_1424 (O_1424,N_19558,N_19029);
and UO_1425 (O_1425,N_19872,N_19056);
nor UO_1426 (O_1426,N_19618,N_19814);
and UO_1427 (O_1427,N_19970,N_19230);
nand UO_1428 (O_1428,N_19035,N_19926);
and UO_1429 (O_1429,N_19420,N_19068);
nand UO_1430 (O_1430,N_19172,N_19637);
and UO_1431 (O_1431,N_19165,N_19423);
nand UO_1432 (O_1432,N_19132,N_19289);
xnor UO_1433 (O_1433,N_19622,N_19065);
nand UO_1434 (O_1434,N_19336,N_19305);
nand UO_1435 (O_1435,N_19032,N_19316);
and UO_1436 (O_1436,N_19411,N_19611);
nor UO_1437 (O_1437,N_19229,N_19830);
xnor UO_1438 (O_1438,N_19091,N_19207);
xnor UO_1439 (O_1439,N_19387,N_19133);
or UO_1440 (O_1440,N_19855,N_19816);
xor UO_1441 (O_1441,N_19921,N_19953);
nand UO_1442 (O_1442,N_19930,N_19995);
nand UO_1443 (O_1443,N_19240,N_19564);
nor UO_1444 (O_1444,N_19256,N_19289);
or UO_1445 (O_1445,N_19349,N_19324);
and UO_1446 (O_1446,N_19944,N_19010);
nor UO_1447 (O_1447,N_19083,N_19046);
xnor UO_1448 (O_1448,N_19266,N_19407);
or UO_1449 (O_1449,N_19311,N_19353);
or UO_1450 (O_1450,N_19756,N_19172);
nand UO_1451 (O_1451,N_19605,N_19193);
xnor UO_1452 (O_1452,N_19542,N_19142);
xnor UO_1453 (O_1453,N_19292,N_19749);
or UO_1454 (O_1454,N_19106,N_19389);
nand UO_1455 (O_1455,N_19234,N_19898);
nand UO_1456 (O_1456,N_19931,N_19005);
nand UO_1457 (O_1457,N_19932,N_19383);
and UO_1458 (O_1458,N_19753,N_19694);
nand UO_1459 (O_1459,N_19752,N_19130);
or UO_1460 (O_1460,N_19114,N_19169);
xor UO_1461 (O_1461,N_19518,N_19315);
xnor UO_1462 (O_1462,N_19503,N_19149);
nand UO_1463 (O_1463,N_19219,N_19784);
or UO_1464 (O_1464,N_19337,N_19682);
nor UO_1465 (O_1465,N_19860,N_19512);
nand UO_1466 (O_1466,N_19491,N_19653);
and UO_1467 (O_1467,N_19952,N_19883);
nor UO_1468 (O_1468,N_19783,N_19437);
nand UO_1469 (O_1469,N_19983,N_19597);
and UO_1470 (O_1470,N_19143,N_19123);
or UO_1471 (O_1471,N_19491,N_19767);
nand UO_1472 (O_1472,N_19649,N_19117);
nor UO_1473 (O_1473,N_19612,N_19720);
or UO_1474 (O_1474,N_19410,N_19251);
xor UO_1475 (O_1475,N_19108,N_19009);
nand UO_1476 (O_1476,N_19974,N_19679);
or UO_1477 (O_1477,N_19700,N_19938);
or UO_1478 (O_1478,N_19506,N_19599);
xor UO_1479 (O_1479,N_19667,N_19586);
xor UO_1480 (O_1480,N_19060,N_19072);
nor UO_1481 (O_1481,N_19500,N_19954);
nor UO_1482 (O_1482,N_19131,N_19344);
and UO_1483 (O_1483,N_19547,N_19292);
or UO_1484 (O_1484,N_19472,N_19768);
nor UO_1485 (O_1485,N_19961,N_19646);
xnor UO_1486 (O_1486,N_19240,N_19430);
nand UO_1487 (O_1487,N_19884,N_19208);
nor UO_1488 (O_1488,N_19505,N_19797);
xor UO_1489 (O_1489,N_19568,N_19945);
xor UO_1490 (O_1490,N_19895,N_19222);
or UO_1491 (O_1491,N_19429,N_19065);
xnor UO_1492 (O_1492,N_19085,N_19918);
and UO_1493 (O_1493,N_19946,N_19409);
and UO_1494 (O_1494,N_19162,N_19356);
and UO_1495 (O_1495,N_19642,N_19968);
or UO_1496 (O_1496,N_19544,N_19952);
and UO_1497 (O_1497,N_19274,N_19135);
or UO_1498 (O_1498,N_19951,N_19497);
and UO_1499 (O_1499,N_19068,N_19508);
and UO_1500 (O_1500,N_19953,N_19037);
or UO_1501 (O_1501,N_19005,N_19388);
and UO_1502 (O_1502,N_19920,N_19394);
nand UO_1503 (O_1503,N_19574,N_19806);
nor UO_1504 (O_1504,N_19753,N_19525);
and UO_1505 (O_1505,N_19999,N_19528);
and UO_1506 (O_1506,N_19618,N_19586);
nand UO_1507 (O_1507,N_19719,N_19918);
and UO_1508 (O_1508,N_19694,N_19631);
xnor UO_1509 (O_1509,N_19738,N_19542);
nand UO_1510 (O_1510,N_19250,N_19621);
or UO_1511 (O_1511,N_19247,N_19461);
or UO_1512 (O_1512,N_19602,N_19464);
and UO_1513 (O_1513,N_19834,N_19062);
and UO_1514 (O_1514,N_19052,N_19976);
and UO_1515 (O_1515,N_19445,N_19098);
and UO_1516 (O_1516,N_19798,N_19351);
and UO_1517 (O_1517,N_19841,N_19910);
nand UO_1518 (O_1518,N_19295,N_19105);
nand UO_1519 (O_1519,N_19385,N_19987);
or UO_1520 (O_1520,N_19486,N_19113);
or UO_1521 (O_1521,N_19624,N_19252);
and UO_1522 (O_1522,N_19400,N_19222);
xnor UO_1523 (O_1523,N_19904,N_19382);
or UO_1524 (O_1524,N_19551,N_19408);
and UO_1525 (O_1525,N_19713,N_19800);
or UO_1526 (O_1526,N_19414,N_19802);
and UO_1527 (O_1527,N_19854,N_19543);
nand UO_1528 (O_1528,N_19001,N_19230);
nor UO_1529 (O_1529,N_19786,N_19589);
nor UO_1530 (O_1530,N_19572,N_19180);
nand UO_1531 (O_1531,N_19040,N_19193);
and UO_1532 (O_1532,N_19542,N_19943);
or UO_1533 (O_1533,N_19755,N_19274);
and UO_1534 (O_1534,N_19260,N_19508);
xor UO_1535 (O_1535,N_19944,N_19397);
nand UO_1536 (O_1536,N_19595,N_19356);
nor UO_1537 (O_1537,N_19563,N_19687);
nand UO_1538 (O_1538,N_19923,N_19340);
or UO_1539 (O_1539,N_19036,N_19423);
xor UO_1540 (O_1540,N_19633,N_19224);
nand UO_1541 (O_1541,N_19494,N_19300);
nand UO_1542 (O_1542,N_19901,N_19050);
or UO_1543 (O_1543,N_19196,N_19961);
nor UO_1544 (O_1544,N_19406,N_19587);
nand UO_1545 (O_1545,N_19500,N_19841);
nand UO_1546 (O_1546,N_19658,N_19832);
or UO_1547 (O_1547,N_19957,N_19535);
nor UO_1548 (O_1548,N_19631,N_19593);
or UO_1549 (O_1549,N_19577,N_19748);
nand UO_1550 (O_1550,N_19641,N_19371);
xnor UO_1551 (O_1551,N_19996,N_19433);
xnor UO_1552 (O_1552,N_19680,N_19236);
nor UO_1553 (O_1553,N_19999,N_19398);
nor UO_1554 (O_1554,N_19443,N_19498);
nand UO_1555 (O_1555,N_19331,N_19928);
and UO_1556 (O_1556,N_19580,N_19810);
nand UO_1557 (O_1557,N_19059,N_19690);
or UO_1558 (O_1558,N_19976,N_19434);
nand UO_1559 (O_1559,N_19729,N_19974);
nor UO_1560 (O_1560,N_19816,N_19196);
nand UO_1561 (O_1561,N_19435,N_19761);
nor UO_1562 (O_1562,N_19834,N_19295);
xor UO_1563 (O_1563,N_19332,N_19749);
and UO_1564 (O_1564,N_19138,N_19110);
xnor UO_1565 (O_1565,N_19608,N_19753);
nor UO_1566 (O_1566,N_19967,N_19042);
nor UO_1567 (O_1567,N_19697,N_19234);
or UO_1568 (O_1568,N_19568,N_19116);
or UO_1569 (O_1569,N_19730,N_19827);
or UO_1570 (O_1570,N_19882,N_19811);
nor UO_1571 (O_1571,N_19269,N_19796);
nand UO_1572 (O_1572,N_19166,N_19535);
or UO_1573 (O_1573,N_19682,N_19602);
or UO_1574 (O_1574,N_19158,N_19707);
nor UO_1575 (O_1575,N_19704,N_19048);
nand UO_1576 (O_1576,N_19109,N_19433);
nor UO_1577 (O_1577,N_19765,N_19006);
nor UO_1578 (O_1578,N_19772,N_19444);
and UO_1579 (O_1579,N_19334,N_19561);
and UO_1580 (O_1580,N_19766,N_19312);
nor UO_1581 (O_1581,N_19980,N_19896);
nor UO_1582 (O_1582,N_19288,N_19750);
and UO_1583 (O_1583,N_19574,N_19270);
nand UO_1584 (O_1584,N_19685,N_19941);
nand UO_1585 (O_1585,N_19787,N_19858);
nand UO_1586 (O_1586,N_19220,N_19358);
and UO_1587 (O_1587,N_19993,N_19429);
and UO_1588 (O_1588,N_19909,N_19662);
nand UO_1589 (O_1589,N_19574,N_19601);
or UO_1590 (O_1590,N_19570,N_19470);
and UO_1591 (O_1591,N_19602,N_19032);
nand UO_1592 (O_1592,N_19694,N_19750);
xor UO_1593 (O_1593,N_19397,N_19765);
or UO_1594 (O_1594,N_19995,N_19318);
nor UO_1595 (O_1595,N_19440,N_19724);
nand UO_1596 (O_1596,N_19731,N_19793);
nand UO_1597 (O_1597,N_19443,N_19212);
and UO_1598 (O_1598,N_19534,N_19050);
nor UO_1599 (O_1599,N_19065,N_19475);
and UO_1600 (O_1600,N_19132,N_19277);
and UO_1601 (O_1601,N_19960,N_19117);
nor UO_1602 (O_1602,N_19491,N_19076);
or UO_1603 (O_1603,N_19107,N_19159);
nand UO_1604 (O_1604,N_19072,N_19676);
and UO_1605 (O_1605,N_19192,N_19605);
xnor UO_1606 (O_1606,N_19619,N_19555);
and UO_1607 (O_1607,N_19162,N_19965);
nor UO_1608 (O_1608,N_19632,N_19420);
nand UO_1609 (O_1609,N_19437,N_19920);
or UO_1610 (O_1610,N_19706,N_19120);
xor UO_1611 (O_1611,N_19514,N_19797);
nor UO_1612 (O_1612,N_19946,N_19210);
xnor UO_1613 (O_1613,N_19653,N_19329);
or UO_1614 (O_1614,N_19734,N_19244);
nor UO_1615 (O_1615,N_19122,N_19391);
and UO_1616 (O_1616,N_19233,N_19990);
or UO_1617 (O_1617,N_19502,N_19019);
or UO_1618 (O_1618,N_19021,N_19102);
xnor UO_1619 (O_1619,N_19308,N_19530);
or UO_1620 (O_1620,N_19128,N_19378);
nor UO_1621 (O_1621,N_19010,N_19947);
xnor UO_1622 (O_1622,N_19702,N_19015);
nor UO_1623 (O_1623,N_19231,N_19307);
xor UO_1624 (O_1624,N_19719,N_19730);
or UO_1625 (O_1625,N_19558,N_19957);
nand UO_1626 (O_1626,N_19186,N_19496);
or UO_1627 (O_1627,N_19377,N_19287);
xor UO_1628 (O_1628,N_19455,N_19691);
xnor UO_1629 (O_1629,N_19409,N_19959);
xor UO_1630 (O_1630,N_19394,N_19241);
and UO_1631 (O_1631,N_19613,N_19928);
nand UO_1632 (O_1632,N_19154,N_19806);
or UO_1633 (O_1633,N_19792,N_19404);
or UO_1634 (O_1634,N_19900,N_19140);
or UO_1635 (O_1635,N_19823,N_19884);
nand UO_1636 (O_1636,N_19137,N_19421);
or UO_1637 (O_1637,N_19472,N_19098);
nor UO_1638 (O_1638,N_19052,N_19602);
nor UO_1639 (O_1639,N_19983,N_19169);
nand UO_1640 (O_1640,N_19283,N_19932);
nand UO_1641 (O_1641,N_19113,N_19036);
nand UO_1642 (O_1642,N_19410,N_19524);
and UO_1643 (O_1643,N_19638,N_19647);
and UO_1644 (O_1644,N_19603,N_19938);
xor UO_1645 (O_1645,N_19784,N_19172);
xor UO_1646 (O_1646,N_19853,N_19608);
and UO_1647 (O_1647,N_19416,N_19795);
nor UO_1648 (O_1648,N_19663,N_19955);
and UO_1649 (O_1649,N_19651,N_19712);
nand UO_1650 (O_1650,N_19069,N_19168);
nor UO_1651 (O_1651,N_19184,N_19191);
nand UO_1652 (O_1652,N_19819,N_19245);
or UO_1653 (O_1653,N_19509,N_19156);
xor UO_1654 (O_1654,N_19381,N_19826);
or UO_1655 (O_1655,N_19219,N_19110);
xor UO_1656 (O_1656,N_19385,N_19435);
nor UO_1657 (O_1657,N_19279,N_19071);
and UO_1658 (O_1658,N_19425,N_19793);
nor UO_1659 (O_1659,N_19723,N_19674);
or UO_1660 (O_1660,N_19533,N_19179);
or UO_1661 (O_1661,N_19597,N_19239);
nor UO_1662 (O_1662,N_19961,N_19936);
xnor UO_1663 (O_1663,N_19378,N_19730);
nor UO_1664 (O_1664,N_19136,N_19103);
xnor UO_1665 (O_1665,N_19629,N_19148);
nand UO_1666 (O_1666,N_19552,N_19859);
or UO_1667 (O_1667,N_19003,N_19910);
nand UO_1668 (O_1668,N_19972,N_19580);
xor UO_1669 (O_1669,N_19564,N_19284);
nand UO_1670 (O_1670,N_19928,N_19939);
nand UO_1671 (O_1671,N_19453,N_19021);
and UO_1672 (O_1672,N_19821,N_19958);
xor UO_1673 (O_1673,N_19147,N_19046);
and UO_1674 (O_1674,N_19807,N_19772);
nor UO_1675 (O_1675,N_19992,N_19652);
nor UO_1676 (O_1676,N_19898,N_19150);
and UO_1677 (O_1677,N_19477,N_19879);
or UO_1678 (O_1678,N_19987,N_19230);
and UO_1679 (O_1679,N_19673,N_19133);
nor UO_1680 (O_1680,N_19572,N_19094);
nand UO_1681 (O_1681,N_19053,N_19141);
xnor UO_1682 (O_1682,N_19561,N_19195);
xor UO_1683 (O_1683,N_19456,N_19273);
and UO_1684 (O_1684,N_19373,N_19952);
nor UO_1685 (O_1685,N_19425,N_19262);
nor UO_1686 (O_1686,N_19621,N_19313);
xor UO_1687 (O_1687,N_19562,N_19521);
and UO_1688 (O_1688,N_19963,N_19402);
xor UO_1689 (O_1689,N_19018,N_19385);
nor UO_1690 (O_1690,N_19194,N_19581);
or UO_1691 (O_1691,N_19895,N_19087);
and UO_1692 (O_1692,N_19476,N_19958);
nor UO_1693 (O_1693,N_19307,N_19111);
or UO_1694 (O_1694,N_19091,N_19546);
or UO_1695 (O_1695,N_19049,N_19329);
nand UO_1696 (O_1696,N_19360,N_19580);
or UO_1697 (O_1697,N_19415,N_19454);
or UO_1698 (O_1698,N_19234,N_19390);
xor UO_1699 (O_1699,N_19832,N_19665);
or UO_1700 (O_1700,N_19617,N_19960);
nor UO_1701 (O_1701,N_19223,N_19711);
nand UO_1702 (O_1702,N_19569,N_19125);
xnor UO_1703 (O_1703,N_19742,N_19989);
xor UO_1704 (O_1704,N_19433,N_19844);
nand UO_1705 (O_1705,N_19484,N_19124);
nor UO_1706 (O_1706,N_19914,N_19598);
or UO_1707 (O_1707,N_19599,N_19311);
nor UO_1708 (O_1708,N_19463,N_19885);
nand UO_1709 (O_1709,N_19221,N_19619);
or UO_1710 (O_1710,N_19465,N_19704);
nor UO_1711 (O_1711,N_19758,N_19138);
xor UO_1712 (O_1712,N_19455,N_19733);
nor UO_1713 (O_1713,N_19962,N_19159);
nand UO_1714 (O_1714,N_19033,N_19507);
xor UO_1715 (O_1715,N_19119,N_19380);
nand UO_1716 (O_1716,N_19441,N_19821);
or UO_1717 (O_1717,N_19374,N_19406);
or UO_1718 (O_1718,N_19773,N_19488);
and UO_1719 (O_1719,N_19659,N_19745);
nand UO_1720 (O_1720,N_19300,N_19710);
nand UO_1721 (O_1721,N_19815,N_19783);
nor UO_1722 (O_1722,N_19679,N_19541);
xor UO_1723 (O_1723,N_19253,N_19946);
nor UO_1724 (O_1724,N_19408,N_19341);
or UO_1725 (O_1725,N_19088,N_19706);
nor UO_1726 (O_1726,N_19360,N_19311);
and UO_1727 (O_1727,N_19484,N_19182);
nand UO_1728 (O_1728,N_19153,N_19906);
or UO_1729 (O_1729,N_19731,N_19158);
xor UO_1730 (O_1730,N_19925,N_19737);
and UO_1731 (O_1731,N_19527,N_19252);
xor UO_1732 (O_1732,N_19819,N_19809);
nand UO_1733 (O_1733,N_19203,N_19196);
or UO_1734 (O_1734,N_19382,N_19906);
xor UO_1735 (O_1735,N_19225,N_19512);
nor UO_1736 (O_1736,N_19082,N_19831);
or UO_1737 (O_1737,N_19751,N_19787);
or UO_1738 (O_1738,N_19981,N_19949);
or UO_1739 (O_1739,N_19189,N_19957);
nor UO_1740 (O_1740,N_19397,N_19031);
or UO_1741 (O_1741,N_19242,N_19257);
xor UO_1742 (O_1742,N_19027,N_19587);
xnor UO_1743 (O_1743,N_19737,N_19483);
nor UO_1744 (O_1744,N_19199,N_19144);
or UO_1745 (O_1745,N_19028,N_19976);
nand UO_1746 (O_1746,N_19136,N_19224);
and UO_1747 (O_1747,N_19279,N_19861);
nor UO_1748 (O_1748,N_19070,N_19140);
or UO_1749 (O_1749,N_19490,N_19885);
and UO_1750 (O_1750,N_19566,N_19398);
xnor UO_1751 (O_1751,N_19789,N_19936);
xnor UO_1752 (O_1752,N_19188,N_19647);
and UO_1753 (O_1753,N_19040,N_19692);
nand UO_1754 (O_1754,N_19047,N_19409);
and UO_1755 (O_1755,N_19880,N_19943);
nand UO_1756 (O_1756,N_19988,N_19962);
nor UO_1757 (O_1757,N_19311,N_19209);
or UO_1758 (O_1758,N_19487,N_19519);
nor UO_1759 (O_1759,N_19445,N_19211);
nor UO_1760 (O_1760,N_19609,N_19566);
nand UO_1761 (O_1761,N_19618,N_19808);
nor UO_1762 (O_1762,N_19770,N_19527);
xor UO_1763 (O_1763,N_19913,N_19342);
nor UO_1764 (O_1764,N_19963,N_19900);
or UO_1765 (O_1765,N_19035,N_19633);
or UO_1766 (O_1766,N_19725,N_19948);
and UO_1767 (O_1767,N_19289,N_19859);
xnor UO_1768 (O_1768,N_19525,N_19302);
or UO_1769 (O_1769,N_19561,N_19070);
and UO_1770 (O_1770,N_19591,N_19211);
xor UO_1771 (O_1771,N_19623,N_19787);
nor UO_1772 (O_1772,N_19774,N_19978);
or UO_1773 (O_1773,N_19484,N_19345);
and UO_1774 (O_1774,N_19081,N_19232);
or UO_1775 (O_1775,N_19053,N_19941);
nor UO_1776 (O_1776,N_19814,N_19929);
nor UO_1777 (O_1777,N_19494,N_19420);
and UO_1778 (O_1778,N_19759,N_19301);
xnor UO_1779 (O_1779,N_19790,N_19381);
nor UO_1780 (O_1780,N_19722,N_19038);
nand UO_1781 (O_1781,N_19114,N_19739);
or UO_1782 (O_1782,N_19810,N_19885);
xor UO_1783 (O_1783,N_19329,N_19510);
nor UO_1784 (O_1784,N_19411,N_19485);
xor UO_1785 (O_1785,N_19955,N_19551);
or UO_1786 (O_1786,N_19766,N_19505);
nor UO_1787 (O_1787,N_19039,N_19769);
or UO_1788 (O_1788,N_19257,N_19516);
nand UO_1789 (O_1789,N_19829,N_19495);
or UO_1790 (O_1790,N_19978,N_19387);
nand UO_1791 (O_1791,N_19426,N_19276);
nor UO_1792 (O_1792,N_19566,N_19222);
nand UO_1793 (O_1793,N_19817,N_19703);
and UO_1794 (O_1794,N_19004,N_19411);
xor UO_1795 (O_1795,N_19411,N_19757);
and UO_1796 (O_1796,N_19057,N_19697);
and UO_1797 (O_1797,N_19896,N_19347);
and UO_1798 (O_1798,N_19049,N_19668);
nand UO_1799 (O_1799,N_19931,N_19802);
and UO_1800 (O_1800,N_19151,N_19380);
xor UO_1801 (O_1801,N_19907,N_19620);
and UO_1802 (O_1802,N_19862,N_19010);
nor UO_1803 (O_1803,N_19556,N_19770);
and UO_1804 (O_1804,N_19244,N_19698);
or UO_1805 (O_1805,N_19373,N_19216);
or UO_1806 (O_1806,N_19937,N_19961);
and UO_1807 (O_1807,N_19130,N_19546);
and UO_1808 (O_1808,N_19095,N_19098);
nor UO_1809 (O_1809,N_19674,N_19087);
xnor UO_1810 (O_1810,N_19727,N_19674);
xnor UO_1811 (O_1811,N_19024,N_19066);
or UO_1812 (O_1812,N_19270,N_19091);
or UO_1813 (O_1813,N_19784,N_19340);
xor UO_1814 (O_1814,N_19308,N_19316);
and UO_1815 (O_1815,N_19090,N_19343);
and UO_1816 (O_1816,N_19667,N_19848);
xor UO_1817 (O_1817,N_19457,N_19012);
and UO_1818 (O_1818,N_19657,N_19495);
xor UO_1819 (O_1819,N_19449,N_19309);
or UO_1820 (O_1820,N_19185,N_19325);
nand UO_1821 (O_1821,N_19068,N_19779);
or UO_1822 (O_1822,N_19074,N_19218);
nor UO_1823 (O_1823,N_19749,N_19628);
or UO_1824 (O_1824,N_19192,N_19780);
nor UO_1825 (O_1825,N_19941,N_19841);
and UO_1826 (O_1826,N_19872,N_19578);
and UO_1827 (O_1827,N_19701,N_19571);
xnor UO_1828 (O_1828,N_19849,N_19612);
nand UO_1829 (O_1829,N_19823,N_19690);
nor UO_1830 (O_1830,N_19536,N_19294);
nor UO_1831 (O_1831,N_19609,N_19864);
nor UO_1832 (O_1832,N_19553,N_19996);
nand UO_1833 (O_1833,N_19852,N_19063);
nand UO_1834 (O_1834,N_19336,N_19088);
or UO_1835 (O_1835,N_19076,N_19046);
xor UO_1836 (O_1836,N_19019,N_19754);
nor UO_1837 (O_1837,N_19509,N_19234);
nor UO_1838 (O_1838,N_19417,N_19046);
nand UO_1839 (O_1839,N_19793,N_19584);
nand UO_1840 (O_1840,N_19586,N_19125);
nor UO_1841 (O_1841,N_19620,N_19801);
or UO_1842 (O_1842,N_19458,N_19856);
nor UO_1843 (O_1843,N_19818,N_19966);
or UO_1844 (O_1844,N_19857,N_19193);
nand UO_1845 (O_1845,N_19395,N_19771);
nand UO_1846 (O_1846,N_19262,N_19575);
or UO_1847 (O_1847,N_19256,N_19782);
nor UO_1848 (O_1848,N_19261,N_19255);
and UO_1849 (O_1849,N_19461,N_19925);
nor UO_1850 (O_1850,N_19199,N_19277);
and UO_1851 (O_1851,N_19689,N_19799);
and UO_1852 (O_1852,N_19890,N_19819);
nor UO_1853 (O_1853,N_19979,N_19369);
or UO_1854 (O_1854,N_19828,N_19384);
or UO_1855 (O_1855,N_19109,N_19717);
nand UO_1856 (O_1856,N_19813,N_19509);
xnor UO_1857 (O_1857,N_19743,N_19249);
or UO_1858 (O_1858,N_19058,N_19175);
nand UO_1859 (O_1859,N_19116,N_19315);
and UO_1860 (O_1860,N_19438,N_19564);
nor UO_1861 (O_1861,N_19212,N_19450);
xnor UO_1862 (O_1862,N_19848,N_19431);
nor UO_1863 (O_1863,N_19935,N_19614);
and UO_1864 (O_1864,N_19565,N_19193);
nor UO_1865 (O_1865,N_19471,N_19192);
nor UO_1866 (O_1866,N_19746,N_19918);
or UO_1867 (O_1867,N_19781,N_19810);
xnor UO_1868 (O_1868,N_19614,N_19768);
nand UO_1869 (O_1869,N_19157,N_19821);
xor UO_1870 (O_1870,N_19462,N_19339);
xor UO_1871 (O_1871,N_19557,N_19677);
and UO_1872 (O_1872,N_19883,N_19265);
xnor UO_1873 (O_1873,N_19198,N_19688);
nor UO_1874 (O_1874,N_19154,N_19816);
and UO_1875 (O_1875,N_19818,N_19532);
and UO_1876 (O_1876,N_19331,N_19086);
nor UO_1877 (O_1877,N_19030,N_19665);
or UO_1878 (O_1878,N_19714,N_19315);
and UO_1879 (O_1879,N_19163,N_19536);
or UO_1880 (O_1880,N_19311,N_19865);
or UO_1881 (O_1881,N_19051,N_19127);
xor UO_1882 (O_1882,N_19145,N_19074);
nand UO_1883 (O_1883,N_19079,N_19258);
nand UO_1884 (O_1884,N_19211,N_19846);
xnor UO_1885 (O_1885,N_19100,N_19422);
nor UO_1886 (O_1886,N_19310,N_19238);
nor UO_1887 (O_1887,N_19781,N_19851);
and UO_1888 (O_1888,N_19978,N_19761);
nand UO_1889 (O_1889,N_19029,N_19315);
xor UO_1890 (O_1890,N_19923,N_19771);
nand UO_1891 (O_1891,N_19255,N_19198);
xnor UO_1892 (O_1892,N_19930,N_19052);
or UO_1893 (O_1893,N_19315,N_19039);
or UO_1894 (O_1894,N_19852,N_19684);
and UO_1895 (O_1895,N_19882,N_19576);
and UO_1896 (O_1896,N_19435,N_19673);
nor UO_1897 (O_1897,N_19077,N_19776);
nor UO_1898 (O_1898,N_19203,N_19867);
and UO_1899 (O_1899,N_19948,N_19942);
and UO_1900 (O_1900,N_19628,N_19524);
nor UO_1901 (O_1901,N_19125,N_19755);
or UO_1902 (O_1902,N_19935,N_19703);
xor UO_1903 (O_1903,N_19378,N_19413);
or UO_1904 (O_1904,N_19247,N_19278);
xnor UO_1905 (O_1905,N_19231,N_19325);
nor UO_1906 (O_1906,N_19699,N_19816);
nor UO_1907 (O_1907,N_19618,N_19889);
nand UO_1908 (O_1908,N_19644,N_19031);
nand UO_1909 (O_1909,N_19088,N_19844);
nand UO_1910 (O_1910,N_19127,N_19498);
and UO_1911 (O_1911,N_19242,N_19367);
nand UO_1912 (O_1912,N_19103,N_19796);
nand UO_1913 (O_1913,N_19035,N_19434);
nor UO_1914 (O_1914,N_19172,N_19854);
nor UO_1915 (O_1915,N_19702,N_19408);
and UO_1916 (O_1916,N_19195,N_19237);
nand UO_1917 (O_1917,N_19931,N_19469);
nand UO_1918 (O_1918,N_19668,N_19927);
xor UO_1919 (O_1919,N_19106,N_19164);
xnor UO_1920 (O_1920,N_19236,N_19643);
xor UO_1921 (O_1921,N_19399,N_19133);
xor UO_1922 (O_1922,N_19969,N_19959);
and UO_1923 (O_1923,N_19055,N_19194);
nand UO_1924 (O_1924,N_19428,N_19927);
nand UO_1925 (O_1925,N_19140,N_19317);
nand UO_1926 (O_1926,N_19608,N_19720);
nor UO_1927 (O_1927,N_19040,N_19984);
nand UO_1928 (O_1928,N_19262,N_19946);
and UO_1929 (O_1929,N_19869,N_19136);
or UO_1930 (O_1930,N_19565,N_19618);
and UO_1931 (O_1931,N_19876,N_19394);
xnor UO_1932 (O_1932,N_19897,N_19022);
xnor UO_1933 (O_1933,N_19701,N_19512);
nand UO_1934 (O_1934,N_19825,N_19676);
nor UO_1935 (O_1935,N_19758,N_19374);
and UO_1936 (O_1936,N_19989,N_19706);
and UO_1937 (O_1937,N_19274,N_19744);
xor UO_1938 (O_1938,N_19610,N_19806);
and UO_1939 (O_1939,N_19740,N_19532);
nand UO_1940 (O_1940,N_19993,N_19111);
nand UO_1941 (O_1941,N_19975,N_19090);
nor UO_1942 (O_1942,N_19687,N_19679);
xor UO_1943 (O_1943,N_19448,N_19894);
xor UO_1944 (O_1944,N_19350,N_19689);
xnor UO_1945 (O_1945,N_19739,N_19838);
xor UO_1946 (O_1946,N_19027,N_19999);
or UO_1947 (O_1947,N_19248,N_19438);
nor UO_1948 (O_1948,N_19683,N_19177);
xor UO_1949 (O_1949,N_19860,N_19333);
nand UO_1950 (O_1950,N_19872,N_19621);
and UO_1951 (O_1951,N_19185,N_19005);
or UO_1952 (O_1952,N_19693,N_19427);
or UO_1953 (O_1953,N_19534,N_19936);
and UO_1954 (O_1954,N_19464,N_19590);
and UO_1955 (O_1955,N_19131,N_19078);
or UO_1956 (O_1956,N_19989,N_19524);
nand UO_1957 (O_1957,N_19476,N_19377);
or UO_1958 (O_1958,N_19090,N_19924);
nor UO_1959 (O_1959,N_19796,N_19998);
or UO_1960 (O_1960,N_19365,N_19854);
or UO_1961 (O_1961,N_19953,N_19382);
and UO_1962 (O_1962,N_19794,N_19954);
or UO_1963 (O_1963,N_19032,N_19365);
nand UO_1964 (O_1964,N_19139,N_19685);
nor UO_1965 (O_1965,N_19601,N_19230);
nor UO_1966 (O_1966,N_19591,N_19760);
and UO_1967 (O_1967,N_19295,N_19263);
and UO_1968 (O_1968,N_19146,N_19043);
xor UO_1969 (O_1969,N_19967,N_19461);
xnor UO_1970 (O_1970,N_19634,N_19689);
nand UO_1971 (O_1971,N_19548,N_19817);
xnor UO_1972 (O_1972,N_19879,N_19957);
xnor UO_1973 (O_1973,N_19543,N_19647);
nor UO_1974 (O_1974,N_19028,N_19849);
or UO_1975 (O_1975,N_19723,N_19169);
or UO_1976 (O_1976,N_19927,N_19638);
xor UO_1977 (O_1977,N_19681,N_19508);
nand UO_1978 (O_1978,N_19687,N_19076);
and UO_1979 (O_1979,N_19021,N_19058);
nand UO_1980 (O_1980,N_19808,N_19409);
xnor UO_1981 (O_1981,N_19364,N_19181);
or UO_1982 (O_1982,N_19208,N_19812);
nand UO_1983 (O_1983,N_19279,N_19740);
xnor UO_1984 (O_1984,N_19623,N_19841);
and UO_1985 (O_1985,N_19012,N_19096);
and UO_1986 (O_1986,N_19344,N_19209);
and UO_1987 (O_1987,N_19479,N_19754);
nand UO_1988 (O_1988,N_19908,N_19156);
nand UO_1989 (O_1989,N_19199,N_19952);
and UO_1990 (O_1990,N_19478,N_19878);
and UO_1991 (O_1991,N_19902,N_19144);
and UO_1992 (O_1992,N_19456,N_19670);
or UO_1993 (O_1993,N_19890,N_19932);
or UO_1994 (O_1994,N_19796,N_19421);
or UO_1995 (O_1995,N_19621,N_19694);
nand UO_1996 (O_1996,N_19900,N_19830);
nor UO_1997 (O_1997,N_19291,N_19975);
nand UO_1998 (O_1998,N_19113,N_19813);
or UO_1999 (O_1999,N_19720,N_19783);
and UO_2000 (O_2000,N_19471,N_19324);
nand UO_2001 (O_2001,N_19906,N_19130);
nand UO_2002 (O_2002,N_19065,N_19679);
or UO_2003 (O_2003,N_19340,N_19491);
and UO_2004 (O_2004,N_19096,N_19659);
or UO_2005 (O_2005,N_19944,N_19381);
nand UO_2006 (O_2006,N_19044,N_19116);
and UO_2007 (O_2007,N_19452,N_19556);
nand UO_2008 (O_2008,N_19918,N_19331);
nand UO_2009 (O_2009,N_19310,N_19566);
nor UO_2010 (O_2010,N_19782,N_19493);
or UO_2011 (O_2011,N_19524,N_19210);
nand UO_2012 (O_2012,N_19558,N_19909);
nand UO_2013 (O_2013,N_19747,N_19004);
nand UO_2014 (O_2014,N_19788,N_19020);
and UO_2015 (O_2015,N_19144,N_19827);
xor UO_2016 (O_2016,N_19434,N_19190);
and UO_2017 (O_2017,N_19190,N_19173);
nor UO_2018 (O_2018,N_19675,N_19631);
nand UO_2019 (O_2019,N_19797,N_19873);
or UO_2020 (O_2020,N_19738,N_19471);
or UO_2021 (O_2021,N_19587,N_19724);
or UO_2022 (O_2022,N_19085,N_19101);
or UO_2023 (O_2023,N_19004,N_19822);
nand UO_2024 (O_2024,N_19069,N_19283);
nor UO_2025 (O_2025,N_19150,N_19440);
nor UO_2026 (O_2026,N_19673,N_19359);
nand UO_2027 (O_2027,N_19100,N_19274);
and UO_2028 (O_2028,N_19992,N_19294);
nor UO_2029 (O_2029,N_19977,N_19442);
nand UO_2030 (O_2030,N_19265,N_19421);
or UO_2031 (O_2031,N_19351,N_19132);
or UO_2032 (O_2032,N_19678,N_19545);
or UO_2033 (O_2033,N_19640,N_19011);
nor UO_2034 (O_2034,N_19198,N_19037);
or UO_2035 (O_2035,N_19670,N_19766);
nand UO_2036 (O_2036,N_19290,N_19888);
and UO_2037 (O_2037,N_19254,N_19528);
or UO_2038 (O_2038,N_19640,N_19857);
and UO_2039 (O_2039,N_19820,N_19830);
nor UO_2040 (O_2040,N_19350,N_19910);
or UO_2041 (O_2041,N_19482,N_19239);
xnor UO_2042 (O_2042,N_19469,N_19990);
nor UO_2043 (O_2043,N_19430,N_19094);
nand UO_2044 (O_2044,N_19853,N_19768);
or UO_2045 (O_2045,N_19388,N_19050);
nand UO_2046 (O_2046,N_19740,N_19271);
and UO_2047 (O_2047,N_19488,N_19087);
xor UO_2048 (O_2048,N_19730,N_19833);
and UO_2049 (O_2049,N_19958,N_19318);
nor UO_2050 (O_2050,N_19778,N_19794);
and UO_2051 (O_2051,N_19782,N_19182);
nor UO_2052 (O_2052,N_19296,N_19532);
nor UO_2053 (O_2053,N_19260,N_19470);
or UO_2054 (O_2054,N_19836,N_19306);
nand UO_2055 (O_2055,N_19591,N_19073);
xnor UO_2056 (O_2056,N_19070,N_19719);
nor UO_2057 (O_2057,N_19651,N_19078);
xnor UO_2058 (O_2058,N_19861,N_19621);
and UO_2059 (O_2059,N_19424,N_19027);
or UO_2060 (O_2060,N_19020,N_19455);
nand UO_2061 (O_2061,N_19579,N_19721);
nand UO_2062 (O_2062,N_19391,N_19628);
and UO_2063 (O_2063,N_19925,N_19469);
nor UO_2064 (O_2064,N_19432,N_19921);
xnor UO_2065 (O_2065,N_19522,N_19209);
xnor UO_2066 (O_2066,N_19849,N_19901);
nor UO_2067 (O_2067,N_19745,N_19327);
or UO_2068 (O_2068,N_19666,N_19110);
nand UO_2069 (O_2069,N_19406,N_19268);
and UO_2070 (O_2070,N_19602,N_19691);
or UO_2071 (O_2071,N_19187,N_19943);
nand UO_2072 (O_2072,N_19528,N_19783);
or UO_2073 (O_2073,N_19173,N_19005);
nand UO_2074 (O_2074,N_19625,N_19399);
and UO_2075 (O_2075,N_19779,N_19648);
nor UO_2076 (O_2076,N_19327,N_19618);
nand UO_2077 (O_2077,N_19563,N_19363);
nor UO_2078 (O_2078,N_19768,N_19935);
xnor UO_2079 (O_2079,N_19685,N_19058);
nor UO_2080 (O_2080,N_19876,N_19573);
nand UO_2081 (O_2081,N_19664,N_19108);
and UO_2082 (O_2082,N_19056,N_19805);
and UO_2083 (O_2083,N_19476,N_19612);
nand UO_2084 (O_2084,N_19219,N_19958);
or UO_2085 (O_2085,N_19381,N_19695);
or UO_2086 (O_2086,N_19207,N_19929);
xnor UO_2087 (O_2087,N_19941,N_19692);
nor UO_2088 (O_2088,N_19525,N_19313);
or UO_2089 (O_2089,N_19478,N_19915);
or UO_2090 (O_2090,N_19155,N_19742);
xnor UO_2091 (O_2091,N_19980,N_19843);
nor UO_2092 (O_2092,N_19039,N_19087);
nor UO_2093 (O_2093,N_19969,N_19670);
nor UO_2094 (O_2094,N_19171,N_19283);
or UO_2095 (O_2095,N_19560,N_19584);
nand UO_2096 (O_2096,N_19789,N_19172);
xor UO_2097 (O_2097,N_19292,N_19044);
and UO_2098 (O_2098,N_19898,N_19840);
xor UO_2099 (O_2099,N_19658,N_19071);
nor UO_2100 (O_2100,N_19798,N_19056);
nor UO_2101 (O_2101,N_19456,N_19787);
nor UO_2102 (O_2102,N_19150,N_19382);
nor UO_2103 (O_2103,N_19154,N_19101);
or UO_2104 (O_2104,N_19684,N_19444);
nor UO_2105 (O_2105,N_19437,N_19991);
nor UO_2106 (O_2106,N_19939,N_19594);
or UO_2107 (O_2107,N_19140,N_19068);
nand UO_2108 (O_2108,N_19324,N_19098);
nand UO_2109 (O_2109,N_19114,N_19950);
and UO_2110 (O_2110,N_19948,N_19982);
xor UO_2111 (O_2111,N_19313,N_19583);
and UO_2112 (O_2112,N_19321,N_19864);
and UO_2113 (O_2113,N_19323,N_19325);
nand UO_2114 (O_2114,N_19113,N_19942);
nand UO_2115 (O_2115,N_19340,N_19577);
xnor UO_2116 (O_2116,N_19327,N_19378);
nand UO_2117 (O_2117,N_19823,N_19882);
nand UO_2118 (O_2118,N_19869,N_19326);
and UO_2119 (O_2119,N_19082,N_19872);
or UO_2120 (O_2120,N_19142,N_19697);
xnor UO_2121 (O_2121,N_19433,N_19024);
and UO_2122 (O_2122,N_19289,N_19761);
xor UO_2123 (O_2123,N_19458,N_19140);
xor UO_2124 (O_2124,N_19742,N_19072);
or UO_2125 (O_2125,N_19025,N_19878);
nor UO_2126 (O_2126,N_19130,N_19195);
and UO_2127 (O_2127,N_19677,N_19730);
nor UO_2128 (O_2128,N_19031,N_19682);
or UO_2129 (O_2129,N_19339,N_19207);
nand UO_2130 (O_2130,N_19514,N_19571);
nand UO_2131 (O_2131,N_19589,N_19197);
xor UO_2132 (O_2132,N_19949,N_19721);
nor UO_2133 (O_2133,N_19053,N_19098);
nand UO_2134 (O_2134,N_19552,N_19258);
and UO_2135 (O_2135,N_19966,N_19701);
nor UO_2136 (O_2136,N_19168,N_19403);
and UO_2137 (O_2137,N_19061,N_19898);
nor UO_2138 (O_2138,N_19302,N_19853);
nor UO_2139 (O_2139,N_19727,N_19851);
or UO_2140 (O_2140,N_19025,N_19703);
xnor UO_2141 (O_2141,N_19951,N_19420);
and UO_2142 (O_2142,N_19197,N_19285);
nand UO_2143 (O_2143,N_19743,N_19787);
and UO_2144 (O_2144,N_19418,N_19309);
and UO_2145 (O_2145,N_19840,N_19967);
xnor UO_2146 (O_2146,N_19933,N_19325);
xnor UO_2147 (O_2147,N_19227,N_19131);
nand UO_2148 (O_2148,N_19384,N_19242);
and UO_2149 (O_2149,N_19655,N_19623);
nand UO_2150 (O_2150,N_19051,N_19722);
nor UO_2151 (O_2151,N_19143,N_19183);
nor UO_2152 (O_2152,N_19786,N_19583);
or UO_2153 (O_2153,N_19073,N_19308);
and UO_2154 (O_2154,N_19259,N_19442);
and UO_2155 (O_2155,N_19501,N_19731);
or UO_2156 (O_2156,N_19441,N_19533);
nor UO_2157 (O_2157,N_19060,N_19905);
and UO_2158 (O_2158,N_19203,N_19508);
nand UO_2159 (O_2159,N_19002,N_19123);
and UO_2160 (O_2160,N_19897,N_19515);
nand UO_2161 (O_2161,N_19522,N_19234);
or UO_2162 (O_2162,N_19024,N_19510);
nand UO_2163 (O_2163,N_19145,N_19083);
or UO_2164 (O_2164,N_19881,N_19316);
and UO_2165 (O_2165,N_19599,N_19828);
or UO_2166 (O_2166,N_19023,N_19698);
or UO_2167 (O_2167,N_19857,N_19788);
nand UO_2168 (O_2168,N_19496,N_19107);
and UO_2169 (O_2169,N_19674,N_19779);
or UO_2170 (O_2170,N_19107,N_19660);
nand UO_2171 (O_2171,N_19113,N_19506);
xnor UO_2172 (O_2172,N_19513,N_19464);
or UO_2173 (O_2173,N_19197,N_19524);
xor UO_2174 (O_2174,N_19901,N_19646);
xor UO_2175 (O_2175,N_19519,N_19206);
nand UO_2176 (O_2176,N_19744,N_19291);
and UO_2177 (O_2177,N_19303,N_19860);
or UO_2178 (O_2178,N_19429,N_19546);
xor UO_2179 (O_2179,N_19490,N_19149);
or UO_2180 (O_2180,N_19534,N_19247);
or UO_2181 (O_2181,N_19982,N_19179);
and UO_2182 (O_2182,N_19737,N_19409);
nand UO_2183 (O_2183,N_19345,N_19991);
nor UO_2184 (O_2184,N_19334,N_19395);
or UO_2185 (O_2185,N_19642,N_19501);
xor UO_2186 (O_2186,N_19557,N_19904);
xnor UO_2187 (O_2187,N_19590,N_19581);
or UO_2188 (O_2188,N_19677,N_19592);
nand UO_2189 (O_2189,N_19454,N_19219);
nor UO_2190 (O_2190,N_19752,N_19178);
nand UO_2191 (O_2191,N_19475,N_19915);
xor UO_2192 (O_2192,N_19994,N_19175);
nor UO_2193 (O_2193,N_19090,N_19131);
nand UO_2194 (O_2194,N_19007,N_19327);
and UO_2195 (O_2195,N_19807,N_19178);
xor UO_2196 (O_2196,N_19205,N_19111);
nor UO_2197 (O_2197,N_19348,N_19212);
and UO_2198 (O_2198,N_19015,N_19825);
xor UO_2199 (O_2199,N_19321,N_19521);
xnor UO_2200 (O_2200,N_19806,N_19564);
and UO_2201 (O_2201,N_19610,N_19402);
nand UO_2202 (O_2202,N_19069,N_19510);
nor UO_2203 (O_2203,N_19254,N_19309);
nor UO_2204 (O_2204,N_19499,N_19092);
nor UO_2205 (O_2205,N_19264,N_19271);
and UO_2206 (O_2206,N_19300,N_19090);
or UO_2207 (O_2207,N_19951,N_19659);
and UO_2208 (O_2208,N_19562,N_19782);
nand UO_2209 (O_2209,N_19170,N_19676);
and UO_2210 (O_2210,N_19105,N_19040);
nand UO_2211 (O_2211,N_19016,N_19849);
or UO_2212 (O_2212,N_19949,N_19503);
and UO_2213 (O_2213,N_19955,N_19328);
xor UO_2214 (O_2214,N_19471,N_19233);
nand UO_2215 (O_2215,N_19918,N_19771);
or UO_2216 (O_2216,N_19904,N_19187);
or UO_2217 (O_2217,N_19244,N_19887);
nand UO_2218 (O_2218,N_19855,N_19698);
nand UO_2219 (O_2219,N_19085,N_19244);
xnor UO_2220 (O_2220,N_19877,N_19717);
xnor UO_2221 (O_2221,N_19115,N_19171);
or UO_2222 (O_2222,N_19189,N_19548);
xnor UO_2223 (O_2223,N_19349,N_19838);
nand UO_2224 (O_2224,N_19319,N_19732);
xor UO_2225 (O_2225,N_19091,N_19990);
or UO_2226 (O_2226,N_19752,N_19403);
and UO_2227 (O_2227,N_19854,N_19238);
nand UO_2228 (O_2228,N_19054,N_19349);
xor UO_2229 (O_2229,N_19451,N_19345);
and UO_2230 (O_2230,N_19318,N_19393);
nor UO_2231 (O_2231,N_19026,N_19711);
or UO_2232 (O_2232,N_19859,N_19654);
or UO_2233 (O_2233,N_19319,N_19321);
nor UO_2234 (O_2234,N_19987,N_19671);
nor UO_2235 (O_2235,N_19209,N_19178);
nor UO_2236 (O_2236,N_19505,N_19246);
xor UO_2237 (O_2237,N_19959,N_19193);
and UO_2238 (O_2238,N_19422,N_19764);
and UO_2239 (O_2239,N_19952,N_19417);
xnor UO_2240 (O_2240,N_19204,N_19559);
or UO_2241 (O_2241,N_19891,N_19215);
nor UO_2242 (O_2242,N_19068,N_19355);
and UO_2243 (O_2243,N_19353,N_19238);
nor UO_2244 (O_2244,N_19897,N_19423);
or UO_2245 (O_2245,N_19644,N_19872);
and UO_2246 (O_2246,N_19574,N_19540);
or UO_2247 (O_2247,N_19485,N_19080);
xor UO_2248 (O_2248,N_19606,N_19176);
nand UO_2249 (O_2249,N_19218,N_19303);
or UO_2250 (O_2250,N_19428,N_19757);
nor UO_2251 (O_2251,N_19010,N_19212);
and UO_2252 (O_2252,N_19787,N_19832);
xnor UO_2253 (O_2253,N_19699,N_19944);
and UO_2254 (O_2254,N_19746,N_19259);
nand UO_2255 (O_2255,N_19292,N_19013);
nor UO_2256 (O_2256,N_19638,N_19981);
nor UO_2257 (O_2257,N_19829,N_19606);
and UO_2258 (O_2258,N_19498,N_19787);
and UO_2259 (O_2259,N_19156,N_19115);
and UO_2260 (O_2260,N_19693,N_19238);
xnor UO_2261 (O_2261,N_19384,N_19107);
nor UO_2262 (O_2262,N_19446,N_19511);
or UO_2263 (O_2263,N_19225,N_19188);
nor UO_2264 (O_2264,N_19823,N_19990);
nor UO_2265 (O_2265,N_19224,N_19832);
and UO_2266 (O_2266,N_19241,N_19132);
or UO_2267 (O_2267,N_19142,N_19647);
and UO_2268 (O_2268,N_19043,N_19993);
nand UO_2269 (O_2269,N_19382,N_19804);
nor UO_2270 (O_2270,N_19689,N_19626);
xnor UO_2271 (O_2271,N_19790,N_19399);
nor UO_2272 (O_2272,N_19157,N_19580);
and UO_2273 (O_2273,N_19216,N_19025);
nand UO_2274 (O_2274,N_19849,N_19054);
nand UO_2275 (O_2275,N_19078,N_19639);
nand UO_2276 (O_2276,N_19849,N_19684);
and UO_2277 (O_2277,N_19634,N_19677);
nor UO_2278 (O_2278,N_19172,N_19264);
nor UO_2279 (O_2279,N_19653,N_19984);
and UO_2280 (O_2280,N_19734,N_19472);
xor UO_2281 (O_2281,N_19167,N_19674);
or UO_2282 (O_2282,N_19026,N_19057);
and UO_2283 (O_2283,N_19922,N_19341);
nand UO_2284 (O_2284,N_19309,N_19138);
or UO_2285 (O_2285,N_19009,N_19531);
nand UO_2286 (O_2286,N_19108,N_19277);
or UO_2287 (O_2287,N_19445,N_19012);
nor UO_2288 (O_2288,N_19079,N_19255);
and UO_2289 (O_2289,N_19362,N_19366);
or UO_2290 (O_2290,N_19392,N_19309);
nand UO_2291 (O_2291,N_19250,N_19437);
xor UO_2292 (O_2292,N_19760,N_19514);
nor UO_2293 (O_2293,N_19966,N_19073);
nor UO_2294 (O_2294,N_19346,N_19420);
or UO_2295 (O_2295,N_19952,N_19927);
nor UO_2296 (O_2296,N_19802,N_19146);
xor UO_2297 (O_2297,N_19959,N_19976);
nor UO_2298 (O_2298,N_19571,N_19465);
nand UO_2299 (O_2299,N_19402,N_19282);
nand UO_2300 (O_2300,N_19970,N_19040);
nand UO_2301 (O_2301,N_19056,N_19086);
and UO_2302 (O_2302,N_19969,N_19578);
nor UO_2303 (O_2303,N_19594,N_19432);
xnor UO_2304 (O_2304,N_19436,N_19816);
or UO_2305 (O_2305,N_19372,N_19656);
nor UO_2306 (O_2306,N_19612,N_19208);
xor UO_2307 (O_2307,N_19426,N_19221);
nand UO_2308 (O_2308,N_19298,N_19669);
xnor UO_2309 (O_2309,N_19861,N_19385);
or UO_2310 (O_2310,N_19518,N_19407);
nand UO_2311 (O_2311,N_19088,N_19823);
or UO_2312 (O_2312,N_19086,N_19625);
nor UO_2313 (O_2313,N_19308,N_19909);
and UO_2314 (O_2314,N_19301,N_19003);
xnor UO_2315 (O_2315,N_19003,N_19108);
nand UO_2316 (O_2316,N_19198,N_19112);
or UO_2317 (O_2317,N_19309,N_19929);
nor UO_2318 (O_2318,N_19774,N_19940);
or UO_2319 (O_2319,N_19857,N_19375);
nand UO_2320 (O_2320,N_19613,N_19565);
and UO_2321 (O_2321,N_19225,N_19914);
or UO_2322 (O_2322,N_19324,N_19905);
xor UO_2323 (O_2323,N_19441,N_19220);
xnor UO_2324 (O_2324,N_19990,N_19385);
or UO_2325 (O_2325,N_19100,N_19961);
or UO_2326 (O_2326,N_19685,N_19024);
nor UO_2327 (O_2327,N_19808,N_19889);
or UO_2328 (O_2328,N_19587,N_19536);
and UO_2329 (O_2329,N_19835,N_19174);
nor UO_2330 (O_2330,N_19324,N_19637);
and UO_2331 (O_2331,N_19913,N_19995);
nand UO_2332 (O_2332,N_19943,N_19811);
or UO_2333 (O_2333,N_19289,N_19228);
or UO_2334 (O_2334,N_19359,N_19015);
and UO_2335 (O_2335,N_19223,N_19203);
xnor UO_2336 (O_2336,N_19253,N_19622);
nand UO_2337 (O_2337,N_19206,N_19788);
xnor UO_2338 (O_2338,N_19154,N_19282);
and UO_2339 (O_2339,N_19036,N_19438);
or UO_2340 (O_2340,N_19681,N_19295);
or UO_2341 (O_2341,N_19822,N_19144);
nand UO_2342 (O_2342,N_19653,N_19946);
and UO_2343 (O_2343,N_19502,N_19549);
or UO_2344 (O_2344,N_19526,N_19941);
nor UO_2345 (O_2345,N_19553,N_19757);
xor UO_2346 (O_2346,N_19016,N_19831);
nor UO_2347 (O_2347,N_19277,N_19681);
nand UO_2348 (O_2348,N_19076,N_19968);
and UO_2349 (O_2349,N_19020,N_19258);
or UO_2350 (O_2350,N_19085,N_19379);
xnor UO_2351 (O_2351,N_19478,N_19157);
xnor UO_2352 (O_2352,N_19823,N_19205);
and UO_2353 (O_2353,N_19074,N_19015);
nor UO_2354 (O_2354,N_19550,N_19027);
or UO_2355 (O_2355,N_19339,N_19331);
xor UO_2356 (O_2356,N_19744,N_19475);
nor UO_2357 (O_2357,N_19194,N_19632);
nor UO_2358 (O_2358,N_19831,N_19928);
nand UO_2359 (O_2359,N_19612,N_19499);
nand UO_2360 (O_2360,N_19631,N_19489);
xnor UO_2361 (O_2361,N_19933,N_19006);
or UO_2362 (O_2362,N_19258,N_19902);
nand UO_2363 (O_2363,N_19636,N_19328);
and UO_2364 (O_2364,N_19447,N_19574);
xor UO_2365 (O_2365,N_19293,N_19248);
or UO_2366 (O_2366,N_19863,N_19304);
or UO_2367 (O_2367,N_19156,N_19539);
xor UO_2368 (O_2368,N_19349,N_19835);
or UO_2369 (O_2369,N_19148,N_19169);
xor UO_2370 (O_2370,N_19533,N_19034);
and UO_2371 (O_2371,N_19366,N_19017);
and UO_2372 (O_2372,N_19105,N_19901);
or UO_2373 (O_2373,N_19092,N_19767);
and UO_2374 (O_2374,N_19705,N_19326);
nor UO_2375 (O_2375,N_19320,N_19647);
nor UO_2376 (O_2376,N_19589,N_19852);
and UO_2377 (O_2377,N_19841,N_19190);
and UO_2378 (O_2378,N_19843,N_19327);
xnor UO_2379 (O_2379,N_19719,N_19247);
nor UO_2380 (O_2380,N_19656,N_19230);
nand UO_2381 (O_2381,N_19645,N_19035);
xnor UO_2382 (O_2382,N_19715,N_19885);
nor UO_2383 (O_2383,N_19046,N_19131);
or UO_2384 (O_2384,N_19759,N_19046);
and UO_2385 (O_2385,N_19395,N_19305);
and UO_2386 (O_2386,N_19117,N_19712);
xnor UO_2387 (O_2387,N_19752,N_19886);
xor UO_2388 (O_2388,N_19058,N_19889);
xor UO_2389 (O_2389,N_19395,N_19538);
and UO_2390 (O_2390,N_19039,N_19587);
nor UO_2391 (O_2391,N_19723,N_19900);
or UO_2392 (O_2392,N_19212,N_19419);
nor UO_2393 (O_2393,N_19158,N_19210);
and UO_2394 (O_2394,N_19997,N_19151);
and UO_2395 (O_2395,N_19384,N_19779);
nor UO_2396 (O_2396,N_19278,N_19601);
and UO_2397 (O_2397,N_19054,N_19194);
or UO_2398 (O_2398,N_19046,N_19154);
or UO_2399 (O_2399,N_19063,N_19276);
xnor UO_2400 (O_2400,N_19130,N_19234);
or UO_2401 (O_2401,N_19705,N_19730);
and UO_2402 (O_2402,N_19279,N_19131);
nor UO_2403 (O_2403,N_19966,N_19438);
or UO_2404 (O_2404,N_19758,N_19207);
xnor UO_2405 (O_2405,N_19814,N_19225);
xnor UO_2406 (O_2406,N_19764,N_19343);
nor UO_2407 (O_2407,N_19886,N_19039);
xor UO_2408 (O_2408,N_19748,N_19369);
nand UO_2409 (O_2409,N_19267,N_19055);
nor UO_2410 (O_2410,N_19751,N_19238);
nor UO_2411 (O_2411,N_19195,N_19811);
xor UO_2412 (O_2412,N_19890,N_19289);
xnor UO_2413 (O_2413,N_19144,N_19805);
or UO_2414 (O_2414,N_19122,N_19593);
xnor UO_2415 (O_2415,N_19299,N_19592);
nand UO_2416 (O_2416,N_19326,N_19429);
and UO_2417 (O_2417,N_19473,N_19174);
and UO_2418 (O_2418,N_19235,N_19807);
xnor UO_2419 (O_2419,N_19889,N_19533);
nor UO_2420 (O_2420,N_19439,N_19191);
nand UO_2421 (O_2421,N_19917,N_19725);
and UO_2422 (O_2422,N_19586,N_19583);
or UO_2423 (O_2423,N_19968,N_19386);
and UO_2424 (O_2424,N_19959,N_19481);
xor UO_2425 (O_2425,N_19309,N_19182);
xor UO_2426 (O_2426,N_19066,N_19914);
nor UO_2427 (O_2427,N_19536,N_19414);
or UO_2428 (O_2428,N_19106,N_19311);
or UO_2429 (O_2429,N_19040,N_19639);
and UO_2430 (O_2430,N_19213,N_19815);
and UO_2431 (O_2431,N_19914,N_19995);
nand UO_2432 (O_2432,N_19471,N_19828);
xnor UO_2433 (O_2433,N_19739,N_19634);
nand UO_2434 (O_2434,N_19360,N_19690);
nor UO_2435 (O_2435,N_19482,N_19553);
or UO_2436 (O_2436,N_19101,N_19667);
xor UO_2437 (O_2437,N_19483,N_19585);
and UO_2438 (O_2438,N_19761,N_19011);
nor UO_2439 (O_2439,N_19048,N_19163);
xnor UO_2440 (O_2440,N_19869,N_19005);
or UO_2441 (O_2441,N_19290,N_19949);
xor UO_2442 (O_2442,N_19059,N_19974);
and UO_2443 (O_2443,N_19166,N_19896);
nand UO_2444 (O_2444,N_19292,N_19285);
or UO_2445 (O_2445,N_19640,N_19783);
nand UO_2446 (O_2446,N_19979,N_19612);
xnor UO_2447 (O_2447,N_19113,N_19245);
nor UO_2448 (O_2448,N_19428,N_19362);
nand UO_2449 (O_2449,N_19780,N_19401);
xnor UO_2450 (O_2450,N_19695,N_19866);
nor UO_2451 (O_2451,N_19114,N_19509);
and UO_2452 (O_2452,N_19199,N_19620);
xnor UO_2453 (O_2453,N_19237,N_19601);
nor UO_2454 (O_2454,N_19294,N_19230);
and UO_2455 (O_2455,N_19008,N_19194);
or UO_2456 (O_2456,N_19893,N_19759);
or UO_2457 (O_2457,N_19564,N_19863);
xor UO_2458 (O_2458,N_19610,N_19613);
or UO_2459 (O_2459,N_19028,N_19900);
nor UO_2460 (O_2460,N_19918,N_19723);
and UO_2461 (O_2461,N_19884,N_19501);
or UO_2462 (O_2462,N_19835,N_19809);
nand UO_2463 (O_2463,N_19350,N_19781);
and UO_2464 (O_2464,N_19222,N_19149);
nand UO_2465 (O_2465,N_19575,N_19478);
nor UO_2466 (O_2466,N_19914,N_19460);
and UO_2467 (O_2467,N_19812,N_19052);
nor UO_2468 (O_2468,N_19591,N_19841);
or UO_2469 (O_2469,N_19655,N_19369);
xnor UO_2470 (O_2470,N_19285,N_19740);
nand UO_2471 (O_2471,N_19111,N_19123);
nand UO_2472 (O_2472,N_19297,N_19504);
nor UO_2473 (O_2473,N_19870,N_19586);
and UO_2474 (O_2474,N_19290,N_19935);
and UO_2475 (O_2475,N_19171,N_19170);
nand UO_2476 (O_2476,N_19736,N_19516);
nor UO_2477 (O_2477,N_19974,N_19172);
xor UO_2478 (O_2478,N_19248,N_19691);
or UO_2479 (O_2479,N_19734,N_19975);
nand UO_2480 (O_2480,N_19098,N_19969);
xor UO_2481 (O_2481,N_19896,N_19250);
nand UO_2482 (O_2482,N_19386,N_19146);
nand UO_2483 (O_2483,N_19927,N_19726);
and UO_2484 (O_2484,N_19435,N_19236);
nor UO_2485 (O_2485,N_19054,N_19373);
or UO_2486 (O_2486,N_19573,N_19723);
nor UO_2487 (O_2487,N_19005,N_19699);
or UO_2488 (O_2488,N_19113,N_19133);
and UO_2489 (O_2489,N_19562,N_19411);
xnor UO_2490 (O_2490,N_19576,N_19779);
nor UO_2491 (O_2491,N_19381,N_19083);
or UO_2492 (O_2492,N_19142,N_19349);
and UO_2493 (O_2493,N_19650,N_19944);
and UO_2494 (O_2494,N_19796,N_19248);
and UO_2495 (O_2495,N_19423,N_19860);
nor UO_2496 (O_2496,N_19423,N_19039);
xor UO_2497 (O_2497,N_19052,N_19139);
nand UO_2498 (O_2498,N_19377,N_19622);
and UO_2499 (O_2499,N_19692,N_19146);
endmodule