module basic_1500_15000_2000_15_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
xnor U0 (N_0,In_376,In_1413);
or U1 (N_1,In_617,In_296);
or U2 (N_2,In_533,In_458);
or U3 (N_3,In_1262,In_61);
and U4 (N_4,In_687,In_993);
nand U5 (N_5,In_1397,In_1098);
or U6 (N_6,In_947,In_1154);
or U7 (N_7,In_1119,In_123);
xnor U8 (N_8,In_36,In_959);
xor U9 (N_9,In_1088,In_148);
xnor U10 (N_10,In_1077,In_900);
and U11 (N_11,In_764,In_1036);
and U12 (N_12,In_1312,In_1275);
xor U13 (N_13,In_1375,In_1206);
xnor U14 (N_14,In_147,In_1247);
xor U15 (N_15,In_1089,In_240);
nor U16 (N_16,In_786,In_1134);
or U17 (N_17,In_840,In_42);
nor U18 (N_18,In_49,In_772);
or U19 (N_19,In_310,In_386);
and U20 (N_20,In_1430,In_1319);
and U21 (N_21,In_856,In_655);
nor U22 (N_22,In_737,In_1014);
nor U23 (N_23,In_428,In_534);
and U24 (N_24,In_849,In_285);
and U25 (N_25,In_940,In_124);
or U26 (N_26,In_1172,In_1015);
xor U27 (N_27,In_438,In_1309);
and U28 (N_28,In_746,In_499);
and U29 (N_29,In_466,In_629);
nor U30 (N_30,In_524,In_835);
xor U31 (N_31,In_1210,In_38);
nand U32 (N_32,In_640,In_468);
nand U33 (N_33,In_185,In_1257);
nand U34 (N_34,In_754,In_1085);
nand U35 (N_35,In_212,In_1341);
nor U36 (N_36,In_1409,In_674);
or U37 (N_37,In_872,In_348);
nand U38 (N_38,In_707,In_1133);
or U39 (N_39,In_908,In_1293);
nor U40 (N_40,In_1388,In_660);
nand U41 (N_41,In_1016,In_99);
and U42 (N_42,In_816,In_1083);
or U43 (N_43,In_383,In_274);
nand U44 (N_44,In_919,In_1436);
nand U45 (N_45,In_1040,In_1153);
xnor U46 (N_46,In_1294,In_1452);
or U47 (N_47,In_1289,In_489);
nor U48 (N_48,In_168,In_1197);
nor U49 (N_49,In_1118,In_836);
nor U50 (N_50,In_1466,In_432);
and U51 (N_51,In_289,In_867);
nor U52 (N_52,In_1403,In_622);
nand U53 (N_53,In_697,In_479);
nand U54 (N_54,In_39,In_1214);
nor U55 (N_55,In_1495,In_1389);
xnor U56 (N_56,In_602,In_437);
xnor U57 (N_57,In_1378,In_1107);
or U58 (N_58,In_630,In_680);
or U59 (N_59,In_1104,In_664);
or U60 (N_60,In_1433,In_619);
xnor U61 (N_61,In_190,In_1062);
xor U62 (N_62,In_1497,In_497);
nand U63 (N_63,In_284,In_1351);
xnor U64 (N_64,In_876,In_1058);
and U65 (N_65,In_1043,In_583);
xor U66 (N_66,In_1039,In_986);
nand U67 (N_67,In_971,In_248);
or U68 (N_68,In_823,In_160);
or U69 (N_69,In_145,In_899);
or U70 (N_70,In_1122,In_1001);
nor U71 (N_71,In_1417,In_1486);
nor U72 (N_72,In_9,In_1229);
or U73 (N_73,In_1344,In_946);
nand U74 (N_74,In_738,In_43);
nand U75 (N_75,In_1434,In_1410);
xnor U76 (N_76,In_396,In_1087);
or U77 (N_77,In_958,In_542);
or U78 (N_78,In_795,In_1463);
and U79 (N_79,In_25,In_588);
or U80 (N_80,In_734,In_684);
and U81 (N_81,In_1281,In_631);
xnor U82 (N_82,In_834,In_1);
nor U83 (N_83,In_1349,In_1221);
nor U84 (N_84,In_1476,In_914);
nor U85 (N_85,In_71,In_1232);
nand U86 (N_86,In_1472,In_311);
nor U87 (N_87,In_865,In_594);
or U88 (N_88,In_564,In_1359);
and U89 (N_89,In_244,In_930);
nor U90 (N_90,In_1330,In_1189);
and U91 (N_91,In_561,In_1475);
xnor U92 (N_92,In_85,In_1228);
nor U93 (N_93,In_554,In_552);
or U94 (N_94,In_1110,In_1424);
xnor U95 (N_95,In_997,In_33);
nand U96 (N_96,In_167,In_1004);
and U97 (N_97,In_643,In_1178);
nor U98 (N_98,In_101,In_1167);
nor U99 (N_99,In_681,In_1314);
xor U100 (N_100,In_863,In_650);
and U101 (N_101,In_722,In_58);
xor U102 (N_102,In_480,In_1018);
or U103 (N_103,In_464,In_339);
nor U104 (N_104,In_1093,In_1169);
xor U105 (N_105,In_418,In_1211);
xnor U106 (N_106,In_105,In_559);
nor U107 (N_107,In_609,In_515);
nor U108 (N_108,In_125,In_106);
nand U109 (N_109,In_1131,In_1129);
or U110 (N_110,In_275,In_1428);
and U111 (N_111,In_201,In_952);
nor U112 (N_112,In_1165,In_478);
or U113 (N_113,In_291,In_1171);
xnor U114 (N_114,In_313,In_1235);
and U115 (N_115,In_424,In_885);
and U116 (N_116,In_12,In_682);
nor U117 (N_117,In_400,In_35);
nor U118 (N_118,In_637,In_365);
nand U119 (N_119,In_693,In_491);
nor U120 (N_120,In_111,In_232);
xor U121 (N_121,In_1261,In_492);
xnor U122 (N_122,In_98,In_255);
nor U123 (N_123,In_1074,In_1381);
or U124 (N_124,In_175,In_522);
nand U125 (N_125,In_1499,In_457);
nand U126 (N_126,In_761,In_937);
or U127 (N_127,In_1082,In_139);
nand U128 (N_128,In_558,In_380);
nor U129 (N_129,In_670,In_1391);
nor U130 (N_130,In_721,In_537);
nand U131 (N_131,In_736,In_1465);
nor U132 (N_132,In_954,In_1163);
xor U133 (N_133,In_186,In_1300);
or U134 (N_134,In_1310,In_1464);
nand U135 (N_135,In_1271,In_368);
or U136 (N_136,In_1138,In_1263);
nor U137 (N_137,In_581,In_352);
nand U138 (N_138,In_525,In_1361);
or U139 (N_139,In_1490,In_505);
nand U140 (N_140,In_1055,In_174);
and U141 (N_141,In_511,In_961);
and U142 (N_142,In_1320,In_1173);
xnor U143 (N_143,In_1485,In_1356);
nand U144 (N_144,In_1045,In_1177);
and U145 (N_145,In_1066,In_1092);
nor U146 (N_146,In_362,In_1205);
and U147 (N_147,In_950,In_1095);
or U148 (N_148,In_226,In_612);
or U149 (N_149,In_749,In_985);
or U150 (N_150,In_370,In_633);
and U151 (N_151,In_116,In_1149);
nand U152 (N_152,In_570,In_213);
nand U153 (N_153,In_502,In_1382);
xor U154 (N_154,In_685,In_820);
xnor U155 (N_155,In_742,In_977);
nand U156 (N_156,In_1373,In_973);
nand U157 (N_157,In_211,In_1064);
nand U158 (N_158,In_1333,In_1393);
or U159 (N_159,In_1362,In_371);
xor U160 (N_160,In_803,In_547);
or U161 (N_161,In_1184,In_936);
nand U162 (N_162,In_50,In_157);
or U163 (N_163,In_938,In_845);
xor U164 (N_164,In_1008,In_812);
xor U165 (N_165,In_328,In_1164);
xnor U166 (N_166,In_253,In_364);
or U167 (N_167,In_51,In_1317);
nand U168 (N_168,In_1020,In_566);
nand U169 (N_169,In_575,In_701);
xnor U170 (N_170,In_421,In_394);
xnor U171 (N_171,In_805,In_273);
or U172 (N_172,In_47,In_102);
nand U173 (N_173,In_1297,In_1038);
nor U174 (N_174,In_1268,In_1299);
nand U175 (N_175,In_735,In_790);
nand U176 (N_176,In_52,In_590);
and U177 (N_177,In_725,In_1226);
or U178 (N_178,In_131,In_1260);
nor U179 (N_179,In_657,In_1421);
xor U180 (N_180,In_1084,In_374);
and U181 (N_181,In_1343,In_819);
nor U182 (N_182,In_994,In_504);
xnor U183 (N_183,In_603,In_1203);
and U184 (N_184,In_409,In_1147);
and U185 (N_185,In_1387,In_196);
nor U186 (N_186,In_327,In_259);
xnor U187 (N_187,In_203,In_1254);
or U188 (N_188,In_1425,In_976);
nor U189 (N_189,In_1030,In_892);
nor U190 (N_190,In_829,In_1304);
or U191 (N_191,In_312,In_119);
xnor U192 (N_192,In_452,In_1029);
and U193 (N_193,In_1049,In_1065);
nor U194 (N_194,In_205,In_903);
or U195 (N_195,In_162,In_960);
nor U196 (N_196,In_426,In_978);
xor U197 (N_197,In_719,In_935);
and U198 (N_198,In_818,In_726);
and U199 (N_199,In_1048,In_349);
or U200 (N_200,In_1477,In_1116);
or U201 (N_201,In_76,In_165);
and U202 (N_202,In_1284,In_995);
or U203 (N_203,In_912,In_1140);
nor U204 (N_204,In_569,In_484);
nor U205 (N_205,In_811,In_614);
and U206 (N_206,In_898,In_1455);
nor U207 (N_207,In_623,In_28);
nor U208 (N_208,In_1287,In_906);
or U209 (N_209,In_733,In_883);
nor U210 (N_210,In_427,In_57);
or U211 (N_211,In_1415,In_846);
or U212 (N_212,In_925,In_5);
and U213 (N_213,In_1017,In_268);
nand U214 (N_214,In_1223,In_783);
nand U215 (N_215,In_359,In_1158);
nor U216 (N_216,In_606,In_546);
nand U217 (N_217,In_460,In_957);
xor U218 (N_218,In_1419,In_269);
nand U219 (N_219,In_708,In_895);
and U220 (N_220,In_228,In_1322);
xnor U221 (N_221,In_1108,In_412);
or U222 (N_222,In_766,In_1059);
nor U223 (N_223,In_1142,In_723);
or U224 (N_224,In_227,In_880);
xnor U225 (N_225,In_1494,In_765);
nand U226 (N_226,In_858,In_1446);
or U227 (N_227,In_875,In_854);
nand U228 (N_228,In_267,In_1234);
or U229 (N_229,In_140,In_222);
and U230 (N_230,In_981,In_1101);
nand U231 (N_231,In_340,In_663);
xnor U232 (N_232,In_709,In_75);
nand U233 (N_233,In_577,In_864);
and U234 (N_234,In_506,In_1240);
nor U235 (N_235,In_369,In_1233);
or U236 (N_236,In_1480,In_449);
xor U237 (N_237,In_16,In_1061);
nor U238 (N_238,In_1220,In_11);
or U239 (N_239,In_990,In_776);
and U240 (N_240,In_1208,In_444);
and U241 (N_241,In_901,In_377);
xnor U242 (N_242,In_473,In_454);
and U243 (N_243,In_481,In_1461);
nor U244 (N_244,In_115,In_679);
nor U245 (N_245,In_399,In_431);
nand U246 (N_246,In_634,In_344);
nand U247 (N_247,In_1236,In_354);
or U248 (N_248,In_367,In_1003);
nand U249 (N_249,In_644,In_4);
nor U250 (N_250,In_214,In_200);
nand U251 (N_251,In_341,In_405);
nor U252 (N_252,In_917,In_87);
nor U253 (N_253,In_1423,In_60);
nor U254 (N_254,In_792,In_172);
xnor U255 (N_255,In_962,In_675);
nor U256 (N_256,In_1002,In_14);
or U257 (N_257,In_455,In_53);
and U258 (N_258,In_249,In_1407);
xnor U259 (N_259,In_1288,In_1292);
nor U260 (N_260,In_1435,In_1347);
or U261 (N_261,In_1286,In_921);
xnor U262 (N_262,In_844,In_1102);
nand U263 (N_263,In_309,In_926);
or U264 (N_264,In_745,In_624);
nand U265 (N_265,In_404,In_1224);
and U266 (N_266,In_668,In_821);
and U267 (N_267,In_616,In_331);
xor U268 (N_268,In_462,In_530);
xor U269 (N_269,In_688,In_1483);
and U270 (N_270,In_218,In_955);
xnor U271 (N_271,In_142,In_1051);
nand U272 (N_272,In_905,In_910);
nand U273 (N_273,In_1367,In_1174);
and U274 (N_274,In_31,In_870);
xnor U275 (N_275,In_1324,In_526);
or U276 (N_276,In_804,In_155);
nor U277 (N_277,In_774,In_611);
nor U278 (N_278,In_389,In_652);
or U279 (N_279,In_1239,In_346);
and U280 (N_280,In_1376,In_326);
nand U281 (N_281,In_563,In_571);
nor U282 (N_282,In_690,In_136);
xor U283 (N_283,In_1075,In_597);
and U284 (N_284,In_689,In_632);
and U285 (N_285,In_81,In_665);
nor U286 (N_286,In_320,In_277);
nand U287 (N_287,In_1068,In_306);
nor U288 (N_288,In_177,In_146);
nand U289 (N_289,In_1241,In_715);
nand U290 (N_290,In_1256,In_621);
nor U291 (N_291,In_841,In_440);
xnor U292 (N_292,In_1010,In_1360);
xor U293 (N_293,In_107,In_265);
and U294 (N_294,In_387,In_314);
xor U295 (N_295,In_860,In_223);
xor U296 (N_296,In_782,In_945);
xnor U297 (N_297,In_1350,In_673);
xor U298 (N_298,In_27,In_448);
nand U299 (N_299,In_984,In_1250);
and U300 (N_300,In_728,In_951);
xor U301 (N_301,In_785,In_839);
nand U302 (N_302,In_1371,In_953);
and U303 (N_303,In_262,In_732);
or U304 (N_304,In_613,In_1069);
nand U305 (N_305,In_1188,In_756);
and U306 (N_306,In_158,In_1469);
or U307 (N_307,In_360,In_23);
and U308 (N_308,In_843,In_392);
xor U309 (N_309,In_797,In_272);
or U310 (N_310,In_1473,In_271);
nand U311 (N_311,In_1230,In_808);
nor U312 (N_312,In_302,In_591);
and U313 (N_313,In_1355,In_1202);
and U314 (N_314,In_996,In_1152);
nand U315 (N_315,In_980,In_1481);
xnor U316 (N_316,In_388,In_292);
or U317 (N_317,In_198,In_800);
and U318 (N_318,In_514,In_2);
nor U319 (N_319,In_894,In_467);
or U320 (N_320,In_1308,In_1144);
nand U321 (N_321,In_104,In_300);
xnor U322 (N_322,In_550,In_618);
and U323 (N_323,In_1328,In_886);
and U324 (N_324,In_784,In_1081);
nand U325 (N_325,In_813,In_403);
and U326 (N_326,In_238,In_1353);
or U327 (N_327,In_1422,In_1471);
nor U328 (N_328,In_1005,In_1246);
and U329 (N_329,In_1162,In_647);
nor U330 (N_330,In_414,In_600);
xor U331 (N_331,In_1487,In_1145);
xnor U332 (N_332,In_827,In_1444);
nor U333 (N_333,In_26,In_1404);
xnor U334 (N_334,In_1035,In_1032);
and U335 (N_335,In_419,In_485);
or U336 (N_336,In_1296,In_197);
nor U337 (N_337,In_1336,In_6);
or U338 (N_338,In_793,In_229);
nor U339 (N_339,In_166,In_615);
xor U340 (N_340,In_199,In_711);
xor U341 (N_341,In_1155,In_1301);
xnor U342 (N_342,In_1225,In_220);
nand U343 (N_343,In_1012,In_1394);
nand U344 (N_344,In_1022,In_1219);
nor U345 (N_345,In_648,In_931);
xnor U346 (N_346,In_178,In_1070);
or U347 (N_347,In_343,In_974);
and U348 (N_348,In_1109,In_97);
and U349 (N_349,In_1318,In_972);
or U350 (N_350,In_117,In_397);
nor U351 (N_351,In_610,In_1390);
xor U352 (N_352,In_280,In_1306);
xor U353 (N_353,In_282,In_420);
nor U354 (N_354,In_948,In_593);
xnor U355 (N_355,In_704,In_1334);
and U356 (N_356,In_1199,In_740);
and U357 (N_357,In_351,In_1440);
nand U358 (N_358,In_549,In_724);
and U359 (N_359,In_17,In_1079);
nand U360 (N_360,In_161,In_127);
and U361 (N_361,In_1496,In_1249);
nand U362 (N_362,In_65,In_1130);
or U363 (N_363,In_1252,In_1195);
or U364 (N_364,In_1139,In_1352);
nand U365 (N_365,In_799,In_246);
and U366 (N_366,In_510,In_1313);
nand U367 (N_367,In_263,In_88);
and U368 (N_368,In_1365,In_1439);
and U369 (N_369,In_699,In_809);
or U370 (N_370,In_90,In_132);
nand U371 (N_371,In_1053,In_970);
or U372 (N_372,In_562,In_338);
and U373 (N_373,In_1372,In_408);
or U374 (N_374,In_254,In_572);
nand U375 (N_375,In_225,In_1290);
xnor U376 (N_376,In_1099,In_788);
nor U377 (N_377,In_944,In_887);
nor U378 (N_378,In_757,In_381);
or U379 (N_379,In_1097,In_1431);
nor U380 (N_380,In_264,In_82);
xor U381 (N_381,In_395,In_916);
and U382 (N_382,In_84,In_415);
xor U383 (N_383,In_398,In_422);
or U384 (N_384,In_1340,In_1259);
nor U385 (N_385,In_1411,In_929);
and U386 (N_386,In_778,In_1454);
nand U387 (N_387,In_752,In_853);
and U388 (N_388,In_601,In_1327);
nand U389 (N_389,In_144,In_323);
or U390 (N_390,In_989,In_763);
or U391 (N_391,In_608,In_1080);
nand U392 (N_392,In_59,In_1212);
and U393 (N_393,In_433,In_560);
nor U394 (N_394,In_869,In_584);
and U395 (N_395,In_436,In_1050);
and U396 (N_396,In_1265,In_181);
xor U397 (N_397,In_406,In_334);
or U398 (N_398,In_545,In_1052);
nand U399 (N_399,In_592,In_91);
xnor U400 (N_400,In_483,In_1445);
or U401 (N_401,In_490,In_293);
or U402 (N_402,In_1479,In_129);
xnor U403 (N_403,In_666,In_787);
and U404 (N_404,In_767,In_283);
and U405 (N_405,In_1456,In_963);
nand U406 (N_406,In_1267,In_112);
or U407 (N_407,In_1370,In_77);
nand U408 (N_408,In_789,In_556);
or U409 (N_409,In_1412,In_318);
xor U410 (N_410,In_1244,In_299);
and U411 (N_411,In_1307,In_95);
xnor U412 (N_412,In_862,In_987);
nand U413 (N_413,In_1492,In_538);
and U414 (N_414,In_1302,In_1056);
and U415 (N_415,In_743,In_692);
xnor U416 (N_416,In_769,In_847);
and U417 (N_417,In_260,In_1321);
and U418 (N_418,In_1316,In_495);
xnor U419 (N_419,In_998,In_250);
xnor U420 (N_420,In_1105,In_206);
nor U421 (N_421,In_1042,In_599);
or U422 (N_422,In_1176,In_850);
nor U423 (N_423,In_645,In_1120);
xor U424 (N_424,In_108,In_1426);
or U425 (N_425,In_1258,In_373);
or U426 (N_426,In_445,In_927);
nor U427 (N_427,In_1157,In_817);
or U428 (N_428,In_1046,In_507);
or U429 (N_429,In_1437,In_1115);
or U430 (N_430,In_964,In_535);
and U431 (N_431,In_453,In_832);
xnor U432 (N_432,In_288,In_1186);
and U433 (N_433,In_638,In_110);
nor U434 (N_434,In_531,In_1126);
and U435 (N_435,In_1121,In_798);
and U436 (N_436,In_1180,In_1366);
nand U437 (N_437,In_64,In_879);
nor U438 (N_438,In_74,In_543);
and U439 (N_439,In_523,In_897);
and U440 (N_440,In_347,In_153);
nor U441 (N_441,In_881,In_700);
nor U442 (N_442,In_332,In_605);
nor U443 (N_443,In_384,In_1054);
or U444 (N_444,In_573,In_1339);
and U445 (N_445,In_1369,In_1027);
or U446 (N_446,In_1493,In_1031);
and U447 (N_447,In_1429,In_1447);
or U448 (N_448,In_1441,In_705);
and U449 (N_449,In_842,In_379);
xor U450 (N_450,In_1380,In_578);
nand U451 (N_451,In_662,In_3);
xnor U452 (N_452,In_128,In_712);
xor U453 (N_453,In_873,In_1414);
nand U454 (N_454,In_992,In_261);
nor U455 (N_455,In_1272,In_410);
nand U456 (N_456,In_1124,In_1013);
xnor U457 (N_457,In_202,In_234);
xor U458 (N_458,In_1457,In_187);
xnor U459 (N_459,In_493,In_194);
and U460 (N_460,In_1096,In_1279);
and U461 (N_461,In_176,In_121);
or U462 (N_462,In_1245,In_1150);
and U463 (N_463,In_83,In_541);
xnor U464 (N_464,In_1026,In_731);
nor U465 (N_465,In_69,In_882);
nor U466 (N_466,In_215,In_889);
and U467 (N_467,In_1200,In_859);
or U468 (N_468,In_29,In_21);
or U469 (N_469,In_156,In_1274);
nor U470 (N_470,In_667,In_768);
or U471 (N_471,In_192,In_1354);
nand U472 (N_472,In_1238,In_1237);
and U473 (N_473,In_730,In_1011);
and U474 (N_474,In_760,In_164);
and U475 (N_475,In_911,In_141);
xor U476 (N_476,In_824,In_1023);
xnor U477 (N_477,In_779,In_1025);
or U478 (N_478,In_1329,In_857);
and U479 (N_479,In_838,In_1111);
nor U480 (N_480,In_1227,In_718);
nor U481 (N_481,In_830,In_520);
or U482 (N_482,In_1315,In_179);
nor U483 (N_483,In_407,In_727);
or U484 (N_484,In_1451,In_773);
or U485 (N_485,In_1392,In_1342);
and U486 (N_486,In_118,In_548);
nand U487 (N_487,In_1041,In_303);
and U488 (N_488,In_1127,In_401);
nand U489 (N_489,In_1311,In_822);
xnor U490 (N_490,In_748,In_298);
nor U491 (N_491,In_527,In_1181);
xor U492 (N_492,In_1418,In_678);
nand U493 (N_493,In_120,In_80);
nor U494 (N_494,In_471,In_967);
nand U495 (N_495,In_1103,In_528);
nor U496 (N_496,In_247,In_130);
nor U497 (N_497,In_1000,In_639);
or U498 (N_498,In_335,In_390);
or U499 (N_499,In_918,In_920);
xor U500 (N_500,In_461,In_163);
and U501 (N_501,In_143,In_1282);
nand U502 (N_502,In_759,In_62);
or U503 (N_503,In_242,In_1146);
nor U504 (N_504,In_235,In_290);
nor U505 (N_505,In_747,In_1462);
nor U506 (N_506,In_595,In_780);
nand U507 (N_507,In_874,In_1086);
nor U508 (N_508,In_848,In_852);
xor U509 (N_509,In_913,In_170);
xnor U510 (N_510,In_717,In_1175);
nand U511 (N_511,In_442,In_557);
and U512 (N_512,In_24,In_1196);
nor U513 (N_513,In_1160,In_1488);
xnor U514 (N_514,In_576,In_92);
or U515 (N_515,In_574,In_851);
xnor U516 (N_516,In_1270,In_184);
nor U517 (N_517,In_171,In_1442);
nor U518 (N_518,In_245,In_230);
or U519 (N_519,In_236,In_1474);
xnor U520 (N_520,In_72,In_55);
and U521 (N_521,In_877,In_659);
or U522 (N_522,In_924,In_182);
nor U523 (N_523,In_350,In_1345);
and U524 (N_524,In_741,In_907);
xnor U525 (N_525,In_286,In_70);
and U526 (N_526,In_1253,In_1395);
nor U527 (N_527,In_425,In_1458);
nor U528 (N_528,In_1047,In_138);
nand U529 (N_529,In_649,In_237);
or U530 (N_530,In_896,In_755);
nand U531 (N_531,In_671,In_579);
and U532 (N_532,In_539,In_221);
nand U533 (N_533,In_517,In_1326);
and U534 (N_534,In_1187,In_189);
nand U535 (N_535,In_372,In_1467);
nand U536 (N_536,In_1453,In_1416);
xor U537 (N_537,In_474,In_382);
and U538 (N_538,In_1459,In_966);
nor U539 (N_539,In_304,In_48);
xor U540 (N_540,In_279,In_1335);
or U541 (N_541,In_751,In_607);
or U542 (N_542,In_1170,In_691);
nor U543 (N_543,In_982,In_565);
or U544 (N_544,In_1277,In_363);
and U545 (N_545,In_317,In_188);
nor U546 (N_546,In_587,In_596);
xnor U547 (N_547,In_258,In_375);
or U548 (N_548,In_434,In_281);
nor U549 (N_549,In_1132,In_336);
and U550 (N_550,In_1357,In_385);
or U551 (N_551,In_1148,In_487);
xnor U552 (N_552,In_477,In_1135);
xnor U553 (N_553,In_744,In_598);
xnor U554 (N_554,In_653,In_1291);
nand U555 (N_555,In_1207,In_1295);
or U556 (N_556,In_625,In_337);
nor U557 (N_557,In_922,In_441);
or U558 (N_558,In_1076,In_126);
xnor U559 (N_559,In_435,In_1179);
and U560 (N_560,In_676,In_472);
nor U561 (N_561,In_68,In_152);
or U562 (N_562,In_89,In_482);
and U563 (N_563,In_555,In_1385);
and U564 (N_564,In_1273,In_41);
nand U565 (N_565,In_703,In_429);
nor U566 (N_566,In_762,In_796);
nor U567 (N_567,In_1305,In_695);
or U568 (N_568,In_1094,In_943);
and U569 (N_569,In_308,In_217);
xnor U570 (N_570,In_814,In_122);
and U571 (N_571,In_208,In_94);
nand U572 (N_572,In_1194,In_781);
and U573 (N_573,In_988,In_100);
or U574 (N_574,In_469,In_580);
and U575 (N_575,In_928,In_775);
xor U576 (N_576,In_1090,In_1243);
xnor U577 (N_577,In_672,In_932);
or U578 (N_578,In_770,In_204);
nor U579 (N_579,In_1185,In_1364);
nor U580 (N_580,In_567,In_1024);
nand U581 (N_581,In_1248,In_1044);
xnor U582 (N_582,In_1449,In_1303);
and U583 (N_583,In_1183,In_378);
nor U584 (N_584,In_13,In_1443);
nand U585 (N_585,In_888,In_1071);
nor U586 (N_586,In_1091,In_706);
nand U587 (N_587,In_1400,In_1491);
and U588 (N_588,In_801,In_18);
nor U589 (N_589,In_1117,In_1191);
or U590 (N_590,In_568,In_983);
nor U591 (N_591,In_1125,In_1338);
nor U592 (N_592,In_503,In_1159);
nand U593 (N_593,In_333,In_1331);
and U594 (N_594,In_1482,In_713);
and U595 (N_595,In_239,In_878);
or U596 (N_596,In_7,In_278);
and U597 (N_597,In_586,In_871);
nand U598 (N_598,In_224,In_1278);
nand U599 (N_599,In_315,In_1190);
nand U600 (N_600,In_46,In_305);
nor U601 (N_601,In_683,In_40);
nand U602 (N_602,In_1358,In_257);
and U603 (N_603,In_322,In_933);
nor U604 (N_604,In_1113,In_513);
nor U605 (N_605,In_301,In_330);
xnor U606 (N_606,In_243,In_698);
xnor U607 (N_607,In_93,In_1123);
and U608 (N_608,In_1006,In_1348);
nand U609 (N_609,In_939,In_1078);
nand U610 (N_610,In_1478,In_219);
xnor U611 (N_611,In_1332,In_20);
or U612 (N_612,In_15,In_710);
nand U613 (N_613,In_325,In_73);
nor U614 (N_614,In_133,In_361);
xor U615 (N_615,In_79,In_1484);
nor U616 (N_616,In_1448,In_295);
and U617 (N_617,In_626,In_447);
nor U618 (N_618,In_1231,In_266);
xnor U619 (N_619,In_771,In_443);
xor U620 (N_620,In_891,In_446);
xor U621 (N_621,In_1405,In_307);
nand U622 (N_622,In_56,In_357);
or U623 (N_623,In_868,In_915);
and U624 (N_624,In_604,In_1009);
xnor U625 (N_625,In_979,In_19);
and U626 (N_626,In_1213,In_890);
and U627 (N_627,In_677,In_22);
nand U628 (N_628,In_451,In_149);
nand U629 (N_629,In_402,In_345);
nand U630 (N_630,In_183,In_553);
or U631 (N_631,In_1468,In_837);
xnor U632 (N_632,In_1057,In_1264);
or U633 (N_633,In_628,In_1072);
or U634 (N_634,In_475,In_114);
nor U635 (N_635,In_321,In_620);
or U636 (N_636,In_1386,In_1215);
and U637 (N_637,In_1201,In_251);
or U638 (N_638,In_658,In_450);
and U639 (N_639,In_806,In_1198);
and U640 (N_640,In_476,In_999);
nor U641 (N_641,In_1067,In_324);
and U642 (N_642,In_1450,In_714);
or U643 (N_643,In_551,In_1021);
xnor U644 (N_644,In_1427,In_904);
or U645 (N_645,In_150,In_1346);
nand U646 (N_646,In_956,In_1377);
and U647 (N_647,In_518,In_1396);
or U648 (N_648,In_1033,In_109);
nand U649 (N_649,In_1161,In_508);
nor U650 (N_650,In_641,In_585);
or U651 (N_651,In_45,In_417);
xnor U652 (N_652,In_1255,In_532);
nor U653 (N_653,In_815,In_416);
nor U654 (N_654,In_758,In_353);
or U655 (N_655,In_1151,In_1489);
nand U656 (N_656,In_1374,In_521);
or U657 (N_657,In_252,In_10);
nor U658 (N_658,In_949,In_498);
or U659 (N_659,In_103,In_802);
nand U660 (N_660,In_191,In_355);
or U661 (N_661,In_1204,In_486);
nand U662 (N_662,In_1073,In_1398);
nand U663 (N_663,In_519,In_656);
nand U664 (N_664,In_1106,In_193);
xnor U665 (N_665,In_463,In_753);
xor U666 (N_666,In_884,In_855);
xor U667 (N_667,In_1298,In_319);
nand U668 (N_668,In_195,In_941);
nor U669 (N_669,In_965,In_137);
nand U670 (N_670,In_1470,In_393);
nand U671 (N_671,In_297,In_1323);
and U672 (N_672,In_207,In_276);
and U673 (N_673,In_439,In_582);
or U674 (N_674,In_456,In_54);
xnor U675 (N_675,In_1193,In_642);
xor U676 (N_676,In_1269,In_1276);
nand U677 (N_677,In_216,In_78);
nor U678 (N_678,In_861,In_134);
and U679 (N_679,In_391,In_627);
nor U680 (N_680,In_1498,In_0);
and U681 (N_681,In_1063,In_536);
nand U682 (N_682,In_651,In_777);
xnor U683 (N_683,In_500,In_151);
and U684 (N_684,In_135,In_1192);
nor U685 (N_685,In_516,In_750);
nand U686 (N_686,In_807,In_1399);
nand U687 (N_687,In_729,In_1283);
nor U688 (N_688,In_716,In_287);
nand U689 (N_689,In_1182,In_1112);
nand U690 (N_690,In_1037,In_1166);
and U691 (N_691,In_686,In_96);
nand U692 (N_692,In_86,In_1337);
or U693 (N_693,In_1218,In_37);
or U694 (N_694,In_1408,In_66);
nand U695 (N_695,In_231,In_1060);
and U696 (N_696,In_1100,In_902);
nor U697 (N_697,In_423,In_669);
nor U698 (N_698,In_1222,In_1128);
xnor U699 (N_699,In_501,In_1368);
nand U700 (N_700,In_496,In_494);
xor U701 (N_701,In_1266,In_636);
or U702 (N_702,In_154,In_180);
and U703 (N_703,In_411,In_366);
or U704 (N_704,In_1217,In_975);
and U705 (N_705,In_1209,In_1402);
and U706 (N_706,In_32,In_909);
xnor U707 (N_707,In_833,In_825);
xnor U708 (N_708,In_241,In_512);
and U709 (N_709,In_540,In_210);
and U710 (N_710,In_1034,In_1137);
and U711 (N_711,In_1438,In_635);
nand U712 (N_712,In_465,In_810);
xor U713 (N_713,In_1432,In_969);
and U714 (N_714,In_1168,In_1007);
or U715 (N_715,In_696,In_44);
or U716 (N_716,In_329,In_356);
and U717 (N_717,In_934,In_654);
nor U718 (N_718,In_430,In_1363);
xor U719 (N_719,In_791,In_942);
nand U720 (N_720,In_826,In_1420);
or U721 (N_721,In_8,In_1384);
nand U722 (N_722,In_1383,In_1028);
xor U723 (N_723,In_589,In_1460);
or U724 (N_724,In_1251,In_113);
xor U725 (N_725,In_1242,In_694);
nor U726 (N_726,In_342,In_739);
nor U727 (N_727,In_1406,In_544);
and U728 (N_728,In_488,In_30);
xnor U729 (N_729,In_991,In_968);
or U730 (N_730,In_209,In_1325);
and U731 (N_731,In_1285,In_459);
nor U732 (N_732,In_270,In_1280);
nor U733 (N_733,In_67,In_34);
or U734 (N_734,In_720,In_1114);
or U735 (N_735,In_358,In_509);
nand U736 (N_736,In_1156,In_702);
or U737 (N_737,In_1141,In_893);
nor U738 (N_738,In_828,In_1136);
nor U739 (N_739,In_413,In_233);
and U740 (N_740,In_173,In_831);
xnor U741 (N_741,In_1019,In_294);
xor U742 (N_742,In_316,In_1379);
xnor U743 (N_743,In_646,In_1143);
xnor U744 (N_744,In_159,In_1401);
xor U745 (N_745,In_470,In_529);
xnor U746 (N_746,In_661,In_923);
or U747 (N_747,In_866,In_63);
and U748 (N_748,In_1216,In_169);
and U749 (N_749,In_794,In_256);
nand U750 (N_750,In_444,In_1449);
nand U751 (N_751,In_1440,In_770);
or U752 (N_752,In_1249,In_553);
xnor U753 (N_753,In_1326,In_385);
nand U754 (N_754,In_731,In_624);
or U755 (N_755,In_319,In_1264);
or U756 (N_756,In_856,In_320);
and U757 (N_757,In_880,In_1265);
or U758 (N_758,In_1175,In_48);
nor U759 (N_759,In_837,In_428);
or U760 (N_760,In_1424,In_1468);
nor U761 (N_761,In_296,In_380);
xnor U762 (N_762,In_308,In_1323);
nor U763 (N_763,In_1369,In_912);
and U764 (N_764,In_750,In_1274);
nor U765 (N_765,In_985,In_873);
or U766 (N_766,In_927,In_843);
nor U767 (N_767,In_1144,In_909);
nor U768 (N_768,In_595,In_436);
xor U769 (N_769,In_267,In_376);
and U770 (N_770,In_1311,In_314);
xor U771 (N_771,In_552,In_2);
and U772 (N_772,In_686,In_195);
xnor U773 (N_773,In_165,In_1209);
and U774 (N_774,In_1397,In_749);
and U775 (N_775,In_947,In_622);
nor U776 (N_776,In_445,In_1060);
nor U777 (N_777,In_588,In_994);
nand U778 (N_778,In_193,In_570);
or U779 (N_779,In_285,In_1315);
nor U780 (N_780,In_1329,In_1321);
nand U781 (N_781,In_682,In_660);
nand U782 (N_782,In_953,In_1385);
xnor U783 (N_783,In_207,In_508);
nand U784 (N_784,In_930,In_232);
and U785 (N_785,In_905,In_1148);
and U786 (N_786,In_1237,In_68);
and U787 (N_787,In_1076,In_350);
nand U788 (N_788,In_195,In_1202);
or U789 (N_789,In_1362,In_388);
xnor U790 (N_790,In_1371,In_1357);
and U791 (N_791,In_346,In_983);
nor U792 (N_792,In_701,In_1395);
nand U793 (N_793,In_1478,In_917);
xor U794 (N_794,In_473,In_328);
or U795 (N_795,In_214,In_1205);
or U796 (N_796,In_842,In_1029);
nor U797 (N_797,In_1021,In_68);
or U798 (N_798,In_801,In_1181);
nor U799 (N_799,In_875,In_575);
xnor U800 (N_800,In_950,In_252);
xor U801 (N_801,In_165,In_727);
xnor U802 (N_802,In_941,In_1296);
xnor U803 (N_803,In_270,In_701);
nor U804 (N_804,In_1492,In_409);
and U805 (N_805,In_324,In_1223);
and U806 (N_806,In_513,In_660);
nor U807 (N_807,In_371,In_87);
and U808 (N_808,In_715,In_746);
nor U809 (N_809,In_1299,In_524);
and U810 (N_810,In_769,In_859);
nor U811 (N_811,In_672,In_395);
xor U812 (N_812,In_142,In_1052);
nand U813 (N_813,In_160,In_386);
xnor U814 (N_814,In_1434,In_811);
and U815 (N_815,In_1201,In_1400);
xnor U816 (N_816,In_720,In_593);
xor U817 (N_817,In_139,In_100);
nor U818 (N_818,In_1266,In_277);
nand U819 (N_819,In_346,In_1118);
nand U820 (N_820,In_159,In_1095);
nor U821 (N_821,In_1405,In_117);
xor U822 (N_822,In_1293,In_1199);
and U823 (N_823,In_141,In_776);
nand U824 (N_824,In_649,In_1408);
xnor U825 (N_825,In_972,In_1057);
nand U826 (N_826,In_1240,In_1122);
nand U827 (N_827,In_673,In_847);
nor U828 (N_828,In_410,In_1458);
nand U829 (N_829,In_838,In_946);
nor U830 (N_830,In_215,In_905);
xnor U831 (N_831,In_1054,In_587);
or U832 (N_832,In_65,In_438);
nor U833 (N_833,In_122,In_1128);
nor U834 (N_834,In_278,In_1435);
and U835 (N_835,In_1404,In_851);
or U836 (N_836,In_1093,In_723);
nand U837 (N_837,In_1067,In_1100);
nand U838 (N_838,In_805,In_1398);
xor U839 (N_839,In_1224,In_864);
or U840 (N_840,In_476,In_1453);
and U841 (N_841,In_1476,In_1253);
nor U842 (N_842,In_736,In_945);
and U843 (N_843,In_1198,In_921);
and U844 (N_844,In_936,In_638);
nand U845 (N_845,In_577,In_631);
nand U846 (N_846,In_887,In_1077);
or U847 (N_847,In_651,In_173);
nor U848 (N_848,In_900,In_461);
nand U849 (N_849,In_1358,In_1128);
or U850 (N_850,In_173,In_92);
nand U851 (N_851,In_1087,In_126);
nor U852 (N_852,In_1121,In_1430);
nand U853 (N_853,In_1151,In_193);
nand U854 (N_854,In_1189,In_637);
nand U855 (N_855,In_1011,In_1108);
xor U856 (N_856,In_1066,In_1077);
xnor U857 (N_857,In_1316,In_98);
xor U858 (N_858,In_1420,In_759);
or U859 (N_859,In_230,In_619);
and U860 (N_860,In_507,In_1375);
xor U861 (N_861,In_391,In_1397);
xor U862 (N_862,In_778,In_1278);
xnor U863 (N_863,In_1259,In_583);
xnor U864 (N_864,In_58,In_1286);
nor U865 (N_865,In_519,In_24);
xor U866 (N_866,In_1321,In_742);
or U867 (N_867,In_772,In_1189);
xnor U868 (N_868,In_613,In_1090);
xor U869 (N_869,In_159,In_224);
and U870 (N_870,In_1110,In_937);
or U871 (N_871,In_962,In_649);
and U872 (N_872,In_1128,In_288);
nand U873 (N_873,In_926,In_632);
nand U874 (N_874,In_1326,In_847);
nand U875 (N_875,In_1361,In_308);
or U876 (N_876,In_1280,In_823);
nand U877 (N_877,In_1343,In_1157);
and U878 (N_878,In_1307,In_803);
or U879 (N_879,In_128,In_1216);
and U880 (N_880,In_1068,In_1217);
nor U881 (N_881,In_836,In_348);
nand U882 (N_882,In_986,In_1143);
nor U883 (N_883,In_1233,In_902);
xnor U884 (N_884,In_550,In_247);
and U885 (N_885,In_365,In_114);
and U886 (N_886,In_207,In_1440);
and U887 (N_887,In_424,In_1434);
or U888 (N_888,In_931,In_741);
nand U889 (N_889,In_19,In_1025);
or U890 (N_890,In_1252,In_363);
and U891 (N_891,In_897,In_70);
and U892 (N_892,In_1081,In_361);
and U893 (N_893,In_541,In_207);
and U894 (N_894,In_903,In_168);
nand U895 (N_895,In_175,In_152);
xor U896 (N_896,In_36,In_1490);
and U897 (N_897,In_1174,In_1322);
nor U898 (N_898,In_1140,In_1335);
xnor U899 (N_899,In_93,In_522);
and U900 (N_900,In_360,In_830);
nor U901 (N_901,In_1198,In_1300);
or U902 (N_902,In_405,In_920);
nand U903 (N_903,In_1483,In_1486);
nand U904 (N_904,In_1347,In_1160);
nor U905 (N_905,In_308,In_27);
xor U906 (N_906,In_1228,In_854);
or U907 (N_907,In_263,In_570);
xnor U908 (N_908,In_230,In_1397);
xnor U909 (N_909,In_1121,In_1284);
xnor U910 (N_910,In_924,In_864);
xnor U911 (N_911,In_241,In_647);
xor U912 (N_912,In_690,In_104);
nand U913 (N_913,In_811,In_325);
xnor U914 (N_914,In_829,In_1489);
and U915 (N_915,In_425,In_75);
xor U916 (N_916,In_1027,In_226);
nor U917 (N_917,In_1145,In_921);
nor U918 (N_918,In_1424,In_1156);
or U919 (N_919,In_707,In_166);
or U920 (N_920,In_740,In_1476);
and U921 (N_921,In_339,In_443);
or U922 (N_922,In_963,In_536);
or U923 (N_923,In_300,In_623);
nand U924 (N_924,In_11,In_1165);
nand U925 (N_925,In_1188,In_326);
xor U926 (N_926,In_982,In_1183);
or U927 (N_927,In_805,In_942);
nand U928 (N_928,In_278,In_17);
nand U929 (N_929,In_1404,In_241);
nor U930 (N_930,In_1202,In_1373);
or U931 (N_931,In_950,In_246);
and U932 (N_932,In_222,In_668);
nor U933 (N_933,In_184,In_836);
nor U934 (N_934,In_429,In_1196);
nor U935 (N_935,In_506,In_1486);
nand U936 (N_936,In_613,In_1360);
and U937 (N_937,In_1371,In_177);
nand U938 (N_938,In_511,In_38);
or U939 (N_939,In_585,In_1260);
and U940 (N_940,In_660,In_306);
and U941 (N_941,In_225,In_1153);
nand U942 (N_942,In_222,In_163);
nand U943 (N_943,In_946,In_419);
nand U944 (N_944,In_299,In_1478);
nor U945 (N_945,In_1026,In_378);
xnor U946 (N_946,In_753,In_1218);
or U947 (N_947,In_348,In_842);
xnor U948 (N_948,In_27,In_1497);
or U949 (N_949,In_1358,In_1499);
or U950 (N_950,In_389,In_1281);
nor U951 (N_951,In_458,In_1181);
nor U952 (N_952,In_371,In_636);
and U953 (N_953,In_823,In_12);
or U954 (N_954,In_1401,In_1076);
nand U955 (N_955,In_1099,In_347);
nand U956 (N_956,In_874,In_798);
or U957 (N_957,In_397,In_622);
nand U958 (N_958,In_780,In_344);
xor U959 (N_959,In_1297,In_206);
or U960 (N_960,In_157,In_302);
nand U961 (N_961,In_1442,In_707);
and U962 (N_962,In_1315,In_342);
or U963 (N_963,In_196,In_1361);
and U964 (N_964,In_207,In_643);
nand U965 (N_965,In_892,In_653);
nor U966 (N_966,In_86,In_980);
and U967 (N_967,In_617,In_545);
nand U968 (N_968,In_139,In_1058);
and U969 (N_969,In_903,In_74);
xnor U970 (N_970,In_1122,In_1091);
and U971 (N_971,In_78,In_1143);
nand U972 (N_972,In_845,In_132);
xnor U973 (N_973,In_754,In_948);
xor U974 (N_974,In_1445,In_728);
and U975 (N_975,In_739,In_874);
or U976 (N_976,In_272,In_523);
xnor U977 (N_977,In_98,In_947);
nand U978 (N_978,In_1078,In_1448);
or U979 (N_979,In_249,In_1089);
nand U980 (N_980,In_223,In_92);
nor U981 (N_981,In_1462,In_875);
xor U982 (N_982,In_61,In_1126);
nor U983 (N_983,In_150,In_7);
or U984 (N_984,In_1137,In_1025);
nor U985 (N_985,In_531,In_1213);
and U986 (N_986,In_1070,In_312);
nor U987 (N_987,In_98,In_534);
or U988 (N_988,In_1124,In_1245);
nand U989 (N_989,In_1245,In_854);
or U990 (N_990,In_351,In_1226);
and U991 (N_991,In_338,In_24);
and U992 (N_992,In_135,In_392);
nor U993 (N_993,In_621,In_1134);
xnor U994 (N_994,In_161,In_499);
nand U995 (N_995,In_309,In_950);
and U996 (N_996,In_63,In_535);
nand U997 (N_997,In_649,In_223);
nand U998 (N_998,In_1477,In_427);
and U999 (N_999,In_605,In_1461);
and U1000 (N_1000,N_543,N_790);
or U1001 (N_1001,N_264,N_432);
nor U1002 (N_1002,N_791,N_254);
xnor U1003 (N_1003,N_525,N_121);
or U1004 (N_1004,N_492,N_125);
or U1005 (N_1005,N_721,N_192);
or U1006 (N_1006,N_953,N_648);
xnor U1007 (N_1007,N_72,N_100);
or U1008 (N_1008,N_684,N_956);
nor U1009 (N_1009,N_268,N_499);
or U1010 (N_1010,N_356,N_411);
xor U1011 (N_1011,N_282,N_448);
xor U1012 (N_1012,N_889,N_623);
and U1013 (N_1013,N_519,N_209);
nand U1014 (N_1014,N_145,N_115);
xnor U1015 (N_1015,N_428,N_248);
and U1016 (N_1016,N_688,N_417);
xnor U1017 (N_1017,N_250,N_224);
nor U1018 (N_1018,N_365,N_553);
xor U1019 (N_1019,N_620,N_157);
xor U1020 (N_1020,N_276,N_691);
or U1021 (N_1021,N_204,N_693);
or U1022 (N_1022,N_540,N_622);
xnor U1023 (N_1023,N_335,N_5);
nor U1024 (N_1024,N_490,N_886);
and U1025 (N_1025,N_781,N_300);
xor U1026 (N_1026,N_345,N_374);
nor U1027 (N_1027,N_109,N_778);
and U1028 (N_1028,N_975,N_487);
xor U1029 (N_1029,N_332,N_714);
xor U1030 (N_1030,N_632,N_615);
nand U1031 (N_1031,N_461,N_407);
or U1032 (N_1032,N_585,N_379);
nand U1033 (N_1033,N_116,N_1);
nand U1034 (N_1034,N_24,N_238);
nor U1035 (N_1035,N_59,N_677);
or U1036 (N_1036,N_851,N_415);
xnor U1037 (N_1037,N_274,N_304);
and U1038 (N_1038,N_748,N_245);
xor U1039 (N_1039,N_897,N_580);
and U1040 (N_1040,N_314,N_194);
nand U1041 (N_1041,N_243,N_172);
or U1042 (N_1042,N_844,N_211);
xor U1043 (N_1043,N_409,N_972);
nand U1044 (N_1044,N_770,N_497);
and U1045 (N_1045,N_366,N_846);
or U1046 (N_1046,N_315,N_261);
nor U1047 (N_1047,N_223,N_403);
nor U1048 (N_1048,N_813,N_960);
nand U1049 (N_1049,N_981,N_854);
nor U1050 (N_1050,N_539,N_431);
nand U1051 (N_1051,N_454,N_303);
and U1052 (N_1052,N_433,N_187);
nor U1053 (N_1053,N_361,N_692);
or U1054 (N_1054,N_970,N_289);
and U1055 (N_1055,N_910,N_530);
nand U1056 (N_1056,N_702,N_545);
and U1057 (N_1057,N_312,N_728);
nor U1058 (N_1058,N_594,N_616);
or U1059 (N_1059,N_232,N_437);
or U1060 (N_1060,N_579,N_932);
or U1061 (N_1061,N_32,N_91);
xnor U1062 (N_1062,N_869,N_52);
nand U1063 (N_1063,N_665,N_928);
and U1064 (N_1064,N_234,N_640);
and U1065 (N_1065,N_658,N_958);
nand U1066 (N_1066,N_440,N_607);
or U1067 (N_1067,N_506,N_763);
xor U1068 (N_1068,N_468,N_758);
nand U1069 (N_1069,N_220,N_200);
and U1070 (N_1070,N_871,N_504);
nand U1071 (N_1071,N_475,N_96);
and U1072 (N_1072,N_17,N_853);
nor U1073 (N_1073,N_759,N_55);
nor U1074 (N_1074,N_350,N_296);
and U1075 (N_1075,N_856,N_973);
xnor U1076 (N_1076,N_795,N_865);
and U1077 (N_1077,N_811,N_765);
xnor U1078 (N_1078,N_771,N_847);
and U1079 (N_1079,N_890,N_652);
and U1080 (N_1080,N_906,N_275);
xor U1081 (N_1081,N_228,N_617);
nor U1082 (N_1082,N_610,N_882);
and U1083 (N_1083,N_399,N_141);
nor U1084 (N_1084,N_36,N_788);
nand U1085 (N_1085,N_241,N_93);
or U1086 (N_1086,N_629,N_33);
or U1087 (N_1087,N_988,N_92);
and U1088 (N_1088,N_435,N_872);
or U1089 (N_1089,N_88,N_152);
nand U1090 (N_1090,N_782,N_239);
or U1091 (N_1091,N_775,N_406);
xor U1092 (N_1092,N_855,N_460);
nand U1093 (N_1093,N_573,N_785);
or U1094 (N_1094,N_820,N_196);
nand U1095 (N_1095,N_783,N_79);
or U1096 (N_1096,N_912,N_509);
and U1097 (N_1097,N_302,N_97);
xor U1098 (N_1098,N_687,N_602);
nand U1099 (N_1099,N_762,N_135);
nand U1100 (N_1100,N_259,N_462);
nand U1101 (N_1101,N_90,N_342);
nand U1102 (N_1102,N_829,N_438);
and U1103 (N_1103,N_705,N_575);
nor U1104 (N_1104,N_527,N_306);
nand U1105 (N_1105,N_707,N_595);
xor U1106 (N_1106,N_182,N_138);
nor U1107 (N_1107,N_309,N_458);
nand U1108 (N_1108,N_596,N_420);
and U1109 (N_1109,N_925,N_201);
nand U1110 (N_1110,N_439,N_959);
and U1111 (N_1111,N_15,N_840);
nand U1112 (N_1112,N_337,N_895);
nor U1113 (N_1113,N_733,N_246);
nand U1114 (N_1114,N_104,N_987);
nand U1115 (N_1115,N_689,N_621);
and U1116 (N_1116,N_747,N_133);
xnor U1117 (N_1117,N_47,N_471);
nand U1118 (N_1118,N_484,N_69);
and U1119 (N_1119,N_367,N_571);
xor U1120 (N_1120,N_681,N_292);
and U1121 (N_1121,N_568,N_107);
nor U1122 (N_1122,N_685,N_963);
nor U1123 (N_1123,N_249,N_908);
nand U1124 (N_1124,N_325,N_348);
nor U1125 (N_1125,N_344,N_741);
and U1126 (N_1126,N_850,N_515);
nor U1127 (N_1127,N_386,N_203);
and U1128 (N_1128,N_542,N_165);
and U1129 (N_1129,N_84,N_675);
and U1130 (N_1130,N_965,N_817);
and U1131 (N_1131,N_108,N_496);
xnor U1132 (N_1132,N_930,N_179);
or U1133 (N_1133,N_819,N_28);
xnor U1134 (N_1134,N_215,N_734);
nor U1135 (N_1135,N_944,N_118);
xnor U1136 (N_1136,N_801,N_10);
nor U1137 (N_1137,N_476,N_336);
and U1138 (N_1138,N_966,N_654);
and U1139 (N_1139,N_478,N_447);
nand U1140 (N_1140,N_551,N_393);
or U1141 (N_1141,N_646,N_395);
nor U1142 (N_1142,N_481,N_662);
nand U1143 (N_1143,N_74,N_311);
nand U1144 (N_1144,N_664,N_673);
or U1145 (N_1145,N_255,N_589);
nor U1146 (N_1146,N_552,N_848);
xnor U1147 (N_1147,N_922,N_301);
nand U1148 (N_1148,N_969,N_548);
nand U1149 (N_1149,N_230,N_559);
and U1150 (N_1150,N_500,N_993);
or U1151 (N_1151,N_700,N_387);
xnor U1152 (N_1152,N_166,N_140);
nor U1153 (N_1153,N_508,N_375);
or U1154 (N_1154,N_150,N_40);
nand U1155 (N_1155,N_666,N_147);
xnor U1156 (N_1156,N_208,N_597);
nor U1157 (N_1157,N_796,N_824);
nand U1158 (N_1158,N_180,N_892);
or U1159 (N_1159,N_715,N_523);
nand U1160 (N_1160,N_881,N_729);
xnor U1161 (N_1161,N_2,N_416);
and U1162 (N_1162,N_560,N_378);
nand U1163 (N_1163,N_43,N_326);
nand U1164 (N_1164,N_916,N_126);
and U1165 (N_1165,N_23,N_940);
xor U1166 (N_1166,N_213,N_308);
nand U1167 (N_1167,N_873,N_343);
xor U1168 (N_1168,N_8,N_441);
and U1169 (N_1169,N_739,N_352);
nor U1170 (N_1170,N_794,N_190);
nor U1171 (N_1171,N_831,N_643);
xnor U1172 (N_1172,N_710,N_544);
or U1173 (N_1173,N_199,N_793);
or U1174 (N_1174,N_372,N_974);
xnor U1175 (N_1175,N_113,N_631);
nor U1176 (N_1176,N_952,N_266);
nand U1177 (N_1177,N_547,N_430);
nand U1178 (N_1178,N_355,N_329);
nor U1179 (N_1179,N_449,N_880);
nor U1180 (N_1180,N_754,N_562);
and U1181 (N_1181,N_34,N_772);
nor U1182 (N_1182,N_584,N_732);
nor U1183 (N_1183,N_722,N_786);
nor U1184 (N_1184,N_26,N_672);
nand U1185 (N_1185,N_514,N_404);
and U1186 (N_1186,N_680,N_465);
nor U1187 (N_1187,N_893,N_608);
xor U1188 (N_1188,N_827,N_64);
xnor U1189 (N_1189,N_983,N_962);
or U1190 (N_1190,N_351,N_751);
and U1191 (N_1191,N_307,N_651);
nor U1192 (N_1192,N_735,N_491);
and U1193 (N_1193,N_334,N_679);
xnor U1194 (N_1194,N_270,N_900);
or U1195 (N_1195,N_236,N_272);
nor U1196 (N_1196,N_67,N_815);
or U1197 (N_1197,N_638,N_843);
or U1198 (N_1198,N_883,N_294);
or U1199 (N_1199,N_945,N_832);
xor U1200 (N_1200,N_434,N_359);
and U1201 (N_1201,N_980,N_875);
and U1202 (N_1202,N_671,N_927);
nor U1203 (N_1203,N_159,N_614);
xor U1204 (N_1204,N_968,N_653);
and U1205 (N_1205,N_0,N_590);
nor U1206 (N_1206,N_66,N_582);
or U1207 (N_1207,N_173,N_825);
or U1208 (N_1208,N_290,N_660);
nor U1209 (N_1209,N_736,N_124);
nand U1210 (N_1210,N_566,N_62);
xnor U1211 (N_1211,N_625,N_546);
xor U1212 (N_1212,N_647,N_798);
or U1213 (N_1213,N_512,N_368);
nand U1214 (N_1214,N_57,N_50);
xor U1215 (N_1215,N_915,N_792);
nand U1216 (N_1216,N_322,N_98);
or U1217 (N_1217,N_61,N_76);
or U1218 (N_1218,N_799,N_533);
nor U1219 (N_1219,N_857,N_907);
nand U1220 (N_1220,N_902,N_577);
nor U1221 (N_1221,N_456,N_740);
or U1222 (N_1222,N_839,N_841);
xor U1223 (N_1223,N_708,N_534);
and U1224 (N_1224,N_341,N_412);
nand U1225 (N_1225,N_737,N_178);
nor U1226 (N_1226,N_130,N_753);
and U1227 (N_1227,N_698,N_455);
nand U1228 (N_1228,N_425,N_174);
nor U1229 (N_1229,N_78,N_750);
or U1230 (N_1230,N_205,N_911);
or U1231 (N_1231,N_995,N_380);
or U1232 (N_1232,N_520,N_258);
nor U1233 (N_1233,N_929,N_526);
nor U1234 (N_1234,N_105,N_556);
or U1235 (N_1235,N_946,N_427);
xor U1236 (N_1236,N_233,N_68);
xnor U1237 (N_1237,N_936,N_943);
and U1238 (N_1238,N_273,N_717);
nand U1239 (N_1239,N_835,N_450);
nand U1240 (N_1240,N_44,N_567);
nor U1241 (N_1241,N_554,N_423);
nor U1242 (N_1242,N_485,N_752);
nor U1243 (N_1243,N_94,N_627);
or U1244 (N_1244,N_787,N_240);
and U1245 (N_1245,N_75,N_588);
nor U1246 (N_1246,N_634,N_466);
nor U1247 (N_1247,N_370,N_931);
nand U1248 (N_1248,N_802,N_516);
and U1249 (N_1249,N_637,N_557);
xnor U1250 (N_1250,N_469,N_726);
nor U1251 (N_1251,N_445,N_320);
and U1252 (N_1252,N_723,N_522);
and U1253 (N_1253,N_86,N_18);
nor U1254 (N_1254,N_400,N_939);
xnor U1255 (N_1255,N_413,N_776);
or U1256 (N_1256,N_253,N_99);
nand U1257 (N_1257,N_19,N_347);
nor U1258 (N_1258,N_202,N_175);
xor U1259 (N_1259,N_868,N_537);
and U1260 (N_1260,N_586,N_690);
xor U1261 (N_1261,N_132,N_587);
nor U1262 (N_1262,N_635,N_976);
nand U1263 (N_1263,N_967,N_926);
or U1264 (N_1264,N_918,N_369);
nor U1265 (N_1265,N_210,N_35);
nand U1266 (N_1266,N_129,N_593);
nand U1267 (N_1267,N_947,N_77);
nor U1268 (N_1268,N_446,N_821);
xnor U1269 (N_1269,N_473,N_191);
xor U1270 (N_1270,N_480,N_877);
xnor U1271 (N_1271,N_11,N_521);
nor U1272 (N_1272,N_826,N_859);
nor U1273 (N_1273,N_459,N_774);
xor U1274 (N_1274,N_382,N_316);
or U1275 (N_1275,N_498,N_299);
nand U1276 (N_1276,N_262,N_697);
nand U1277 (N_1277,N_661,N_574);
xor U1278 (N_1278,N_151,N_49);
nand U1279 (N_1279,N_331,N_295);
nor U1280 (N_1280,N_488,N_992);
nand U1281 (N_1281,N_950,N_764);
nand U1282 (N_1282,N_780,N_453);
nand U1283 (N_1283,N_961,N_444);
xor U1284 (N_1284,N_87,N_719);
nand U1285 (N_1285,N_878,N_879);
and U1286 (N_1286,N_624,N_267);
and U1287 (N_1287,N_618,N_720);
or U1288 (N_1288,N_168,N_206);
or U1289 (N_1289,N_749,N_106);
xnor U1290 (N_1290,N_221,N_467);
and U1291 (N_1291,N_866,N_58);
and U1292 (N_1292,N_169,N_163);
nand U1293 (N_1293,N_313,N_287);
nand U1294 (N_1294,N_20,N_701);
or U1295 (N_1295,N_373,N_807);
or U1296 (N_1296,N_251,N_513);
or U1297 (N_1297,N_102,N_442);
xor U1298 (N_1298,N_396,N_195);
xnor U1299 (N_1299,N_131,N_518);
and U1300 (N_1300,N_21,N_167);
xor U1301 (N_1301,N_153,N_110);
and U1302 (N_1302,N_860,N_392);
nor U1303 (N_1303,N_156,N_641);
or U1304 (N_1304,N_604,N_247);
or U1305 (N_1305,N_704,N_887);
or U1306 (N_1306,N_164,N_738);
nand U1307 (N_1307,N_128,N_838);
nor U1308 (N_1308,N_283,N_60);
xor U1309 (N_1309,N_894,N_402);
nand U1310 (N_1310,N_845,N_142);
xnor U1311 (N_1311,N_134,N_71);
nor U1312 (N_1312,N_991,N_612);
or U1313 (N_1313,N_123,N_111);
or U1314 (N_1314,N_127,N_193);
nand U1315 (N_1315,N_324,N_694);
or U1316 (N_1316,N_979,N_833);
and U1317 (N_1317,N_649,N_360);
nor U1318 (N_1318,N_605,N_531);
nand U1319 (N_1319,N_482,N_362);
or U1320 (N_1320,N_122,N_388);
xor U1321 (N_1321,N_184,N_176);
or U1322 (N_1322,N_421,N_528);
and U1323 (N_1323,N_898,N_330);
xor U1324 (N_1324,N_600,N_41);
xor U1325 (N_1325,N_609,N_933);
nor U1326 (N_1326,N_377,N_842);
xor U1327 (N_1327,N_212,N_14);
and U1328 (N_1328,N_30,N_381);
xor U1329 (N_1329,N_227,N_674);
or U1330 (N_1330,N_226,N_185);
xnor U1331 (N_1331,N_328,N_657);
or U1332 (N_1332,N_148,N_257);
or U1333 (N_1333,N_809,N_998);
or U1334 (N_1334,N_494,N_996);
nor U1335 (N_1335,N_999,N_570);
or U1336 (N_1336,N_598,N_565);
xor U1337 (N_1337,N_37,N_155);
nand U1338 (N_1338,N_864,N_921);
and U1339 (N_1339,N_564,N_278);
nand U1340 (N_1340,N_644,N_323);
nand U1341 (N_1341,N_80,N_712);
nand U1342 (N_1342,N_293,N_581);
or U1343 (N_1343,N_806,N_231);
nor U1344 (N_1344,N_744,N_112);
xnor U1345 (N_1345,N_538,N_663);
or U1346 (N_1346,N_834,N_464);
nor U1347 (N_1347,N_816,N_948);
xor U1348 (N_1348,N_884,N_746);
nand U1349 (N_1349,N_83,N_479);
or U1350 (N_1350,N_830,N_954);
nand U1351 (N_1351,N_891,N_12);
and U1352 (N_1352,N_477,N_867);
and U1353 (N_1353,N_683,N_310);
nor U1354 (N_1354,N_682,N_25);
xnor U1355 (N_1355,N_773,N_904);
and U1356 (N_1356,N_656,N_760);
nor U1357 (N_1357,N_288,N_22);
and U1358 (N_1358,N_63,N_924);
nand U1359 (N_1359,N_862,N_483);
or U1360 (N_1360,N_216,N_298);
xnor U1361 (N_1361,N_917,N_54);
and U1362 (N_1362,N_951,N_990);
nor U1363 (N_1363,N_463,N_376);
nand U1364 (N_1364,N_144,N_804);
nand U1365 (N_1365,N_13,N_899);
and U1366 (N_1366,N_810,N_572);
nand U1367 (N_1367,N_645,N_285);
nand U1368 (N_1368,N_286,N_655);
nor U1369 (N_1369,N_977,N_923);
nand U1370 (N_1370,N_162,N_507);
nor U1371 (N_1371,N_767,N_903);
xor U1372 (N_1372,N_628,N_452);
nor U1373 (N_1373,N_852,N_65);
nor U1374 (N_1374,N_822,N_158);
or U1375 (N_1375,N_909,N_457);
nor U1376 (N_1376,N_364,N_143);
xnor U1377 (N_1377,N_327,N_699);
nand U1378 (N_1378,N_919,N_994);
or U1379 (N_1379,N_474,N_170);
or U1380 (N_1380,N_235,N_858);
and U1381 (N_1381,N_743,N_529);
xnor U1382 (N_1382,N_385,N_139);
xor U1383 (N_1383,N_667,N_422);
or U1384 (N_1384,N_670,N_451);
nand U1385 (N_1385,N_384,N_363);
xor U1386 (N_1386,N_920,N_229);
nor U1387 (N_1387,N_934,N_219);
nor U1388 (N_1388,N_812,N_46);
nand U1389 (N_1389,N_354,N_742);
xnor U1390 (N_1390,N_524,N_284);
and U1391 (N_1391,N_89,N_837);
xor U1392 (N_1392,N_814,N_768);
nand U1393 (N_1393,N_414,N_70);
xnor U1394 (N_1394,N_136,N_561);
nor U1395 (N_1395,N_777,N_189);
or U1396 (N_1396,N_281,N_613);
nand U1397 (N_1397,N_731,N_42);
or U1398 (N_1398,N_935,N_755);
xor U1399 (N_1399,N_695,N_181);
and U1400 (N_1400,N_340,N_419);
and U1401 (N_1401,N_318,N_317);
nor U1402 (N_1402,N_319,N_885);
and U1403 (N_1403,N_45,N_103);
and U1404 (N_1404,N_601,N_730);
xor U1405 (N_1405,N_997,N_495);
nand U1406 (N_1406,N_177,N_676);
xor U1407 (N_1407,N_984,N_756);
nor U1408 (N_1408,N_727,N_630);
xor U1409 (N_1409,N_828,N_532);
xnor U1410 (N_1410,N_650,N_703);
and U1411 (N_1411,N_592,N_146);
or U1412 (N_1412,N_905,N_51);
and U1413 (N_1413,N_16,N_718);
nand U1414 (N_1414,N_263,N_279);
nand U1415 (N_1415,N_502,N_611);
nor U1416 (N_1416,N_53,N_160);
nor U1417 (N_1417,N_383,N_277);
nor U1418 (N_1418,N_686,N_297);
nand U1419 (N_1419,N_636,N_149);
nor U1420 (N_1420,N_603,N_510);
nor U1421 (N_1421,N_217,N_390);
nand U1422 (N_1422,N_823,N_619);
or U1423 (N_1423,N_985,N_222);
nor U1424 (N_1424,N_244,N_346);
xnor U1425 (N_1425,N_724,N_633);
nor U1426 (N_1426,N_7,N_349);
or U1427 (N_1427,N_511,N_321);
nor U1428 (N_1428,N_849,N_913);
or U1429 (N_1429,N_4,N_358);
xnor U1430 (N_1430,N_541,N_252);
nor U1431 (N_1431,N_3,N_563);
and U1432 (N_1432,N_576,N_38);
or U1433 (N_1433,N_642,N_265);
nand U1434 (N_1434,N_668,N_938);
xnor U1435 (N_1435,N_808,N_914);
nand U1436 (N_1436,N_218,N_766);
nand U1437 (N_1437,N_888,N_39);
xor U1438 (N_1438,N_874,N_408);
xor U1439 (N_1439,N_73,N_339);
and U1440 (N_1440,N_183,N_986);
nand U1441 (N_1441,N_949,N_599);
and U1442 (N_1442,N_443,N_410);
xnor U1443 (N_1443,N_493,N_501);
xnor U1444 (N_1444,N_558,N_357);
and U1445 (N_1445,N_535,N_797);
and U1446 (N_1446,N_260,N_725);
xor U1447 (N_1447,N_237,N_119);
or U1448 (N_1448,N_578,N_154);
nand U1449 (N_1449,N_333,N_81);
nor U1450 (N_1450,N_896,N_942);
nor U1451 (N_1451,N_418,N_669);
nand U1452 (N_1452,N_398,N_591);
or U1453 (N_1453,N_803,N_101);
nand U1454 (N_1454,N_9,N_555);
nor U1455 (N_1455,N_137,N_941);
nor U1456 (N_1456,N_517,N_186);
nor U1457 (N_1457,N_503,N_486);
or U1458 (N_1458,N_769,N_394);
nand U1459 (N_1459,N_716,N_626);
nand U1460 (N_1460,N_711,N_971);
nand U1461 (N_1461,N_569,N_391);
and U1462 (N_1462,N_120,N_955);
nand U1463 (N_1463,N_29,N_256);
and U1464 (N_1464,N_606,N_371);
and U1465 (N_1465,N_964,N_957);
nor U1466 (N_1466,N_757,N_405);
nor U1467 (N_1467,N_214,N_27);
or U1468 (N_1468,N_784,N_779);
nand U1469 (N_1469,N_436,N_805);
and U1470 (N_1470,N_305,N_280);
xor U1471 (N_1471,N_401,N_161);
xnor U1472 (N_1472,N_639,N_85);
nand U1473 (N_1473,N_225,N_863);
nand U1474 (N_1474,N_800,N_550);
nand U1475 (N_1475,N_82,N_114);
nand U1476 (N_1476,N_876,N_659);
nor U1477 (N_1477,N_271,N_117);
or U1478 (N_1478,N_745,N_470);
or U1479 (N_1479,N_549,N_583);
or U1480 (N_1480,N_48,N_761);
nor U1481 (N_1481,N_489,N_429);
nand U1482 (N_1482,N_197,N_818);
nand U1483 (N_1483,N_424,N_989);
and U1484 (N_1484,N_6,N_505);
and U1485 (N_1485,N_95,N_31);
xor U1486 (N_1486,N_269,N_171);
or U1487 (N_1487,N_198,N_426);
and U1488 (N_1488,N_678,N_937);
or U1489 (N_1489,N_242,N_706);
and U1490 (N_1490,N_713,N_696);
nor U1491 (N_1491,N_709,N_836);
and U1492 (N_1492,N_901,N_207);
nor U1493 (N_1493,N_789,N_353);
nor U1494 (N_1494,N_861,N_291);
or U1495 (N_1495,N_338,N_536);
xor U1496 (N_1496,N_188,N_978);
and U1497 (N_1497,N_870,N_56);
nand U1498 (N_1498,N_982,N_397);
nand U1499 (N_1499,N_472,N_389);
xnor U1500 (N_1500,N_35,N_406);
nand U1501 (N_1501,N_896,N_100);
nand U1502 (N_1502,N_323,N_310);
nor U1503 (N_1503,N_461,N_206);
and U1504 (N_1504,N_53,N_444);
nand U1505 (N_1505,N_330,N_113);
nand U1506 (N_1506,N_112,N_610);
nand U1507 (N_1507,N_51,N_237);
nor U1508 (N_1508,N_890,N_484);
nand U1509 (N_1509,N_225,N_470);
xor U1510 (N_1510,N_787,N_259);
nand U1511 (N_1511,N_446,N_263);
nand U1512 (N_1512,N_783,N_357);
nand U1513 (N_1513,N_655,N_291);
xor U1514 (N_1514,N_206,N_729);
nand U1515 (N_1515,N_75,N_186);
nor U1516 (N_1516,N_134,N_340);
xnor U1517 (N_1517,N_572,N_435);
xor U1518 (N_1518,N_932,N_912);
or U1519 (N_1519,N_601,N_542);
and U1520 (N_1520,N_723,N_502);
xnor U1521 (N_1521,N_668,N_936);
nor U1522 (N_1522,N_276,N_690);
nand U1523 (N_1523,N_714,N_359);
or U1524 (N_1524,N_766,N_436);
and U1525 (N_1525,N_544,N_859);
nand U1526 (N_1526,N_518,N_897);
nand U1527 (N_1527,N_472,N_453);
nor U1528 (N_1528,N_782,N_454);
or U1529 (N_1529,N_727,N_545);
xnor U1530 (N_1530,N_33,N_838);
xnor U1531 (N_1531,N_50,N_953);
nand U1532 (N_1532,N_429,N_620);
xnor U1533 (N_1533,N_824,N_569);
nor U1534 (N_1534,N_237,N_505);
nand U1535 (N_1535,N_684,N_114);
nor U1536 (N_1536,N_160,N_159);
and U1537 (N_1537,N_534,N_727);
xnor U1538 (N_1538,N_831,N_975);
nand U1539 (N_1539,N_745,N_381);
and U1540 (N_1540,N_662,N_819);
and U1541 (N_1541,N_851,N_663);
or U1542 (N_1542,N_487,N_397);
nor U1543 (N_1543,N_14,N_710);
and U1544 (N_1544,N_366,N_43);
xor U1545 (N_1545,N_643,N_226);
nand U1546 (N_1546,N_694,N_784);
nor U1547 (N_1547,N_61,N_602);
or U1548 (N_1548,N_861,N_205);
nand U1549 (N_1549,N_135,N_939);
nor U1550 (N_1550,N_142,N_160);
nand U1551 (N_1551,N_860,N_928);
xor U1552 (N_1552,N_215,N_296);
xnor U1553 (N_1553,N_689,N_750);
or U1554 (N_1554,N_760,N_160);
nor U1555 (N_1555,N_750,N_243);
xnor U1556 (N_1556,N_183,N_42);
nor U1557 (N_1557,N_648,N_36);
and U1558 (N_1558,N_177,N_62);
xor U1559 (N_1559,N_456,N_216);
nand U1560 (N_1560,N_619,N_195);
nand U1561 (N_1561,N_327,N_172);
or U1562 (N_1562,N_851,N_1);
nand U1563 (N_1563,N_773,N_448);
nor U1564 (N_1564,N_550,N_60);
xnor U1565 (N_1565,N_146,N_342);
or U1566 (N_1566,N_147,N_57);
xnor U1567 (N_1567,N_608,N_207);
or U1568 (N_1568,N_208,N_136);
xor U1569 (N_1569,N_787,N_923);
nor U1570 (N_1570,N_489,N_6);
and U1571 (N_1571,N_249,N_302);
nor U1572 (N_1572,N_948,N_2);
nand U1573 (N_1573,N_91,N_966);
or U1574 (N_1574,N_437,N_35);
or U1575 (N_1575,N_888,N_499);
and U1576 (N_1576,N_407,N_655);
or U1577 (N_1577,N_216,N_687);
xor U1578 (N_1578,N_372,N_659);
xnor U1579 (N_1579,N_755,N_24);
xnor U1580 (N_1580,N_619,N_243);
xnor U1581 (N_1581,N_411,N_796);
or U1582 (N_1582,N_131,N_157);
and U1583 (N_1583,N_500,N_962);
and U1584 (N_1584,N_520,N_460);
or U1585 (N_1585,N_192,N_848);
nor U1586 (N_1586,N_385,N_322);
and U1587 (N_1587,N_635,N_751);
xor U1588 (N_1588,N_688,N_264);
and U1589 (N_1589,N_122,N_301);
xor U1590 (N_1590,N_545,N_830);
or U1591 (N_1591,N_792,N_808);
nor U1592 (N_1592,N_284,N_279);
xor U1593 (N_1593,N_533,N_488);
xor U1594 (N_1594,N_954,N_186);
xor U1595 (N_1595,N_258,N_709);
or U1596 (N_1596,N_416,N_124);
xor U1597 (N_1597,N_879,N_592);
nand U1598 (N_1598,N_696,N_227);
or U1599 (N_1599,N_126,N_551);
nand U1600 (N_1600,N_654,N_836);
xor U1601 (N_1601,N_436,N_804);
nand U1602 (N_1602,N_397,N_311);
nand U1603 (N_1603,N_689,N_897);
and U1604 (N_1604,N_612,N_567);
or U1605 (N_1605,N_374,N_614);
nand U1606 (N_1606,N_221,N_446);
and U1607 (N_1607,N_75,N_610);
xnor U1608 (N_1608,N_772,N_587);
nand U1609 (N_1609,N_472,N_251);
or U1610 (N_1610,N_207,N_652);
or U1611 (N_1611,N_914,N_541);
nand U1612 (N_1612,N_919,N_591);
xor U1613 (N_1613,N_816,N_285);
nand U1614 (N_1614,N_433,N_945);
nor U1615 (N_1615,N_985,N_207);
and U1616 (N_1616,N_751,N_945);
nand U1617 (N_1617,N_323,N_474);
nand U1618 (N_1618,N_50,N_197);
xor U1619 (N_1619,N_801,N_8);
nor U1620 (N_1620,N_716,N_977);
xnor U1621 (N_1621,N_21,N_278);
and U1622 (N_1622,N_354,N_770);
xnor U1623 (N_1623,N_946,N_136);
nor U1624 (N_1624,N_240,N_644);
nor U1625 (N_1625,N_221,N_228);
or U1626 (N_1626,N_445,N_985);
xor U1627 (N_1627,N_764,N_570);
or U1628 (N_1628,N_457,N_436);
or U1629 (N_1629,N_354,N_888);
or U1630 (N_1630,N_746,N_45);
or U1631 (N_1631,N_786,N_233);
nand U1632 (N_1632,N_77,N_188);
nand U1633 (N_1633,N_442,N_707);
nor U1634 (N_1634,N_451,N_170);
xnor U1635 (N_1635,N_92,N_37);
or U1636 (N_1636,N_353,N_296);
nor U1637 (N_1637,N_823,N_363);
and U1638 (N_1638,N_748,N_781);
and U1639 (N_1639,N_456,N_370);
and U1640 (N_1640,N_66,N_32);
or U1641 (N_1641,N_517,N_886);
nor U1642 (N_1642,N_955,N_401);
and U1643 (N_1643,N_166,N_442);
or U1644 (N_1644,N_107,N_684);
nor U1645 (N_1645,N_49,N_910);
nor U1646 (N_1646,N_780,N_459);
and U1647 (N_1647,N_114,N_298);
xnor U1648 (N_1648,N_839,N_880);
nor U1649 (N_1649,N_347,N_76);
and U1650 (N_1650,N_399,N_414);
or U1651 (N_1651,N_572,N_76);
nand U1652 (N_1652,N_829,N_437);
nor U1653 (N_1653,N_499,N_326);
and U1654 (N_1654,N_90,N_813);
nand U1655 (N_1655,N_602,N_140);
nand U1656 (N_1656,N_926,N_902);
and U1657 (N_1657,N_570,N_358);
nand U1658 (N_1658,N_739,N_499);
nand U1659 (N_1659,N_180,N_478);
or U1660 (N_1660,N_487,N_202);
and U1661 (N_1661,N_799,N_506);
or U1662 (N_1662,N_905,N_467);
nand U1663 (N_1663,N_122,N_14);
nand U1664 (N_1664,N_643,N_412);
or U1665 (N_1665,N_688,N_49);
nor U1666 (N_1666,N_231,N_595);
nand U1667 (N_1667,N_615,N_801);
xnor U1668 (N_1668,N_19,N_318);
or U1669 (N_1669,N_782,N_810);
and U1670 (N_1670,N_104,N_985);
or U1671 (N_1671,N_986,N_291);
or U1672 (N_1672,N_406,N_502);
or U1673 (N_1673,N_10,N_856);
or U1674 (N_1674,N_683,N_376);
nand U1675 (N_1675,N_19,N_1);
or U1676 (N_1676,N_68,N_530);
nand U1677 (N_1677,N_546,N_381);
xnor U1678 (N_1678,N_561,N_139);
and U1679 (N_1679,N_225,N_79);
and U1680 (N_1680,N_243,N_83);
or U1681 (N_1681,N_786,N_967);
nand U1682 (N_1682,N_658,N_893);
and U1683 (N_1683,N_654,N_203);
and U1684 (N_1684,N_404,N_216);
nand U1685 (N_1685,N_47,N_381);
and U1686 (N_1686,N_737,N_447);
and U1687 (N_1687,N_449,N_870);
and U1688 (N_1688,N_386,N_562);
nand U1689 (N_1689,N_71,N_554);
nand U1690 (N_1690,N_701,N_297);
nor U1691 (N_1691,N_701,N_960);
or U1692 (N_1692,N_910,N_376);
nand U1693 (N_1693,N_122,N_318);
xnor U1694 (N_1694,N_486,N_828);
xnor U1695 (N_1695,N_104,N_126);
nor U1696 (N_1696,N_683,N_788);
xor U1697 (N_1697,N_558,N_309);
nor U1698 (N_1698,N_29,N_37);
nand U1699 (N_1699,N_162,N_790);
nand U1700 (N_1700,N_572,N_766);
and U1701 (N_1701,N_117,N_635);
nor U1702 (N_1702,N_50,N_128);
nand U1703 (N_1703,N_375,N_649);
nand U1704 (N_1704,N_160,N_6);
or U1705 (N_1705,N_128,N_718);
or U1706 (N_1706,N_503,N_826);
xnor U1707 (N_1707,N_52,N_101);
xor U1708 (N_1708,N_953,N_671);
nand U1709 (N_1709,N_809,N_385);
xnor U1710 (N_1710,N_960,N_904);
or U1711 (N_1711,N_237,N_838);
nor U1712 (N_1712,N_217,N_183);
nor U1713 (N_1713,N_861,N_276);
and U1714 (N_1714,N_234,N_116);
or U1715 (N_1715,N_790,N_625);
xnor U1716 (N_1716,N_145,N_958);
nor U1717 (N_1717,N_618,N_235);
nand U1718 (N_1718,N_828,N_886);
or U1719 (N_1719,N_71,N_829);
xnor U1720 (N_1720,N_370,N_197);
nand U1721 (N_1721,N_597,N_617);
or U1722 (N_1722,N_921,N_645);
or U1723 (N_1723,N_95,N_958);
and U1724 (N_1724,N_265,N_854);
or U1725 (N_1725,N_721,N_460);
and U1726 (N_1726,N_35,N_281);
or U1727 (N_1727,N_245,N_182);
xnor U1728 (N_1728,N_214,N_386);
nand U1729 (N_1729,N_975,N_7);
or U1730 (N_1730,N_587,N_651);
nor U1731 (N_1731,N_225,N_835);
and U1732 (N_1732,N_324,N_38);
xor U1733 (N_1733,N_558,N_498);
nand U1734 (N_1734,N_652,N_658);
nor U1735 (N_1735,N_207,N_822);
xor U1736 (N_1736,N_388,N_564);
nor U1737 (N_1737,N_297,N_724);
and U1738 (N_1738,N_31,N_415);
and U1739 (N_1739,N_996,N_560);
nand U1740 (N_1740,N_563,N_700);
and U1741 (N_1741,N_766,N_516);
or U1742 (N_1742,N_88,N_520);
nor U1743 (N_1743,N_421,N_939);
nand U1744 (N_1744,N_840,N_557);
nor U1745 (N_1745,N_777,N_4);
and U1746 (N_1746,N_103,N_198);
or U1747 (N_1747,N_620,N_948);
or U1748 (N_1748,N_878,N_378);
and U1749 (N_1749,N_39,N_71);
xnor U1750 (N_1750,N_250,N_251);
or U1751 (N_1751,N_927,N_229);
xnor U1752 (N_1752,N_271,N_940);
or U1753 (N_1753,N_461,N_252);
or U1754 (N_1754,N_610,N_324);
nand U1755 (N_1755,N_32,N_306);
nand U1756 (N_1756,N_385,N_719);
nor U1757 (N_1757,N_951,N_556);
and U1758 (N_1758,N_350,N_825);
xnor U1759 (N_1759,N_915,N_371);
or U1760 (N_1760,N_167,N_385);
xor U1761 (N_1761,N_738,N_92);
nor U1762 (N_1762,N_606,N_882);
and U1763 (N_1763,N_619,N_626);
nand U1764 (N_1764,N_222,N_864);
and U1765 (N_1765,N_47,N_55);
xnor U1766 (N_1766,N_724,N_693);
nor U1767 (N_1767,N_598,N_726);
xor U1768 (N_1768,N_400,N_545);
xnor U1769 (N_1769,N_110,N_486);
and U1770 (N_1770,N_137,N_639);
nand U1771 (N_1771,N_521,N_594);
and U1772 (N_1772,N_854,N_837);
or U1773 (N_1773,N_47,N_404);
xnor U1774 (N_1774,N_313,N_452);
and U1775 (N_1775,N_931,N_764);
nor U1776 (N_1776,N_608,N_297);
or U1777 (N_1777,N_322,N_277);
nor U1778 (N_1778,N_378,N_680);
nor U1779 (N_1779,N_801,N_700);
nand U1780 (N_1780,N_733,N_539);
nand U1781 (N_1781,N_440,N_770);
nand U1782 (N_1782,N_916,N_670);
xnor U1783 (N_1783,N_876,N_730);
xor U1784 (N_1784,N_818,N_81);
nand U1785 (N_1785,N_304,N_652);
nand U1786 (N_1786,N_498,N_670);
nand U1787 (N_1787,N_518,N_704);
nand U1788 (N_1788,N_58,N_811);
nor U1789 (N_1789,N_90,N_276);
xor U1790 (N_1790,N_421,N_213);
xor U1791 (N_1791,N_251,N_951);
xor U1792 (N_1792,N_94,N_799);
nand U1793 (N_1793,N_814,N_145);
nand U1794 (N_1794,N_594,N_554);
nor U1795 (N_1795,N_382,N_76);
nand U1796 (N_1796,N_515,N_275);
nor U1797 (N_1797,N_906,N_954);
nand U1798 (N_1798,N_842,N_87);
xor U1799 (N_1799,N_262,N_875);
and U1800 (N_1800,N_414,N_592);
nand U1801 (N_1801,N_442,N_787);
and U1802 (N_1802,N_355,N_704);
or U1803 (N_1803,N_370,N_528);
or U1804 (N_1804,N_147,N_190);
xor U1805 (N_1805,N_638,N_954);
nor U1806 (N_1806,N_458,N_350);
xnor U1807 (N_1807,N_467,N_862);
and U1808 (N_1808,N_643,N_119);
or U1809 (N_1809,N_856,N_611);
xor U1810 (N_1810,N_421,N_289);
and U1811 (N_1811,N_92,N_414);
nor U1812 (N_1812,N_238,N_618);
and U1813 (N_1813,N_798,N_222);
nor U1814 (N_1814,N_313,N_484);
nand U1815 (N_1815,N_356,N_612);
and U1816 (N_1816,N_318,N_117);
nand U1817 (N_1817,N_259,N_27);
and U1818 (N_1818,N_157,N_154);
and U1819 (N_1819,N_801,N_424);
xnor U1820 (N_1820,N_921,N_115);
or U1821 (N_1821,N_191,N_108);
or U1822 (N_1822,N_720,N_401);
nor U1823 (N_1823,N_790,N_399);
or U1824 (N_1824,N_622,N_569);
or U1825 (N_1825,N_880,N_388);
or U1826 (N_1826,N_474,N_479);
nor U1827 (N_1827,N_158,N_128);
and U1828 (N_1828,N_119,N_985);
or U1829 (N_1829,N_822,N_662);
nor U1830 (N_1830,N_765,N_660);
nand U1831 (N_1831,N_33,N_209);
nor U1832 (N_1832,N_481,N_982);
or U1833 (N_1833,N_771,N_595);
or U1834 (N_1834,N_672,N_240);
nand U1835 (N_1835,N_904,N_148);
nand U1836 (N_1836,N_52,N_878);
xnor U1837 (N_1837,N_198,N_151);
nand U1838 (N_1838,N_976,N_654);
or U1839 (N_1839,N_201,N_376);
and U1840 (N_1840,N_0,N_723);
and U1841 (N_1841,N_131,N_185);
nand U1842 (N_1842,N_523,N_890);
and U1843 (N_1843,N_381,N_727);
and U1844 (N_1844,N_914,N_419);
nor U1845 (N_1845,N_868,N_932);
xor U1846 (N_1846,N_596,N_570);
nor U1847 (N_1847,N_929,N_721);
nand U1848 (N_1848,N_939,N_614);
xor U1849 (N_1849,N_49,N_91);
nand U1850 (N_1850,N_70,N_494);
nand U1851 (N_1851,N_610,N_179);
nor U1852 (N_1852,N_622,N_680);
or U1853 (N_1853,N_502,N_776);
nand U1854 (N_1854,N_862,N_308);
nor U1855 (N_1855,N_483,N_758);
xor U1856 (N_1856,N_803,N_184);
and U1857 (N_1857,N_519,N_435);
and U1858 (N_1858,N_606,N_289);
nor U1859 (N_1859,N_656,N_349);
nand U1860 (N_1860,N_158,N_531);
nand U1861 (N_1861,N_608,N_288);
nor U1862 (N_1862,N_912,N_456);
xnor U1863 (N_1863,N_863,N_993);
or U1864 (N_1864,N_600,N_520);
nor U1865 (N_1865,N_828,N_294);
and U1866 (N_1866,N_298,N_10);
and U1867 (N_1867,N_318,N_661);
nor U1868 (N_1868,N_426,N_919);
xnor U1869 (N_1869,N_145,N_949);
nand U1870 (N_1870,N_284,N_482);
xor U1871 (N_1871,N_819,N_719);
xor U1872 (N_1872,N_731,N_222);
and U1873 (N_1873,N_257,N_222);
and U1874 (N_1874,N_566,N_939);
xnor U1875 (N_1875,N_176,N_533);
xnor U1876 (N_1876,N_683,N_638);
nor U1877 (N_1877,N_777,N_556);
and U1878 (N_1878,N_107,N_147);
or U1879 (N_1879,N_260,N_436);
nor U1880 (N_1880,N_302,N_994);
nand U1881 (N_1881,N_230,N_844);
nor U1882 (N_1882,N_116,N_149);
nand U1883 (N_1883,N_401,N_148);
xnor U1884 (N_1884,N_638,N_996);
and U1885 (N_1885,N_695,N_718);
xor U1886 (N_1886,N_482,N_780);
nor U1887 (N_1887,N_120,N_237);
and U1888 (N_1888,N_833,N_918);
or U1889 (N_1889,N_130,N_41);
xor U1890 (N_1890,N_190,N_449);
nand U1891 (N_1891,N_307,N_73);
and U1892 (N_1892,N_180,N_67);
and U1893 (N_1893,N_782,N_276);
or U1894 (N_1894,N_772,N_911);
and U1895 (N_1895,N_10,N_13);
xor U1896 (N_1896,N_977,N_396);
nor U1897 (N_1897,N_417,N_775);
and U1898 (N_1898,N_516,N_474);
nor U1899 (N_1899,N_690,N_710);
nor U1900 (N_1900,N_802,N_815);
nor U1901 (N_1901,N_662,N_912);
nand U1902 (N_1902,N_668,N_137);
nand U1903 (N_1903,N_323,N_324);
nand U1904 (N_1904,N_206,N_662);
nor U1905 (N_1905,N_829,N_359);
nand U1906 (N_1906,N_872,N_425);
nand U1907 (N_1907,N_266,N_869);
xnor U1908 (N_1908,N_198,N_165);
nor U1909 (N_1909,N_27,N_394);
or U1910 (N_1910,N_114,N_528);
or U1911 (N_1911,N_936,N_900);
or U1912 (N_1912,N_285,N_778);
nand U1913 (N_1913,N_498,N_575);
nor U1914 (N_1914,N_580,N_975);
xnor U1915 (N_1915,N_228,N_234);
or U1916 (N_1916,N_630,N_573);
nor U1917 (N_1917,N_517,N_190);
xor U1918 (N_1918,N_718,N_386);
or U1919 (N_1919,N_215,N_60);
nor U1920 (N_1920,N_348,N_548);
xor U1921 (N_1921,N_791,N_332);
nand U1922 (N_1922,N_898,N_54);
or U1923 (N_1923,N_154,N_600);
or U1924 (N_1924,N_112,N_932);
nand U1925 (N_1925,N_721,N_248);
and U1926 (N_1926,N_555,N_44);
nor U1927 (N_1927,N_333,N_245);
xnor U1928 (N_1928,N_992,N_812);
xnor U1929 (N_1929,N_90,N_319);
nand U1930 (N_1930,N_473,N_773);
or U1931 (N_1931,N_913,N_890);
and U1932 (N_1932,N_453,N_128);
nand U1933 (N_1933,N_865,N_926);
xor U1934 (N_1934,N_683,N_985);
nand U1935 (N_1935,N_686,N_465);
and U1936 (N_1936,N_902,N_220);
nand U1937 (N_1937,N_483,N_304);
nand U1938 (N_1938,N_543,N_972);
or U1939 (N_1939,N_49,N_231);
and U1940 (N_1940,N_714,N_476);
nand U1941 (N_1941,N_259,N_486);
nor U1942 (N_1942,N_173,N_574);
nor U1943 (N_1943,N_120,N_747);
or U1944 (N_1944,N_518,N_66);
xnor U1945 (N_1945,N_229,N_2);
or U1946 (N_1946,N_502,N_378);
and U1947 (N_1947,N_147,N_298);
and U1948 (N_1948,N_468,N_604);
or U1949 (N_1949,N_199,N_575);
nand U1950 (N_1950,N_767,N_946);
nand U1951 (N_1951,N_54,N_340);
or U1952 (N_1952,N_755,N_155);
nand U1953 (N_1953,N_773,N_820);
nor U1954 (N_1954,N_443,N_294);
and U1955 (N_1955,N_307,N_936);
xnor U1956 (N_1956,N_642,N_985);
nor U1957 (N_1957,N_298,N_234);
and U1958 (N_1958,N_614,N_862);
nor U1959 (N_1959,N_257,N_638);
xor U1960 (N_1960,N_562,N_614);
xor U1961 (N_1961,N_444,N_422);
and U1962 (N_1962,N_37,N_279);
or U1963 (N_1963,N_845,N_104);
nor U1964 (N_1964,N_515,N_547);
xor U1965 (N_1965,N_209,N_597);
nor U1966 (N_1966,N_208,N_509);
xor U1967 (N_1967,N_110,N_483);
or U1968 (N_1968,N_373,N_174);
nand U1969 (N_1969,N_309,N_382);
and U1970 (N_1970,N_183,N_613);
nand U1971 (N_1971,N_449,N_719);
nand U1972 (N_1972,N_656,N_97);
and U1973 (N_1973,N_64,N_18);
and U1974 (N_1974,N_712,N_826);
and U1975 (N_1975,N_598,N_186);
nor U1976 (N_1976,N_283,N_102);
nand U1977 (N_1977,N_665,N_520);
and U1978 (N_1978,N_733,N_409);
xor U1979 (N_1979,N_583,N_881);
nor U1980 (N_1980,N_988,N_421);
or U1981 (N_1981,N_820,N_781);
nor U1982 (N_1982,N_790,N_756);
or U1983 (N_1983,N_245,N_632);
or U1984 (N_1984,N_842,N_788);
xnor U1985 (N_1985,N_132,N_654);
xor U1986 (N_1986,N_43,N_522);
xnor U1987 (N_1987,N_779,N_656);
nand U1988 (N_1988,N_428,N_756);
nor U1989 (N_1989,N_193,N_521);
xor U1990 (N_1990,N_539,N_323);
and U1991 (N_1991,N_931,N_116);
and U1992 (N_1992,N_517,N_438);
or U1993 (N_1993,N_435,N_411);
xnor U1994 (N_1994,N_356,N_83);
and U1995 (N_1995,N_787,N_742);
nor U1996 (N_1996,N_956,N_177);
and U1997 (N_1997,N_483,N_305);
xnor U1998 (N_1998,N_111,N_810);
nand U1999 (N_1999,N_947,N_930);
nor U2000 (N_2000,N_1382,N_1214);
or U2001 (N_2001,N_1275,N_1208);
xnor U2002 (N_2002,N_1190,N_1433);
xor U2003 (N_2003,N_1745,N_1731);
and U2004 (N_2004,N_1762,N_1060);
or U2005 (N_2005,N_1933,N_1193);
nand U2006 (N_2006,N_1801,N_1141);
xnor U2007 (N_2007,N_1550,N_1901);
xor U2008 (N_2008,N_1918,N_1029);
or U2009 (N_2009,N_1604,N_1172);
nor U2010 (N_2010,N_1832,N_1635);
nor U2011 (N_2011,N_1370,N_1578);
nor U2012 (N_2012,N_1870,N_1000);
nand U2013 (N_2013,N_1508,N_1676);
nand U2014 (N_2014,N_1037,N_1450);
xor U2015 (N_2015,N_1605,N_1129);
nand U2016 (N_2016,N_1943,N_1534);
nand U2017 (N_2017,N_1634,N_1632);
and U2018 (N_2018,N_1527,N_1880);
xnor U2019 (N_2019,N_1455,N_1505);
nand U2020 (N_2020,N_1182,N_1102);
nand U2021 (N_2021,N_1706,N_1893);
xor U2022 (N_2022,N_1445,N_1813);
xor U2023 (N_2023,N_1669,N_1916);
and U2024 (N_2024,N_1337,N_1197);
nor U2025 (N_2025,N_1216,N_1793);
and U2026 (N_2026,N_1758,N_1617);
or U2027 (N_2027,N_1059,N_1820);
nand U2028 (N_2028,N_1904,N_1816);
nor U2029 (N_2029,N_1046,N_1392);
nand U2030 (N_2030,N_1856,N_1618);
and U2031 (N_2031,N_1951,N_1664);
xor U2032 (N_2032,N_1448,N_1308);
xnor U2033 (N_2033,N_1369,N_1792);
nor U2034 (N_2034,N_1571,N_1311);
nand U2035 (N_2035,N_1285,N_1969);
and U2036 (N_2036,N_1101,N_1986);
or U2037 (N_2037,N_1939,N_1887);
and U2038 (N_2038,N_1688,N_1614);
or U2039 (N_2039,N_1021,N_1325);
xnor U2040 (N_2040,N_1631,N_1707);
nor U2041 (N_2041,N_1967,N_1388);
and U2042 (N_2042,N_1122,N_1406);
xor U2043 (N_2043,N_1068,N_1695);
or U2044 (N_2044,N_1858,N_1401);
or U2045 (N_2045,N_1373,N_1464);
and U2046 (N_2046,N_1948,N_1767);
or U2047 (N_2047,N_1850,N_1330);
nor U2048 (N_2048,N_1211,N_1553);
nor U2049 (N_2049,N_1570,N_1541);
xnor U2050 (N_2050,N_1528,N_1278);
and U2051 (N_2051,N_1081,N_1807);
nand U2052 (N_2052,N_1657,N_1804);
nor U2053 (N_2053,N_1746,N_1394);
nor U2054 (N_2054,N_1867,N_1425);
xnor U2055 (N_2055,N_1023,N_1449);
nand U2056 (N_2056,N_1339,N_1823);
and U2057 (N_2057,N_1261,N_1366);
xor U2058 (N_2058,N_1775,N_1935);
or U2059 (N_2059,N_1824,N_1321);
and U2060 (N_2060,N_1010,N_1420);
and U2061 (N_2061,N_1130,N_1032);
and U2062 (N_2062,N_1502,N_1266);
xor U2063 (N_2063,N_1902,N_1350);
or U2064 (N_2064,N_1964,N_1298);
xor U2065 (N_2065,N_1223,N_1552);
xnor U2066 (N_2066,N_1472,N_1621);
nor U2067 (N_2067,N_1545,N_1761);
nor U2068 (N_2068,N_1771,N_1312);
xor U2069 (N_2069,N_1763,N_1929);
or U2070 (N_2070,N_1993,N_1728);
or U2071 (N_2071,N_1280,N_1682);
nand U2072 (N_2072,N_1999,N_1753);
nor U2073 (N_2073,N_1555,N_1778);
and U2074 (N_2074,N_1187,N_1334);
and U2075 (N_2075,N_1093,N_1825);
nor U2076 (N_2076,N_1355,N_1959);
nor U2077 (N_2077,N_1599,N_1191);
or U2078 (N_2078,N_1096,N_1517);
and U2079 (N_2079,N_1720,N_1784);
and U2080 (N_2080,N_1205,N_1836);
or U2081 (N_2081,N_1594,N_1882);
xor U2082 (N_2082,N_1936,N_1646);
nand U2083 (N_2083,N_1700,N_1254);
or U2084 (N_2084,N_1227,N_1252);
nand U2085 (N_2085,N_1041,N_1466);
or U2086 (N_2086,N_1835,N_1259);
and U2087 (N_2087,N_1347,N_1241);
nor U2088 (N_2088,N_1297,N_1198);
nand U2089 (N_2089,N_1219,N_1760);
nor U2090 (N_2090,N_1245,N_1195);
or U2091 (N_2091,N_1301,N_1158);
xor U2092 (N_2092,N_1487,N_1846);
xor U2093 (N_2093,N_1616,N_1884);
or U2094 (N_2094,N_1381,N_1317);
or U2095 (N_2095,N_1643,N_1495);
xnor U2096 (N_2096,N_1652,N_1611);
xor U2097 (N_2097,N_1708,N_1623);
nand U2098 (N_2098,N_1100,N_1459);
nand U2099 (N_2099,N_1210,N_1496);
and U2100 (N_2100,N_1307,N_1180);
xnor U2101 (N_2101,N_1989,N_1670);
xnor U2102 (N_2102,N_1480,N_1869);
xnor U2103 (N_2103,N_1583,N_1966);
xnor U2104 (N_2104,N_1145,N_1136);
nor U2105 (N_2105,N_1351,N_1926);
nand U2106 (N_2106,N_1209,N_1659);
xor U2107 (N_2107,N_1713,N_1465);
nor U2108 (N_2108,N_1542,N_1803);
and U2109 (N_2109,N_1300,N_1976);
or U2110 (N_2110,N_1919,N_1019);
xnor U2111 (N_2111,N_1460,N_1645);
and U2112 (N_2112,N_1769,N_1133);
nor U2113 (N_2113,N_1403,N_1033);
nand U2114 (N_2114,N_1743,N_1680);
and U2115 (N_2115,N_1162,N_1538);
nor U2116 (N_2116,N_1173,N_1353);
or U2117 (N_2117,N_1446,N_1927);
nand U2118 (N_2118,N_1485,N_1957);
xnor U2119 (N_2119,N_1977,N_1685);
or U2120 (N_2120,N_1013,N_1965);
xor U2121 (N_2121,N_1015,N_1510);
and U2122 (N_2122,N_1315,N_1636);
xnor U2123 (N_2123,N_1609,N_1426);
nor U2124 (N_2124,N_1886,N_1383);
nand U2125 (N_2125,N_1112,N_1547);
nand U2126 (N_2126,N_1672,N_1045);
nand U2127 (N_2127,N_1126,N_1110);
nand U2128 (N_2128,N_1949,N_1452);
nand U2129 (N_2129,N_1106,N_1717);
and U2130 (N_2130,N_1196,N_1954);
or U2131 (N_2131,N_1386,N_1437);
nand U2132 (N_2132,N_1387,N_1840);
xnor U2133 (N_2133,N_1267,N_1741);
and U2134 (N_2134,N_1549,N_1482);
and U2135 (N_2135,N_1170,N_1932);
xnor U2136 (N_2136,N_1090,N_1722);
nand U2137 (N_2137,N_1828,N_1078);
nand U2138 (N_2138,N_1584,N_1883);
or U2139 (N_2139,N_1212,N_1735);
and U2140 (N_2140,N_1087,N_1585);
nand U2141 (N_2141,N_1475,N_1814);
xor U2142 (N_2142,N_1498,N_1593);
nand U2143 (N_2143,N_1247,N_1917);
and U2144 (N_2144,N_1027,N_1898);
nand U2145 (N_2145,N_1503,N_1303);
and U2146 (N_2146,N_1432,N_1914);
or U2147 (N_2147,N_1159,N_1513);
and U2148 (N_2148,N_1730,N_1515);
xnor U2149 (N_2149,N_1233,N_1716);
xnor U2150 (N_2150,N_1451,N_1907);
nor U2151 (N_2151,N_1218,N_1001);
and U2152 (N_2152,N_1567,N_1625);
xor U2153 (N_2153,N_1668,N_1915);
or U2154 (N_2154,N_1160,N_1895);
nand U2155 (N_2155,N_1866,N_1782);
nand U2156 (N_2156,N_1074,N_1596);
or U2157 (N_2157,N_1072,N_1759);
and U2158 (N_2158,N_1613,N_1615);
nor U2159 (N_2159,N_1945,N_1031);
nand U2160 (N_2160,N_1328,N_1765);
or U2161 (N_2161,N_1690,N_1808);
and U2162 (N_2162,N_1429,N_1253);
or U2163 (N_2163,N_1281,N_1127);
nand U2164 (N_2164,N_1131,N_1372);
or U2165 (N_2165,N_1470,N_1819);
nand U2166 (N_2166,N_1691,N_1903);
and U2167 (N_2167,N_1140,N_1338);
nand U2168 (N_2168,N_1794,N_1120);
nand U2169 (N_2169,N_1491,N_1171);
nor U2170 (N_2170,N_1248,N_1105);
xnor U2171 (N_2171,N_1294,N_1327);
and U2172 (N_2172,N_1411,N_1453);
xnor U2173 (N_2173,N_1357,N_1342);
nor U2174 (N_2174,N_1367,N_1841);
nor U2175 (N_2175,N_1016,N_1269);
xor U2176 (N_2176,N_1930,N_1899);
and U2177 (N_2177,N_1718,N_1085);
nor U2178 (N_2178,N_1390,N_1540);
or U2179 (N_2179,N_1582,N_1155);
and U2180 (N_2180,N_1079,N_1863);
or U2181 (N_2181,N_1526,N_1335);
and U2182 (N_2182,N_1662,N_1568);
xnor U2183 (N_2183,N_1833,N_1048);
xor U2184 (N_2184,N_1065,N_1088);
nor U2185 (N_2185,N_1514,N_1953);
nor U2186 (N_2186,N_1810,N_1537);
nor U2187 (N_2187,N_1226,N_1979);
nor U2188 (N_2188,N_1991,N_1062);
xor U2189 (N_2189,N_1457,N_1572);
nor U2190 (N_2190,N_1737,N_1650);
xor U2191 (N_2191,N_1274,N_1675);
nor U2192 (N_2192,N_1711,N_1473);
and U2193 (N_2193,N_1444,N_1142);
and U2194 (N_2194,N_1629,N_1220);
or U2195 (N_2195,N_1256,N_1982);
or U2196 (N_2196,N_1815,N_1217);
and U2197 (N_2197,N_1358,N_1064);
xnor U2198 (N_2198,N_1034,N_1323);
nand U2199 (N_2199,N_1356,N_1407);
nand U2200 (N_2200,N_1360,N_1602);
xnor U2201 (N_2201,N_1830,N_1569);
and U2202 (N_2202,N_1781,N_1017);
xnor U2203 (N_2203,N_1299,N_1573);
nand U2204 (N_2204,N_1073,N_1871);
or U2205 (N_2205,N_1075,N_1415);
and U2206 (N_2206,N_1590,N_1861);
or U2207 (N_2207,N_1644,N_1674);
nand U2208 (N_2208,N_1282,N_1500);
nor U2209 (N_2209,N_1222,N_1519);
nor U2210 (N_2210,N_1413,N_1003);
or U2211 (N_2211,N_1974,N_1119);
nor U2212 (N_2212,N_1789,N_1891);
or U2213 (N_2213,N_1612,N_1752);
nand U2214 (N_2214,N_1928,N_1864);
and U2215 (N_2215,N_1071,N_1847);
xnor U2216 (N_2216,N_1975,N_1525);
nor U2217 (N_2217,N_1011,N_1694);
xnor U2218 (N_2218,N_1852,N_1408);
and U2219 (N_2219,N_1468,N_1359);
xnor U2220 (N_2220,N_1134,N_1742);
and U2221 (N_2221,N_1958,N_1516);
or U2222 (N_2222,N_1234,N_1755);
and U2223 (N_2223,N_1047,N_1257);
nor U2224 (N_2224,N_1441,N_1346);
and U2225 (N_2225,N_1619,N_1293);
or U2226 (N_2226,N_1361,N_1264);
nor U2227 (N_2227,N_1391,N_1207);
nor U2228 (N_2228,N_1238,N_1364);
nand U2229 (N_2229,N_1521,N_1409);
and U2230 (N_2230,N_1947,N_1302);
or U2231 (N_2231,N_1042,N_1270);
nand U2232 (N_2232,N_1086,N_1506);
or U2233 (N_2233,N_1798,N_1859);
nand U2234 (N_2234,N_1287,N_1362);
or U2235 (N_2235,N_1960,N_1633);
and U2236 (N_2236,N_1067,N_1564);
xor U2237 (N_2237,N_1421,N_1271);
xnor U2238 (N_2238,N_1559,N_1138);
xnor U2239 (N_2239,N_1591,N_1580);
xnor U2240 (N_2240,N_1934,N_1284);
nand U2241 (N_2241,N_1561,N_1598);
and U2242 (N_2242,N_1546,N_1913);
xor U2243 (N_2243,N_1289,N_1440);
xnor U2244 (N_2244,N_1990,N_1002);
or U2245 (N_2245,N_1427,N_1821);
or U2246 (N_2246,N_1660,N_1262);
xor U2247 (N_2247,N_1203,N_1970);
or U2248 (N_2248,N_1082,N_1149);
nand U2249 (N_2249,N_1844,N_1486);
nand U2250 (N_2250,N_1434,N_1194);
and U2251 (N_2251,N_1683,N_1597);
or U2252 (N_2252,N_1479,N_1838);
or U2253 (N_2253,N_1463,N_1076);
or U2254 (N_2254,N_1354,N_1512);
or U2255 (N_2255,N_1749,N_1493);
xnor U2256 (N_2256,N_1398,N_1729);
nand U2257 (N_2257,N_1704,N_1157);
nor U2258 (N_2258,N_1378,N_1199);
nand U2259 (N_2259,N_1848,N_1908);
and U2260 (N_2260,N_1036,N_1404);
xnor U2261 (N_2261,N_1471,N_1181);
nand U2262 (N_2262,N_1879,N_1697);
xnor U2263 (N_2263,N_1900,N_1575);
xor U2264 (N_2264,N_1851,N_1875);
and U2265 (N_2265,N_1843,N_1462);
or U2266 (N_2266,N_1324,N_1049);
nand U2267 (N_2267,N_1419,N_1375);
nand U2268 (N_2268,N_1925,N_1831);
xnor U2269 (N_2269,N_1296,N_1030);
nor U2270 (N_2270,N_1981,N_1009);
xor U2271 (N_2271,N_1962,N_1215);
nand U2272 (N_2272,N_1961,N_1152);
nor U2273 (N_2273,N_1658,N_1978);
nand U2274 (N_2274,N_1050,N_1345);
xor U2275 (N_2275,N_1114,N_1905);
or U2276 (N_2276,N_1380,N_1007);
nand U2277 (N_2277,N_1754,N_1051);
nor U2278 (N_2278,N_1876,N_1649);
and U2279 (N_2279,N_1822,N_1996);
and U2280 (N_2280,N_1972,N_1175);
nor U2281 (N_2281,N_1995,N_1028);
or U2282 (N_2282,N_1014,N_1497);
nand U2283 (N_2283,N_1371,N_1777);
nand U2284 (N_2284,N_1053,N_1200);
nor U2285 (N_2285,N_1349,N_1586);
and U2286 (N_2286,N_1796,N_1243);
and U2287 (N_2287,N_1236,N_1225);
nand U2288 (N_2288,N_1250,N_1678);
xor U2289 (N_2289,N_1221,N_1107);
or U2290 (N_2290,N_1544,N_1698);
xnor U2291 (N_2291,N_1428,N_1488);
nand U2292 (N_2292,N_1509,N_1083);
or U2293 (N_2293,N_1185,N_1201);
or U2294 (N_2294,N_1397,N_1476);
or U2295 (N_2295,N_1834,N_1890);
nor U2296 (N_2296,N_1532,N_1522);
nor U2297 (N_2297,N_1288,N_1922);
nor U2298 (N_2298,N_1565,N_1551);
xor U2299 (N_2299,N_1806,N_1277);
nand U2300 (N_2300,N_1376,N_1724);
nand U2301 (N_2301,N_1921,N_1484);
nand U2302 (N_2302,N_1539,N_1679);
nand U2303 (N_2303,N_1291,N_1098);
xor U2304 (N_2304,N_1118,N_1103);
or U2305 (N_2305,N_1304,N_1530);
and U2306 (N_2306,N_1889,N_1574);
nor U2307 (N_2307,N_1723,N_1699);
xor U2308 (N_2308,N_1601,N_1436);
nand U2309 (N_2309,N_1089,N_1229);
xnor U2310 (N_2310,N_1092,N_1447);
or U2311 (N_2311,N_1143,N_1693);
nor U2312 (N_2312,N_1837,N_1374);
nor U2313 (N_2313,N_1703,N_1084);
nand U2314 (N_2314,N_1290,N_1940);
or U2315 (N_2315,N_1123,N_1520);
nand U2316 (N_2316,N_1422,N_1165);
xnor U2317 (N_2317,N_1795,N_1012);
nor U2318 (N_2318,N_1230,N_1857);
nor U2319 (N_2319,N_1687,N_1414);
and U2320 (N_2320,N_1405,N_1595);
nor U2321 (N_2321,N_1710,N_1121);
nand U2322 (N_2322,N_1412,N_1654);
nand U2323 (N_2323,N_1579,N_1108);
xor U2324 (N_2324,N_1454,N_1556);
nand U2325 (N_2325,N_1128,N_1091);
or U2326 (N_2326,N_1400,N_1554);
and U2327 (N_2327,N_1314,N_1860);
or U2328 (N_2328,N_1008,N_1620);
or U2329 (N_2329,N_1562,N_1424);
and U2330 (N_2330,N_1956,N_1310);
or U2331 (N_2331,N_1770,N_1111);
and U2332 (N_2332,N_1139,N_1783);
nor U2333 (N_2333,N_1577,N_1344);
and U2334 (N_2334,N_1326,N_1791);
and U2335 (N_2335,N_1524,N_1726);
xnor U2336 (N_2336,N_1184,N_1987);
or U2337 (N_2337,N_1786,N_1709);
xor U2338 (N_2338,N_1167,N_1418);
or U2339 (N_2339,N_1779,N_1909);
nor U2340 (N_2340,N_1511,N_1639);
or U2341 (N_2341,N_1776,N_1799);
or U2342 (N_2342,N_1603,N_1666);
nor U2343 (N_2343,N_1038,N_1240);
nand U2344 (N_2344,N_1166,N_1183);
and U2345 (N_2345,N_1153,N_1712);
and U2346 (N_2346,N_1906,N_1156);
xnor U2347 (N_2347,N_1224,N_1396);
and U2348 (N_2348,N_1757,N_1651);
and U2349 (N_2349,N_1461,N_1018);
and U2350 (N_2350,N_1624,N_1097);
nand U2351 (N_2351,N_1787,N_1279);
xor U2352 (N_2352,N_1104,N_1377);
nand U2353 (N_2353,N_1174,N_1732);
nand U2354 (N_2354,N_1035,N_1557);
xor U2355 (N_2355,N_1438,N_1780);
nand U2356 (N_2356,N_1333,N_1309);
xor U2357 (N_2357,N_1747,N_1179);
and U2358 (N_2358,N_1077,N_1316);
or U2359 (N_2359,N_1116,N_1842);
and U2360 (N_2360,N_1507,N_1677);
xor U2361 (N_2361,N_1738,N_1576);
nand U2362 (N_2362,N_1237,N_1764);
nor U2363 (N_2363,N_1950,N_1653);
and U2364 (N_2364,N_1715,N_1589);
nor U2365 (N_2365,N_1971,N_1286);
xnor U2366 (N_2366,N_1058,N_1751);
xor U2367 (N_2367,N_1494,N_1385);
nand U2368 (N_2368,N_1006,N_1740);
nor U2369 (N_2369,N_1812,N_1276);
or U2370 (N_2370,N_1176,N_1878);
or U2371 (N_2371,N_1606,N_1040);
nand U2372 (N_2372,N_1692,N_1774);
or U2373 (N_2373,N_1931,N_1946);
or U2374 (N_2374,N_1696,N_1721);
xnor U2375 (N_2375,N_1983,N_1161);
nor U2376 (N_2376,N_1817,N_1628);
xnor U2377 (N_2377,N_1827,N_1642);
and U2378 (N_2378,N_1249,N_1384);
nor U2379 (N_2379,N_1331,N_1826);
nand U2380 (N_2380,N_1489,N_1566);
or U2381 (N_2381,N_1938,N_1151);
or U2382 (N_2382,N_1744,N_1163);
xnor U2383 (N_2383,N_1458,N_1283);
or U2384 (N_2384,N_1655,N_1719);
xor U2385 (N_2385,N_1057,N_1188);
or U2386 (N_2386,N_1431,N_1305);
or U2387 (N_2387,N_1206,N_1910);
and U2388 (N_2388,N_1942,N_1069);
nor U2389 (N_2389,N_1474,N_1004);
xor U2390 (N_2390,N_1020,N_1477);
nor U2391 (N_2391,N_1439,N_1168);
nand U2392 (N_2392,N_1873,N_1733);
xnor U2393 (N_2393,N_1169,N_1984);
xnor U2394 (N_2394,N_1056,N_1117);
or U2395 (N_2395,N_1363,N_1080);
xor U2396 (N_2396,N_1231,N_1109);
nand U2397 (N_2397,N_1150,N_1968);
nand U2398 (N_2398,N_1788,N_1395);
nand U2399 (N_2399,N_1490,N_1607);
and U2400 (N_2400,N_1802,N_1024);
xnor U2401 (N_2401,N_1504,N_1885);
and U2402 (N_2402,N_1626,N_1483);
or U2403 (N_2403,N_1393,N_1805);
or U2404 (N_2404,N_1980,N_1026);
nor U2405 (N_2405,N_1994,N_1952);
nand U2406 (N_2406,N_1671,N_1268);
nor U2407 (N_2407,N_1923,N_1992);
and U2408 (N_2408,N_1531,N_1313);
or U2409 (N_2409,N_1306,N_1896);
nor U2410 (N_2410,N_1845,N_1963);
nor U2411 (N_2411,N_1272,N_1499);
and U2412 (N_2412,N_1600,N_1924);
nor U2413 (N_2413,N_1178,N_1095);
and U2414 (N_2414,N_1849,N_1329);
and U2415 (N_2415,N_1663,N_1588);
xnor U2416 (N_2416,N_1467,N_1242);
nand U2417 (N_2417,N_1768,N_1608);
nor U2418 (N_2418,N_1937,N_1022);
and U2419 (N_2419,N_1790,N_1340);
nor U2420 (N_2420,N_1322,N_1368);
nand U2421 (N_2421,N_1684,N_1877);
xnor U2422 (N_2422,N_1423,N_1973);
xor U2423 (N_2423,N_1988,N_1137);
and U2424 (N_2424,N_1204,N_1052);
xor U2425 (N_2425,N_1627,N_1343);
or U2426 (N_2426,N_1558,N_1320);
nor U2427 (N_2427,N_1529,N_1039);
and U2428 (N_2428,N_1435,N_1025);
nand U2429 (N_2429,N_1478,N_1536);
xor U2430 (N_2430,N_1702,N_1640);
or U2431 (N_2431,N_1661,N_1592);
xnor U2432 (N_2432,N_1443,N_1251);
and U2433 (N_2433,N_1985,N_1518);
and U2434 (N_2434,N_1535,N_1862);
nand U2435 (N_2435,N_1263,N_1686);
nand U2436 (N_2436,N_1800,N_1319);
and U2437 (N_2437,N_1273,N_1336);
and U2438 (N_2438,N_1154,N_1872);
nor U2439 (N_2439,N_1725,N_1701);
xor U2440 (N_2440,N_1874,N_1881);
or U2441 (N_2441,N_1352,N_1258);
nand U2442 (N_2442,N_1235,N_1099);
and U2443 (N_2443,N_1773,N_1292);
xnor U2444 (N_2444,N_1348,N_1295);
xnor U2445 (N_2445,N_1442,N_1239);
xor U2446 (N_2446,N_1610,N_1055);
or U2447 (N_2447,N_1063,N_1647);
nand U2448 (N_2448,N_1638,N_1402);
and U2449 (N_2449,N_1417,N_1581);
xor U2450 (N_2450,N_1894,N_1736);
nand U2451 (N_2451,N_1734,N_1865);
nand U2452 (N_2452,N_1186,N_1132);
nand U2453 (N_2453,N_1868,N_1135);
nand U2454 (N_2454,N_1637,N_1318);
or U2455 (N_2455,N_1673,N_1853);
nor U2456 (N_2456,N_1667,N_1656);
xnor U2457 (N_2457,N_1630,N_1341);
nand U2458 (N_2458,N_1622,N_1410);
nor U2459 (N_2459,N_1054,N_1255);
and U2460 (N_2460,N_1766,N_1094);
nand U2461 (N_2461,N_1587,N_1501);
nand U2462 (N_2462,N_1146,N_1955);
or U2463 (N_2463,N_1492,N_1005);
nand U2464 (N_2464,N_1113,N_1389);
nor U2465 (N_2465,N_1854,N_1365);
or U2466 (N_2466,N_1379,N_1855);
nor U2467 (N_2467,N_1124,N_1399);
xnor U2468 (N_2468,N_1727,N_1892);
xnor U2469 (N_2469,N_1705,N_1665);
xor U2470 (N_2470,N_1548,N_1560);
nand U2471 (N_2471,N_1115,N_1944);
xor U2472 (N_2472,N_1818,N_1523);
xnor U2473 (N_2473,N_1066,N_1148);
xor U2474 (N_2474,N_1714,N_1681);
nand U2475 (N_2475,N_1265,N_1044);
nand U2476 (N_2476,N_1648,N_1213);
xnor U2477 (N_2477,N_1911,N_1232);
xnor U2478 (N_2478,N_1244,N_1246);
or U2479 (N_2479,N_1228,N_1797);
nor U2480 (N_2480,N_1202,N_1164);
nand U2481 (N_2481,N_1641,N_1785);
nand U2482 (N_2482,N_1941,N_1416);
nand U2483 (N_2483,N_1125,N_1689);
nor U2484 (N_2484,N_1811,N_1897);
xor U2485 (N_2485,N_1043,N_1144);
and U2486 (N_2486,N_1756,N_1920);
and U2487 (N_2487,N_1469,N_1430);
and U2488 (N_2488,N_1750,N_1543);
and U2489 (N_2489,N_1997,N_1192);
and U2490 (N_2490,N_1070,N_1456);
xor U2491 (N_2491,N_1912,N_1998);
and U2492 (N_2492,N_1829,N_1748);
or U2493 (N_2493,N_1739,N_1533);
and U2494 (N_2494,N_1260,N_1839);
nor U2495 (N_2495,N_1177,N_1772);
nor U2496 (N_2496,N_1563,N_1888);
xor U2497 (N_2497,N_1809,N_1189);
nand U2498 (N_2498,N_1481,N_1332);
nor U2499 (N_2499,N_1061,N_1147);
xnor U2500 (N_2500,N_1931,N_1744);
nand U2501 (N_2501,N_1623,N_1921);
nand U2502 (N_2502,N_1997,N_1836);
nand U2503 (N_2503,N_1968,N_1360);
nor U2504 (N_2504,N_1315,N_1415);
or U2505 (N_2505,N_1090,N_1633);
nor U2506 (N_2506,N_1003,N_1563);
or U2507 (N_2507,N_1588,N_1120);
nor U2508 (N_2508,N_1057,N_1283);
and U2509 (N_2509,N_1100,N_1799);
xor U2510 (N_2510,N_1453,N_1393);
and U2511 (N_2511,N_1957,N_1748);
and U2512 (N_2512,N_1529,N_1034);
nor U2513 (N_2513,N_1429,N_1091);
or U2514 (N_2514,N_1846,N_1441);
xor U2515 (N_2515,N_1424,N_1809);
nand U2516 (N_2516,N_1124,N_1729);
and U2517 (N_2517,N_1683,N_1168);
nor U2518 (N_2518,N_1407,N_1244);
and U2519 (N_2519,N_1888,N_1486);
and U2520 (N_2520,N_1906,N_1651);
nand U2521 (N_2521,N_1109,N_1874);
xnor U2522 (N_2522,N_1305,N_1432);
and U2523 (N_2523,N_1854,N_1561);
and U2524 (N_2524,N_1273,N_1833);
or U2525 (N_2525,N_1981,N_1376);
or U2526 (N_2526,N_1650,N_1773);
xor U2527 (N_2527,N_1703,N_1401);
nor U2528 (N_2528,N_1633,N_1742);
and U2529 (N_2529,N_1841,N_1122);
nor U2530 (N_2530,N_1403,N_1856);
xnor U2531 (N_2531,N_1417,N_1099);
and U2532 (N_2532,N_1042,N_1049);
nor U2533 (N_2533,N_1590,N_1236);
xor U2534 (N_2534,N_1458,N_1875);
nor U2535 (N_2535,N_1988,N_1675);
nor U2536 (N_2536,N_1166,N_1169);
nor U2537 (N_2537,N_1671,N_1933);
and U2538 (N_2538,N_1496,N_1979);
nor U2539 (N_2539,N_1787,N_1821);
nand U2540 (N_2540,N_1961,N_1692);
or U2541 (N_2541,N_1348,N_1402);
nand U2542 (N_2542,N_1588,N_1823);
xor U2543 (N_2543,N_1252,N_1533);
or U2544 (N_2544,N_1756,N_1427);
xnor U2545 (N_2545,N_1878,N_1366);
nor U2546 (N_2546,N_1892,N_1599);
nor U2547 (N_2547,N_1654,N_1637);
xnor U2548 (N_2548,N_1979,N_1007);
nand U2549 (N_2549,N_1602,N_1664);
nand U2550 (N_2550,N_1768,N_1738);
nand U2551 (N_2551,N_1340,N_1614);
nor U2552 (N_2552,N_1524,N_1511);
nand U2553 (N_2553,N_1816,N_1392);
and U2554 (N_2554,N_1851,N_1980);
nand U2555 (N_2555,N_1061,N_1288);
or U2556 (N_2556,N_1546,N_1049);
or U2557 (N_2557,N_1932,N_1957);
and U2558 (N_2558,N_1094,N_1798);
xor U2559 (N_2559,N_1488,N_1911);
nand U2560 (N_2560,N_1129,N_1997);
xor U2561 (N_2561,N_1521,N_1413);
xor U2562 (N_2562,N_1791,N_1465);
xor U2563 (N_2563,N_1185,N_1986);
xnor U2564 (N_2564,N_1485,N_1330);
nor U2565 (N_2565,N_1835,N_1576);
or U2566 (N_2566,N_1974,N_1789);
xor U2567 (N_2567,N_1700,N_1830);
nor U2568 (N_2568,N_1282,N_1050);
xnor U2569 (N_2569,N_1437,N_1959);
nor U2570 (N_2570,N_1396,N_1214);
xor U2571 (N_2571,N_1655,N_1523);
nand U2572 (N_2572,N_1541,N_1799);
nand U2573 (N_2573,N_1162,N_1679);
nand U2574 (N_2574,N_1513,N_1610);
nor U2575 (N_2575,N_1837,N_1526);
nor U2576 (N_2576,N_1790,N_1439);
and U2577 (N_2577,N_1296,N_1462);
or U2578 (N_2578,N_1082,N_1067);
xnor U2579 (N_2579,N_1292,N_1118);
or U2580 (N_2580,N_1236,N_1418);
or U2581 (N_2581,N_1706,N_1730);
nor U2582 (N_2582,N_1897,N_1280);
nor U2583 (N_2583,N_1074,N_1709);
xor U2584 (N_2584,N_1616,N_1562);
or U2585 (N_2585,N_1974,N_1583);
and U2586 (N_2586,N_1825,N_1153);
or U2587 (N_2587,N_1920,N_1003);
xnor U2588 (N_2588,N_1587,N_1889);
nand U2589 (N_2589,N_1208,N_1259);
or U2590 (N_2590,N_1139,N_1238);
nor U2591 (N_2591,N_1076,N_1751);
nor U2592 (N_2592,N_1365,N_1884);
nand U2593 (N_2593,N_1992,N_1581);
and U2594 (N_2594,N_1899,N_1892);
and U2595 (N_2595,N_1762,N_1629);
nor U2596 (N_2596,N_1113,N_1287);
nand U2597 (N_2597,N_1098,N_1137);
and U2598 (N_2598,N_1834,N_1869);
and U2599 (N_2599,N_1919,N_1017);
and U2600 (N_2600,N_1971,N_1202);
xnor U2601 (N_2601,N_1881,N_1113);
nand U2602 (N_2602,N_1248,N_1951);
xor U2603 (N_2603,N_1866,N_1522);
and U2604 (N_2604,N_1577,N_1122);
and U2605 (N_2605,N_1079,N_1113);
or U2606 (N_2606,N_1456,N_1912);
nand U2607 (N_2607,N_1106,N_1902);
and U2608 (N_2608,N_1581,N_1050);
nand U2609 (N_2609,N_1571,N_1198);
xor U2610 (N_2610,N_1235,N_1437);
and U2611 (N_2611,N_1879,N_1002);
nand U2612 (N_2612,N_1023,N_1225);
or U2613 (N_2613,N_1529,N_1640);
nand U2614 (N_2614,N_1995,N_1164);
or U2615 (N_2615,N_1595,N_1015);
nor U2616 (N_2616,N_1806,N_1235);
and U2617 (N_2617,N_1324,N_1079);
xor U2618 (N_2618,N_1668,N_1737);
nor U2619 (N_2619,N_1222,N_1549);
nand U2620 (N_2620,N_1595,N_1986);
xnor U2621 (N_2621,N_1334,N_1854);
nor U2622 (N_2622,N_1522,N_1738);
xnor U2623 (N_2623,N_1258,N_1073);
nor U2624 (N_2624,N_1314,N_1537);
or U2625 (N_2625,N_1893,N_1760);
xnor U2626 (N_2626,N_1436,N_1616);
or U2627 (N_2627,N_1364,N_1392);
and U2628 (N_2628,N_1764,N_1162);
nand U2629 (N_2629,N_1977,N_1007);
nor U2630 (N_2630,N_1456,N_1648);
nor U2631 (N_2631,N_1039,N_1143);
xor U2632 (N_2632,N_1725,N_1445);
nand U2633 (N_2633,N_1349,N_1238);
xnor U2634 (N_2634,N_1807,N_1791);
or U2635 (N_2635,N_1402,N_1916);
nor U2636 (N_2636,N_1754,N_1692);
or U2637 (N_2637,N_1066,N_1655);
nand U2638 (N_2638,N_1950,N_1176);
nor U2639 (N_2639,N_1106,N_1077);
nand U2640 (N_2640,N_1942,N_1034);
and U2641 (N_2641,N_1661,N_1982);
or U2642 (N_2642,N_1432,N_1789);
nand U2643 (N_2643,N_1713,N_1088);
nand U2644 (N_2644,N_1695,N_1350);
nor U2645 (N_2645,N_1230,N_1031);
xnor U2646 (N_2646,N_1446,N_1564);
nand U2647 (N_2647,N_1719,N_1924);
nand U2648 (N_2648,N_1054,N_1098);
nand U2649 (N_2649,N_1970,N_1506);
xnor U2650 (N_2650,N_1474,N_1514);
or U2651 (N_2651,N_1533,N_1664);
xor U2652 (N_2652,N_1942,N_1417);
nand U2653 (N_2653,N_1023,N_1964);
and U2654 (N_2654,N_1170,N_1333);
and U2655 (N_2655,N_1510,N_1928);
xor U2656 (N_2656,N_1996,N_1672);
nor U2657 (N_2657,N_1512,N_1327);
nor U2658 (N_2658,N_1467,N_1796);
nand U2659 (N_2659,N_1925,N_1537);
xnor U2660 (N_2660,N_1809,N_1114);
and U2661 (N_2661,N_1632,N_1047);
nand U2662 (N_2662,N_1098,N_1704);
or U2663 (N_2663,N_1965,N_1543);
and U2664 (N_2664,N_1197,N_1475);
and U2665 (N_2665,N_1706,N_1068);
xor U2666 (N_2666,N_1294,N_1631);
or U2667 (N_2667,N_1971,N_1144);
xnor U2668 (N_2668,N_1086,N_1356);
xor U2669 (N_2669,N_1375,N_1567);
nand U2670 (N_2670,N_1468,N_1883);
xnor U2671 (N_2671,N_1103,N_1024);
or U2672 (N_2672,N_1811,N_1590);
nand U2673 (N_2673,N_1564,N_1838);
nand U2674 (N_2674,N_1289,N_1087);
xor U2675 (N_2675,N_1944,N_1622);
xnor U2676 (N_2676,N_1347,N_1043);
or U2677 (N_2677,N_1534,N_1520);
nand U2678 (N_2678,N_1064,N_1242);
nor U2679 (N_2679,N_1243,N_1563);
xnor U2680 (N_2680,N_1963,N_1109);
xor U2681 (N_2681,N_1250,N_1467);
nor U2682 (N_2682,N_1439,N_1224);
and U2683 (N_2683,N_1667,N_1708);
or U2684 (N_2684,N_1547,N_1612);
xnor U2685 (N_2685,N_1132,N_1921);
or U2686 (N_2686,N_1084,N_1162);
nand U2687 (N_2687,N_1489,N_1819);
xnor U2688 (N_2688,N_1853,N_1308);
and U2689 (N_2689,N_1878,N_1379);
and U2690 (N_2690,N_1330,N_1052);
and U2691 (N_2691,N_1282,N_1573);
or U2692 (N_2692,N_1066,N_1115);
nor U2693 (N_2693,N_1980,N_1550);
xnor U2694 (N_2694,N_1989,N_1220);
or U2695 (N_2695,N_1577,N_1797);
xnor U2696 (N_2696,N_1260,N_1328);
nor U2697 (N_2697,N_1563,N_1974);
or U2698 (N_2698,N_1262,N_1481);
nand U2699 (N_2699,N_1894,N_1048);
nor U2700 (N_2700,N_1178,N_1569);
nand U2701 (N_2701,N_1456,N_1659);
xor U2702 (N_2702,N_1878,N_1637);
nor U2703 (N_2703,N_1111,N_1202);
or U2704 (N_2704,N_1586,N_1726);
and U2705 (N_2705,N_1463,N_1205);
nand U2706 (N_2706,N_1257,N_1010);
nor U2707 (N_2707,N_1269,N_1643);
or U2708 (N_2708,N_1939,N_1580);
or U2709 (N_2709,N_1703,N_1605);
xnor U2710 (N_2710,N_1087,N_1571);
or U2711 (N_2711,N_1827,N_1012);
nor U2712 (N_2712,N_1523,N_1615);
xor U2713 (N_2713,N_1659,N_1895);
nor U2714 (N_2714,N_1665,N_1788);
xor U2715 (N_2715,N_1282,N_1864);
nand U2716 (N_2716,N_1902,N_1245);
and U2717 (N_2717,N_1429,N_1562);
nand U2718 (N_2718,N_1313,N_1233);
nor U2719 (N_2719,N_1230,N_1782);
or U2720 (N_2720,N_1034,N_1268);
xnor U2721 (N_2721,N_1158,N_1928);
xor U2722 (N_2722,N_1617,N_1013);
or U2723 (N_2723,N_1243,N_1947);
nor U2724 (N_2724,N_1871,N_1938);
nand U2725 (N_2725,N_1548,N_1156);
nand U2726 (N_2726,N_1922,N_1805);
or U2727 (N_2727,N_1933,N_1083);
and U2728 (N_2728,N_1183,N_1916);
or U2729 (N_2729,N_1244,N_1955);
nand U2730 (N_2730,N_1674,N_1771);
or U2731 (N_2731,N_1878,N_1297);
and U2732 (N_2732,N_1664,N_1708);
or U2733 (N_2733,N_1770,N_1243);
and U2734 (N_2734,N_1614,N_1105);
nand U2735 (N_2735,N_1142,N_1679);
xnor U2736 (N_2736,N_1757,N_1799);
nor U2737 (N_2737,N_1671,N_1074);
and U2738 (N_2738,N_1821,N_1192);
nand U2739 (N_2739,N_1174,N_1317);
or U2740 (N_2740,N_1924,N_1376);
or U2741 (N_2741,N_1360,N_1801);
nor U2742 (N_2742,N_1727,N_1736);
or U2743 (N_2743,N_1801,N_1629);
xor U2744 (N_2744,N_1412,N_1205);
nor U2745 (N_2745,N_1174,N_1199);
nor U2746 (N_2746,N_1537,N_1662);
nor U2747 (N_2747,N_1480,N_1316);
or U2748 (N_2748,N_1082,N_1516);
nand U2749 (N_2749,N_1397,N_1269);
nand U2750 (N_2750,N_1186,N_1968);
or U2751 (N_2751,N_1739,N_1775);
nor U2752 (N_2752,N_1224,N_1566);
and U2753 (N_2753,N_1346,N_1139);
or U2754 (N_2754,N_1040,N_1533);
nand U2755 (N_2755,N_1721,N_1925);
or U2756 (N_2756,N_1368,N_1229);
nand U2757 (N_2757,N_1061,N_1748);
nor U2758 (N_2758,N_1749,N_1308);
and U2759 (N_2759,N_1050,N_1222);
or U2760 (N_2760,N_1320,N_1613);
xor U2761 (N_2761,N_1929,N_1114);
and U2762 (N_2762,N_1993,N_1652);
nand U2763 (N_2763,N_1226,N_1574);
and U2764 (N_2764,N_1990,N_1318);
nor U2765 (N_2765,N_1357,N_1866);
and U2766 (N_2766,N_1665,N_1148);
or U2767 (N_2767,N_1119,N_1654);
and U2768 (N_2768,N_1046,N_1635);
nand U2769 (N_2769,N_1103,N_1697);
xnor U2770 (N_2770,N_1337,N_1964);
or U2771 (N_2771,N_1637,N_1038);
and U2772 (N_2772,N_1222,N_1376);
or U2773 (N_2773,N_1525,N_1945);
xnor U2774 (N_2774,N_1069,N_1505);
and U2775 (N_2775,N_1742,N_1645);
xor U2776 (N_2776,N_1630,N_1213);
nand U2777 (N_2777,N_1995,N_1529);
and U2778 (N_2778,N_1452,N_1411);
xnor U2779 (N_2779,N_1956,N_1013);
nor U2780 (N_2780,N_1046,N_1435);
xnor U2781 (N_2781,N_1496,N_1539);
xor U2782 (N_2782,N_1205,N_1197);
nor U2783 (N_2783,N_1553,N_1009);
xor U2784 (N_2784,N_1966,N_1762);
nand U2785 (N_2785,N_1512,N_1333);
or U2786 (N_2786,N_1189,N_1302);
nand U2787 (N_2787,N_1621,N_1204);
nand U2788 (N_2788,N_1595,N_1832);
nand U2789 (N_2789,N_1784,N_1822);
nand U2790 (N_2790,N_1815,N_1037);
nor U2791 (N_2791,N_1752,N_1203);
or U2792 (N_2792,N_1037,N_1582);
nand U2793 (N_2793,N_1636,N_1800);
nor U2794 (N_2794,N_1763,N_1907);
nor U2795 (N_2795,N_1755,N_1771);
or U2796 (N_2796,N_1491,N_1360);
and U2797 (N_2797,N_1028,N_1033);
or U2798 (N_2798,N_1430,N_1493);
or U2799 (N_2799,N_1313,N_1608);
and U2800 (N_2800,N_1823,N_1150);
nand U2801 (N_2801,N_1982,N_1373);
and U2802 (N_2802,N_1936,N_1361);
nor U2803 (N_2803,N_1485,N_1087);
and U2804 (N_2804,N_1285,N_1854);
or U2805 (N_2805,N_1057,N_1621);
and U2806 (N_2806,N_1703,N_1149);
and U2807 (N_2807,N_1118,N_1747);
nor U2808 (N_2808,N_1143,N_1459);
nor U2809 (N_2809,N_1517,N_1195);
nor U2810 (N_2810,N_1462,N_1549);
and U2811 (N_2811,N_1748,N_1325);
and U2812 (N_2812,N_1330,N_1303);
xnor U2813 (N_2813,N_1883,N_1852);
nand U2814 (N_2814,N_1745,N_1740);
or U2815 (N_2815,N_1207,N_1799);
nand U2816 (N_2816,N_1980,N_1972);
and U2817 (N_2817,N_1240,N_1727);
or U2818 (N_2818,N_1877,N_1375);
or U2819 (N_2819,N_1264,N_1449);
and U2820 (N_2820,N_1913,N_1027);
xnor U2821 (N_2821,N_1103,N_1330);
and U2822 (N_2822,N_1694,N_1017);
nor U2823 (N_2823,N_1049,N_1827);
nor U2824 (N_2824,N_1416,N_1609);
xor U2825 (N_2825,N_1096,N_1222);
nand U2826 (N_2826,N_1261,N_1282);
xor U2827 (N_2827,N_1102,N_1110);
nand U2828 (N_2828,N_1012,N_1473);
nand U2829 (N_2829,N_1756,N_1235);
and U2830 (N_2830,N_1887,N_1499);
and U2831 (N_2831,N_1874,N_1459);
or U2832 (N_2832,N_1411,N_1749);
xnor U2833 (N_2833,N_1148,N_1188);
or U2834 (N_2834,N_1405,N_1185);
and U2835 (N_2835,N_1255,N_1624);
and U2836 (N_2836,N_1268,N_1338);
nor U2837 (N_2837,N_1207,N_1299);
or U2838 (N_2838,N_1388,N_1575);
xor U2839 (N_2839,N_1635,N_1114);
and U2840 (N_2840,N_1946,N_1069);
and U2841 (N_2841,N_1730,N_1800);
and U2842 (N_2842,N_1439,N_1977);
and U2843 (N_2843,N_1844,N_1674);
and U2844 (N_2844,N_1375,N_1472);
xnor U2845 (N_2845,N_1235,N_1732);
or U2846 (N_2846,N_1563,N_1368);
xor U2847 (N_2847,N_1186,N_1978);
and U2848 (N_2848,N_1848,N_1870);
or U2849 (N_2849,N_1829,N_1488);
nor U2850 (N_2850,N_1870,N_1748);
or U2851 (N_2851,N_1280,N_1565);
xnor U2852 (N_2852,N_1955,N_1891);
xor U2853 (N_2853,N_1781,N_1274);
nor U2854 (N_2854,N_1002,N_1261);
nor U2855 (N_2855,N_1860,N_1671);
nand U2856 (N_2856,N_1894,N_1041);
and U2857 (N_2857,N_1459,N_1693);
and U2858 (N_2858,N_1846,N_1621);
or U2859 (N_2859,N_1985,N_1170);
or U2860 (N_2860,N_1945,N_1246);
or U2861 (N_2861,N_1441,N_1883);
nor U2862 (N_2862,N_1371,N_1047);
xor U2863 (N_2863,N_1611,N_1227);
or U2864 (N_2864,N_1056,N_1772);
nand U2865 (N_2865,N_1515,N_1100);
and U2866 (N_2866,N_1586,N_1483);
xnor U2867 (N_2867,N_1066,N_1548);
xor U2868 (N_2868,N_1831,N_1563);
nor U2869 (N_2869,N_1939,N_1267);
xnor U2870 (N_2870,N_1555,N_1883);
nor U2871 (N_2871,N_1544,N_1948);
xnor U2872 (N_2872,N_1001,N_1770);
and U2873 (N_2873,N_1025,N_1627);
or U2874 (N_2874,N_1677,N_1171);
nand U2875 (N_2875,N_1411,N_1576);
xnor U2876 (N_2876,N_1161,N_1115);
nand U2877 (N_2877,N_1560,N_1061);
nand U2878 (N_2878,N_1588,N_1395);
nand U2879 (N_2879,N_1700,N_1331);
or U2880 (N_2880,N_1482,N_1409);
xnor U2881 (N_2881,N_1261,N_1062);
nor U2882 (N_2882,N_1567,N_1052);
nor U2883 (N_2883,N_1988,N_1113);
and U2884 (N_2884,N_1822,N_1625);
nor U2885 (N_2885,N_1521,N_1887);
and U2886 (N_2886,N_1252,N_1472);
or U2887 (N_2887,N_1323,N_1941);
or U2888 (N_2888,N_1118,N_1410);
nand U2889 (N_2889,N_1561,N_1630);
or U2890 (N_2890,N_1972,N_1989);
and U2891 (N_2891,N_1579,N_1700);
or U2892 (N_2892,N_1391,N_1622);
or U2893 (N_2893,N_1432,N_1488);
nand U2894 (N_2894,N_1804,N_1581);
nor U2895 (N_2895,N_1971,N_1417);
or U2896 (N_2896,N_1297,N_1512);
and U2897 (N_2897,N_1125,N_1838);
nor U2898 (N_2898,N_1038,N_1898);
and U2899 (N_2899,N_1886,N_1846);
and U2900 (N_2900,N_1532,N_1599);
or U2901 (N_2901,N_1065,N_1068);
nor U2902 (N_2902,N_1824,N_1874);
nand U2903 (N_2903,N_1970,N_1774);
nand U2904 (N_2904,N_1289,N_1426);
nor U2905 (N_2905,N_1004,N_1216);
or U2906 (N_2906,N_1963,N_1833);
or U2907 (N_2907,N_1164,N_1258);
xnor U2908 (N_2908,N_1573,N_1184);
nor U2909 (N_2909,N_1164,N_1363);
nand U2910 (N_2910,N_1612,N_1758);
or U2911 (N_2911,N_1434,N_1953);
nand U2912 (N_2912,N_1933,N_1984);
or U2913 (N_2913,N_1434,N_1844);
nand U2914 (N_2914,N_1361,N_1999);
and U2915 (N_2915,N_1323,N_1918);
and U2916 (N_2916,N_1591,N_1445);
nand U2917 (N_2917,N_1798,N_1392);
nor U2918 (N_2918,N_1670,N_1739);
nand U2919 (N_2919,N_1204,N_1671);
nand U2920 (N_2920,N_1487,N_1344);
nand U2921 (N_2921,N_1749,N_1113);
xor U2922 (N_2922,N_1855,N_1873);
nand U2923 (N_2923,N_1077,N_1331);
nor U2924 (N_2924,N_1455,N_1715);
and U2925 (N_2925,N_1540,N_1246);
xnor U2926 (N_2926,N_1309,N_1211);
nor U2927 (N_2927,N_1741,N_1008);
nand U2928 (N_2928,N_1070,N_1862);
xnor U2929 (N_2929,N_1826,N_1863);
nor U2930 (N_2930,N_1766,N_1008);
nor U2931 (N_2931,N_1436,N_1984);
or U2932 (N_2932,N_1187,N_1096);
and U2933 (N_2933,N_1510,N_1939);
or U2934 (N_2934,N_1713,N_1859);
and U2935 (N_2935,N_1090,N_1985);
nand U2936 (N_2936,N_1682,N_1989);
nand U2937 (N_2937,N_1769,N_1502);
and U2938 (N_2938,N_1202,N_1358);
nor U2939 (N_2939,N_1277,N_1790);
nand U2940 (N_2940,N_1053,N_1479);
nand U2941 (N_2941,N_1731,N_1022);
or U2942 (N_2942,N_1950,N_1728);
and U2943 (N_2943,N_1402,N_1594);
and U2944 (N_2944,N_1341,N_1508);
nor U2945 (N_2945,N_1380,N_1396);
nand U2946 (N_2946,N_1667,N_1071);
and U2947 (N_2947,N_1478,N_1919);
nand U2948 (N_2948,N_1517,N_1001);
nand U2949 (N_2949,N_1855,N_1894);
and U2950 (N_2950,N_1760,N_1683);
and U2951 (N_2951,N_1008,N_1509);
or U2952 (N_2952,N_1019,N_1225);
or U2953 (N_2953,N_1376,N_1315);
nor U2954 (N_2954,N_1486,N_1128);
nor U2955 (N_2955,N_1398,N_1589);
xor U2956 (N_2956,N_1969,N_1613);
xnor U2957 (N_2957,N_1891,N_1061);
nor U2958 (N_2958,N_1538,N_1810);
or U2959 (N_2959,N_1922,N_1551);
and U2960 (N_2960,N_1758,N_1069);
xor U2961 (N_2961,N_1514,N_1290);
nor U2962 (N_2962,N_1383,N_1567);
xor U2963 (N_2963,N_1653,N_1336);
and U2964 (N_2964,N_1763,N_1678);
or U2965 (N_2965,N_1076,N_1921);
xnor U2966 (N_2966,N_1357,N_1341);
or U2967 (N_2967,N_1619,N_1775);
nand U2968 (N_2968,N_1432,N_1195);
and U2969 (N_2969,N_1723,N_1286);
xor U2970 (N_2970,N_1524,N_1194);
xnor U2971 (N_2971,N_1794,N_1052);
nand U2972 (N_2972,N_1582,N_1191);
nor U2973 (N_2973,N_1809,N_1571);
nor U2974 (N_2974,N_1236,N_1238);
or U2975 (N_2975,N_1954,N_1971);
and U2976 (N_2976,N_1584,N_1369);
and U2977 (N_2977,N_1067,N_1809);
or U2978 (N_2978,N_1760,N_1119);
and U2979 (N_2979,N_1238,N_1536);
nand U2980 (N_2980,N_1709,N_1678);
nor U2981 (N_2981,N_1688,N_1933);
xnor U2982 (N_2982,N_1971,N_1354);
nor U2983 (N_2983,N_1187,N_1727);
and U2984 (N_2984,N_1083,N_1179);
xor U2985 (N_2985,N_1073,N_1307);
nand U2986 (N_2986,N_1004,N_1797);
nor U2987 (N_2987,N_1322,N_1312);
and U2988 (N_2988,N_1547,N_1400);
nand U2989 (N_2989,N_1596,N_1914);
and U2990 (N_2990,N_1695,N_1001);
nor U2991 (N_2991,N_1168,N_1444);
nand U2992 (N_2992,N_1086,N_1899);
xnor U2993 (N_2993,N_1790,N_1040);
or U2994 (N_2994,N_1250,N_1899);
nand U2995 (N_2995,N_1883,N_1483);
or U2996 (N_2996,N_1774,N_1948);
nor U2997 (N_2997,N_1735,N_1697);
or U2998 (N_2998,N_1628,N_1318);
and U2999 (N_2999,N_1696,N_1124);
nand U3000 (N_3000,N_2079,N_2349);
xor U3001 (N_3001,N_2387,N_2723);
and U3002 (N_3002,N_2166,N_2154);
and U3003 (N_3003,N_2578,N_2132);
and U3004 (N_3004,N_2089,N_2605);
nand U3005 (N_3005,N_2117,N_2244);
and U3006 (N_3006,N_2034,N_2688);
nand U3007 (N_3007,N_2914,N_2122);
and U3008 (N_3008,N_2844,N_2682);
nand U3009 (N_3009,N_2307,N_2480);
xor U3010 (N_3010,N_2736,N_2748);
nand U3011 (N_3011,N_2608,N_2583);
xor U3012 (N_3012,N_2932,N_2103);
and U3013 (N_3013,N_2717,N_2820);
xor U3014 (N_3014,N_2477,N_2162);
nand U3015 (N_3015,N_2807,N_2242);
nor U3016 (N_3016,N_2160,N_2450);
or U3017 (N_3017,N_2173,N_2335);
xor U3018 (N_3018,N_2017,N_2804);
or U3019 (N_3019,N_2975,N_2239);
and U3020 (N_3020,N_2272,N_2327);
xnor U3021 (N_3021,N_2436,N_2212);
xor U3022 (N_3022,N_2520,N_2850);
and U3023 (N_3023,N_2250,N_2375);
and U3024 (N_3024,N_2359,N_2793);
nand U3025 (N_3025,N_2991,N_2740);
nand U3026 (N_3026,N_2464,N_2847);
nor U3027 (N_3027,N_2594,N_2626);
and U3028 (N_3028,N_2245,N_2935);
xor U3029 (N_3029,N_2083,N_2111);
nand U3030 (N_3030,N_2779,N_2942);
xnor U3031 (N_3031,N_2445,N_2574);
nand U3032 (N_3032,N_2725,N_2255);
xor U3033 (N_3033,N_2398,N_2300);
xor U3034 (N_3034,N_2551,N_2232);
nor U3035 (N_3035,N_2163,N_2903);
nor U3036 (N_3036,N_2802,N_2159);
or U3037 (N_3037,N_2179,N_2518);
xnor U3038 (N_3038,N_2858,N_2192);
nor U3039 (N_3039,N_2050,N_2822);
nand U3040 (N_3040,N_2823,N_2509);
nor U3041 (N_3041,N_2277,N_2086);
or U3042 (N_3042,N_2229,N_2714);
and U3043 (N_3043,N_2483,N_2333);
nand U3044 (N_3044,N_2074,N_2648);
nand U3045 (N_3045,N_2488,N_2718);
or U3046 (N_3046,N_2266,N_2954);
xor U3047 (N_3047,N_2175,N_2440);
and U3048 (N_3048,N_2362,N_2121);
nand U3049 (N_3049,N_2618,N_2478);
nand U3050 (N_3050,N_2129,N_2555);
xnor U3051 (N_3051,N_2262,N_2570);
nand U3052 (N_3052,N_2655,N_2285);
nor U3053 (N_3053,N_2875,N_2538);
or U3054 (N_3054,N_2061,N_2247);
nor U3055 (N_3055,N_2028,N_2634);
nand U3056 (N_3056,N_2781,N_2884);
xor U3057 (N_3057,N_2891,N_2692);
and U3058 (N_3058,N_2747,N_2241);
xnor U3059 (N_3059,N_2306,N_2434);
and U3060 (N_3060,N_2169,N_2243);
xnor U3061 (N_3061,N_2762,N_2356);
and U3062 (N_3062,N_2170,N_2818);
and U3063 (N_3063,N_2185,N_2224);
xnor U3064 (N_3064,N_2339,N_2135);
or U3065 (N_3065,N_2941,N_2430);
nor U3066 (N_3066,N_2102,N_2067);
xnor U3067 (N_3067,N_2722,N_2829);
nand U3068 (N_3068,N_2222,N_2680);
and U3069 (N_3069,N_2646,N_2894);
or U3070 (N_3070,N_2649,N_2857);
xor U3071 (N_3071,N_2856,N_2145);
and U3072 (N_3072,N_2967,N_2606);
xor U3073 (N_3073,N_2075,N_2908);
nand U3074 (N_3074,N_2305,N_2656);
xor U3075 (N_3075,N_2883,N_2407);
xnor U3076 (N_3076,N_2238,N_2627);
nor U3077 (N_3077,N_2824,N_2734);
or U3078 (N_3078,N_2261,N_2280);
nand U3079 (N_3079,N_2458,N_2237);
or U3080 (N_3080,N_2293,N_2429);
xnor U3081 (N_3081,N_2350,N_2156);
xnor U3082 (N_3082,N_2052,N_2615);
or U3083 (N_3083,N_2765,N_2022);
nor U3084 (N_3084,N_2629,N_2841);
xnor U3085 (N_3085,N_2998,N_2855);
or U3086 (N_3086,N_2108,N_2544);
xor U3087 (N_3087,N_2826,N_2183);
nand U3088 (N_3088,N_2667,N_2755);
nand U3089 (N_3089,N_2233,N_2336);
and U3090 (N_3090,N_2417,N_2757);
nor U3091 (N_3091,N_2677,N_2180);
nand U3092 (N_3092,N_2959,N_2985);
nand U3093 (N_3093,N_2936,N_2716);
xnor U3094 (N_3094,N_2563,N_2146);
xor U3095 (N_3095,N_2465,N_2738);
nand U3096 (N_3096,N_2453,N_2413);
xor U3097 (N_3097,N_2663,N_2548);
and U3098 (N_3098,N_2670,N_2957);
or U3099 (N_3099,N_2486,N_2106);
or U3100 (N_3100,N_2813,N_2298);
xnor U3101 (N_3101,N_2977,N_2726);
nand U3102 (N_3102,N_2004,N_2438);
or U3103 (N_3103,N_2585,N_2961);
or U3104 (N_3104,N_2796,N_2611);
or U3105 (N_3105,N_2968,N_2878);
and U3106 (N_3106,N_2988,N_2294);
xnor U3107 (N_3107,N_2376,N_2926);
nor U3108 (N_3108,N_2918,N_2066);
and U3109 (N_3109,N_2475,N_2158);
xnor U3110 (N_3110,N_2130,N_2027);
xnor U3111 (N_3111,N_2925,N_2337);
nand U3112 (N_3112,N_2938,N_2297);
xor U3113 (N_3113,N_2927,N_2068);
nor U3114 (N_3114,N_2654,N_2764);
and U3115 (N_3115,N_2309,N_2502);
nor U3116 (N_3116,N_2225,N_2744);
nor U3117 (N_3117,N_2361,N_2395);
xnor U3118 (N_3118,N_2310,N_2394);
nand U3119 (N_3119,N_2142,N_2949);
or U3120 (N_3120,N_2834,N_2821);
nand U3121 (N_3121,N_2476,N_2901);
nand U3122 (N_3122,N_2276,N_2481);
and U3123 (N_3123,N_2202,N_2960);
nand U3124 (N_3124,N_2288,N_2887);
nor U3125 (N_3125,N_2099,N_2474);
or U3126 (N_3126,N_2040,N_2426);
or U3127 (N_3127,N_2193,N_2390);
nand U3128 (N_3128,N_2246,N_2161);
or U3129 (N_3129,N_2473,N_2269);
or U3130 (N_3130,N_2489,N_2787);
and U3131 (N_3131,N_2705,N_2389);
nand U3132 (N_3132,N_2549,N_2187);
xor U3133 (N_3133,N_2852,N_2871);
xnor U3134 (N_3134,N_2562,N_2093);
xor U3135 (N_3135,N_2018,N_2080);
nand U3136 (N_3136,N_2599,N_2775);
nor U3137 (N_3137,N_2650,N_2505);
nand U3138 (N_3138,N_2283,N_2076);
or U3139 (N_3139,N_2902,N_2660);
and U3140 (N_3140,N_2172,N_2900);
nor U3141 (N_3141,N_2569,N_2200);
or U3142 (N_3142,N_2109,N_2437);
and U3143 (N_3143,N_2746,N_2571);
nor U3144 (N_3144,N_2905,N_2439);
or U3145 (N_3145,N_2444,N_2866);
nand U3146 (N_3146,N_2418,N_2196);
and U3147 (N_3147,N_2321,N_2637);
nand U3148 (N_3148,N_2055,N_2534);
and U3149 (N_3149,N_2707,N_2147);
or U3150 (N_3150,N_2435,N_2039);
nor U3151 (N_3151,N_2256,N_2817);
or U3152 (N_3152,N_2979,N_2059);
nor U3153 (N_3153,N_2021,N_2839);
nand U3154 (N_3154,N_2492,N_2165);
xnor U3155 (N_3155,N_2433,N_2946);
nand U3156 (N_3156,N_2547,N_2064);
nand U3157 (N_3157,N_2745,N_2816);
nor U3158 (N_3158,N_2380,N_2600);
nand U3159 (N_3159,N_2522,N_2273);
xnor U3160 (N_3160,N_2621,N_2030);
xor U3161 (N_3161,N_2385,N_2009);
and U3162 (N_3162,N_2780,N_2760);
nor U3163 (N_3163,N_2207,N_2937);
or U3164 (N_3164,N_2046,N_2743);
nor U3165 (N_3165,N_2545,N_2733);
and U3166 (N_3166,N_2536,N_2194);
nor U3167 (N_3167,N_2907,N_2580);
xor U3168 (N_3168,N_2543,N_2416);
nor U3169 (N_3169,N_2057,N_2119);
and U3170 (N_3170,N_2964,N_2054);
or U3171 (N_3171,N_2730,N_2572);
xor U3172 (N_3172,N_2258,N_2124);
nor U3173 (N_3173,N_2636,N_2999);
and U3174 (N_3174,N_2329,N_2454);
xor U3175 (N_3175,N_2065,N_2609);
nand U3176 (N_3176,N_2996,N_2195);
xor U3177 (N_3177,N_2410,N_2217);
and U3178 (N_3178,N_2876,N_2507);
nand U3179 (N_3179,N_2593,N_2610);
nor U3180 (N_3180,N_2377,N_2213);
and U3181 (N_3181,N_2084,N_2976);
xnor U3182 (N_3182,N_2782,N_2323);
nand U3183 (N_3183,N_2916,N_2324);
nand U3184 (N_3184,N_2368,N_2719);
nand U3185 (N_3185,N_2687,N_2542);
and U3186 (N_3186,N_2992,N_2565);
nand U3187 (N_3187,N_2370,N_2056);
xnor U3188 (N_3188,N_2939,N_2047);
nand U3189 (N_3189,N_2251,N_2789);
or U3190 (N_3190,N_2471,N_2012);
nor U3191 (N_3191,N_2457,N_2091);
xor U3192 (N_3192,N_2487,N_2859);
and U3193 (N_3193,N_2911,N_2346);
and U3194 (N_3194,N_2943,N_2556);
or U3195 (N_3195,N_2644,N_2851);
or U3196 (N_3196,N_2763,N_2713);
nor U3197 (N_3197,N_2397,N_2498);
nand U3198 (N_3198,N_2402,N_2651);
or U3199 (N_3199,N_2930,N_2421);
nand U3200 (N_3200,N_2137,N_2128);
or U3201 (N_3201,N_2024,N_2803);
xor U3202 (N_3202,N_2786,N_2189);
or U3203 (N_3203,N_2809,N_2100);
or U3204 (N_3204,N_2973,N_2101);
nand U3205 (N_3205,N_2553,N_2302);
and U3206 (N_3206,N_2208,N_2231);
xnor U3207 (N_3207,N_2533,N_2861);
nand U3208 (N_3208,N_2299,N_2770);
and U3209 (N_3209,N_2127,N_2882);
nand U3210 (N_3210,N_2374,N_2291);
nor U3211 (N_3211,N_2446,N_2353);
nor U3212 (N_3212,N_2675,N_2575);
and U3213 (N_3213,N_2931,N_2835);
nand U3214 (N_3214,N_2422,N_2092);
nand U3215 (N_3215,N_2761,N_2315);
nor U3216 (N_3216,N_2920,N_2110);
or U3217 (N_3217,N_2097,N_2026);
and U3218 (N_3218,N_2589,N_2167);
nand U3219 (N_3219,N_2559,N_2073);
or U3220 (N_3220,N_2383,N_2051);
nand U3221 (N_3221,N_2983,N_2463);
xor U3222 (N_3222,N_2501,N_2703);
or U3223 (N_3223,N_2788,N_2567);
xor U3224 (N_3224,N_2699,N_2708);
and U3225 (N_3225,N_2526,N_2149);
or U3226 (N_3226,N_2778,N_2077);
nor U3227 (N_3227,N_2000,N_2114);
nor U3228 (N_3228,N_2624,N_2423);
nand U3229 (N_3229,N_2592,N_2304);
and U3230 (N_3230,N_2517,N_2521);
nor U3231 (N_3231,N_2071,N_2358);
or U3232 (N_3232,N_2922,N_2118);
nand U3233 (N_3233,N_2428,N_2371);
nor U3234 (N_3234,N_2322,N_2774);
or U3235 (N_3235,N_2317,N_2406);
nand U3236 (N_3236,N_2843,N_2155);
nor U3237 (N_3237,N_2546,N_2331);
nor U3238 (N_3238,N_2581,N_2525);
nor U3239 (N_3239,N_2105,N_2326);
or U3240 (N_3240,N_2287,N_2303);
and U3241 (N_3241,N_2772,N_2537);
xnor U3242 (N_3242,N_2993,N_2221);
xor U3243 (N_3243,N_2365,N_2750);
and U3244 (N_3244,N_2532,N_2603);
and U3245 (N_3245,N_2801,N_2669);
or U3246 (N_3246,N_2314,N_2769);
nand U3247 (N_3247,N_2341,N_2472);
nor U3248 (N_3248,N_2897,N_2484);
or U3249 (N_3249,N_2497,N_2947);
xnor U3250 (N_3250,N_2679,N_2424);
xor U3251 (N_3251,N_2657,N_2403);
nand U3252 (N_3252,N_2830,N_2831);
nor U3253 (N_3253,N_2598,N_2735);
nor U3254 (N_3254,N_2143,N_2928);
xnor U3255 (N_3255,N_2863,N_2284);
or U3256 (N_3256,N_2898,N_2819);
nor U3257 (N_3257,N_2720,N_2209);
nand U3258 (N_3258,N_2633,N_2016);
or U3259 (N_3259,N_2854,N_2301);
xnor U3260 (N_3260,N_2226,N_2728);
nand U3261 (N_3261,N_2904,N_2527);
nor U3262 (N_3262,N_2460,N_2812);
or U3263 (N_3263,N_2591,N_2539);
nor U3264 (N_3264,N_2678,N_2561);
nand U3265 (N_3265,N_2253,N_2493);
nor U3266 (N_3266,N_2205,N_2290);
nand U3267 (N_3267,N_2500,N_2666);
nand U3268 (N_3268,N_2771,N_2776);
or U3269 (N_3269,N_2252,N_2401);
nand U3270 (N_3270,N_2013,N_2447);
or U3271 (N_3271,N_2759,N_2254);
or U3272 (N_3272,N_2895,N_2204);
nand U3273 (N_3273,N_2178,N_2003);
nand U3274 (N_3274,N_2741,N_2363);
nor U3275 (N_3275,N_2892,N_2686);
or U3276 (N_3276,N_2710,N_2419);
and U3277 (N_3277,N_2257,N_2950);
xor U3278 (N_3278,N_2441,N_2994);
xnor U3279 (N_3279,N_2511,N_2836);
or U3280 (N_3280,N_2072,N_2602);
xnor U3281 (N_3281,N_2466,N_2384);
or U3282 (N_3282,N_2674,N_2576);
and U3283 (N_3283,N_2613,N_2148);
or U3284 (N_3284,N_2910,N_2035);
xnor U3285 (N_3285,N_2671,N_2877);
xnor U3286 (N_3286,N_2825,N_2963);
nand U3287 (N_3287,N_2095,N_2325);
or U3288 (N_3288,N_2015,N_2354);
or U3289 (N_3289,N_2643,N_2558);
nor U3290 (N_3290,N_2382,N_2062);
nand U3291 (N_3291,N_2853,N_2529);
xnor U3292 (N_3292,N_2404,N_2414);
or U3293 (N_3293,N_2347,N_2978);
nand U3294 (N_3294,N_2783,N_2890);
xor U3295 (N_3295,N_2739,N_2658);
nor U3296 (N_3296,N_2945,N_2279);
xnor U3297 (N_3297,N_2917,N_2881);
or U3298 (N_3298,N_2889,N_2867);
nor U3299 (N_3299,N_2690,N_2391);
nand U3300 (N_3300,N_2094,N_2982);
and U3301 (N_3301,N_2987,N_2431);
xnor U3302 (N_3302,N_2742,N_2702);
and U3303 (N_3303,N_2879,N_2485);
nand U3304 (N_3304,N_2704,N_2524);
xnor U3305 (N_3305,N_2001,N_2944);
nand U3306 (N_3306,N_2340,N_2312);
nand U3307 (N_3307,N_2698,N_2566);
nand U3308 (N_3308,N_2997,N_2442);
or U3309 (N_3309,N_2186,N_2259);
and U3310 (N_3310,N_2827,N_2685);
and U3311 (N_3311,N_2845,N_2727);
xor U3312 (N_3312,N_2448,N_2381);
nand U3313 (N_3313,N_2320,N_2712);
or U3314 (N_3314,N_2921,N_2459);
and U3315 (N_3315,N_2115,N_2098);
and U3316 (N_3316,N_2625,N_2230);
and U3317 (N_3317,N_2136,N_2794);
nor U3318 (N_3318,N_2623,N_2168);
nand U3319 (N_3319,N_2282,N_2612);
nor U3320 (N_3320,N_2838,N_2496);
nand U3321 (N_3321,N_2639,N_2316);
nand U3322 (N_3322,N_2409,N_2491);
nand U3323 (N_3323,N_2721,N_2711);
or U3324 (N_3324,N_2494,N_2519);
nand U3325 (N_3325,N_2271,N_2886);
or U3326 (N_3326,N_2635,N_2216);
nor U3327 (N_3327,N_2184,N_2125);
nand U3328 (N_3328,N_2456,N_2795);
or U3329 (N_3329,N_2510,N_2528);
nor U3330 (N_3330,N_2053,N_2096);
nand U3331 (N_3331,N_2134,N_2029);
xnor U3332 (N_3332,N_2694,N_2150);
nand U3333 (N_3333,N_2328,N_2800);
and U3334 (N_3334,N_2729,N_2564);
and U3335 (N_3335,N_2360,N_2405);
or U3336 (N_3336,N_2811,N_2351);
nand U3337 (N_3337,N_2181,N_2219);
nand U3338 (N_3338,N_2508,N_2955);
nand U3339 (N_3339,N_2929,N_2248);
and U3340 (N_3340,N_2151,N_2392);
or U3341 (N_3341,N_2171,N_2792);
nand U3342 (N_3342,N_2632,N_2995);
nand U3343 (N_3343,N_2768,N_2915);
nand U3344 (N_3344,N_2664,N_2638);
nand U3345 (N_3345,N_2379,N_2215);
and U3346 (N_3346,N_2467,N_2133);
xnor U3347 (N_3347,N_2345,N_2211);
or U3348 (N_3348,N_2116,N_2270);
nand U3349 (N_3349,N_2751,N_2724);
and U3350 (N_3350,N_2366,N_2120);
or U3351 (N_3351,N_2620,N_2749);
xnor U3352 (N_3352,N_2590,N_2701);
nand U3353 (N_3353,N_2278,N_2504);
or U3354 (N_3354,N_2037,N_2828);
and U3355 (N_3355,N_2235,N_2668);
nand U3356 (N_3356,N_2924,N_2791);
or U3357 (N_3357,N_2631,N_2846);
and U3358 (N_3358,N_2777,N_2731);
and U3359 (N_3359,N_2338,N_2989);
and U3360 (N_3360,N_2378,N_2281);
or U3361 (N_3361,N_2948,N_2953);
nand U3362 (N_3362,N_2236,N_2152);
nor U3363 (N_3363,N_2596,N_2899);
xnor U3364 (N_3364,N_2058,N_2700);
and U3365 (N_3365,N_2090,N_2043);
nand U3366 (N_3366,N_2234,N_2396);
and U3367 (N_3367,N_2506,N_2642);
nand U3368 (N_3368,N_2286,N_2342);
and U3369 (N_3369,N_2140,N_2176);
or U3370 (N_3370,N_2837,N_2573);
and U3371 (N_3371,N_2069,N_2044);
and U3372 (N_3372,N_2785,N_2364);
nor U3373 (N_3373,N_2676,N_2641);
nor U3374 (N_3374,N_2174,N_2808);
xnor U3375 (N_3375,N_2031,N_2958);
xnor U3376 (N_3376,N_2601,N_2372);
nand U3377 (N_3377,N_2607,N_2032);
and U3378 (N_3378,N_2190,N_2972);
or U3379 (N_3379,N_2990,N_2334);
xnor U3380 (N_3380,N_2706,N_2874);
and U3381 (N_3381,N_2191,N_2832);
and U3382 (N_3382,N_2662,N_2512);
nand U3383 (N_3383,N_2138,N_2318);
nor U3384 (N_3384,N_2557,N_2799);
or U3385 (N_3385,N_2514,N_2449);
and U3386 (N_3386,N_2956,N_2131);
nor U3387 (N_3387,N_2499,N_2344);
nor U3388 (N_3388,N_2696,N_2451);
nand U3389 (N_3389,N_2868,N_2348);
or U3390 (N_3390,N_2516,N_2595);
nor U3391 (N_3391,N_2971,N_2974);
nand U3392 (N_3392,N_2490,N_2737);
and U3393 (N_3393,N_2530,N_2070);
and U3394 (N_3394,N_2087,N_2470);
or U3395 (N_3395,N_2038,N_2008);
xnor U3396 (N_3396,N_2797,N_2645);
nand U3397 (N_3397,N_2014,N_2665);
or U3398 (N_3398,N_2684,N_2264);
and U3399 (N_3399,N_2647,N_2541);
or U3400 (N_3400,N_2554,N_2373);
or U3401 (N_3401,N_2869,N_2617);
nor U3402 (N_3402,N_2367,N_2860);
xor U3403 (N_3403,N_2153,N_2754);
nand U3404 (N_3404,N_2672,N_2420);
or U3405 (N_3405,N_2552,N_2319);
xnor U3406 (N_3406,N_2113,N_2653);
nor U3407 (N_3407,N_2584,N_2940);
nand U3408 (N_3408,N_2872,N_2412);
nand U3409 (N_3409,N_2011,N_2228);
nand U3410 (N_3410,N_2036,N_2970);
or U3411 (N_3411,N_2411,N_2962);
xor U3412 (N_3412,N_2683,N_2753);
or U3413 (N_3413,N_2078,N_2986);
xnor U3414 (N_3414,N_2332,N_2865);
nand U3415 (N_3415,N_2604,N_2019);
nand U3416 (N_3416,N_2199,N_2023);
nand U3417 (N_3417,N_2063,N_2123);
xor U3418 (N_3418,N_2295,N_2531);
xor U3419 (N_3419,N_2311,N_2462);
xor U3420 (N_3420,N_2984,N_2144);
xnor U3421 (N_3421,N_2218,N_2535);
and U3422 (N_3422,N_2614,N_2885);
nand U3423 (N_3423,N_2249,N_2214);
nor U3424 (N_3424,N_2197,N_2833);
nor U3425 (N_3425,N_2443,N_2756);
or U3426 (N_3426,N_2308,N_2805);
nand U3427 (N_3427,N_2427,N_2619);
nor U3428 (N_3428,N_2355,N_2432);
and U3429 (N_3429,N_2275,N_2400);
nand U3430 (N_3430,N_2815,N_2909);
xnor U3431 (N_3431,N_2888,N_2296);
xnor U3432 (N_3432,N_2042,N_2227);
nand U3433 (N_3433,N_2870,N_2386);
and U3434 (N_3434,N_2452,N_2715);
xnor U3435 (N_3435,N_2265,N_2896);
nand U3436 (N_3436,N_2085,N_2263);
or U3437 (N_3437,N_2223,N_2126);
nor U3438 (N_3438,N_2873,N_2913);
or U3439 (N_3439,N_2640,N_2966);
and U3440 (N_3440,N_2049,N_2002);
or U3441 (N_3441,N_2582,N_2659);
and U3442 (N_3442,N_2586,N_2513);
or U3443 (N_3443,N_2082,N_2880);
nand U3444 (N_3444,N_2482,N_2007);
or U3445 (N_3445,N_2399,N_2025);
and U3446 (N_3446,N_2164,N_2630);
nor U3447 (N_3447,N_2622,N_2661);
nand U3448 (N_3448,N_2709,N_2206);
or U3449 (N_3449,N_2107,N_2628);
nor U3450 (N_3450,N_2864,N_2357);
xnor U3451 (N_3451,N_2289,N_2503);
nor U3452 (N_3452,N_2523,N_2455);
xor U3453 (N_3453,N_2408,N_2767);
nand U3454 (N_3454,N_2965,N_2893);
xnor U3455 (N_3455,N_2790,N_2141);
nor U3456 (N_3456,N_2515,N_2210);
and U3457 (N_3457,N_2010,N_2352);
or U3458 (N_3458,N_2969,N_2810);
or U3459 (N_3459,N_2550,N_2912);
and U3460 (N_3460,N_2923,N_2041);
nor U3461 (N_3461,N_2906,N_2188);
xnor U3462 (N_3462,N_2934,N_2951);
and U3463 (N_3463,N_2203,N_2697);
or U3464 (N_3464,N_2806,N_2798);
nor U3465 (N_3465,N_2814,N_2758);
or U3466 (N_3466,N_2177,N_2020);
xor U3467 (N_3467,N_2673,N_2919);
nand U3468 (N_3468,N_2766,N_2980);
or U3469 (N_3469,N_2695,N_2292);
nand U3470 (N_3470,N_2048,N_2752);
xor U3471 (N_3471,N_2220,N_2840);
nand U3472 (N_3472,N_2560,N_2693);
and U3473 (N_3473,N_2579,N_2597);
nor U3474 (N_3474,N_2267,N_2060);
nor U3475 (N_3475,N_2495,N_2274);
xor U3476 (N_3476,N_2343,N_2689);
and U3477 (N_3477,N_2330,N_2691);
or U3478 (N_3478,N_2198,N_2652);
xor U3479 (N_3479,N_2461,N_2112);
nand U3480 (N_3480,N_2479,N_2201);
xnor U3481 (N_3481,N_2369,N_2842);
nor U3482 (N_3482,N_2588,N_2933);
and U3483 (N_3483,N_2577,N_2268);
nor U3484 (N_3484,N_2732,N_2182);
nand U3485 (N_3485,N_2088,N_2862);
nor U3486 (N_3486,N_2981,N_2045);
and U3487 (N_3487,N_2157,N_2033);
or U3488 (N_3488,N_2568,N_2681);
nor U3489 (N_3489,N_2784,N_2005);
xor U3490 (N_3490,N_2616,N_2773);
nor U3491 (N_3491,N_2393,N_2468);
nand U3492 (N_3492,N_2587,N_2260);
xnor U3493 (N_3493,N_2540,N_2240);
nand U3494 (N_3494,N_2388,N_2415);
xnor U3495 (N_3495,N_2469,N_2313);
xor U3496 (N_3496,N_2006,N_2848);
or U3497 (N_3497,N_2849,N_2081);
and U3498 (N_3498,N_2425,N_2104);
nand U3499 (N_3499,N_2952,N_2139);
nand U3500 (N_3500,N_2289,N_2104);
xor U3501 (N_3501,N_2705,N_2101);
nand U3502 (N_3502,N_2103,N_2093);
and U3503 (N_3503,N_2929,N_2065);
or U3504 (N_3504,N_2631,N_2927);
nor U3505 (N_3505,N_2957,N_2794);
nand U3506 (N_3506,N_2096,N_2239);
xnor U3507 (N_3507,N_2852,N_2730);
xnor U3508 (N_3508,N_2460,N_2393);
xor U3509 (N_3509,N_2574,N_2978);
or U3510 (N_3510,N_2769,N_2757);
or U3511 (N_3511,N_2178,N_2475);
nor U3512 (N_3512,N_2738,N_2388);
or U3513 (N_3513,N_2328,N_2196);
nand U3514 (N_3514,N_2955,N_2653);
and U3515 (N_3515,N_2783,N_2153);
xor U3516 (N_3516,N_2945,N_2395);
nor U3517 (N_3517,N_2197,N_2042);
nor U3518 (N_3518,N_2991,N_2160);
nor U3519 (N_3519,N_2039,N_2299);
nand U3520 (N_3520,N_2810,N_2033);
xnor U3521 (N_3521,N_2091,N_2082);
nor U3522 (N_3522,N_2165,N_2790);
nor U3523 (N_3523,N_2618,N_2411);
or U3524 (N_3524,N_2747,N_2533);
nand U3525 (N_3525,N_2933,N_2048);
nand U3526 (N_3526,N_2913,N_2865);
xor U3527 (N_3527,N_2556,N_2939);
and U3528 (N_3528,N_2448,N_2081);
xnor U3529 (N_3529,N_2794,N_2335);
or U3530 (N_3530,N_2836,N_2092);
nor U3531 (N_3531,N_2704,N_2602);
and U3532 (N_3532,N_2234,N_2681);
xnor U3533 (N_3533,N_2480,N_2584);
xnor U3534 (N_3534,N_2917,N_2802);
nor U3535 (N_3535,N_2020,N_2305);
and U3536 (N_3536,N_2727,N_2480);
or U3537 (N_3537,N_2835,N_2061);
nor U3538 (N_3538,N_2925,N_2079);
nor U3539 (N_3539,N_2480,N_2469);
xor U3540 (N_3540,N_2360,N_2130);
xor U3541 (N_3541,N_2751,N_2595);
and U3542 (N_3542,N_2421,N_2083);
xnor U3543 (N_3543,N_2126,N_2072);
xor U3544 (N_3544,N_2433,N_2081);
and U3545 (N_3545,N_2216,N_2089);
nor U3546 (N_3546,N_2271,N_2910);
xor U3547 (N_3547,N_2015,N_2685);
nor U3548 (N_3548,N_2598,N_2696);
nor U3549 (N_3549,N_2753,N_2356);
or U3550 (N_3550,N_2934,N_2939);
xnor U3551 (N_3551,N_2668,N_2971);
nor U3552 (N_3552,N_2528,N_2174);
nand U3553 (N_3553,N_2051,N_2267);
xnor U3554 (N_3554,N_2983,N_2192);
xor U3555 (N_3555,N_2496,N_2209);
and U3556 (N_3556,N_2269,N_2847);
nor U3557 (N_3557,N_2454,N_2858);
or U3558 (N_3558,N_2102,N_2992);
nand U3559 (N_3559,N_2174,N_2801);
xnor U3560 (N_3560,N_2890,N_2154);
nand U3561 (N_3561,N_2973,N_2855);
nand U3562 (N_3562,N_2768,N_2382);
nand U3563 (N_3563,N_2123,N_2021);
xnor U3564 (N_3564,N_2687,N_2912);
or U3565 (N_3565,N_2186,N_2840);
or U3566 (N_3566,N_2037,N_2870);
xor U3567 (N_3567,N_2134,N_2595);
xnor U3568 (N_3568,N_2370,N_2936);
nor U3569 (N_3569,N_2508,N_2123);
nand U3570 (N_3570,N_2476,N_2623);
nand U3571 (N_3571,N_2175,N_2515);
or U3572 (N_3572,N_2220,N_2207);
and U3573 (N_3573,N_2110,N_2670);
nor U3574 (N_3574,N_2789,N_2878);
nand U3575 (N_3575,N_2949,N_2261);
nor U3576 (N_3576,N_2259,N_2084);
and U3577 (N_3577,N_2793,N_2612);
nor U3578 (N_3578,N_2150,N_2940);
nand U3579 (N_3579,N_2969,N_2451);
nand U3580 (N_3580,N_2131,N_2673);
nand U3581 (N_3581,N_2920,N_2529);
xor U3582 (N_3582,N_2293,N_2450);
nand U3583 (N_3583,N_2738,N_2786);
nor U3584 (N_3584,N_2712,N_2496);
xnor U3585 (N_3585,N_2589,N_2077);
nor U3586 (N_3586,N_2966,N_2987);
and U3587 (N_3587,N_2641,N_2936);
or U3588 (N_3588,N_2259,N_2867);
or U3589 (N_3589,N_2288,N_2703);
or U3590 (N_3590,N_2409,N_2267);
nor U3591 (N_3591,N_2823,N_2332);
or U3592 (N_3592,N_2504,N_2913);
xor U3593 (N_3593,N_2513,N_2435);
or U3594 (N_3594,N_2012,N_2667);
xor U3595 (N_3595,N_2876,N_2114);
nor U3596 (N_3596,N_2570,N_2297);
nor U3597 (N_3597,N_2614,N_2632);
nor U3598 (N_3598,N_2421,N_2954);
xnor U3599 (N_3599,N_2517,N_2113);
and U3600 (N_3600,N_2276,N_2881);
nand U3601 (N_3601,N_2089,N_2221);
xor U3602 (N_3602,N_2164,N_2368);
nand U3603 (N_3603,N_2039,N_2408);
xor U3604 (N_3604,N_2942,N_2623);
xnor U3605 (N_3605,N_2655,N_2427);
nand U3606 (N_3606,N_2124,N_2893);
or U3607 (N_3607,N_2837,N_2700);
and U3608 (N_3608,N_2309,N_2065);
and U3609 (N_3609,N_2134,N_2905);
xor U3610 (N_3610,N_2869,N_2835);
nor U3611 (N_3611,N_2837,N_2720);
and U3612 (N_3612,N_2567,N_2203);
and U3613 (N_3613,N_2890,N_2250);
xor U3614 (N_3614,N_2364,N_2534);
xor U3615 (N_3615,N_2615,N_2419);
and U3616 (N_3616,N_2057,N_2736);
or U3617 (N_3617,N_2418,N_2335);
xnor U3618 (N_3618,N_2933,N_2091);
nand U3619 (N_3619,N_2811,N_2072);
or U3620 (N_3620,N_2226,N_2089);
and U3621 (N_3621,N_2957,N_2591);
xor U3622 (N_3622,N_2215,N_2289);
nor U3623 (N_3623,N_2321,N_2964);
xor U3624 (N_3624,N_2629,N_2918);
xnor U3625 (N_3625,N_2663,N_2512);
and U3626 (N_3626,N_2808,N_2700);
xnor U3627 (N_3627,N_2641,N_2544);
and U3628 (N_3628,N_2052,N_2282);
and U3629 (N_3629,N_2758,N_2170);
nand U3630 (N_3630,N_2697,N_2923);
or U3631 (N_3631,N_2256,N_2786);
nand U3632 (N_3632,N_2185,N_2776);
xnor U3633 (N_3633,N_2646,N_2254);
xnor U3634 (N_3634,N_2984,N_2123);
or U3635 (N_3635,N_2072,N_2565);
xnor U3636 (N_3636,N_2363,N_2747);
nand U3637 (N_3637,N_2195,N_2731);
and U3638 (N_3638,N_2455,N_2535);
xor U3639 (N_3639,N_2095,N_2352);
or U3640 (N_3640,N_2227,N_2525);
and U3641 (N_3641,N_2384,N_2432);
and U3642 (N_3642,N_2354,N_2997);
xnor U3643 (N_3643,N_2808,N_2189);
xnor U3644 (N_3644,N_2193,N_2709);
xnor U3645 (N_3645,N_2925,N_2088);
xnor U3646 (N_3646,N_2310,N_2540);
nand U3647 (N_3647,N_2383,N_2257);
nor U3648 (N_3648,N_2616,N_2111);
xnor U3649 (N_3649,N_2612,N_2976);
or U3650 (N_3650,N_2524,N_2503);
nor U3651 (N_3651,N_2985,N_2299);
or U3652 (N_3652,N_2721,N_2457);
or U3653 (N_3653,N_2312,N_2537);
nand U3654 (N_3654,N_2701,N_2446);
nand U3655 (N_3655,N_2834,N_2607);
and U3656 (N_3656,N_2540,N_2197);
nand U3657 (N_3657,N_2301,N_2829);
and U3658 (N_3658,N_2327,N_2309);
and U3659 (N_3659,N_2288,N_2777);
nand U3660 (N_3660,N_2005,N_2543);
nor U3661 (N_3661,N_2427,N_2051);
xor U3662 (N_3662,N_2283,N_2224);
nand U3663 (N_3663,N_2312,N_2496);
and U3664 (N_3664,N_2160,N_2344);
xor U3665 (N_3665,N_2272,N_2827);
and U3666 (N_3666,N_2969,N_2577);
or U3667 (N_3667,N_2941,N_2723);
and U3668 (N_3668,N_2527,N_2178);
or U3669 (N_3669,N_2212,N_2838);
and U3670 (N_3670,N_2420,N_2008);
or U3671 (N_3671,N_2941,N_2086);
or U3672 (N_3672,N_2949,N_2977);
nand U3673 (N_3673,N_2031,N_2423);
nand U3674 (N_3674,N_2359,N_2685);
nor U3675 (N_3675,N_2533,N_2728);
or U3676 (N_3676,N_2156,N_2850);
nand U3677 (N_3677,N_2065,N_2621);
xnor U3678 (N_3678,N_2103,N_2648);
or U3679 (N_3679,N_2973,N_2918);
nand U3680 (N_3680,N_2581,N_2213);
xor U3681 (N_3681,N_2794,N_2915);
and U3682 (N_3682,N_2225,N_2547);
xor U3683 (N_3683,N_2565,N_2150);
nand U3684 (N_3684,N_2103,N_2071);
xor U3685 (N_3685,N_2981,N_2638);
nand U3686 (N_3686,N_2113,N_2278);
xnor U3687 (N_3687,N_2027,N_2278);
nor U3688 (N_3688,N_2847,N_2226);
or U3689 (N_3689,N_2909,N_2735);
nor U3690 (N_3690,N_2706,N_2530);
xor U3691 (N_3691,N_2988,N_2089);
or U3692 (N_3692,N_2420,N_2662);
and U3693 (N_3693,N_2979,N_2252);
or U3694 (N_3694,N_2632,N_2322);
nand U3695 (N_3695,N_2445,N_2791);
nor U3696 (N_3696,N_2250,N_2856);
nor U3697 (N_3697,N_2069,N_2419);
xor U3698 (N_3698,N_2870,N_2876);
and U3699 (N_3699,N_2970,N_2641);
xor U3700 (N_3700,N_2046,N_2296);
nor U3701 (N_3701,N_2426,N_2812);
nor U3702 (N_3702,N_2840,N_2534);
nor U3703 (N_3703,N_2133,N_2832);
or U3704 (N_3704,N_2807,N_2275);
xnor U3705 (N_3705,N_2805,N_2046);
or U3706 (N_3706,N_2479,N_2388);
nor U3707 (N_3707,N_2744,N_2341);
xor U3708 (N_3708,N_2547,N_2721);
nor U3709 (N_3709,N_2411,N_2434);
or U3710 (N_3710,N_2736,N_2082);
nand U3711 (N_3711,N_2186,N_2473);
xnor U3712 (N_3712,N_2362,N_2237);
nor U3713 (N_3713,N_2436,N_2941);
or U3714 (N_3714,N_2288,N_2937);
or U3715 (N_3715,N_2553,N_2378);
or U3716 (N_3716,N_2204,N_2858);
xor U3717 (N_3717,N_2281,N_2219);
nand U3718 (N_3718,N_2652,N_2840);
xnor U3719 (N_3719,N_2331,N_2186);
or U3720 (N_3720,N_2233,N_2016);
and U3721 (N_3721,N_2217,N_2961);
xnor U3722 (N_3722,N_2191,N_2762);
xor U3723 (N_3723,N_2470,N_2628);
or U3724 (N_3724,N_2545,N_2689);
and U3725 (N_3725,N_2923,N_2609);
and U3726 (N_3726,N_2174,N_2718);
or U3727 (N_3727,N_2839,N_2105);
nor U3728 (N_3728,N_2177,N_2120);
nor U3729 (N_3729,N_2587,N_2707);
and U3730 (N_3730,N_2184,N_2898);
or U3731 (N_3731,N_2825,N_2117);
or U3732 (N_3732,N_2103,N_2007);
or U3733 (N_3733,N_2139,N_2376);
nand U3734 (N_3734,N_2710,N_2985);
nor U3735 (N_3735,N_2117,N_2938);
and U3736 (N_3736,N_2715,N_2101);
nand U3737 (N_3737,N_2979,N_2917);
xor U3738 (N_3738,N_2034,N_2506);
xor U3739 (N_3739,N_2733,N_2009);
or U3740 (N_3740,N_2343,N_2003);
and U3741 (N_3741,N_2759,N_2989);
or U3742 (N_3742,N_2886,N_2316);
nand U3743 (N_3743,N_2077,N_2437);
and U3744 (N_3744,N_2479,N_2636);
nor U3745 (N_3745,N_2233,N_2957);
nor U3746 (N_3746,N_2329,N_2885);
xnor U3747 (N_3747,N_2216,N_2882);
and U3748 (N_3748,N_2327,N_2354);
nor U3749 (N_3749,N_2513,N_2815);
or U3750 (N_3750,N_2869,N_2042);
nand U3751 (N_3751,N_2000,N_2647);
nand U3752 (N_3752,N_2945,N_2674);
or U3753 (N_3753,N_2137,N_2026);
xor U3754 (N_3754,N_2295,N_2246);
or U3755 (N_3755,N_2011,N_2839);
or U3756 (N_3756,N_2010,N_2940);
or U3757 (N_3757,N_2126,N_2731);
nor U3758 (N_3758,N_2154,N_2936);
nor U3759 (N_3759,N_2294,N_2010);
and U3760 (N_3760,N_2282,N_2587);
nor U3761 (N_3761,N_2057,N_2882);
or U3762 (N_3762,N_2757,N_2626);
nand U3763 (N_3763,N_2244,N_2854);
nand U3764 (N_3764,N_2355,N_2768);
nor U3765 (N_3765,N_2056,N_2883);
nand U3766 (N_3766,N_2833,N_2626);
and U3767 (N_3767,N_2209,N_2544);
or U3768 (N_3768,N_2477,N_2908);
nand U3769 (N_3769,N_2504,N_2894);
and U3770 (N_3770,N_2950,N_2027);
nor U3771 (N_3771,N_2723,N_2286);
nand U3772 (N_3772,N_2735,N_2022);
nand U3773 (N_3773,N_2604,N_2646);
xnor U3774 (N_3774,N_2518,N_2741);
xor U3775 (N_3775,N_2983,N_2017);
xnor U3776 (N_3776,N_2631,N_2008);
xnor U3777 (N_3777,N_2167,N_2380);
xnor U3778 (N_3778,N_2809,N_2844);
or U3779 (N_3779,N_2458,N_2441);
or U3780 (N_3780,N_2501,N_2525);
nand U3781 (N_3781,N_2420,N_2298);
nor U3782 (N_3782,N_2674,N_2873);
xnor U3783 (N_3783,N_2566,N_2202);
or U3784 (N_3784,N_2548,N_2121);
xnor U3785 (N_3785,N_2019,N_2295);
and U3786 (N_3786,N_2826,N_2290);
nor U3787 (N_3787,N_2056,N_2993);
and U3788 (N_3788,N_2770,N_2708);
and U3789 (N_3789,N_2930,N_2146);
nor U3790 (N_3790,N_2253,N_2810);
xor U3791 (N_3791,N_2486,N_2753);
nor U3792 (N_3792,N_2330,N_2273);
nor U3793 (N_3793,N_2551,N_2484);
nor U3794 (N_3794,N_2319,N_2301);
nand U3795 (N_3795,N_2950,N_2781);
and U3796 (N_3796,N_2255,N_2772);
and U3797 (N_3797,N_2202,N_2099);
or U3798 (N_3798,N_2789,N_2363);
and U3799 (N_3799,N_2091,N_2565);
xor U3800 (N_3800,N_2637,N_2754);
xnor U3801 (N_3801,N_2965,N_2369);
nor U3802 (N_3802,N_2963,N_2821);
nor U3803 (N_3803,N_2962,N_2709);
and U3804 (N_3804,N_2606,N_2986);
and U3805 (N_3805,N_2662,N_2227);
nor U3806 (N_3806,N_2434,N_2042);
or U3807 (N_3807,N_2754,N_2010);
nor U3808 (N_3808,N_2330,N_2006);
xor U3809 (N_3809,N_2521,N_2840);
nor U3810 (N_3810,N_2745,N_2496);
or U3811 (N_3811,N_2958,N_2071);
nand U3812 (N_3812,N_2408,N_2488);
or U3813 (N_3813,N_2500,N_2491);
and U3814 (N_3814,N_2871,N_2935);
or U3815 (N_3815,N_2915,N_2379);
nor U3816 (N_3816,N_2565,N_2180);
nand U3817 (N_3817,N_2507,N_2085);
nand U3818 (N_3818,N_2003,N_2652);
and U3819 (N_3819,N_2450,N_2071);
nor U3820 (N_3820,N_2405,N_2162);
nor U3821 (N_3821,N_2560,N_2037);
nor U3822 (N_3822,N_2678,N_2477);
and U3823 (N_3823,N_2818,N_2115);
nand U3824 (N_3824,N_2096,N_2967);
or U3825 (N_3825,N_2288,N_2233);
nor U3826 (N_3826,N_2532,N_2798);
xnor U3827 (N_3827,N_2198,N_2777);
and U3828 (N_3828,N_2213,N_2512);
nor U3829 (N_3829,N_2201,N_2796);
xnor U3830 (N_3830,N_2489,N_2633);
or U3831 (N_3831,N_2782,N_2934);
and U3832 (N_3832,N_2009,N_2458);
or U3833 (N_3833,N_2116,N_2521);
nand U3834 (N_3834,N_2148,N_2021);
nor U3835 (N_3835,N_2398,N_2134);
nor U3836 (N_3836,N_2079,N_2586);
nor U3837 (N_3837,N_2709,N_2107);
nor U3838 (N_3838,N_2126,N_2921);
nand U3839 (N_3839,N_2278,N_2810);
nand U3840 (N_3840,N_2098,N_2328);
nor U3841 (N_3841,N_2707,N_2705);
nand U3842 (N_3842,N_2396,N_2093);
and U3843 (N_3843,N_2158,N_2737);
or U3844 (N_3844,N_2117,N_2699);
and U3845 (N_3845,N_2326,N_2190);
or U3846 (N_3846,N_2310,N_2081);
nand U3847 (N_3847,N_2962,N_2890);
nor U3848 (N_3848,N_2857,N_2218);
and U3849 (N_3849,N_2380,N_2168);
or U3850 (N_3850,N_2989,N_2590);
nor U3851 (N_3851,N_2894,N_2947);
or U3852 (N_3852,N_2720,N_2076);
xnor U3853 (N_3853,N_2575,N_2240);
nor U3854 (N_3854,N_2101,N_2345);
and U3855 (N_3855,N_2119,N_2962);
nand U3856 (N_3856,N_2543,N_2064);
nor U3857 (N_3857,N_2090,N_2520);
nand U3858 (N_3858,N_2818,N_2475);
nor U3859 (N_3859,N_2228,N_2384);
nor U3860 (N_3860,N_2996,N_2295);
or U3861 (N_3861,N_2843,N_2859);
and U3862 (N_3862,N_2351,N_2872);
xnor U3863 (N_3863,N_2975,N_2595);
xor U3864 (N_3864,N_2344,N_2850);
and U3865 (N_3865,N_2043,N_2679);
xnor U3866 (N_3866,N_2286,N_2321);
xnor U3867 (N_3867,N_2490,N_2159);
or U3868 (N_3868,N_2084,N_2764);
and U3869 (N_3869,N_2193,N_2480);
nand U3870 (N_3870,N_2736,N_2535);
nor U3871 (N_3871,N_2575,N_2105);
and U3872 (N_3872,N_2185,N_2570);
xnor U3873 (N_3873,N_2578,N_2107);
nand U3874 (N_3874,N_2944,N_2764);
xnor U3875 (N_3875,N_2021,N_2571);
and U3876 (N_3876,N_2219,N_2831);
nand U3877 (N_3877,N_2314,N_2146);
nand U3878 (N_3878,N_2313,N_2933);
xnor U3879 (N_3879,N_2676,N_2736);
nand U3880 (N_3880,N_2238,N_2086);
or U3881 (N_3881,N_2043,N_2409);
or U3882 (N_3882,N_2115,N_2382);
nor U3883 (N_3883,N_2290,N_2737);
nor U3884 (N_3884,N_2431,N_2149);
and U3885 (N_3885,N_2756,N_2041);
or U3886 (N_3886,N_2325,N_2160);
nand U3887 (N_3887,N_2825,N_2991);
nand U3888 (N_3888,N_2521,N_2510);
nor U3889 (N_3889,N_2561,N_2177);
and U3890 (N_3890,N_2797,N_2785);
and U3891 (N_3891,N_2883,N_2305);
xnor U3892 (N_3892,N_2973,N_2228);
nor U3893 (N_3893,N_2832,N_2335);
or U3894 (N_3894,N_2079,N_2617);
nand U3895 (N_3895,N_2509,N_2149);
nor U3896 (N_3896,N_2505,N_2671);
and U3897 (N_3897,N_2447,N_2433);
or U3898 (N_3898,N_2335,N_2127);
xnor U3899 (N_3899,N_2988,N_2465);
nand U3900 (N_3900,N_2513,N_2723);
nor U3901 (N_3901,N_2448,N_2696);
and U3902 (N_3902,N_2469,N_2509);
nand U3903 (N_3903,N_2184,N_2637);
nor U3904 (N_3904,N_2979,N_2525);
nor U3905 (N_3905,N_2187,N_2753);
or U3906 (N_3906,N_2963,N_2531);
nand U3907 (N_3907,N_2620,N_2293);
nor U3908 (N_3908,N_2678,N_2074);
or U3909 (N_3909,N_2785,N_2760);
nand U3910 (N_3910,N_2472,N_2310);
or U3911 (N_3911,N_2076,N_2682);
or U3912 (N_3912,N_2680,N_2218);
nor U3913 (N_3913,N_2982,N_2361);
xor U3914 (N_3914,N_2119,N_2639);
or U3915 (N_3915,N_2143,N_2521);
and U3916 (N_3916,N_2376,N_2215);
and U3917 (N_3917,N_2765,N_2925);
xnor U3918 (N_3918,N_2517,N_2779);
or U3919 (N_3919,N_2077,N_2559);
nand U3920 (N_3920,N_2130,N_2180);
nor U3921 (N_3921,N_2055,N_2238);
or U3922 (N_3922,N_2006,N_2174);
nor U3923 (N_3923,N_2255,N_2397);
xor U3924 (N_3924,N_2412,N_2410);
and U3925 (N_3925,N_2452,N_2967);
or U3926 (N_3926,N_2087,N_2931);
or U3927 (N_3927,N_2365,N_2821);
and U3928 (N_3928,N_2923,N_2316);
and U3929 (N_3929,N_2078,N_2302);
nand U3930 (N_3930,N_2402,N_2383);
nand U3931 (N_3931,N_2126,N_2949);
nor U3932 (N_3932,N_2371,N_2579);
nor U3933 (N_3933,N_2473,N_2910);
or U3934 (N_3934,N_2036,N_2199);
and U3935 (N_3935,N_2371,N_2832);
and U3936 (N_3936,N_2549,N_2755);
nor U3937 (N_3937,N_2576,N_2683);
nor U3938 (N_3938,N_2014,N_2188);
nor U3939 (N_3939,N_2307,N_2044);
or U3940 (N_3940,N_2847,N_2436);
and U3941 (N_3941,N_2337,N_2398);
and U3942 (N_3942,N_2776,N_2634);
or U3943 (N_3943,N_2448,N_2924);
xnor U3944 (N_3944,N_2712,N_2304);
nor U3945 (N_3945,N_2080,N_2802);
nor U3946 (N_3946,N_2613,N_2216);
nand U3947 (N_3947,N_2683,N_2901);
or U3948 (N_3948,N_2515,N_2189);
nand U3949 (N_3949,N_2607,N_2203);
and U3950 (N_3950,N_2460,N_2742);
nand U3951 (N_3951,N_2124,N_2778);
or U3952 (N_3952,N_2616,N_2483);
nand U3953 (N_3953,N_2658,N_2181);
and U3954 (N_3954,N_2074,N_2944);
nor U3955 (N_3955,N_2599,N_2361);
nor U3956 (N_3956,N_2380,N_2258);
nor U3957 (N_3957,N_2697,N_2572);
nor U3958 (N_3958,N_2639,N_2484);
nor U3959 (N_3959,N_2505,N_2384);
or U3960 (N_3960,N_2577,N_2556);
nand U3961 (N_3961,N_2389,N_2552);
nand U3962 (N_3962,N_2938,N_2905);
and U3963 (N_3963,N_2114,N_2002);
and U3964 (N_3964,N_2552,N_2152);
or U3965 (N_3965,N_2222,N_2705);
xor U3966 (N_3966,N_2265,N_2535);
or U3967 (N_3967,N_2689,N_2458);
nand U3968 (N_3968,N_2045,N_2940);
xnor U3969 (N_3969,N_2817,N_2769);
xor U3970 (N_3970,N_2770,N_2682);
and U3971 (N_3971,N_2591,N_2817);
xnor U3972 (N_3972,N_2210,N_2479);
or U3973 (N_3973,N_2223,N_2484);
or U3974 (N_3974,N_2546,N_2333);
xnor U3975 (N_3975,N_2735,N_2112);
nand U3976 (N_3976,N_2645,N_2922);
nand U3977 (N_3977,N_2699,N_2105);
nand U3978 (N_3978,N_2089,N_2599);
or U3979 (N_3979,N_2232,N_2683);
nor U3980 (N_3980,N_2513,N_2594);
nor U3981 (N_3981,N_2093,N_2961);
or U3982 (N_3982,N_2851,N_2765);
or U3983 (N_3983,N_2807,N_2999);
or U3984 (N_3984,N_2624,N_2206);
xor U3985 (N_3985,N_2849,N_2723);
nor U3986 (N_3986,N_2966,N_2675);
or U3987 (N_3987,N_2679,N_2298);
and U3988 (N_3988,N_2989,N_2970);
nand U3989 (N_3989,N_2114,N_2627);
nor U3990 (N_3990,N_2103,N_2067);
nor U3991 (N_3991,N_2284,N_2090);
and U3992 (N_3992,N_2719,N_2941);
xnor U3993 (N_3993,N_2570,N_2134);
nand U3994 (N_3994,N_2824,N_2110);
and U3995 (N_3995,N_2875,N_2950);
xnor U3996 (N_3996,N_2288,N_2835);
nor U3997 (N_3997,N_2887,N_2511);
or U3998 (N_3998,N_2835,N_2482);
and U3999 (N_3999,N_2353,N_2943);
xnor U4000 (N_4000,N_3104,N_3959);
and U4001 (N_4001,N_3246,N_3746);
nand U4002 (N_4002,N_3795,N_3545);
nor U4003 (N_4003,N_3972,N_3574);
or U4004 (N_4004,N_3001,N_3568);
nand U4005 (N_4005,N_3283,N_3344);
xor U4006 (N_4006,N_3306,N_3629);
and U4007 (N_4007,N_3887,N_3288);
nor U4008 (N_4008,N_3882,N_3496);
and U4009 (N_4009,N_3782,N_3880);
xor U4010 (N_4010,N_3708,N_3889);
or U4011 (N_4011,N_3093,N_3033);
or U4012 (N_4012,N_3627,N_3360);
or U4013 (N_4013,N_3830,N_3829);
xor U4014 (N_4014,N_3314,N_3244);
and U4015 (N_4015,N_3696,N_3346);
xor U4016 (N_4016,N_3162,N_3793);
xnor U4017 (N_4017,N_3113,N_3318);
and U4018 (N_4018,N_3185,N_3247);
nor U4019 (N_4019,N_3906,N_3676);
or U4020 (N_4020,N_3991,N_3564);
and U4021 (N_4021,N_3460,N_3662);
nor U4022 (N_4022,N_3119,N_3920);
nor U4023 (N_4023,N_3692,N_3488);
nor U4024 (N_4024,N_3573,N_3144);
nor U4025 (N_4025,N_3068,N_3265);
and U4026 (N_4026,N_3624,N_3058);
xor U4027 (N_4027,N_3831,N_3100);
xnor U4028 (N_4028,N_3341,N_3459);
nor U4029 (N_4029,N_3267,N_3851);
and U4030 (N_4030,N_3653,N_3383);
nand U4031 (N_4031,N_3110,N_3726);
xnor U4032 (N_4032,N_3710,N_3222);
xor U4033 (N_4033,N_3397,N_3802);
nand U4034 (N_4034,N_3857,N_3021);
nand U4035 (N_4035,N_3912,N_3027);
nand U4036 (N_4036,N_3749,N_3052);
nor U4037 (N_4037,N_3184,N_3965);
xor U4038 (N_4038,N_3720,N_3403);
and U4039 (N_4039,N_3131,N_3442);
or U4040 (N_4040,N_3492,N_3894);
and U4041 (N_4041,N_3177,N_3172);
or U4042 (N_4042,N_3481,N_3757);
nor U4043 (N_4043,N_3210,N_3217);
nand U4044 (N_4044,N_3084,N_3311);
nor U4045 (N_4045,N_3260,N_3039);
xor U4046 (N_4046,N_3159,N_3468);
and U4047 (N_4047,N_3562,N_3538);
nor U4048 (N_4048,N_3194,N_3005);
and U4049 (N_4049,N_3335,N_3097);
nor U4050 (N_4050,N_3719,N_3211);
or U4051 (N_4051,N_3425,N_3841);
or U4052 (N_4052,N_3038,N_3495);
or U4053 (N_4053,N_3284,N_3542);
or U4054 (N_4054,N_3613,N_3728);
nor U4055 (N_4055,N_3229,N_3571);
xnor U4056 (N_4056,N_3685,N_3096);
xor U4057 (N_4057,N_3953,N_3654);
or U4058 (N_4058,N_3473,N_3674);
and U4059 (N_4059,N_3839,N_3480);
nand U4060 (N_4060,N_3150,N_3598);
and U4061 (N_4061,N_3560,N_3811);
or U4062 (N_4062,N_3905,N_3242);
xnor U4063 (N_4063,N_3273,N_3255);
nor U4064 (N_4064,N_3312,N_3703);
nor U4065 (N_4065,N_3364,N_3234);
xor U4066 (N_4066,N_3069,N_3324);
nor U4067 (N_4067,N_3816,N_3704);
and U4068 (N_4068,N_3414,N_3680);
xor U4069 (N_4069,N_3171,N_3952);
nand U4070 (N_4070,N_3277,N_3075);
or U4071 (N_4071,N_3577,N_3553);
or U4072 (N_4072,N_3987,N_3569);
and U4073 (N_4073,N_3818,N_3711);
nor U4074 (N_4074,N_3020,N_3489);
and U4075 (N_4075,N_3156,N_3517);
or U4076 (N_4076,N_3715,N_3585);
xor U4077 (N_4077,N_3734,N_3541);
or U4078 (N_4078,N_3619,N_3437);
xnor U4079 (N_4079,N_3432,N_3471);
xnor U4080 (N_4080,N_3503,N_3511);
or U4081 (N_4081,N_3126,N_3633);
xnor U4082 (N_4082,N_3621,N_3589);
xor U4083 (N_4083,N_3752,N_3307);
and U4084 (N_4084,N_3165,N_3588);
nor U4085 (N_4085,N_3855,N_3048);
and U4086 (N_4086,N_3451,N_3739);
nand U4087 (N_4087,N_3901,N_3645);
nor U4088 (N_4088,N_3874,N_3607);
and U4089 (N_4089,N_3979,N_3958);
and U4090 (N_4090,N_3315,N_3865);
xor U4091 (N_4091,N_3722,N_3153);
or U4092 (N_4092,N_3103,N_3092);
and U4093 (N_4093,N_3504,N_3130);
and U4094 (N_4094,N_3008,N_3259);
nand U4095 (N_4095,N_3693,N_3561);
and U4096 (N_4096,N_3056,N_3822);
nand U4097 (N_4097,N_3984,N_3820);
and U4098 (N_4098,N_3399,N_3376);
and U4099 (N_4099,N_3407,N_3929);
and U4100 (N_4100,N_3173,N_3840);
nor U4101 (N_4101,N_3679,N_3374);
nor U4102 (N_4102,N_3155,N_3011);
nor U4103 (N_4103,N_3114,N_3934);
nand U4104 (N_4104,N_3913,N_3365);
xor U4105 (N_4105,N_3850,N_3723);
nand U4106 (N_4106,N_3799,N_3579);
or U4107 (N_4107,N_3102,N_3922);
and U4108 (N_4108,N_3189,N_3474);
or U4109 (N_4109,N_3724,N_3744);
xnor U4110 (N_4110,N_3815,N_3673);
and U4111 (N_4111,N_3866,N_3998);
nand U4112 (N_4112,N_3129,N_3237);
and U4113 (N_4113,N_3384,N_3817);
or U4114 (N_4114,N_3042,N_3493);
or U4115 (N_4115,N_3753,N_3225);
or U4116 (N_4116,N_3707,N_3532);
or U4117 (N_4117,N_3806,N_3389);
nor U4118 (N_4118,N_3978,N_3748);
and U4119 (N_4119,N_3738,N_3472);
nand U4120 (N_4120,N_3940,N_3566);
or U4121 (N_4121,N_3235,N_3651);
or U4122 (N_4122,N_3529,N_3907);
xnor U4123 (N_4123,N_3208,N_3232);
or U4124 (N_4124,N_3028,N_3256);
nor U4125 (N_4125,N_3963,N_3047);
nand U4126 (N_4126,N_3076,N_3647);
and U4127 (N_4127,N_3054,N_3132);
or U4128 (N_4128,N_3043,N_3623);
xnor U4129 (N_4129,N_3316,N_3390);
xnor U4130 (N_4130,N_3993,N_3071);
nand U4131 (N_4131,N_3226,N_3643);
nor U4132 (N_4132,N_3745,N_3550);
nand U4133 (N_4133,N_3060,N_3310);
nor U4134 (N_4134,N_3160,N_3632);
and U4135 (N_4135,N_3618,N_3982);
nand U4136 (N_4136,N_3691,N_3124);
xor U4137 (N_4137,N_3617,N_3427);
nor U4138 (N_4138,N_3911,N_3832);
or U4139 (N_4139,N_3044,N_3756);
and U4140 (N_4140,N_3123,N_3903);
xnor U4141 (N_4141,N_3608,N_3218);
xor U4142 (N_4142,N_3422,N_3995);
or U4143 (N_4143,N_3435,N_3333);
nand U4144 (N_4144,N_3438,N_3891);
and U4145 (N_4145,N_3197,N_3801);
and U4146 (N_4146,N_3385,N_3271);
nor U4147 (N_4147,N_3484,N_3781);
and U4148 (N_4148,N_3361,N_3292);
or U4149 (N_4149,N_3101,N_3309);
or U4150 (N_4150,N_3406,N_3461);
nor U4151 (N_4151,N_3849,N_3329);
nand U4152 (N_4152,N_3338,N_3078);
xor U4153 (N_4153,N_3698,N_3702);
nand U4154 (N_4154,N_3666,N_3605);
nor U4155 (N_4155,N_3603,N_3164);
and U4156 (N_4156,N_3828,N_3320);
or U4157 (N_4157,N_3559,N_3875);
nand U4158 (N_4158,N_3766,N_3649);
and U4159 (N_4159,N_3732,N_3419);
nor U4160 (N_4160,N_3371,N_3721);
and U4161 (N_4161,N_3506,N_3883);
and U4162 (N_4162,N_3678,N_3771);
or U4163 (N_4163,N_3475,N_3441);
or U4164 (N_4164,N_3548,N_3227);
nand U4165 (N_4165,N_3467,N_3899);
and U4166 (N_4166,N_3445,N_3367);
nand U4167 (N_4167,N_3423,N_3876);
xor U4168 (N_4168,N_3926,N_3928);
nand U4169 (N_4169,N_3400,N_3392);
nor U4170 (N_4170,N_3668,N_3956);
nor U4171 (N_4171,N_3885,N_3090);
nand U4172 (N_4172,N_3622,N_3764);
or U4173 (N_4173,N_3712,N_3515);
nor U4174 (N_4174,N_3366,N_3526);
nor U4175 (N_4175,N_3688,N_3148);
xor U4176 (N_4176,N_3513,N_3729);
xor U4177 (N_4177,N_3302,N_3943);
nor U4178 (N_4178,N_3699,N_3951);
nor U4179 (N_4179,N_3250,N_3626);
or U4180 (N_4180,N_3827,N_3188);
xor U4181 (N_4181,N_3682,N_3375);
nand U4182 (N_4182,N_3490,N_3199);
nor U4183 (N_4183,N_3193,N_3594);
xor U4184 (N_4184,N_3558,N_3181);
and U4185 (N_4185,N_3740,N_3836);
and U4186 (N_4186,N_3677,N_3105);
xnor U4187 (N_4187,N_3456,N_3258);
nand U4188 (N_4188,N_3700,N_3631);
nor U4189 (N_4189,N_3733,N_3362);
nand U4190 (N_4190,N_3287,N_3486);
and U4191 (N_4191,N_3294,N_3847);
or U4192 (N_4192,N_3767,N_3863);
nand U4193 (N_4193,N_3270,N_3285);
or U4194 (N_4194,N_3025,N_3833);
or U4195 (N_4195,N_3636,N_3040);
nor U4196 (N_4196,N_3635,N_3578);
or U4197 (N_4197,N_3557,N_3821);
and U4198 (N_4198,N_3154,N_3379);
nor U4199 (N_4199,N_3029,N_3862);
xor U4200 (N_4200,N_3522,N_3118);
nor U4201 (N_4201,N_3669,N_3494);
nor U4202 (N_4202,N_3814,N_3773);
nor U4203 (N_4203,N_3602,N_3228);
nor U4204 (N_4204,N_3336,N_3004);
or U4205 (N_4205,N_3971,N_3465);
nor U4206 (N_4206,N_3168,N_3945);
xnor U4207 (N_4207,N_3931,N_3440);
xor U4208 (N_4208,N_3786,N_3634);
nand U4209 (N_4209,N_3937,N_3140);
or U4210 (N_4210,N_3002,N_3378);
nand U4211 (N_4211,N_3599,N_3293);
and U4212 (N_4212,N_3065,N_3051);
nor U4213 (N_4213,N_3055,N_3094);
xnor U4214 (N_4214,N_3418,N_3053);
and U4215 (N_4215,N_3994,N_3800);
nor U4216 (N_4216,N_3582,N_3415);
xor U4217 (N_4217,N_3923,N_3339);
and U4218 (N_4218,N_3334,N_3252);
xor U4219 (N_4219,N_3737,N_3133);
nor U4220 (N_4220,N_3368,N_3347);
nand U4221 (N_4221,N_3176,N_3448);
and U4222 (N_4222,N_3884,N_3463);
and U4223 (N_4223,N_3637,N_3409);
nor U4224 (N_4224,N_3290,N_3031);
or U4225 (N_4225,N_3308,N_3508);
or U4226 (N_4226,N_3661,N_3567);
or U4227 (N_4227,N_3837,N_3416);
nor U4228 (N_4228,N_3591,N_3067);
nor U4229 (N_4229,N_3219,N_3135);
xor U4230 (N_4230,N_3037,N_3996);
or U4231 (N_4231,N_3000,N_3041);
and U4232 (N_4232,N_3079,N_3596);
or U4233 (N_4233,N_3879,N_3877);
or U4234 (N_4234,N_3300,N_3650);
xnor U4235 (N_4235,N_3032,N_3981);
nor U4236 (N_4236,N_3547,N_3554);
nand U4237 (N_4237,N_3396,N_3202);
nand U4238 (N_4238,N_3892,N_3112);
nand U4239 (N_4239,N_3278,N_3625);
xor U4240 (N_4240,N_3439,N_3083);
nor U4241 (N_4241,N_3600,N_3136);
or U4242 (N_4242,N_3803,N_3867);
nand U4243 (N_4243,N_3961,N_3015);
and U4244 (N_4244,N_3976,N_3291);
nor U4245 (N_4245,N_3022,N_3340);
nand U4246 (N_4246,N_3754,N_3759);
and U4247 (N_4247,N_3487,N_3497);
nand U4248 (N_4248,N_3245,N_3147);
nand U4249 (N_4249,N_3797,N_3269);
nor U4250 (N_4250,N_3717,N_3500);
or U4251 (N_4251,N_3174,N_3016);
xnor U4252 (N_4252,N_3747,N_3659);
and U4253 (N_4253,N_3687,N_3763);
nor U4254 (N_4254,N_3412,N_3281);
and U4255 (N_4255,N_3443,N_3476);
and U4256 (N_4256,N_3706,N_3109);
nand U4257 (N_4257,N_3939,N_3483);
and U4258 (N_4258,N_3580,N_3531);
nor U4259 (N_4259,N_3718,N_3337);
or U4260 (N_4260,N_3854,N_3466);
nand U4261 (N_4261,N_3904,N_3207);
or U4262 (N_4262,N_3977,N_3220);
or U4263 (N_4263,N_3684,N_3354);
nand U4264 (N_4264,N_3825,N_3784);
nor U4265 (N_4265,N_3804,N_3452);
xnor U4266 (N_4266,N_3145,N_3236);
xnor U4267 (N_4267,N_3070,N_3421);
nor U4268 (N_4268,N_3238,N_3498);
nand U4269 (N_4269,N_3914,N_3611);
nand U4270 (N_4270,N_3358,N_3380);
xor U4271 (N_4271,N_3970,N_3697);
and U4272 (N_4272,N_3186,N_3356);
nor U4273 (N_4273,N_3158,N_3127);
nor U4274 (N_4274,N_3248,N_3587);
xor U4275 (N_4275,N_3464,N_3775);
nand U4276 (N_4276,N_3122,N_3080);
and U4277 (N_4277,N_3012,N_3897);
or U4278 (N_4278,N_3507,N_3166);
nand U4279 (N_4279,N_3985,N_3597);
nor U4280 (N_4280,N_3295,N_3974);
nor U4281 (N_4281,N_3410,N_3019);
xor U4282 (N_4282,N_3231,N_3064);
nand U4283 (N_4283,N_3790,N_3402);
nor U4284 (N_4284,N_3592,N_3167);
xnor U4285 (N_4285,N_3233,N_3206);
nor U4286 (N_4286,N_3555,N_3537);
or U4287 (N_4287,N_3642,N_3809);
and U4288 (N_4288,N_3570,N_3652);
xnor U4289 (N_4289,N_3139,N_3180);
xnor U4290 (N_4290,N_3453,N_3686);
or U4291 (N_4291,N_3683,N_3387);
or U4292 (N_4292,N_3896,N_3462);
or U4293 (N_4293,N_3735,N_3968);
nor U4294 (N_4294,N_3915,N_3111);
nand U4295 (N_4295,N_3013,N_3469);
nor U4296 (N_4296,N_3405,N_3581);
or U4297 (N_4297,N_3216,N_3152);
nor U4298 (N_4298,N_3411,N_3482);
nor U4299 (N_4299,N_3089,N_3325);
or U4300 (N_4300,N_3736,N_3321);
nand U4301 (N_4301,N_3116,N_3108);
and U4302 (N_4302,N_3230,N_3796);
and U4303 (N_4303,N_3485,N_3343);
nand U4304 (N_4304,N_3030,N_3919);
nor U4305 (N_4305,N_3964,N_3794);
or U4306 (N_4306,N_3878,N_3169);
and U4307 (N_4307,N_3099,N_3434);
and U4308 (N_4308,N_3224,N_3552);
nand U4309 (N_4309,N_3212,N_3137);
nor U4310 (N_4310,N_3835,N_3656);
and U4311 (N_4311,N_3727,N_3813);
nand U4312 (N_4312,N_3433,N_3351);
or U4313 (N_4313,N_3916,N_3115);
xnor U4314 (N_4314,N_3446,N_3536);
or U4315 (N_4315,N_3017,N_3762);
nand U4316 (N_4316,N_3296,N_3950);
and U4317 (N_4317,N_3125,N_3253);
and U4318 (N_4318,N_3264,N_3997);
xor U4319 (N_4319,N_3936,N_3755);
nand U4320 (N_4320,N_3450,N_3539);
and U4321 (N_4321,N_3516,N_3195);
xnor U4322 (N_4322,N_3774,N_3898);
nor U4323 (N_4323,N_3860,N_3436);
or U4324 (N_4324,N_3812,N_3563);
xor U4325 (N_4325,N_3644,N_3275);
xnor U4326 (N_4326,N_3332,N_3785);
or U4327 (N_4327,N_3714,N_3163);
or U4328 (N_4328,N_3886,N_3518);
or U4329 (N_4329,N_3063,N_3298);
nor U4330 (N_4330,N_3888,N_3908);
or U4331 (N_4331,N_3944,N_3120);
or U4332 (N_4332,N_3930,N_3061);
xor U4333 (N_4333,N_3535,N_3282);
xor U4334 (N_4334,N_3593,N_3823);
nand U4335 (N_4335,N_3671,N_3470);
xnor U4336 (N_4336,N_3612,N_3454);
and U4337 (N_4337,N_3525,N_3969);
and U4338 (N_4338,N_3792,N_3086);
nand U4339 (N_4339,N_3778,N_3190);
xnor U4340 (N_4340,N_3609,N_3861);
nand U4341 (N_4341,N_3352,N_3741);
nor U4342 (N_4342,N_3575,N_3192);
nand U4343 (N_4343,N_3512,N_3777);
or U4344 (N_4344,N_3509,N_3938);
and U4345 (N_4345,N_3765,N_3059);
xor U4346 (N_4346,N_3447,N_3357);
nor U4347 (N_4347,N_3657,N_3750);
nor U4348 (N_4348,N_3276,N_3946);
and U4349 (N_4349,N_3121,N_3890);
and U4350 (N_4350,N_3606,N_3838);
xor U4351 (N_4351,N_3009,N_3909);
and U4352 (N_4352,N_3957,N_3942);
nor U4353 (N_4353,N_3204,N_3858);
nand U4354 (N_4354,N_3081,N_3791);
xnor U4355 (N_4355,N_3313,N_3955);
nand U4356 (N_4356,N_3342,N_3393);
nand U4357 (N_4357,N_3254,N_3690);
or U4358 (N_4358,N_3262,N_3455);
or U4359 (N_4359,N_3085,N_3664);
nor U4360 (N_4360,N_3370,N_3864);
nor U4361 (N_4361,N_3299,N_3694);
and U4362 (N_4362,N_3667,N_3304);
or U4363 (N_4363,N_3209,N_3117);
nor U4364 (N_4364,N_3034,N_3758);
nor U4365 (N_4365,N_3725,N_3305);
and U4366 (N_4366,N_3221,N_3932);
xnor U4367 (N_4367,N_3353,N_3014);
nand U4368 (N_4368,N_3243,N_3491);
xnor U4369 (N_4369,N_3134,N_3280);
nand U4370 (N_4370,N_3395,N_3091);
xnor U4371 (N_4371,N_3615,N_3429);
xor U4372 (N_4372,N_3268,N_3035);
xnor U4373 (N_4373,N_3373,N_3331);
nand U4374 (N_4374,N_3178,N_3322);
nand U4375 (N_4375,N_3363,N_3533);
nor U4376 (N_4376,N_3869,N_3372);
nand U4377 (N_4377,N_3297,N_3730);
nor U4378 (N_4378,N_3917,N_3431);
and U4379 (N_4379,N_3323,N_3983);
and U4380 (N_4380,N_3326,N_3772);
and U4381 (N_4381,N_3933,N_3106);
nor U4382 (N_4382,N_3523,N_3924);
xor U4383 (N_4383,N_3805,N_3143);
nor U4384 (N_4384,N_3595,N_3910);
xnor U4385 (N_4385,N_3583,N_3408);
and U4386 (N_4386,N_3214,N_3641);
xor U4387 (N_4387,N_3330,N_3263);
and U4388 (N_4388,N_3842,N_3973);
nand U4389 (N_4389,N_3941,N_3731);
xor U4390 (N_4390,N_3544,N_3935);
nor U4391 (N_4391,N_3798,N_3648);
xor U4392 (N_4392,N_3388,N_3239);
or U4393 (N_4393,N_3141,N_3881);
or U4394 (N_4394,N_3279,N_3179);
nor U4395 (N_4395,N_3528,N_3382);
nand U4396 (N_4396,N_3992,N_3925);
xor U4397 (N_4397,N_3424,N_3045);
or U4398 (N_4398,N_3203,N_3317);
or U4399 (N_4399,N_3066,N_3191);
nor U4400 (N_4400,N_3426,N_3843);
nor U4401 (N_4401,N_3663,N_3534);
nor U4402 (N_4402,N_3665,N_3272);
and U4403 (N_4403,N_3182,N_3157);
nor U4404 (N_4404,N_3074,N_3675);
nand U4405 (N_4405,N_3499,N_3527);
nor U4406 (N_4406,N_3660,N_3010);
nand U4407 (N_4407,N_3986,N_3989);
nor U4408 (N_4408,N_3848,N_3640);
xor U4409 (N_4409,N_3921,N_3026);
and U4410 (N_4410,N_3601,N_3543);
xnor U4411 (N_4411,N_3709,N_3701);
and U4412 (N_4412,N_3369,N_3565);
xor U4413 (N_4413,N_3057,N_3240);
or U4414 (N_4414,N_3689,N_3128);
or U4415 (N_4415,N_3266,N_3834);
nand U4416 (N_4416,N_3810,N_3151);
xor U4417 (N_4417,N_3988,N_3824);
nand U4418 (N_4418,N_3519,N_3681);
nor U4419 (N_4419,N_3576,N_3510);
nand U4420 (N_4420,N_3457,N_3003);
and U4421 (N_4421,N_3514,N_3458);
or U4422 (N_4422,N_3398,N_3551);
or U4423 (N_4423,N_3107,N_3349);
xor U4424 (N_4424,N_3853,N_3530);
nor U4425 (N_4425,N_3073,N_3479);
xor U4426 (N_4426,N_3018,N_3428);
nor U4427 (N_4427,N_3980,N_3359);
and U4428 (N_4428,N_3394,N_3175);
nor U4429 (N_4429,N_3819,N_3604);
nand U4430 (N_4430,N_3780,N_3949);
or U4431 (N_4431,N_3261,N_3095);
xnor U4432 (N_4432,N_3477,N_3776);
nor U4433 (N_4433,N_3807,N_3751);
nor U4434 (N_4434,N_3007,N_3873);
or U4435 (N_4435,N_3902,N_3556);
nor U4436 (N_4436,N_3161,N_3521);
and U4437 (N_4437,N_3630,N_3586);
nor U4438 (N_4438,N_3856,N_3098);
xor U4439 (N_4439,N_3761,N_3655);
or U4440 (N_4440,N_3241,N_3572);
and U4441 (N_4441,N_3350,N_3077);
or U4442 (N_4442,N_3846,N_3146);
xor U4443 (N_4443,N_3672,N_3223);
nor U4444 (N_4444,N_3670,N_3872);
and U4445 (N_4445,N_3639,N_3377);
nand U4446 (N_4446,N_3549,N_3417);
nor U4447 (N_4447,N_3501,N_3524);
and U4448 (N_4448,N_3695,N_3355);
nor U4449 (N_4449,N_3142,N_3614);
nor U4450 (N_4450,N_3546,N_3024);
xor U4451 (N_4451,N_3859,N_3960);
nand U4452 (N_4452,N_3975,N_3743);
and U4453 (N_4453,N_3844,N_3046);
nand U4454 (N_4454,N_3893,N_3900);
nand U4455 (N_4455,N_3328,N_3401);
xor U4456 (N_4456,N_3999,N_3213);
or U4457 (N_4457,N_3584,N_3947);
or U4458 (N_4458,N_3138,N_3716);
or U4459 (N_4459,N_3638,N_3620);
nor U4460 (N_4460,N_3386,N_3183);
and U4461 (N_4461,N_3062,N_3257);
xnor U4462 (N_4462,N_3478,N_3768);
nor U4463 (N_4463,N_3705,N_3072);
and U4464 (N_4464,N_3870,N_3251);
xnor U4465 (N_4465,N_3201,N_3962);
or U4466 (N_4466,N_3788,N_3215);
nand U4467 (N_4467,N_3769,N_3948);
nor U4468 (N_4468,N_3303,N_3200);
xnor U4469 (N_4469,N_3449,N_3345);
nor U4470 (N_4470,N_3187,N_3023);
xnor U4471 (N_4471,N_3196,N_3713);
nand U4472 (N_4472,N_3868,N_3616);
xor U4473 (N_4473,N_3787,N_3742);
and U4474 (N_4474,N_3520,N_3852);
and U4475 (N_4475,N_3327,N_3540);
or U4476 (N_4476,N_3954,N_3348);
and U4477 (N_4477,N_3381,N_3646);
and U4478 (N_4478,N_3301,N_3088);
nand U4479 (N_4479,N_3808,N_3170);
nor U4480 (N_4480,N_3826,N_3404);
nand U4481 (N_4481,N_3918,N_3967);
nand U4482 (N_4482,N_3087,N_3205);
or U4483 (N_4483,N_3198,N_3783);
nand U4484 (N_4484,N_3274,N_3770);
nor U4485 (N_4485,N_3628,N_3658);
nor U4486 (N_4486,N_3590,N_3789);
or U4487 (N_4487,N_3049,N_3319);
or U4488 (N_4488,N_3082,N_3289);
xor U4489 (N_4489,N_3444,N_3050);
nor U4490 (N_4490,N_3249,N_3413);
and U4491 (N_4491,N_3391,N_3505);
or U4492 (N_4492,N_3845,N_3990);
and U4493 (N_4493,N_3430,N_3610);
and U4494 (N_4494,N_3502,N_3779);
or U4495 (N_4495,N_3966,N_3286);
or U4496 (N_4496,N_3006,N_3895);
or U4497 (N_4497,N_3760,N_3149);
nand U4498 (N_4498,N_3420,N_3036);
or U4499 (N_4499,N_3871,N_3927);
and U4500 (N_4500,N_3350,N_3686);
and U4501 (N_4501,N_3828,N_3974);
and U4502 (N_4502,N_3027,N_3358);
nand U4503 (N_4503,N_3279,N_3581);
nand U4504 (N_4504,N_3284,N_3283);
nor U4505 (N_4505,N_3679,N_3654);
nand U4506 (N_4506,N_3211,N_3984);
nand U4507 (N_4507,N_3964,N_3560);
and U4508 (N_4508,N_3063,N_3041);
nand U4509 (N_4509,N_3470,N_3255);
nand U4510 (N_4510,N_3471,N_3240);
nor U4511 (N_4511,N_3294,N_3043);
or U4512 (N_4512,N_3571,N_3146);
or U4513 (N_4513,N_3691,N_3075);
nand U4514 (N_4514,N_3153,N_3214);
nand U4515 (N_4515,N_3389,N_3115);
and U4516 (N_4516,N_3464,N_3950);
nand U4517 (N_4517,N_3300,N_3770);
or U4518 (N_4518,N_3224,N_3964);
or U4519 (N_4519,N_3507,N_3086);
and U4520 (N_4520,N_3471,N_3028);
nand U4521 (N_4521,N_3601,N_3439);
xnor U4522 (N_4522,N_3983,N_3413);
or U4523 (N_4523,N_3676,N_3778);
and U4524 (N_4524,N_3422,N_3077);
nand U4525 (N_4525,N_3300,N_3625);
nor U4526 (N_4526,N_3560,N_3575);
and U4527 (N_4527,N_3045,N_3761);
nor U4528 (N_4528,N_3220,N_3839);
nand U4529 (N_4529,N_3238,N_3107);
xnor U4530 (N_4530,N_3917,N_3921);
nor U4531 (N_4531,N_3839,N_3382);
nand U4532 (N_4532,N_3559,N_3560);
nand U4533 (N_4533,N_3598,N_3040);
nand U4534 (N_4534,N_3458,N_3867);
and U4535 (N_4535,N_3548,N_3716);
xor U4536 (N_4536,N_3829,N_3533);
nand U4537 (N_4537,N_3008,N_3748);
nand U4538 (N_4538,N_3833,N_3012);
or U4539 (N_4539,N_3579,N_3548);
nand U4540 (N_4540,N_3015,N_3039);
nand U4541 (N_4541,N_3710,N_3914);
nor U4542 (N_4542,N_3934,N_3424);
xor U4543 (N_4543,N_3142,N_3170);
xor U4544 (N_4544,N_3619,N_3531);
xnor U4545 (N_4545,N_3777,N_3496);
nor U4546 (N_4546,N_3064,N_3042);
xor U4547 (N_4547,N_3132,N_3191);
nor U4548 (N_4548,N_3091,N_3587);
nand U4549 (N_4549,N_3623,N_3768);
and U4550 (N_4550,N_3597,N_3523);
xnor U4551 (N_4551,N_3851,N_3402);
and U4552 (N_4552,N_3243,N_3627);
or U4553 (N_4553,N_3030,N_3867);
nor U4554 (N_4554,N_3462,N_3213);
nand U4555 (N_4555,N_3273,N_3343);
and U4556 (N_4556,N_3588,N_3151);
or U4557 (N_4557,N_3658,N_3111);
or U4558 (N_4558,N_3168,N_3045);
and U4559 (N_4559,N_3468,N_3996);
and U4560 (N_4560,N_3081,N_3684);
nand U4561 (N_4561,N_3579,N_3665);
nor U4562 (N_4562,N_3228,N_3748);
xor U4563 (N_4563,N_3853,N_3927);
nand U4564 (N_4564,N_3111,N_3430);
xnor U4565 (N_4565,N_3637,N_3462);
or U4566 (N_4566,N_3531,N_3334);
and U4567 (N_4567,N_3068,N_3901);
nor U4568 (N_4568,N_3437,N_3298);
nor U4569 (N_4569,N_3013,N_3199);
or U4570 (N_4570,N_3099,N_3752);
and U4571 (N_4571,N_3370,N_3749);
or U4572 (N_4572,N_3162,N_3962);
xnor U4573 (N_4573,N_3515,N_3377);
and U4574 (N_4574,N_3104,N_3242);
nand U4575 (N_4575,N_3025,N_3575);
xor U4576 (N_4576,N_3796,N_3926);
nor U4577 (N_4577,N_3043,N_3502);
nor U4578 (N_4578,N_3023,N_3551);
nand U4579 (N_4579,N_3130,N_3025);
or U4580 (N_4580,N_3137,N_3528);
and U4581 (N_4581,N_3024,N_3714);
xnor U4582 (N_4582,N_3790,N_3540);
or U4583 (N_4583,N_3156,N_3400);
xnor U4584 (N_4584,N_3695,N_3027);
nand U4585 (N_4585,N_3286,N_3667);
or U4586 (N_4586,N_3431,N_3525);
nor U4587 (N_4587,N_3455,N_3673);
nand U4588 (N_4588,N_3042,N_3207);
nor U4589 (N_4589,N_3244,N_3172);
xor U4590 (N_4590,N_3061,N_3130);
nor U4591 (N_4591,N_3634,N_3817);
and U4592 (N_4592,N_3893,N_3443);
xor U4593 (N_4593,N_3826,N_3956);
or U4594 (N_4594,N_3026,N_3773);
and U4595 (N_4595,N_3360,N_3670);
nand U4596 (N_4596,N_3386,N_3439);
or U4597 (N_4597,N_3432,N_3918);
nor U4598 (N_4598,N_3807,N_3563);
nand U4599 (N_4599,N_3015,N_3122);
and U4600 (N_4600,N_3562,N_3961);
and U4601 (N_4601,N_3039,N_3189);
and U4602 (N_4602,N_3924,N_3851);
nand U4603 (N_4603,N_3342,N_3221);
nand U4604 (N_4604,N_3896,N_3546);
and U4605 (N_4605,N_3646,N_3686);
or U4606 (N_4606,N_3784,N_3049);
xnor U4607 (N_4607,N_3837,N_3386);
nor U4608 (N_4608,N_3577,N_3588);
and U4609 (N_4609,N_3333,N_3943);
xnor U4610 (N_4610,N_3544,N_3815);
xnor U4611 (N_4611,N_3085,N_3566);
nand U4612 (N_4612,N_3108,N_3085);
nor U4613 (N_4613,N_3580,N_3420);
or U4614 (N_4614,N_3950,N_3575);
or U4615 (N_4615,N_3440,N_3703);
nand U4616 (N_4616,N_3289,N_3252);
or U4617 (N_4617,N_3450,N_3537);
xnor U4618 (N_4618,N_3527,N_3112);
nor U4619 (N_4619,N_3682,N_3565);
nand U4620 (N_4620,N_3901,N_3888);
nor U4621 (N_4621,N_3620,N_3047);
or U4622 (N_4622,N_3541,N_3464);
or U4623 (N_4623,N_3304,N_3356);
and U4624 (N_4624,N_3690,N_3481);
and U4625 (N_4625,N_3097,N_3361);
nand U4626 (N_4626,N_3653,N_3472);
xnor U4627 (N_4627,N_3131,N_3258);
or U4628 (N_4628,N_3353,N_3345);
and U4629 (N_4629,N_3110,N_3819);
or U4630 (N_4630,N_3383,N_3025);
and U4631 (N_4631,N_3879,N_3080);
xor U4632 (N_4632,N_3459,N_3875);
xnor U4633 (N_4633,N_3922,N_3852);
and U4634 (N_4634,N_3923,N_3723);
or U4635 (N_4635,N_3086,N_3366);
xor U4636 (N_4636,N_3161,N_3662);
and U4637 (N_4637,N_3433,N_3122);
nor U4638 (N_4638,N_3461,N_3599);
and U4639 (N_4639,N_3603,N_3097);
nand U4640 (N_4640,N_3454,N_3892);
xnor U4641 (N_4641,N_3496,N_3656);
xnor U4642 (N_4642,N_3347,N_3185);
nor U4643 (N_4643,N_3318,N_3989);
nor U4644 (N_4644,N_3640,N_3118);
nand U4645 (N_4645,N_3659,N_3459);
xnor U4646 (N_4646,N_3853,N_3252);
nand U4647 (N_4647,N_3895,N_3231);
xnor U4648 (N_4648,N_3451,N_3962);
xnor U4649 (N_4649,N_3923,N_3759);
xnor U4650 (N_4650,N_3824,N_3746);
nand U4651 (N_4651,N_3449,N_3166);
and U4652 (N_4652,N_3020,N_3929);
xnor U4653 (N_4653,N_3664,N_3929);
and U4654 (N_4654,N_3151,N_3636);
or U4655 (N_4655,N_3098,N_3254);
nand U4656 (N_4656,N_3562,N_3315);
nor U4657 (N_4657,N_3440,N_3392);
nor U4658 (N_4658,N_3852,N_3617);
or U4659 (N_4659,N_3205,N_3653);
nor U4660 (N_4660,N_3124,N_3803);
and U4661 (N_4661,N_3728,N_3311);
xor U4662 (N_4662,N_3180,N_3521);
nand U4663 (N_4663,N_3811,N_3728);
nor U4664 (N_4664,N_3095,N_3021);
nand U4665 (N_4665,N_3592,N_3458);
and U4666 (N_4666,N_3759,N_3120);
nor U4667 (N_4667,N_3919,N_3977);
xor U4668 (N_4668,N_3381,N_3920);
and U4669 (N_4669,N_3935,N_3615);
and U4670 (N_4670,N_3811,N_3304);
or U4671 (N_4671,N_3773,N_3013);
nand U4672 (N_4672,N_3814,N_3934);
xor U4673 (N_4673,N_3890,N_3294);
and U4674 (N_4674,N_3149,N_3853);
or U4675 (N_4675,N_3891,N_3200);
nor U4676 (N_4676,N_3310,N_3938);
xnor U4677 (N_4677,N_3277,N_3221);
nand U4678 (N_4678,N_3857,N_3821);
or U4679 (N_4679,N_3911,N_3929);
nor U4680 (N_4680,N_3364,N_3194);
xor U4681 (N_4681,N_3531,N_3777);
or U4682 (N_4682,N_3448,N_3841);
nor U4683 (N_4683,N_3792,N_3772);
and U4684 (N_4684,N_3184,N_3723);
or U4685 (N_4685,N_3895,N_3371);
nand U4686 (N_4686,N_3052,N_3336);
nor U4687 (N_4687,N_3135,N_3512);
nand U4688 (N_4688,N_3435,N_3491);
nor U4689 (N_4689,N_3679,N_3903);
and U4690 (N_4690,N_3566,N_3945);
or U4691 (N_4691,N_3145,N_3455);
or U4692 (N_4692,N_3034,N_3102);
xnor U4693 (N_4693,N_3188,N_3181);
xnor U4694 (N_4694,N_3906,N_3682);
xor U4695 (N_4695,N_3890,N_3945);
and U4696 (N_4696,N_3884,N_3835);
nand U4697 (N_4697,N_3235,N_3487);
and U4698 (N_4698,N_3941,N_3879);
xor U4699 (N_4699,N_3477,N_3445);
or U4700 (N_4700,N_3330,N_3483);
or U4701 (N_4701,N_3355,N_3947);
nor U4702 (N_4702,N_3569,N_3487);
and U4703 (N_4703,N_3242,N_3195);
nand U4704 (N_4704,N_3146,N_3887);
nand U4705 (N_4705,N_3547,N_3436);
or U4706 (N_4706,N_3725,N_3592);
xor U4707 (N_4707,N_3278,N_3319);
nor U4708 (N_4708,N_3569,N_3983);
nand U4709 (N_4709,N_3740,N_3234);
and U4710 (N_4710,N_3719,N_3486);
nand U4711 (N_4711,N_3373,N_3409);
xor U4712 (N_4712,N_3228,N_3821);
nand U4713 (N_4713,N_3991,N_3982);
nand U4714 (N_4714,N_3807,N_3028);
and U4715 (N_4715,N_3931,N_3466);
and U4716 (N_4716,N_3727,N_3337);
nand U4717 (N_4717,N_3775,N_3785);
nor U4718 (N_4718,N_3758,N_3085);
nor U4719 (N_4719,N_3628,N_3193);
xnor U4720 (N_4720,N_3168,N_3260);
nor U4721 (N_4721,N_3549,N_3290);
nor U4722 (N_4722,N_3520,N_3987);
and U4723 (N_4723,N_3927,N_3608);
and U4724 (N_4724,N_3696,N_3721);
and U4725 (N_4725,N_3969,N_3450);
xor U4726 (N_4726,N_3486,N_3107);
or U4727 (N_4727,N_3084,N_3002);
nand U4728 (N_4728,N_3249,N_3140);
nor U4729 (N_4729,N_3199,N_3800);
or U4730 (N_4730,N_3782,N_3591);
or U4731 (N_4731,N_3963,N_3685);
nand U4732 (N_4732,N_3287,N_3955);
nand U4733 (N_4733,N_3107,N_3185);
xnor U4734 (N_4734,N_3789,N_3735);
or U4735 (N_4735,N_3233,N_3777);
nor U4736 (N_4736,N_3076,N_3178);
nand U4737 (N_4737,N_3279,N_3674);
nand U4738 (N_4738,N_3223,N_3011);
nor U4739 (N_4739,N_3572,N_3590);
nor U4740 (N_4740,N_3071,N_3671);
nand U4741 (N_4741,N_3646,N_3889);
nor U4742 (N_4742,N_3198,N_3164);
nand U4743 (N_4743,N_3552,N_3499);
or U4744 (N_4744,N_3992,N_3358);
nor U4745 (N_4745,N_3068,N_3994);
and U4746 (N_4746,N_3256,N_3791);
nor U4747 (N_4747,N_3353,N_3727);
and U4748 (N_4748,N_3048,N_3440);
and U4749 (N_4749,N_3284,N_3895);
nand U4750 (N_4750,N_3545,N_3459);
xor U4751 (N_4751,N_3522,N_3041);
or U4752 (N_4752,N_3664,N_3211);
xnor U4753 (N_4753,N_3518,N_3221);
nor U4754 (N_4754,N_3986,N_3010);
nor U4755 (N_4755,N_3903,N_3190);
and U4756 (N_4756,N_3506,N_3709);
xnor U4757 (N_4757,N_3284,N_3853);
xnor U4758 (N_4758,N_3349,N_3599);
nor U4759 (N_4759,N_3692,N_3524);
or U4760 (N_4760,N_3817,N_3682);
nand U4761 (N_4761,N_3960,N_3813);
nor U4762 (N_4762,N_3250,N_3255);
xor U4763 (N_4763,N_3453,N_3858);
xnor U4764 (N_4764,N_3558,N_3174);
nor U4765 (N_4765,N_3672,N_3159);
and U4766 (N_4766,N_3797,N_3465);
nand U4767 (N_4767,N_3257,N_3279);
and U4768 (N_4768,N_3491,N_3698);
nand U4769 (N_4769,N_3522,N_3411);
and U4770 (N_4770,N_3477,N_3826);
nor U4771 (N_4771,N_3292,N_3230);
xor U4772 (N_4772,N_3420,N_3494);
and U4773 (N_4773,N_3883,N_3373);
nor U4774 (N_4774,N_3442,N_3509);
nor U4775 (N_4775,N_3507,N_3486);
and U4776 (N_4776,N_3859,N_3302);
or U4777 (N_4777,N_3223,N_3177);
or U4778 (N_4778,N_3725,N_3321);
or U4779 (N_4779,N_3944,N_3097);
nand U4780 (N_4780,N_3640,N_3346);
xnor U4781 (N_4781,N_3093,N_3730);
nand U4782 (N_4782,N_3713,N_3488);
and U4783 (N_4783,N_3649,N_3506);
nor U4784 (N_4784,N_3336,N_3534);
or U4785 (N_4785,N_3581,N_3691);
or U4786 (N_4786,N_3577,N_3322);
xnor U4787 (N_4787,N_3997,N_3353);
nand U4788 (N_4788,N_3602,N_3410);
and U4789 (N_4789,N_3754,N_3652);
and U4790 (N_4790,N_3995,N_3205);
and U4791 (N_4791,N_3930,N_3171);
nand U4792 (N_4792,N_3439,N_3654);
and U4793 (N_4793,N_3719,N_3034);
nor U4794 (N_4794,N_3861,N_3413);
xor U4795 (N_4795,N_3420,N_3034);
nand U4796 (N_4796,N_3946,N_3739);
xnor U4797 (N_4797,N_3011,N_3423);
and U4798 (N_4798,N_3552,N_3811);
xor U4799 (N_4799,N_3270,N_3271);
or U4800 (N_4800,N_3695,N_3747);
nor U4801 (N_4801,N_3298,N_3882);
nor U4802 (N_4802,N_3054,N_3288);
nor U4803 (N_4803,N_3855,N_3740);
and U4804 (N_4804,N_3319,N_3149);
nand U4805 (N_4805,N_3498,N_3050);
and U4806 (N_4806,N_3904,N_3042);
nand U4807 (N_4807,N_3542,N_3136);
xor U4808 (N_4808,N_3060,N_3014);
nand U4809 (N_4809,N_3416,N_3085);
xor U4810 (N_4810,N_3207,N_3532);
and U4811 (N_4811,N_3712,N_3025);
xnor U4812 (N_4812,N_3737,N_3147);
or U4813 (N_4813,N_3357,N_3118);
nand U4814 (N_4814,N_3090,N_3634);
or U4815 (N_4815,N_3414,N_3917);
or U4816 (N_4816,N_3440,N_3442);
xor U4817 (N_4817,N_3826,N_3964);
xor U4818 (N_4818,N_3545,N_3942);
nand U4819 (N_4819,N_3725,N_3546);
xnor U4820 (N_4820,N_3064,N_3372);
nand U4821 (N_4821,N_3896,N_3541);
and U4822 (N_4822,N_3218,N_3661);
nand U4823 (N_4823,N_3414,N_3644);
and U4824 (N_4824,N_3703,N_3474);
or U4825 (N_4825,N_3254,N_3001);
and U4826 (N_4826,N_3304,N_3255);
and U4827 (N_4827,N_3401,N_3101);
or U4828 (N_4828,N_3047,N_3176);
or U4829 (N_4829,N_3721,N_3015);
nor U4830 (N_4830,N_3316,N_3670);
xnor U4831 (N_4831,N_3079,N_3500);
and U4832 (N_4832,N_3271,N_3177);
nor U4833 (N_4833,N_3182,N_3046);
xor U4834 (N_4834,N_3785,N_3753);
xor U4835 (N_4835,N_3854,N_3479);
nand U4836 (N_4836,N_3580,N_3769);
nand U4837 (N_4837,N_3749,N_3768);
nand U4838 (N_4838,N_3099,N_3486);
xnor U4839 (N_4839,N_3489,N_3646);
or U4840 (N_4840,N_3571,N_3012);
and U4841 (N_4841,N_3392,N_3056);
nand U4842 (N_4842,N_3405,N_3560);
or U4843 (N_4843,N_3907,N_3592);
nand U4844 (N_4844,N_3887,N_3155);
nor U4845 (N_4845,N_3554,N_3929);
nand U4846 (N_4846,N_3324,N_3962);
nor U4847 (N_4847,N_3439,N_3279);
nand U4848 (N_4848,N_3600,N_3908);
nor U4849 (N_4849,N_3033,N_3026);
nor U4850 (N_4850,N_3756,N_3973);
or U4851 (N_4851,N_3548,N_3385);
and U4852 (N_4852,N_3251,N_3002);
and U4853 (N_4853,N_3900,N_3035);
xnor U4854 (N_4854,N_3816,N_3534);
nor U4855 (N_4855,N_3052,N_3401);
nand U4856 (N_4856,N_3710,N_3898);
xnor U4857 (N_4857,N_3047,N_3965);
and U4858 (N_4858,N_3572,N_3608);
nand U4859 (N_4859,N_3698,N_3065);
and U4860 (N_4860,N_3208,N_3235);
nor U4861 (N_4861,N_3509,N_3868);
xnor U4862 (N_4862,N_3217,N_3061);
xor U4863 (N_4863,N_3699,N_3094);
xnor U4864 (N_4864,N_3474,N_3493);
nor U4865 (N_4865,N_3663,N_3757);
and U4866 (N_4866,N_3117,N_3384);
xor U4867 (N_4867,N_3176,N_3471);
or U4868 (N_4868,N_3455,N_3315);
xnor U4869 (N_4869,N_3101,N_3230);
xor U4870 (N_4870,N_3366,N_3113);
nand U4871 (N_4871,N_3166,N_3896);
or U4872 (N_4872,N_3545,N_3759);
xor U4873 (N_4873,N_3376,N_3121);
nor U4874 (N_4874,N_3429,N_3531);
and U4875 (N_4875,N_3648,N_3678);
nand U4876 (N_4876,N_3183,N_3692);
nor U4877 (N_4877,N_3756,N_3905);
xnor U4878 (N_4878,N_3374,N_3829);
nand U4879 (N_4879,N_3333,N_3178);
and U4880 (N_4880,N_3331,N_3317);
or U4881 (N_4881,N_3783,N_3364);
xor U4882 (N_4882,N_3078,N_3194);
and U4883 (N_4883,N_3527,N_3202);
or U4884 (N_4884,N_3713,N_3628);
nand U4885 (N_4885,N_3626,N_3542);
nor U4886 (N_4886,N_3173,N_3020);
and U4887 (N_4887,N_3056,N_3941);
or U4888 (N_4888,N_3630,N_3549);
nand U4889 (N_4889,N_3022,N_3331);
and U4890 (N_4890,N_3975,N_3550);
and U4891 (N_4891,N_3906,N_3719);
nor U4892 (N_4892,N_3200,N_3047);
nor U4893 (N_4893,N_3169,N_3910);
and U4894 (N_4894,N_3786,N_3368);
and U4895 (N_4895,N_3989,N_3773);
or U4896 (N_4896,N_3670,N_3046);
nor U4897 (N_4897,N_3094,N_3276);
nor U4898 (N_4898,N_3289,N_3114);
nor U4899 (N_4899,N_3182,N_3641);
xor U4900 (N_4900,N_3694,N_3627);
xor U4901 (N_4901,N_3872,N_3312);
nor U4902 (N_4902,N_3585,N_3184);
or U4903 (N_4903,N_3773,N_3212);
or U4904 (N_4904,N_3383,N_3491);
nand U4905 (N_4905,N_3421,N_3602);
xor U4906 (N_4906,N_3534,N_3325);
or U4907 (N_4907,N_3931,N_3549);
and U4908 (N_4908,N_3354,N_3147);
or U4909 (N_4909,N_3196,N_3192);
and U4910 (N_4910,N_3352,N_3113);
nor U4911 (N_4911,N_3929,N_3731);
nor U4912 (N_4912,N_3523,N_3824);
nor U4913 (N_4913,N_3780,N_3886);
nand U4914 (N_4914,N_3891,N_3413);
nor U4915 (N_4915,N_3465,N_3887);
and U4916 (N_4916,N_3546,N_3693);
nand U4917 (N_4917,N_3713,N_3556);
nand U4918 (N_4918,N_3491,N_3852);
xnor U4919 (N_4919,N_3853,N_3012);
or U4920 (N_4920,N_3706,N_3221);
and U4921 (N_4921,N_3923,N_3018);
nor U4922 (N_4922,N_3090,N_3886);
or U4923 (N_4923,N_3352,N_3651);
xor U4924 (N_4924,N_3801,N_3051);
xnor U4925 (N_4925,N_3927,N_3781);
or U4926 (N_4926,N_3898,N_3754);
nor U4927 (N_4927,N_3578,N_3177);
xor U4928 (N_4928,N_3416,N_3683);
nor U4929 (N_4929,N_3151,N_3976);
nand U4930 (N_4930,N_3277,N_3955);
xor U4931 (N_4931,N_3946,N_3428);
nand U4932 (N_4932,N_3119,N_3292);
or U4933 (N_4933,N_3981,N_3932);
and U4934 (N_4934,N_3944,N_3767);
xnor U4935 (N_4935,N_3511,N_3887);
nand U4936 (N_4936,N_3932,N_3728);
nor U4937 (N_4937,N_3894,N_3741);
nor U4938 (N_4938,N_3461,N_3939);
xor U4939 (N_4939,N_3665,N_3685);
nand U4940 (N_4940,N_3673,N_3924);
and U4941 (N_4941,N_3086,N_3261);
and U4942 (N_4942,N_3529,N_3240);
or U4943 (N_4943,N_3481,N_3498);
xor U4944 (N_4944,N_3386,N_3112);
nor U4945 (N_4945,N_3330,N_3640);
nor U4946 (N_4946,N_3206,N_3804);
nand U4947 (N_4947,N_3073,N_3546);
or U4948 (N_4948,N_3468,N_3265);
and U4949 (N_4949,N_3150,N_3376);
or U4950 (N_4950,N_3561,N_3932);
or U4951 (N_4951,N_3676,N_3201);
xnor U4952 (N_4952,N_3143,N_3189);
nand U4953 (N_4953,N_3012,N_3467);
or U4954 (N_4954,N_3602,N_3741);
nand U4955 (N_4955,N_3649,N_3378);
or U4956 (N_4956,N_3190,N_3479);
nor U4957 (N_4957,N_3682,N_3429);
nand U4958 (N_4958,N_3165,N_3750);
nor U4959 (N_4959,N_3320,N_3175);
or U4960 (N_4960,N_3346,N_3922);
nand U4961 (N_4961,N_3153,N_3852);
nand U4962 (N_4962,N_3713,N_3254);
nand U4963 (N_4963,N_3765,N_3622);
xor U4964 (N_4964,N_3683,N_3130);
or U4965 (N_4965,N_3121,N_3721);
nor U4966 (N_4966,N_3062,N_3751);
nor U4967 (N_4967,N_3574,N_3287);
and U4968 (N_4968,N_3219,N_3495);
xnor U4969 (N_4969,N_3894,N_3864);
nand U4970 (N_4970,N_3419,N_3229);
nor U4971 (N_4971,N_3607,N_3291);
xor U4972 (N_4972,N_3270,N_3822);
xnor U4973 (N_4973,N_3921,N_3813);
nand U4974 (N_4974,N_3329,N_3795);
or U4975 (N_4975,N_3271,N_3545);
and U4976 (N_4976,N_3675,N_3716);
and U4977 (N_4977,N_3143,N_3277);
or U4978 (N_4978,N_3702,N_3391);
nand U4979 (N_4979,N_3800,N_3954);
xor U4980 (N_4980,N_3304,N_3387);
xor U4981 (N_4981,N_3448,N_3260);
nand U4982 (N_4982,N_3112,N_3818);
and U4983 (N_4983,N_3021,N_3694);
or U4984 (N_4984,N_3667,N_3580);
nor U4985 (N_4985,N_3814,N_3450);
nor U4986 (N_4986,N_3260,N_3253);
nor U4987 (N_4987,N_3584,N_3138);
nor U4988 (N_4988,N_3476,N_3559);
xor U4989 (N_4989,N_3180,N_3032);
nor U4990 (N_4990,N_3660,N_3012);
xnor U4991 (N_4991,N_3695,N_3405);
and U4992 (N_4992,N_3071,N_3337);
and U4993 (N_4993,N_3089,N_3521);
nor U4994 (N_4994,N_3419,N_3650);
or U4995 (N_4995,N_3858,N_3827);
xor U4996 (N_4996,N_3891,N_3742);
or U4997 (N_4997,N_3810,N_3031);
xnor U4998 (N_4998,N_3279,N_3805);
xor U4999 (N_4999,N_3557,N_3206);
or U5000 (N_5000,N_4809,N_4644);
and U5001 (N_5001,N_4839,N_4291);
or U5002 (N_5002,N_4777,N_4606);
nor U5003 (N_5003,N_4878,N_4334);
and U5004 (N_5004,N_4072,N_4690);
and U5005 (N_5005,N_4896,N_4026);
and U5006 (N_5006,N_4941,N_4985);
xor U5007 (N_5007,N_4421,N_4721);
xnor U5008 (N_5008,N_4104,N_4278);
xor U5009 (N_5009,N_4715,N_4868);
xor U5010 (N_5010,N_4163,N_4780);
nor U5011 (N_5011,N_4028,N_4645);
nor U5012 (N_5012,N_4182,N_4654);
xor U5013 (N_5013,N_4348,N_4097);
xor U5014 (N_5014,N_4245,N_4456);
xnor U5015 (N_5015,N_4442,N_4788);
or U5016 (N_5016,N_4725,N_4712);
xnor U5017 (N_5017,N_4710,N_4661);
nor U5018 (N_5018,N_4870,N_4750);
nor U5019 (N_5019,N_4186,N_4521);
xor U5020 (N_5020,N_4300,N_4465);
or U5021 (N_5021,N_4063,N_4293);
or U5022 (N_5022,N_4894,N_4524);
and U5023 (N_5023,N_4541,N_4543);
or U5024 (N_5024,N_4167,N_4717);
nand U5025 (N_5025,N_4169,N_4608);
nor U5026 (N_5026,N_4085,N_4216);
or U5027 (N_5027,N_4116,N_4526);
and U5028 (N_5028,N_4437,N_4301);
nand U5029 (N_5029,N_4774,N_4693);
nand U5030 (N_5030,N_4108,N_4002);
nor U5031 (N_5031,N_4588,N_4631);
nor U5032 (N_5032,N_4555,N_4770);
nand U5033 (N_5033,N_4461,N_4473);
nor U5034 (N_5034,N_4538,N_4280);
nand U5035 (N_5035,N_4975,N_4227);
nor U5036 (N_5036,N_4741,N_4203);
nor U5037 (N_5037,N_4785,N_4700);
or U5038 (N_5038,N_4350,N_4923);
and U5039 (N_5039,N_4578,N_4614);
and U5040 (N_5040,N_4393,N_4472);
nor U5041 (N_5041,N_4957,N_4748);
xor U5042 (N_5042,N_4586,N_4241);
nor U5043 (N_5043,N_4080,N_4045);
nor U5044 (N_5044,N_4575,N_4905);
and U5045 (N_5045,N_4112,N_4920);
nor U5046 (N_5046,N_4556,N_4434);
and U5047 (N_5047,N_4239,N_4722);
or U5048 (N_5048,N_4830,N_4598);
nor U5049 (N_5049,N_4643,N_4775);
nand U5050 (N_5050,N_4795,N_4796);
and U5051 (N_5051,N_4056,N_4219);
or U5052 (N_5052,N_4423,N_4288);
xnor U5053 (N_5053,N_4967,N_4211);
xor U5054 (N_5054,N_4847,N_4044);
nor U5055 (N_5055,N_4490,N_4345);
xnor U5056 (N_5056,N_4639,N_4043);
xnor U5057 (N_5057,N_4455,N_4095);
and U5058 (N_5058,N_4409,N_4294);
and U5059 (N_5059,N_4477,N_4435);
nand U5060 (N_5060,N_4867,N_4931);
or U5061 (N_5061,N_4733,N_4582);
nand U5062 (N_5062,N_4745,N_4600);
and U5063 (N_5063,N_4726,N_4162);
xnor U5064 (N_5064,N_4235,N_4206);
and U5065 (N_5065,N_4752,N_4798);
xnor U5066 (N_5066,N_4264,N_4910);
nand U5067 (N_5067,N_4836,N_4694);
and U5068 (N_5068,N_4376,N_4248);
nand U5069 (N_5069,N_4518,N_4340);
and U5070 (N_5070,N_4765,N_4478);
and U5071 (N_5071,N_4170,N_4512);
and U5072 (N_5072,N_4533,N_4572);
nor U5073 (N_5073,N_4189,N_4779);
and U5074 (N_5074,N_4630,N_4445);
nor U5075 (N_5075,N_4035,N_4713);
nand U5076 (N_5076,N_4401,N_4823);
or U5077 (N_5077,N_4115,N_4122);
xnor U5078 (N_5078,N_4411,N_4751);
nor U5079 (N_5079,N_4876,N_4328);
or U5080 (N_5080,N_4290,N_4962);
and U5081 (N_5081,N_4811,N_4386);
nand U5082 (N_5082,N_4025,N_4226);
xnor U5083 (N_5083,N_4793,N_4707);
and U5084 (N_5084,N_4164,N_4091);
or U5085 (N_5085,N_4205,N_4991);
nor U5086 (N_5086,N_4209,N_4902);
nor U5087 (N_5087,N_4316,N_4674);
and U5088 (N_5088,N_4269,N_4535);
or U5089 (N_5089,N_4503,N_4622);
nor U5090 (N_5090,N_4486,N_4958);
or U5091 (N_5091,N_4439,N_4354);
xnor U5092 (N_5092,N_4580,N_4621);
or U5093 (N_5093,N_4816,N_4760);
and U5094 (N_5094,N_4739,N_4545);
or U5095 (N_5095,N_4319,N_4221);
or U5096 (N_5096,N_4947,N_4948);
nor U5097 (N_5097,N_4031,N_4994);
and U5098 (N_5098,N_4367,N_4305);
and U5099 (N_5099,N_4375,N_4046);
and U5100 (N_5100,N_4799,N_4038);
nand U5101 (N_5101,N_4196,N_4756);
nand U5102 (N_5102,N_4051,N_4786);
xnor U5103 (N_5103,N_4980,N_4907);
or U5104 (N_5104,N_4866,N_4388);
xor U5105 (N_5105,N_4037,N_4475);
and U5106 (N_5106,N_4998,N_4520);
xnor U5107 (N_5107,N_4415,N_4502);
xor U5108 (N_5108,N_4881,N_4926);
nand U5109 (N_5109,N_4193,N_4360);
nand U5110 (N_5110,N_4605,N_4766);
nor U5111 (N_5111,N_4142,N_4986);
xor U5112 (N_5112,N_4691,N_4813);
or U5113 (N_5113,N_4394,N_4659);
and U5114 (N_5114,N_4029,N_4257);
nor U5115 (N_5115,N_4508,N_4871);
nand U5116 (N_5116,N_4671,N_4332);
nor U5117 (N_5117,N_4238,N_4889);
nor U5118 (N_5118,N_4047,N_4900);
and U5119 (N_5119,N_4454,N_4826);
nand U5120 (N_5120,N_4018,N_4109);
and U5121 (N_5121,N_4794,N_4297);
nand U5122 (N_5122,N_4769,N_4507);
or U5123 (N_5123,N_4424,N_4527);
and U5124 (N_5124,N_4407,N_4124);
nor U5125 (N_5125,N_4879,N_4113);
nor U5126 (N_5126,N_4107,N_4254);
nand U5127 (N_5127,N_4075,N_4010);
nand U5128 (N_5128,N_4458,N_4172);
nor U5129 (N_5129,N_4467,N_4174);
nor U5130 (N_5130,N_4596,N_4778);
or U5131 (N_5131,N_4074,N_4433);
and U5132 (N_5132,N_4247,N_4460);
nor U5133 (N_5133,N_4850,N_4464);
nor U5134 (N_5134,N_4098,N_4466);
or U5135 (N_5135,N_4997,N_4077);
nor U5136 (N_5136,N_4819,N_4152);
or U5137 (N_5137,N_4151,N_4263);
and U5138 (N_5138,N_4853,N_4976);
nor U5139 (N_5139,N_4706,N_4567);
xnor U5140 (N_5140,N_4494,N_4563);
xor U5141 (N_5141,N_4984,N_4338);
xor U5142 (N_5142,N_4824,N_4032);
and U5143 (N_5143,N_4383,N_4679);
or U5144 (N_5144,N_4062,N_4728);
nor U5145 (N_5145,N_4242,N_4703);
or U5146 (N_5146,N_4525,N_4365);
xor U5147 (N_5147,N_4451,N_4546);
and U5148 (N_5148,N_4228,N_4176);
nand U5149 (N_5149,N_4073,N_4325);
xnor U5150 (N_5150,N_4759,N_4523);
nor U5151 (N_5151,N_4347,N_4470);
and U5152 (N_5152,N_4559,N_4049);
nand U5153 (N_5153,N_4965,N_4898);
xor U5154 (N_5154,N_4719,N_4761);
nand U5155 (N_5155,N_4724,N_4873);
and U5156 (N_5156,N_4492,N_4207);
and U5157 (N_5157,N_4505,N_4530);
nor U5158 (N_5158,N_4515,N_4619);
or U5159 (N_5159,N_4822,N_4651);
and U5160 (N_5160,N_4253,N_4140);
and U5161 (N_5161,N_4202,N_4052);
nand U5162 (N_5162,N_4872,N_4323);
and U5163 (N_5163,N_4657,N_4021);
xnor U5164 (N_5164,N_4611,N_4625);
nor U5165 (N_5165,N_4704,N_4312);
and U5166 (N_5166,N_4033,N_4637);
nand U5167 (N_5167,N_4810,N_4531);
nand U5168 (N_5168,N_4379,N_4749);
nor U5169 (N_5169,N_4601,N_4971);
nor U5170 (N_5170,N_4865,N_4904);
nor U5171 (N_5171,N_4071,N_4925);
and U5172 (N_5172,N_4837,N_4584);
or U5173 (N_5173,N_4743,N_4491);
or U5174 (N_5174,N_4015,N_4855);
nand U5175 (N_5175,N_4141,N_4757);
nand U5176 (N_5176,N_4634,N_4061);
and U5177 (N_5177,N_4680,N_4883);
or U5178 (N_5178,N_4429,N_4337);
xor U5179 (N_5179,N_4101,N_4772);
and U5180 (N_5180,N_4534,N_4100);
nand U5181 (N_5181,N_4418,N_4689);
nand U5182 (N_5182,N_4720,N_4553);
nor U5183 (N_5183,N_4921,N_4309);
nor U5184 (N_5184,N_4979,N_4315);
or U5185 (N_5185,N_4673,N_4358);
xnor U5186 (N_5186,N_4457,N_4258);
nand U5187 (N_5187,N_4763,N_4060);
nor U5188 (N_5188,N_4686,N_4181);
xor U5189 (N_5189,N_4942,N_4413);
nor U5190 (N_5190,N_4016,N_4368);
nand U5191 (N_5191,N_4616,N_4642);
or U5192 (N_5192,N_4938,N_4117);
xor U5193 (N_5193,N_4560,N_4851);
xor U5194 (N_5194,N_4090,N_4735);
or U5195 (N_5195,N_4082,N_4310);
and U5196 (N_5196,N_4131,N_4989);
nor U5197 (N_5197,N_4862,N_4057);
nor U5198 (N_5198,N_4916,N_4506);
and U5199 (N_5199,N_4173,N_4628);
or U5200 (N_5200,N_4381,N_4869);
nor U5201 (N_5201,N_4908,N_4573);
and U5202 (N_5202,N_4183,N_4444);
xor U5203 (N_5203,N_4753,N_4498);
nand U5204 (N_5204,N_4385,N_4399);
and U5205 (N_5205,N_4988,N_4660);
xnor U5206 (N_5206,N_4877,N_4968);
or U5207 (N_5207,N_4274,N_4705);
nand U5208 (N_5208,N_4955,N_4331);
xor U5209 (N_5209,N_4570,N_4561);
or U5210 (N_5210,N_4913,N_4326);
nor U5211 (N_5211,N_4146,N_4727);
nor U5212 (N_5212,N_4237,N_4814);
nor U5213 (N_5213,N_4945,N_4564);
or U5214 (N_5214,N_4519,N_4893);
nand U5215 (N_5215,N_4463,N_4943);
or U5216 (N_5216,N_4180,N_4964);
and U5217 (N_5217,N_4177,N_4592);
nor U5218 (N_5218,N_4476,N_4542);
nor U5219 (N_5219,N_4079,N_4656);
nand U5220 (N_5220,N_4929,N_4144);
xor U5221 (N_5221,N_4504,N_4539);
or U5222 (N_5222,N_4511,N_4844);
nor U5223 (N_5223,N_4577,N_4776);
xnor U5224 (N_5224,N_4487,N_4011);
nor U5225 (N_5225,N_4800,N_4134);
xnor U5226 (N_5226,N_4436,N_4603);
xor U5227 (N_5227,N_4554,N_4155);
nor U5228 (N_5228,N_4184,N_4192);
nor U5229 (N_5229,N_4136,N_4672);
xor U5230 (N_5230,N_4357,N_4602);
and U5231 (N_5231,N_4001,N_4270);
or U5232 (N_5232,N_4302,N_4019);
nand U5233 (N_5233,N_4922,N_4903);
or U5234 (N_5234,N_4391,N_4396);
xnor U5235 (N_5235,N_4389,N_4303);
and U5236 (N_5236,N_4420,N_4479);
nand U5237 (N_5237,N_4150,N_4552);
nand U5238 (N_5238,N_4742,N_4311);
nand U5239 (N_5239,N_4935,N_4818);
nor U5240 (N_5240,N_4852,N_4158);
and U5241 (N_5241,N_4138,N_4084);
and U5242 (N_5242,N_4730,N_4392);
nand U5243 (N_5243,N_4683,N_4204);
or U5244 (N_5244,N_4857,N_4304);
nor U5245 (N_5245,N_4408,N_4884);
and U5246 (N_5246,N_4569,N_4398);
or U5247 (N_5247,N_4343,N_4432);
xnor U5248 (N_5248,N_4681,N_4911);
xnor U5249 (N_5249,N_4990,N_4327);
xnor U5250 (N_5250,N_4017,N_4547);
xor U5251 (N_5251,N_4145,N_4863);
nand U5252 (N_5252,N_4428,N_4118);
xor U5253 (N_5253,N_4450,N_4734);
nor U5254 (N_5254,N_4023,N_4736);
nor U5255 (N_5255,N_4027,N_4917);
or U5256 (N_5256,N_4246,N_4230);
and U5257 (N_5257,N_4522,N_4664);
xor U5258 (N_5258,N_4285,N_4251);
xnor U5259 (N_5259,N_4738,N_4212);
xnor U5260 (N_5260,N_4933,N_4528);
and U5261 (N_5261,N_4185,N_4532);
nor U5262 (N_5262,N_4792,N_4675);
nand U5263 (N_5263,N_4156,N_4537);
xnor U5264 (N_5264,N_4655,N_4557);
xnor U5265 (N_5265,N_4781,N_4784);
and U5266 (N_5266,N_4906,N_4314);
or U5267 (N_5267,N_4448,N_4787);
nand U5268 (N_5268,N_4609,N_4972);
xnor U5269 (N_5269,N_4571,N_4154);
and U5270 (N_5270,N_4832,N_4973);
xnor U5271 (N_5271,N_4668,N_4279);
and U5272 (N_5272,N_4509,N_4897);
nand U5273 (N_5273,N_4481,N_4566);
and U5274 (N_5274,N_4482,N_4669);
or U5275 (N_5275,N_4854,N_4562);
nand U5276 (N_5276,N_4344,N_4802);
nand U5277 (N_5277,N_4373,N_4648);
nor U5278 (N_5278,N_4208,N_4848);
nor U5279 (N_5279,N_4210,N_4036);
xor U5280 (N_5280,N_4013,N_4159);
or U5281 (N_5281,N_4791,N_4133);
or U5282 (N_5282,N_4803,N_4059);
and U5283 (N_5283,N_4058,N_4342);
or U5284 (N_5284,N_4692,N_4320);
and U5285 (N_5285,N_4252,N_4899);
and U5286 (N_5286,N_4308,N_4548);
or U5287 (N_5287,N_4970,N_4633);
nor U5288 (N_5288,N_4307,N_4882);
and U5289 (N_5289,N_4918,N_4747);
and U5290 (N_5290,N_4333,N_4652);
xor U5291 (N_5291,N_4371,N_4583);
nand U5292 (N_5292,N_4716,N_4828);
xnor U5293 (N_5293,N_4233,N_4352);
and U5294 (N_5294,N_4377,N_4773);
and U5295 (N_5295,N_4914,N_4081);
nor U5296 (N_5296,N_4623,N_4499);
nor U5297 (N_5297,N_4066,N_4587);
or U5298 (N_5298,N_4963,N_4374);
and U5299 (N_5299,N_4983,N_4153);
and U5300 (N_5300,N_4372,N_4771);
nand U5301 (N_5301,N_4624,N_4888);
nor U5302 (N_5302,N_4629,N_4111);
nor U5303 (N_5303,N_4483,N_4610);
nor U5304 (N_5304,N_4646,N_4093);
xor U5305 (N_5305,N_4329,N_4874);
nor U5306 (N_5306,N_4215,N_4821);
or U5307 (N_5307,N_4272,N_4083);
nor U5308 (N_5308,N_4198,N_4232);
xor U5309 (N_5309,N_4070,N_4147);
and U5310 (N_5310,N_4662,N_4324);
xor U5311 (N_5311,N_4143,N_4737);
or U5312 (N_5312,N_4382,N_4488);
or U5313 (N_5313,N_4149,N_4223);
or U5314 (N_5314,N_4982,N_4236);
nand U5315 (N_5315,N_4480,N_4006);
or U5316 (N_5316,N_4403,N_4485);
nor U5317 (N_5317,N_4412,N_4353);
and U5318 (N_5318,N_4168,N_4089);
or U5319 (N_5319,N_4321,N_4709);
and U5320 (N_5320,N_4020,N_4714);
xor U5321 (N_5321,N_4283,N_4449);
nand U5322 (N_5322,N_4260,N_4369);
nand U5323 (N_5323,N_4128,N_4201);
and U5324 (N_5324,N_4322,N_4797);
nand U5325 (N_5325,N_4387,N_4231);
or U5326 (N_5326,N_4318,N_4262);
xor U5327 (N_5327,N_4953,N_4723);
and U5328 (N_5328,N_4670,N_4240);
or U5329 (N_5329,N_4936,N_4946);
nor U5330 (N_5330,N_4419,N_4175);
nor U5331 (N_5331,N_4806,N_4361);
xnor U5332 (N_5332,N_4627,N_4699);
xnor U5333 (N_5333,N_4362,N_4256);
and U5334 (N_5334,N_4468,N_4767);
or U5335 (N_5335,N_4484,N_4042);
or U5336 (N_5336,N_4313,N_4834);
xor U5337 (N_5337,N_4607,N_4617);
and U5338 (N_5338,N_4453,N_4000);
and U5339 (N_5339,N_4992,N_4827);
or U5340 (N_5340,N_4397,N_4551);
xnor U5341 (N_5341,N_4249,N_4860);
or U5342 (N_5342,N_4641,N_4978);
nand U5343 (N_5343,N_4114,N_4076);
nor U5344 (N_5344,N_4593,N_4363);
and U5345 (N_5345,N_4840,N_4430);
nor U5346 (N_5346,N_4086,N_4842);
and U5347 (N_5347,N_4349,N_4462);
xor U5348 (N_5348,N_4431,N_4514);
or U5349 (N_5349,N_4030,N_4157);
xnor U5350 (N_5350,N_4843,N_4536);
nor U5351 (N_5351,N_4999,N_4078);
xnor U5352 (N_5352,N_4296,N_4804);
xnor U5353 (N_5353,N_4649,N_4041);
nor U5354 (N_5354,N_4171,N_4579);
nor U5355 (N_5355,N_4224,N_4495);
nor U5356 (N_5356,N_4267,N_4817);
xor U5357 (N_5357,N_4783,N_4426);
xnor U5358 (N_5358,N_4459,N_4335);
and U5359 (N_5359,N_4474,N_4489);
xor U5360 (N_5360,N_4590,N_4048);
nor U5361 (N_5361,N_4271,N_4934);
nor U5362 (N_5362,N_4831,N_4259);
xnor U5363 (N_5363,N_4808,N_4885);
xor U5364 (N_5364,N_4053,N_4613);
and U5365 (N_5365,N_4125,N_4195);
xnor U5366 (N_5366,N_4008,N_4165);
xor U5367 (N_5367,N_4764,N_4568);
nor U5368 (N_5368,N_4287,N_4234);
nand U5369 (N_5369,N_4054,N_4864);
nand U5370 (N_5370,N_4126,N_4944);
nand U5371 (N_5371,N_4050,N_4135);
nand U5372 (N_5372,N_4517,N_4178);
nor U5373 (N_5373,N_4589,N_4820);
nand U5374 (N_5374,N_4166,N_4443);
nor U5375 (N_5375,N_4404,N_4665);
and U5376 (N_5376,N_4218,N_4410);
nor U5377 (N_5377,N_4981,N_4427);
xor U5378 (N_5378,N_4996,N_4447);
xnor U5379 (N_5379,N_4446,N_4441);
nor U5380 (N_5380,N_4677,N_4012);
nand U5381 (N_5381,N_4891,N_4951);
nor U5382 (N_5382,N_4754,N_4604);
and U5383 (N_5383,N_4132,N_4406);
xor U5384 (N_5384,N_4284,N_4317);
or U5385 (N_5385,N_4250,N_4103);
or U5386 (N_5386,N_4214,N_4243);
xnor U5387 (N_5387,N_4650,N_4364);
nand U5388 (N_5388,N_4217,N_4179);
nand U5389 (N_5389,N_4678,N_4640);
or U5390 (N_5390,N_4977,N_4121);
xor U5391 (N_5391,N_4960,N_4886);
or U5392 (N_5392,N_4336,N_4758);
or U5393 (N_5393,N_4356,N_4956);
or U5394 (N_5394,N_4928,N_4647);
nand U5395 (N_5395,N_4299,N_4127);
and U5396 (N_5396,N_4915,N_4684);
xnor U5397 (N_5397,N_4695,N_4003);
nand U5398 (N_5398,N_4636,N_4746);
xnor U5399 (N_5399,N_4007,N_4940);
nor U5400 (N_5400,N_4096,N_4768);
xnor U5401 (N_5401,N_4969,N_4615);
xor U5402 (N_5402,N_4510,N_4974);
or U5403 (N_5403,N_4416,N_4846);
or U5404 (N_5404,N_4068,N_4581);
or U5405 (N_5405,N_4229,N_4618);
nor U5406 (N_5406,N_4856,N_4711);
xor U5407 (N_5407,N_4950,N_4222);
nor U5408 (N_5408,N_4841,N_4346);
and U5409 (N_5409,N_4493,N_4663);
xor U5410 (N_5410,N_4801,N_4281);
nand U5411 (N_5411,N_4927,N_4295);
nor U5412 (N_5412,N_4330,N_4064);
nand U5413 (N_5413,N_4440,N_4400);
xnor U5414 (N_5414,N_4009,N_4701);
nor U5415 (N_5415,N_4932,N_4959);
or U5416 (N_5416,N_4040,N_4731);
or U5417 (N_5417,N_4402,N_4626);
nor U5418 (N_5418,N_4191,N_4014);
xor U5419 (N_5419,N_4835,N_4366);
or U5420 (N_5420,N_4405,N_4762);
nor U5421 (N_5421,N_4190,N_4500);
nand U5422 (N_5422,N_4858,N_4924);
or U5423 (N_5423,N_4638,N_4937);
nand U5424 (N_5424,N_4698,N_4123);
nor U5425 (N_5425,N_4597,N_4298);
nand U5426 (N_5426,N_4261,N_4496);
or U5427 (N_5427,N_4110,N_4708);
xor U5428 (N_5428,N_4092,N_4292);
or U5429 (N_5429,N_4595,N_4501);
or U5430 (N_5430,N_4952,N_4740);
or U5431 (N_5431,N_4685,N_4676);
xnor U5432 (N_5432,N_4805,N_4591);
xnor U5433 (N_5433,N_4004,N_4667);
and U5434 (N_5434,N_4789,N_4875);
or U5435 (N_5435,N_4188,N_4351);
xnor U5436 (N_5436,N_4688,N_4544);
or U5437 (N_5437,N_4620,N_4892);
or U5438 (N_5438,N_4729,N_4102);
nor U5439 (N_5439,N_4024,N_4119);
or U5440 (N_5440,N_4067,N_4306);
and U5441 (N_5441,N_4666,N_4549);
xor U5442 (N_5442,N_4160,N_4909);
and U5443 (N_5443,N_4282,N_4120);
or U5444 (N_5444,N_4452,N_4161);
and U5445 (N_5445,N_4732,N_4148);
nor U5446 (N_5446,N_4930,N_4378);
xor U5447 (N_5447,N_4471,N_4187);
xnor U5448 (N_5448,N_4696,N_4022);
or U5449 (N_5449,N_4594,N_4390);
or U5450 (N_5450,N_4612,N_4635);
nand U5451 (N_5451,N_4632,N_4995);
and U5452 (N_5452,N_4782,N_4276);
xor U5453 (N_5453,N_4954,N_4919);
nand U5454 (N_5454,N_4755,N_4812);
xnor U5455 (N_5455,N_4065,N_4417);
nor U5456 (N_5456,N_4558,N_4697);
xnor U5457 (N_5457,N_4422,N_4744);
or U5458 (N_5458,N_4702,N_4244);
xor U5459 (N_5459,N_4895,N_4137);
or U5460 (N_5460,N_4380,N_4289);
nor U5461 (N_5461,N_4194,N_4576);
nor U5462 (N_5462,N_4890,N_4961);
or U5463 (N_5463,N_4497,N_4277);
nand U5464 (N_5464,N_4268,N_4833);
or U5465 (N_5465,N_4069,N_4825);
and U5466 (N_5466,N_4469,N_4106);
nor U5467 (N_5467,N_4341,N_4845);
nand U5468 (N_5468,N_4425,N_4585);
and U5469 (N_5469,N_4105,N_4087);
and U5470 (N_5470,N_4273,N_4265);
and U5471 (N_5471,N_4200,N_4034);
xnor U5472 (N_5472,N_4414,N_4966);
and U5473 (N_5473,N_4339,N_4199);
nand U5474 (N_5474,N_4225,N_4094);
and U5475 (N_5475,N_4987,N_4359);
or U5476 (N_5476,N_4807,N_4682);
and U5477 (N_5477,N_4255,N_4540);
nor U5478 (N_5478,N_4718,N_4880);
and U5479 (N_5479,N_4550,N_4912);
xnor U5480 (N_5480,N_4213,N_4574);
and U5481 (N_5481,N_4838,N_4130);
or U5482 (N_5482,N_4829,N_4653);
or U5483 (N_5483,N_4529,N_4599);
xor U5484 (N_5484,N_4993,N_4949);
nor U5485 (N_5485,N_4939,N_4790);
nor U5486 (N_5486,N_4005,N_4139);
nor U5487 (N_5487,N_4039,N_4055);
nand U5488 (N_5488,N_4861,N_4887);
or U5489 (N_5489,N_4687,N_4901);
xor U5490 (N_5490,N_4516,N_4438);
and U5491 (N_5491,N_4197,N_4513);
nand U5492 (N_5492,N_4266,N_4815);
or U5493 (N_5493,N_4088,N_4658);
xnor U5494 (N_5494,N_4565,N_4355);
and U5495 (N_5495,N_4220,N_4275);
or U5496 (N_5496,N_4129,N_4849);
xnor U5497 (N_5497,N_4370,N_4384);
nor U5498 (N_5498,N_4286,N_4099);
nand U5499 (N_5499,N_4859,N_4395);
nand U5500 (N_5500,N_4886,N_4640);
and U5501 (N_5501,N_4348,N_4161);
xnor U5502 (N_5502,N_4391,N_4806);
nor U5503 (N_5503,N_4373,N_4076);
and U5504 (N_5504,N_4994,N_4963);
and U5505 (N_5505,N_4510,N_4579);
xor U5506 (N_5506,N_4033,N_4904);
or U5507 (N_5507,N_4683,N_4780);
or U5508 (N_5508,N_4852,N_4730);
xor U5509 (N_5509,N_4961,N_4038);
and U5510 (N_5510,N_4961,N_4572);
nor U5511 (N_5511,N_4376,N_4901);
or U5512 (N_5512,N_4549,N_4495);
nor U5513 (N_5513,N_4803,N_4051);
xnor U5514 (N_5514,N_4017,N_4699);
nor U5515 (N_5515,N_4506,N_4231);
xnor U5516 (N_5516,N_4601,N_4998);
or U5517 (N_5517,N_4618,N_4293);
nor U5518 (N_5518,N_4058,N_4117);
nor U5519 (N_5519,N_4538,N_4777);
nand U5520 (N_5520,N_4824,N_4718);
xor U5521 (N_5521,N_4753,N_4219);
nor U5522 (N_5522,N_4641,N_4799);
xor U5523 (N_5523,N_4656,N_4318);
xor U5524 (N_5524,N_4086,N_4146);
xnor U5525 (N_5525,N_4596,N_4932);
and U5526 (N_5526,N_4004,N_4131);
xor U5527 (N_5527,N_4100,N_4459);
nand U5528 (N_5528,N_4889,N_4666);
and U5529 (N_5529,N_4639,N_4909);
nor U5530 (N_5530,N_4007,N_4734);
and U5531 (N_5531,N_4566,N_4537);
and U5532 (N_5532,N_4262,N_4109);
xor U5533 (N_5533,N_4270,N_4327);
xor U5534 (N_5534,N_4070,N_4478);
and U5535 (N_5535,N_4343,N_4147);
nand U5536 (N_5536,N_4728,N_4583);
nor U5537 (N_5537,N_4429,N_4417);
xor U5538 (N_5538,N_4119,N_4432);
nor U5539 (N_5539,N_4150,N_4982);
xnor U5540 (N_5540,N_4644,N_4616);
and U5541 (N_5541,N_4265,N_4347);
nor U5542 (N_5542,N_4498,N_4316);
or U5543 (N_5543,N_4141,N_4792);
xnor U5544 (N_5544,N_4139,N_4254);
xnor U5545 (N_5545,N_4104,N_4836);
xnor U5546 (N_5546,N_4213,N_4381);
and U5547 (N_5547,N_4221,N_4828);
nand U5548 (N_5548,N_4490,N_4777);
xor U5549 (N_5549,N_4569,N_4295);
nor U5550 (N_5550,N_4037,N_4006);
and U5551 (N_5551,N_4846,N_4011);
and U5552 (N_5552,N_4989,N_4615);
or U5553 (N_5553,N_4853,N_4226);
or U5554 (N_5554,N_4608,N_4643);
nand U5555 (N_5555,N_4830,N_4038);
xor U5556 (N_5556,N_4397,N_4401);
xnor U5557 (N_5557,N_4642,N_4299);
and U5558 (N_5558,N_4781,N_4752);
xor U5559 (N_5559,N_4939,N_4706);
nand U5560 (N_5560,N_4560,N_4799);
nor U5561 (N_5561,N_4921,N_4245);
nor U5562 (N_5562,N_4693,N_4759);
nand U5563 (N_5563,N_4049,N_4631);
nor U5564 (N_5564,N_4282,N_4369);
nor U5565 (N_5565,N_4385,N_4348);
or U5566 (N_5566,N_4051,N_4264);
xor U5567 (N_5567,N_4401,N_4881);
nor U5568 (N_5568,N_4674,N_4868);
nor U5569 (N_5569,N_4438,N_4418);
xor U5570 (N_5570,N_4867,N_4972);
and U5571 (N_5571,N_4674,N_4203);
nand U5572 (N_5572,N_4452,N_4889);
nor U5573 (N_5573,N_4840,N_4292);
or U5574 (N_5574,N_4813,N_4427);
or U5575 (N_5575,N_4723,N_4299);
xor U5576 (N_5576,N_4105,N_4707);
and U5577 (N_5577,N_4638,N_4571);
xor U5578 (N_5578,N_4510,N_4518);
nand U5579 (N_5579,N_4962,N_4429);
nand U5580 (N_5580,N_4022,N_4093);
or U5581 (N_5581,N_4039,N_4550);
nor U5582 (N_5582,N_4767,N_4521);
or U5583 (N_5583,N_4937,N_4210);
or U5584 (N_5584,N_4081,N_4812);
nor U5585 (N_5585,N_4271,N_4755);
nand U5586 (N_5586,N_4014,N_4290);
or U5587 (N_5587,N_4739,N_4664);
and U5588 (N_5588,N_4537,N_4380);
nand U5589 (N_5589,N_4167,N_4249);
or U5590 (N_5590,N_4294,N_4615);
nand U5591 (N_5591,N_4234,N_4986);
or U5592 (N_5592,N_4894,N_4239);
nand U5593 (N_5593,N_4925,N_4650);
or U5594 (N_5594,N_4754,N_4757);
or U5595 (N_5595,N_4178,N_4497);
and U5596 (N_5596,N_4076,N_4484);
or U5597 (N_5597,N_4198,N_4828);
or U5598 (N_5598,N_4008,N_4537);
nor U5599 (N_5599,N_4500,N_4977);
nand U5600 (N_5600,N_4235,N_4944);
nand U5601 (N_5601,N_4752,N_4817);
and U5602 (N_5602,N_4766,N_4341);
and U5603 (N_5603,N_4489,N_4007);
nor U5604 (N_5604,N_4819,N_4567);
nand U5605 (N_5605,N_4792,N_4721);
nor U5606 (N_5606,N_4429,N_4257);
nor U5607 (N_5607,N_4472,N_4940);
nand U5608 (N_5608,N_4295,N_4913);
xnor U5609 (N_5609,N_4715,N_4351);
or U5610 (N_5610,N_4316,N_4262);
nor U5611 (N_5611,N_4212,N_4865);
and U5612 (N_5612,N_4479,N_4379);
xnor U5613 (N_5613,N_4300,N_4403);
nand U5614 (N_5614,N_4560,N_4919);
nor U5615 (N_5615,N_4174,N_4722);
or U5616 (N_5616,N_4123,N_4037);
or U5617 (N_5617,N_4344,N_4991);
or U5618 (N_5618,N_4839,N_4965);
and U5619 (N_5619,N_4627,N_4402);
xor U5620 (N_5620,N_4802,N_4353);
xor U5621 (N_5621,N_4247,N_4025);
nand U5622 (N_5622,N_4219,N_4516);
and U5623 (N_5623,N_4302,N_4625);
xnor U5624 (N_5624,N_4851,N_4712);
and U5625 (N_5625,N_4701,N_4886);
nor U5626 (N_5626,N_4086,N_4227);
and U5627 (N_5627,N_4338,N_4620);
xor U5628 (N_5628,N_4739,N_4239);
nor U5629 (N_5629,N_4283,N_4302);
nor U5630 (N_5630,N_4602,N_4839);
or U5631 (N_5631,N_4873,N_4439);
and U5632 (N_5632,N_4702,N_4890);
xnor U5633 (N_5633,N_4406,N_4817);
or U5634 (N_5634,N_4287,N_4062);
and U5635 (N_5635,N_4702,N_4457);
or U5636 (N_5636,N_4645,N_4708);
nand U5637 (N_5637,N_4945,N_4418);
xor U5638 (N_5638,N_4965,N_4202);
nand U5639 (N_5639,N_4845,N_4730);
or U5640 (N_5640,N_4264,N_4296);
or U5641 (N_5641,N_4242,N_4072);
or U5642 (N_5642,N_4808,N_4564);
and U5643 (N_5643,N_4880,N_4500);
or U5644 (N_5644,N_4552,N_4689);
and U5645 (N_5645,N_4373,N_4424);
and U5646 (N_5646,N_4869,N_4534);
xnor U5647 (N_5647,N_4138,N_4163);
or U5648 (N_5648,N_4003,N_4121);
or U5649 (N_5649,N_4358,N_4336);
or U5650 (N_5650,N_4786,N_4490);
or U5651 (N_5651,N_4618,N_4766);
nor U5652 (N_5652,N_4204,N_4015);
nor U5653 (N_5653,N_4701,N_4463);
nor U5654 (N_5654,N_4671,N_4188);
and U5655 (N_5655,N_4111,N_4447);
xnor U5656 (N_5656,N_4658,N_4203);
nand U5657 (N_5657,N_4475,N_4225);
xor U5658 (N_5658,N_4676,N_4199);
nand U5659 (N_5659,N_4548,N_4259);
or U5660 (N_5660,N_4488,N_4199);
and U5661 (N_5661,N_4937,N_4753);
and U5662 (N_5662,N_4256,N_4668);
or U5663 (N_5663,N_4729,N_4436);
xor U5664 (N_5664,N_4975,N_4866);
xnor U5665 (N_5665,N_4502,N_4190);
nand U5666 (N_5666,N_4374,N_4552);
xnor U5667 (N_5667,N_4533,N_4683);
nand U5668 (N_5668,N_4574,N_4934);
nand U5669 (N_5669,N_4910,N_4281);
and U5670 (N_5670,N_4369,N_4771);
nand U5671 (N_5671,N_4802,N_4039);
and U5672 (N_5672,N_4871,N_4465);
nand U5673 (N_5673,N_4807,N_4391);
nor U5674 (N_5674,N_4878,N_4119);
and U5675 (N_5675,N_4385,N_4451);
or U5676 (N_5676,N_4860,N_4416);
nand U5677 (N_5677,N_4068,N_4182);
xor U5678 (N_5678,N_4873,N_4217);
or U5679 (N_5679,N_4491,N_4389);
nor U5680 (N_5680,N_4323,N_4210);
xor U5681 (N_5681,N_4115,N_4598);
and U5682 (N_5682,N_4538,N_4717);
nor U5683 (N_5683,N_4272,N_4657);
and U5684 (N_5684,N_4608,N_4488);
nor U5685 (N_5685,N_4292,N_4667);
or U5686 (N_5686,N_4564,N_4654);
or U5687 (N_5687,N_4196,N_4810);
xor U5688 (N_5688,N_4587,N_4668);
nand U5689 (N_5689,N_4523,N_4554);
xnor U5690 (N_5690,N_4131,N_4789);
nor U5691 (N_5691,N_4308,N_4816);
nand U5692 (N_5692,N_4632,N_4145);
and U5693 (N_5693,N_4438,N_4286);
xor U5694 (N_5694,N_4652,N_4298);
or U5695 (N_5695,N_4612,N_4068);
xor U5696 (N_5696,N_4282,N_4157);
xor U5697 (N_5697,N_4204,N_4091);
or U5698 (N_5698,N_4828,N_4123);
and U5699 (N_5699,N_4809,N_4077);
nor U5700 (N_5700,N_4564,N_4289);
or U5701 (N_5701,N_4853,N_4130);
nand U5702 (N_5702,N_4808,N_4669);
nor U5703 (N_5703,N_4635,N_4251);
and U5704 (N_5704,N_4725,N_4103);
nor U5705 (N_5705,N_4911,N_4850);
xor U5706 (N_5706,N_4597,N_4203);
nand U5707 (N_5707,N_4628,N_4709);
nor U5708 (N_5708,N_4496,N_4963);
or U5709 (N_5709,N_4812,N_4800);
or U5710 (N_5710,N_4317,N_4696);
nor U5711 (N_5711,N_4949,N_4452);
and U5712 (N_5712,N_4966,N_4611);
and U5713 (N_5713,N_4609,N_4964);
nor U5714 (N_5714,N_4064,N_4633);
or U5715 (N_5715,N_4031,N_4444);
nand U5716 (N_5716,N_4185,N_4103);
nand U5717 (N_5717,N_4370,N_4588);
and U5718 (N_5718,N_4983,N_4772);
xnor U5719 (N_5719,N_4537,N_4988);
nor U5720 (N_5720,N_4273,N_4551);
nor U5721 (N_5721,N_4227,N_4053);
nor U5722 (N_5722,N_4989,N_4106);
and U5723 (N_5723,N_4068,N_4646);
nand U5724 (N_5724,N_4975,N_4013);
xor U5725 (N_5725,N_4040,N_4038);
nand U5726 (N_5726,N_4007,N_4382);
nand U5727 (N_5727,N_4480,N_4978);
xor U5728 (N_5728,N_4492,N_4338);
nor U5729 (N_5729,N_4984,N_4852);
nor U5730 (N_5730,N_4442,N_4661);
and U5731 (N_5731,N_4048,N_4344);
xnor U5732 (N_5732,N_4823,N_4789);
xor U5733 (N_5733,N_4908,N_4913);
or U5734 (N_5734,N_4418,N_4150);
or U5735 (N_5735,N_4329,N_4385);
and U5736 (N_5736,N_4807,N_4771);
xor U5737 (N_5737,N_4684,N_4800);
or U5738 (N_5738,N_4316,N_4525);
and U5739 (N_5739,N_4632,N_4125);
or U5740 (N_5740,N_4703,N_4836);
xnor U5741 (N_5741,N_4432,N_4257);
nor U5742 (N_5742,N_4025,N_4849);
and U5743 (N_5743,N_4384,N_4696);
nor U5744 (N_5744,N_4886,N_4312);
and U5745 (N_5745,N_4721,N_4506);
and U5746 (N_5746,N_4196,N_4423);
and U5747 (N_5747,N_4270,N_4380);
or U5748 (N_5748,N_4555,N_4154);
nor U5749 (N_5749,N_4596,N_4413);
and U5750 (N_5750,N_4964,N_4188);
nand U5751 (N_5751,N_4752,N_4320);
or U5752 (N_5752,N_4709,N_4333);
nand U5753 (N_5753,N_4285,N_4145);
nor U5754 (N_5754,N_4990,N_4985);
nand U5755 (N_5755,N_4111,N_4722);
and U5756 (N_5756,N_4897,N_4439);
xnor U5757 (N_5757,N_4336,N_4839);
xnor U5758 (N_5758,N_4619,N_4395);
and U5759 (N_5759,N_4626,N_4207);
and U5760 (N_5760,N_4720,N_4638);
nor U5761 (N_5761,N_4326,N_4496);
or U5762 (N_5762,N_4230,N_4182);
or U5763 (N_5763,N_4376,N_4175);
nand U5764 (N_5764,N_4156,N_4795);
or U5765 (N_5765,N_4016,N_4343);
or U5766 (N_5766,N_4061,N_4705);
and U5767 (N_5767,N_4343,N_4369);
nor U5768 (N_5768,N_4274,N_4891);
nor U5769 (N_5769,N_4380,N_4886);
and U5770 (N_5770,N_4840,N_4057);
nor U5771 (N_5771,N_4077,N_4735);
xnor U5772 (N_5772,N_4314,N_4046);
nand U5773 (N_5773,N_4490,N_4833);
or U5774 (N_5774,N_4101,N_4024);
xor U5775 (N_5775,N_4086,N_4147);
nand U5776 (N_5776,N_4414,N_4359);
xor U5777 (N_5777,N_4961,N_4328);
nand U5778 (N_5778,N_4443,N_4198);
nand U5779 (N_5779,N_4782,N_4936);
or U5780 (N_5780,N_4816,N_4595);
nor U5781 (N_5781,N_4390,N_4499);
nor U5782 (N_5782,N_4047,N_4568);
xnor U5783 (N_5783,N_4360,N_4307);
and U5784 (N_5784,N_4306,N_4352);
xor U5785 (N_5785,N_4654,N_4829);
and U5786 (N_5786,N_4843,N_4559);
xor U5787 (N_5787,N_4309,N_4325);
xnor U5788 (N_5788,N_4931,N_4101);
xor U5789 (N_5789,N_4945,N_4457);
nand U5790 (N_5790,N_4539,N_4473);
nand U5791 (N_5791,N_4307,N_4520);
xnor U5792 (N_5792,N_4797,N_4920);
xnor U5793 (N_5793,N_4225,N_4502);
nand U5794 (N_5794,N_4676,N_4902);
nand U5795 (N_5795,N_4235,N_4665);
or U5796 (N_5796,N_4313,N_4271);
or U5797 (N_5797,N_4242,N_4950);
xnor U5798 (N_5798,N_4331,N_4086);
nor U5799 (N_5799,N_4685,N_4860);
and U5800 (N_5800,N_4130,N_4171);
nor U5801 (N_5801,N_4653,N_4695);
or U5802 (N_5802,N_4771,N_4909);
nand U5803 (N_5803,N_4359,N_4749);
nand U5804 (N_5804,N_4385,N_4804);
nor U5805 (N_5805,N_4960,N_4430);
nand U5806 (N_5806,N_4571,N_4897);
nand U5807 (N_5807,N_4319,N_4686);
or U5808 (N_5808,N_4557,N_4724);
nor U5809 (N_5809,N_4549,N_4314);
nand U5810 (N_5810,N_4197,N_4294);
and U5811 (N_5811,N_4956,N_4071);
nor U5812 (N_5812,N_4550,N_4821);
or U5813 (N_5813,N_4226,N_4262);
or U5814 (N_5814,N_4344,N_4386);
or U5815 (N_5815,N_4681,N_4025);
and U5816 (N_5816,N_4982,N_4647);
nand U5817 (N_5817,N_4511,N_4289);
xor U5818 (N_5818,N_4833,N_4025);
nand U5819 (N_5819,N_4285,N_4629);
and U5820 (N_5820,N_4477,N_4595);
nand U5821 (N_5821,N_4769,N_4271);
and U5822 (N_5822,N_4159,N_4766);
xnor U5823 (N_5823,N_4590,N_4469);
or U5824 (N_5824,N_4471,N_4806);
xnor U5825 (N_5825,N_4834,N_4369);
nor U5826 (N_5826,N_4471,N_4165);
or U5827 (N_5827,N_4971,N_4637);
nand U5828 (N_5828,N_4034,N_4681);
and U5829 (N_5829,N_4133,N_4428);
or U5830 (N_5830,N_4222,N_4100);
xnor U5831 (N_5831,N_4269,N_4452);
nand U5832 (N_5832,N_4053,N_4095);
nor U5833 (N_5833,N_4476,N_4687);
nand U5834 (N_5834,N_4397,N_4297);
nor U5835 (N_5835,N_4690,N_4921);
and U5836 (N_5836,N_4184,N_4276);
nor U5837 (N_5837,N_4269,N_4469);
xor U5838 (N_5838,N_4109,N_4647);
nor U5839 (N_5839,N_4497,N_4672);
xnor U5840 (N_5840,N_4548,N_4640);
or U5841 (N_5841,N_4596,N_4509);
and U5842 (N_5842,N_4688,N_4873);
xnor U5843 (N_5843,N_4325,N_4408);
nand U5844 (N_5844,N_4683,N_4337);
xor U5845 (N_5845,N_4814,N_4907);
or U5846 (N_5846,N_4196,N_4643);
and U5847 (N_5847,N_4308,N_4280);
xor U5848 (N_5848,N_4448,N_4204);
nand U5849 (N_5849,N_4704,N_4003);
nor U5850 (N_5850,N_4969,N_4977);
nand U5851 (N_5851,N_4656,N_4125);
or U5852 (N_5852,N_4866,N_4206);
and U5853 (N_5853,N_4710,N_4712);
nor U5854 (N_5854,N_4035,N_4640);
nor U5855 (N_5855,N_4992,N_4206);
and U5856 (N_5856,N_4599,N_4183);
and U5857 (N_5857,N_4665,N_4947);
or U5858 (N_5858,N_4033,N_4592);
and U5859 (N_5859,N_4111,N_4199);
and U5860 (N_5860,N_4818,N_4426);
or U5861 (N_5861,N_4108,N_4847);
nand U5862 (N_5862,N_4789,N_4263);
nor U5863 (N_5863,N_4771,N_4192);
nor U5864 (N_5864,N_4463,N_4632);
and U5865 (N_5865,N_4394,N_4030);
xnor U5866 (N_5866,N_4160,N_4141);
nand U5867 (N_5867,N_4199,N_4685);
nand U5868 (N_5868,N_4255,N_4235);
nand U5869 (N_5869,N_4840,N_4120);
or U5870 (N_5870,N_4604,N_4117);
and U5871 (N_5871,N_4739,N_4751);
and U5872 (N_5872,N_4063,N_4845);
xnor U5873 (N_5873,N_4067,N_4521);
and U5874 (N_5874,N_4300,N_4804);
nor U5875 (N_5875,N_4244,N_4784);
nand U5876 (N_5876,N_4697,N_4165);
or U5877 (N_5877,N_4122,N_4665);
nand U5878 (N_5878,N_4319,N_4133);
and U5879 (N_5879,N_4252,N_4516);
nand U5880 (N_5880,N_4798,N_4364);
nand U5881 (N_5881,N_4849,N_4260);
xor U5882 (N_5882,N_4654,N_4986);
nor U5883 (N_5883,N_4033,N_4756);
nand U5884 (N_5884,N_4637,N_4242);
nand U5885 (N_5885,N_4545,N_4015);
nor U5886 (N_5886,N_4891,N_4846);
and U5887 (N_5887,N_4965,N_4482);
nor U5888 (N_5888,N_4806,N_4132);
or U5889 (N_5889,N_4712,N_4954);
nor U5890 (N_5890,N_4570,N_4926);
nand U5891 (N_5891,N_4242,N_4248);
xor U5892 (N_5892,N_4142,N_4651);
and U5893 (N_5893,N_4407,N_4267);
or U5894 (N_5894,N_4240,N_4001);
or U5895 (N_5895,N_4506,N_4620);
nand U5896 (N_5896,N_4095,N_4300);
nand U5897 (N_5897,N_4098,N_4278);
nor U5898 (N_5898,N_4421,N_4626);
and U5899 (N_5899,N_4122,N_4681);
and U5900 (N_5900,N_4542,N_4296);
nand U5901 (N_5901,N_4514,N_4881);
or U5902 (N_5902,N_4093,N_4404);
nor U5903 (N_5903,N_4159,N_4339);
xnor U5904 (N_5904,N_4650,N_4681);
and U5905 (N_5905,N_4131,N_4573);
and U5906 (N_5906,N_4375,N_4042);
or U5907 (N_5907,N_4300,N_4296);
nor U5908 (N_5908,N_4037,N_4213);
or U5909 (N_5909,N_4531,N_4130);
xnor U5910 (N_5910,N_4548,N_4916);
and U5911 (N_5911,N_4591,N_4131);
and U5912 (N_5912,N_4123,N_4361);
nand U5913 (N_5913,N_4868,N_4332);
or U5914 (N_5914,N_4339,N_4907);
and U5915 (N_5915,N_4163,N_4460);
xor U5916 (N_5916,N_4710,N_4369);
xor U5917 (N_5917,N_4356,N_4431);
nor U5918 (N_5918,N_4417,N_4289);
xnor U5919 (N_5919,N_4882,N_4019);
or U5920 (N_5920,N_4222,N_4930);
xor U5921 (N_5921,N_4795,N_4684);
nand U5922 (N_5922,N_4798,N_4883);
and U5923 (N_5923,N_4999,N_4466);
xnor U5924 (N_5924,N_4812,N_4636);
or U5925 (N_5925,N_4100,N_4752);
or U5926 (N_5926,N_4459,N_4284);
nand U5927 (N_5927,N_4318,N_4443);
nand U5928 (N_5928,N_4227,N_4953);
nand U5929 (N_5929,N_4266,N_4937);
xnor U5930 (N_5930,N_4192,N_4096);
nand U5931 (N_5931,N_4509,N_4978);
nor U5932 (N_5932,N_4076,N_4837);
nand U5933 (N_5933,N_4803,N_4770);
and U5934 (N_5934,N_4492,N_4009);
and U5935 (N_5935,N_4128,N_4650);
xor U5936 (N_5936,N_4681,N_4526);
or U5937 (N_5937,N_4344,N_4362);
and U5938 (N_5938,N_4539,N_4475);
xor U5939 (N_5939,N_4907,N_4817);
or U5940 (N_5940,N_4335,N_4152);
nand U5941 (N_5941,N_4640,N_4616);
and U5942 (N_5942,N_4115,N_4765);
or U5943 (N_5943,N_4688,N_4171);
nor U5944 (N_5944,N_4838,N_4369);
nand U5945 (N_5945,N_4152,N_4389);
or U5946 (N_5946,N_4790,N_4012);
and U5947 (N_5947,N_4197,N_4221);
nor U5948 (N_5948,N_4359,N_4566);
and U5949 (N_5949,N_4789,N_4655);
nor U5950 (N_5950,N_4396,N_4325);
or U5951 (N_5951,N_4902,N_4282);
xor U5952 (N_5952,N_4474,N_4827);
or U5953 (N_5953,N_4493,N_4010);
nand U5954 (N_5954,N_4529,N_4090);
nor U5955 (N_5955,N_4310,N_4865);
nor U5956 (N_5956,N_4253,N_4387);
nor U5957 (N_5957,N_4158,N_4318);
nand U5958 (N_5958,N_4011,N_4736);
xor U5959 (N_5959,N_4536,N_4394);
and U5960 (N_5960,N_4987,N_4118);
nor U5961 (N_5961,N_4096,N_4141);
nand U5962 (N_5962,N_4640,N_4577);
xnor U5963 (N_5963,N_4240,N_4170);
or U5964 (N_5964,N_4202,N_4755);
or U5965 (N_5965,N_4556,N_4285);
xor U5966 (N_5966,N_4675,N_4200);
nand U5967 (N_5967,N_4955,N_4685);
nor U5968 (N_5968,N_4054,N_4146);
and U5969 (N_5969,N_4065,N_4082);
nor U5970 (N_5970,N_4446,N_4770);
xnor U5971 (N_5971,N_4233,N_4633);
nor U5972 (N_5972,N_4518,N_4381);
nor U5973 (N_5973,N_4919,N_4476);
nand U5974 (N_5974,N_4723,N_4822);
or U5975 (N_5975,N_4391,N_4509);
nand U5976 (N_5976,N_4677,N_4633);
nor U5977 (N_5977,N_4734,N_4586);
and U5978 (N_5978,N_4011,N_4991);
nand U5979 (N_5979,N_4312,N_4974);
xnor U5980 (N_5980,N_4497,N_4550);
and U5981 (N_5981,N_4006,N_4436);
xnor U5982 (N_5982,N_4316,N_4853);
and U5983 (N_5983,N_4334,N_4985);
xor U5984 (N_5984,N_4202,N_4389);
or U5985 (N_5985,N_4855,N_4487);
xor U5986 (N_5986,N_4923,N_4041);
and U5987 (N_5987,N_4348,N_4809);
nor U5988 (N_5988,N_4363,N_4218);
nor U5989 (N_5989,N_4887,N_4191);
nand U5990 (N_5990,N_4519,N_4729);
nand U5991 (N_5991,N_4969,N_4522);
and U5992 (N_5992,N_4457,N_4741);
nand U5993 (N_5993,N_4673,N_4563);
nand U5994 (N_5994,N_4178,N_4598);
or U5995 (N_5995,N_4185,N_4749);
or U5996 (N_5996,N_4422,N_4500);
xor U5997 (N_5997,N_4726,N_4483);
xnor U5998 (N_5998,N_4403,N_4818);
or U5999 (N_5999,N_4829,N_4388);
nand U6000 (N_6000,N_5748,N_5606);
and U6001 (N_6001,N_5876,N_5611);
or U6002 (N_6002,N_5805,N_5739);
nor U6003 (N_6003,N_5548,N_5459);
and U6004 (N_6004,N_5615,N_5492);
nand U6005 (N_6005,N_5896,N_5682);
nand U6006 (N_6006,N_5849,N_5484);
nor U6007 (N_6007,N_5861,N_5730);
xnor U6008 (N_6008,N_5160,N_5802);
nand U6009 (N_6009,N_5393,N_5737);
or U6010 (N_6010,N_5817,N_5267);
and U6011 (N_6011,N_5237,N_5708);
xnor U6012 (N_6012,N_5847,N_5519);
nor U6013 (N_6013,N_5518,N_5418);
and U6014 (N_6014,N_5116,N_5703);
or U6015 (N_6015,N_5029,N_5061);
nor U6016 (N_6016,N_5932,N_5069);
nor U6017 (N_6017,N_5774,N_5115);
nand U6018 (N_6018,N_5996,N_5335);
or U6019 (N_6019,N_5507,N_5389);
xor U6020 (N_6020,N_5401,N_5362);
nor U6021 (N_6021,N_5411,N_5537);
nor U6022 (N_6022,N_5469,N_5063);
or U6023 (N_6023,N_5946,N_5030);
or U6024 (N_6024,N_5648,N_5617);
nand U6025 (N_6025,N_5587,N_5008);
nand U6026 (N_6026,N_5625,N_5435);
xnor U6027 (N_6027,N_5300,N_5917);
nand U6028 (N_6028,N_5409,N_5341);
nor U6029 (N_6029,N_5099,N_5466);
xnor U6030 (N_6030,N_5463,N_5542);
xor U6031 (N_6031,N_5428,N_5727);
nand U6032 (N_6032,N_5568,N_5779);
xnor U6033 (N_6033,N_5177,N_5743);
nor U6034 (N_6034,N_5833,N_5502);
nand U6035 (N_6035,N_5759,N_5270);
nor U6036 (N_6036,N_5578,N_5642);
nor U6037 (N_6037,N_5051,N_5485);
nand U6038 (N_6038,N_5747,N_5071);
or U6039 (N_6039,N_5574,N_5208);
and U6040 (N_6040,N_5266,N_5149);
nor U6041 (N_6041,N_5910,N_5718);
nand U6042 (N_6042,N_5624,N_5764);
nor U6043 (N_6043,N_5607,N_5262);
and U6044 (N_6044,N_5991,N_5369);
or U6045 (N_6045,N_5470,N_5550);
and U6046 (N_6046,N_5480,N_5877);
or U6047 (N_6047,N_5514,N_5521);
or U6048 (N_6048,N_5738,N_5289);
xnor U6049 (N_6049,N_5556,N_5448);
xor U6050 (N_6050,N_5155,N_5186);
or U6051 (N_6051,N_5583,N_5807);
and U6052 (N_6052,N_5082,N_5026);
nand U6053 (N_6053,N_5422,N_5723);
nand U6054 (N_6054,N_5992,N_5894);
nor U6055 (N_6055,N_5602,N_5250);
nor U6056 (N_6056,N_5698,N_5693);
or U6057 (N_6057,N_5049,N_5908);
and U6058 (N_6058,N_5786,N_5742);
or U6059 (N_6059,N_5076,N_5810);
xor U6060 (N_6060,N_5150,N_5661);
nor U6061 (N_6061,N_5206,N_5925);
xor U6062 (N_6062,N_5856,N_5359);
nand U6063 (N_6063,N_5001,N_5596);
nand U6064 (N_6064,N_5103,N_5032);
nand U6065 (N_6065,N_5784,N_5880);
and U6066 (N_6066,N_5950,N_5702);
nand U6067 (N_6067,N_5223,N_5960);
nor U6068 (N_6068,N_5151,N_5651);
xnor U6069 (N_6069,N_5399,N_5348);
nor U6070 (N_6070,N_5656,N_5553);
or U6071 (N_6071,N_5516,N_5719);
nand U6072 (N_6072,N_5573,N_5357);
nor U6073 (N_6073,N_5888,N_5456);
and U6074 (N_6074,N_5654,N_5226);
or U6075 (N_6075,N_5512,N_5923);
or U6076 (N_6076,N_5787,N_5387);
xnor U6077 (N_6077,N_5557,N_5334);
xor U6078 (N_6078,N_5249,N_5709);
and U6079 (N_6079,N_5394,N_5102);
nand U6080 (N_6080,N_5958,N_5373);
xnor U6081 (N_6081,N_5461,N_5294);
and U6082 (N_6082,N_5004,N_5318);
nand U6083 (N_6083,N_5586,N_5258);
nor U6084 (N_6084,N_5870,N_5215);
nand U6085 (N_6085,N_5581,N_5424);
and U6086 (N_6086,N_5660,N_5707);
nor U6087 (N_6087,N_5655,N_5980);
nand U6088 (N_6088,N_5343,N_5280);
or U6089 (N_6089,N_5657,N_5639);
nor U6090 (N_6090,N_5506,N_5672);
and U6091 (N_6091,N_5021,N_5563);
nor U6092 (N_6092,N_5153,N_5798);
nor U6093 (N_6093,N_5644,N_5228);
nor U6094 (N_6094,N_5746,N_5057);
and U6095 (N_6095,N_5229,N_5033);
nand U6096 (N_6096,N_5475,N_5489);
nor U6097 (N_6097,N_5398,N_5246);
nor U6098 (N_6098,N_5388,N_5821);
and U6099 (N_6099,N_5257,N_5814);
nand U6100 (N_6100,N_5011,N_5264);
nand U6101 (N_6101,N_5451,N_5086);
or U6102 (N_6102,N_5575,N_5791);
xnor U6103 (N_6103,N_5652,N_5555);
or U6104 (N_6104,N_5241,N_5909);
nand U6105 (N_6105,N_5536,N_5981);
nor U6106 (N_6106,N_5332,N_5097);
or U6107 (N_6107,N_5945,N_5193);
nand U6108 (N_6108,N_5982,N_5538);
or U6109 (N_6109,N_5533,N_5181);
or U6110 (N_6110,N_5785,N_5064);
nand U6111 (N_6111,N_5647,N_5970);
nand U6112 (N_6112,N_5105,N_5751);
and U6113 (N_6113,N_5315,N_5460);
nand U6114 (N_6114,N_5919,N_5618);
xor U6115 (N_6115,N_5288,N_5783);
and U6116 (N_6116,N_5975,N_5331);
nor U6117 (N_6117,N_5501,N_5118);
and U6118 (N_6118,N_5454,N_5998);
xnor U6119 (N_6119,N_5349,N_5361);
xnor U6120 (N_6120,N_5132,N_5094);
xor U6121 (N_6121,N_5564,N_5733);
or U6122 (N_6122,N_5230,N_5579);
or U6123 (N_6123,N_5715,N_5859);
or U6124 (N_6124,N_5952,N_5036);
xor U6125 (N_6125,N_5614,N_5570);
nor U6126 (N_6126,N_5845,N_5217);
or U6127 (N_6127,N_5942,N_5420);
or U6128 (N_6128,N_5993,N_5732);
xor U6129 (N_6129,N_5199,N_5117);
and U6130 (N_6130,N_5902,N_5872);
nor U6131 (N_6131,N_5951,N_5749);
nor U6132 (N_6132,N_5178,N_5121);
and U6133 (N_6133,N_5678,N_5884);
and U6134 (N_6134,N_5256,N_5493);
nor U6135 (N_6135,N_5754,N_5515);
xnor U6136 (N_6136,N_5308,N_5436);
nor U6137 (N_6137,N_5559,N_5297);
xor U6138 (N_6138,N_5056,N_5898);
nor U6139 (N_6139,N_5948,N_5365);
nand U6140 (N_6140,N_5292,N_5142);
nor U6141 (N_6141,N_5963,N_5277);
or U6142 (N_6142,N_5628,N_5453);
xor U6143 (N_6143,N_5402,N_5773);
nand U6144 (N_6144,N_5758,N_5200);
nor U6145 (N_6145,N_5159,N_5728);
xor U6146 (N_6146,N_5174,N_5584);
or U6147 (N_6147,N_5854,N_5075);
and U6148 (N_6148,N_5320,N_5949);
xnor U6149 (N_6149,N_5106,N_5846);
or U6150 (N_6150,N_5700,N_5901);
nor U6151 (N_6151,N_5911,N_5552);
nor U6152 (N_6152,N_5310,N_5216);
nand U6153 (N_6153,N_5044,N_5120);
and U6154 (N_6154,N_5377,N_5168);
xnor U6155 (N_6155,N_5471,N_5676);
nand U6156 (N_6156,N_5410,N_5491);
nand U6157 (N_6157,N_5209,N_5313);
or U6158 (N_6158,N_5601,N_5458);
nand U6159 (N_6159,N_5776,N_5190);
or U6160 (N_6160,N_5858,N_5825);
nand U6161 (N_6161,N_5598,N_5195);
xnor U6162 (N_6162,N_5765,N_5412);
nor U6163 (N_6163,N_5650,N_5176);
or U6164 (N_6164,N_5885,N_5772);
or U6165 (N_6165,N_5148,N_5081);
or U6166 (N_6166,N_5203,N_5599);
or U6167 (N_6167,N_5572,N_5353);
nor U6168 (N_6168,N_5287,N_5042);
nand U6169 (N_6169,N_5452,N_5824);
nand U6170 (N_6170,N_5760,N_5182);
and U6171 (N_6171,N_5561,N_5281);
xnor U6172 (N_6172,N_5803,N_5843);
or U6173 (N_6173,N_5173,N_5595);
or U6174 (N_6174,N_5590,N_5705);
xor U6175 (N_6175,N_5073,N_5558);
xor U6176 (N_6176,N_5517,N_5423);
nand U6177 (N_6177,N_5272,N_5851);
nor U6178 (N_6178,N_5816,N_5804);
and U6179 (N_6179,N_5878,N_5594);
nor U6180 (N_6180,N_5867,N_5696);
and U6181 (N_6181,N_5122,N_5988);
and U6182 (N_6182,N_5285,N_5974);
xnor U6183 (N_6183,N_5721,N_5665);
and U6184 (N_6184,N_5442,N_5311);
nand U6185 (N_6185,N_5457,N_5662);
or U6186 (N_6186,N_5140,N_5890);
or U6187 (N_6187,N_5383,N_5834);
or U6188 (N_6188,N_5937,N_5395);
nor U6189 (N_6189,N_5408,N_5242);
or U6190 (N_6190,N_5013,N_5669);
or U6191 (N_6191,N_5392,N_5130);
nor U6192 (N_6192,N_5571,N_5585);
or U6193 (N_6193,N_5244,N_5014);
xor U6194 (N_6194,N_5124,N_5670);
xor U6195 (N_6195,N_5767,N_5995);
nor U6196 (N_6196,N_5068,N_5179);
and U6197 (N_6197,N_5938,N_5936);
nor U6198 (N_6198,N_5712,N_5820);
nor U6199 (N_6199,N_5694,N_5447);
nor U6200 (N_6200,N_5350,N_5808);
xnor U6201 (N_6201,N_5291,N_5110);
nor U6202 (N_6202,N_5797,N_5508);
nand U6203 (N_6203,N_5455,N_5218);
nand U6204 (N_6204,N_5905,N_5915);
and U6205 (N_6205,N_5464,N_5054);
and U6206 (N_6206,N_5616,N_5818);
or U6207 (N_6207,N_5080,N_5416);
and U6208 (N_6208,N_5681,N_5828);
xor U6209 (N_6209,N_5725,N_5243);
xnor U6210 (N_6210,N_5795,N_5089);
nor U6211 (N_6211,N_5701,N_5074);
or U6212 (N_6212,N_5539,N_5477);
nand U6213 (N_6213,N_5969,N_5328);
nand U6214 (N_6214,N_5697,N_5158);
xor U6215 (N_6215,N_5207,N_5303);
and U6216 (N_6216,N_5113,N_5037);
nand U6217 (N_6217,N_5873,N_5293);
xnor U6218 (N_6218,N_5695,N_5830);
xnor U6219 (N_6219,N_5138,N_5222);
xnor U6220 (N_6220,N_5666,N_5378);
and U6221 (N_6221,N_5630,N_5340);
xnor U6222 (N_6222,N_5147,N_5683);
xor U6223 (N_6223,N_5520,N_5576);
and U6224 (N_6224,N_5108,N_5253);
nand U6225 (N_6225,N_5490,N_5112);
xor U6226 (N_6226,N_5835,N_5499);
nor U6227 (N_6227,N_5675,N_5941);
xnor U6228 (N_6228,N_5005,N_5994);
or U6229 (N_6229,N_5417,N_5819);
nand U6230 (N_6230,N_5944,N_5227);
or U6231 (N_6231,N_5545,N_5511);
xor U6232 (N_6232,N_5114,N_5312);
and U6233 (N_6233,N_5871,N_5525);
xor U6234 (N_6234,N_5922,N_5636);
or U6235 (N_6235,N_5734,N_5437);
xor U6236 (N_6236,N_5531,N_5523);
xor U6237 (N_6237,N_5726,N_5175);
xor U6238 (N_6238,N_5473,N_5360);
and U6239 (N_6239,N_5366,N_5146);
and U6240 (N_6240,N_5079,N_5775);
xor U6241 (N_6241,N_5481,N_5342);
xnor U6242 (N_6242,N_5986,N_5035);
and U6243 (N_6243,N_5107,N_5060);
and U6244 (N_6244,N_5263,N_5663);
and U6245 (N_6245,N_5188,N_5326);
or U6246 (N_6246,N_5842,N_5918);
nand U6247 (N_6247,N_5164,N_5434);
xor U6248 (N_6248,N_5391,N_5192);
xor U6249 (N_6249,N_5157,N_5731);
or U6250 (N_6250,N_5716,N_5488);
and U6251 (N_6251,N_5770,N_5866);
and U6252 (N_6252,N_5649,N_5900);
xor U6253 (N_6253,N_5282,N_5827);
or U6254 (N_6254,N_5848,N_5893);
xor U6255 (N_6255,N_5510,N_5962);
nand U6256 (N_6256,N_5184,N_5381);
nand U6257 (N_6257,N_5926,N_5686);
nand U6258 (N_6258,N_5319,N_5710);
nor U6259 (N_6259,N_5083,N_5432);
xor U6260 (N_6260,N_5677,N_5997);
and U6261 (N_6261,N_5687,N_5643);
nand U6262 (N_6262,N_5100,N_5912);
and U6263 (N_6263,N_5966,N_5498);
nand U6264 (N_6264,N_5284,N_5714);
and U6265 (N_6265,N_5443,N_5012);
and U6266 (N_6266,N_5474,N_5674);
nand U6267 (N_6267,N_5736,N_5028);
nand U6268 (N_6268,N_5935,N_5528);
xor U6269 (N_6269,N_5892,N_5055);
nand U6270 (N_6270,N_5375,N_5251);
nor U6271 (N_6271,N_5141,N_5245);
and U6272 (N_6272,N_5761,N_5809);
nand U6273 (N_6273,N_5792,N_5296);
and U6274 (N_6274,N_5123,N_5125);
nand U6275 (N_6275,N_5831,N_5367);
nand U6276 (N_6276,N_5968,N_5077);
nor U6277 (N_6277,N_5009,N_5449);
or U6278 (N_6278,N_5431,N_5608);
nor U6279 (N_6279,N_5047,N_5984);
and U6280 (N_6280,N_5302,N_5019);
xnor U6281 (N_6281,N_5371,N_5172);
nor U6282 (N_6282,N_5439,N_5865);
nand U6283 (N_6283,N_5713,N_5956);
xor U6284 (N_6284,N_5541,N_5104);
nor U6285 (N_6285,N_5039,N_5622);
xnor U6286 (N_6286,N_5560,N_5197);
and U6287 (N_6287,N_5554,N_5777);
xnor U6288 (N_6288,N_5165,N_5605);
and U6289 (N_6289,N_5863,N_5619);
nor U6290 (N_6290,N_5330,N_5487);
nor U6291 (N_6291,N_5384,N_5862);
nand U6292 (N_6292,N_5352,N_5048);
or U6293 (N_6293,N_5635,N_5221);
nand U6294 (N_6294,N_5040,N_5626);
or U6295 (N_6295,N_5852,N_5279);
nand U6296 (N_6296,N_5347,N_5129);
xnor U6297 (N_6297,N_5839,N_5766);
xnor U6298 (N_6298,N_5806,N_5868);
xnor U6299 (N_6299,N_5844,N_5641);
or U6300 (N_6300,N_5170,N_5569);
xor U6301 (N_6301,N_5610,N_5390);
xnor U6302 (N_6302,N_5904,N_5465);
or U6303 (N_6303,N_5685,N_5419);
nand U6304 (N_6304,N_5066,N_5756);
nand U6305 (N_6305,N_5653,N_5058);
and U6306 (N_6306,N_5143,N_5532);
and U6307 (N_6307,N_5495,N_5017);
nand U6308 (N_6308,N_5169,N_5881);
nor U6309 (N_6309,N_5977,N_5233);
nand U6310 (N_6310,N_5278,N_5396);
xnor U6311 (N_6311,N_5634,N_5087);
and U6312 (N_6312,N_5000,N_5788);
nor U6313 (N_6313,N_5438,N_5943);
xnor U6314 (N_6314,N_5162,N_5692);
or U6315 (N_6315,N_5065,N_5078);
xnor U6316 (N_6316,N_5236,N_5961);
nand U6317 (N_6317,N_5750,N_5543);
and U6318 (N_6318,N_5582,N_5689);
and U6319 (N_6319,N_5631,N_5535);
nor U6320 (N_6320,N_5126,N_5400);
or U6321 (N_6321,N_5358,N_5680);
xor U6322 (N_6322,N_5038,N_5671);
nand U6323 (N_6323,N_5346,N_5240);
or U6324 (N_6324,N_5811,N_5603);
and U6325 (N_6325,N_5006,N_5658);
xor U6326 (N_6326,N_5837,N_5397);
or U6327 (N_6327,N_5214,N_5052);
and U6328 (N_6328,N_5462,N_5796);
xor U6329 (N_6329,N_5500,N_5530);
xor U6330 (N_6330,N_5134,N_5668);
and U6331 (N_6331,N_5740,N_5762);
and U6332 (N_6332,N_5972,N_5540);
nand U6333 (N_6333,N_5374,N_5566);
or U6334 (N_6334,N_5957,N_5815);
or U6335 (N_6335,N_5985,N_5920);
and U6336 (N_6336,N_5025,N_5735);
or U6337 (N_6337,N_5522,N_5385);
nor U6338 (N_6338,N_5154,N_5415);
nor U6339 (N_6339,N_5973,N_5916);
and U6340 (N_6340,N_5684,N_5934);
xnor U6341 (N_6341,N_5212,N_5646);
and U6342 (N_6342,N_5053,N_5673);
nor U6343 (N_6343,N_5483,N_5370);
or U6344 (N_6344,N_5494,N_5265);
nand U6345 (N_6345,N_5092,N_5043);
or U6346 (N_6346,N_5664,N_5260);
nand U6347 (N_6347,N_5829,N_5298);
and U6348 (N_6348,N_5379,N_5185);
nand U6349 (N_6349,N_5794,N_5131);
or U6350 (N_6350,N_5755,N_5597);
or U6351 (N_6351,N_5426,N_5799);
and U6352 (N_6352,N_5007,N_5269);
nand U6353 (N_6353,N_5921,N_5273);
xor U6354 (N_6354,N_5304,N_5156);
or U6355 (N_6355,N_5355,N_5745);
xor U6356 (N_6356,N_5505,N_5429);
xor U6357 (N_6357,N_5826,N_5836);
and U6358 (N_6358,N_5874,N_5382);
nor U6359 (N_6359,N_5201,N_5857);
or U6360 (N_6360,N_5204,N_5580);
nor U6361 (N_6361,N_5577,N_5592);
nor U6362 (N_6362,N_5220,N_5768);
xnor U6363 (N_6363,N_5299,N_5210);
nor U6364 (N_6364,N_5720,N_5235);
and U6365 (N_6365,N_5440,N_5368);
nor U6366 (N_6366,N_5546,N_5327);
and U6367 (N_6367,N_5386,N_5933);
and U6368 (N_6368,N_5274,N_5213);
xnor U6369 (N_6369,N_5699,N_5329);
nor U6370 (N_6370,N_5659,N_5822);
nor U6371 (N_6371,N_5899,N_5345);
xor U6372 (N_6372,N_5813,N_5119);
nor U6373 (N_6373,N_5414,N_5072);
or U6374 (N_6374,N_5152,N_5476);
nand U6375 (N_6375,N_5959,N_5321);
nand U6376 (N_6376,N_5145,N_5224);
nor U6377 (N_6377,N_5163,N_5180);
xnor U6378 (N_6378,N_5316,N_5838);
or U6379 (N_6379,N_5351,N_5924);
nor U6380 (N_6380,N_5513,N_5724);
and U6381 (N_6381,N_5137,N_5247);
nor U6382 (N_6382,N_5363,N_5046);
or U6383 (N_6383,N_5887,N_5623);
or U6384 (N_6384,N_5613,N_5248);
nor U6385 (N_6385,N_5301,N_5782);
or U6386 (N_6386,N_5380,N_5059);
xor U6387 (N_6387,N_5015,N_5403);
nor U6388 (N_6388,N_5927,N_5612);
or U6389 (N_6389,N_5620,N_5627);
xnor U6390 (N_6390,N_5551,N_5679);
and U6391 (N_6391,N_5793,N_5196);
xor U6392 (N_6392,N_5914,N_5407);
xnor U6393 (N_6393,N_5205,N_5339);
xor U6394 (N_6394,N_5840,N_5913);
or U6395 (N_6395,N_5855,N_5161);
or U6396 (N_6396,N_5085,N_5018);
nor U6397 (N_6397,N_5166,N_5978);
nor U6398 (N_6398,N_5589,N_5729);
xnor U6399 (N_6399,N_5479,N_5769);
nor U6400 (N_6400,N_5633,N_5562);
or U6401 (N_6401,N_5882,N_5259);
or U6402 (N_6402,N_5929,N_5691);
nor U6403 (N_6403,N_5983,N_5413);
nand U6404 (N_6404,N_5433,N_5955);
and U6405 (N_6405,N_5144,N_5023);
xor U6406 (N_6406,N_5717,N_5780);
and U6407 (N_6407,N_5534,N_5690);
and U6408 (N_6408,N_5907,N_5964);
or U6409 (N_6409,N_5781,N_5979);
nand U6410 (N_6410,N_5041,N_5305);
xnor U6411 (N_6411,N_5869,N_5632);
or U6412 (N_6412,N_5020,N_5090);
or U6413 (N_6413,N_5875,N_5275);
or U6414 (N_6414,N_5128,N_5939);
xnor U6415 (N_6415,N_5406,N_5045);
nor U6416 (N_6416,N_5812,N_5325);
xnor U6417 (N_6417,N_5999,N_5763);
or U6418 (N_6418,N_5309,N_5093);
xnor U6419 (N_6419,N_5832,N_5372);
and U6420 (N_6420,N_5976,N_5771);
and U6421 (N_6421,N_5135,N_5096);
nand U6422 (N_6422,N_5971,N_5405);
nor U6423 (N_6423,N_5593,N_5640);
and U6424 (N_6424,N_5027,N_5290);
nand U6425 (N_6425,N_5283,N_5084);
xnor U6426 (N_6426,N_5404,N_5527);
nor U6427 (N_6427,N_5189,N_5338);
or U6428 (N_6428,N_5268,N_5789);
xnor U6429 (N_6429,N_5091,N_5940);
nand U6430 (N_6430,N_5688,N_5198);
nand U6431 (N_6431,N_5895,N_5778);
and U6432 (N_6432,N_5741,N_5127);
xor U6433 (N_6433,N_5050,N_5067);
xnor U6434 (N_6434,N_5600,N_5286);
xor U6435 (N_6435,N_5194,N_5202);
or U6436 (N_6436,N_5211,N_5706);
nor U6437 (N_6437,N_5823,N_5930);
or U6438 (N_6438,N_5095,N_5232);
nand U6439 (N_6439,N_5482,N_5897);
or U6440 (N_6440,N_5790,N_5171);
xnor U6441 (N_6441,N_5990,N_5967);
and U6442 (N_6442,N_5234,N_5864);
nand U6443 (N_6443,N_5139,N_5883);
nor U6444 (N_6444,N_5609,N_5003);
nor U6445 (N_6445,N_5167,N_5191);
nand U6446 (N_6446,N_5239,N_5101);
and U6447 (N_6447,N_5133,N_5800);
or U6448 (N_6448,N_5062,N_5906);
or U6449 (N_6449,N_5421,N_5376);
and U6450 (N_6450,N_5031,N_5989);
nor U6451 (N_6451,N_5509,N_5441);
and U6452 (N_6452,N_5987,N_5947);
nor U6453 (N_6453,N_5010,N_5891);
nand U6454 (N_6454,N_5588,N_5444);
nand U6455 (N_6455,N_5954,N_5529);
xor U6456 (N_6456,N_5344,N_5238);
or U6457 (N_6457,N_5604,N_5276);
or U6458 (N_6458,N_5109,N_5931);
xor U6459 (N_6459,N_5497,N_5629);
nor U6460 (N_6460,N_5478,N_5903);
nor U6461 (N_6461,N_5841,N_5472);
and U6462 (N_6462,N_5356,N_5953);
and U6463 (N_6463,N_5889,N_5853);
nor U6464 (N_6464,N_5324,N_5486);
or U6465 (N_6465,N_5621,N_5098);
or U6466 (N_6466,N_5744,N_5752);
nand U6467 (N_6467,N_5757,N_5722);
or U6468 (N_6468,N_5271,N_5425);
xor U6469 (N_6469,N_5524,N_5504);
nor U6470 (N_6470,N_5022,N_5430);
nor U6471 (N_6471,N_5704,N_5070);
or U6472 (N_6472,N_5468,N_5591);
nand U6473 (N_6473,N_5467,N_5252);
or U6474 (N_6474,N_5231,N_5337);
nand U6475 (N_6475,N_5547,N_5333);
xor U6476 (N_6476,N_5567,N_5496);
nor U6477 (N_6477,N_5034,N_5450);
xnor U6478 (N_6478,N_5753,N_5427);
and U6479 (N_6479,N_5336,N_5850);
nor U6480 (N_6480,N_5354,N_5801);
nand U6481 (N_6481,N_5645,N_5317);
nand U6482 (N_6482,N_5183,N_5024);
and U6483 (N_6483,N_5323,N_5886);
xor U6484 (N_6484,N_5965,N_5503);
or U6485 (N_6485,N_5261,N_5219);
xnor U6486 (N_6486,N_5637,N_5136);
or U6487 (N_6487,N_5565,N_5016);
or U6488 (N_6488,N_5002,N_5306);
and U6489 (N_6489,N_5111,N_5314);
or U6490 (N_6490,N_5860,N_5446);
or U6491 (N_6491,N_5928,N_5307);
nand U6492 (N_6492,N_5445,N_5544);
xnor U6493 (N_6493,N_5879,N_5187);
xnor U6494 (N_6494,N_5254,N_5711);
or U6495 (N_6495,N_5225,N_5526);
or U6496 (N_6496,N_5667,N_5088);
or U6497 (N_6497,N_5255,N_5295);
xor U6498 (N_6498,N_5364,N_5322);
and U6499 (N_6499,N_5638,N_5549);
nor U6500 (N_6500,N_5934,N_5825);
nand U6501 (N_6501,N_5733,N_5888);
or U6502 (N_6502,N_5695,N_5397);
nor U6503 (N_6503,N_5273,N_5073);
nand U6504 (N_6504,N_5817,N_5729);
or U6505 (N_6505,N_5947,N_5135);
and U6506 (N_6506,N_5615,N_5433);
xor U6507 (N_6507,N_5389,N_5116);
and U6508 (N_6508,N_5190,N_5223);
nor U6509 (N_6509,N_5627,N_5764);
nand U6510 (N_6510,N_5611,N_5323);
and U6511 (N_6511,N_5772,N_5120);
xnor U6512 (N_6512,N_5455,N_5803);
and U6513 (N_6513,N_5505,N_5717);
or U6514 (N_6514,N_5289,N_5181);
and U6515 (N_6515,N_5169,N_5264);
nand U6516 (N_6516,N_5005,N_5368);
nor U6517 (N_6517,N_5323,N_5412);
and U6518 (N_6518,N_5857,N_5139);
nor U6519 (N_6519,N_5918,N_5620);
nor U6520 (N_6520,N_5388,N_5859);
nor U6521 (N_6521,N_5687,N_5974);
and U6522 (N_6522,N_5084,N_5202);
nor U6523 (N_6523,N_5549,N_5273);
xor U6524 (N_6524,N_5537,N_5253);
and U6525 (N_6525,N_5204,N_5284);
nor U6526 (N_6526,N_5162,N_5995);
or U6527 (N_6527,N_5392,N_5969);
xnor U6528 (N_6528,N_5497,N_5043);
nand U6529 (N_6529,N_5930,N_5235);
or U6530 (N_6530,N_5431,N_5179);
nand U6531 (N_6531,N_5387,N_5209);
or U6532 (N_6532,N_5427,N_5990);
and U6533 (N_6533,N_5208,N_5180);
xnor U6534 (N_6534,N_5293,N_5390);
or U6535 (N_6535,N_5248,N_5566);
xor U6536 (N_6536,N_5677,N_5800);
or U6537 (N_6537,N_5871,N_5530);
nand U6538 (N_6538,N_5980,N_5005);
xor U6539 (N_6539,N_5046,N_5337);
or U6540 (N_6540,N_5075,N_5454);
xnor U6541 (N_6541,N_5870,N_5657);
nand U6542 (N_6542,N_5836,N_5046);
nor U6543 (N_6543,N_5373,N_5621);
nand U6544 (N_6544,N_5560,N_5687);
and U6545 (N_6545,N_5409,N_5636);
or U6546 (N_6546,N_5348,N_5043);
nor U6547 (N_6547,N_5442,N_5586);
xor U6548 (N_6548,N_5121,N_5248);
and U6549 (N_6549,N_5423,N_5365);
xnor U6550 (N_6550,N_5240,N_5078);
nor U6551 (N_6551,N_5108,N_5839);
and U6552 (N_6552,N_5684,N_5222);
and U6553 (N_6553,N_5649,N_5864);
and U6554 (N_6554,N_5554,N_5219);
nand U6555 (N_6555,N_5460,N_5481);
nand U6556 (N_6556,N_5778,N_5789);
xor U6557 (N_6557,N_5030,N_5660);
nand U6558 (N_6558,N_5865,N_5459);
and U6559 (N_6559,N_5404,N_5418);
xnor U6560 (N_6560,N_5882,N_5126);
nor U6561 (N_6561,N_5990,N_5810);
or U6562 (N_6562,N_5841,N_5972);
or U6563 (N_6563,N_5763,N_5727);
nand U6564 (N_6564,N_5536,N_5623);
and U6565 (N_6565,N_5343,N_5498);
nand U6566 (N_6566,N_5520,N_5414);
nor U6567 (N_6567,N_5888,N_5423);
or U6568 (N_6568,N_5575,N_5321);
or U6569 (N_6569,N_5388,N_5504);
or U6570 (N_6570,N_5712,N_5294);
nand U6571 (N_6571,N_5290,N_5742);
nor U6572 (N_6572,N_5809,N_5196);
and U6573 (N_6573,N_5904,N_5017);
nand U6574 (N_6574,N_5120,N_5900);
or U6575 (N_6575,N_5382,N_5506);
or U6576 (N_6576,N_5725,N_5445);
nor U6577 (N_6577,N_5798,N_5583);
xor U6578 (N_6578,N_5266,N_5938);
and U6579 (N_6579,N_5093,N_5703);
or U6580 (N_6580,N_5365,N_5903);
nand U6581 (N_6581,N_5273,N_5655);
and U6582 (N_6582,N_5005,N_5691);
nor U6583 (N_6583,N_5838,N_5515);
nor U6584 (N_6584,N_5688,N_5637);
nand U6585 (N_6585,N_5622,N_5970);
and U6586 (N_6586,N_5477,N_5064);
nor U6587 (N_6587,N_5897,N_5614);
xor U6588 (N_6588,N_5253,N_5880);
nor U6589 (N_6589,N_5918,N_5494);
or U6590 (N_6590,N_5378,N_5633);
nor U6591 (N_6591,N_5818,N_5233);
xnor U6592 (N_6592,N_5745,N_5361);
xor U6593 (N_6593,N_5344,N_5025);
or U6594 (N_6594,N_5570,N_5158);
and U6595 (N_6595,N_5241,N_5575);
nand U6596 (N_6596,N_5626,N_5561);
nand U6597 (N_6597,N_5431,N_5279);
nand U6598 (N_6598,N_5467,N_5242);
nor U6599 (N_6599,N_5762,N_5784);
or U6600 (N_6600,N_5364,N_5833);
nor U6601 (N_6601,N_5940,N_5851);
xnor U6602 (N_6602,N_5225,N_5898);
or U6603 (N_6603,N_5613,N_5136);
or U6604 (N_6604,N_5537,N_5428);
nand U6605 (N_6605,N_5736,N_5149);
nand U6606 (N_6606,N_5192,N_5153);
xnor U6607 (N_6607,N_5708,N_5497);
xor U6608 (N_6608,N_5461,N_5376);
and U6609 (N_6609,N_5511,N_5843);
nand U6610 (N_6610,N_5946,N_5941);
xnor U6611 (N_6611,N_5838,N_5665);
or U6612 (N_6612,N_5993,N_5819);
xnor U6613 (N_6613,N_5943,N_5311);
xnor U6614 (N_6614,N_5200,N_5601);
or U6615 (N_6615,N_5387,N_5380);
nand U6616 (N_6616,N_5991,N_5973);
nand U6617 (N_6617,N_5134,N_5400);
or U6618 (N_6618,N_5644,N_5420);
nand U6619 (N_6619,N_5958,N_5847);
xnor U6620 (N_6620,N_5513,N_5092);
nor U6621 (N_6621,N_5936,N_5790);
and U6622 (N_6622,N_5479,N_5070);
nand U6623 (N_6623,N_5906,N_5138);
or U6624 (N_6624,N_5647,N_5568);
xnor U6625 (N_6625,N_5693,N_5674);
xor U6626 (N_6626,N_5240,N_5732);
nor U6627 (N_6627,N_5323,N_5687);
or U6628 (N_6628,N_5628,N_5902);
nor U6629 (N_6629,N_5180,N_5401);
nand U6630 (N_6630,N_5730,N_5576);
nand U6631 (N_6631,N_5372,N_5611);
nand U6632 (N_6632,N_5519,N_5332);
nand U6633 (N_6633,N_5440,N_5291);
or U6634 (N_6634,N_5065,N_5235);
nor U6635 (N_6635,N_5385,N_5075);
nand U6636 (N_6636,N_5462,N_5132);
nor U6637 (N_6637,N_5248,N_5474);
and U6638 (N_6638,N_5457,N_5289);
and U6639 (N_6639,N_5396,N_5871);
and U6640 (N_6640,N_5530,N_5526);
nor U6641 (N_6641,N_5863,N_5449);
nand U6642 (N_6642,N_5520,N_5994);
and U6643 (N_6643,N_5030,N_5614);
nand U6644 (N_6644,N_5910,N_5998);
nand U6645 (N_6645,N_5027,N_5311);
xnor U6646 (N_6646,N_5977,N_5680);
nor U6647 (N_6647,N_5663,N_5655);
nand U6648 (N_6648,N_5824,N_5869);
xor U6649 (N_6649,N_5753,N_5740);
and U6650 (N_6650,N_5490,N_5474);
xor U6651 (N_6651,N_5151,N_5733);
and U6652 (N_6652,N_5300,N_5129);
xnor U6653 (N_6653,N_5517,N_5826);
nand U6654 (N_6654,N_5199,N_5878);
or U6655 (N_6655,N_5920,N_5680);
xnor U6656 (N_6656,N_5062,N_5662);
xnor U6657 (N_6657,N_5817,N_5458);
nand U6658 (N_6658,N_5220,N_5815);
or U6659 (N_6659,N_5280,N_5992);
xor U6660 (N_6660,N_5095,N_5759);
nand U6661 (N_6661,N_5817,N_5870);
nor U6662 (N_6662,N_5798,N_5393);
nor U6663 (N_6663,N_5547,N_5863);
nand U6664 (N_6664,N_5074,N_5806);
nor U6665 (N_6665,N_5297,N_5624);
xor U6666 (N_6666,N_5368,N_5846);
and U6667 (N_6667,N_5557,N_5282);
and U6668 (N_6668,N_5822,N_5581);
nand U6669 (N_6669,N_5714,N_5024);
nand U6670 (N_6670,N_5442,N_5451);
and U6671 (N_6671,N_5741,N_5156);
xor U6672 (N_6672,N_5423,N_5989);
nand U6673 (N_6673,N_5620,N_5571);
nand U6674 (N_6674,N_5262,N_5357);
xnor U6675 (N_6675,N_5364,N_5488);
nand U6676 (N_6676,N_5732,N_5986);
or U6677 (N_6677,N_5875,N_5330);
nand U6678 (N_6678,N_5344,N_5505);
xnor U6679 (N_6679,N_5944,N_5745);
xor U6680 (N_6680,N_5476,N_5193);
or U6681 (N_6681,N_5510,N_5606);
or U6682 (N_6682,N_5518,N_5731);
nor U6683 (N_6683,N_5257,N_5902);
nor U6684 (N_6684,N_5655,N_5234);
nand U6685 (N_6685,N_5027,N_5875);
or U6686 (N_6686,N_5866,N_5834);
nor U6687 (N_6687,N_5835,N_5621);
xnor U6688 (N_6688,N_5846,N_5046);
nand U6689 (N_6689,N_5524,N_5055);
and U6690 (N_6690,N_5109,N_5116);
nor U6691 (N_6691,N_5407,N_5051);
or U6692 (N_6692,N_5236,N_5449);
or U6693 (N_6693,N_5094,N_5353);
xnor U6694 (N_6694,N_5309,N_5268);
nand U6695 (N_6695,N_5433,N_5053);
nor U6696 (N_6696,N_5967,N_5880);
or U6697 (N_6697,N_5095,N_5523);
or U6698 (N_6698,N_5380,N_5818);
nand U6699 (N_6699,N_5719,N_5023);
or U6700 (N_6700,N_5486,N_5025);
or U6701 (N_6701,N_5895,N_5568);
nor U6702 (N_6702,N_5842,N_5363);
or U6703 (N_6703,N_5830,N_5714);
nor U6704 (N_6704,N_5913,N_5019);
nor U6705 (N_6705,N_5824,N_5305);
nand U6706 (N_6706,N_5304,N_5703);
nand U6707 (N_6707,N_5952,N_5447);
or U6708 (N_6708,N_5009,N_5102);
and U6709 (N_6709,N_5500,N_5228);
or U6710 (N_6710,N_5245,N_5087);
nor U6711 (N_6711,N_5526,N_5381);
and U6712 (N_6712,N_5801,N_5229);
xor U6713 (N_6713,N_5037,N_5624);
nor U6714 (N_6714,N_5809,N_5859);
nor U6715 (N_6715,N_5033,N_5924);
nand U6716 (N_6716,N_5652,N_5489);
or U6717 (N_6717,N_5410,N_5865);
and U6718 (N_6718,N_5919,N_5852);
or U6719 (N_6719,N_5282,N_5992);
and U6720 (N_6720,N_5002,N_5725);
nand U6721 (N_6721,N_5221,N_5968);
or U6722 (N_6722,N_5472,N_5791);
and U6723 (N_6723,N_5283,N_5740);
and U6724 (N_6724,N_5844,N_5355);
nor U6725 (N_6725,N_5407,N_5752);
xor U6726 (N_6726,N_5367,N_5562);
and U6727 (N_6727,N_5904,N_5325);
nand U6728 (N_6728,N_5881,N_5000);
and U6729 (N_6729,N_5113,N_5330);
and U6730 (N_6730,N_5680,N_5571);
and U6731 (N_6731,N_5983,N_5288);
and U6732 (N_6732,N_5161,N_5008);
nor U6733 (N_6733,N_5446,N_5344);
or U6734 (N_6734,N_5255,N_5490);
or U6735 (N_6735,N_5607,N_5927);
nand U6736 (N_6736,N_5732,N_5997);
or U6737 (N_6737,N_5042,N_5103);
nand U6738 (N_6738,N_5759,N_5094);
xnor U6739 (N_6739,N_5446,N_5761);
and U6740 (N_6740,N_5284,N_5349);
nor U6741 (N_6741,N_5113,N_5123);
nor U6742 (N_6742,N_5711,N_5739);
xor U6743 (N_6743,N_5069,N_5005);
nand U6744 (N_6744,N_5444,N_5058);
nand U6745 (N_6745,N_5779,N_5420);
and U6746 (N_6746,N_5316,N_5479);
or U6747 (N_6747,N_5304,N_5932);
nor U6748 (N_6748,N_5534,N_5766);
and U6749 (N_6749,N_5764,N_5536);
nor U6750 (N_6750,N_5401,N_5508);
or U6751 (N_6751,N_5275,N_5618);
xnor U6752 (N_6752,N_5260,N_5721);
nand U6753 (N_6753,N_5626,N_5663);
and U6754 (N_6754,N_5216,N_5485);
or U6755 (N_6755,N_5900,N_5070);
xnor U6756 (N_6756,N_5634,N_5385);
and U6757 (N_6757,N_5784,N_5066);
nand U6758 (N_6758,N_5780,N_5419);
nand U6759 (N_6759,N_5489,N_5612);
or U6760 (N_6760,N_5942,N_5108);
xnor U6761 (N_6761,N_5424,N_5093);
nor U6762 (N_6762,N_5611,N_5375);
nand U6763 (N_6763,N_5932,N_5186);
or U6764 (N_6764,N_5790,N_5995);
xor U6765 (N_6765,N_5022,N_5087);
or U6766 (N_6766,N_5071,N_5331);
or U6767 (N_6767,N_5723,N_5471);
nor U6768 (N_6768,N_5052,N_5251);
and U6769 (N_6769,N_5903,N_5667);
and U6770 (N_6770,N_5550,N_5788);
nand U6771 (N_6771,N_5098,N_5493);
xor U6772 (N_6772,N_5785,N_5463);
nand U6773 (N_6773,N_5020,N_5567);
xnor U6774 (N_6774,N_5473,N_5336);
and U6775 (N_6775,N_5328,N_5427);
nor U6776 (N_6776,N_5956,N_5105);
or U6777 (N_6777,N_5288,N_5406);
nand U6778 (N_6778,N_5061,N_5830);
and U6779 (N_6779,N_5057,N_5613);
and U6780 (N_6780,N_5557,N_5319);
xor U6781 (N_6781,N_5113,N_5299);
or U6782 (N_6782,N_5671,N_5893);
and U6783 (N_6783,N_5251,N_5959);
or U6784 (N_6784,N_5106,N_5327);
nor U6785 (N_6785,N_5595,N_5640);
nor U6786 (N_6786,N_5506,N_5331);
or U6787 (N_6787,N_5624,N_5377);
nand U6788 (N_6788,N_5580,N_5124);
nand U6789 (N_6789,N_5920,N_5115);
nand U6790 (N_6790,N_5403,N_5069);
nor U6791 (N_6791,N_5048,N_5353);
nor U6792 (N_6792,N_5295,N_5976);
or U6793 (N_6793,N_5359,N_5212);
nor U6794 (N_6794,N_5789,N_5466);
xor U6795 (N_6795,N_5680,N_5268);
nand U6796 (N_6796,N_5912,N_5219);
nor U6797 (N_6797,N_5662,N_5617);
and U6798 (N_6798,N_5168,N_5202);
nand U6799 (N_6799,N_5762,N_5706);
and U6800 (N_6800,N_5818,N_5476);
and U6801 (N_6801,N_5837,N_5235);
nor U6802 (N_6802,N_5472,N_5474);
nor U6803 (N_6803,N_5274,N_5204);
nand U6804 (N_6804,N_5459,N_5654);
nand U6805 (N_6805,N_5761,N_5453);
xnor U6806 (N_6806,N_5541,N_5674);
nand U6807 (N_6807,N_5912,N_5150);
nand U6808 (N_6808,N_5159,N_5532);
xor U6809 (N_6809,N_5180,N_5581);
and U6810 (N_6810,N_5255,N_5412);
xor U6811 (N_6811,N_5755,N_5953);
nand U6812 (N_6812,N_5288,N_5086);
or U6813 (N_6813,N_5888,N_5467);
or U6814 (N_6814,N_5300,N_5223);
and U6815 (N_6815,N_5787,N_5689);
and U6816 (N_6816,N_5921,N_5634);
or U6817 (N_6817,N_5099,N_5005);
nand U6818 (N_6818,N_5902,N_5837);
nor U6819 (N_6819,N_5731,N_5604);
or U6820 (N_6820,N_5236,N_5180);
nand U6821 (N_6821,N_5696,N_5350);
or U6822 (N_6822,N_5048,N_5529);
or U6823 (N_6823,N_5343,N_5604);
nor U6824 (N_6824,N_5538,N_5809);
nand U6825 (N_6825,N_5119,N_5299);
or U6826 (N_6826,N_5831,N_5108);
nor U6827 (N_6827,N_5354,N_5712);
nor U6828 (N_6828,N_5976,N_5732);
xor U6829 (N_6829,N_5661,N_5238);
and U6830 (N_6830,N_5203,N_5878);
nand U6831 (N_6831,N_5339,N_5903);
nand U6832 (N_6832,N_5638,N_5878);
xor U6833 (N_6833,N_5592,N_5063);
nor U6834 (N_6834,N_5813,N_5243);
xor U6835 (N_6835,N_5082,N_5994);
nand U6836 (N_6836,N_5263,N_5857);
and U6837 (N_6837,N_5672,N_5903);
nand U6838 (N_6838,N_5025,N_5173);
nand U6839 (N_6839,N_5833,N_5801);
nand U6840 (N_6840,N_5630,N_5634);
and U6841 (N_6841,N_5435,N_5995);
nor U6842 (N_6842,N_5496,N_5793);
and U6843 (N_6843,N_5772,N_5510);
nor U6844 (N_6844,N_5384,N_5998);
or U6845 (N_6845,N_5887,N_5151);
and U6846 (N_6846,N_5058,N_5231);
nor U6847 (N_6847,N_5749,N_5441);
nand U6848 (N_6848,N_5362,N_5731);
or U6849 (N_6849,N_5185,N_5089);
nand U6850 (N_6850,N_5617,N_5499);
or U6851 (N_6851,N_5854,N_5268);
xor U6852 (N_6852,N_5853,N_5352);
and U6853 (N_6853,N_5800,N_5311);
or U6854 (N_6854,N_5803,N_5565);
xnor U6855 (N_6855,N_5742,N_5461);
nand U6856 (N_6856,N_5048,N_5186);
xor U6857 (N_6857,N_5453,N_5270);
xor U6858 (N_6858,N_5217,N_5885);
nand U6859 (N_6859,N_5577,N_5303);
xor U6860 (N_6860,N_5288,N_5014);
and U6861 (N_6861,N_5169,N_5363);
and U6862 (N_6862,N_5029,N_5730);
and U6863 (N_6863,N_5635,N_5434);
or U6864 (N_6864,N_5541,N_5577);
or U6865 (N_6865,N_5572,N_5204);
or U6866 (N_6866,N_5135,N_5658);
xnor U6867 (N_6867,N_5820,N_5227);
or U6868 (N_6868,N_5698,N_5545);
nand U6869 (N_6869,N_5344,N_5452);
and U6870 (N_6870,N_5585,N_5257);
and U6871 (N_6871,N_5871,N_5005);
and U6872 (N_6872,N_5424,N_5817);
or U6873 (N_6873,N_5234,N_5260);
or U6874 (N_6874,N_5957,N_5775);
xnor U6875 (N_6875,N_5133,N_5872);
nor U6876 (N_6876,N_5630,N_5363);
or U6877 (N_6877,N_5046,N_5937);
nor U6878 (N_6878,N_5410,N_5184);
and U6879 (N_6879,N_5772,N_5829);
nor U6880 (N_6880,N_5109,N_5512);
nand U6881 (N_6881,N_5085,N_5963);
nor U6882 (N_6882,N_5467,N_5623);
nand U6883 (N_6883,N_5018,N_5521);
or U6884 (N_6884,N_5262,N_5670);
nand U6885 (N_6885,N_5517,N_5744);
nor U6886 (N_6886,N_5754,N_5695);
nor U6887 (N_6887,N_5814,N_5613);
nand U6888 (N_6888,N_5963,N_5058);
xnor U6889 (N_6889,N_5125,N_5579);
or U6890 (N_6890,N_5918,N_5250);
nand U6891 (N_6891,N_5728,N_5036);
or U6892 (N_6892,N_5121,N_5411);
nand U6893 (N_6893,N_5139,N_5091);
nand U6894 (N_6894,N_5428,N_5845);
and U6895 (N_6895,N_5296,N_5057);
and U6896 (N_6896,N_5385,N_5890);
or U6897 (N_6897,N_5219,N_5295);
xnor U6898 (N_6898,N_5233,N_5528);
and U6899 (N_6899,N_5897,N_5728);
or U6900 (N_6900,N_5562,N_5445);
xor U6901 (N_6901,N_5614,N_5965);
nand U6902 (N_6902,N_5835,N_5752);
and U6903 (N_6903,N_5878,N_5057);
nand U6904 (N_6904,N_5458,N_5385);
or U6905 (N_6905,N_5513,N_5050);
nor U6906 (N_6906,N_5026,N_5152);
nor U6907 (N_6907,N_5258,N_5611);
and U6908 (N_6908,N_5008,N_5918);
nand U6909 (N_6909,N_5931,N_5892);
or U6910 (N_6910,N_5338,N_5748);
xor U6911 (N_6911,N_5094,N_5688);
xnor U6912 (N_6912,N_5453,N_5456);
nor U6913 (N_6913,N_5596,N_5513);
and U6914 (N_6914,N_5953,N_5066);
or U6915 (N_6915,N_5613,N_5418);
nand U6916 (N_6916,N_5822,N_5633);
nor U6917 (N_6917,N_5566,N_5498);
xor U6918 (N_6918,N_5697,N_5241);
or U6919 (N_6919,N_5106,N_5947);
xor U6920 (N_6920,N_5077,N_5552);
xor U6921 (N_6921,N_5913,N_5694);
nor U6922 (N_6922,N_5570,N_5390);
nor U6923 (N_6923,N_5730,N_5819);
nand U6924 (N_6924,N_5152,N_5188);
and U6925 (N_6925,N_5155,N_5890);
xnor U6926 (N_6926,N_5835,N_5914);
nor U6927 (N_6927,N_5304,N_5982);
or U6928 (N_6928,N_5192,N_5495);
or U6929 (N_6929,N_5761,N_5333);
nand U6930 (N_6930,N_5286,N_5727);
nor U6931 (N_6931,N_5955,N_5661);
xor U6932 (N_6932,N_5075,N_5660);
xor U6933 (N_6933,N_5245,N_5417);
and U6934 (N_6934,N_5199,N_5383);
or U6935 (N_6935,N_5880,N_5075);
and U6936 (N_6936,N_5115,N_5759);
or U6937 (N_6937,N_5388,N_5261);
nand U6938 (N_6938,N_5147,N_5037);
xnor U6939 (N_6939,N_5552,N_5692);
nand U6940 (N_6940,N_5956,N_5197);
nor U6941 (N_6941,N_5550,N_5388);
and U6942 (N_6942,N_5172,N_5979);
xnor U6943 (N_6943,N_5381,N_5333);
or U6944 (N_6944,N_5807,N_5719);
and U6945 (N_6945,N_5981,N_5125);
or U6946 (N_6946,N_5446,N_5569);
nand U6947 (N_6947,N_5804,N_5819);
xnor U6948 (N_6948,N_5587,N_5702);
xor U6949 (N_6949,N_5751,N_5647);
and U6950 (N_6950,N_5965,N_5270);
nor U6951 (N_6951,N_5225,N_5484);
nor U6952 (N_6952,N_5693,N_5585);
nand U6953 (N_6953,N_5955,N_5541);
nand U6954 (N_6954,N_5955,N_5799);
and U6955 (N_6955,N_5952,N_5815);
or U6956 (N_6956,N_5424,N_5490);
nor U6957 (N_6957,N_5059,N_5419);
nand U6958 (N_6958,N_5201,N_5130);
xnor U6959 (N_6959,N_5064,N_5389);
or U6960 (N_6960,N_5926,N_5181);
and U6961 (N_6961,N_5774,N_5702);
xnor U6962 (N_6962,N_5405,N_5586);
and U6963 (N_6963,N_5072,N_5324);
nand U6964 (N_6964,N_5784,N_5734);
xnor U6965 (N_6965,N_5941,N_5619);
nor U6966 (N_6966,N_5639,N_5112);
and U6967 (N_6967,N_5546,N_5117);
nand U6968 (N_6968,N_5233,N_5984);
or U6969 (N_6969,N_5104,N_5901);
and U6970 (N_6970,N_5203,N_5808);
xor U6971 (N_6971,N_5871,N_5769);
nand U6972 (N_6972,N_5679,N_5366);
nor U6973 (N_6973,N_5689,N_5992);
or U6974 (N_6974,N_5834,N_5831);
xor U6975 (N_6975,N_5401,N_5052);
nor U6976 (N_6976,N_5855,N_5342);
or U6977 (N_6977,N_5062,N_5511);
and U6978 (N_6978,N_5363,N_5096);
nand U6979 (N_6979,N_5686,N_5819);
nand U6980 (N_6980,N_5761,N_5884);
or U6981 (N_6981,N_5889,N_5597);
nor U6982 (N_6982,N_5344,N_5231);
and U6983 (N_6983,N_5168,N_5570);
nand U6984 (N_6984,N_5423,N_5510);
xnor U6985 (N_6985,N_5685,N_5621);
nor U6986 (N_6986,N_5398,N_5253);
and U6987 (N_6987,N_5489,N_5097);
xor U6988 (N_6988,N_5778,N_5784);
nor U6989 (N_6989,N_5115,N_5134);
nand U6990 (N_6990,N_5550,N_5419);
xor U6991 (N_6991,N_5820,N_5006);
and U6992 (N_6992,N_5015,N_5338);
or U6993 (N_6993,N_5248,N_5367);
and U6994 (N_6994,N_5458,N_5941);
nor U6995 (N_6995,N_5903,N_5831);
nor U6996 (N_6996,N_5728,N_5854);
nand U6997 (N_6997,N_5182,N_5381);
and U6998 (N_6998,N_5544,N_5949);
or U6999 (N_6999,N_5497,N_5618);
nand U7000 (N_7000,N_6195,N_6743);
nand U7001 (N_7001,N_6486,N_6671);
or U7002 (N_7002,N_6439,N_6634);
and U7003 (N_7003,N_6932,N_6350);
xnor U7004 (N_7004,N_6167,N_6248);
nand U7005 (N_7005,N_6741,N_6191);
or U7006 (N_7006,N_6044,N_6641);
xnor U7007 (N_7007,N_6446,N_6319);
and U7008 (N_7008,N_6669,N_6731);
and U7009 (N_7009,N_6636,N_6421);
or U7010 (N_7010,N_6948,N_6818);
nor U7011 (N_7011,N_6656,N_6036);
or U7012 (N_7012,N_6012,N_6241);
and U7013 (N_7013,N_6691,N_6535);
nor U7014 (N_7014,N_6298,N_6884);
nor U7015 (N_7015,N_6740,N_6040);
nor U7016 (N_7016,N_6806,N_6702);
nand U7017 (N_7017,N_6349,N_6847);
and U7018 (N_7018,N_6147,N_6686);
xor U7019 (N_7019,N_6412,N_6005);
nor U7020 (N_7020,N_6114,N_6067);
and U7021 (N_7021,N_6417,N_6336);
and U7022 (N_7022,N_6986,N_6247);
and U7023 (N_7023,N_6840,N_6532);
or U7024 (N_7024,N_6978,N_6983);
xor U7025 (N_7025,N_6124,N_6815);
and U7026 (N_7026,N_6888,N_6768);
xor U7027 (N_7027,N_6259,N_6724);
nand U7028 (N_7028,N_6726,N_6299);
nand U7029 (N_7029,N_6400,N_6221);
nor U7030 (N_7030,N_6531,N_6592);
or U7031 (N_7031,N_6562,N_6771);
or U7032 (N_7032,N_6396,N_6182);
and U7033 (N_7033,N_6008,N_6950);
nor U7034 (N_7034,N_6503,N_6628);
xnor U7035 (N_7035,N_6921,N_6719);
nor U7036 (N_7036,N_6386,N_6540);
and U7037 (N_7037,N_6677,N_6618);
nor U7038 (N_7038,N_6523,N_6845);
xnor U7039 (N_7039,N_6727,N_6559);
or U7040 (N_7040,N_6693,N_6514);
nand U7041 (N_7041,N_6829,N_6240);
and U7042 (N_7042,N_6415,N_6896);
xor U7043 (N_7043,N_6870,N_6251);
and U7044 (N_7044,N_6632,N_6046);
xor U7045 (N_7045,N_6141,N_6228);
or U7046 (N_7046,N_6521,N_6395);
or U7047 (N_7047,N_6613,N_6546);
xnor U7048 (N_7048,N_6650,N_6112);
or U7049 (N_7049,N_6738,N_6916);
nor U7050 (N_7050,N_6068,N_6313);
nand U7051 (N_7051,N_6157,N_6770);
nor U7052 (N_7052,N_6858,N_6301);
or U7053 (N_7053,N_6679,N_6994);
nor U7054 (N_7054,N_6057,N_6934);
or U7055 (N_7055,N_6452,N_6123);
nor U7056 (N_7056,N_6831,N_6069);
and U7057 (N_7057,N_6583,N_6661);
xnor U7058 (N_7058,N_6164,N_6939);
nor U7059 (N_7059,N_6537,N_6051);
xnor U7060 (N_7060,N_6672,N_6370);
nor U7061 (N_7061,N_6220,N_6111);
or U7062 (N_7062,N_6070,N_6625);
or U7063 (N_7063,N_6754,N_6784);
xnor U7064 (N_7064,N_6472,N_6424);
or U7065 (N_7065,N_6683,N_6128);
or U7066 (N_7066,N_6718,N_6365);
and U7067 (N_7067,N_6042,N_6804);
and U7068 (N_7068,N_6122,N_6226);
xor U7069 (N_7069,N_6675,N_6881);
nor U7070 (N_7070,N_6876,N_6029);
nor U7071 (N_7071,N_6183,N_6515);
nand U7072 (N_7072,N_6021,N_6561);
xor U7073 (N_7073,N_6843,N_6031);
nor U7074 (N_7074,N_6458,N_6149);
nand U7075 (N_7075,N_6734,N_6019);
or U7076 (N_7076,N_6755,N_6603);
nand U7077 (N_7077,N_6293,N_6316);
or U7078 (N_7078,N_6893,N_6127);
nand U7079 (N_7079,N_6476,N_6886);
nand U7080 (N_7080,N_6109,N_6974);
xor U7081 (N_7081,N_6020,N_6468);
and U7082 (N_7082,N_6721,N_6587);
and U7083 (N_7083,N_6168,N_6223);
xor U7084 (N_7084,N_6832,N_6200);
or U7085 (N_7085,N_6591,N_6491);
xnor U7086 (N_7086,N_6817,N_6694);
nand U7087 (N_7087,N_6972,N_6204);
nor U7088 (N_7088,N_6507,N_6563);
and U7089 (N_7089,N_6134,N_6139);
and U7090 (N_7090,N_6579,N_6857);
xnor U7091 (N_7091,N_6254,N_6580);
xnor U7092 (N_7092,N_6805,N_6558);
or U7093 (N_7093,N_6457,N_6766);
nand U7094 (N_7094,N_6135,N_6272);
xnor U7095 (N_7095,N_6668,N_6552);
or U7096 (N_7096,N_6748,N_6374);
nor U7097 (N_7097,N_6436,N_6667);
nor U7098 (N_7098,N_6793,N_6607);
nor U7099 (N_7099,N_6504,N_6955);
nor U7100 (N_7100,N_6369,N_6826);
xor U7101 (N_7101,N_6553,N_6985);
nand U7102 (N_7102,N_6414,N_6665);
xnor U7103 (N_7103,N_6957,N_6953);
and U7104 (N_7104,N_6496,N_6991);
and U7105 (N_7105,N_6216,N_6614);
xnor U7106 (N_7106,N_6066,N_6398);
nor U7107 (N_7107,N_6889,N_6851);
or U7108 (N_7108,N_6930,N_6894);
or U7109 (N_7109,N_6163,N_6624);
nor U7110 (N_7110,N_6153,N_6078);
and U7111 (N_7111,N_6494,N_6742);
or U7112 (N_7112,N_6030,N_6918);
or U7113 (N_7113,N_6002,N_6119);
nand U7114 (N_7114,N_6391,N_6217);
or U7115 (N_7115,N_6383,N_6509);
and U7116 (N_7116,N_6411,N_6685);
xnor U7117 (N_7117,N_6185,N_6321);
nor U7118 (N_7118,N_6730,N_6423);
and U7119 (N_7119,N_6354,N_6534);
xor U7120 (N_7120,N_6666,N_6642);
nand U7121 (N_7121,N_6648,N_6483);
nand U7122 (N_7122,N_6441,N_6337);
xor U7123 (N_7123,N_6343,N_6943);
nand U7124 (N_7124,N_6035,N_6853);
nor U7125 (N_7125,N_6173,N_6381);
nand U7126 (N_7126,N_6500,N_6309);
xnor U7127 (N_7127,N_6287,N_6631);
nor U7128 (N_7128,N_6184,N_6705);
nor U7129 (N_7129,N_6203,N_6404);
and U7130 (N_7130,N_6692,N_6456);
or U7131 (N_7131,N_6490,N_6033);
and U7132 (N_7132,N_6987,N_6497);
or U7133 (N_7133,N_6297,N_6659);
nor U7134 (N_7134,N_6998,N_6087);
and U7135 (N_7135,N_6879,N_6915);
nand U7136 (N_7136,N_6023,N_6593);
nor U7137 (N_7137,N_6001,N_6289);
and U7138 (N_7138,N_6442,N_6338);
xor U7139 (N_7139,N_6760,N_6110);
and U7140 (N_7140,N_6901,N_6554);
or U7141 (N_7141,N_6202,N_6467);
nor U7142 (N_7142,N_6864,N_6113);
nand U7143 (N_7143,N_6126,N_6431);
xnor U7144 (N_7144,N_6158,N_6096);
nand U7145 (N_7145,N_6043,N_6557);
xor U7146 (N_7146,N_6571,N_6024);
and U7147 (N_7147,N_6660,N_6092);
and U7148 (N_7148,N_6544,N_6419);
xor U7149 (N_7149,N_6574,N_6695);
nand U7150 (N_7150,N_6795,N_6697);
nor U7151 (N_7151,N_6746,N_6358);
nor U7152 (N_7152,N_6469,N_6739);
or U7153 (N_7153,N_6339,N_6984);
nor U7154 (N_7154,N_6891,N_6282);
nand U7155 (N_7155,N_6786,N_6264);
nor U7156 (N_7156,N_6682,N_6639);
xor U7157 (N_7157,N_6708,N_6175);
nand U7158 (N_7158,N_6551,N_6645);
nor U7159 (N_7159,N_6942,N_6244);
xor U7160 (N_7160,N_6867,N_6004);
xnor U7161 (N_7161,N_6288,N_6209);
and U7162 (N_7162,N_6849,N_6599);
nor U7163 (N_7163,N_6931,N_6397);
nor U7164 (N_7164,N_6969,N_6790);
nor U7165 (N_7165,N_6522,N_6283);
nor U7166 (N_7166,N_6025,N_6059);
nand U7167 (N_7167,N_6261,N_6905);
xor U7168 (N_7168,N_6410,N_6154);
nor U7169 (N_7169,N_6996,N_6951);
and U7170 (N_7170,N_6302,N_6049);
nand U7171 (N_7171,N_6756,N_6892);
xor U7172 (N_7172,N_6187,N_6802);
nor U7173 (N_7173,N_6954,N_6758);
nor U7174 (N_7174,N_6463,N_6373);
nor U7175 (N_7175,N_6461,N_6041);
nand U7176 (N_7176,N_6435,N_6052);
nand U7177 (N_7177,N_6792,N_6062);
xor U7178 (N_7178,N_6108,N_6919);
or U7179 (N_7179,N_6159,N_6909);
nor U7180 (N_7180,N_6594,N_6451);
nand U7181 (N_7181,N_6081,N_6376);
xor U7182 (N_7182,N_6478,N_6578);
and U7183 (N_7183,N_6524,N_6810);
xnor U7184 (N_7184,N_6920,N_6017);
or U7185 (N_7185,N_6085,N_6866);
or U7186 (N_7186,N_6207,N_6459);
and U7187 (N_7187,N_6883,N_6151);
nor U7188 (N_7188,N_6312,N_6824);
nor U7189 (N_7189,N_6575,N_6097);
xor U7190 (N_7190,N_6638,N_6455);
xnor U7191 (N_7191,N_6873,N_6773);
nor U7192 (N_7192,N_6246,N_6305);
and U7193 (N_7193,N_6772,N_6935);
nor U7194 (N_7194,N_6627,N_6406);
nor U7195 (N_7195,N_6308,N_6077);
nor U7196 (N_7196,N_6902,N_6505);
and U7197 (N_7197,N_6785,N_6809);
nand U7198 (N_7198,N_6517,N_6556);
nor U7199 (N_7199,N_6712,N_6479);
or U7200 (N_7200,N_6555,N_6545);
nand U7201 (N_7201,N_6156,N_6854);
and U7202 (N_7202,N_6484,N_6060);
and U7203 (N_7203,N_6944,N_6566);
or U7204 (N_7204,N_6131,N_6965);
or U7205 (N_7205,N_6968,N_6116);
nand U7206 (N_7206,N_6776,N_6949);
nor U7207 (N_7207,N_6630,N_6732);
or U7208 (N_7208,N_6995,N_6527);
nand U7209 (N_7209,N_6003,N_6573);
nand U7210 (N_7210,N_6160,N_6009);
nand U7211 (N_7211,N_6977,N_6703);
and U7212 (N_7212,N_6433,N_6728);
xnor U7213 (N_7213,N_6617,N_6878);
nor U7214 (N_7214,N_6783,N_6382);
or U7215 (N_7215,N_6198,N_6488);
xor U7216 (N_7216,N_6234,N_6595);
or U7217 (N_7217,N_6268,N_6895);
nor U7218 (N_7218,N_6304,N_6233);
nor U7219 (N_7219,N_6992,N_6814);
and U7220 (N_7220,N_6064,N_6150);
nor U7221 (N_7221,N_6447,N_6063);
xor U7222 (N_7222,N_6684,N_6178);
or U7223 (N_7223,N_6820,N_6605);
and U7224 (N_7224,N_6260,N_6711);
nor U7225 (N_7225,N_6794,N_6481);
nor U7226 (N_7226,N_6637,N_6306);
and U7227 (N_7227,N_6769,N_6189);
nor U7228 (N_7228,N_6989,N_6144);
nand U7229 (N_7229,N_6101,N_6148);
or U7230 (N_7230,N_6401,N_6560);
or U7231 (N_7231,N_6947,N_6493);
nand U7232 (N_7232,N_6443,N_6548);
nand U7233 (N_7233,N_6192,N_6292);
and U7234 (N_7234,N_6520,N_6420);
nand U7235 (N_7235,N_6232,N_6162);
nand U7236 (N_7236,N_6880,N_6936);
xnor U7237 (N_7237,N_6577,N_6499);
nand U7238 (N_7238,N_6710,N_6698);
xor U7239 (N_7239,N_6225,N_6913);
nor U7240 (N_7240,N_6361,N_6762);
or U7241 (N_7241,N_6345,N_6926);
nand U7242 (N_7242,N_6798,N_6117);
or U7243 (N_7243,N_6425,N_6837);
xnor U7244 (N_7244,N_6655,N_6775);
nor U7245 (N_7245,N_6541,N_6498);
xnor U7246 (N_7246,N_6564,N_6196);
nand U7247 (N_7247,N_6501,N_6871);
xor U7248 (N_7248,N_6725,N_6797);
nor U7249 (N_7249,N_6016,N_6598);
nand U7250 (N_7250,N_6485,N_6372);
and U7251 (N_7251,N_6588,N_6224);
or U7252 (N_7252,N_6568,N_6807);
xnor U7253 (N_7253,N_6589,N_6388);
or U7254 (N_7254,N_6611,N_6080);
or U7255 (N_7255,N_6946,N_6174);
or U7256 (N_7256,N_6529,N_6856);
and U7257 (N_7257,N_6502,N_6342);
nor U7258 (N_7258,N_6327,N_6166);
nand U7259 (N_7259,N_6427,N_6600);
or U7260 (N_7260,N_6767,N_6800);
nand U7261 (N_7261,N_6214,N_6480);
nor U7262 (N_7262,N_6887,N_6231);
xnor U7263 (N_7263,N_6704,N_6328);
nand U7264 (N_7264,N_6229,N_6606);
or U7265 (N_7265,N_6190,N_6914);
nor U7266 (N_7266,N_6547,N_6238);
nor U7267 (N_7267,N_6280,N_6872);
and U7268 (N_7268,N_6542,N_6054);
xor U7269 (N_7269,N_6177,N_6674);
and U7270 (N_7270,N_6621,N_6543);
xor U7271 (N_7271,N_6859,N_6812);
nand U7272 (N_7272,N_6927,N_6171);
and U7273 (N_7273,N_6910,N_6917);
or U7274 (N_7274,N_6565,N_6394);
or U7275 (N_7275,N_6375,N_6314);
nand U7276 (N_7276,N_6699,N_6828);
xnor U7277 (N_7277,N_6324,N_6295);
or U7278 (N_7278,N_6133,N_6359);
nor U7279 (N_7279,N_6093,N_6610);
nand U7280 (N_7280,N_6351,N_6700);
nor U7281 (N_7281,N_6982,N_6519);
nand U7282 (N_7282,N_6550,N_6549);
and U7283 (N_7283,N_6102,N_6687);
nand U7284 (N_7284,N_6048,N_6356);
nor U7285 (N_7285,N_6958,N_6201);
xor U7286 (N_7286,N_6975,N_6011);
and U7287 (N_7287,N_6367,N_6651);
nand U7288 (N_7288,N_6530,N_6208);
nor U7289 (N_7289,N_6952,N_6979);
nand U7290 (N_7290,N_6130,N_6010);
nand U7291 (N_7291,N_6205,N_6027);
and U7292 (N_7292,N_6334,N_6170);
nor U7293 (N_7293,N_6852,N_6609);
xor U7294 (N_7294,N_6363,N_6875);
nand U7295 (N_7295,N_6765,N_6999);
nand U7296 (N_7296,N_6058,N_6475);
and U7297 (N_7297,N_6325,N_6352);
or U7298 (N_7298,N_6581,N_6779);
xor U7299 (N_7299,N_6990,N_6567);
nand U7300 (N_7300,N_6258,N_6335);
nand U7301 (N_7301,N_6877,N_6569);
xnor U7302 (N_7302,N_6644,N_6848);
xor U7303 (N_7303,N_6715,N_6657);
and U7304 (N_7304,N_6923,N_6836);
or U7305 (N_7305,N_6409,N_6083);
nor U7306 (N_7306,N_6941,N_6125);
nor U7307 (N_7307,N_6846,N_6448);
or U7308 (N_7308,N_6347,N_6688);
nor U7309 (N_7309,N_6937,N_6819);
nand U7310 (N_7310,N_6658,N_6047);
nand U7311 (N_7311,N_6281,N_6825);
and U7312 (N_7312,N_6830,N_6462);
nand U7313 (N_7313,N_6318,N_6713);
xnor U7314 (N_7314,N_6906,N_6744);
xnor U7315 (N_7315,N_6082,N_6371);
nor U7316 (N_7316,N_6407,N_6752);
or U7317 (N_7317,N_6393,N_6422);
nand U7318 (N_7318,N_6640,N_6464);
and U7319 (N_7319,N_6761,N_6115);
nor U7320 (N_7320,N_6215,N_6267);
or U7321 (N_7321,N_6445,N_6716);
xnor U7322 (N_7322,N_6249,N_6473);
xnor U7323 (N_7323,N_6105,N_6291);
or U7324 (N_7324,N_6834,N_6899);
nor U7325 (N_7325,N_6053,N_6253);
nor U7326 (N_7326,N_6094,N_6323);
xnor U7327 (N_7327,N_6993,N_6787);
or U7328 (N_7328,N_6311,N_6188);
or U7329 (N_7329,N_6516,N_6907);
xor U7330 (N_7330,N_6865,N_6492);
nor U7331 (N_7331,N_6495,N_6180);
nor U7332 (N_7332,N_6643,N_6956);
and U7333 (N_7333,N_6850,N_6256);
or U7334 (N_7334,N_6266,N_6444);
or U7335 (N_7335,N_6277,N_6320);
nor U7336 (N_7336,N_6526,N_6827);
xor U7337 (N_7337,N_6142,N_6405);
xnor U7338 (N_7338,N_6106,N_6000);
and U7339 (N_7339,N_6402,N_6315);
nor U7340 (N_7340,N_6416,N_6964);
or U7341 (N_7341,N_6353,N_6013);
xnor U7342 (N_7342,N_6757,N_6924);
nor U7343 (N_7343,N_6511,N_6132);
and U7344 (N_7344,N_6034,N_6026);
xor U7345 (N_7345,N_6822,N_6525);
nor U7346 (N_7346,N_6165,N_6874);
or U7347 (N_7347,N_6399,N_6265);
or U7348 (N_7348,N_6426,N_6152);
xnor U7349 (N_7349,N_6222,N_6844);
or U7350 (N_7350,N_6155,N_6169);
nor U7351 (N_7351,N_6273,N_6676);
nor U7352 (N_7352,N_6211,N_6100);
nor U7353 (N_7353,N_6582,N_6300);
and U7354 (N_7354,N_6392,N_6032);
or U7355 (N_7355,N_6720,N_6533);
xnor U7356 (N_7356,N_6791,N_6868);
or U7357 (N_7357,N_6833,N_6018);
nor U7358 (N_7358,N_6487,N_6938);
xnor U7359 (N_7359,N_6821,N_6257);
xnor U7360 (N_7360,N_6237,N_6673);
xor U7361 (N_7361,N_6090,N_6489);
and U7362 (N_7362,N_6570,N_6103);
nor U7363 (N_7363,N_6799,N_6903);
nor U7364 (N_7364,N_6737,N_6193);
or U7365 (N_7365,N_6513,N_6310);
nor U7366 (N_7366,N_6709,N_6245);
nand U7367 (N_7367,N_6186,N_6270);
or U7368 (N_7368,N_6616,N_6678);
nor U7369 (N_7369,N_6908,N_6075);
or U7370 (N_7370,N_6007,N_6121);
xor U7371 (N_7371,N_6839,N_6646);
nor U7372 (N_7372,N_6197,N_6729);
nor U7373 (N_7373,N_6140,N_6777);
nand U7374 (N_7374,N_6065,N_6970);
or U7375 (N_7375,N_6466,N_6681);
nand U7376 (N_7376,N_6317,N_6782);
nor U7377 (N_7377,N_6344,N_6107);
and U7378 (N_7378,N_6680,N_6922);
and U7379 (N_7379,N_6963,N_6835);
xor U7380 (N_7380,N_6945,N_6199);
or U7381 (N_7381,N_6285,N_6988);
nand U7382 (N_7382,N_6763,N_6961);
nor U7383 (N_7383,N_6104,N_6294);
nand U7384 (N_7384,N_6898,N_6663);
xnor U7385 (N_7385,N_6296,N_6389);
nand U7386 (N_7386,N_6213,N_6745);
and U7387 (N_7387,N_6252,N_6633);
and U7388 (N_7388,N_6378,N_6454);
xor U7389 (N_7389,N_6022,N_6808);
and U7390 (N_7390,N_6028,N_6366);
or U7391 (N_7391,N_6512,N_6084);
xor U7392 (N_7392,N_6778,N_6967);
or U7393 (N_7393,N_6604,N_6911);
nand U7394 (N_7394,N_6622,N_6477);
or U7395 (N_7395,N_6377,N_6747);
nand U7396 (N_7396,N_6368,N_6037);
or U7397 (N_7397,N_6664,N_6418);
nand U7398 (N_7398,N_6780,N_6360);
nor U7399 (N_7399,N_6750,N_6855);
xnor U7400 (N_7400,N_6331,N_6962);
nand U7401 (N_7401,N_6278,N_6143);
xor U7402 (N_7402,N_6863,N_6789);
and U7403 (N_7403,N_6933,N_6882);
and U7404 (N_7404,N_6006,N_6434);
nand U7405 (N_7405,N_6437,N_6652);
or U7406 (N_7406,N_6269,N_6654);
nand U7407 (N_7407,N_6061,N_6074);
xnor U7408 (N_7408,N_6218,N_6960);
nor U7409 (N_7409,N_6286,N_6242);
xor U7410 (N_7410,N_6120,N_6227);
nor U7411 (N_7411,N_6073,N_6980);
nand U7412 (N_7412,N_6429,N_6813);
and U7413 (N_7413,N_6584,N_6751);
nor U7414 (N_7414,N_6385,N_6136);
nand U7415 (N_7415,N_6925,N_6689);
nor U7416 (N_7416,N_6384,N_6438);
and U7417 (N_7417,N_6091,N_6212);
xnor U7418 (N_7418,N_6619,N_6355);
or U7419 (N_7419,N_6340,N_6981);
xor U7420 (N_7420,N_6528,N_6210);
nor U7421 (N_7421,N_6390,N_6088);
nand U7422 (N_7422,N_6236,N_6346);
nand U7423 (N_7423,N_6647,N_6239);
xnor U7424 (N_7424,N_6250,N_6602);
or U7425 (N_7425,N_6403,N_6973);
nor U7426 (N_7426,N_6076,N_6735);
or U7427 (N_7427,N_6255,N_6460);
and U7428 (N_7428,N_6940,N_6620);
nor U7429 (N_7429,N_6841,N_6307);
or U7430 (N_7430,N_6161,N_6089);
nand U7431 (N_7431,N_6172,N_6869);
nor U7432 (N_7432,N_6050,N_6271);
or U7433 (N_7433,N_6736,N_6722);
and U7434 (N_7434,N_6072,N_6518);
and U7435 (N_7435,N_6508,N_6408);
xor U7436 (N_7436,N_6904,N_6219);
or U7437 (N_7437,N_6179,N_6099);
and U7438 (N_7438,N_6230,N_6332);
or U7439 (N_7439,N_6538,N_6243);
or U7440 (N_7440,N_6056,N_6430);
nor U7441 (N_7441,N_6601,N_6900);
nor U7442 (N_7442,N_6626,N_6181);
xnor U7443 (N_7443,N_6539,N_6861);
nor U7444 (N_7444,N_6753,N_6788);
or U7445 (N_7445,N_6118,N_6774);
nor U7446 (N_7446,N_6585,N_6290);
and U7447 (N_7447,N_6597,N_6303);
or U7448 (N_7448,N_6206,N_6428);
nor U7449 (N_7449,N_6629,N_6959);
nand U7450 (N_7450,N_6928,N_6357);
xnor U7451 (N_7451,N_6701,N_6796);
and U7452 (N_7452,N_6362,N_6816);
xor U7453 (N_7453,N_6379,N_6038);
and U7454 (N_7454,N_6971,N_6842);
and U7455 (N_7455,N_6333,N_6707);
and U7456 (N_7456,N_6482,N_6838);
and U7457 (N_7457,N_6860,N_6138);
nor U7458 (N_7458,N_6055,N_6862);
or U7459 (N_7459,N_6284,N_6714);
nor U7460 (N_7460,N_6039,N_6470);
and U7461 (N_7461,N_6471,N_6706);
or U7462 (N_7462,N_6576,N_6275);
nand U7463 (N_7463,N_6976,N_6764);
nand U7464 (N_7464,N_6326,N_6885);
nor U7465 (N_7465,N_6440,N_6098);
nand U7466 (N_7466,N_6586,N_6723);
nor U7467 (N_7467,N_6095,N_6274);
nand U7468 (N_7468,N_6387,N_6510);
xnor U7469 (N_7469,N_6014,N_6474);
nor U7470 (N_7470,N_6635,N_6596);
and U7471 (N_7471,N_6670,N_6966);
or U7472 (N_7472,N_6235,N_6145);
or U7473 (N_7473,N_6717,N_6453);
nand U7474 (N_7474,N_6653,N_6194);
or U7475 (N_7475,N_6506,N_6572);
and U7476 (N_7476,N_6781,N_6623);
nor U7477 (N_7477,N_6137,N_6465);
nand U7478 (N_7478,N_6086,N_6330);
or U7479 (N_7479,N_6329,N_6279);
nand U7480 (N_7480,N_6322,N_6432);
nand U7481 (N_7481,N_6612,N_6696);
xnor U7482 (N_7482,N_6749,N_6662);
nor U7483 (N_7483,N_6649,N_6997);
and U7484 (N_7484,N_6929,N_6733);
and U7485 (N_7485,N_6262,N_6912);
or U7486 (N_7486,N_6801,N_6079);
xor U7487 (N_7487,N_6176,N_6803);
xnor U7488 (N_7488,N_6897,N_6890);
xor U7489 (N_7489,N_6348,N_6536);
xor U7490 (N_7490,N_6263,N_6608);
and U7491 (N_7491,N_6146,N_6380);
nand U7492 (N_7492,N_6590,N_6811);
nor U7493 (N_7493,N_6045,N_6823);
xnor U7494 (N_7494,N_6615,N_6364);
nor U7495 (N_7495,N_6341,N_6071);
or U7496 (N_7496,N_6759,N_6413);
nor U7497 (N_7497,N_6129,N_6015);
xnor U7498 (N_7498,N_6450,N_6690);
nand U7499 (N_7499,N_6276,N_6449);
nor U7500 (N_7500,N_6592,N_6093);
nand U7501 (N_7501,N_6512,N_6785);
xnor U7502 (N_7502,N_6955,N_6176);
and U7503 (N_7503,N_6424,N_6071);
and U7504 (N_7504,N_6325,N_6821);
nor U7505 (N_7505,N_6589,N_6171);
nand U7506 (N_7506,N_6781,N_6476);
nor U7507 (N_7507,N_6762,N_6643);
nor U7508 (N_7508,N_6264,N_6363);
and U7509 (N_7509,N_6438,N_6038);
or U7510 (N_7510,N_6793,N_6737);
nand U7511 (N_7511,N_6221,N_6993);
xor U7512 (N_7512,N_6344,N_6608);
nor U7513 (N_7513,N_6721,N_6087);
or U7514 (N_7514,N_6504,N_6636);
xor U7515 (N_7515,N_6230,N_6284);
xnor U7516 (N_7516,N_6935,N_6462);
and U7517 (N_7517,N_6702,N_6756);
nor U7518 (N_7518,N_6284,N_6036);
xnor U7519 (N_7519,N_6914,N_6065);
and U7520 (N_7520,N_6406,N_6432);
nand U7521 (N_7521,N_6776,N_6483);
xor U7522 (N_7522,N_6003,N_6540);
and U7523 (N_7523,N_6629,N_6322);
xor U7524 (N_7524,N_6369,N_6164);
and U7525 (N_7525,N_6930,N_6233);
or U7526 (N_7526,N_6558,N_6277);
and U7527 (N_7527,N_6119,N_6139);
and U7528 (N_7528,N_6634,N_6498);
xnor U7529 (N_7529,N_6621,N_6820);
nor U7530 (N_7530,N_6226,N_6763);
nand U7531 (N_7531,N_6189,N_6220);
xnor U7532 (N_7532,N_6315,N_6931);
and U7533 (N_7533,N_6409,N_6718);
and U7534 (N_7534,N_6862,N_6132);
and U7535 (N_7535,N_6182,N_6814);
and U7536 (N_7536,N_6513,N_6126);
xnor U7537 (N_7537,N_6743,N_6820);
and U7538 (N_7538,N_6377,N_6429);
nand U7539 (N_7539,N_6450,N_6419);
nor U7540 (N_7540,N_6038,N_6468);
xnor U7541 (N_7541,N_6968,N_6329);
xnor U7542 (N_7542,N_6374,N_6024);
nor U7543 (N_7543,N_6234,N_6708);
xnor U7544 (N_7544,N_6456,N_6498);
and U7545 (N_7545,N_6261,N_6978);
nand U7546 (N_7546,N_6152,N_6429);
nor U7547 (N_7547,N_6044,N_6319);
nand U7548 (N_7548,N_6457,N_6054);
and U7549 (N_7549,N_6091,N_6689);
and U7550 (N_7550,N_6285,N_6410);
or U7551 (N_7551,N_6306,N_6264);
or U7552 (N_7552,N_6874,N_6923);
nor U7553 (N_7553,N_6028,N_6971);
nand U7554 (N_7554,N_6658,N_6867);
or U7555 (N_7555,N_6647,N_6849);
or U7556 (N_7556,N_6365,N_6134);
nor U7557 (N_7557,N_6284,N_6461);
and U7558 (N_7558,N_6309,N_6429);
xor U7559 (N_7559,N_6873,N_6200);
xor U7560 (N_7560,N_6266,N_6479);
xor U7561 (N_7561,N_6014,N_6491);
nor U7562 (N_7562,N_6518,N_6195);
nor U7563 (N_7563,N_6555,N_6095);
and U7564 (N_7564,N_6747,N_6693);
or U7565 (N_7565,N_6426,N_6988);
and U7566 (N_7566,N_6473,N_6813);
and U7567 (N_7567,N_6798,N_6766);
xor U7568 (N_7568,N_6723,N_6136);
and U7569 (N_7569,N_6358,N_6562);
nand U7570 (N_7570,N_6391,N_6633);
xnor U7571 (N_7571,N_6444,N_6148);
or U7572 (N_7572,N_6063,N_6292);
and U7573 (N_7573,N_6157,N_6656);
nor U7574 (N_7574,N_6839,N_6019);
nor U7575 (N_7575,N_6304,N_6697);
nand U7576 (N_7576,N_6124,N_6158);
and U7577 (N_7577,N_6768,N_6849);
xor U7578 (N_7578,N_6402,N_6733);
and U7579 (N_7579,N_6609,N_6330);
or U7580 (N_7580,N_6409,N_6211);
xnor U7581 (N_7581,N_6335,N_6984);
or U7582 (N_7582,N_6842,N_6083);
nand U7583 (N_7583,N_6297,N_6933);
or U7584 (N_7584,N_6296,N_6877);
or U7585 (N_7585,N_6735,N_6605);
nand U7586 (N_7586,N_6855,N_6473);
nor U7587 (N_7587,N_6478,N_6249);
and U7588 (N_7588,N_6275,N_6816);
xor U7589 (N_7589,N_6130,N_6524);
or U7590 (N_7590,N_6115,N_6033);
nand U7591 (N_7591,N_6565,N_6218);
xnor U7592 (N_7592,N_6935,N_6436);
or U7593 (N_7593,N_6002,N_6110);
nand U7594 (N_7594,N_6451,N_6453);
xnor U7595 (N_7595,N_6855,N_6557);
xnor U7596 (N_7596,N_6600,N_6132);
nor U7597 (N_7597,N_6985,N_6649);
nand U7598 (N_7598,N_6298,N_6593);
nand U7599 (N_7599,N_6927,N_6958);
nor U7600 (N_7600,N_6450,N_6624);
or U7601 (N_7601,N_6364,N_6645);
or U7602 (N_7602,N_6019,N_6821);
nor U7603 (N_7603,N_6807,N_6878);
nor U7604 (N_7604,N_6191,N_6455);
nand U7605 (N_7605,N_6684,N_6935);
nor U7606 (N_7606,N_6470,N_6549);
xor U7607 (N_7607,N_6349,N_6897);
xnor U7608 (N_7608,N_6986,N_6028);
nor U7609 (N_7609,N_6571,N_6349);
xnor U7610 (N_7610,N_6126,N_6919);
xor U7611 (N_7611,N_6054,N_6022);
or U7612 (N_7612,N_6152,N_6380);
xnor U7613 (N_7613,N_6687,N_6799);
nand U7614 (N_7614,N_6630,N_6588);
and U7615 (N_7615,N_6830,N_6102);
and U7616 (N_7616,N_6681,N_6316);
and U7617 (N_7617,N_6285,N_6247);
xnor U7618 (N_7618,N_6347,N_6007);
nor U7619 (N_7619,N_6902,N_6527);
nor U7620 (N_7620,N_6160,N_6050);
and U7621 (N_7621,N_6273,N_6554);
nor U7622 (N_7622,N_6394,N_6868);
nor U7623 (N_7623,N_6380,N_6636);
nand U7624 (N_7624,N_6404,N_6768);
nor U7625 (N_7625,N_6983,N_6387);
nand U7626 (N_7626,N_6551,N_6277);
nor U7627 (N_7627,N_6547,N_6435);
xor U7628 (N_7628,N_6490,N_6025);
nor U7629 (N_7629,N_6912,N_6944);
nand U7630 (N_7630,N_6838,N_6164);
nor U7631 (N_7631,N_6726,N_6957);
or U7632 (N_7632,N_6263,N_6709);
or U7633 (N_7633,N_6351,N_6431);
xnor U7634 (N_7634,N_6725,N_6359);
xor U7635 (N_7635,N_6389,N_6431);
nand U7636 (N_7636,N_6664,N_6304);
nand U7637 (N_7637,N_6650,N_6087);
nor U7638 (N_7638,N_6058,N_6052);
xnor U7639 (N_7639,N_6944,N_6471);
nor U7640 (N_7640,N_6194,N_6988);
xnor U7641 (N_7641,N_6436,N_6388);
and U7642 (N_7642,N_6909,N_6375);
nand U7643 (N_7643,N_6621,N_6849);
and U7644 (N_7644,N_6479,N_6587);
nand U7645 (N_7645,N_6287,N_6000);
nor U7646 (N_7646,N_6569,N_6109);
and U7647 (N_7647,N_6474,N_6566);
xnor U7648 (N_7648,N_6545,N_6319);
nand U7649 (N_7649,N_6091,N_6294);
nand U7650 (N_7650,N_6618,N_6190);
and U7651 (N_7651,N_6833,N_6291);
nand U7652 (N_7652,N_6055,N_6343);
xnor U7653 (N_7653,N_6625,N_6451);
nand U7654 (N_7654,N_6837,N_6475);
xor U7655 (N_7655,N_6227,N_6387);
or U7656 (N_7656,N_6825,N_6903);
nor U7657 (N_7657,N_6635,N_6033);
and U7658 (N_7658,N_6417,N_6107);
xnor U7659 (N_7659,N_6493,N_6916);
nand U7660 (N_7660,N_6612,N_6990);
and U7661 (N_7661,N_6330,N_6507);
and U7662 (N_7662,N_6517,N_6417);
nor U7663 (N_7663,N_6103,N_6793);
xnor U7664 (N_7664,N_6337,N_6479);
xor U7665 (N_7665,N_6046,N_6610);
nor U7666 (N_7666,N_6335,N_6951);
nor U7667 (N_7667,N_6339,N_6229);
xor U7668 (N_7668,N_6789,N_6929);
xnor U7669 (N_7669,N_6161,N_6534);
xor U7670 (N_7670,N_6106,N_6708);
and U7671 (N_7671,N_6925,N_6973);
nand U7672 (N_7672,N_6821,N_6674);
nor U7673 (N_7673,N_6171,N_6660);
xor U7674 (N_7674,N_6116,N_6396);
xnor U7675 (N_7675,N_6941,N_6234);
nor U7676 (N_7676,N_6676,N_6518);
xnor U7677 (N_7677,N_6061,N_6382);
xor U7678 (N_7678,N_6668,N_6703);
and U7679 (N_7679,N_6806,N_6569);
nor U7680 (N_7680,N_6831,N_6021);
xor U7681 (N_7681,N_6988,N_6461);
or U7682 (N_7682,N_6627,N_6323);
nand U7683 (N_7683,N_6257,N_6939);
and U7684 (N_7684,N_6653,N_6723);
xor U7685 (N_7685,N_6412,N_6056);
or U7686 (N_7686,N_6142,N_6971);
or U7687 (N_7687,N_6805,N_6839);
or U7688 (N_7688,N_6272,N_6176);
and U7689 (N_7689,N_6818,N_6636);
and U7690 (N_7690,N_6223,N_6509);
nand U7691 (N_7691,N_6774,N_6145);
and U7692 (N_7692,N_6606,N_6749);
nor U7693 (N_7693,N_6205,N_6056);
nand U7694 (N_7694,N_6060,N_6122);
nand U7695 (N_7695,N_6598,N_6817);
and U7696 (N_7696,N_6885,N_6123);
nor U7697 (N_7697,N_6966,N_6544);
nor U7698 (N_7698,N_6291,N_6228);
nand U7699 (N_7699,N_6388,N_6029);
nor U7700 (N_7700,N_6735,N_6983);
nand U7701 (N_7701,N_6018,N_6427);
nand U7702 (N_7702,N_6380,N_6287);
xor U7703 (N_7703,N_6990,N_6078);
nor U7704 (N_7704,N_6414,N_6784);
or U7705 (N_7705,N_6947,N_6399);
nor U7706 (N_7706,N_6592,N_6834);
xnor U7707 (N_7707,N_6676,N_6057);
and U7708 (N_7708,N_6376,N_6752);
and U7709 (N_7709,N_6373,N_6596);
xnor U7710 (N_7710,N_6577,N_6866);
and U7711 (N_7711,N_6593,N_6227);
nor U7712 (N_7712,N_6888,N_6245);
xor U7713 (N_7713,N_6804,N_6255);
xnor U7714 (N_7714,N_6558,N_6791);
or U7715 (N_7715,N_6757,N_6715);
nor U7716 (N_7716,N_6271,N_6827);
nor U7717 (N_7717,N_6435,N_6999);
xor U7718 (N_7718,N_6083,N_6241);
nand U7719 (N_7719,N_6278,N_6886);
nand U7720 (N_7720,N_6788,N_6859);
xor U7721 (N_7721,N_6501,N_6975);
nor U7722 (N_7722,N_6765,N_6254);
or U7723 (N_7723,N_6707,N_6125);
xor U7724 (N_7724,N_6088,N_6656);
xnor U7725 (N_7725,N_6821,N_6673);
nand U7726 (N_7726,N_6124,N_6168);
nor U7727 (N_7727,N_6122,N_6972);
nand U7728 (N_7728,N_6913,N_6884);
xnor U7729 (N_7729,N_6467,N_6949);
xnor U7730 (N_7730,N_6988,N_6128);
and U7731 (N_7731,N_6835,N_6078);
nand U7732 (N_7732,N_6062,N_6962);
and U7733 (N_7733,N_6976,N_6542);
or U7734 (N_7734,N_6865,N_6183);
nand U7735 (N_7735,N_6943,N_6314);
nand U7736 (N_7736,N_6481,N_6666);
nor U7737 (N_7737,N_6070,N_6280);
xnor U7738 (N_7738,N_6640,N_6702);
xnor U7739 (N_7739,N_6779,N_6815);
nand U7740 (N_7740,N_6515,N_6274);
and U7741 (N_7741,N_6734,N_6686);
nor U7742 (N_7742,N_6607,N_6058);
nand U7743 (N_7743,N_6287,N_6103);
or U7744 (N_7744,N_6076,N_6274);
nand U7745 (N_7745,N_6794,N_6787);
nand U7746 (N_7746,N_6368,N_6614);
and U7747 (N_7747,N_6076,N_6703);
nand U7748 (N_7748,N_6046,N_6974);
and U7749 (N_7749,N_6739,N_6209);
or U7750 (N_7750,N_6979,N_6088);
nor U7751 (N_7751,N_6441,N_6447);
nor U7752 (N_7752,N_6091,N_6996);
and U7753 (N_7753,N_6783,N_6141);
or U7754 (N_7754,N_6244,N_6054);
and U7755 (N_7755,N_6818,N_6444);
and U7756 (N_7756,N_6430,N_6424);
xnor U7757 (N_7757,N_6118,N_6519);
and U7758 (N_7758,N_6396,N_6194);
and U7759 (N_7759,N_6230,N_6082);
or U7760 (N_7760,N_6646,N_6508);
nor U7761 (N_7761,N_6058,N_6094);
and U7762 (N_7762,N_6671,N_6351);
nor U7763 (N_7763,N_6673,N_6885);
nor U7764 (N_7764,N_6096,N_6157);
xor U7765 (N_7765,N_6423,N_6307);
or U7766 (N_7766,N_6625,N_6346);
nor U7767 (N_7767,N_6099,N_6175);
nor U7768 (N_7768,N_6182,N_6129);
xor U7769 (N_7769,N_6028,N_6407);
nand U7770 (N_7770,N_6152,N_6615);
and U7771 (N_7771,N_6728,N_6565);
and U7772 (N_7772,N_6786,N_6841);
xnor U7773 (N_7773,N_6709,N_6319);
xnor U7774 (N_7774,N_6064,N_6352);
nor U7775 (N_7775,N_6082,N_6984);
xnor U7776 (N_7776,N_6988,N_6247);
xor U7777 (N_7777,N_6464,N_6724);
nor U7778 (N_7778,N_6596,N_6142);
and U7779 (N_7779,N_6727,N_6672);
or U7780 (N_7780,N_6107,N_6189);
nand U7781 (N_7781,N_6127,N_6095);
or U7782 (N_7782,N_6010,N_6883);
nor U7783 (N_7783,N_6114,N_6887);
and U7784 (N_7784,N_6975,N_6592);
xnor U7785 (N_7785,N_6348,N_6113);
xor U7786 (N_7786,N_6537,N_6980);
nand U7787 (N_7787,N_6492,N_6649);
nand U7788 (N_7788,N_6138,N_6524);
xnor U7789 (N_7789,N_6672,N_6837);
nand U7790 (N_7790,N_6296,N_6630);
or U7791 (N_7791,N_6033,N_6790);
or U7792 (N_7792,N_6914,N_6984);
and U7793 (N_7793,N_6213,N_6137);
nor U7794 (N_7794,N_6839,N_6017);
and U7795 (N_7795,N_6605,N_6448);
nand U7796 (N_7796,N_6783,N_6060);
or U7797 (N_7797,N_6968,N_6908);
or U7798 (N_7798,N_6413,N_6124);
and U7799 (N_7799,N_6101,N_6316);
nor U7800 (N_7800,N_6658,N_6251);
xnor U7801 (N_7801,N_6970,N_6771);
and U7802 (N_7802,N_6904,N_6746);
nor U7803 (N_7803,N_6985,N_6701);
nor U7804 (N_7804,N_6706,N_6426);
or U7805 (N_7805,N_6363,N_6544);
and U7806 (N_7806,N_6206,N_6897);
and U7807 (N_7807,N_6106,N_6773);
nor U7808 (N_7808,N_6567,N_6967);
and U7809 (N_7809,N_6937,N_6913);
nor U7810 (N_7810,N_6531,N_6701);
nand U7811 (N_7811,N_6713,N_6472);
nor U7812 (N_7812,N_6826,N_6476);
nor U7813 (N_7813,N_6376,N_6381);
nand U7814 (N_7814,N_6371,N_6718);
nor U7815 (N_7815,N_6575,N_6249);
and U7816 (N_7816,N_6791,N_6267);
nand U7817 (N_7817,N_6039,N_6696);
nand U7818 (N_7818,N_6322,N_6850);
nand U7819 (N_7819,N_6327,N_6649);
or U7820 (N_7820,N_6703,N_6300);
and U7821 (N_7821,N_6566,N_6750);
nor U7822 (N_7822,N_6876,N_6343);
nor U7823 (N_7823,N_6911,N_6428);
nor U7824 (N_7824,N_6596,N_6756);
or U7825 (N_7825,N_6870,N_6095);
nand U7826 (N_7826,N_6069,N_6864);
xnor U7827 (N_7827,N_6506,N_6660);
nand U7828 (N_7828,N_6090,N_6937);
nand U7829 (N_7829,N_6807,N_6723);
or U7830 (N_7830,N_6681,N_6436);
nand U7831 (N_7831,N_6648,N_6199);
and U7832 (N_7832,N_6868,N_6478);
and U7833 (N_7833,N_6168,N_6027);
nand U7834 (N_7834,N_6832,N_6685);
or U7835 (N_7835,N_6478,N_6965);
xor U7836 (N_7836,N_6869,N_6422);
or U7837 (N_7837,N_6194,N_6642);
xnor U7838 (N_7838,N_6075,N_6917);
or U7839 (N_7839,N_6458,N_6366);
nand U7840 (N_7840,N_6086,N_6745);
nand U7841 (N_7841,N_6406,N_6621);
or U7842 (N_7842,N_6948,N_6363);
xor U7843 (N_7843,N_6478,N_6998);
nor U7844 (N_7844,N_6919,N_6327);
nand U7845 (N_7845,N_6756,N_6044);
and U7846 (N_7846,N_6100,N_6676);
nand U7847 (N_7847,N_6989,N_6207);
nor U7848 (N_7848,N_6548,N_6184);
nor U7849 (N_7849,N_6917,N_6575);
xor U7850 (N_7850,N_6576,N_6258);
nor U7851 (N_7851,N_6333,N_6733);
nand U7852 (N_7852,N_6635,N_6421);
or U7853 (N_7853,N_6845,N_6056);
nor U7854 (N_7854,N_6362,N_6824);
or U7855 (N_7855,N_6137,N_6686);
xnor U7856 (N_7856,N_6551,N_6396);
nand U7857 (N_7857,N_6992,N_6529);
nand U7858 (N_7858,N_6734,N_6360);
or U7859 (N_7859,N_6159,N_6051);
and U7860 (N_7860,N_6367,N_6199);
or U7861 (N_7861,N_6240,N_6581);
xor U7862 (N_7862,N_6647,N_6593);
nand U7863 (N_7863,N_6191,N_6200);
nand U7864 (N_7864,N_6904,N_6538);
nor U7865 (N_7865,N_6100,N_6301);
nand U7866 (N_7866,N_6256,N_6491);
xor U7867 (N_7867,N_6484,N_6328);
and U7868 (N_7868,N_6186,N_6933);
xnor U7869 (N_7869,N_6903,N_6569);
nor U7870 (N_7870,N_6643,N_6365);
nor U7871 (N_7871,N_6339,N_6803);
nand U7872 (N_7872,N_6526,N_6427);
nor U7873 (N_7873,N_6163,N_6618);
and U7874 (N_7874,N_6502,N_6330);
nor U7875 (N_7875,N_6725,N_6486);
nand U7876 (N_7876,N_6152,N_6784);
or U7877 (N_7877,N_6105,N_6725);
nor U7878 (N_7878,N_6887,N_6632);
xor U7879 (N_7879,N_6818,N_6559);
nand U7880 (N_7880,N_6798,N_6608);
nand U7881 (N_7881,N_6591,N_6025);
xor U7882 (N_7882,N_6881,N_6062);
nor U7883 (N_7883,N_6102,N_6522);
nor U7884 (N_7884,N_6625,N_6716);
nand U7885 (N_7885,N_6913,N_6645);
or U7886 (N_7886,N_6053,N_6000);
nor U7887 (N_7887,N_6113,N_6396);
and U7888 (N_7888,N_6452,N_6853);
or U7889 (N_7889,N_6204,N_6748);
or U7890 (N_7890,N_6612,N_6001);
and U7891 (N_7891,N_6600,N_6762);
and U7892 (N_7892,N_6281,N_6483);
or U7893 (N_7893,N_6104,N_6784);
xor U7894 (N_7894,N_6222,N_6478);
nand U7895 (N_7895,N_6266,N_6100);
nor U7896 (N_7896,N_6782,N_6086);
xnor U7897 (N_7897,N_6438,N_6537);
or U7898 (N_7898,N_6148,N_6726);
nand U7899 (N_7899,N_6626,N_6486);
and U7900 (N_7900,N_6229,N_6646);
nor U7901 (N_7901,N_6739,N_6027);
nor U7902 (N_7902,N_6257,N_6412);
nor U7903 (N_7903,N_6621,N_6885);
nand U7904 (N_7904,N_6623,N_6272);
and U7905 (N_7905,N_6304,N_6151);
nand U7906 (N_7906,N_6536,N_6493);
xnor U7907 (N_7907,N_6521,N_6320);
xnor U7908 (N_7908,N_6456,N_6751);
nor U7909 (N_7909,N_6420,N_6957);
and U7910 (N_7910,N_6531,N_6764);
nand U7911 (N_7911,N_6548,N_6294);
xor U7912 (N_7912,N_6684,N_6314);
and U7913 (N_7913,N_6556,N_6483);
and U7914 (N_7914,N_6230,N_6238);
and U7915 (N_7915,N_6959,N_6180);
or U7916 (N_7916,N_6541,N_6458);
nor U7917 (N_7917,N_6332,N_6753);
nand U7918 (N_7918,N_6972,N_6006);
nor U7919 (N_7919,N_6566,N_6780);
xor U7920 (N_7920,N_6396,N_6211);
and U7921 (N_7921,N_6851,N_6470);
nand U7922 (N_7922,N_6593,N_6453);
or U7923 (N_7923,N_6914,N_6934);
nand U7924 (N_7924,N_6398,N_6278);
or U7925 (N_7925,N_6992,N_6612);
or U7926 (N_7926,N_6524,N_6578);
and U7927 (N_7927,N_6311,N_6045);
xnor U7928 (N_7928,N_6958,N_6239);
xor U7929 (N_7929,N_6602,N_6793);
nand U7930 (N_7930,N_6519,N_6293);
xnor U7931 (N_7931,N_6514,N_6731);
or U7932 (N_7932,N_6261,N_6335);
and U7933 (N_7933,N_6314,N_6364);
or U7934 (N_7934,N_6469,N_6765);
nor U7935 (N_7935,N_6241,N_6629);
and U7936 (N_7936,N_6173,N_6840);
nor U7937 (N_7937,N_6643,N_6925);
nand U7938 (N_7938,N_6986,N_6621);
nand U7939 (N_7939,N_6683,N_6734);
and U7940 (N_7940,N_6200,N_6313);
or U7941 (N_7941,N_6338,N_6522);
and U7942 (N_7942,N_6934,N_6999);
nor U7943 (N_7943,N_6801,N_6007);
nor U7944 (N_7944,N_6187,N_6075);
and U7945 (N_7945,N_6519,N_6899);
and U7946 (N_7946,N_6051,N_6269);
xnor U7947 (N_7947,N_6399,N_6856);
and U7948 (N_7948,N_6391,N_6186);
nand U7949 (N_7949,N_6881,N_6045);
xnor U7950 (N_7950,N_6960,N_6491);
nor U7951 (N_7951,N_6071,N_6684);
xor U7952 (N_7952,N_6473,N_6566);
and U7953 (N_7953,N_6693,N_6510);
nand U7954 (N_7954,N_6797,N_6447);
and U7955 (N_7955,N_6014,N_6449);
nand U7956 (N_7956,N_6409,N_6891);
nand U7957 (N_7957,N_6813,N_6273);
nand U7958 (N_7958,N_6836,N_6473);
or U7959 (N_7959,N_6702,N_6487);
nand U7960 (N_7960,N_6635,N_6983);
nand U7961 (N_7961,N_6334,N_6709);
or U7962 (N_7962,N_6105,N_6041);
and U7963 (N_7963,N_6747,N_6504);
nor U7964 (N_7964,N_6129,N_6080);
xor U7965 (N_7965,N_6177,N_6578);
xor U7966 (N_7966,N_6267,N_6524);
nand U7967 (N_7967,N_6810,N_6577);
and U7968 (N_7968,N_6138,N_6382);
xor U7969 (N_7969,N_6133,N_6375);
nand U7970 (N_7970,N_6968,N_6914);
nand U7971 (N_7971,N_6219,N_6123);
or U7972 (N_7972,N_6950,N_6104);
or U7973 (N_7973,N_6547,N_6201);
nand U7974 (N_7974,N_6253,N_6023);
nor U7975 (N_7975,N_6502,N_6276);
nor U7976 (N_7976,N_6880,N_6645);
xnor U7977 (N_7977,N_6745,N_6372);
or U7978 (N_7978,N_6219,N_6389);
xnor U7979 (N_7979,N_6630,N_6307);
and U7980 (N_7980,N_6761,N_6317);
nand U7981 (N_7981,N_6732,N_6050);
xnor U7982 (N_7982,N_6653,N_6495);
xnor U7983 (N_7983,N_6661,N_6499);
xnor U7984 (N_7984,N_6557,N_6393);
nor U7985 (N_7985,N_6240,N_6747);
nand U7986 (N_7986,N_6152,N_6569);
nand U7987 (N_7987,N_6304,N_6157);
xor U7988 (N_7988,N_6421,N_6619);
xnor U7989 (N_7989,N_6092,N_6297);
and U7990 (N_7990,N_6981,N_6698);
nor U7991 (N_7991,N_6156,N_6437);
nand U7992 (N_7992,N_6482,N_6884);
nand U7993 (N_7993,N_6558,N_6354);
xor U7994 (N_7994,N_6258,N_6036);
and U7995 (N_7995,N_6678,N_6586);
nand U7996 (N_7996,N_6054,N_6313);
nor U7997 (N_7997,N_6218,N_6395);
and U7998 (N_7998,N_6763,N_6540);
nand U7999 (N_7999,N_6790,N_6133);
nor U8000 (N_8000,N_7267,N_7486);
xnor U8001 (N_8001,N_7118,N_7078);
nand U8002 (N_8002,N_7769,N_7091);
and U8003 (N_8003,N_7908,N_7972);
xnor U8004 (N_8004,N_7669,N_7414);
or U8005 (N_8005,N_7058,N_7152);
nand U8006 (N_8006,N_7348,N_7060);
or U8007 (N_8007,N_7073,N_7300);
or U8008 (N_8008,N_7625,N_7920);
nor U8009 (N_8009,N_7638,N_7210);
and U8010 (N_8010,N_7855,N_7956);
and U8011 (N_8011,N_7911,N_7951);
or U8012 (N_8012,N_7453,N_7420);
or U8013 (N_8013,N_7179,N_7438);
xnor U8014 (N_8014,N_7359,N_7460);
or U8015 (N_8015,N_7514,N_7699);
nor U8016 (N_8016,N_7935,N_7484);
and U8017 (N_8017,N_7451,N_7431);
or U8018 (N_8018,N_7067,N_7954);
nor U8019 (N_8019,N_7435,N_7527);
nand U8020 (N_8020,N_7618,N_7955);
nor U8021 (N_8021,N_7286,N_7900);
xnor U8022 (N_8022,N_7469,N_7182);
and U8023 (N_8023,N_7052,N_7779);
xnor U8024 (N_8024,N_7958,N_7965);
nor U8025 (N_8025,N_7086,N_7532);
or U8026 (N_8026,N_7545,N_7026);
nand U8027 (N_8027,N_7500,N_7934);
nor U8028 (N_8028,N_7032,N_7491);
nor U8029 (N_8029,N_7044,N_7045);
or U8030 (N_8030,N_7553,N_7903);
xnor U8031 (N_8031,N_7861,N_7998);
or U8032 (N_8032,N_7054,N_7860);
nor U8033 (N_8033,N_7439,N_7391);
or U8034 (N_8034,N_7971,N_7433);
xor U8035 (N_8035,N_7876,N_7108);
xnor U8036 (N_8036,N_7242,N_7105);
nand U8037 (N_8037,N_7726,N_7866);
and U8038 (N_8038,N_7477,N_7253);
and U8039 (N_8039,N_7331,N_7260);
and U8040 (N_8040,N_7762,N_7790);
or U8041 (N_8041,N_7795,N_7661);
xor U8042 (N_8042,N_7436,N_7016);
xnor U8043 (N_8043,N_7133,N_7275);
or U8044 (N_8044,N_7796,N_7813);
and U8045 (N_8045,N_7266,N_7428);
nor U8046 (N_8046,N_7290,N_7150);
or U8047 (N_8047,N_7333,N_7881);
and U8048 (N_8048,N_7406,N_7776);
and U8049 (N_8049,N_7894,N_7544);
and U8050 (N_8050,N_7159,N_7383);
or U8051 (N_8051,N_7684,N_7847);
xnor U8052 (N_8052,N_7364,N_7960);
nor U8053 (N_8053,N_7330,N_7172);
or U8054 (N_8054,N_7385,N_7691);
and U8055 (N_8055,N_7094,N_7234);
nor U8056 (N_8056,N_7768,N_7719);
and U8057 (N_8057,N_7495,N_7791);
xnor U8058 (N_8058,N_7156,N_7176);
nand U8059 (N_8059,N_7656,N_7307);
nand U8060 (N_8060,N_7799,N_7189);
nand U8061 (N_8061,N_7465,N_7205);
nand U8062 (N_8062,N_7830,N_7015);
xnor U8063 (N_8063,N_7147,N_7593);
nor U8064 (N_8064,N_7503,N_7072);
nor U8065 (N_8065,N_7419,N_7539);
or U8066 (N_8066,N_7734,N_7758);
and U8067 (N_8067,N_7910,N_7884);
nand U8068 (N_8068,N_7224,N_7896);
xor U8069 (N_8069,N_7890,N_7766);
and U8070 (N_8070,N_7740,N_7035);
xnor U8071 (N_8071,N_7280,N_7327);
xor U8072 (N_8072,N_7301,N_7243);
and U8073 (N_8073,N_7009,N_7181);
or U8074 (N_8074,N_7975,N_7631);
or U8075 (N_8075,N_7562,N_7113);
and U8076 (N_8076,N_7199,N_7195);
xnor U8077 (N_8077,N_7706,N_7028);
nor U8078 (N_8078,N_7867,N_7774);
and U8079 (N_8079,N_7238,N_7640);
nor U8080 (N_8080,N_7013,N_7744);
xor U8081 (N_8081,N_7427,N_7747);
nand U8082 (N_8082,N_7127,N_7843);
nand U8083 (N_8083,N_7621,N_7980);
nand U8084 (N_8084,N_7175,N_7422);
or U8085 (N_8085,N_7240,N_7700);
and U8086 (N_8086,N_7184,N_7627);
nand U8087 (N_8087,N_7565,N_7952);
xnor U8088 (N_8088,N_7670,N_7467);
xor U8089 (N_8089,N_7763,N_7639);
and U8090 (N_8090,N_7668,N_7513);
nand U8091 (N_8091,N_7851,N_7564);
nor U8092 (N_8092,N_7711,N_7114);
xor U8093 (N_8093,N_7720,N_7589);
nand U8094 (N_8094,N_7079,N_7745);
or U8095 (N_8095,N_7981,N_7966);
xor U8096 (N_8096,N_7308,N_7987);
nor U8097 (N_8097,N_7212,N_7628);
nor U8098 (N_8098,N_7658,N_7029);
nor U8099 (N_8099,N_7852,N_7213);
nand U8100 (N_8100,N_7268,N_7722);
nand U8101 (N_8101,N_7974,N_7694);
or U8102 (N_8102,N_7686,N_7917);
nor U8103 (N_8103,N_7816,N_7347);
xnor U8104 (N_8104,N_7022,N_7757);
or U8105 (N_8105,N_7546,N_7374);
nand U8106 (N_8106,N_7755,N_7217);
and U8107 (N_8107,N_7794,N_7613);
or U8108 (N_8108,N_7927,N_7895);
and U8109 (N_8109,N_7397,N_7031);
nand U8110 (N_8110,N_7899,N_7509);
or U8111 (N_8111,N_7069,N_7925);
nor U8112 (N_8112,N_7050,N_7919);
nand U8113 (N_8113,N_7575,N_7186);
and U8114 (N_8114,N_7723,N_7116);
nor U8115 (N_8115,N_7271,N_7001);
and U8116 (N_8116,N_7842,N_7992);
and U8117 (N_8117,N_7311,N_7335);
xor U8118 (N_8118,N_7528,N_7141);
or U8119 (N_8119,N_7521,N_7402);
or U8120 (N_8120,N_7106,N_7540);
nor U8121 (N_8121,N_7939,N_7529);
or U8122 (N_8122,N_7440,N_7426);
or U8123 (N_8123,N_7702,N_7446);
xnor U8124 (N_8124,N_7797,N_7246);
and U8125 (N_8125,N_7211,N_7568);
xor U8126 (N_8126,N_7735,N_7407);
or U8127 (N_8127,N_7019,N_7125);
xor U8128 (N_8128,N_7024,N_7101);
and U8129 (N_8129,N_7765,N_7090);
and U8130 (N_8130,N_7056,N_7368);
xnor U8131 (N_8131,N_7134,N_7983);
nand U8132 (N_8132,N_7321,N_7635);
nand U8133 (N_8133,N_7102,N_7148);
or U8134 (N_8134,N_7778,N_7736);
or U8135 (N_8135,N_7355,N_7690);
nand U8136 (N_8136,N_7077,N_7360);
nand U8137 (N_8137,N_7023,N_7109);
and U8138 (N_8138,N_7817,N_7695);
nor U8139 (N_8139,N_7390,N_7315);
or U8140 (N_8140,N_7902,N_7815);
or U8141 (N_8141,N_7168,N_7284);
xor U8142 (N_8142,N_7493,N_7689);
and U8143 (N_8143,N_7076,N_7898);
xor U8144 (N_8144,N_7207,N_7456);
nor U8145 (N_8145,N_7993,N_7709);
nand U8146 (N_8146,N_7558,N_7443);
nor U8147 (N_8147,N_7226,N_7617);
nand U8148 (N_8148,N_7649,N_7957);
or U8149 (N_8149,N_7976,N_7646);
nor U8150 (N_8150,N_7637,N_7345);
xor U8151 (N_8151,N_7384,N_7142);
or U8152 (N_8152,N_7128,N_7615);
nor U8153 (N_8153,N_7018,N_7276);
nor U8154 (N_8154,N_7551,N_7804);
xnor U8155 (N_8155,N_7346,N_7025);
and U8156 (N_8156,N_7888,N_7525);
xor U8157 (N_8157,N_7233,N_7490);
or U8158 (N_8158,N_7724,N_7258);
nor U8159 (N_8159,N_7798,N_7096);
nand U8160 (N_8160,N_7550,N_7279);
or U8161 (N_8161,N_7732,N_7319);
nor U8162 (N_8162,N_7288,N_7496);
or U8163 (N_8163,N_7962,N_7468);
xnor U8164 (N_8164,N_7120,N_7512);
and U8165 (N_8165,N_7294,N_7809);
xor U8166 (N_8166,N_7961,N_7985);
nand U8167 (N_8167,N_7892,N_7098);
and U8168 (N_8168,N_7097,N_7413);
xnor U8169 (N_8169,N_7715,N_7472);
nor U8170 (N_8170,N_7520,N_7158);
nand U8171 (N_8171,N_7585,N_7714);
xnor U8172 (N_8172,N_7357,N_7606);
or U8173 (N_8173,N_7020,N_7561);
and U8174 (N_8174,N_7633,N_7208);
nor U8175 (N_8175,N_7004,N_7062);
xnor U8176 (N_8176,N_7990,N_7704);
or U8177 (N_8177,N_7832,N_7773);
or U8178 (N_8178,N_7857,N_7746);
nor U8179 (N_8179,N_7377,N_7683);
or U8180 (N_8180,N_7573,N_7143);
and U8181 (N_8181,N_7375,N_7862);
nor U8182 (N_8182,N_7687,N_7787);
or U8183 (N_8183,N_7250,N_7257);
nand U8184 (N_8184,N_7169,N_7249);
xnor U8185 (N_8185,N_7444,N_7567);
and U8186 (N_8186,N_7873,N_7466);
or U8187 (N_8187,N_7655,N_7201);
and U8188 (N_8188,N_7111,N_7400);
nor U8189 (N_8189,N_7767,N_7449);
and U8190 (N_8190,N_7929,N_7808);
nand U8191 (N_8191,N_7821,N_7274);
nand U8192 (N_8192,N_7382,N_7534);
xnor U8193 (N_8193,N_7964,N_7818);
or U8194 (N_8194,N_7581,N_7462);
nor U8195 (N_8195,N_7164,N_7997);
nor U8196 (N_8196,N_7916,N_7886);
nand U8197 (N_8197,N_7314,N_7144);
xnor U8198 (N_8198,N_7488,N_7342);
nor U8199 (N_8199,N_7410,N_7296);
and U8200 (N_8200,N_7068,N_7930);
xnor U8201 (N_8201,N_7666,N_7577);
and U8202 (N_8202,N_7829,N_7423);
xnor U8203 (N_8203,N_7063,N_7629);
xnor U8204 (N_8204,N_7188,N_7877);
nor U8205 (N_8205,N_7672,N_7584);
xor U8206 (N_8206,N_7252,N_7070);
xor U8207 (N_8207,N_7351,N_7064);
nand U8208 (N_8208,N_7826,N_7283);
nor U8209 (N_8209,N_7474,N_7675);
nor U8210 (N_8210,N_7075,N_7986);
nand U8211 (N_8211,N_7285,N_7479);
and U8212 (N_8212,N_7445,N_7055);
and U8213 (N_8213,N_7576,N_7918);
nor U8214 (N_8214,N_7478,N_7858);
nand U8215 (N_8215,N_7729,N_7800);
and U8216 (N_8216,N_7601,N_7340);
and U8217 (N_8217,N_7667,N_7921);
nor U8218 (N_8218,N_7865,N_7953);
xnor U8219 (N_8219,N_7708,N_7730);
or U8220 (N_8220,N_7978,N_7557);
or U8221 (N_8221,N_7543,N_7489);
nand U8222 (N_8222,N_7552,N_7620);
and U8223 (N_8223,N_7149,N_7781);
nor U8224 (N_8224,N_7185,N_7053);
xnor U8225 (N_8225,N_7115,N_7614);
xnor U8226 (N_8226,N_7942,N_7030);
nand U8227 (N_8227,N_7306,N_7662);
and U8228 (N_8228,N_7739,N_7681);
nand U8229 (N_8229,N_7411,N_7136);
xor U8230 (N_8230,N_7559,N_7356);
or U8231 (N_8231,N_7157,N_7932);
and U8232 (N_8232,N_7713,N_7906);
or U8233 (N_8233,N_7705,N_7872);
xor U8234 (N_8234,N_7220,N_7623);
nand U8235 (N_8235,N_7047,N_7678);
or U8236 (N_8236,N_7295,N_7820);
and U8237 (N_8237,N_7508,N_7569);
or U8238 (N_8238,N_7756,N_7727);
xor U8239 (N_8239,N_7177,N_7570);
nand U8240 (N_8240,N_7760,N_7262);
nor U8241 (N_8241,N_7297,N_7261);
and U8242 (N_8242,N_7145,N_7178);
or U8243 (N_8243,N_7256,N_7470);
or U8244 (N_8244,N_7594,N_7441);
nand U8245 (N_8245,N_7793,N_7463);
nand U8246 (N_8246,N_7416,N_7963);
and U8247 (N_8247,N_7448,N_7783);
nand U8248 (N_8248,N_7671,N_7556);
nor U8249 (N_8249,N_7092,N_7547);
nor U8250 (N_8250,N_7278,N_7772);
xor U8251 (N_8251,N_7352,N_7037);
nor U8252 (N_8252,N_7457,N_7395);
and U8253 (N_8253,N_7313,N_7322);
and U8254 (N_8254,N_7560,N_7324);
or U8255 (N_8255,N_7535,N_7389);
and U8256 (N_8256,N_7394,N_7247);
xnor U8257 (N_8257,N_7138,N_7982);
nand U8258 (N_8258,N_7653,N_7000);
nor U8259 (N_8259,N_7583,N_7650);
xor U8260 (N_8260,N_7905,N_7874);
and U8261 (N_8261,N_7945,N_7541);
nor U8262 (N_8262,N_7840,N_7648);
nand U8263 (N_8263,N_7354,N_7447);
nand U8264 (N_8264,N_7731,N_7586);
nand U8265 (N_8265,N_7046,N_7819);
nand U8266 (N_8266,N_7785,N_7225);
and U8267 (N_8267,N_7464,N_7007);
or U8268 (N_8268,N_7844,N_7519);
nor U8269 (N_8269,N_7043,N_7329);
xor U8270 (N_8270,N_7891,N_7598);
xor U8271 (N_8271,N_7511,N_7538);
xnor U8272 (N_8272,N_7434,N_7171);
or U8273 (N_8273,N_7458,N_7880);
xor U8274 (N_8274,N_7636,N_7893);
or U8275 (N_8275,N_7728,N_7362);
nor U8276 (N_8276,N_7856,N_7337);
xor U8277 (N_8277,N_7265,N_7599);
or U8278 (N_8278,N_7017,N_7163);
or U8279 (N_8279,N_7282,N_7619);
nand U8280 (N_8280,N_7034,N_7518);
and U8281 (N_8281,N_7170,N_7167);
xnor U8282 (N_8282,N_7198,N_7940);
xnor U8283 (N_8283,N_7721,N_7802);
or U8284 (N_8284,N_7970,N_7782);
xor U8285 (N_8285,N_7595,N_7753);
nand U8286 (N_8286,N_7379,N_7775);
nand U8287 (N_8287,N_7200,N_7483);
nand U8288 (N_8288,N_7973,N_7049);
xnor U8289 (N_8289,N_7269,N_7372);
nor U8290 (N_8290,N_7151,N_7679);
xor U8291 (N_8291,N_7692,N_7165);
xor U8292 (N_8292,N_7287,N_7823);
xnor U8293 (N_8293,N_7602,N_7701);
and U8294 (N_8294,N_7989,N_7237);
xnor U8295 (N_8295,N_7580,N_7089);
or U8296 (N_8296,N_7381,N_7574);
nand U8297 (N_8297,N_7155,N_7825);
xnor U8298 (N_8298,N_7688,N_7241);
xor U8299 (N_8299,N_7251,N_7338);
nand U8300 (N_8300,N_7771,N_7473);
nand U8301 (N_8301,N_7291,N_7475);
and U8302 (N_8302,N_7792,N_7239);
and U8303 (N_8303,N_7537,N_7343);
nand U8304 (N_8304,N_7572,N_7405);
nand U8305 (N_8305,N_7641,N_7471);
and U8306 (N_8306,N_7751,N_7011);
nand U8307 (N_8307,N_7350,N_7310);
or U8308 (N_8308,N_7871,N_7897);
and U8309 (N_8309,N_7303,N_7624);
and U8310 (N_8310,N_7353,N_7612);
or U8311 (N_8311,N_7376,N_7845);
xor U8312 (N_8312,N_7707,N_7947);
or U8313 (N_8313,N_7870,N_7716);
xnor U8314 (N_8314,N_7616,N_7008);
and U8315 (N_8315,N_7859,N_7923);
nand U8316 (N_8316,N_7677,N_7270);
and U8317 (N_8317,N_7733,N_7788);
nor U8318 (N_8318,N_7487,N_7454);
and U8319 (N_8319,N_7418,N_7033);
xor U8320 (N_8320,N_7481,N_7632);
nand U8321 (N_8321,N_7273,N_7216);
xor U8322 (N_8322,N_7083,N_7183);
or U8323 (N_8323,N_7010,N_7834);
or U8324 (N_8324,N_7305,N_7074);
nor U8325 (N_8325,N_7944,N_7991);
xor U8326 (N_8326,N_7837,N_7373);
nor U8327 (N_8327,N_7725,N_7254);
xnor U8328 (N_8328,N_7588,N_7380);
nand U8329 (N_8329,N_7741,N_7281);
nor U8330 (N_8330,N_7759,N_7318);
nand U8331 (N_8331,N_7738,N_7194);
nor U8332 (N_8332,N_7071,N_7665);
nor U8333 (N_8333,N_7430,N_7367);
nor U8334 (N_8334,N_7365,N_7664);
and U8335 (N_8335,N_7084,N_7603);
or U8336 (N_8336,N_7309,N_7742);
nand U8337 (N_8337,N_7810,N_7928);
or U8338 (N_8338,N_7875,N_7085);
or U8339 (N_8339,N_7680,N_7949);
xnor U8340 (N_8340,N_7126,N_7780);
xor U8341 (N_8341,N_7931,N_7304);
xor U8342 (N_8342,N_7979,N_7135);
nand U8343 (N_8343,N_7036,N_7263);
nor U8344 (N_8344,N_7203,N_7663);
xnor U8345 (N_8345,N_7103,N_7597);
nor U8346 (N_8346,N_7968,N_7137);
nand U8347 (N_8347,N_7432,N_7801);
xor U8348 (N_8348,N_7039,N_7107);
nor U8349 (N_8349,N_7232,N_7904);
nor U8350 (N_8350,N_7202,N_7429);
nor U8351 (N_8351,N_7501,N_7235);
nand U8352 (N_8352,N_7849,N_7227);
or U8353 (N_8353,N_7206,N_7222);
or U8354 (N_8354,N_7421,N_7196);
nand U8355 (N_8355,N_7048,N_7644);
and U8356 (N_8356,N_7839,N_7082);
nor U8357 (N_8357,N_7388,N_7600);
nor U8358 (N_8358,N_7409,N_7937);
xor U8359 (N_8359,N_7673,N_7889);
xnor U8360 (N_8360,N_7634,N_7698);
xor U8361 (N_8361,N_7882,N_7883);
nand U8362 (N_8362,N_7230,N_7061);
nand U8363 (N_8363,N_7166,N_7838);
or U8364 (N_8364,N_7909,N_7292);
nor U8365 (N_8365,N_7850,N_7228);
nor U8366 (N_8366,N_7566,N_7450);
nor U8367 (N_8367,N_7153,N_7645);
or U8368 (N_8368,N_7459,N_7610);
nand U8369 (N_8369,N_7626,N_7912);
nor U8370 (N_8370,N_7363,N_7946);
and U8371 (N_8371,N_7192,N_7885);
and U8372 (N_8372,N_7130,N_7807);
xor U8373 (N_8373,N_7869,N_7334);
nand U8374 (N_8374,N_7786,N_7517);
xnor U8375 (N_8375,N_7272,N_7293);
or U8376 (N_8376,N_7104,N_7948);
xor U8377 (N_8377,N_7219,N_7370);
nand U8378 (N_8378,N_7160,N_7504);
nand U8379 (N_8379,N_7914,N_7879);
and U8380 (N_8380,N_7651,N_7323);
nand U8381 (N_8381,N_7643,N_7361);
and U8382 (N_8382,N_7339,N_7591);
nor U8383 (N_8383,N_7093,N_7396);
nand U8384 (N_8384,N_7642,N_7831);
nand U8385 (N_8385,N_7784,N_7320);
xnor U8386 (N_8386,N_7833,N_7259);
or U8387 (N_8387,N_7789,N_7401);
or U8388 (N_8388,N_7326,N_7516);
nand U8389 (N_8389,N_7002,N_7846);
nand U8390 (N_8390,N_7289,N_7492);
nand U8391 (N_8391,N_7040,N_7041);
or U8392 (N_8392,N_7828,N_7996);
and U8393 (N_8393,N_7827,N_7922);
or U8394 (N_8394,N_7554,N_7542);
and U8395 (N_8395,N_7012,N_7341);
or U8396 (N_8396,N_7131,N_7386);
xnor U8397 (N_8397,N_7737,N_7592);
or U8398 (N_8398,N_7197,N_7424);
nand U8399 (N_8399,N_7387,N_7915);
xnor U8400 (N_8400,N_7485,N_7298);
and U8401 (N_8401,N_7657,N_7999);
and U8402 (N_8402,N_7578,N_7214);
nand U8403 (N_8403,N_7836,N_7536);
xnor U8404 (N_8404,N_7605,N_7607);
nor U8405 (N_8405,N_7476,N_7506);
nor U8406 (N_8406,N_7878,N_7452);
nand U8407 (N_8407,N_7674,N_7193);
or U8408 (N_8408,N_7676,N_7480);
nand U8409 (N_8409,N_7812,N_7995);
and U8410 (N_8410,N_7712,N_7693);
and U8411 (N_8411,N_7938,N_7393);
nand U8412 (N_8412,N_7984,N_7317);
and U8413 (N_8413,N_7173,N_7936);
xor U8414 (N_8414,N_7523,N_7571);
or U8415 (N_8415,N_7209,N_7924);
nor U8416 (N_8416,N_7630,N_7926);
and U8417 (N_8417,N_7191,N_7065);
xnor U8418 (N_8418,N_7455,N_7498);
and U8419 (N_8419,N_7682,N_7822);
nor U8420 (N_8420,N_7132,N_7121);
nand U8421 (N_8421,N_7579,N_7215);
nor U8422 (N_8422,N_7277,N_7392);
xnor U8423 (N_8423,N_7764,N_7081);
xor U8424 (N_8424,N_7110,N_7187);
xnor U8425 (N_8425,N_7328,N_7522);
or U8426 (N_8426,N_7750,N_7358);
nand U8427 (N_8427,N_7408,N_7398);
and U8428 (N_8428,N_7425,N_7505);
or U8429 (N_8429,N_7442,N_7122);
nor U8430 (N_8430,N_7752,N_7696);
xor U8431 (N_8431,N_7006,N_7814);
nor U8432 (N_8432,N_7119,N_7190);
or U8433 (N_8433,N_7369,N_7229);
and U8434 (N_8434,N_7057,N_7336);
xor U8435 (N_8435,N_7042,N_7231);
nand U8436 (N_8436,N_7497,N_7112);
or U8437 (N_8437,N_7703,N_7654);
nor U8438 (N_8438,N_7563,N_7848);
xor U8439 (N_8439,N_7038,N_7959);
nand U8440 (N_8440,N_7587,N_7059);
and U8441 (N_8441,N_7245,N_7549);
or U8442 (N_8442,N_7853,N_7236);
or U8443 (N_8443,N_7066,N_7003);
nand U8444 (N_8444,N_7531,N_7095);
xnor U8445 (N_8445,N_7652,N_7660);
nand U8446 (N_8446,N_7988,N_7332);
and U8447 (N_8447,N_7590,N_7913);
nor U8448 (N_8448,N_7622,N_7099);
nand U8449 (N_8449,N_7510,N_7868);
xnor U8450 (N_8450,N_7461,N_7854);
or U8451 (N_8451,N_7901,N_7754);
nand U8452 (N_8452,N_7977,N_7161);
or U8453 (N_8453,N_7950,N_7088);
and U8454 (N_8454,N_7717,N_7806);
nor U8455 (N_8455,N_7967,N_7051);
or U8456 (N_8456,N_7117,N_7811);
and U8457 (N_8457,N_7941,N_7146);
nand U8458 (N_8458,N_7969,N_7710);
xnor U8459 (N_8459,N_7611,N_7994);
and U8460 (N_8460,N_7604,N_7697);
and U8461 (N_8461,N_7399,N_7749);
and U8462 (N_8462,N_7404,N_7123);
nor U8463 (N_8463,N_7933,N_7533);
nor U8464 (N_8464,N_7582,N_7803);
or U8465 (N_8465,N_7255,N_7526);
nor U8466 (N_8466,N_7080,N_7863);
xnor U8467 (N_8467,N_7366,N_7087);
nor U8468 (N_8468,N_7403,N_7264);
xor U8469 (N_8469,N_7417,N_7344);
nor U8470 (N_8470,N_7378,N_7349);
and U8471 (N_8471,N_7223,N_7743);
nand U8472 (N_8472,N_7302,N_7777);
nand U8473 (N_8473,N_7596,N_7415);
and U8474 (N_8474,N_7805,N_7499);
xnor U8475 (N_8475,N_7021,N_7180);
and U8476 (N_8476,N_7835,N_7014);
nor U8477 (N_8477,N_7530,N_7371);
xnor U8478 (N_8478,N_7139,N_7412);
nand U8479 (N_8479,N_7943,N_7907);
nand U8480 (N_8480,N_7027,N_7129);
xor U8481 (N_8481,N_7312,N_7005);
nor U8482 (N_8482,N_7162,N_7548);
or U8483 (N_8483,N_7609,N_7316);
nor U8484 (N_8484,N_7524,N_7244);
and U8485 (N_8485,N_7770,N_7718);
and U8486 (N_8486,N_7124,N_7299);
or U8487 (N_8487,N_7824,N_7748);
xor U8488 (N_8488,N_7647,N_7659);
xnor U8489 (N_8489,N_7502,N_7437);
or U8490 (N_8490,N_7325,N_7174);
nand U8491 (N_8491,N_7221,N_7864);
nand U8492 (N_8492,N_7100,N_7218);
xnor U8493 (N_8493,N_7154,N_7608);
or U8494 (N_8494,N_7555,N_7515);
nor U8495 (N_8495,N_7248,N_7685);
nand U8496 (N_8496,N_7204,N_7482);
nand U8497 (N_8497,N_7140,N_7841);
nor U8498 (N_8498,N_7887,N_7507);
nand U8499 (N_8499,N_7761,N_7494);
nor U8500 (N_8500,N_7153,N_7429);
nor U8501 (N_8501,N_7514,N_7941);
nor U8502 (N_8502,N_7360,N_7004);
xnor U8503 (N_8503,N_7487,N_7181);
nor U8504 (N_8504,N_7185,N_7308);
nor U8505 (N_8505,N_7177,N_7846);
or U8506 (N_8506,N_7874,N_7632);
xnor U8507 (N_8507,N_7167,N_7141);
nor U8508 (N_8508,N_7057,N_7948);
nor U8509 (N_8509,N_7470,N_7541);
and U8510 (N_8510,N_7352,N_7134);
xor U8511 (N_8511,N_7974,N_7781);
nand U8512 (N_8512,N_7092,N_7060);
nor U8513 (N_8513,N_7481,N_7454);
or U8514 (N_8514,N_7628,N_7053);
nor U8515 (N_8515,N_7542,N_7407);
xor U8516 (N_8516,N_7964,N_7424);
or U8517 (N_8517,N_7097,N_7454);
nor U8518 (N_8518,N_7029,N_7981);
or U8519 (N_8519,N_7147,N_7447);
xor U8520 (N_8520,N_7159,N_7636);
and U8521 (N_8521,N_7076,N_7522);
nor U8522 (N_8522,N_7622,N_7546);
or U8523 (N_8523,N_7352,N_7950);
or U8524 (N_8524,N_7266,N_7585);
and U8525 (N_8525,N_7817,N_7826);
nand U8526 (N_8526,N_7082,N_7751);
nand U8527 (N_8527,N_7335,N_7488);
or U8528 (N_8528,N_7201,N_7803);
xnor U8529 (N_8529,N_7704,N_7270);
xnor U8530 (N_8530,N_7911,N_7990);
and U8531 (N_8531,N_7643,N_7394);
or U8532 (N_8532,N_7845,N_7430);
nor U8533 (N_8533,N_7390,N_7169);
xnor U8534 (N_8534,N_7199,N_7565);
or U8535 (N_8535,N_7745,N_7191);
or U8536 (N_8536,N_7707,N_7003);
nor U8537 (N_8537,N_7453,N_7559);
and U8538 (N_8538,N_7902,N_7822);
nor U8539 (N_8539,N_7974,N_7557);
xnor U8540 (N_8540,N_7913,N_7810);
nor U8541 (N_8541,N_7959,N_7310);
or U8542 (N_8542,N_7964,N_7715);
and U8543 (N_8543,N_7021,N_7100);
and U8544 (N_8544,N_7863,N_7343);
and U8545 (N_8545,N_7144,N_7658);
nand U8546 (N_8546,N_7869,N_7676);
nand U8547 (N_8547,N_7424,N_7725);
nor U8548 (N_8548,N_7222,N_7467);
xnor U8549 (N_8549,N_7556,N_7572);
nor U8550 (N_8550,N_7588,N_7239);
and U8551 (N_8551,N_7601,N_7356);
nor U8552 (N_8552,N_7435,N_7193);
nand U8553 (N_8553,N_7584,N_7848);
nand U8554 (N_8554,N_7093,N_7120);
and U8555 (N_8555,N_7709,N_7959);
nor U8556 (N_8556,N_7080,N_7322);
and U8557 (N_8557,N_7895,N_7320);
xnor U8558 (N_8558,N_7682,N_7481);
and U8559 (N_8559,N_7297,N_7407);
or U8560 (N_8560,N_7414,N_7973);
nand U8561 (N_8561,N_7160,N_7143);
nand U8562 (N_8562,N_7638,N_7031);
nand U8563 (N_8563,N_7151,N_7378);
nor U8564 (N_8564,N_7367,N_7149);
and U8565 (N_8565,N_7403,N_7946);
nand U8566 (N_8566,N_7581,N_7896);
and U8567 (N_8567,N_7540,N_7108);
and U8568 (N_8568,N_7978,N_7897);
and U8569 (N_8569,N_7030,N_7134);
and U8570 (N_8570,N_7651,N_7541);
or U8571 (N_8571,N_7946,N_7455);
nor U8572 (N_8572,N_7010,N_7353);
and U8573 (N_8573,N_7274,N_7188);
or U8574 (N_8574,N_7994,N_7199);
or U8575 (N_8575,N_7287,N_7840);
xnor U8576 (N_8576,N_7635,N_7190);
nand U8577 (N_8577,N_7580,N_7943);
nand U8578 (N_8578,N_7099,N_7350);
nor U8579 (N_8579,N_7717,N_7753);
and U8580 (N_8580,N_7331,N_7485);
or U8581 (N_8581,N_7818,N_7840);
and U8582 (N_8582,N_7487,N_7107);
xor U8583 (N_8583,N_7506,N_7926);
nor U8584 (N_8584,N_7336,N_7654);
nand U8585 (N_8585,N_7522,N_7302);
nand U8586 (N_8586,N_7073,N_7789);
xor U8587 (N_8587,N_7737,N_7338);
nand U8588 (N_8588,N_7820,N_7237);
xnor U8589 (N_8589,N_7912,N_7783);
and U8590 (N_8590,N_7236,N_7235);
xor U8591 (N_8591,N_7517,N_7087);
nor U8592 (N_8592,N_7862,N_7509);
and U8593 (N_8593,N_7715,N_7746);
or U8594 (N_8594,N_7730,N_7103);
xnor U8595 (N_8595,N_7540,N_7810);
nor U8596 (N_8596,N_7748,N_7556);
xnor U8597 (N_8597,N_7713,N_7217);
nand U8598 (N_8598,N_7077,N_7647);
and U8599 (N_8599,N_7561,N_7973);
or U8600 (N_8600,N_7624,N_7210);
nor U8601 (N_8601,N_7643,N_7511);
xor U8602 (N_8602,N_7650,N_7651);
or U8603 (N_8603,N_7557,N_7356);
or U8604 (N_8604,N_7214,N_7216);
nor U8605 (N_8605,N_7683,N_7847);
xor U8606 (N_8606,N_7629,N_7788);
nand U8607 (N_8607,N_7258,N_7464);
xnor U8608 (N_8608,N_7842,N_7680);
or U8609 (N_8609,N_7923,N_7553);
xnor U8610 (N_8610,N_7658,N_7325);
and U8611 (N_8611,N_7683,N_7151);
or U8612 (N_8612,N_7176,N_7382);
and U8613 (N_8613,N_7668,N_7454);
or U8614 (N_8614,N_7227,N_7812);
nor U8615 (N_8615,N_7155,N_7087);
or U8616 (N_8616,N_7300,N_7775);
and U8617 (N_8617,N_7885,N_7162);
nand U8618 (N_8618,N_7200,N_7062);
and U8619 (N_8619,N_7668,N_7423);
nor U8620 (N_8620,N_7007,N_7599);
xnor U8621 (N_8621,N_7964,N_7321);
xor U8622 (N_8622,N_7886,N_7506);
and U8623 (N_8623,N_7690,N_7074);
nor U8624 (N_8624,N_7692,N_7465);
nor U8625 (N_8625,N_7860,N_7842);
or U8626 (N_8626,N_7365,N_7325);
nand U8627 (N_8627,N_7305,N_7470);
or U8628 (N_8628,N_7286,N_7842);
or U8629 (N_8629,N_7693,N_7750);
or U8630 (N_8630,N_7493,N_7983);
and U8631 (N_8631,N_7773,N_7170);
and U8632 (N_8632,N_7866,N_7174);
xnor U8633 (N_8633,N_7107,N_7458);
and U8634 (N_8634,N_7492,N_7442);
or U8635 (N_8635,N_7404,N_7080);
and U8636 (N_8636,N_7461,N_7222);
or U8637 (N_8637,N_7793,N_7346);
or U8638 (N_8638,N_7187,N_7174);
nand U8639 (N_8639,N_7968,N_7672);
xor U8640 (N_8640,N_7781,N_7257);
and U8641 (N_8641,N_7101,N_7638);
or U8642 (N_8642,N_7520,N_7746);
xnor U8643 (N_8643,N_7160,N_7747);
nor U8644 (N_8644,N_7214,N_7010);
or U8645 (N_8645,N_7697,N_7206);
xnor U8646 (N_8646,N_7212,N_7739);
nor U8647 (N_8647,N_7060,N_7313);
or U8648 (N_8648,N_7355,N_7036);
nor U8649 (N_8649,N_7336,N_7369);
and U8650 (N_8650,N_7231,N_7254);
and U8651 (N_8651,N_7232,N_7675);
nor U8652 (N_8652,N_7026,N_7195);
and U8653 (N_8653,N_7690,N_7794);
nand U8654 (N_8654,N_7073,N_7476);
xnor U8655 (N_8655,N_7509,N_7823);
nor U8656 (N_8656,N_7196,N_7730);
xnor U8657 (N_8657,N_7070,N_7999);
or U8658 (N_8658,N_7932,N_7750);
or U8659 (N_8659,N_7658,N_7064);
nor U8660 (N_8660,N_7792,N_7415);
nor U8661 (N_8661,N_7613,N_7295);
xor U8662 (N_8662,N_7266,N_7503);
nand U8663 (N_8663,N_7028,N_7653);
nor U8664 (N_8664,N_7916,N_7933);
and U8665 (N_8665,N_7942,N_7356);
and U8666 (N_8666,N_7823,N_7964);
and U8667 (N_8667,N_7600,N_7521);
nand U8668 (N_8668,N_7929,N_7233);
and U8669 (N_8669,N_7324,N_7243);
and U8670 (N_8670,N_7926,N_7496);
or U8671 (N_8671,N_7697,N_7608);
nand U8672 (N_8672,N_7742,N_7552);
nand U8673 (N_8673,N_7350,N_7409);
xor U8674 (N_8674,N_7395,N_7053);
nand U8675 (N_8675,N_7065,N_7700);
nand U8676 (N_8676,N_7008,N_7579);
and U8677 (N_8677,N_7455,N_7104);
and U8678 (N_8678,N_7132,N_7749);
or U8679 (N_8679,N_7057,N_7390);
and U8680 (N_8680,N_7961,N_7832);
nand U8681 (N_8681,N_7340,N_7615);
nand U8682 (N_8682,N_7156,N_7402);
nor U8683 (N_8683,N_7865,N_7489);
nand U8684 (N_8684,N_7366,N_7045);
nand U8685 (N_8685,N_7494,N_7872);
or U8686 (N_8686,N_7050,N_7868);
xnor U8687 (N_8687,N_7802,N_7254);
or U8688 (N_8688,N_7053,N_7665);
nor U8689 (N_8689,N_7580,N_7652);
xnor U8690 (N_8690,N_7823,N_7034);
nand U8691 (N_8691,N_7303,N_7635);
and U8692 (N_8692,N_7408,N_7511);
xor U8693 (N_8693,N_7572,N_7788);
and U8694 (N_8694,N_7975,N_7621);
and U8695 (N_8695,N_7596,N_7430);
or U8696 (N_8696,N_7906,N_7582);
or U8697 (N_8697,N_7911,N_7310);
nor U8698 (N_8698,N_7564,N_7718);
nor U8699 (N_8699,N_7133,N_7050);
xor U8700 (N_8700,N_7443,N_7437);
nor U8701 (N_8701,N_7503,N_7629);
nand U8702 (N_8702,N_7545,N_7620);
nor U8703 (N_8703,N_7383,N_7767);
nor U8704 (N_8704,N_7195,N_7329);
xor U8705 (N_8705,N_7598,N_7671);
nor U8706 (N_8706,N_7445,N_7682);
nand U8707 (N_8707,N_7677,N_7226);
or U8708 (N_8708,N_7153,N_7776);
or U8709 (N_8709,N_7991,N_7539);
nor U8710 (N_8710,N_7728,N_7647);
nand U8711 (N_8711,N_7010,N_7340);
or U8712 (N_8712,N_7405,N_7940);
or U8713 (N_8713,N_7679,N_7935);
and U8714 (N_8714,N_7945,N_7540);
or U8715 (N_8715,N_7982,N_7306);
and U8716 (N_8716,N_7510,N_7952);
xnor U8717 (N_8717,N_7166,N_7501);
xor U8718 (N_8718,N_7940,N_7034);
nor U8719 (N_8719,N_7398,N_7967);
nand U8720 (N_8720,N_7531,N_7376);
and U8721 (N_8721,N_7360,N_7772);
nor U8722 (N_8722,N_7589,N_7547);
xnor U8723 (N_8723,N_7990,N_7678);
and U8724 (N_8724,N_7910,N_7933);
and U8725 (N_8725,N_7996,N_7678);
or U8726 (N_8726,N_7120,N_7594);
nand U8727 (N_8727,N_7386,N_7933);
nor U8728 (N_8728,N_7077,N_7976);
nand U8729 (N_8729,N_7280,N_7996);
xor U8730 (N_8730,N_7541,N_7976);
nor U8731 (N_8731,N_7107,N_7124);
or U8732 (N_8732,N_7701,N_7358);
or U8733 (N_8733,N_7757,N_7166);
nor U8734 (N_8734,N_7974,N_7765);
and U8735 (N_8735,N_7042,N_7394);
xor U8736 (N_8736,N_7680,N_7987);
xor U8737 (N_8737,N_7198,N_7486);
nor U8738 (N_8738,N_7710,N_7492);
nand U8739 (N_8739,N_7878,N_7743);
nand U8740 (N_8740,N_7366,N_7061);
and U8741 (N_8741,N_7039,N_7197);
nor U8742 (N_8742,N_7299,N_7274);
nor U8743 (N_8743,N_7035,N_7212);
nand U8744 (N_8744,N_7286,N_7765);
nor U8745 (N_8745,N_7162,N_7176);
or U8746 (N_8746,N_7281,N_7480);
nor U8747 (N_8747,N_7391,N_7500);
nand U8748 (N_8748,N_7405,N_7503);
nand U8749 (N_8749,N_7971,N_7747);
xnor U8750 (N_8750,N_7771,N_7238);
nand U8751 (N_8751,N_7936,N_7233);
nand U8752 (N_8752,N_7833,N_7529);
and U8753 (N_8753,N_7286,N_7148);
or U8754 (N_8754,N_7518,N_7553);
xor U8755 (N_8755,N_7223,N_7570);
nor U8756 (N_8756,N_7482,N_7392);
nand U8757 (N_8757,N_7479,N_7916);
and U8758 (N_8758,N_7396,N_7726);
xnor U8759 (N_8759,N_7973,N_7513);
nand U8760 (N_8760,N_7344,N_7014);
or U8761 (N_8761,N_7887,N_7203);
and U8762 (N_8762,N_7944,N_7765);
or U8763 (N_8763,N_7798,N_7544);
nor U8764 (N_8764,N_7651,N_7012);
and U8765 (N_8765,N_7350,N_7204);
nor U8766 (N_8766,N_7647,N_7220);
or U8767 (N_8767,N_7261,N_7580);
nor U8768 (N_8768,N_7885,N_7013);
and U8769 (N_8769,N_7669,N_7141);
or U8770 (N_8770,N_7242,N_7836);
and U8771 (N_8771,N_7927,N_7920);
and U8772 (N_8772,N_7650,N_7442);
xor U8773 (N_8773,N_7378,N_7944);
nand U8774 (N_8774,N_7293,N_7635);
and U8775 (N_8775,N_7494,N_7107);
nor U8776 (N_8776,N_7070,N_7515);
or U8777 (N_8777,N_7069,N_7830);
xor U8778 (N_8778,N_7123,N_7411);
nor U8779 (N_8779,N_7559,N_7004);
or U8780 (N_8780,N_7359,N_7719);
nand U8781 (N_8781,N_7409,N_7043);
nor U8782 (N_8782,N_7521,N_7524);
nand U8783 (N_8783,N_7535,N_7649);
xor U8784 (N_8784,N_7128,N_7408);
nor U8785 (N_8785,N_7278,N_7127);
xnor U8786 (N_8786,N_7801,N_7383);
xor U8787 (N_8787,N_7265,N_7314);
nand U8788 (N_8788,N_7172,N_7938);
nand U8789 (N_8789,N_7124,N_7283);
and U8790 (N_8790,N_7473,N_7057);
or U8791 (N_8791,N_7356,N_7310);
nor U8792 (N_8792,N_7941,N_7806);
nand U8793 (N_8793,N_7036,N_7109);
xnor U8794 (N_8794,N_7749,N_7850);
and U8795 (N_8795,N_7084,N_7335);
and U8796 (N_8796,N_7644,N_7541);
xnor U8797 (N_8797,N_7127,N_7432);
xnor U8798 (N_8798,N_7946,N_7295);
or U8799 (N_8799,N_7285,N_7759);
xor U8800 (N_8800,N_7093,N_7450);
or U8801 (N_8801,N_7952,N_7552);
nor U8802 (N_8802,N_7845,N_7897);
or U8803 (N_8803,N_7520,N_7446);
or U8804 (N_8804,N_7846,N_7987);
nand U8805 (N_8805,N_7882,N_7169);
and U8806 (N_8806,N_7742,N_7856);
xnor U8807 (N_8807,N_7561,N_7614);
xnor U8808 (N_8808,N_7585,N_7401);
xor U8809 (N_8809,N_7336,N_7471);
nor U8810 (N_8810,N_7768,N_7196);
nor U8811 (N_8811,N_7928,N_7921);
nand U8812 (N_8812,N_7094,N_7314);
or U8813 (N_8813,N_7268,N_7230);
nor U8814 (N_8814,N_7019,N_7899);
nand U8815 (N_8815,N_7455,N_7189);
nand U8816 (N_8816,N_7303,N_7427);
and U8817 (N_8817,N_7522,N_7966);
or U8818 (N_8818,N_7713,N_7009);
and U8819 (N_8819,N_7917,N_7265);
xor U8820 (N_8820,N_7235,N_7626);
nand U8821 (N_8821,N_7043,N_7153);
and U8822 (N_8822,N_7167,N_7594);
or U8823 (N_8823,N_7468,N_7161);
nand U8824 (N_8824,N_7592,N_7237);
nor U8825 (N_8825,N_7193,N_7825);
nor U8826 (N_8826,N_7923,N_7936);
nor U8827 (N_8827,N_7097,N_7181);
or U8828 (N_8828,N_7524,N_7357);
xnor U8829 (N_8829,N_7436,N_7117);
xor U8830 (N_8830,N_7616,N_7492);
and U8831 (N_8831,N_7385,N_7534);
nor U8832 (N_8832,N_7309,N_7172);
nand U8833 (N_8833,N_7098,N_7070);
nor U8834 (N_8834,N_7449,N_7948);
xnor U8835 (N_8835,N_7831,N_7499);
nor U8836 (N_8836,N_7747,N_7646);
xor U8837 (N_8837,N_7620,N_7328);
or U8838 (N_8838,N_7624,N_7463);
nand U8839 (N_8839,N_7850,N_7741);
and U8840 (N_8840,N_7406,N_7479);
nor U8841 (N_8841,N_7103,N_7489);
nor U8842 (N_8842,N_7199,N_7159);
or U8843 (N_8843,N_7022,N_7056);
or U8844 (N_8844,N_7046,N_7572);
and U8845 (N_8845,N_7753,N_7377);
nor U8846 (N_8846,N_7369,N_7691);
xor U8847 (N_8847,N_7545,N_7380);
xnor U8848 (N_8848,N_7364,N_7281);
nand U8849 (N_8849,N_7639,N_7288);
and U8850 (N_8850,N_7937,N_7144);
or U8851 (N_8851,N_7025,N_7824);
xnor U8852 (N_8852,N_7371,N_7713);
xnor U8853 (N_8853,N_7408,N_7281);
xnor U8854 (N_8854,N_7504,N_7748);
xnor U8855 (N_8855,N_7196,N_7908);
xor U8856 (N_8856,N_7939,N_7401);
nor U8857 (N_8857,N_7064,N_7750);
or U8858 (N_8858,N_7255,N_7164);
nand U8859 (N_8859,N_7968,N_7893);
or U8860 (N_8860,N_7100,N_7349);
nor U8861 (N_8861,N_7824,N_7947);
or U8862 (N_8862,N_7833,N_7387);
nor U8863 (N_8863,N_7764,N_7754);
or U8864 (N_8864,N_7985,N_7148);
xor U8865 (N_8865,N_7866,N_7897);
or U8866 (N_8866,N_7855,N_7064);
and U8867 (N_8867,N_7477,N_7439);
nor U8868 (N_8868,N_7959,N_7975);
or U8869 (N_8869,N_7810,N_7873);
nand U8870 (N_8870,N_7525,N_7493);
nor U8871 (N_8871,N_7379,N_7502);
and U8872 (N_8872,N_7413,N_7155);
xor U8873 (N_8873,N_7336,N_7995);
and U8874 (N_8874,N_7741,N_7371);
and U8875 (N_8875,N_7922,N_7076);
or U8876 (N_8876,N_7973,N_7357);
nor U8877 (N_8877,N_7392,N_7235);
and U8878 (N_8878,N_7326,N_7401);
and U8879 (N_8879,N_7460,N_7215);
or U8880 (N_8880,N_7642,N_7594);
and U8881 (N_8881,N_7299,N_7042);
and U8882 (N_8882,N_7084,N_7058);
nand U8883 (N_8883,N_7176,N_7424);
xnor U8884 (N_8884,N_7025,N_7931);
and U8885 (N_8885,N_7934,N_7127);
xor U8886 (N_8886,N_7064,N_7603);
xor U8887 (N_8887,N_7819,N_7537);
or U8888 (N_8888,N_7743,N_7031);
nand U8889 (N_8889,N_7702,N_7874);
or U8890 (N_8890,N_7352,N_7692);
nand U8891 (N_8891,N_7181,N_7568);
and U8892 (N_8892,N_7432,N_7633);
and U8893 (N_8893,N_7579,N_7243);
or U8894 (N_8894,N_7834,N_7238);
and U8895 (N_8895,N_7937,N_7406);
or U8896 (N_8896,N_7560,N_7126);
nor U8897 (N_8897,N_7763,N_7397);
or U8898 (N_8898,N_7660,N_7115);
xnor U8899 (N_8899,N_7580,N_7387);
or U8900 (N_8900,N_7948,N_7261);
or U8901 (N_8901,N_7607,N_7488);
or U8902 (N_8902,N_7149,N_7811);
xnor U8903 (N_8903,N_7683,N_7512);
or U8904 (N_8904,N_7398,N_7056);
or U8905 (N_8905,N_7014,N_7083);
and U8906 (N_8906,N_7560,N_7941);
nand U8907 (N_8907,N_7268,N_7163);
xor U8908 (N_8908,N_7379,N_7275);
or U8909 (N_8909,N_7734,N_7356);
nor U8910 (N_8910,N_7354,N_7586);
and U8911 (N_8911,N_7196,N_7794);
xor U8912 (N_8912,N_7154,N_7382);
and U8913 (N_8913,N_7408,N_7118);
nand U8914 (N_8914,N_7673,N_7320);
nor U8915 (N_8915,N_7805,N_7114);
xnor U8916 (N_8916,N_7336,N_7862);
or U8917 (N_8917,N_7903,N_7061);
or U8918 (N_8918,N_7905,N_7832);
nand U8919 (N_8919,N_7419,N_7820);
or U8920 (N_8920,N_7523,N_7201);
or U8921 (N_8921,N_7025,N_7160);
xor U8922 (N_8922,N_7274,N_7028);
nand U8923 (N_8923,N_7677,N_7369);
and U8924 (N_8924,N_7758,N_7705);
and U8925 (N_8925,N_7365,N_7928);
xor U8926 (N_8926,N_7536,N_7861);
and U8927 (N_8927,N_7643,N_7868);
nand U8928 (N_8928,N_7364,N_7269);
and U8929 (N_8929,N_7559,N_7877);
and U8930 (N_8930,N_7376,N_7286);
and U8931 (N_8931,N_7623,N_7507);
nor U8932 (N_8932,N_7157,N_7080);
nand U8933 (N_8933,N_7120,N_7295);
xnor U8934 (N_8934,N_7846,N_7315);
and U8935 (N_8935,N_7800,N_7293);
nor U8936 (N_8936,N_7641,N_7775);
or U8937 (N_8937,N_7092,N_7480);
nand U8938 (N_8938,N_7971,N_7486);
xor U8939 (N_8939,N_7675,N_7352);
nand U8940 (N_8940,N_7278,N_7168);
nand U8941 (N_8941,N_7104,N_7604);
nor U8942 (N_8942,N_7306,N_7925);
nor U8943 (N_8943,N_7274,N_7752);
xnor U8944 (N_8944,N_7595,N_7702);
nand U8945 (N_8945,N_7246,N_7569);
and U8946 (N_8946,N_7254,N_7945);
or U8947 (N_8947,N_7129,N_7092);
nand U8948 (N_8948,N_7858,N_7161);
xnor U8949 (N_8949,N_7208,N_7052);
xor U8950 (N_8950,N_7204,N_7824);
nor U8951 (N_8951,N_7949,N_7452);
and U8952 (N_8952,N_7485,N_7344);
xor U8953 (N_8953,N_7750,N_7362);
xnor U8954 (N_8954,N_7964,N_7623);
nor U8955 (N_8955,N_7413,N_7141);
xor U8956 (N_8956,N_7462,N_7561);
nand U8957 (N_8957,N_7524,N_7721);
and U8958 (N_8958,N_7205,N_7993);
xnor U8959 (N_8959,N_7197,N_7733);
nor U8960 (N_8960,N_7748,N_7580);
xor U8961 (N_8961,N_7426,N_7294);
nor U8962 (N_8962,N_7238,N_7005);
and U8963 (N_8963,N_7351,N_7432);
nand U8964 (N_8964,N_7519,N_7791);
and U8965 (N_8965,N_7409,N_7222);
nand U8966 (N_8966,N_7800,N_7430);
or U8967 (N_8967,N_7129,N_7627);
and U8968 (N_8968,N_7936,N_7822);
nor U8969 (N_8969,N_7965,N_7916);
nand U8970 (N_8970,N_7263,N_7326);
xnor U8971 (N_8971,N_7835,N_7915);
nand U8972 (N_8972,N_7222,N_7451);
or U8973 (N_8973,N_7671,N_7559);
or U8974 (N_8974,N_7719,N_7421);
and U8975 (N_8975,N_7750,N_7394);
nor U8976 (N_8976,N_7710,N_7361);
nor U8977 (N_8977,N_7284,N_7160);
nand U8978 (N_8978,N_7620,N_7430);
or U8979 (N_8979,N_7095,N_7777);
and U8980 (N_8980,N_7996,N_7951);
or U8981 (N_8981,N_7609,N_7109);
or U8982 (N_8982,N_7839,N_7100);
nor U8983 (N_8983,N_7849,N_7725);
nor U8984 (N_8984,N_7277,N_7312);
nor U8985 (N_8985,N_7403,N_7925);
nor U8986 (N_8986,N_7519,N_7479);
nor U8987 (N_8987,N_7600,N_7482);
and U8988 (N_8988,N_7002,N_7569);
nor U8989 (N_8989,N_7248,N_7371);
nor U8990 (N_8990,N_7125,N_7621);
xnor U8991 (N_8991,N_7359,N_7311);
xor U8992 (N_8992,N_7861,N_7411);
nor U8993 (N_8993,N_7486,N_7383);
nand U8994 (N_8994,N_7054,N_7997);
nand U8995 (N_8995,N_7990,N_7645);
or U8996 (N_8996,N_7801,N_7723);
nor U8997 (N_8997,N_7238,N_7251);
nand U8998 (N_8998,N_7448,N_7184);
and U8999 (N_8999,N_7695,N_7523);
or U9000 (N_9000,N_8449,N_8646);
or U9001 (N_9001,N_8340,N_8565);
or U9002 (N_9002,N_8009,N_8768);
xor U9003 (N_9003,N_8307,N_8226);
and U9004 (N_9004,N_8848,N_8200);
nor U9005 (N_9005,N_8096,N_8130);
and U9006 (N_9006,N_8358,N_8855);
and U9007 (N_9007,N_8338,N_8567);
or U9008 (N_9008,N_8081,N_8936);
nand U9009 (N_9009,N_8209,N_8949);
nor U9010 (N_9010,N_8968,N_8624);
nand U9011 (N_9011,N_8765,N_8259);
and U9012 (N_9012,N_8019,N_8817);
and U9013 (N_9013,N_8020,N_8759);
nand U9014 (N_9014,N_8502,N_8649);
or U9015 (N_9015,N_8382,N_8676);
xor U9016 (N_9016,N_8432,N_8182);
and U9017 (N_9017,N_8147,N_8870);
nor U9018 (N_9018,N_8863,N_8722);
nor U9019 (N_9019,N_8254,N_8396);
nand U9020 (N_9020,N_8906,N_8588);
nand U9021 (N_9021,N_8654,N_8472);
nand U9022 (N_9022,N_8157,N_8665);
nor U9023 (N_9023,N_8005,N_8123);
nor U9024 (N_9024,N_8711,N_8135);
and U9025 (N_9025,N_8206,N_8710);
nor U9026 (N_9026,N_8370,N_8648);
or U9027 (N_9027,N_8141,N_8046);
xnor U9028 (N_9028,N_8414,N_8947);
nor U9029 (N_9029,N_8609,N_8680);
nand U9030 (N_9030,N_8470,N_8416);
xnor U9031 (N_9031,N_8994,N_8294);
or U9032 (N_9032,N_8637,N_8023);
or U9033 (N_9033,N_8858,N_8129);
or U9034 (N_9034,N_8011,N_8308);
nor U9035 (N_9035,N_8555,N_8729);
xor U9036 (N_9036,N_8986,N_8140);
or U9037 (N_9037,N_8544,N_8539);
and U9038 (N_9038,N_8821,N_8508);
nor U9039 (N_9039,N_8709,N_8643);
xor U9040 (N_9040,N_8280,N_8439);
or U9041 (N_9041,N_8916,N_8160);
and U9042 (N_9042,N_8910,N_8530);
nor U9043 (N_9043,N_8720,N_8374);
nand U9044 (N_9044,N_8059,N_8929);
nor U9045 (N_9045,N_8301,N_8060);
nand U9046 (N_9046,N_8976,N_8049);
and U9047 (N_9047,N_8190,N_8881);
or U9048 (N_9048,N_8133,N_8660);
nand U9049 (N_9049,N_8996,N_8314);
nor U9050 (N_9050,N_8224,N_8792);
and U9051 (N_9051,N_8635,N_8510);
nor U9052 (N_9052,N_8112,N_8726);
nand U9053 (N_9053,N_8569,N_8772);
or U9054 (N_9054,N_8069,N_8550);
xor U9055 (N_9055,N_8708,N_8935);
or U9056 (N_9056,N_8311,N_8335);
nand U9057 (N_9057,N_8877,N_8867);
nand U9058 (N_9058,N_8445,N_8261);
nand U9059 (N_9059,N_8106,N_8528);
or U9060 (N_9060,N_8807,N_8953);
or U9061 (N_9061,N_8601,N_8412);
xor U9062 (N_9062,N_8698,N_8094);
and U9063 (N_9063,N_8437,N_8002);
nor U9064 (N_9064,N_8498,N_8853);
or U9065 (N_9065,N_8477,N_8557);
or U9066 (N_9066,N_8107,N_8796);
nand U9067 (N_9067,N_8885,N_8343);
nor U9068 (N_9068,N_8405,N_8869);
and U9069 (N_9069,N_8795,N_8741);
nand U9070 (N_9070,N_8578,N_8706);
nand U9071 (N_9071,N_8511,N_8850);
xnor U9072 (N_9072,N_8442,N_8605);
and U9073 (N_9073,N_8950,N_8526);
and U9074 (N_9074,N_8355,N_8989);
and U9075 (N_9075,N_8198,N_8967);
nor U9076 (N_9076,N_8612,N_8856);
or U9077 (N_9077,N_8375,N_8455);
and U9078 (N_9078,N_8043,N_8684);
and U9079 (N_9079,N_8415,N_8801);
nand U9080 (N_9080,N_8516,N_8004);
or U9081 (N_9081,N_8529,N_8840);
and U9082 (N_9082,N_8621,N_8841);
nand U9083 (N_9083,N_8017,N_8938);
nor U9084 (N_9084,N_8583,N_8608);
or U9085 (N_9085,N_8816,N_8234);
and U9086 (N_9086,N_8315,N_8580);
or U9087 (N_9087,N_8762,N_8440);
xnor U9088 (N_9088,N_8247,N_8925);
nand U9089 (N_9089,N_8667,N_8100);
xor U9090 (N_9090,N_8851,N_8479);
xnor U9091 (N_9091,N_8407,N_8255);
and U9092 (N_9092,N_8427,N_8907);
and U9093 (N_9093,N_8101,N_8551);
or U9094 (N_9094,N_8393,N_8592);
nand U9095 (N_9095,N_8776,N_8153);
nor U9096 (N_9096,N_8118,N_8073);
nand U9097 (N_9097,N_8493,N_8217);
nand U9098 (N_9098,N_8634,N_8724);
nand U9099 (N_9099,N_8451,N_8657);
nand U9100 (N_9100,N_8804,N_8620);
nand U9101 (N_9101,N_8482,N_8156);
nand U9102 (N_9102,N_8626,N_8097);
nand U9103 (N_9103,N_8878,N_8290);
and U9104 (N_9104,N_8337,N_8025);
and U9105 (N_9105,N_8227,N_8436);
and U9106 (N_9106,N_8114,N_8467);
nand U9107 (N_9107,N_8196,N_8181);
nand U9108 (N_9108,N_8973,N_8536);
and U9109 (N_9109,N_8201,N_8015);
xor U9110 (N_9110,N_8622,N_8447);
and U9111 (N_9111,N_8981,N_8653);
xnor U9112 (N_9112,N_8538,N_8235);
nor U9113 (N_9113,N_8492,N_8959);
nand U9114 (N_9114,N_8596,N_8942);
nor U9115 (N_9115,N_8347,N_8007);
xnor U9116 (N_9116,N_8572,N_8832);
and U9117 (N_9117,N_8532,N_8168);
nor U9118 (N_9118,N_8974,N_8456);
nand U9119 (N_9119,N_8363,N_8260);
nor U9120 (N_9120,N_8633,N_8194);
nor U9121 (N_9121,N_8272,N_8253);
and U9122 (N_9122,N_8589,N_8566);
or U9123 (N_9123,N_8281,N_8638);
nand U9124 (N_9124,N_8733,N_8604);
nor U9125 (N_9125,N_8798,N_8320);
xnor U9126 (N_9126,N_8429,N_8418);
and U9127 (N_9127,N_8599,N_8222);
and U9128 (N_9128,N_8831,N_8758);
nand U9129 (N_9129,N_8179,N_8509);
and U9130 (N_9130,N_8763,N_8564);
nand U9131 (N_9131,N_8948,N_8339);
nor U9132 (N_9132,N_8450,N_8186);
nand U9133 (N_9133,N_8868,N_8458);
xnor U9134 (N_9134,N_8408,N_8505);
xor U9135 (N_9135,N_8924,N_8813);
xnor U9136 (N_9136,N_8754,N_8388);
or U9137 (N_9137,N_8171,N_8242);
xor U9138 (N_9138,N_8327,N_8675);
nor U9139 (N_9139,N_8379,N_8122);
nor U9140 (N_9140,N_8812,N_8700);
nor U9141 (N_9141,N_8854,N_8735);
and U9142 (N_9142,N_8613,N_8518);
xnor U9143 (N_9143,N_8302,N_8541);
nand U9144 (N_9144,N_8045,N_8717);
nor U9145 (N_9145,N_8992,N_8494);
nand U9146 (N_9146,N_8263,N_8984);
xor U9147 (N_9147,N_8785,N_8752);
xor U9148 (N_9148,N_8083,N_8233);
xor U9149 (N_9149,N_8095,N_8677);
and U9150 (N_9150,N_8210,N_8443);
xnor U9151 (N_9151,N_8462,N_8282);
or U9152 (N_9152,N_8406,N_8425);
xor U9153 (N_9153,N_8890,N_8997);
nor U9154 (N_9154,N_8000,N_8628);
or U9155 (N_9155,N_8399,N_8092);
and U9156 (N_9156,N_8420,N_8430);
nand U9157 (N_9157,N_8842,N_8586);
or U9158 (N_9158,N_8829,N_8356);
nor U9159 (N_9159,N_8040,N_8962);
nand U9160 (N_9160,N_8471,N_8696);
and U9161 (N_9161,N_8317,N_8312);
or U9162 (N_9162,N_8299,N_8672);
or U9163 (N_9163,N_8348,N_8811);
nor U9164 (N_9164,N_8940,N_8423);
nand U9165 (N_9165,N_8287,N_8266);
nor U9166 (N_9166,N_8360,N_8614);
nor U9167 (N_9167,N_8006,N_8740);
and U9168 (N_9168,N_8678,N_8264);
nor U9169 (N_9169,N_8610,N_8435);
and U9170 (N_9170,N_8286,N_8368);
xnor U9171 (N_9171,N_8714,N_8283);
nand U9172 (N_9172,N_8333,N_8563);
xnor U9173 (N_9173,N_8945,N_8731);
xor U9174 (N_9174,N_8035,N_8359);
nand U9175 (N_9175,N_8386,N_8051);
nor U9176 (N_9176,N_8262,N_8775);
and U9177 (N_9177,N_8365,N_8350);
nor U9178 (N_9178,N_8164,N_8560);
nor U9179 (N_9179,N_8229,N_8499);
and U9180 (N_9180,N_8380,N_8372);
nor U9181 (N_9181,N_8158,N_8076);
nand U9182 (N_9182,N_8876,N_8618);
nand U9183 (N_9183,N_8982,N_8694);
nand U9184 (N_9184,N_8595,N_8269);
xor U9185 (N_9185,N_8993,N_8930);
nor U9186 (N_9186,N_8826,N_8738);
xor U9187 (N_9187,N_8279,N_8513);
nor U9188 (N_9188,N_8244,N_8884);
nor U9189 (N_9189,N_8561,N_8417);
and U9190 (N_9190,N_8579,N_8783);
or U9191 (N_9191,N_8422,N_8943);
xor U9192 (N_9192,N_8914,N_8237);
nand U9193 (N_9193,N_8652,N_8822);
xor U9194 (N_9194,N_8901,N_8491);
nand U9195 (N_9195,N_8354,N_8662);
nand U9196 (N_9196,N_8468,N_8611);
or U9197 (N_9197,N_8788,N_8245);
nor U9198 (N_9198,N_8008,N_8593);
nor U9199 (N_9199,N_8362,N_8463);
nor U9200 (N_9200,N_8641,N_8223);
xor U9201 (N_9201,N_8366,N_8514);
and U9202 (N_9202,N_8297,N_8220);
nand U9203 (N_9203,N_8138,N_8166);
or U9204 (N_9204,N_8257,N_8747);
and U9205 (N_9205,N_8137,N_8072);
nor U9206 (N_9206,N_8871,N_8161);
xnor U9207 (N_9207,N_8378,N_8033);
xnor U9208 (N_9208,N_8584,N_8679);
and U9209 (N_9209,N_8815,N_8324);
nand U9210 (N_9210,N_8705,N_8212);
nor U9211 (N_9211,N_8545,N_8438);
nand U9212 (N_9212,N_8799,N_8170);
nor U9213 (N_9213,N_8629,N_8316);
nor U9214 (N_9214,N_8861,N_8689);
xor U9215 (N_9215,N_8488,N_8903);
nor U9216 (N_9216,N_8787,N_8603);
nor U9217 (N_9217,N_8003,N_8766);
and U9218 (N_9218,N_8411,N_8904);
and U9219 (N_9219,N_8117,N_8955);
xnor U9220 (N_9220,N_8873,N_8784);
nand U9221 (N_9221,N_8460,N_8484);
and U9222 (N_9222,N_8902,N_8547);
and U9223 (N_9223,N_8666,N_8797);
or U9224 (N_9224,N_8699,N_8573);
nor U9225 (N_9225,N_8042,N_8808);
or U9226 (N_9226,N_8975,N_8805);
and U9227 (N_9227,N_8300,N_8330);
nand U9228 (N_9228,N_8295,N_8941);
nor U9229 (N_9229,N_8977,N_8207);
xor U9230 (N_9230,N_8139,N_8650);
or U9231 (N_9231,N_8401,N_8998);
or U9232 (N_9232,N_8068,N_8178);
nor U9233 (N_9233,N_8814,N_8755);
nand U9234 (N_9234,N_8892,N_8037);
nand U9235 (N_9235,N_8748,N_8630);
nor U9236 (N_9236,N_8431,N_8148);
nor U9237 (N_9237,N_8497,N_8719);
or U9238 (N_9238,N_8022,N_8651);
nor U9239 (N_9239,N_8419,N_8453);
and U9240 (N_9240,N_8669,N_8865);
or U9241 (N_9241,N_8154,N_8256);
xnor U9242 (N_9242,N_8697,N_8964);
nand U9243 (N_9243,N_8506,N_8732);
nand U9244 (N_9244,N_8014,N_8127);
or U9245 (N_9245,N_8376,N_8329);
nor U9246 (N_9246,N_8512,N_8857);
and U9247 (N_9247,N_8520,N_8185);
and U9248 (N_9248,N_8001,N_8552);
nand U9249 (N_9249,N_8079,N_8152);
and U9250 (N_9250,N_8957,N_8639);
nand U9251 (N_9251,N_8318,N_8522);
and U9252 (N_9252,N_8052,N_8028);
and U9253 (N_9253,N_8131,N_8562);
xor U9254 (N_9254,N_8761,N_8958);
or U9255 (N_9255,N_8844,N_8369);
nor U9256 (N_9256,N_8760,N_8278);
or U9257 (N_9257,N_8024,N_8970);
nor U9258 (N_9258,N_8771,N_8575);
and U9259 (N_9259,N_8288,N_8144);
nor U9260 (N_9260,N_8543,N_8021);
xor U9261 (N_9261,N_8485,N_8238);
nor U9262 (N_9262,N_8012,N_8277);
nand U9263 (N_9263,N_8995,N_8062);
and U9264 (N_9264,N_8361,N_8742);
or U9265 (N_9265,N_8010,N_8803);
xnor U9266 (N_9266,N_8134,N_8313);
xnor U9267 (N_9267,N_8167,N_8728);
xnor U9268 (N_9268,N_8837,N_8751);
xnor U9269 (N_9269,N_8197,N_8128);
nor U9270 (N_9270,N_8917,N_8250);
xor U9271 (N_9271,N_8559,N_8843);
xnor U9272 (N_9272,N_8847,N_8725);
and U9273 (N_9273,N_8839,N_8570);
or U9274 (N_9274,N_8270,N_8132);
xor U9275 (N_9275,N_8424,N_8616);
or U9276 (N_9276,N_8746,N_8954);
and U9277 (N_9277,N_8764,N_8099);
nor U9278 (N_9278,N_8490,N_8218);
and U9279 (N_9279,N_8480,N_8331);
or U9280 (N_9280,N_8632,N_8057);
and U9281 (N_9281,N_8743,N_8126);
or U9282 (N_9282,N_8923,N_8860);
or U9283 (N_9283,N_8888,N_8600);
nor U9284 (N_9284,N_8172,N_8292);
xnor U9285 (N_9285,N_8251,N_8150);
nor U9286 (N_9286,N_8880,N_8809);
nor U9287 (N_9287,N_8875,N_8483);
nand U9288 (N_9288,N_8304,N_8770);
nand U9289 (N_9289,N_8585,N_8554);
nor U9290 (N_9290,N_8574,N_8428);
nor U9291 (N_9291,N_8125,N_8756);
nor U9292 (N_9292,N_8546,N_8531);
xnor U9293 (N_9293,N_8750,N_8221);
and U9294 (N_9294,N_8819,N_8602);
and U9295 (N_9295,N_8064,N_8162);
xnor U9296 (N_9296,N_8778,N_8031);
and U9297 (N_9297,N_8535,N_8736);
nor U9298 (N_9298,N_8219,N_8695);
and U9299 (N_9299,N_8400,N_8188);
nand U9300 (N_9300,N_8882,N_8800);
nor U9301 (N_9301,N_8478,N_8791);
and U9302 (N_9302,N_8061,N_8874);
nor U9303 (N_9303,N_8521,N_8619);
xnor U9304 (N_9304,N_8155,N_8659);
nand U9305 (N_9305,N_8136,N_8457);
nand U9306 (N_9306,N_8500,N_8905);
and U9307 (N_9307,N_8204,N_8988);
or U9308 (N_9308,N_8745,N_8284);
nor U9309 (N_9309,N_8780,N_8845);
nand U9310 (N_9310,N_8786,N_8448);
and U9311 (N_9311,N_8961,N_8631);
xnor U9312 (N_9312,N_8030,N_8063);
xnor U9313 (N_9313,N_8991,N_8103);
or U9314 (N_9314,N_8390,N_8937);
xor U9315 (N_9315,N_8149,N_8034);
nor U9316 (N_9316,N_8607,N_8305);
nor U9317 (N_9317,N_8645,N_8082);
and U9318 (N_9318,N_8757,N_8987);
or U9319 (N_9319,N_8712,N_8656);
or U9320 (N_9320,N_8922,N_8474);
or U9321 (N_9321,N_8075,N_8838);
nor U9322 (N_9322,N_8306,N_8960);
or U9323 (N_9323,N_8644,N_8897);
nand U9324 (N_9324,N_8018,N_8887);
or U9325 (N_9325,N_8367,N_8625);
nor U9326 (N_9326,N_8093,N_8124);
xor U9327 (N_9327,N_8215,N_8091);
or U9328 (N_9328,N_8661,N_8927);
xor U9329 (N_9329,N_8252,N_8965);
nand U9330 (N_9330,N_8794,N_8055);
nand U9331 (N_9331,N_8990,N_8029);
or U9332 (N_9332,N_8926,N_8828);
or U9333 (N_9333,N_8184,N_8793);
or U9334 (N_9334,N_8704,N_8243);
or U9335 (N_9335,N_8016,N_8920);
xor U9336 (N_9336,N_8446,N_8169);
nand U9337 (N_9337,N_8351,N_8703);
nor U9338 (N_9338,N_8322,N_8032);
and U9339 (N_9339,N_8323,N_8889);
nand U9340 (N_9340,N_8963,N_8663);
or U9341 (N_9341,N_8265,N_8473);
nand U9342 (N_9342,N_8782,N_8334);
nor U9343 (N_9343,N_8192,N_8886);
nand U9344 (N_9344,N_8108,N_8402);
nor U9345 (N_9345,N_8674,N_8895);
or U9346 (N_9346,N_8341,N_8971);
and U9347 (N_9347,N_8146,N_8345);
and U9348 (N_9348,N_8387,N_8391);
xor U9349 (N_9349,N_8193,N_8026);
nor U9350 (N_9350,N_8504,N_8199);
xnor U9351 (N_9351,N_8598,N_8866);
or U9352 (N_9352,N_8836,N_8972);
xnor U9353 (N_9353,N_8395,N_8534);
nor U9354 (N_9354,N_8214,N_8248);
nor U9355 (N_9355,N_8298,N_8342);
or U9356 (N_9356,N_8163,N_8978);
and U9357 (N_9357,N_8979,N_8558);
xnor U9358 (N_9358,N_8085,N_8475);
nand U9359 (N_9359,N_8145,N_8683);
nand U9360 (N_9360,N_8883,N_8409);
and U9361 (N_9361,N_8383,N_8228);
nor U9362 (N_9362,N_8056,N_8896);
nor U9363 (N_9363,N_8187,N_8501);
or U9364 (N_9364,N_8357,N_8293);
nand U9365 (N_9365,N_8273,N_8693);
nand U9366 (N_9366,N_8173,N_8525);
or U9367 (N_9367,N_8549,N_8615);
and U9368 (N_9368,N_8670,N_8274);
nor U9369 (N_9369,N_8344,N_8258);
xnor U9370 (N_9370,N_8090,N_8377);
or U9371 (N_9371,N_8176,N_8332);
and U9372 (N_9372,N_8495,N_8898);
nand U9373 (N_9373,N_8673,N_8753);
nor U9374 (N_9374,N_8980,N_8681);
nand U9375 (N_9375,N_8113,N_8918);
or U9376 (N_9376,N_8859,N_8737);
nor U9377 (N_9377,N_8054,N_8789);
nand U9378 (N_9378,N_8951,N_8328);
and U9379 (N_9379,N_8452,N_8921);
and U9380 (N_9380,N_8180,N_8594);
xor U9381 (N_9381,N_8834,N_8053);
xor U9382 (N_9382,N_8110,N_8668);
nor U9383 (N_9383,N_8734,N_8321);
nand U9384 (N_9384,N_8098,N_8285);
or U9385 (N_9385,N_8050,N_8537);
nor U9386 (N_9386,N_8739,N_8267);
and U9387 (N_9387,N_8749,N_8213);
xnor U9388 (N_9388,N_8909,N_8486);
nor U9389 (N_9389,N_8105,N_8894);
xnor U9390 (N_9390,N_8174,N_8582);
nor U9391 (N_9391,N_8088,N_8825);
and U9392 (N_9392,N_8540,N_8403);
xor U9393 (N_9393,N_8202,N_8296);
xor U9394 (N_9394,N_8489,N_8275);
nand U9395 (N_9395,N_8820,N_8730);
and U9396 (N_9396,N_8769,N_8177);
xor U9397 (N_9397,N_8142,N_8086);
and U9398 (N_9398,N_8038,N_8524);
xnor U9399 (N_9399,N_8392,N_8115);
nor U9400 (N_9400,N_8225,N_8928);
nand U9401 (N_9401,N_8381,N_8818);
nor U9402 (N_9402,N_8398,N_8827);
nand U9403 (N_9403,N_8835,N_8241);
or U9404 (N_9404,N_8476,N_8915);
or U9405 (N_9405,N_8617,N_8919);
xnor U9406 (N_9406,N_8433,N_8542);
or U9407 (N_9407,N_8872,N_8627);
and U9408 (N_9408,N_8325,N_8686);
nor U9409 (N_9409,N_8189,N_8833);
xnor U9410 (N_9410,N_8774,N_8671);
and U9411 (N_9411,N_8577,N_8707);
xnor U9412 (N_9412,N_8240,N_8533);
or U9413 (N_9413,N_8077,N_8371);
xor U9414 (N_9414,N_8773,N_8688);
or U9415 (N_9415,N_8385,N_8908);
or U9416 (N_9416,N_8718,N_8946);
nor U9417 (N_9417,N_8121,N_8727);
nand U9418 (N_9418,N_8806,N_8952);
xor U9419 (N_9419,N_8421,N_8087);
xnor U9420 (N_9420,N_8568,N_8464);
nor U9421 (N_9421,N_8310,N_8336);
or U9422 (N_9422,N_8623,N_8576);
nand U9423 (N_9423,N_8956,N_8647);
nor U9424 (N_9424,N_8692,N_8891);
nand U9425 (N_9425,N_8723,N_8899);
nor U9426 (N_9426,N_8426,N_8268);
or U9427 (N_9427,N_8319,N_8900);
nor U9428 (N_9428,N_8830,N_8058);
or U9429 (N_9429,N_8587,N_8879);
xor U9430 (N_9430,N_8303,N_8503);
and U9431 (N_9431,N_8519,N_8346);
xor U9432 (N_9432,N_8159,N_8823);
xnor U9433 (N_9433,N_8461,N_8389);
xnor U9434 (N_9434,N_8691,N_8713);
and U9435 (N_9435,N_8932,N_8353);
or U9436 (N_9436,N_8216,N_8779);
or U9437 (N_9437,N_8655,N_8271);
nand U9438 (N_9438,N_8496,N_8934);
or U9439 (N_9439,N_8893,N_8434);
or U9440 (N_9440,N_8413,N_8702);
xor U9441 (N_9441,N_8556,N_8658);
nand U9442 (N_9442,N_8039,N_8507);
or U9443 (N_9443,N_8548,N_8289);
nand U9444 (N_9444,N_8523,N_8715);
nand U9445 (N_9445,N_8701,N_8404);
or U9446 (N_9446,N_8078,N_8230);
and U9447 (N_9447,N_8767,N_8802);
and U9448 (N_9448,N_8790,N_8067);
nor U9449 (N_9449,N_8143,N_8036);
xnor U9450 (N_9450,N_8852,N_8966);
nor U9451 (N_9451,N_8203,N_8912);
xor U9452 (N_9452,N_8911,N_8664);
or U9453 (N_9453,N_8469,N_8939);
or U9454 (N_9454,N_8944,N_8211);
xnor U9455 (N_9455,N_8571,N_8102);
and U9456 (N_9456,N_8441,N_8397);
nand U9457 (N_9457,N_8089,N_8864);
or U9458 (N_9458,N_8205,N_8208);
xnor U9459 (N_9459,N_8044,N_8999);
or U9460 (N_9460,N_8373,N_8810);
or U9461 (N_9461,N_8515,N_8466);
nand U9462 (N_9462,N_8047,N_8239);
xor U9463 (N_9463,N_8175,N_8183);
or U9464 (N_9464,N_8394,N_8410);
nand U9465 (N_9465,N_8120,N_8276);
nand U9466 (N_9466,N_8597,N_8640);
xnor U9467 (N_9467,N_8459,N_8465);
xor U9468 (N_9468,N_8384,N_8236);
or U9469 (N_9469,N_8151,N_8291);
nor U9470 (N_9470,N_8985,N_8104);
nand U9471 (N_9471,N_8364,N_8682);
xor U9472 (N_9472,N_8824,N_8581);
and U9473 (N_9473,N_8191,N_8231);
and U9474 (N_9474,N_8744,N_8913);
and U9475 (N_9475,N_8349,N_8249);
and U9476 (N_9476,N_8636,N_8690);
and U9477 (N_9477,N_8111,N_8041);
or U9478 (N_9478,N_8553,N_8846);
nor U9479 (N_9479,N_8590,N_8232);
and U9480 (N_9480,N_8481,N_8080);
or U9481 (N_9481,N_8119,N_8048);
and U9482 (N_9482,N_8027,N_8074);
and U9483 (N_9483,N_8933,N_8931);
or U9484 (N_9484,N_8444,N_8721);
and U9485 (N_9485,N_8591,N_8777);
xnor U9486 (N_9486,N_8862,N_8983);
or U9487 (N_9487,N_8070,N_8109);
nand U9488 (N_9488,N_8454,N_8066);
nor U9489 (N_9489,N_8487,N_8309);
and U9490 (N_9490,N_8687,N_8165);
nor U9491 (N_9491,N_8849,N_8716);
nor U9492 (N_9492,N_8065,N_8116);
or U9493 (N_9493,N_8013,N_8517);
nor U9494 (N_9494,N_8246,N_8195);
xnor U9495 (N_9495,N_8352,N_8781);
nor U9496 (N_9496,N_8606,N_8527);
or U9497 (N_9497,N_8969,N_8326);
and U9498 (N_9498,N_8685,N_8071);
and U9499 (N_9499,N_8084,N_8642);
nand U9500 (N_9500,N_8565,N_8378);
xor U9501 (N_9501,N_8615,N_8849);
nor U9502 (N_9502,N_8728,N_8099);
nand U9503 (N_9503,N_8944,N_8378);
nand U9504 (N_9504,N_8303,N_8027);
nor U9505 (N_9505,N_8857,N_8075);
or U9506 (N_9506,N_8482,N_8827);
xor U9507 (N_9507,N_8787,N_8594);
or U9508 (N_9508,N_8020,N_8536);
or U9509 (N_9509,N_8460,N_8081);
xor U9510 (N_9510,N_8596,N_8779);
nand U9511 (N_9511,N_8484,N_8876);
nor U9512 (N_9512,N_8477,N_8168);
xnor U9513 (N_9513,N_8881,N_8874);
nor U9514 (N_9514,N_8527,N_8543);
nand U9515 (N_9515,N_8619,N_8372);
nand U9516 (N_9516,N_8875,N_8839);
nor U9517 (N_9517,N_8061,N_8081);
nand U9518 (N_9518,N_8409,N_8538);
xor U9519 (N_9519,N_8861,N_8600);
nor U9520 (N_9520,N_8872,N_8461);
nand U9521 (N_9521,N_8155,N_8000);
xnor U9522 (N_9522,N_8779,N_8435);
xnor U9523 (N_9523,N_8620,N_8946);
xnor U9524 (N_9524,N_8627,N_8801);
or U9525 (N_9525,N_8992,N_8309);
and U9526 (N_9526,N_8303,N_8853);
nand U9527 (N_9527,N_8022,N_8276);
nor U9528 (N_9528,N_8616,N_8803);
and U9529 (N_9529,N_8593,N_8878);
and U9530 (N_9530,N_8922,N_8526);
nand U9531 (N_9531,N_8510,N_8744);
or U9532 (N_9532,N_8774,N_8732);
or U9533 (N_9533,N_8997,N_8308);
xor U9534 (N_9534,N_8845,N_8346);
nand U9535 (N_9535,N_8284,N_8994);
or U9536 (N_9536,N_8090,N_8102);
and U9537 (N_9537,N_8432,N_8575);
nor U9538 (N_9538,N_8584,N_8566);
nor U9539 (N_9539,N_8734,N_8597);
and U9540 (N_9540,N_8378,N_8005);
or U9541 (N_9541,N_8842,N_8065);
nor U9542 (N_9542,N_8668,N_8760);
xor U9543 (N_9543,N_8463,N_8140);
nor U9544 (N_9544,N_8715,N_8020);
xor U9545 (N_9545,N_8675,N_8383);
nand U9546 (N_9546,N_8158,N_8869);
and U9547 (N_9547,N_8057,N_8931);
nand U9548 (N_9548,N_8534,N_8491);
or U9549 (N_9549,N_8768,N_8794);
nor U9550 (N_9550,N_8898,N_8416);
and U9551 (N_9551,N_8544,N_8029);
xor U9552 (N_9552,N_8636,N_8614);
nand U9553 (N_9553,N_8854,N_8641);
or U9554 (N_9554,N_8806,N_8390);
nor U9555 (N_9555,N_8220,N_8356);
nand U9556 (N_9556,N_8839,N_8982);
nor U9557 (N_9557,N_8972,N_8716);
and U9558 (N_9558,N_8298,N_8758);
nor U9559 (N_9559,N_8432,N_8549);
nand U9560 (N_9560,N_8086,N_8219);
and U9561 (N_9561,N_8935,N_8603);
xor U9562 (N_9562,N_8228,N_8324);
or U9563 (N_9563,N_8667,N_8479);
or U9564 (N_9564,N_8642,N_8361);
nor U9565 (N_9565,N_8656,N_8722);
and U9566 (N_9566,N_8614,N_8106);
xnor U9567 (N_9567,N_8680,N_8888);
and U9568 (N_9568,N_8597,N_8729);
or U9569 (N_9569,N_8830,N_8389);
xor U9570 (N_9570,N_8562,N_8336);
and U9571 (N_9571,N_8691,N_8890);
or U9572 (N_9572,N_8154,N_8718);
xor U9573 (N_9573,N_8559,N_8216);
or U9574 (N_9574,N_8259,N_8413);
and U9575 (N_9575,N_8612,N_8679);
nor U9576 (N_9576,N_8191,N_8823);
xor U9577 (N_9577,N_8366,N_8694);
nor U9578 (N_9578,N_8578,N_8640);
or U9579 (N_9579,N_8758,N_8163);
nor U9580 (N_9580,N_8418,N_8226);
nor U9581 (N_9581,N_8133,N_8171);
xor U9582 (N_9582,N_8795,N_8009);
nor U9583 (N_9583,N_8670,N_8542);
and U9584 (N_9584,N_8463,N_8890);
xnor U9585 (N_9585,N_8990,N_8017);
xnor U9586 (N_9586,N_8319,N_8224);
xor U9587 (N_9587,N_8121,N_8827);
and U9588 (N_9588,N_8709,N_8703);
or U9589 (N_9589,N_8902,N_8876);
xor U9590 (N_9590,N_8399,N_8494);
nor U9591 (N_9591,N_8534,N_8167);
and U9592 (N_9592,N_8757,N_8025);
nor U9593 (N_9593,N_8842,N_8246);
xor U9594 (N_9594,N_8892,N_8236);
xor U9595 (N_9595,N_8191,N_8533);
or U9596 (N_9596,N_8104,N_8377);
xnor U9597 (N_9597,N_8074,N_8929);
or U9598 (N_9598,N_8291,N_8573);
or U9599 (N_9599,N_8413,N_8101);
or U9600 (N_9600,N_8403,N_8593);
or U9601 (N_9601,N_8023,N_8828);
and U9602 (N_9602,N_8500,N_8243);
or U9603 (N_9603,N_8288,N_8638);
nor U9604 (N_9604,N_8342,N_8403);
and U9605 (N_9605,N_8805,N_8375);
or U9606 (N_9606,N_8033,N_8687);
nand U9607 (N_9607,N_8758,N_8053);
nor U9608 (N_9608,N_8595,N_8697);
nand U9609 (N_9609,N_8293,N_8059);
and U9610 (N_9610,N_8176,N_8501);
and U9611 (N_9611,N_8837,N_8530);
nor U9612 (N_9612,N_8855,N_8643);
or U9613 (N_9613,N_8652,N_8759);
xor U9614 (N_9614,N_8474,N_8428);
nand U9615 (N_9615,N_8282,N_8166);
xnor U9616 (N_9616,N_8824,N_8873);
nor U9617 (N_9617,N_8869,N_8972);
or U9618 (N_9618,N_8684,N_8121);
or U9619 (N_9619,N_8603,N_8129);
xor U9620 (N_9620,N_8322,N_8541);
and U9621 (N_9621,N_8882,N_8668);
and U9622 (N_9622,N_8510,N_8898);
xnor U9623 (N_9623,N_8842,N_8231);
and U9624 (N_9624,N_8124,N_8070);
or U9625 (N_9625,N_8214,N_8677);
and U9626 (N_9626,N_8178,N_8437);
nor U9627 (N_9627,N_8765,N_8965);
or U9628 (N_9628,N_8760,N_8877);
and U9629 (N_9629,N_8559,N_8793);
xnor U9630 (N_9630,N_8799,N_8537);
xnor U9631 (N_9631,N_8481,N_8427);
nand U9632 (N_9632,N_8337,N_8133);
nor U9633 (N_9633,N_8170,N_8841);
nor U9634 (N_9634,N_8548,N_8721);
nor U9635 (N_9635,N_8608,N_8831);
and U9636 (N_9636,N_8723,N_8634);
or U9637 (N_9637,N_8542,N_8645);
nor U9638 (N_9638,N_8096,N_8732);
nand U9639 (N_9639,N_8966,N_8783);
nor U9640 (N_9640,N_8061,N_8038);
xor U9641 (N_9641,N_8367,N_8613);
or U9642 (N_9642,N_8505,N_8652);
xnor U9643 (N_9643,N_8466,N_8465);
and U9644 (N_9644,N_8189,N_8215);
nand U9645 (N_9645,N_8632,N_8513);
or U9646 (N_9646,N_8132,N_8807);
and U9647 (N_9647,N_8877,N_8231);
or U9648 (N_9648,N_8429,N_8219);
nand U9649 (N_9649,N_8842,N_8686);
nor U9650 (N_9650,N_8667,N_8401);
xnor U9651 (N_9651,N_8875,N_8885);
nand U9652 (N_9652,N_8571,N_8700);
and U9653 (N_9653,N_8416,N_8698);
nor U9654 (N_9654,N_8441,N_8029);
nor U9655 (N_9655,N_8622,N_8875);
xnor U9656 (N_9656,N_8652,N_8720);
and U9657 (N_9657,N_8161,N_8517);
nand U9658 (N_9658,N_8277,N_8813);
or U9659 (N_9659,N_8736,N_8318);
or U9660 (N_9660,N_8369,N_8412);
and U9661 (N_9661,N_8435,N_8320);
nor U9662 (N_9662,N_8166,N_8463);
and U9663 (N_9663,N_8613,N_8293);
and U9664 (N_9664,N_8085,N_8033);
xor U9665 (N_9665,N_8659,N_8957);
and U9666 (N_9666,N_8764,N_8794);
and U9667 (N_9667,N_8434,N_8439);
nor U9668 (N_9668,N_8862,N_8545);
xor U9669 (N_9669,N_8251,N_8552);
and U9670 (N_9670,N_8870,N_8716);
and U9671 (N_9671,N_8301,N_8444);
xnor U9672 (N_9672,N_8285,N_8065);
nor U9673 (N_9673,N_8495,N_8957);
and U9674 (N_9674,N_8699,N_8373);
and U9675 (N_9675,N_8724,N_8779);
or U9676 (N_9676,N_8531,N_8656);
and U9677 (N_9677,N_8710,N_8249);
xnor U9678 (N_9678,N_8824,N_8861);
nor U9679 (N_9679,N_8223,N_8518);
nor U9680 (N_9680,N_8991,N_8625);
nand U9681 (N_9681,N_8951,N_8373);
nor U9682 (N_9682,N_8401,N_8257);
or U9683 (N_9683,N_8313,N_8193);
and U9684 (N_9684,N_8141,N_8245);
nand U9685 (N_9685,N_8470,N_8219);
or U9686 (N_9686,N_8550,N_8381);
or U9687 (N_9687,N_8365,N_8413);
and U9688 (N_9688,N_8449,N_8563);
and U9689 (N_9689,N_8986,N_8600);
nor U9690 (N_9690,N_8445,N_8622);
and U9691 (N_9691,N_8928,N_8005);
and U9692 (N_9692,N_8418,N_8730);
nor U9693 (N_9693,N_8632,N_8179);
or U9694 (N_9694,N_8213,N_8804);
or U9695 (N_9695,N_8470,N_8656);
and U9696 (N_9696,N_8195,N_8436);
and U9697 (N_9697,N_8224,N_8499);
and U9698 (N_9698,N_8364,N_8066);
nand U9699 (N_9699,N_8965,N_8714);
nor U9700 (N_9700,N_8782,N_8561);
nand U9701 (N_9701,N_8751,N_8303);
or U9702 (N_9702,N_8814,N_8659);
xnor U9703 (N_9703,N_8897,N_8347);
nand U9704 (N_9704,N_8058,N_8492);
and U9705 (N_9705,N_8716,N_8293);
or U9706 (N_9706,N_8708,N_8674);
or U9707 (N_9707,N_8306,N_8006);
xor U9708 (N_9708,N_8245,N_8627);
and U9709 (N_9709,N_8482,N_8284);
nand U9710 (N_9710,N_8400,N_8224);
nor U9711 (N_9711,N_8219,N_8492);
nor U9712 (N_9712,N_8509,N_8156);
nor U9713 (N_9713,N_8601,N_8297);
and U9714 (N_9714,N_8868,N_8570);
nand U9715 (N_9715,N_8964,N_8053);
nand U9716 (N_9716,N_8117,N_8826);
nand U9717 (N_9717,N_8611,N_8694);
nor U9718 (N_9718,N_8352,N_8820);
or U9719 (N_9719,N_8849,N_8260);
and U9720 (N_9720,N_8275,N_8808);
nand U9721 (N_9721,N_8671,N_8743);
xnor U9722 (N_9722,N_8016,N_8718);
and U9723 (N_9723,N_8774,N_8698);
nor U9724 (N_9724,N_8811,N_8937);
xnor U9725 (N_9725,N_8283,N_8619);
nor U9726 (N_9726,N_8435,N_8729);
nand U9727 (N_9727,N_8526,N_8586);
xnor U9728 (N_9728,N_8282,N_8915);
and U9729 (N_9729,N_8786,N_8323);
nor U9730 (N_9730,N_8297,N_8446);
nand U9731 (N_9731,N_8770,N_8787);
nor U9732 (N_9732,N_8820,N_8039);
nor U9733 (N_9733,N_8519,N_8515);
nor U9734 (N_9734,N_8660,N_8969);
nand U9735 (N_9735,N_8076,N_8433);
or U9736 (N_9736,N_8721,N_8955);
nor U9737 (N_9737,N_8804,N_8718);
nand U9738 (N_9738,N_8436,N_8522);
and U9739 (N_9739,N_8156,N_8522);
nand U9740 (N_9740,N_8546,N_8960);
xor U9741 (N_9741,N_8839,N_8808);
xnor U9742 (N_9742,N_8637,N_8959);
nor U9743 (N_9743,N_8534,N_8102);
nand U9744 (N_9744,N_8627,N_8802);
nor U9745 (N_9745,N_8607,N_8254);
or U9746 (N_9746,N_8298,N_8055);
and U9747 (N_9747,N_8925,N_8517);
xor U9748 (N_9748,N_8674,N_8205);
or U9749 (N_9749,N_8293,N_8392);
nor U9750 (N_9750,N_8607,N_8782);
and U9751 (N_9751,N_8213,N_8029);
nor U9752 (N_9752,N_8419,N_8406);
nor U9753 (N_9753,N_8290,N_8473);
nand U9754 (N_9754,N_8262,N_8223);
xnor U9755 (N_9755,N_8592,N_8113);
xor U9756 (N_9756,N_8180,N_8409);
xnor U9757 (N_9757,N_8395,N_8413);
nand U9758 (N_9758,N_8775,N_8867);
or U9759 (N_9759,N_8618,N_8403);
xnor U9760 (N_9760,N_8278,N_8413);
and U9761 (N_9761,N_8904,N_8764);
nor U9762 (N_9762,N_8502,N_8519);
and U9763 (N_9763,N_8483,N_8730);
xnor U9764 (N_9764,N_8461,N_8117);
and U9765 (N_9765,N_8452,N_8714);
nand U9766 (N_9766,N_8361,N_8780);
and U9767 (N_9767,N_8178,N_8622);
or U9768 (N_9768,N_8660,N_8641);
xor U9769 (N_9769,N_8319,N_8476);
xnor U9770 (N_9770,N_8327,N_8204);
nor U9771 (N_9771,N_8492,N_8834);
and U9772 (N_9772,N_8516,N_8336);
and U9773 (N_9773,N_8500,N_8471);
nor U9774 (N_9774,N_8696,N_8084);
or U9775 (N_9775,N_8626,N_8115);
nand U9776 (N_9776,N_8548,N_8070);
nand U9777 (N_9777,N_8980,N_8430);
or U9778 (N_9778,N_8837,N_8133);
nor U9779 (N_9779,N_8916,N_8301);
xnor U9780 (N_9780,N_8295,N_8294);
or U9781 (N_9781,N_8505,N_8818);
xor U9782 (N_9782,N_8020,N_8056);
and U9783 (N_9783,N_8171,N_8506);
xnor U9784 (N_9784,N_8794,N_8524);
or U9785 (N_9785,N_8517,N_8141);
or U9786 (N_9786,N_8793,N_8390);
nand U9787 (N_9787,N_8650,N_8967);
xor U9788 (N_9788,N_8130,N_8410);
or U9789 (N_9789,N_8480,N_8199);
nor U9790 (N_9790,N_8619,N_8155);
or U9791 (N_9791,N_8988,N_8173);
and U9792 (N_9792,N_8684,N_8400);
nor U9793 (N_9793,N_8572,N_8778);
or U9794 (N_9794,N_8153,N_8992);
xnor U9795 (N_9795,N_8737,N_8408);
nor U9796 (N_9796,N_8986,N_8640);
xor U9797 (N_9797,N_8464,N_8390);
nor U9798 (N_9798,N_8372,N_8497);
and U9799 (N_9799,N_8720,N_8747);
xnor U9800 (N_9800,N_8805,N_8115);
or U9801 (N_9801,N_8973,N_8648);
and U9802 (N_9802,N_8304,N_8245);
nand U9803 (N_9803,N_8766,N_8542);
or U9804 (N_9804,N_8185,N_8101);
and U9805 (N_9805,N_8562,N_8692);
nand U9806 (N_9806,N_8753,N_8269);
or U9807 (N_9807,N_8191,N_8394);
nor U9808 (N_9808,N_8784,N_8762);
and U9809 (N_9809,N_8295,N_8648);
nor U9810 (N_9810,N_8283,N_8031);
nor U9811 (N_9811,N_8086,N_8983);
or U9812 (N_9812,N_8664,N_8465);
or U9813 (N_9813,N_8473,N_8836);
nand U9814 (N_9814,N_8936,N_8973);
xor U9815 (N_9815,N_8940,N_8345);
nand U9816 (N_9816,N_8038,N_8848);
and U9817 (N_9817,N_8897,N_8806);
nor U9818 (N_9818,N_8251,N_8769);
nand U9819 (N_9819,N_8502,N_8601);
nand U9820 (N_9820,N_8223,N_8464);
and U9821 (N_9821,N_8703,N_8530);
xnor U9822 (N_9822,N_8538,N_8885);
and U9823 (N_9823,N_8704,N_8222);
and U9824 (N_9824,N_8326,N_8730);
or U9825 (N_9825,N_8122,N_8638);
nand U9826 (N_9826,N_8321,N_8642);
and U9827 (N_9827,N_8559,N_8178);
nand U9828 (N_9828,N_8507,N_8963);
or U9829 (N_9829,N_8897,N_8632);
or U9830 (N_9830,N_8104,N_8840);
xnor U9831 (N_9831,N_8182,N_8063);
xnor U9832 (N_9832,N_8808,N_8510);
nor U9833 (N_9833,N_8464,N_8727);
xor U9834 (N_9834,N_8324,N_8178);
nand U9835 (N_9835,N_8185,N_8148);
xnor U9836 (N_9836,N_8813,N_8636);
nor U9837 (N_9837,N_8632,N_8929);
nor U9838 (N_9838,N_8469,N_8883);
or U9839 (N_9839,N_8812,N_8152);
xnor U9840 (N_9840,N_8244,N_8845);
and U9841 (N_9841,N_8339,N_8407);
xor U9842 (N_9842,N_8674,N_8749);
or U9843 (N_9843,N_8984,N_8694);
and U9844 (N_9844,N_8319,N_8070);
and U9845 (N_9845,N_8878,N_8439);
and U9846 (N_9846,N_8155,N_8594);
and U9847 (N_9847,N_8509,N_8487);
or U9848 (N_9848,N_8892,N_8013);
nor U9849 (N_9849,N_8371,N_8440);
and U9850 (N_9850,N_8867,N_8191);
nor U9851 (N_9851,N_8163,N_8061);
nor U9852 (N_9852,N_8989,N_8795);
and U9853 (N_9853,N_8672,N_8578);
nor U9854 (N_9854,N_8696,N_8196);
or U9855 (N_9855,N_8158,N_8392);
nor U9856 (N_9856,N_8764,N_8132);
or U9857 (N_9857,N_8075,N_8988);
and U9858 (N_9858,N_8142,N_8965);
xor U9859 (N_9859,N_8445,N_8933);
xor U9860 (N_9860,N_8515,N_8989);
or U9861 (N_9861,N_8917,N_8136);
xor U9862 (N_9862,N_8503,N_8912);
nor U9863 (N_9863,N_8624,N_8464);
or U9864 (N_9864,N_8252,N_8469);
or U9865 (N_9865,N_8642,N_8650);
xnor U9866 (N_9866,N_8078,N_8602);
and U9867 (N_9867,N_8860,N_8029);
nand U9868 (N_9868,N_8902,N_8690);
nor U9869 (N_9869,N_8749,N_8794);
nand U9870 (N_9870,N_8374,N_8739);
and U9871 (N_9871,N_8375,N_8165);
nand U9872 (N_9872,N_8698,N_8587);
xnor U9873 (N_9873,N_8030,N_8318);
nor U9874 (N_9874,N_8132,N_8507);
nand U9875 (N_9875,N_8798,N_8755);
xor U9876 (N_9876,N_8180,N_8715);
or U9877 (N_9877,N_8246,N_8432);
and U9878 (N_9878,N_8844,N_8704);
xor U9879 (N_9879,N_8173,N_8489);
nand U9880 (N_9880,N_8410,N_8530);
or U9881 (N_9881,N_8251,N_8748);
nand U9882 (N_9882,N_8889,N_8429);
xnor U9883 (N_9883,N_8085,N_8192);
or U9884 (N_9884,N_8783,N_8232);
nor U9885 (N_9885,N_8409,N_8327);
nor U9886 (N_9886,N_8333,N_8497);
nand U9887 (N_9887,N_8872,N_8825);
or U9888 (N_9888,N_8018,N_8754);
or U9889 (N_9889,N_8249,N_8848);
or U9890 (N_9890,N_8756,N_8422);
or U9891 (N_9891,N_8646,N_8086);
and U9892 (N_9892,N_8059,N_8743);
xnor U9893 (N_9893,N_8842,N_8708);
and U9894 (N_9894,N_8881,N_8479);
nand U9895 (N_9895,N_8418,N_8621);
xor U9896 (N_9896,N_8377,N_8568);
xor U9897 (N_9897,N_8932,N_8708);
and U9898 (N_9898,N_8447,N_8198);
and U9899 (N_9899,N_8538,N_8467);
nand U9900 (N_9900,N_8712,N_8192);
xnor U9901 (N_9901,N_8632,N_8980);
xor U9902 (N_9902,N_8868,N_8050);
or U9903 (N_9903,N_8219,N_8775);
and U9904 (N_9904,N_8154,N_8638);
or U9905 (N_9905,N_8700,N_8460);
or U9906 (N_9906,N_8046,N_8558);
xor U9907 (N_9907,N_8900,N_8764);
nand U9908 (N_9908,N_8415,N_8064);
or U9909 (N_9909,N_8667,N_8918);
xor U9910 (N_9910,N_8277,N_8724);
or U9911 (N_9911,N_8597,N_8399);
nor U9912 (N_9912,N_8937,N_8063);
or U9913 (N_9913,N_8171,N_8493);
and U9914 (N_9914,N_8752,N_8196);
nor U9915 (N_9915,N_8164,N_8442);
nand U9916 (N_9916,N_8167,N_8391);
nand U9917 (N_9917,N_8638,N_8769);
nand U9918 (N_9918,N_8072,N_8666);
xnor U9919 (N_9919,N_8460,N_8876);
xor U9920 (N_9920,N_8480,N_8693);
or U9921 (N_9921,N_8229,N_8284);
or U9922 (N_9922,N_8357,N_8323);
or U9923 (N_9923,N_8383,N_8586);
xnor U9924 (N_9924,N_8334,N_8959);
xnor U9925 (N_9925,N_8784,N_8754);
and U9926 (N_9926,N_8025,N_8522);
nor U9927 (N_9927,N_8813,N_8955);
nand U9928 (N_9928,N_8454,N_8332);
nor U9929 (N_9929,N_8166,N_8664);
or U9930 (N_9930,N_8926,N_8790);
xor U9931 (N_9931,N_8282,N_8983);
nor U9932 (N_9932,N_8620,N_8926);
nor U9933 (N_9933,N_8060,N_8005);
xnor U9934 (N_9934,N_8349,N_8066);
nand U9935 (N_9935,N_8977,N_8179);
and U9936 (N_9936,N_8659,N_8478);
or U9937 (N_9937,N_8796,N_8292);
xnor U9938 (N_9938,N_8930,N_8833);
xnor U9939 (N_9939,N_8666,N_8398);
nor U9940 (N_9940,N_8918,N_8220);
or U9941 (N_9941,N_8910,N_8671);
nand U9942 (N_9942,N_8581,N_8905);
nand U9943 (N_9943,N_8274,N_8548);
xor U9944 (N_9944,N_8439,N_8033);
nor U9945 (N_9945,N_8163,N_8091);
and U9946 (N_9946,N_8174,N_8522);
or U9947 (N_9947,N_8357,N_8272);
nor U9948 (N_9948,N_8725,N_8117);
xnor U9949 (N_9949,N_8119,N_8323);
and U9950 (N_9950,N_8999,N_8455);
nor U9951 (N_9951,N_8464,N_8447);
or U9952 (N_9952,N_8460,N_8818);
or U9953 (N_9953,N_8708,N_8211);
and U9954 (N_9954,N_8385,N_8458);
xor U9955 (N_9955,N_8848,N_8029);
xnor U9956 (N_9956,N_8743,N_8078);
nor U9957 (N_9957,N_8355,N_8652);
nor U9958 (N_9958,N_8470,N_8217);
or U9959 (N_9959,N_8945,N_8106);
nor U9960 (N_9960,N_8668,N_8469);
and U9961 (N_9961,N_8856,N_8682);
and U9962 (N_9962,N_8702,N_8336);
and U9963 (N_9963,N_8828,N_8732);
and U9964 (N_9964,N_8654,N_8156);
nor U9965 (N_9965,N_8545,N_8869);
and U9966 (N_9966,N_8763,N_8894);
nor U9967 (N_9967,N_8736,N_8587);
xnor U9968 (N_9968,N_8758,N_8507);
nand U9969 (N_9969,N_8934,N_8272);
and U9970 (N_9970,N_8429,N_8103);
xor U9971 (N_9971,N_8882,N_8805);
or U9972 (N_9972,N_8461,N_8996);
and U9973 (N_9973,N_8906,N_8728);
xor U9974 (N_9974,N_8938,N_8582);
or U9975 (N_9975,N_8598,N_8441);
or U9976 (N_9976,N_8350,N_8797);
nor U9977 (N_9977,N_8651,N_8682);
nor U9978 (N_9978,N_8543,N_8467);
nand U9979 (N_9979,N_8875,N_8091);
or U9980 (N_9980,N_8298,N_8072);
xnor U9981 (N_9981,N_8182,N_8520);
and U9982 (N_9982,N_8352,N_8675);
or U9983 (N_9983,N_8748,N_8221);
and U9984 (N_9984,N_8825,N_8991);
nand U9985 (N_9985,N_8550,N_8415);
xor U9986 (N_9986,N_8957,N_8423);
xnor U9987 (N_9987,N_8440,N_8036);
nor U9988 (N_9988,N_8827,N_8138);
nand U9989 (N_9989,N_8644,N_8403);
xnor U9990 (N_9990,N_8901,N_8575);
and U9991 (N_9991,N_8889,N_8018);
xnor U9992 (N_9992,N_8180,N_8520);
or U9993 (N_9993,N_8253,N_8425);
or U9994 (N_9994,N_8573,N_8856);
xor U9995 (N_9995,N_8239,N_8941);
or U9996 (N_9996,N_8838,N_8090);
or U9997 (N_9997,N_8272,N_8146);
nor U9998 (N_9998,N_8784,N_8373);
nor U9999 (N_9999,N_8349,N_8388);
nor U10000 (N_10000,N_9832,N_9779);
xnor U10001 (N_10001,N_9331,N_9949);
xnor U10002 (N_10002,N_9287,N_9786);
and U10003 (N_10003,N_9788,N_9935);
and U10004 (N_10004,N_9611,N_9849);
and U10005 (N_10005,N_9439,N_9640);
xnor U10006 (N_10006,N_9704,N_9534);
nand U10007 (N_10007,N_9279,N_9450);
nand U10008 (N_10008,N_9032,N_9666);
and U10009 (N_10009,N_9566,N_9511);
nand U10010 (N_10010,N_9000,N_9319);
or U10011 (N_10011,N_9738,N_9440);
and U10012 (N_10012,N_9307,N_9193);
xor U10013 (N_10013,N_9767,N_9321);
nor U10014 (N_10014,N_9557,N_9376);
xnor U10015 (N_10015,N_9838,N_9172);
nand U10016 (N_10016,N_9411,N_9750);
or U10017 (N_10017,N_9651,N_9845);
nand U10018 (N_10018,N_9985,N_9424);
nand U10019 (N_10019,N_9427,N_9490);
nand U10020 (N_10020,N_9066,N_9471);
nor U10021 (N_10021,N_9434,N_9360);
nand U10022 (N_10022,N_9273,N_9400);
nor U10023 (N_10023,N_9748,N_9372);
and U10024 (N_10024,N_9100,N_9844);
nor U10025 (N_10025,N_9834,N_9665);
xor U10026 (N_10026,N_9910,N_9064);
nand U10027 (N_10027,N_9368,N_9054);
and U10028 (N_10028,N_9098,N_9495);
nor U10029 (N_10029,N_9728,N_9037);
nor U10030 (N_10030,N_9409,N_9455);
xnor U10031 (N_10031,N_9686,N_9426);
and U10032 (N_10032,N_9795,N_9463);
nand U10033 (N_10033,N_9960,N_9417);
or U10034 (N_10034,N_9496,N_9751);
nand U10035 (N_10035,N_9710,N_9248);
xor U10036 (N_10036,N_9310,N_9452);
nor U10037 (N_10037,N_9599,N_9225);
nor U10038 (N_10038,N_9993,N_9161);
and U10039 (N_10039,N_9585,N_9291);
or U10040 (N_10040,N_9829,N_9071);
nor U10041 (N_10041,N_9873,N_9869);
nor U10042 (N_10042,N_9370,N_9460);
nor U10043 (N_10043,N_9027,N_9092);
xor U10044 (N_10044,N_9796,N_9862);
xnor U10045 (N_10045,N_9604,N_9180);
nor U10046 (N_10046,N_9264,N_9652);
nand U10047 (N_10047,N_9997,N_9777);
nand U10048 (N_10048,N_9893,N_9923);
nor U10049 (N_10049,N_9358,N_9648);
xor U10050 (N_10050,N_9116,N_9811);
or U10051 (N_10051,N_9079,N_9660);
nor U10052 (N_10052,N_9941,N_9057);
nand U10053 (N_10053,N_9277,N_9323);
xor U10054 (N_10054,N_9864,N_9617);
and U10055 (N_10055,N_9663,N_9999);
and U10056 (N_10056,N_9930,N_9252);
and U10057 (N_10057,N_9076,N_9715);
nor U10058 (N_10058,N_9757,N_9645);
nand U10059 (N_10059,N_9612,N_9888);
and U10060 (N_10060,N_9669,N_9018);
nor U10061 (N_10061,N_9934,N_9764);
or U10062 (N_10062,N_9355,N_9654);
xnor U10063 (N_10063,N_9972,N_9322);
or U10064 (N_10064,N_9553,N_9241);
and U10065 (N_10065,N_9123,N_9026);
or U10066 (N_10066,N_9905,N_9254);
or U10067 (N_10067,N_9384,N_9213);
and U10068 (N_10068,N_9973,N_9635);
nand U10069 (N_10069,N_9224,N_9084);
nand U10070 (N_10070,N_9632,N_9919);
and U10071 (N_10071,N_9695,N_9314);
xor U10072 (N_10072,N_9031,N_9001);
nand U10073 (N_10073,N_9379,N_9573);
or U10074 (N_10074,N_9181,N_9917);
nand U10075 (N_10075,N_9067,N_9402);
or U10076 (N_10076,N_9294,N_9883);
and U10077 (N_10077,N_9647,N_9984);
nand U10078 (N_10078,N_9774,N_9721);
and U10079 (N_10079,N_9624,N_9005);
nor U10080 (N_10080,N_9349,N_9684);
or U10081 (N_10081,N_9746,N_9316);
xor U10082 (N_10082,N_9190,N_9664);
and U10083 (N_10083,N_9244,N_9661);
xnor U10084 (N_10084,N_9170,N_9741);
nand U10085 (N_10085,N_9073,N_9565);
and U10086 (N_10086,N_9288,N_9994);
xor U10087 (N_10087,N_9982,N_9311);
xor U10088 (N_10088,N_9404,N_9183);
or U10089 (N_10089,N_9709,N_9546);
and U10090 (N_10090,N_9278,N_9544);
nand U10091 (N_10091,N_9465,N_9812);
nand U10092 (N_10092,N_9242,N_9348);
nand U10093 (N_10093,N_9870,N_9211);
and U10094 (N_10094,N_9769,N_9313);
or U10095 (N_10095,N_9035,N_9149);
or U10096 (N_10096,N_9503,N_9042);
or U10097 (N_10097,N_9050,N_9334);
or U10098 (N_10098,N_9520,N_9247);
and U10099 (N_10099,N_9043,N_9970);
xor U10100 (N_10100,N_9898,N_9979);
and U10101 (N_10101,N_9320,N_9399);
nand U10102 (N_10102,N_9528,N_9276);
nand U10103 (N_10103,N_9229,N_9397);
or U10104 (N_10104,N_9878,N_9095);
and U10105 (N_10105,N_9706,N_9594);
xnor U10106 (N_10106,N_9406,N_9938);
nor U10107 (N_10107,N_9713,N_9430);
nor U10108 (N_10108,N_9539,N_9782);
and U10109 (N_10109,N_9559,N_9950);
and U10110 (N_10110,N_9822,N_9630);
and U10111 (N_10111,N_9292,N_9639);
xnor U10112 (N_10112,N_9340,N_9998);
xor U10113 (N_10113,N_9965,N_9816);
nor U10114 (N_10114,N_9185,N_9256);
nor U10115 (N_10115,N_9049,N_9041);
nand U10116 (N_10116,N_9521,N_9964);
or U10117 (N_10117,N_9489,N_9238);
nand U10118 (N_10118,N_9201,N_9343);
nor U10119 (N_10119,N_9628,N_9234);
nand U10120 (N_10120,N_9672,N_9129);
xor U10121 (N_10121,N_9494,N_9646);
and U10122 (N_10122,N_9702,N_9415);
or U10123 (N_10123,N_9515,N_9009);
xnor U10124 (N_10124,N_9936,N_9697);
nand U10125 (N_10125,N_9872,N_9270);
and U10126 (N_10126,N_9016,N_9740);
nand U10127 (N_10127,N_9700,N_9033);
or U10128 (N_10128,N_9516,N_9570);
and U10129 (N_10129,N_9086,N_9433);
xnor U10130 (N_10130,N_9462,N_9363);
and U10131 (N_10131,N_9112,N_9113);
xor U10132 (N_10132,N_9863,N_9887);
and U10133 (N_10133,N_9538,N_9852);
and U10134 (N_10134,N_9479,N_9030);
xor U10135 (N_10135,N_9194,N_9192);
nand U10136 (N_10136,N_9051,N_9861);
or U10137 (N_10137,N_9217,N_9290);
and U10138 (N_10138,N_9703,N_9245);
nor U10139 (N_10139,N_9961,N_9535);
and U10140 (N_10140,N_9140,N_9874);
xor U10141 (N_10141,N_9246,N_9563);
xnor U10142 (N_10142,N_9596,N_9304);
or U10143 (N_10143,N_9168,N_9882);
xor U10144 (N_10144,N_9745,N_9135);
nand U10145 (N_10145,N_9359,N_9101);
or U10146 (N_10146,N_9002,N_9267);
and U10147 (N_10147,N_9357,N_9945);
xor U10148 (N_10148,N_9527,N_9601);
xnor U10149 (N_10149,N_9877,N_9326);
and U10150 (N_10150,N_9231,N_9127);
nand U10151 (N_10151,N_9044,N_9678);
or U10152 (N_10152,N_9093,N_9283);
and U10153 (N_10153,N_9674,N_9590);
nand U10154 (N_10154,N_9235,N_9815);
nand U10155 (N_10155,N_9744,N_9581);
nor U10156 (N_10156,N_9731,N_9164);
and U10157 (N_10157,N_9913,N_9166);
xnor U10158 (N_10158,N_9301,N_9438);
or U10159 (N_10159,N_9912,N_9218);
nor U10160 (N_10160,N_9345,N_9775);
xor U10161 (N_10161,N_9159,N_9146);
and U10162 (N_10162,N_9856,N_9006);
nand U10163 (N_10163,N_9371,N_9160);
and U10164 (N_10164,N_9668,N_9395);
xnor U10165 (N_10165,N_9980,N_9763);
xnor U10166 (N_10166,N_9853,N_9029);
xor U10167 (N_10167,N_9134,N_9837);
or U10168 (N_10168,N_9718,N_9924);
xor U10169 (N_10169,N_9077,N_9588);
nand U10170 (N_10170,N_9981,N_9631);
nand U10171 (N_10171,N_9352,N_9391);
and U10172 (N_10172,N_9720,N_9121);
nand U10173 (N_10173,N_9658,N_9023);
nor U10174 (N_10174,N_9650,N_9875);
xor U10175 (N_10175,N_9955,N_9475);
nand U10176 (N_10176,N_9039,N_9068);
xor U10177 (N_10177,N_9346,N_9509);
xnor U10178 (N_10178,N_9797,N_9541);
nand U10179 (N_10179,N_9677,N_9813);
xnor U10180 (N_10180,N_9714,N_9025);
or U10181 (N_10181,N_9470,N_9827);
and U10182 (N_10182,N_9673,N_9550);
and U10183 (N_10183,N_9036,N_9459);
nand U10184 (N_10184,N_9132,N_9342);
nand U10185 (N_10185,N_9469,N_9947);
nor U10186 (N_10186,N_9727,N_9881);
nand U10187 (N_10187,N_9808,N_9966);
nand U10188 (N_10188,N_9493,N_9333);
nor U10189 (N_10189,N_9420,N_9447);
nor U10190 (N_10190,N_9189,N_9591);
nor U10191 (N_10191,N_9053,N_9724);
nor U10192 (N_10192,N_9885,N_9806);
and U10193 (N_10193,N_9472,N_9986);
and U10194 (N_10194,N_9569,N_9173);
and U10195 (N_10195,N_9297,N_9922);
nor U10196 (N_10196,N_9605,N_9125);
nand U10197 (N_10197,N_9094,N_9843);
and U10198 (N_10198,N_9303,N_9776);
nor U10199 (N_10199,N_9103,N_9486);
nand U10200 (N_10200,N_9906,N_9070);
and U10201 (N_10201,N_9722,N_9477);
nand U10202 (N_10202,N_9943,N_9162);
or U10203 (N_10203,N_9389,N_9122);
or U10204 (N_10204,N_9377,N_9328);
xor U10205 (N_10205,N_9904,N_9339);
and U10206 (N_10206,N_9099,N_9756);
and U10207 (N_10207,N_9848,N_9753);
xnor U10208 (N_10208,N_9963,N_9586);
nand U10209 (N_10209,N_9988,N_9532);
xnor U10210 (N_10210,N_9265,N_9158);
xnor U10211 (N_10211,N_9369,N_9800);
nor U10212 (N_10212,N_9012,N_9860);
nor U10213 (N_10213,N_9271,N_9719);
nand U10214 (N_10214,N_9131,N_9380);
nand U10215 (N_10215,N_9268,N_9991);
and U10216 (N_10216,N_9641,N_9188);
xnor U10217 (N_10217,N_9754,N_9560);
nor U10218 (N_10218,N_9858,N_9995);
nand U10219 (N_10219,N_9350,N_9736);
and U10220 (N_10220,N_9024,N_9770);
and U10221 (N_10221,N_9280,N_9046);
nand U10222 (N_10222,N_9083,N_9347);
and U10223 (N_10223,N_9208,N_9743);
xnor U10224 (N_10224,N_9968,N_9216);
and U10225 (N_10225,N_9701,N_9107);
nand U10226 (N_10226,N_9990,N_9859);
or U10227 (N_10227,N_9381,N_9284);
or U10228 (N_10228,N_9790,N_9236);
nor U10229 (N_10229,N_9065,N_9078);
and U10230 (N_10230,N_9466,N_9257);
nand U10231 (N_10231,N_9413,N_9143);
nand U10232 (N_10232,N_9820,N_9163);
xor U10233 (N_10233,N_9846,N_9761);
xor U10234 (N_10234,N_9890,N_9351);
xnor U10235 (N_10235,N_9087,N_9004);
or U10236 (N_10236,N_9567,N_9821);
and U10237 (N_10237,N_9962,N_9155);
or U10238 (N_10238,N_9689,N_9847);
and U10239 (N_10239,N_9136,N_9772);
and U10240 (N_10240,N_9682,N_9457);
nor U10241 (N_10241,N_9819,N_9491);
and U10242 (N_10242,N_9732,N_9212);
xor U10243 (N_10243,N_9536,N_9197);
xor U10244 (N_10244,N_9809,N_9220);
xor U10245 (N_10245,N_9778,N_9914);
nand U10246 (N_10246,N_9974,N_9106);
or U10247 (N_10247,N_9971,N_9476);
xnor U10248 (N_10248,N_9685,N_9047);
and U10249 (N_10249,N_9556,N_9531);
or U10250 (N_10250,N_9336,N_9382);
or U10251 (N_10251,N_9946,N_9393);
nor U10252 (N_10252,N_9854,N_9603);
and U10253 (N_10253,N_9221,N_9422);
nand U10254 (N_10254,N_9442,N_9865);
xnor U10255 (N_10255,N_9783,N_9487);
or U10256 (N_10256,N_9387,N_9354);
nor U10257 (N_10257,N_9976,N_9554);
nor U10258 (N_10258,N_9578,N_9766);
nor U10259 (N_10259,N_9620,N_9437);
and U10260 (N_10260,N_9742,N_9329);
or U10261 (N_10261,N_9187,N_9826);
nor U10262 (N_10262,N_9418,N_9525);
nand U10263 (N_10263,N_9894,N_9571);
and U10264 (N_10264,N_9667,N_9014);
nand U10265 (N_10265,N_9281,N_9622);
xor U10266 (N_10266,N_9299,N_9653);
nor U10267 (N_10267,N_9088,N_9337);
nand U10268 (N_10268,N_9482,N_9773);
nor U10269 (N_10269,N_9332,N_9072);
xor U10270 (N_10270,N_9671,N_9587);
nor U10271 (N_10271,N_9705,N_9925);
or U10272 (N_10272,N_9805,N_9927);
nor U10273 (N_10273,N_9633,N_9260);
or U10274 (N_10274,N_9219,N_9451);
nand U10275 (N_10275,N_9958,N_9504);
and U10276 (N_10276,N_9801,N_9978);
nand U10277 (N_10277,N_9169,N_9537);
or U10278 (N_10278,N_9010,N_9110);
or U10279 (N_10279,N_9954,N_9687);
and U10280 (N_10280,N_9052,N_9931);
nand U10281 (N_10281,N_9282,N_9759);
and U10282 (N_10282,N_9214,N_9405);
or U10283 (N_10283,N_9419,N_9215);
nand U10284 (N_10284,N_9614,N_9484);
nand U10285 (N_10285,N_9226,N_9200);
nand U10286 (N_10286,N_9823,N_9597);
and U10287 (N_10287,N_9325,N_9108);
nand U10288 (N_10288,N_9388,N_9436);
and U10289 (N_10289,N_9081,N_9755);
nand U10290 (N_10290,N_9517,N_9341);
xor U10291 (N_10291,N_9824,N_9485);
nor U10292 (N_10292,N_9063,N_9488);
or U10293 (N_10293,N_9627,N_9921);
nor U10294 (N_10294,N_9825,N_9787);
nand U10295 (N_10295,N_9625,N_9643);
and U10296 (N_10296,N_9866,N_9940);
nand U10297 (N_10297,N_9562,N_9114);
and U10298 (N_10298,N_9842,N_9996);
or U10299 (N_10299,N_9186,N_9969);
or U10300 (N_10300,N_9891,N_9302);
and U10301 (N_10301,N_9799,N_9120);
xor U10302 (N_10302,N_9977,N_9207);
nand U10303 (N_10303,N_9261,N_9007);
and U10304 (N_10304,N_9711,N_9792);
or U10305 (N_10305,N_9681,N_9045);
nand U10306 (N_10306,N_9416,N_9202);
nor U10307 (N_10307,N_9378,N_9659);
xnor U10308 (N_10308,N_9456,N_9552);
xnor U10309 (N_10309,N_9916,N_9109);
and U10310 (N_10310,N_9699,N_9523);
xor U10311 (N_10311,N_9895,N_9240);
nor U10312 (N_10312,N_9274,N_9884);
or U10313 (N_10313,N_9028,N_9621);
or U10314 (N_10314,N_9729,N_9174);
nor U10315 (N_10315,N_9577,N_9992);
and U10316 (N_10316,N_9431,N_9983);
nand U10317 (N_10317,N_9871,N_9555);
nor U10318 (N_10318,N_9008,N_9747);
nand U10319 (N_10319,N_9879,N_9153);
or U10320 (N_10320,N_9385,N_9074);
or U10321 (N_10321,N_9952,N_9449);
xor U10322 (N_10322,N_9785,N_9392);
nand U10323 (N_10323,N_9735,N_9119);
xor U10324 (N_10324,N_9752,N_9549);
or U10325 (N_10325,N_9768,N_9897);
nor U10326 (N_10326,N_9580,N_9227);
nand U10327 (N_10327,N_9269,N_9414);
and U10328 (N_10328,N_9263,N_9429);
nand U10329 (N_10329,N_9144,N_9038);
nor U10330 (N_10330,N_9019,N_9831);
nand U10331 (N_10331,N_9529,N_9467);
and U10332 (N_10332,N_9835,N_9435);
or U10333 (N_10333,N_9317,N_9505);
xor U10334 (N_10334,N_9111,N_9330);
nand U10335 (N_10335,N_9423,N_9444);
nor U10336 (N_10336,N_9126,N_9059);
or U10337 (N_10337,N_9583,N_9448);
and U10338 (N_10338,N_9089,N_9683);
nor U10339 (N_10339,N_9315,N_9902);
and U10340 (N_10340,N_9441,N_9814);
xnor U10341 (N_10341,N_9401,N_9803);
nand U10342 (N_10342,N_9696,N_9530);
xnor U10343 (N_10343,N_9306,N_9157);
or U10344 (N_10344,N_9483,N_9454);
nor U10345 (N_10345,N_9533,N_9506);
nand U10346 (N_10346,N_9137,N_9607);
nor U10347 (N_10347,N_9867,N_9500);
nand U10348 (N_10348,N_9626,N_9575);
xnor U10349 (N_10349,N_9147,N_9545);
xnor U10350 (N_10350,N_9512,N_9616);
and U10351 (N_10351,N_9464,N_9474);
or U10352 (N_10352,N_9944,N_9758);
and U10353 (N_10353,N_9600,N_9656);
nor U10354 (N_10354,N_9289,N_9818);
xor U10355 (N_10355,N_9295,N_9361);
nand U10356 (N_10356,N_9177,N_9518);
nor U10357 (N_10357,N_9501,N_9375);
xor U10358 (N_10358,N_9903,N_9104);
and U10359 (N_10359,N_9892,N_9386);
and U10360 (N_10360,N_9610,N_9929);
or U10361 (N_10361,N_9508,N_9676);
or U10362 (N_10362,N_9062,N_9876);
or U10363 (N_10363,N_9739,N_9344);
xnor U10364 (N_10364,N_9206,N_9817);
or U10365 (N_10365,N_9445,N_9712);
or U10366 (N_10366,N_9850,N_9096);
xor U10367 (N_10367,N_9021,N_9760);
and U10368 (N_10368,N_9595,N_9765);
nand U10369 (N_10369,N_9151,N_9296);
xor U10370 (N_10370,N_9942,N_9734);
and U10371 (N_10371,N_9698,N_9362);
nor U10372 (N_10372,N_9156,N_9139);
xnor U10373 (N_10373,N_9182,N_9421);
and U10374 (N_10374,N_9398,N_9498);
or U10375 (N_10375,N_9918,N_9353);
nor U10376 (N_10376,N_9239,N_9142);
xnor U10377 (N_10377,N_9896,N_9060);
xor U10378 (N_10378,N_9011,N_9058);
nand U10379 (N_10379,N_9308,N_9798);
or U10380 (N_10380,N_9513,N_9636);
xnor U10381 (N_10381,N_9262,N_9840);
xor U10382 (N_10382,N_9285,N_9613);
and U10383 (N_10383,N_9629,N_9199);
and U10384 (N_10384,N_9547,N_9644);
nand U10385 (N_10385,N_9880,N_9618);
nand U10386 (N_10386,N_9733,N_9967);
nand U10387 (N_10387,N_9075,N_9324);
nand U10388 (N_10388,N_9105,N_9195);
nor U10389 (N_10389,N_9839,N_9243);
and U10390 (N_10390,N_9598,N_9097);
nor U10391 (N_10391,N_9230,N_9022);
or U10392 (N_10392,N_9179,N_9615);
or U10393 (N_10393,N_9374,N_9222);
and U10394 (N_10394,N_9975,N_9857);
and U10395 (N_10395,N_9804,N_9899);
or U10396 (N_10396,N_9040,N_9502);
and U10397 (N_10397,N_9130,N_9507);
nand U10398 (N_10398,N_9953,N_9642);
or U10399 (N_10399,N_9272,N_9886);
nor U10400 (N_10400,N_9499,N_9410);
or U10401 (N_10401,N_9510,N_9841);
nor U10402 (N_10402,N_9184,N_9020);
or U10403 (N_10403,N_9657,N_9138);
xnor U10404 (N_10404,N_9481,N_9249);
or U10405 (N_10405,N_9602,N_9810);
or U10406 (N_10406,N_9367,N_9789);
nor U10407 (N_10407,N_9634,N_9196);
xor U10408 (N_10408,N_9959,N_9055);
and U10409 (N_10409,N_9589,N_9085);
or U10410 (N_10410,N_9572,N_9338);
or U10411 (N_10411,N_9649,N_9833);
or U10412 (N_10412,N_9791,N_9253);
xor U10413 (N_10413,N_9176,N_9623);
nand U10414 (N_10414,N_9128,N_9167);
and U10415 (N_10415,N_9793,N_9048);
nand U10416 (N_10416,N_9606,N_9655);
xnor U10417 (N_10417,N_9209,N_9694);
and U10418 (N_10418,N_9191,N_9900);
and U10419 (N_10419,N_9275,N_9937);
xor U10420 (N_10420,N_9233,N_9412);
and U10421 (N_10421,N_9255,N_9061);
nand U10422 (N_10422,N_9432,N_9150);
and U10423 (N_10423,N_9312,N_9364);
nor U10424 (N_10424,N_9115,N_9680);
nor U10425 (N_10425,N_9383,N_9015);
nor U10426 (N_10426,N_9619,N_9609);
or U10427 (N_10427,N_9939,N_9069);
or U10428 (N_10428,N_9519,N_9210);
and U10429 (N_10429,N_9901,N_9492);
nor U10430 (N_10430,N_9582,N_9118);
nor U10431 (N_10431,N_9670,N_9258);
nor U10432 (N_10432,N_9141,N_9522);
nand U10433 (N_10433,N_9390,N_9468);
nor U10434 (N_10434,N_9920,N_9576);
or U10435 (N_10435,N_9692,N_9707);
and U10436 (N_10436,N_9473,N_9165);
and U10437 (N_10437,N_9951,N_9178);
or U10438 (N_10438,N_9443,N_9828);
or U10439 (N_10439,N_9428,N_9293);
xor U10440 (N_10440,N_9723,N_9458);
or U10441 (N_10441,N_9956,N_9148);
or U10442 (N_10442,N_9584,N_9514);
nor U10443 (N_10443,N_9366,N_9638);
nor U10444 (N_10444,N_9784,N_9855);
and U10445 (N_10445,N_9568,N_9133);
nor U10446 (N_10446,N_9124,N_9730);
nand U10447 (N_10447,N_9781,N_9205);
nand U10448 (N_10448,N_9675,N_9725);
and U10449 (N_10449,N_9228,N_9082);
or U10450 (N_10450,N_9091,N_9989);
nor U10451 (N_10451,N_9551,N_9300);
nor U10452 (N_10452,N_9807,N_9286);
xor U10453 (N_10453,N_9145,N_9356);
xnor U10454 (N_10454,N_9526,N_9851);
nor U10455 (N_10455,N_9453,N_9911);
nor U10456 (N_10456,N_9693,N_9154);
or U10457 (N_10457,N_9592,N_9608);
and U10458 (N_10458,N_9446,N_9497);
or U10459 (N_10459,N_9593,N_9564);
nor U10460 (N_10460,N_9688,N_9933);
or U10461 (N_10461,N_9259,N_9175);
nor U10462 (N_10462,N_9717,N_9034);
nor U10463 (N_10463,N_9558,N_9802);
and U10464 (N_10464,N_9679,N_9203);
and U10465 (N_10465,N_9542,N_9394);
nor U10466 (N_10466,N_9396,N_9726);
and U10467 (N_10467,N_9637,N_9948);
or U10468 (N_10468,N_9232,N_9543);
and U10469 (N_10469,N_9561,N_9928);
xor U10470 (N_10470,N_9762,N_9889);
nand U10471 (N_10471,N_9915,N_9250);
xnor U10472 (N_10472,N_9171,N_9013);
or U10473 (N_10473,N_9780,N_9117);
or U10474 (N_10474,N_9425,N_9056);
nand U10475 (N_10475,N_9908,N_9716);
nor U10476 (N_10476,N_9691,N_9708);
or U10477 (N_10477,N_9868,N_9266);
xnor U10478 (N_10478,N_9926,N_9251);
xnor U10479 (N_10479,N_9403,N_9836);
and U10480 (N_10480,N_9335,N_9461);
nor U10481 (N_10481,N_9080,N_9907);
xor U10482 (N_10482,N_9204,N_9548);
or U10483 (N_10483,N_9771,N_9237);
xor U10484 (N_10484,N_9987,N_9524);
or U10485 (N_10485,N_9152,N_9327);
xor U10486 (N_10486,N_9223,N_9579);
or U10487 (N_10487,N_9309,N_9407);
nand U10488 (N_10488,N_9737,N_9365);
nand U10489 (N_10489,N_9305,N_9090);
nand U10490 (N_10490,N_9690,N_9198);
xnor U10491 (N_10491,N_9408,N_9574);
xnor U10492 (N_10492,N_9480,N_9794);
nand U10493 (N_10493,N_9373,N_9749);
xor U10494 (N_10494,N_9540,N_9830);
xnor U10495 (N_10495,N_9662,N_9318);
and U10496 (N_10496,N_9478,N_9298);
nand U10497 (N_10497,N_9909,N_9017);
or U10498 (N_10498,N_9003,N_9102);
or U10499 (N_10499,N_9932,N_9957);
and U10500 (N_10500,N_9121,N_9911);
nor U10501 (N_10501,N_9573,N_9387);
nor U10502 (N_10502,N_9866,N_9861);
and U10503 (N_10503,N_9824,N_9550);
nand U10504 (N_10504,N_9158,N_9367);
or U10505 (N_10505,N_9417,N_9248);
nor U10506 (N_10506,N_9047,N_9961);
xor U10507 (N_10507,N_9792,N_9362);
nand U10508 (N_10508,N_9630,N_9434);
or U10509 (N_10509,N_9833,N_9530);
and U10510 (N_10510,N_9438,N_9510);
or U10511 (N_10511,N_9674,N_9121);
xnor U10512 (N_10512,N_9269,N_9522);
and U10513 (N_10513,N_9309,N_9797);
or U10514 (N_10514,N_9689,N_9368);
nand U10515 (N_10515,N_9761,N_9895);
nand U10516 (N_10516,N_9505,N_9025);
or U10517 (N_10517,N_9926,N_9353);
nand U10518 (N_10518,N_9372,N_9345);
and U10519 (N_10519,N_9694,N_9500);
xor U10520 (N_10520,N_9681,N_9837);
and U10521 (N_10521,N_9854,N_9308);
and U10522 (N_10522,N_9836,N_9064);
nor U10523 (N_10523,N_9503,N_9056);
or U10524 (N_10524,N_9058,N_9552);
or U10525 (N_10525,N_9602,N_9466);
or U10526 (N_10526,N_9386,N_9431);
and U10527 (N_10527,N_9641,N_9882);
or U10528 (N_10528,N_9315,N_9155);
nand U10529 (N_10529,N_9253,N_9105);
and U10530 (N_10530,N_9828,N_9559);
nand U10531 (N_10531,N_9889,N_9225);
nor U10532 (N_10532,N_9329,N_9500);
xor U10533 (N_10533,N_9728,N_9084);
nand U10534 (N_10534,N_9282,N_9964);
nand U10535 (N_10535,N_9693,N_9043);
xnor U10536 (N_10536,N_9640,N_9782);
and U10537 (N_10537,N_9252,N_9432);
nand U10538 (N_10538,N_9493,N_9532);
and U10539 (N_10539,N_9797,N_9933);
or U10540 (N_10540,N_9174,N_9845);
nand U10541 (N_10541,N_9217,N_9442);
and U10542 (N_10542,N_9435,N_9126);
nor U10543 (N_10543,N_9641,N_9314);
or U10544 (N_10544,N_9673,N_9692);
nor U10545 (N_10545,N_9306,N_9935);
and U10546 (N_10546,N_9427,N_9383);
nor U10547 (N_10547,N_9971,N_9589);
nor U10548 (N_10548,N_9056,N_9891);
or U10549 (N_10549,N_9084,N_9121);
and U10550 (N_10550,N_9207,N_9686);
or U10551 (N_10551,N_9746,N_9479);
or U10552 (N_10552,N_9919,N_9259);
xnor U10553 (N_10553,N_9306,N_9053);
nor U10554 (N_10554,N_9278,N_9800);
xor U10555 (N_10555,N_9726,N_9201);
nor U10556 (N_10556,N_9047,N_9715);
and U10557 (N_10557,N_9120,N_9342);
or U10558 (N_10558,N_9433,N_9006);
or U10559 (N_10559,N_9462,N_9762);
and U10560 (N_10560,N_9846,N_9585);
or U10561 (N_10561,N_9353,N_9526);
or U10562 (N_10562,N_9506,N_9266);
and U10563 (N_10563,N_9437,N_9612);
nor U10564 (N_10564,N_9323,N_9092);
or U10565 (N_10565,N_9821,N_9388);
and U10566 (N_10566,N_9900,N_9218);
nor U10567 (N_10567,N_9324,N_9397);
or U10568 (N_10568,N_9230,N_9494);
nor U10569 (N_10569,N_9158,N_9888);
or U10570 (N_10570,N_9710,N_9354);
and U10571 (N_10571,N_9884,N_9089);
xnor U10572 (N_10572,N_9864,N_9474);
nor U10573 (N_10573,N_9592,N_9536);
nand U10574 (N_10574,N_9478,N_9041);
nor U10575 (N_10575,N_9758,N_9817);
or U10576 (N_10576,N_9145,N_9373);
or U10577 (N_10577,N_9878,N_9435);
nand U10578 (N_10578,N_9050,N_9402);
and U10579 (N_10579,N_9293,N_9702);
or U10580 (N_10580,N_9744,N_9733);
xor U10581 (N_10581,N_9192,N_9661);
or U10582 (N_10582,N_9444,N_9849);
or U10583 (N_10583,N_9150,N_9631);
nor U10584 (N_10584,N_9326,N_9434);
or U10585 (N_10585,N_9770,N_9516);
and U10586 (N_10586,N_9321,N_9435);
nand U10587 (N_10587,N_9586,N_9073);
and U10588 (N_10588,N_9605,N_9847);
and U10589 (N_10589,N_9819,N_9244);
or U10590 (N_10590,N_9104,N_9858);
nand U10591 (N_10591,N_9620,N_9911);
and U10592 (N_10592,N_9860,N_9898);
and U10593 (N_10593,N_9531,N_9389);
or U10594 (N_10594,N_9798,N_9878);
nor U10595 (N_10595,N_9823,N_9580);
xnor U10596 (N_10596,N_9995,N_9866);
xnor U10597 (N_10597,N_9107,N_9455);
nor U10598 (N_10598,N_9025,N_9239);
and U10599 (N_10599,N_9082,N_9815);
nand U10600 (N_10600,N_9796,N_9528);
nor U10601 (N_10601,N_9898,N_9599);
xor U10602 (N_10602,N_9800,N_9322);
nand U10603 (N_10603,N_9274,N_9544);
nand U10604 (N_10604,N_9693,N_9476);
xnor U10605 (N_10605,N_9420,N_9490);
or U10606 (N_10606,N_9370,N_9239);
xor U10607 (N_10607,N_9469,N_9057);
nor U10608 (N_10608,N_9958,N_9191);
nor U10609 (N_10609,N_9679,N_9712);
nor U10610 (N_10610,N_9654,N_9713);
nor U10611 (N_10611,N_9062,N_9998);
xnor U10612 (N_10612,N_9351,N_9882);
and U10613 (N_10613,N_9142,N_9139);
and U10614 (N_10614,N_9605,N_9197);
and U10615 (N_10615,N_9512,N_9916);
nand U10616 (N_10616,N_9256,N_9336);
xnor U10617 (N_10617,N_9346,N_9225);
nor U10618 (N_10618,N_9441,N_9366);
nand U10619 (N_10619,N_9663,N_9895);
or U10620 (N_10620,N_9988,N_9733);
nand U10621 (N_10621,N_9347,N_9163);
and U10622 (N_10622,N_9532,N_9883);
nor U10623 (N_10623,N_9149,N_9234);
nor U10624 (N_10624,N_9091,N_9513);
or U10625 (N_10625,N_9090,N_9793);
nor U10626 (N_10626,N_9513,N_9800);
nor U10627 (N_10627,N_9801,N_9419);
nand U10628 (N_10628,N_9720,N_9972);
xnor U10629 (N_10629,N_9502,N_9867);
xnor U10630 (N_10630,N_9559,N_9254);
or U10631 (N_10631,N_9215,N_9144);
or U10632 (N_10632,N_9013,N_9800);
nand U10633 (N_10633,N_9295,N_9107);
or U10634 (N_10634,N_9110,N_9888);
nor U10635 (N_10635,N_9915,N_9607);
nand U10636 (N_10636,N_9196,N_9200);
xor U10637 (N_10637,N_9587,N_9184);
nand U10638 (N_10638,N_9606,N_9071);
xor U10639 (N_10639,N_9863,N_9895);
nor U10640 (N_10640,N_9659,N_9388);
nand U10641 (N_10641,N_9513,N_9086);
nand U10642 (N_10642,N_9832,N_9208);
nand U10643 (N_10643,N_9001,N_9634);
nand U10644 (N_10644,N_9862,N_9063);
and U10645 (N_10645,N_9889,N_9816);
nor U10646 (N_10646,N_9956,N_9654);
nor U10647 (N_10647,N_9476,N_9998);
or U10648 (N_10648,N_9791,N_9080);
or U10649 (N_10649,N_9273,N_9242);
and U10650 (N_10650,N_9352,N_9209);
xnor U10651 (N_10651,N_9783,N_9714);
nor U10652 (N_10652,N_9096,N_9103);
and U10653 (N_10653,N_9786,N_9364);
and U10654 (N_10654,N_9402,N_9806);
or U10655 (N_10655,N_9552,N_9964);
nor U10656 (N_10656,N_9445,N_9893);
xor U10657 (N_10657,N_9892,N_9223);
nor U10658 (N_10658,N_9874,N_9849);
or U10659 (N_10659,N_9090,N_9503);
nand U10660 (N_10660,N_9299,N_9008);
nand U10661 (N_10661,N_9894,N_9486);
or U10662 (N_10662,N_9373,N_9035);
or U10663 (N_10663,N_9810,N_9635);
nand U10664 (N_10664,N_9932,N_9413);
or U10665 (N_10665,N_9154,N_9052);
nand U10666 (N_10666,N_9437,N_9062);
nor U10667 (N_10667,N_9032,N_9908);
and U10668 (N_10668,N_9110,N_9727);
nor U10669 (N_10669,N_9132,N_9210);
and U10670 (N_10670,N_9732,N_9461);
xor U10671 (N_10671,N_9784,N_9913);
or U10672 (N_10672,N_9631,N_9148);
nand U10673 (N_10673,N_9096,N_9945);
or U10674 (N_10674,N_9980,N_9927);
nor U10675 (N_10675,N_9490,N_9287);
nor U10676 (N_10676,N_9824,N_9162);
nand U10677 (N_10677,N_9285,N_9751);
nand U10678 (N_10678,N_9593,N_9531);
nor U10679 (N_10679,N_9379,N_9676);
nand U10680 (N_10680,N_9166,N_9656);
and U10681 (N_10681,N_9073,N_9890);
nand U10682 (N_10682,N_9040,N_9006);
nand U10683 (N_10683,N_9441,N_9861);
nor U10684 (N_10684,N_9485,N_9655);
nand U10685 (N_10685,N_9862,N_9972);
nor U10686 (N_10686,N_9763,N_9527);
nand U10687 (N_10687,N_9301,N_9333);
nor U10688 (N_10688,N_9618,N_9104);
or U10689 (N_10689,N_9027,N_9198);
nand U10690 (N_10690,N_9890,N_9629);
xor U10691 (N_10691,N_9912,N_9670);
xnor U10692 (N_10692,N_9969,N_9115);
xor U10693 (N_10693,N_9865,N_9408);
or U10694 (N_10694,N_9240,N_9457);
nor U10695 (N_10695,N_9382,N_9722);
xnor U10696 (N_10696,N_9830,N_9472);
nand U10697 (N_10697,N_9684,N_9723);
nand U10698 (N_10698,N_9683,N_9174);
nor U10699 (N_10699,N_9311,N_9801);
xnor U10700 (N_10700,N_9583,N_9184);
nand U10701 (N_10701,N_9220,N_9613);
nand U10702 (N_10702,N_9174,N_9100);
nor U10703 (N_10703,N_9620,N_9632);
or U10704 (N_10704,N_9645,N_9443);
nor U10705 (N_10705,N_9283,N_9410);
nand U10706 (N_10706,N_9235,N_9083);
nor U10707 (N_10707,N_9708,N_9874);
xnor U10708 (N_10708,N_9715,N_9481);
nand U10709 (N_10709,N_9188,N_9273);
nor U10710 (N_10710,N_9481,N_9447);
nand U10711 (N_10711,N_9246,N_9354);
xor U10712 (N_10712,N_9115,N_9073);
nor U10713 (N_10713,N_9276,N_9455);
nor U10714 (N_10714,N_9903,N_9405);
or U10715 (N_10715,N_9282,N_9866);
or U10716 (N_10716,N_9410,N_9664);
nor U10717 (N_10717,N_9705,N_9830);
or U10718 (N_10718,N_9187,N_9003);
xor U10719 (N_10719,N_9029,N_9352);
and U10720 (N_10720,N_9785,N_9989);
or U10721 (N_10721,N_9635,N_9223);
or U10722 (N_10722,N_9965,N_9794);
xnor U10723 (N_10723,N_9515,N_9446);
and U10724 (N_10724,N_9979,N_9491);
xnor U10725 (N_10725,N_9492,N_9553);
nand U10726 (N_10726,N_9636,N_9666);
nor U10727 (N_10727,N_9493,N_9742);
or U10728 (N_10728,N_9492,N_9670);
or U10729 (N_10729,N_9023,N_9281);
xor U10730 (N_10730,N_9870,N_9453);
and U10731 (N_10731,N_9188,N_9027);
nor U10732 (N_10732,N_9043,N_9100);
nand U10733 (N_10733,N_9288,N_9575);
nor U10734 (N_10734,N_9994,N_9323);
nor U10735 (N_10735,N_9565,N_9334);
nor U10736 (N_10736,N_9795,N_9033);
xor U10737 (N_10737,N_9147,N_9604);
nor U10738 (N_10738,N_9191,N_9197);
xnor U10739 (N_10739,N_9069,N_9049);
xor U10740 (N_10740,N_9605,N_9676);
xnor U10741 (N_10741,N_9835,N_9999);
xor U10742 (N_10742,N_9157,N_9551);
or U10743 (N_10743,N_9622,N_9802);
nand U10744 (N_10744,N_9375,N_9865);
nor U10745 (N_10745,N_9692,N_9381);
and U10746 (N_10746,N_9953,N_9788);
xor U10747 (N_10747,N_9914,N_9442);
or U10748 (N_10748,N_9791,N_9989);
or U10749 (N_10749,N_9479,N_9234);
nor U10750 (N_10750,N_9679,N_9686);
nor U10751 (N_10751,N_9816,N_9596);
nand U10752 (N_10752,N_9086,N_9606);
nor U10753 (N_10753,N_9316,N_9092);
and U10754 (N_10754,N_9222,N_9442);
or U10755 (N_10755,N_9664,N_9863);
or U10756 (N_10756,N_9699,N_9765);
or U10757 (N_10757,N_9652,N_9492);
and U10758 (N_10758,N_9094,N_9463);
and U10759 (N_10759,N_9920,N_9300);
or U10760 (N_10760,N_9113,N_9440);
or U10761 (N_10761,N_9671,N_9745);
or U10762 (N_10762,N_9154,N_9144);
nor U10763 (N_10763,N_9079,N_9308);
or U10764 (N_10764,N_9649,N_9942);
and U10765 (N_10765,N_9121,N_9900);
xor U10766 (N_10766,N_9317,N_9903);
nor U10767 (N_10767,N_9315,N_9113);
xnor U10768 (N_10768,N_9610,N_9650);
nor U10769 (N_10769,N_9052,N_9924);
nand U10770 (N_10770,N_9686,N_9017);
and U10771 (N_10771,N_9180,N_9259);
or U10772 (N_10772,N_9681,N_9065);
nand U10773 (N_10773,N_9596,N_9073);
or U10774 (N_10774,N_9884,N_9846);
and U10775 (N_10775,N_9894,N_9202);
and U10776 (N_10776,N_9680,N_9217);
nor U10777 (N_10777,N_9686,N_9233);
nand U10778 (N_10778,N_9588,N_9374);
or U10779 (N_10779,N_9240,N_9674);
and U10780 (N_10780,N_9391,N_9103);
nand U10781 (N_10781,N_9764,N_9528);
or U10782 (N_10782,N_9427,N_9589);
and U10783 (N_10783,N_9386,N_9150);
or U10784 (N_10784,N_9675,N_9753);
xnor U10785 (N_10785,N_9962,N_9447);
xor U10786 (N_10786,N_9936,N_9620);
nor U10787 (N_10787,N_9590,N_9942);
nor U10788 (N_10788,N_9256,N_9539);
nand U10789 (N_10789,N_9864,N_9059);
and U10790 (N_10790,N_9878,N_9614);
xor U10791 (N_10791,N_9225,N_9034);
xnor U10792 (N_10792,N_9172,N_9988);
nand U10793 (N_10793,N_9378,N_9073);
xnor U10794 (N_10794,N_9719,N_9024);
nor U10795 (N_10795,N_9685,N_9605);
xor U10796 (N_10796,N_9636,N_9520);
nor U10797 (N_10797,N_9895,N_9683);
nand U10798 (N_10798,N_9531,N_9326);
or U10799 (N_10799,N_9234,N_9457);
or U10800 (N_10800,N_9289,N_9693);
and U10801 (N_10801,N_9109,N_9853);
and U10802 (N_10802,N_9006,N_9615);
or U10803 (N_10803,N_9636,N_9568);
nand U10804 (N_10804,N_9610,N_9371);
xor U10805 (N_10805,N_9098,N_9298);
xor U10806 (N_10806,N_9980,N_9211);
nor U10807 (N_10807,N_9512,N_9385);
xor U10808 (N_10808,N_9080,N_9805);
nand U10809 (N_10809,N_9857,N_9278);
or U10810 (N_10810,N_9753,N_9400);
nand U10811 (N_10811,N_9960,N_9577);
or U10812 (N_10812,N_9255,N_9675);
or U10813 (N_10813,N_9046,N_9789);
nand U10814 (N_10814,N_9622,N_9075);
xor U10815 (N_10815,N_9466,N_9838);
or U10816 (N_10816,N_9528,N_9769);
xnor U10817 (N_10817,N_9384,N_9095);
xor U10818 (N_10818,N_9164,N_9013);
nor U10819 (N_10819,N_9154,N_9806);
nand U10820 (N_10820,N_9373,N_9328);
nand U10821 (N_10821,N_9919,N_9424);
and U10822 (N_10822,N_9868,N_9730);
xor U10823 (N_10823,N_9762,N_9136);
nor U10824 (N_10824,N_9078,N_9130);
xor U10825 (N_10825,N_9019,N_9749);
nand U10826 (N_10826,N_9288,N_9944);
nand U10827 (N_10827,N_9319,N_9999);
nor U10828 (N_10828,N_9508,N_9967);
xor U10829 (N_10829,N_9205,N_9464);
nand U10830 (N_10830,N_9748,N_9636);
nand U10831 (N_10831,N_9808,N_9687);
xnor U10832 (N_10832,N_9776,N_9536);
or U10833 (N_10833,N_9330,N_9689);
nand U10834 (N_10834,N_9676,N_9383);
nor U10835 (N_10835,N_9770,N_9458);
or U10836 (N_10836,N_9391,N_9186);
xor U10837 (N_10837,N_9027,N_9967);
or U10838 (N_10838,N_9391,N_9591);
nor U10839 (N_10839,N_9629,N_9433);
or U10840 (N_10840,N_9214,N_9365);
nand U10841 (N_10841,N_9678,N_9507);
nand U10842 (N_10842,N_9805,N_9419);
and U10843 (N_10843,N_9259,N_9086);
nor U10844 (N_10844,N_9075,N_9961);
nor U10845 (N_10845,N_9586,N_9155);
or U10846 (N_10846,N_9671,N_9754);
nand U10847 (N_10847,N_9918,N_9721);
nand U10848 (N_10848,N_9687,N_9415);
nor U10849 (N_10849,N_9566,N_9847);
or U10850 (N_10850,N_9283,N_9863);
nand U10851 (N_10851,N_9895,N_9224);
or U10852 (N_10852,N_9293,N_9877);
and U10853 (N_10853,N_9022,N_9820);
xor U10854 (N_10854,N_9281,N_9037);
xnor U10855 (N_10855,N_9326,N_9933);
or U10856 (N_10856,N_9857,N_9397);
or U10857 (N_10857,N_9544,N_9677);
or U10858 (N_10858,N_9708,N_9925);
nand U10859 (N_10859,N_9692,N_9262);
or U10860 (N_10860,N_9328,N_9977);
and U10861 (N_10861,N_9617,N_9856);
or U10862 (N_10862,N_9963,N_9976);
or U10863 (N_10863,N_9659,N_9549);
nand U10864 (N_10864,N_9095,N_9967);
or U10865 (N_10865,N_9337,N_9518);
nor U10866 (N_10866,N_9299,N_9610);
nand U10867 (N_10867,N_9032,N_9434);
nand U10868 (N_10868,N_9630,N_9890);
nor U10869 (N_10869,N_9212,N_9234);
nand U10870 (N_10870,N_9553,N_9549);
and U10871 (N_10871,N_9628,N_9936);
nor U10872 (N_10872,N_9415,N_9068);
and U10873 (N_10873,N_9249,N_9135);
and U10874 (N_10874,N_9503,N_9193);
and U10875 (N_10875,N_9397,N_9746);
nor U10876 (N_10876,N_9107,N_9054);
xor U10877 (N_10877,N_9821,N_9393);
and U10878 (N_10878,N_9883,N_9351);
xnor U10879 (N_10879,N_9629,N_9144);
xnor U10880 (N_10880,N_9712,N_9585);
nor U10881 (N_10881,N_9853,N_9547);
xnor U10882 (N_10882,N_9951,N_9220);
nor U10883 (N_10883,N_9556,N_9438);
or U10884 (N_10884,N_9169,N_9863);
nor U10885 (N_10885,N_9043,N_9055);
xor U10886 (N_10886,N_9222,N_9496);
and U10887 (N_10887,N_9702,N_9548);
nand U10888 (N_10888,N_9154,N_9386);
or U10889 (N_10889,N_9021,N_9951);
and U10890 (N_10890,N_9209,N_9022);
or U10891 (N_10891,N_9182,N_9419);
nand U10892 (N_10892,N_9194,N_9395);
nand U10893 (N_10893,N_9418,N_9210);
nor U10894 (N_10894,N_9381,N_9170);
xor U10895 (N_10895,N_9781,N_9065);
and U10896 (N_10896,N_9056,N_9994);
nor U10897 (N_10897,N_9285,N_9575);
and U10898 (N_10898,N_9330,N_9376);
or U10899 (N_10899,N_9031,N_9741);
nand U10900 (N_10900,N_9705,N_9810);
nand U10901 (N_10901,N_9727,N_9192);
xor U10902 (N_10902,N_9528,N_9834);
nor U10903 (N_10903,N_9377,N_9587);
or U10904 (N_10904,N_9608,N_9409);
and U10905 (N_10905,N_9304,N_9649);
xnor U10906 (N_10906,N_9383,N_9752);
xnor U10907 (N_10907,N_9967,N_9740);
nor U10908 (N_10908,N_9457,N_9366);
or U10909 (N_10909,N_9357,N_9226);
nor U10910 (N_10910,N_9691,N_9898);
nor U10911 (N_10911,N_9056,N_9967);
and U10912 (N_10912,N_9194,N_9359);
xnor U10913 (N_10913,N_9142,N_9919);
nor U10914 (N_10914,N_9056,N_9284);
or U10915 (N_10915,N_9300,N_9125);
nor U10916 (N_10916,N_9951,N_9770);
and U10917 (N_10917,N_9798,N_9795);
xor U10918 (N_10918,N_9259,N_9310);
nand U10919 (N_10919,N_9578,N_9611);
nor U10920 (N_10920,N_9926,N_9743);
or U10921 (N_10921,N_9403,N_9301);
xnor U10922 (N_10922,N_9772,N_9143);
and U10923 (N_10923,N_9640,N_9302);
nand U10924 (N_10924,N_9621,N_9526);
nor U10925 (N_10925,N_9187,N_9518);
xnor U10926 (N_10926,N_9841,N_9908);
nor U10927 (N_10927,N_9297,N_9319);
or U10928 (N_10928,N_9917,N_9650);
nand U10929 (N_10929,N_9083,N_9100);
and U10930 (N_10930,N_9554,N_9105);
xnor U10931 (N_10931,N_9872,N_9248);
nor U10932 (N_10932,N_9395,N_9549);
nand U10933 (N_10933,N_9496,N_9517);
or U10934 (N_10934,N_9639,N_9839);
or U10935 (N_10935,N_9241,N_9887);
and U10936 (N_10936,N_9709,N_9862);
xor U10937 (N_10937,N_9235,N_9379);
nand U10938 (N_10938,N_9787,N_9198);
nand U10939 (N_10939,N_9211,N_9812);
xnor U10940 (N_10940,N_9372,N_9781);
or U10941 (N_10941,N_9245,N_9086);
nor U10942 (N_10942,N_9275,N_9479);
nor U10943 (N_10943,N_9605,N_9859);
xnor U10944 (N_10944,N_9239,N_9706);
nor U10945 (N_10945,N_9920,N_9989);
nand U10946 (N_10946,N_9449,N_9080);
xnor U10947 (N_10947,N_9161,N_9727);
and U10948 (N_10948,N_9144,N_9522);
or U10949 (N_10949,N_9919,N_9682);
xor U10950 (N_10950,N_9870,N_9935);
nor U10951 (N_10951,N_9906,N_9193);
and U10952 (N_10952,N_9123,N_9431);
nor U10953 (N_10953,N_9933,N_9042);
nand U10954 (N_10954,N_9172,N_9012);
and U10955 (N_10955,N_9771,N_9759);
nand U10956 (N_10956,N_9892,N_9212);
nand U10957 (N_10957,N_9314,N_9281);
or U10958 (N_10958,N_9918,N_9472);
nor U10959 (N_10959,N_9167,N_9330);
xor U10960 (N_10960,N_9477,N_9676);
nand U10961 (N_10961,N_9511,N_9211);
xnor U10962 (N_10962,N_9213,N_9207);
or U10963 (N_10963,N_9355,N_9360);
xnor U10964 (N_10964,N_9442,N_9367);
nor U10965 (N_10965,N_9204,N_9669);
or U10966 (N_10966,N_9132,N_9370);
nand U10967 (N_10967,N_9988,N_9826);
xnor U10968 (N_10968,N_9419,N_9587);
xor U10969 (N_10969,N_9249,N_9906);
or U10970 (N_10970,N_9160,N_9557);
and U10971 (N_10971,N_9306,N_9091);
and U10972 (N_10972,N_9474,N_9295);
xor U10973 (N_10973,N_9095,N_9679);
or U10974 (N_10974,N_9425,N_9682);
or U10975 (N_10975,N_9275,N_9268);
or U10976 (N_10976,N_9484,N_9111);
and U10977 (N_10977,N_9012,N_9257);
nand U10978 (N_10978,N_9820,N_9673);
and U10979 (N_10979,N_9279,N_9847);
nor U10980 (N_10980,N_9010,N_9966);
xor U10981 (N_10981,N_9919,N_9870);
or U10982 (N_10982,N_9060,N_9255);
xnor U10983 (N_10983,N_9569,N_9050);
xor U10984 (N_10984,N_9857,N_9794);
and U10985 (N_10985,N_9690,N_9011);
xor U10986 (N_10986,N_9039,N_9647);
nor U10987 (N_10987,N_9355,N_9528);
xnor U10988 (N_10988,N_9391,N_9646);
nand U10989 (N_10989,N_9872,N_9919);
and U10990 (N_10990,N_9150,N_9262);
xnor U10991 (N_10991,N_9985,N_9489);
and U10992 (N_10992,N_9768,N_9187);
nor U10993 (N_10993,N_9781,N_9603);
or U10994 (N_10994,N_9510,N_9630);
nand U10995 (N_10995,N_9329,N_9112);
and U10996 (N_10996,N_9945,N_9673);
and U10997 (N_10997,N_9479,N_9086);
and U10998 (N_10998,N_9021,N_9137);
and U10999 (N_10999,N_9235,N_9647);
xor U11000 (N_11000,N_10844,N_10155);
or U11001 (N_11001,N_10629,N_10433);
nand U11002 (N_11002,N_10478,N_10733);
nor U11003 (N_11003,N_10590,N_10619);
and U11004 (N_11004,N_10896,N_10525);
xnor U11005 (N_11005,N_10931,N_10225);
or U11006 (N_11006,N_10543,N_10819);
or U11007 (N_11007,N_10982,N_10820);
nor U11008 (N_11008,N_10517,N_10624);
or U11009 (N_11009,N_10273,N_10279);
nand U11010 (N_11010,N_10384,N_10388);
nor U11011 (N_11011,N_10675,N_10887);
or U11012 (N_11012,N_10937,N_10008);
or U11013 (N_11013,N_10255,N_10642);
xor U11014 (N_11014,N_10371,N_10337);
nor U11015 (N_11015,N_10065,N_10060);
or U11016 (N_11016,N_10266,N_10278);
and U11017 (N_11017,N_10929,N_10934);
nand U11018 (N_11018,N_10913,N_10342);
and U11019 (N_11019,N_10951,N_10545);
xnor U11020 (N_11020,N_10723,N_10295);
nor U11021 (N_11021,N_10021,N_10565);
or U11022 (N_11022,N_10980,N_10506);
xnor U11023 (N_11023,N_10219,N_10217);
xnor U11024 (N_11024,N_10987,N_10585);
nand U11025 (N_11025,N_10183,N_10960);
nand U11026 (N_11026,N_10835,N_10631);
nor U11027 (N_11027,N_10877,N_10370);
xor U11028 (N_11028,N_10632,N_10664);
nor U11029 (N_11029,N_10808,N_10591);
nand U11030 (N_11030,N_10976,N_10330);
nand U11031 (N_11031,N_10326,N_10275);
and U11032 (N_11032,N_10159,N_10638);
xor U11033 (N_11033,N_10407,N_10324);
or U11034 (N_11034,N_10164,N_10564);
or U11035 (N_11035,N_10571,N_10686);
or U11036 (N_11036,N_10837,N_10623);
nand U11037 (N_11037,N_10464,N_10730);
nand U11038 (N_11038,N_10666,N_10191);
and U11039 (N_11039,N_10607,N_10173);
xnor U11040 (N_11040,N_10716,N_10169);
xnor U11041 (N_11041,N_10651,N_10568);
nand U11042 (N_11042,N_10160,N_10542);
nand U11043 (N_11043,N_10296,N_10643);
and U11044 (N_11044,N_10910,N_10866);
or U11045 (N_11045,N_10802,N_10030);
or U11046 (N_11046,N_10510,N_10452);
and U11047 (N_11047,N_10298,N_10272);
and U11048 (N_11048,N_10769,N_10831);
xor U11049 (N_11049,N_10434,N_10046);
nand U11050 (N_11050,N_10778,N_10577);
nor U11051 (N_11051,N_10840,N_10036);
nand U11052 (N_11052,N_10810,N_10582);
or U11053 (N_11053,N_10446,N_10906);
or U11054 (N_11054,N_10772,N_10578);
xnor U11055 (N_11055,N_10075,N_10395);
or U11056 (N_11056,N_10533,N_10277);
and U11057 (N_11057,N_10637,N_10768);
xnor U11058 (N_11058,N_10989,N_10941);
nor U11059 (N_11059,N_10552,N_10396);
or U11060 (N_11060,N_10703,N_10226);
and U11061 (N_11061,N_10824,N_10660);
xor U11062 (N_11062,N_10974,N_10421);
nand U11063 (N_11063,N_10857,N_10055);
nor U11064 (N_11064,N_10812,N_10059);
xor U11065 (N_11065,N_10293,N_10676);
and U11066 (N_11066,N_10107,N_10181);
nor U11067 (N_11067,N_10064,N_10770);
nand U11068 (N_11068,N_10786,N_10015);
or U11069 (N_11069,N_10102,N_10701);
xor U11070 (N_11070,N_10400,N_10507);
or U11071 (N_11071,N_10113,N_10265);
nor U11072 (N_11072,N_10357,N_10628);
or U11073 (N_11073,N_10302,N_10054);
or U11074 (N_11074,N_10860,N_10430);
nor U11075 (N_11075,N_10214,N_10815);
or U11076 (N_11076,N_10520,N_10901);
xor U11077 (N_11077,N_10926,N_10668);
xnor U11078 (N_11078,N_10161,N_10473);
nand U11079 (N_11079,N_10805,N_10086);
or U11080 (N_11080,N_10244,N_10366);
or U11081 (N_11081,N_10340,N_10771);
or U11082 (N_11082,N_10401,N_10750);
and U11083 (N_11083,N_10163,N_10080);
nor U11084 (N_11084,N_10853,N_10609);
nor U11085 (N_11085,N_10353,N_10119);
nor U11086 (N_11086,N_10954,N_10338);
xor U11087 (N_11087,N_10882,N_10438);
or U11088 (N_11088,N_10476,N_10232);
nor U11089 (N_11089,N_10014,N_10618);
nor U11090 (N_11090,N_10177,N_10634);
xor U11091 (N_11091,N_10462,N_10082);
nor U11092 (N_11092,N_10763,N_10515);
nor U11093 (N_11093,N_10207,N_10202);
nor U11094 (N_11094,N_10404,N_10774);
nand U11095 (N_11095,N_10873,N_10678);
and U11096 (N_11096,N_10540,N_10408);
nand U11097 (N_11097,N_10653,N_10461);
xnor U11098 (N_11098,N_10000,N_10953);
or U11099 (N_11099,N_10459,N_10697);
nand U11100 (N_11100,N_10004,N_10372);
nor U11101 (N_11101,N_10007,N_10304);
nand U11102 (N_11102,N_10363,N_10997);
or U11103 (N_11103,N_10672,N_10792);
nand U11104 (N_11104,N_10373,N_10549);
or U11105 (N_11105,N_10123,N_10416);
and U11106 (N_11106,N_10178,N_10383);
nor U11107 (N_11107,N_10814,N_10253);
nand U11108 (N_11108,N_10496,N_10442);
or U11109 (N_11109,N_10908,N_10696);
or U11110 (N_11110,N_10156,N_10635);
or U11111 (N_11111,N_10988,N_10174);
nor U11112 (N_11112,N_10871,N_10816);
nor U11113 (N_11113,N_10482,N_10185);
nand U11114 (N_11114,N_10091,N_10310);
xnor U11115 (N_11115,N_10912,N_10600);
nor U11116 (N_11116,N_10027,N_10131);
nor U11117 (N_11117,N_10876,N_10024);
nor U11118 (N_11118,N_10268,N_10503);
and U11119 (N_11119,N_10621,N_10115);
xnor U11120 (N_11120,N_10405,N_10789);
and U11121 (N_11121,N_10700,N_10248);
nor U11122 (N_11122,N_10579,N_10151);
nand U11123 (N_11123,N_10572,N_10811);
nand U11124 (N_11124,N_10237,N_10134);
or U11125 (N_11125,N_10299,N_10186);
and U11126 (N_11126,N_10252,N_10677);
xnor U11127 (N_11127,N_10133,N_10331);
nor U11128 (N_11128,N_10426,N_10335);
nor U11129 (N_11129,N_10254,N_10785);
or U11130 (N_11130,N_10041,N_10345);
nor U11131 (N_11131,N_10247,N_10606);
and U11132 (N_11132,N_10058,N_10414);
nand U11133 (N_11133,N_10221,N_10449);
and U11134 (N_11134,N_10198,N_10106);
xor U11135 (N_11135,N_10402,N_10881);
nand U11136 (N_11136,N_10839,N_10754);
xor U11137 (N_11137,N_10625,N_10052);
xor U11138 (N_11138,N_10524,N_10016);
or U11139 (N_11139,N_10467,N_10380);
nor U11140 (N_11140,N_10514,N_10137);
xnor U11141 (N_11141,N_10386,N_10270);
xor U11142 (N_11142,N_10604,N_10350);
or U11143 (N_11143,N_10967,N_10243);
xnor U11144 (N_11144,N_10130,N_10508);
and U11145 (N_11145,N_10787,N_10559);
nor U11146 (N_11146,N_10339,N_10294);
nor U11147 (N_11147,N_10368,N_10587);
or U11148 (N_11148,N_10627,N_10708);
and U11149 (N_11149,N_10895,N_10126);
or U11150 (N_11150,N_10419,N_10048);
or U11151 (N_11151,N_10576,N_10020);
or U11152 (N_11152,N_10229,N_10705);
nand U11153 (N_11153,N_10317,N_10072);
nand U11154 (N_11154,N_10842,N_10961);
or U11155 (N_11155,N_10109,N_10532);
or U11156 (N_11156,N_10586,N_10209);
xnor U11157 (N_11157,N_10238,N_10135);
nand U11158 (N_11158,N_10655,N_10965);
and U11159 (N_11159,N_10403,N_10028);
nor U11160 (N_11160,N_10479,N_10352);
nand U11161 (N_11161,N_10658,N_10736);
or U11162 (N_11162,N_10610,N_10818);
nand U11163 (N_11163,N_10759,N_10474);
or U11164 (N_11164,N_10725,N_10746);
nand U11165 (N_11165,N_10829,N_10611);
xnor U11166 (N_11166,N_10788,N_10732);
and U11167 (N_11167,N_10307,N_10136);
nor U11168 (N_11168,N_10722,N_10475);
or U11169 (N_11169,N_10040,N_10715);
xnor U11170 (N_11170,N_10071,N_10455);
nor U11171 (N_11171,N_10468,N_10749);
and U11172 (N_11172,N_10051,N_10779);
nor U11173 (N_11173,N_10833,N_10985);
nor U11174 (N_11174,N_10349,N_10448);
and U11175 (N_11175,N_10504,N_10859);
and U11176 (N_11176,N_10488,N_10240);
or U11177 (N_11177,N_10923,N_10096);
nor U11178 (N_11178,N_10344,N_10555);
xor U11179 (N_11179,N_10612,N_10952);
nor U11180 (N_11180,N_10614,N_10261);
and U11181 (N_11181,N_10494,N_10827);
nand U11182 (N_11182,N_10035,N_10850);
or U11183 (N_11183,N_10673,N_10057);
or U11184 (N_11184,N_10063,N_10088);
nor U11185 (N_11185,N_10918,N_10129);
nor U11186 (N_11186,N_10681,N_10470);
or U11187 (N_11187,N_10146,N_10043);
nand U11188 (N_11188,N_10535,N_10728);
and U11189 (N_11189,N_10153,N_10726);
and U11190 (N_11190,N_10547,N_10132);
and U11191 (N_11191,N_10704,N_10143);
nand U11192 (N_11192,N_10457,N_10190);
and U11193 (N_11193,N_10224,N_10721);
nor U11194 (N_11194,N_10499,N_10731);
nand U11195 (N_11195,N_10199,N_10592);
xnor U11196 (N_11196,N_10879,N_10411);
nor U11197 (N_11197,N_10200,N_10394);
xor U11198 (N_11198,N_10147,N_10447);
or U11199 (N_11199,N_10083,N_10530);
and U11200 (N_11200,N_10925,N_10561);
and U11201 (N_11201,N_10907,N_10581);
and U11202 (N_11202,N_10546,N_10188);
and U11203 (N_11203,N_10359,N_10356);
or U11204 (N_11204,N_10935,N_10258);
and U11205 (N_11205,N_10099,N_10256);
nand U11206 (N_11206,N_10617,N_10795);
or U11207 (N_11207,N_10847,N_10919);
nand U11208 (N_11208,N_10999,N_10699);
nor U11209 (N_11209,N_10662,N_10365);
nor U11210 (N_11210,N_10720,N_10215);
nor U11211 (N_11211,N_10593,N_10195);
nand U11212 (N_11212,N_10886,N_10874);
or U11213 (N_11213,N_10836,N_10179);
nand U11214 (N_11214,N_10897,N_10456);
nand U11215 (N_11215,N_10117,N_10392);
or U11216 (N_11216,N_10242,N_10813);
xnor U11217 (N_11217,N_10529,N_10724);
and U11218 (N_11218,N_10290,N_10991);
xor U11219 (N_11219,N_10927,N_10501);
nor U11220 (N_11220,N_10127,N_10103);
or U11221 (N_11221,N_10996,N_10553);
nor U11222 (N_11222,N_10116,N_10741);
nand U11223 (N_11223,N_10595,N_10271);
xnor U11224 (N_11224,N_10782,N_10206);
xor U11225 (N_11225,N_10740,N_10427);
nor U11226 (N_11226,N_10230,N_10005);
nand U11227 (N_11227,N_10431,N_10804);
and U11228 (N_11228,N_10981,N_10570);
and U11229 (N_11229,N_10544,N_10009);
or U11230 (N_11230,N_10262,N_10484);
or U11231 (N_11231,N_10930,N_10320);
nor U11232 (N_11232,N_10167,N_10626);
xnor U11233 (N_11233,N_10880,N_10846);
nor U11234 (N_11234,N_10321,N_10241);
and U11235 (N_11235,N_10745,N_10502);
xnor U11236 (N_11236,N_10114,N_10914);
or U11237 (N_11237,N_10718,N_10825);
nor U11238 (N_11238,N_10640,N_10087);
nor U11239 (N_11239,N_10776,N_10001);
nor U11240 (N_11240,N_10758,N_10081);
or U11241 (N_11241,N_10233,N_10061);
xor U11242 (N_11242,N_10432,N_10712);
xor U11243 (N_11243,N_10674,N_10026);
nand U11244 (N_11244,N_10693,N_10076);
xnor U11245 (N_11245,N_10382,N_10193);
nand U11246 (N_11246,N_10560,N_10223);
nor U11247 (N_11247,N_10947,N_10276);
or U11248 (N_11248,N_10867,N_10212);
nand U11249 (N_11249,N_10070,N_10092);
xnor U11250 (N_11250,N_10334,N_10305);
nor U11251 (N_11251,N_10713,N_10379);
nand U11252 (N_11252,N_10033,N_10319);
xor U11253 (N_11253,N_10019,N_10841);
nor U11254 (N_11254,N_10869,N_10097);
nor U11255 (N_11255,N_10111,N_10870);
or U11256 (N_11256,N_10493,N_10894);
and U11257 (N_11257,N_10729,N_10390);
or U11258 (N_11258,N_10429,N_10936);
nand U11259 (N_11259,N_10291,N_10616);
nand U11260 (N_11260,N_10053,N_10955);
and U11261 (N_11261,N_10584,N_10773);
and U11262 (N_11262,N_10142,N_10239);
xor U11263 (N_11263,N_10671,N_10231);
xnor U11264 (N_11264,N_10002,N_10781);
xnor U11265 (N_11265,N_10393,N_10848);
xor U11266 (N_11266,N_10037,N_10978);
or U11267 (N_11267,N_10205,N_10343);
xnor U11268 (N_11268,N_10039,N_10667);
xor U11269 (N_11269,N_10184,N_10050);
or U11270 (N_11270,N_10605,N_10192);
nand U11271 (N_11271,N_10957,N_10670);
nor U11272 (N_11272,N_10491,N_10306);
xor U11273 (N_11273,N_10665,N_10645);
nor U11274 (N_11274,N_10641,N_10523);
xor U11275 (N_11275,N_10888,N_10854);
nand U11276 (N_11276,N_10398,N_10423);
xor U11277 (N_11277,N_10211,N_10717);
and U11278 (N_11278,N_10257,N_10216);
or U11279 (N_11279,N_10264,N_10527);
nand U11280 (N_11280,N_10329,N_10562);
nor U11281 (N_11281,N_10639,N_10045);
nor U11282 (N_11282,N_10068,N_10790);
xor U11283 (N_11283,N_10924,N_10358);
xnor U11284 (N_11284,N_10367,N_10056);
nand U11285 (N_11285,N_10596,N_10783);
or U11286 (N_11286,N_10702,N_10694);
nand U11287 (N_11287,N_10236,N_10110);
xnor U11288 (N_11288,N_10902,N_10049);
or U11289 (N_11289,N_10916,N_10748);
or U11290 (N_11290,N_10922,N_10399);
xnor U11291 (N_11291,N_10436,N_10148);
nor U11292 (N_11292,N_10509,N_10450);
or U11293 (N_11293,N_10558,N_10010);
nor U11294 (N_11294,N_10968,N_10743);
xor U11295 (N_11295,N_10100,N_10417);
or U11296 (N_11296,N_10485,N_10511);
and U11297 (N_11297,N_10453,N_10439);
or U11298 (N_11298,N_10798,N_10312);
or U11299 (N_11299,N_10554,N_10682);
and U11300 (N_11300,N_10636,N_10139);
xnor U11301 (N_11301,N_10706,N_10118);
nor U11302 (N_11302,N_10864,N_10522);
and U11303 (N_11303,N_10044,N_10830);
nor U11304 (N_11304,N_10196,N_10737);
nand U11305 (N_11305,N_10300,N_10656);
xnor U11306 (N_11306,N_10471,N_10128);
nor U11307 (N_11307,N_10140,N_10917);
or U11308 (N_11308,N_10104,N_10280);
nand U11309 (N_11309,N_10851,N_10249);
and U11310 (N_11310,N_10537,N_10998);
and U11311 (N_11311,N_10679,N_10424);
xor U11312 (N_11312,N_10435,N_10466);
and U11313 (N_11313,N_10495,N_10176);
and U11314 (N_11314,N_10066,N_10852);
nor U11315 (N_11315,N_10751,N_10440);
or U11316 (N_11316,N_10101,N_10210);
nor U11317 (N_11317,N_10865,N_10784);
nand U11318 (N_11318,N_10316,N_10539);
or U11319 (N_11319,N_10943,N_10903);
and U11320 (N_11320,N_10227,N_10369);
or U11321 (N_11321,N_10890,N_10441);
xnor U11322 (N_11322,N_10172,N_10757);
nand U11323 (N_11323,N_10480,N_10165);
xor U11324 (N_11324,N_10397,N_10516);
and U11325 (N_11325,N_10622,N_10284);
nor U11326 (N_11326,N_10806,N_10940);
or U11327 (N_11327,N_10719,N_10166);
nand U11328 (N_11328,N_10287,N_10422);
nand U11329 (N_11329,N_10460,N_10972);
nand U11330 (N_11330,N_10566,N_10003);
xnor U11331 (N_11331,N_10801,N_10067);
or U11332 (N_11332,N_10822,N_10078);
nand U11333 (N_11333,N_10282,N_10807);
and U11334 (N_11334,N_10993,N_10269);
or U11335 (N_11335,N_10698,N_10351);
nor U11336 (N_11336,N_10695,N_10898);
and U11337 (N_11337,N_10410,N_10597);
xnor U11338 (N_11338,N_10767,N_10197);
xor U11339 (N_11339,N_10531,N_10328);
nand U11340 (N_11340,N_10283,N_10762);
xnor U11341 (N_11341,N_10093,N_10025);
xor U11342 (N_11342,N_10332,N_10512);
nand U11343 (N_11343,N_10158,N_10311);
nand U11344 (N_11344,N_10012,N_10680);
or U11345 (N_11345,N_10038,N_10428);
nand U11346 (N_11346,N_10376,N_10444);
nand U11347 (N_11347,N_10228,N_10187);
and U11348 (N_11348,N_10654,N_10800);
nand U11349 (N_11349,N_10138,N_10944);
nand U11350 (N_11350,N_10950,N_10029);
nand U11351 (N_11351,N_10883,N_10661);
nor U11352 (N_11352,N_10855,N_10569);
or U11353 (N_11353,N_10309,N_10753);
nand U11354 (N_11354,N_10928,N_10498);
nand U11355 (N_11355,N_10990,N_10084);
nand U11356 (N_11356,N_10420,N_10125);
xor U11357 (N_11357,N_10690,N_10201);
and U11358 (N_11358,N_10970,N_10152);
and U11359 (N_11359,N_10220,N_10023);
and U11360 (N_11360,N_10477,N_10218);
or U11361 (N_11361,N_10175,N_10945);
and U11362 (N_11362,N_10251,N_10465);
nand U11363 (N_11363,N_10599,N_10245);
xor U11364 (N_11364,N_10747,N_10031);
nand U11365 (N_11365,N_10355,N_10964);
or U11366 (N_11366,N_10451,N_10189);
and U11367 (N_11367,N_10022,N_10878);
nand U11368 (N_11368,N_10872,N_10630);
xnor U11369 (N_11369,N_10490,N_10834);
or U11370 (N_11370,N_10891,N_10354);
nor U11371 (N_11371,N_10443,N_10803);
nand U11372 (N_11372,N_10322,N_10760);
nand U11373 (N_11373,N_10500,N_10683);
nor U11374 (N_11374,N_10650,N_10689);
xor U11375 (N_11375,N_10588,N_10687);
xnor U11376 (N_11376,N_10979,N_10647);
and U11377 (N_11377,N_10378,N_10594);
xor U11378 (N_11378,N_10018,N_10203);
or U11379 (N_11379,N_10374,N_10141);
nand U11380 (N_11380,N_10845,N_10652);
nor U11381 (N_11381,N_10095,N_10727);
and U11382 (N_11382,N_10108,N_10958);
xnor U11383 (N_11383,N_10691,N_10971);
or U11384 (N_11384,N_10303,N_10911);
and U11385 (N_11385,N_10333,N_10905);
nand U11386 (N_11386,N_10208,N_10263);
xor U11387 (N_11387,N_10863,N_10323);
nand U11388 (N_11388,N_10124,N_10246);
nor U11389 (N_11389,N_10885,N_10856);
nor U11390 (N_11390,N_10613,N_10889);
and U11391 (N_11391,N_10992,N_10412);
or U11392 (N_11392,N_10222,N_10315);
nand U11393 (N_11393,N_10764,N_10437);
xor U11394 (N_11394,N_10487,N_10973);
and U11395 (N_11395,N_10893,N_10458);
nand U11396 (N_11396,N_10013,N_10550);
nand U11397 (N_11397,N_10168,N_10289);
nor U11398 (N_11398,N_10809,N_10977);
and U11399 (N_11399,N_10821,N_10521);
xor U11400 (N_11400,N_10548,N_10659);
and U11401 (N_11401,N_10826,N_10062);
and U11402 (N_11402,N_10144,N_10793);
nand U11403 (N_11403,N_10341,N_10346);
or U11404 (N_11404,N_10649,N_10170);
xnor U11405 (N_11405,N_10085,N_10995);
xnor U11406 (N_11406,N_10994,N_10551);
and U11407 (N_11407,N_10047,N_10946);
nor U11408 (N_11408,N_10949,N_10418);
xor U11409 (N_11409,N_10094,N_10098);
and U11410 (N_11410,N_10939,N_10154);
xor U11411 (N_11411,N_10348,N_10361);
xor U11412 (N_11412,N_10513,N_10489);
nor U11413 (N_11413,N_10285,N_10556);
and U11414 (N_11414,N_10909,N_10526);
nand U11415 (N_11415,N_10259,N_10648);
xnor U11416 (N_11416,N_10112,N_10608);
or U11417 (N_11417,N_10381,N_10391);
nand U11418 (N_11418,N_10387,N_10744);
nand U11419 (N_11419,N_10603,N_10445);
or U11420 (N_11420,N_10986,N_10286);
or U11421 (N_11421,N_10120,N_10794);
or U11422 (N_11422,N_10297,N_10375);
xor U11423 (N_11423,N_10011,N_10235);
nand U11424 (N_11424,N_10042,N_10090);
nand U11425 (N_11425,N_10413,N_10580);
nand U11426 (N_11426,N_10145,N_10620);
nand U11427 (N_11427,N_10574,N_10079);
xnor U11428 (N_11428,N_10360,N_10862);
nor U11429 (N_11429,N_10069,N_10074);
and U11430 (N_11430,N_10663,N_10267);
nor U11431 (N_11431,N_10861,N_10884);
or U11432 (N_11432,N_10557,N_10150);
xnor U11433 (N_11433,N_10709,N_10260);
xnor U11434 (N_11434,N_10921,N_10959);
nor U11435 (N_11435,N_10377,N_10541);
nor U11436 (N_11436,N_10105,N_10646);
nand U11437 (N_11437,N_10969,N_10162);
or U11438 (N_11438,N_10077,N_10347);
nor U11439 (N_11439,N_10528,N_10314);
nor U11440 (N_11440,N_10032,N_10644);
and U11441 (N_11441,N_10336,N_10932);
nor U11442 (N_11442,N_10755,N_10017);
or U11443 (N_11443,N_10707,N_10602);
and U11444 (N_11444,N_10006,N_10318);
and U11445 (N_11445,N_10797,N_10288);
nor U11446 (N_11446,N_10313,N_10389);
nand U11447 (N_11447,N_10121,N_10601);
or U11448 (N_11448,N_10325,N_10984);
and U11449 (N_11449,N_10975,N_10832);
nor U11450 (N_11450,N_10963,N_10292);
nor U11451 (N_11451,N_10274,N_10875);
nand U11452 (N_11452,N_10734,N_10122);
nor U11453 (N_11453,N_10633,N_10583);
xnor U11454 (N_11454,N_10684,N_10838);
xnor U11455 (N_11455,N_10669,N_10454);
xnor U11456 (N_11456,N_10739,N_10756);
and U11457 (N_11457,N_10519,N_10234);
nand U11458 (N_11458,N_10796,N_10481);
nor U11459 (N_11459,N_10688,N_10791);
nand U11460 (N_11460,N_10904,N_10308);
nand U11461 (N_11461,N_10892,N_10765);
and U11462 (N_11462,N_10573,N_10171);
nor U11463 (N_11463,N_10948,N_10505);
or U11464 (N_11464,N_10899,N_10657);
and U11465 (N_11465,N_10942,N_10180);
nor U11466 (N_11466,N_10538,N_10149);
nor U11467 (N_11467,N_10563,N_10843);
xor U11468 (N_11468,N_10766,N_10472);
xor U11469 (N_11469,N_10777,N_10799);
nand U11470 (N_11470,N_10589,N_10281);
nand U11471 (N_11471,N_10685,N_10483);
nand U11472 (N_11472,N_10486,N_10327);
or U11473 (N_11473,N_10497,N_10536);
nor U11474 (N_11474,N_10567,N_10933);
nor U11475 (N_11475,N_10752,N_10735);
and U11476 (N_11476,N_10817,N_10364);
or U11477 (N_11477,N_10463,N_10409);
nand U11478 (N_11478,N_10469,N_10157);
and U11479 (N_11479,N_10711,N_10089);
or U11480 (N_11480,N_10761,N_10742);
nand U11481 (N_11481,N_10775,N_10966);
xnor U11482 (N_11482,N_10204,N_10575);
xnor U11483 (N_11483,N_10983,N_10250);
or U11484 (N_11484,N_10692,N_10534);
nand U11485 (N_11485,N_10615,N_10182);
or U11486 (N_11486,N_10849,N_10714);
nor U11487 (N_11487,N_10194,N_10710);
nand U11488 (N_11488,N_10868,N_10823);
or U11489 (N_11489,N_10956,N_10780);
xnor U11490 (N_11490,N_10920,N_10598);
nor U11491 (N_11491,N_10828,N_10425);
and U11492 (N_11492,N_10738,N_10385);
nand U11493 (N_11493,N_10962,N_10301);
nor U11494 (N_11494,N_10213,N_10900);
xor U11495 (N_11495,N_10034,N_10858);
and U11496 (N_11496,N_10362,N_10073);
nor U11497 (N_11497,N_10938,N_10492);
and U11498 (N_11498,N_10915,N_10415);
nand U11499 (N_11499,N_10406,N_10518);
xnor U11500 (N_11500,N_10020,N_10890);
and U11501 (N_11501,N_10669,N_10439);
xor U11502 (N_11502,N_10757,N_10937);
and U11503 (N_11503,N_10111,N_10328);
or U11504 (N_11504,N_10350,N_10371);
and U11505 (N_11505,N_10527,N_10366);
xnor U11506 (N_11506,N_10188,N_10200);
and U11507 (N_11507,N_10141,N_10185);
or U11508 (N_11508,N_10849,N_10244);
nand U11509 (N_11509,N_10372,N_10497);
nor U11510 (N_11510,N_10650,N_10752);
and U11511 (N_11511,N_10687,N_10532);
or U11512 (N_11512,N_10263,N_10610);
nand U11513 (N_11513,N_10057,N_10901);
nor U11514 (N_11514,N_10351,N_10902);
and U11515 (N_11515,N_10788,N_10175);
or U11516 (N_11516,N_10156,N_10511);
or U11517 (N_11517,N_10330,N_10729);
or U11518 (N_11518,N_10433,N_10063);
xor U11519 (N_11519,N_10818,N_10516);
xnor U11520 (N_11520,N_10094,N_10727);
nand U11521 (N_11521,N_10564,N_10290);
and U11522 (N_11522,N_10431,N_10485);
and U11523 (N_11523,N_10150,N_10673);
nor U11524 (N_11524,N_10910,N_10903);
nor U11525 (N_11525,N_10911,N_10149);
and U11526 (N_11526,N_10120,N_10330);
or U11527 (N_11527,N_10344,N_10074);
nand U11528 (N_11528,N_10777,N_10129);
nor U11529 (N_11529,N_10539,N_10701);
or U11530 (N_11530,N_10983,N_10570);
or U11531 (N_11531,N_10628,N_10742);
nand U11532 (N_11532,N_10715,N_10683);
nand U11533 (N_11533,N_10164,N_10588);
xor U11534 (N_11534,N_10915,N_10272);
and U11535 (N_11535,N_10330,N_10421);
xor U11536 (N_11536,N_10062,N_10800);
or U11537 (N_11537,N_10875,N_10491);
and U11538 (N_11538,N_10911,N_10479);
xnor U11539 (N_11539,N_10267,N_10112);
nor U11540 (N_11540,N_10718,N_10837);
xnor U11541 (N_11541,N_10467,N_10369);
or U11542 (N_11542,N_10602,N_10042);
xor U11543 (N_11543,N_10064,N_10231);
and U11544 (N_11544,N_10459,N_10999);
and U11545 (N_11545,N_10520,N_10399);
nor U11546 (N_11546,N_10607,N_10367);
nand U11547 (N_11547,N_10430,N_10434);
and U11548 (N_11548,N_10254,N_10992);
or U11549 (N_11549,N_10418,N_10935);
nor U11550 (N_11550,N_10893,N_10131);
xnor U11551 (N_11551,N_10207,N_10325);
nor U11552 (N_11552,N_10668,N_10150);
or U11553 (N_11553,N_10680,N_10482);
xnor U11554 (N_11554,N_10723,N_10196);
xnor U11555 (N_11555,N_10482,N_10188);
nor U11556 (N_11556,N_10111,N_10778);
and U11557 (N_11557,N_10091,N_10745);
nor U11558 (N_11558,N_10890,N_10533);
and U11559 (N_11559,N_10309,N_10419);
xnor U11560 (N_11560,N_10444,N_10275);
nand U11561 (N_11561,N_10696,N_10459);
nor U11562 (N_11562,N_10102,N_10961);
or U11563 (N_11563,N_10175,N_10561);
and U11564 (N_11564,N_10734,N_10127);
or U11565 (N_11565,N_10610,N_10039);
xor U11566 (N_11566,N_10196,N_10063);
xor U11567 (N_11567,N_10623,N_10799);
or U11568 (N_11568,N_10955,N_10737);
or U11569 (N_11569,N_10393,N_10387);
xnor U11570 (N_11570,N_10773,N_10837);
and U11571 (N_11571,N_10223,N_10774);
nor U11572 (N_11572,N_10448,N_10339);
nor U11573 (N_11573,N_10977,N_10334);
and U11574 (N_11574,N_10348,N_10911);
and U11575 (N_11575,N_10986,N_10753);
nor U11576 (N_11576,N_10629,N_10439);
nand U11577 (N_11577,N_10390,N_10090);
xnor U11578 (N_11578,N_10819,N_10939);
and U11579 (N_11579,N_10713,N_10822);
or U11580 (N_11580,N_10664,N_10105);
and U11581 (N_11581,N_10186,N_10419);
or U11582 (N_11582,N_10699,N_10402);
nand U11583 (N_11583,N_10990,N_10252);
xnor U11584 (N_11584,N_10116,N_10795);
nor U11585 (N_11585,N_10249,N_10837);
xor U11586 (N_11586,N_10499,N_10955);
nand U11587 (N_11587,N_10966,N_10383);
and U11588 (N_11588,N_10037,N_10599);
or U11589 (N_11589,N_10590,N_10460);
xor U11590 (N_11590,N_10399,N_10243);
xor U11591 (N_11591,N_10839,N_10212);
nand U11592 (N_11592,N_10107,N_10977);
or U11593 (N_11593,N_10838,N_10278);
nand U11594 (N_11594,N_10513,N_10956);
nand U11595 (N_11595,N_10418,N_10171);
and U11596 (N_11596,N_10687,N_10377);
and U11597 (N_11597,N_10190,N_10767);
xor U11598 (N_11598,N_10200,N_10407);
xnor U11599 (N_11599,N_10632,N_10044);
nor U11600 (N_11600,N_10495,N_10998);
nand U11601 (N_11601,N_10486,N_10428);
xor U11602 (N_11602,N_10545,N_10146);
or U11603 (N_11603,N_10376,N_10027);
and U11604 (N_11604,N_10224,N_10312);
nand U11605 (N_11605,N_10975,N_10344);
nor U11606 (N_11606,N_10106,N_10037);
nand U11607 (N_11607,N_10903,N_10375);
nand U11608 (N_11608,N_10162,N_10489);
or U11609 (N_11609,N_10189,N_10555);
nor U11610 (N_11610,N_10838,N_10409);
nand U11611 (N_11611,N_10750,N_10117);
xor U11612 (N_11612,N_10155,N_10063);
or U11613 (N_11613,N_10278,N_10010);
nor U11614 (N_11614,N_10220,N_10673);
xor U11615 (N_11615,N_10251,N_10551);
or U11616 (N_11616,N_10376,N_10488);
nand U11617 (N_11617,N_10234,N_10258);
and U11618 (N_11618,N_10075,N_10204);
xor U11619 (N_11619,N_10479,N_10570);
nand U11620 (N_11620,N_10841,N_10591);
xnor U11621 (N_11621,N_10886,N_10431);
and U11622 (N_11622,N_10864,N_10069);
nand U11623 (N_11623,N_10772,N_10219);
or U11624 (N_11624,N_10684,N_10426);
nand U11625 (N_11625,N_10430,N_10996);
xor U11626 (N_11626,N_10420,N_10200);
nand U11627 (N_11627,N_10067,N_10879);
nand U11628 (N_11628,N_10602,N_10928);
nand U11629 (N_11629,N_10564,N_10386);
and U11630 (N_11630,N_10027,N_10471);
and U11631 (N_11631,N_10923,N_10029);
or U11632 (N_11632,N_10648,N_10700);
nor U11633 (N_11633,N_10122,N_10033);
xnor U11634 (N_11634,N_10097,N_10839);
nand U11635 (N_11635,N_10452,N_10507);
nand U11636 (N_11636,N_10206,N_10875);
nor U11637 (N_11637,N_10176,N_10916);
and U11638 (N_11638,N_10635,N_10317);
nand U11639 (N_11639,N_10819,N_10251);
or U11640 (N_11640,N_10442,N_10602);
nand U11641 (N_11641,N_10305,N_10389);
or U11642 (N_11642,N_10348,N_10307);
or U11643 (N_11643,N_10298,N_10439);
nand U11644 (N_11644,N_10849,N_10405);
nor U11645 (N_11645,N_10272,N_10205);
and U11646 (N_11646,N_10526,N_10967);
and U11647 (N_11647,N_10212,N_10972);
nor U11648 (N_11648,N_10591,N_10487);
xor U11649 (N_11649,N_10452,N_10867);
nor U11650 (N_11650,N_10008,N_10966);
and U11651 (N_11651,N_10973,N_10252);
or U11652 (N_11652,N_10821,N_10233);
nand U11653 (N_11653,N_10682,N_10797);
nor U11654 (N_11654,N_10751,N_10386);
nor U11655 (N_11655,N_10246,N_10419);
or U11656 (N_11656,N_10134,N_10069);
and U11657 (N_11657,N_10708,N_10121);
nor U11658 (N_11658,N_10193,N_10416);
xnor U11659 (N_11659,N_10306,N_10250);
or U11660 (N_11660,N_10810,N_10640);
xor U11661 (N_11661,N_10509,N_10378);
xnor U11662 (N_11662,N_10397,N_10944);
xor U11663 (N_11663,N_10523,N_10295);
nand U11664 (N_11664,N_10184,N_10842);
and U11665 (N_11665,N_10625,N_10332);
xor U11666 (N_11666,N_10452,N_10753);
nand U11667 (N_11667,N_10399,N_10278);
nor U11668 (N_11668,N_10138,N_10221);
nand U11669 (N_11669,N_10541,N_10483);
and U11670 (N_11670,N_10029,N_10136);
xnor U11671 (N_11671,N_10055,N_10323);
xnor U11672 (N_11672,N_10114,N_10746);
and U11673 (N_11673,N_10782,N_10945);
nor U11674 (N_11674,N_10013,N_10679);
or U11675 (N_11675,N_10080,N_10082);
xnor U11676 (N_11676,N_10069,N_10614);
or U11677 (N_11677,N_10631,N_10416);
and U11678 (N_11678,N_10000,N_10805);
and U11679 (N_11679,N_10775,N_10991);
or U11680 (N_11680,N_10967,N_10080);
or U11681 (N_11681,N_10088,N_10455);
nand U11682 (N_11682,N_10953,N_10178);
nor U11683 (N_11683,N_10844,N_10774);
or U11684 (N_11684,N_10570,N_10113);
nand U11685 (N_11685,N_10455,N_10509);
xnor U11686 (N_11686,N_10884,N_10428);
xnor U11687 (N_11687,N_10180,N_10718);
and U11688 (N_11688,N_10894,N_10965);
nor U11689 (N_11689,N_10541,N_10420);
xnor U11690 (N_11690,N_10287,N_10811);
and U11691 (N_11691,N_10634,N_10161);
or U11692 (N_11692,N_10398,N_10016);
or U11693 (N_11693,N_10475,N_10599);
or U11694 (N_11694,N_10983,N_10949);
nand U11695 (N_11695,N_10458,N_10099);
nand U11696 (N_11696,N_10410,N_10655);
nor U11697 (N_11697,N_10813,N_10807);
xor U11698 (N_11698,N_10081,N_10086);
and U11699 (N_11699,N_10379,N_10288);
and U11700 (N_11700,N_10556,N_10578);
xnor U11701 (N_11701,N_10590,N_10507);
nand U11702 (N_11702,N_10431,N_10333);
and U11703 (N_11703,N_10732,N_10099);
xor U11704 (N_11704,N_10826,N_10932);
and U11705 (N_11705,N_10251,N_10254);
or U11706 (N_11706,N_10577,N_10674);
nor U11707 (N_11707,N_10563,N_10652);
or U11708 (N_11708,N_10565,N_10785);
or U11709 (N_11709,N_10651,N_10710);
nand U11710 (N_11710,N_10519,N_10491);
nand U11711 (N_11711,N_10012,N_10468);
or U11712 (N_11712,N_10856,N_10353);
nor U11713 (N_11713,N_10222,N_10378);
xor U11714 (N_11714,N_10984,N_10597);
xor U11715 (N_11715,N_10286,N_10328);
or U11716 (N_11716,N_10201,N_10860);
nor U11717 (N_11717,N_10837,N_10218);
nor U11718 (N_11718,N_10074,N_10690);
nand U11719 (N_11719,N_10680,N_10839);
xor U11720 (N_11720,N_10446,N_10545);
xnor U11721 (N_11721,N_10125,N_10275);
nand U11722 (N_11722,N_10669,N_10969);
or U11723 (N_11723,N_10926,N_10444);
xor U11724 (N_11724,N_10156,N_10309);
nand U11725 (N_11725,N_10593,N_10907);
nor U11726 (N_11726,N_10534,N_10470);
nor U11727 (N_11727,N_10517,N_10092);
and U11728 (N_11728,N_10099,N_10018);
xnor U11729 (N_11729,N_10133,N_10655);
and U11730 (N_11730,N_10616,N_10064);
or U11731 (N_11731,N_10102,N_10699);
nand U11732 (N_11732,N_10729,N_10920);
and U11733 (N_11733,N_10080,N_10190);
or U11734 (N_11734,N_10984,N_10463);
nor U11735 (N_11735,N_10281,N_10184);
and U11736 (N_11736,N_10808,N_10350);
or U11737 (N_11737,N_10811,N_10540);
and U11738 (N_11738,N_10723,N_10934);
nor U11739 (N_11739,N_10606,N_10375);
xor U11740 (N_11740,N_10391,N_10117);
or U11741 (N_11741,N_10583,N_10289);
nand U11742 (N_11742,N_10994,N_10641);
or U11743 (N_11743,N_10900,N_10336);
xnor U11744 (N_11744,N_10251,N_10502);
or U11745 (N_11745,N_10800,N_10024);
xor U11746 (N_11746,N_10783,N_10286);
xnor U11747 (N_11747,N_10059,N_10807);
or U11748 (N_11748,N_10400,N_10910);
nand U11749 (N_11749,N_10956,N_10254);
nand U11750 (N_11750,N_10984,N_10938);
and U11751 (N_11751,N_10361,N_10859);
xor U11752 (N_11752,N_10936,N_10784);
nor U11753 (N_11753,N_10477,N_10239);
or U11754 (N_11754,N_10386,N_10291);
nand U11755 (N_11755,N_10566,N_10143);
nor U11756 (N_11756,N_10768,N_10249);
xnor U11757 (N_11757,N_10437,N_10634);
nand U11758 (N_11758,N_10798,N_10757);
xnor U11759 (N_11759,N_10653,N_10597);
or U11760 (N_11760,N_10915,N_10293);
and U11761 (N_11761,N_10084,N_10136);
nand U11762 (N_11762,N_10060,N_10666);
and U11763 (N_11763,N_10719,N_10003);
nand U11764 (N_11764,N_10792,N_10897);
xor U11765 (N_11765,N_10635,N_10355);
nor U11766 (N_11766,N_10932,N_10272);
or U11767 (N_11767,N_10351,N_10179);
nand U11768 (N_11768,N_10199,N_10438);
nand U11769 (N_11769,N_10505,N_10100);
and U11770 (N_11770,N_10978,N_10668);
or U11771 (N_11771,N_10748,N_10438);
nor U11772 (N_11772,N_10748,N_10701);
nand U11773 (N_11773,N_10395,N_10037);
nor U11774 (N_11774,N_10461,N_10744);
xnor U11775 (N_11775,N_10187,N_10981);
and U11776 (N_11776,N_10922,N_10479);
and U11777 (N_11777,N_10280,N_10715);
nand U11778 (N_11778,N_10515,N_10610);
and U11779 (N_11779,N_10073,N_10280);
or U11780 (N_11780,N_10343,N_10796);
or U11781 (N_11781,N_10735,N_10025);
nor U11782 (N_11782,N_10757,N_10167);
nor U11783 (N_11783,N_10813,N_10157);
or U11784 (N_11784,N_10800,N_10798);
and U11785 (N_11785,N_10716,N_10403);
and U11786 (N_11786,N_10939,N_10513);
xnor U11787 (N_11787,N_10942,N_10963);
or U11788 (N_11788,N_10226,N_10642);
nor U11789 (N_11789,N_10207,N_10037);
and U11790 (N_11790,N_10689,N_10473);
and U11791 (N_11791,N_10585,N_10124);
nor U11792 (N_11792,N_10428,N_10595);
and U11793 (N_11793,N_10511,N_10987);
and U11794 (N_11794,N_10925,N_10538);
nand U11795 (N_11795,N_10596,N_10244);
nor U11796 (N_11796,N_10190,N_10142);
nor U11797 (N_11797,N_10631,N_10223);
nor U11798 (N_11798,N_10601,N_10069);
nor U11799 (N_11799,N_10049,N_10942);
and U11800 (N_11800,N_10593,N_10978);
nor U11801 (N_11801,N_10153,N_10194);
nand U11802 (N_11802,N_10934,N_10904);
or U11803 (N_11803,N_10650,N_10080);
or U11804 (N_11804,N_10430,N_10358);
nand U11805 (N_11805,N_10814,N_10481);
and U11806 (N_11806,N_10814,N_10091);
and U11807 (N_11807,N_10084,N_10531);
nor U11808 (N_11808,N_10282,N_10005);
or U11809 (N_11809,N_10033,N_10370);
nand U11810 (N_11810,N_10859,N_10931);
or U11811 (N_11811,N_10233,N_10089);
or U11812 (N_11812,N_10234,N_10069);
nor U11813 (N_11813,N_10354,N_10911);
or U11814 (N_11814,N_10938,N_10344);
and U11815 (N_11815,N_10775,N_10245);
or U11816 (N_11816,N_10534,N_10582);
nor U11817 (N_11817,N_10284,N_10788);
xnor U11818 (N_11818,N_10165,N_10412);
and U11819 (N_11819,N_10745,N_10171);
nor U11820 (N_11820,N_10580,N_10029);
nand U11821 (N_11821,N_10465,N_10958);
or U11822 (N_11822,N_10869,N_10557);
nand U11823 (N_11823,N_10430,N_10887);
xor U11824 (N_11824,N_10469,N_10080);
or U11825 (N_11825,N_10512,N_10485);
nand U11826 (N_11826,N_10756,N_10728);
and U11827 (N_11827,N_10707,N_10697);
nor U11828 (N_11828,N_10492,N_10418);
xnor U11829 (N_11829,N_10931,N_10068);
xnor U11830 (N_11830,N_10109,N_10502);
or U11831 (N_11831,N_10666,N_10701);
nor U11832 (N_11832,N_10975,N_10560);
or U11833 (N_11833,N_10002,N_10684);
and U11834 (N_11834,N_10444,N_10144);
and U11835 (N_11835,N_10250,N_10193);
and U11836 (N_11836,N_10942,N_10895);
nand U11837 (N_11837,N_10547,N_10181);
xnor U11838 (N_11838,N_10244,N_10153);
and U11839 (N_11839,N_10892,N_10153);
nand U11840 (N_11840,N_10197,N_10116);
and U11841 (N_11841,N_10410,N_10687);
or U11842 (N_11842,N_10668,N_10567);
nand U11843 (N_11843,N_10802,N_10760);
nor U11844 (N_11844,N_10951,N_10277);
and U11845 (N_11845,N_10313,N_10450);
or U11846 (N_11846,N_10142,N_10981);
and U11847 (N_11847,N_10236,N_10185);
and U11848 (N_11848,N_10009,N_10447);
nor U11849 (N_11849,N_10210,N_10357);
xnor U11850 (N_11850,N_10887,N_10474);
and U11851 (N_11851,N_10361,N_10130);
and U11852 (N_11852,N_10571,N_10826);
and U11853 (N_11853,N_10799,N_10153);
xnor U11854 (N_11854,N_10957,N_10768);
nand U11855 (N_11855,N_10979,N_10320);
or U11856 (N_11856,N_10268,N_10870);
nor U11857 (N_11857,N_10071,N_10288);
or U11858 (N_11858,N_10531,N_10991);
xnor U11859 (N_11859,N_10337,N_10573);
nor U11860 (N_11860,N_10587,N_10435);
xor U11861 (N_11861,N_10289,N_10437);
xnor U11862 (N_11862,N_10501,N_10787);
xor U11863 (N_11863,N_10960,N_10875);
nand U11864 (N_11864,N_10232,N_10419);
xor U11865 (N_11865,N_10120,N_10733);
nand U11866 (N_11866,N_10243,N_10724);
nor U11867 (N_11867,N_10191,N_10501);
nor U11868 (N_11868,N_10431,N_10609);
nor U11869 (N_11869,N_10263,N_10839);
nand U11870 (N_11870,N_10160,N_10261);
nand U11871 (N_11871,N_10557,N_10066);
and U11872 (N_11872,N_10329,N_10166);
nand U11873 (N_11873,N_10655,N_10248);
xor U11874 (N_11874,N_10538,N_10988);
xnor U11875 (N_11875,N_10136,N_10863);
nand U11876 (N_11876,N_10566,N_10038);
and U11877 (N_11877,N_10152,N_10717);
nor U11878 (N_11878,N_10910,N_10222);
xor U11879 (N_11879,N_10132,N_10434);
or U11880 (N_11880,N_10462,N_10311);
nand U11881 (N_11881,N_10675,N_10419);
and U11882 (N_11882,N_10411,N_10960);
nand U11883 (N_11883,N_10312,N_10432);
nor U11884 (N_11884,N_10056,N_10820);
nor U11885 (N_11885,N_10814,N_10703);
nand U11886 (N_11886,N_10709,N_10346);
nor U11887 (N_11887,N_10605,N_10054);
or U11888 (N_11888,N_10261,N_10243);
nand U11889 (N_11889,N_10247,N_10911);
xnor U11890 (N_11890,N_10513,N_10999);
nor U11891 (N_11891,N_10310,N_10741);
nor U11892 (N_11892,N_10836,N_10208);
or U11893 (N_11893,N_10225,N_10114);
and U11894 (N_11894,N_10454,N_10672);
xor U11895 (N_11895,N_10424,N_10685);
xor U11896 (N_11896,N_10399,N_10215);
and U11897 (N_11897,N_10141,N_10538);
nor U11898 (N_11898,N_10771,N_10582);
nand U11899 (N_11899,N_10403,N_10313);
and U11900 (N_11900,N_10584,N_10258);
nand U11901 (N_11901,N_10188,N_10360);
xor U11902 (N_11902,N_10039,N_10964);
and U11903 (N_11903,N_10918,N_10454);
and U11904 (N_11904,N_10063,N_10358);
and U11905 (N_11905,N_10545,N_10021);
nand U11906 (N_11906,N_10847,N_10727);
nand U11907 (N_11907,N_10669,N_10966);
xnor U11908 (N_11908,N_10553,N_10666);
and U11909 (N_11909,N_10738,N_10330);
nor U11910 (N_11910,N_10061,N_10457);
xor U11911 (N_11911,N_10028,N_10471);
and U11912 (N_11912,N_10881,N_10932);
or U11913 (N_11913,N_10874,N_10757);
nand U11914 (N_11914,N_10447,N_10495);
or U11915 (N_11915,N_10407,N_10399);
nand U11916 (N_11916,N_10460,N_10938);
nor U11917 (N_11917,N_10509,N_10099);
nor U11918 (N_11918,N_10515,N_10862);
nand U11919 (N_11919,N_10071,N_10770);
and U11920 (N_11920,N_10941,N_10587);
or U11921 (N_11921,N_10459,N_10492);
nor U11922 (N_11922,N_10202,N_10509);
or U11923 (N_11923,N_10296,N_10752);
or U11924 (N_11924,N_10660,N_10731);
nand U11925 (N_11925,N_10668,N_10941);
xor U11926 (N_11926,N_10597,N_10723);
and U11927 (N_11927,N_10246,N_10250);
or U11928 (N_11928,N_10057,N_10379);
nor U11929 (N_11929,N_10262,N_10581);
or U11930 (N_11930,N_10036,N_10675);
nand U11931 (N_11931,N_10891,N_10660);
nor U11932 (N_11932,N_10420,N_10897);
nand U11933 (N_11933,N_10625,N_10866);
and U11934 (N_11934,N_10302,N_10393);
nor U11935 (N_11935,N_10864,N_10990);
or U11936 (N_11936,N_10317,N_10799);
nand U11937 (N_11937,N_10814,N_10691);
nand U11938 (N_11938,N_10070,N_10487);
or U11939 (N_11939,N_10774,N_10291);
xnor U11940 (N_11940,N_10362,N_10036);
xnor U11941 (N_11941,N_10780,N_10203);
nor U11942 (N_11942,N_10225,N_10004);
nor U11943 (N_11943,N_10195,N_10874);
nand U11944 (N_11944,N_10896,N_10146);
nand U11945 (N_11945,N_10347,N_10895);
xnor U11946 (N_11946,N_10969,N_10502);
or U11947 (N_11947,N_10110,N_10027);
nor U11948 (N_11948,N_10413,N_10172);
or U11949 (N_11949,N_10152,N_10974);
nor U11950 (N_11950,N_10360,N_10915);
or U11951 (N_11951,N_10194,N_10588);
xnor U11952 (N_11952,N_10820,N_10853);
or U11953 (N_11953,N_10221,N_10429);
xnor U11954 (N_11954,N_10811,N_10606);
or U11955 (N_11955,N_10777,N_10729);
and U11956 (N_11956,N_10712,N_10108);
and U11957 (N_11957,N_10095,N_10596);
and U11958 (N_11958,N_10614,N_10597);
or U11959 (N_11959,N_10674,N_10488);
nand U11960 (N_11960,N_10635,N_10013);
and U11961 (N_11961,N_10277,N_10338);
or U11962 (N_11962,N_10700,N_10683);
nand U11963 (N_11963,N_10894,N_10078);
or U11964 (N_11964,N_10051,N_10452);
or U11965 (N_11965,N_10674,N_10043);
and U11966 (N_11966,N_10678,N_10320);
xnor U11967 (N_11967,N_10393,N_10045);
nand U11968 (N_11968,N_10870,N_10159);
nor U11969 (N_11969,N_10757,N_10563);
and U11970 (N_11970,N_10236,N_10723);
or U11971 (N_11971,N_10654,N_10574);
nor U11972 (N_11972,N_10294,N_10250);
xnor U11973 (N_11973,N_10000,N_10529);
and U11974 (N_11974,N_10711,N_10560);
xnor U11975 (N_11975,N_10468,N_10545);
or U11976 (N_11976,N_10981,N_10217);
and U11977 (N_11977,N_10316,N_10894);
nand U11978 (N_11978,N_10906,N_10284);
or U11979 (N_11979,N_10871,N_10905);
or U11980 (N_11980,N_10697,N_10227);
or U11981 (N_11981,N_10859,N_10772);
nand U11982 (N_11982,N_10000,N_10621);
nor U11983 (N_11983,N_10787,N_10746);
and U11984 (N_11984,N_10793,N_10896);
nand U11985 (N_11985,N_10046,N_10767);
and U11986 (N_11986,N_10034,N_10835);
and U11987 (N_11987,N_10193,N_10402);
and U11988 (N_11988,N_10408,N_10521);
or U11989 (N_11989,N_10507,N_10878);
nor U11990 (N_11990,N_10043,N_10184);
nand U11991 (N_11991,N_10661,N_10875);
and U11992 (N_11992,N_10056,N_10470);
xor U11993 (N_11993,N_10424,N_10144);
and U11994 (N_11994,N_10403,N_10782);
nand U11995 (N_11995,N_10788,N_10576);
nand U11996 (N_11996,N_10233,N_10564);
and U11997 (N_11997,N_10992,N_10897);
xor U11998 (N_11998,N_10648,N_10932);
and U11999 (N_11999,N_10597,N_10804);
and U12000 (N_12000,N_11029,N_11967);
nor U12001 (N_12001,N_11020,N_11389);
or U12002 (N_12002,N_11616,N_11207);
or U12003 (N_12003,N_11147,N_11933);
nand U12004 (N_12004,N_11945,N_11709);
or U12005 (N_12005,N_11805,N_11747);
nor U12006 (N_12006,N_11537,N_11507);
nand U12007 (N_12007,N_11232,N_11190);
or U12008 (N_12008,N_11339,N_11305);
and U12009 (N_12009,N_11285,N_11535);
nor U12010 (N_12010,N_11669,N_11549);
nor U12011 (N_12011,N_11929,N_11873);
nor U12012 (N_12012,N_11003,N_11472);
nand U12013 (N_12013,N_11772,N_11824);
nand U12014 (N_12014,N_11785,N_11219);
xor U12015 (N_12015,N_11303,N_11144);
or U12016 (N_12016,N_11782,N_11658);
nand U12017 (N_12017,N_11295,N_11229);
or U12018 (N_12018,N_11088,N_11018);
xnor U12019 (N_12019,N_11813,N_11275);
or U12020 (N_12020,N_11071,N_11524);
or U12021 (N_12021,N_11917,N_11919);
and U12022 (N_12022,N_11613,N_11134);
or U12023 (N_12023,N_11469,N_11889);
or U12024 (N_12024,N_11490,N_11256);
xor U12025 (N_12025,N_11653,N_11848);
nor U12026 (N_12026,N_11804,N_11587);
nor U12027 (N_12027,N_11569,N_11575);
nand U12028 (N_12028,N_11337,N_11854);
nor U12029 (N_12029,N_11129,N_11744);
nand U12030 (N_12030,N_11547,N_11151);
and U12031 (N_12031,N_11157,N_11483);
nor U12032 (N_12032,N_11221,N_11960);
nand U12033 (N_12033,N_11066,N_11054);
nor U12034 (N_12034,N_11489,N_11815);
xnor U12035 (N_12035,N_11384,N_11769);
xor U12036 (N_12036,N_11936,N_11609);
or U12037 (N_12037,N_11555,N_11974);
or U12038 (N_12038,N_11953,N_11801);
or U12039 (N_12039,N_11468,N_11876);
nand U12040 (N_12040,N_11736,N_11301);
xnor U12041 (N_12041,N_11759,N_11154);
or U12042 (N_12042,N_11955,N_11198);
and U12043 (N_12043,N_11450,N_11139);
or U12044 (N_12044,N_11189,N_11006);
nand U12045 (N_12045,N_11973,N_11979);
or U12046 (N_12046,N_11556,N_11745);
nor U12047 (N_12047,N_11534,N_11619);
xor U12048 (N_12048,N_11734,N_11114);
xor U12049 (N_12049,N_11090,N_11526);
nand U12050 (N_12050,N_11203,N_11227);
nand U12051 (N_12051,N_11880,N_11529);
and U12052 (N_12052,N_11493,N_11320);
nand U12053 (N_12053,N_11372,N_11254);
or U12054 (N_12054,N_11317,N_11686);
nand U12055 (N_12055,N_11228,N_11521);
xor U12056 (N_12056,N_11716,N_11268);
xnor U12057 (N_12057,N_11459,N_11480);
xor U12058 (N_12058,N_11969,N_11554);
nor U12059 (N_12059,N_11695,N_11205);
nand U12060 (N_12060,N_11059,N_11302);
nand U12061 (N_12061,N_11046,N_11342);
xor U12062 (N_12062,N_11853,N_11774);
nand U12063 (N_12063,N_11290,N_11764);
xor U12064 (N_12064,N_11859,N_11894);
and U12065 (N_12065,N_11588,N_11570);
xor U12066 (N_12066,N_11288,N_11340);
nand U12067 (N_12067,N_11623,N_11777);
and U12068 (N_12068,N_11610,N_11742);
nor U12069 (N_12069,N_11437,N_11428);
nor U12070 (N_12070,N_11064,N_11358);
nor U12071 (N_12071,N_11829,N_11943);
nor U12072 (N_12072,N_11224,N_11075);
nand U12073 (N_12073,N_11362,N_11706);
or U12074 (N_12074,N_11366,N_11976);
and U12075 (N_12075,N_11142,N_11211);
or U12076 (N_12076,N_11625,N_11084);
xor U12077 (N_12077,N_11400,N_11098);
and U12078 (N_12078,N_11385,N_11741);
xnor U12079 (N_12079,N_11944,N_11025);
nor U12080 (N_12080,N_11286,N_11171);
nor U12081 (N_12081,N_11710,N_11421);
xnor U12082 (N_12082,N_11835,N_11940);
nand U12083 (N_12083,N_11107,N_11466);
nor U12084 (N_12084,N_11430,N_11872);
nor U12085 (N_12085,N_11886,N_11331);
nor U12086 (N_12086,N_11831,N_11603);
or U12087 (N_12087,N_11380,N_11453);
nor U12088 (N_12088,N_11418,N_11394);
nand U12089 (N_12089,N_11530,N_11773);
or U12090 (N_12090,N_11344,N_11345);
and U12091 (N_12091,N_11776,N_11986);
or U12092 (N_12092,N_11907,N_11921);
xor U12093 (N_12093,N_11849,N_11137);
nand U12094 (N_12094,N_11012,N_11665);
and U12095 (N_12095,N_11553,N_11467);
nor U12096 (N_12096,N_11998,N_11648);
and U12097 (N_12097,N_11370,N_11070);
and U12098 (N_12098,N_11594,N_11024);
xor U12099 (N_12099,N_11324,N_11712);
xor U12100 (N_12100,N_11009,N_11840);
xnor U12101 (N_12101,N_11100,N_11057);
nand U12102 (N_12102,N_11338,N_11375);
nor U12103 (N_12103,N_11404,N_11896);
and U12104 (N_12104,N_11749,N_11335);
and U12105 (N_12105,N_11265,N_11138);
nand U12106 (N_12106,N_11667,N_11373);
or U12107 (N_12107,N_11272,N_11714);
xor U12108 (N_12108,N_11146,N_11803);
nor U12109 (N_12109,N_11433,N_11935);
nand U12110 (N_12110,N_11761,N_11562);
xnor U12111 (N_12111,N_11270,N_11898);
and U12112 (N_12112,N_11497,N_11760);
nand U12113 (N_12113,N_11304,N_11184);
nand U12114 (N_12114,N_11197,N_11503);
xnor U12115 (N_12115,N_11635,N_11685);
xnor U12116 (N_12116,N_11456,N_11532);
nor U12117 (N_12117,N_11826,N_11014);
xnor U12118 (N_12118,N_11789,N_11308);
or U12119 (N_12119,N_11023,N_11730);
xor U12120 (N_12120,N_11850,N_11168);
nand U12121 (N_12121,N_11405,N_11802);
or U12122 (N_12122,N_11444,N_11699);
nor U12123 (N_12123,N_11432,N_11688);
nor U12124 (N_12124,N_11266,N_11527);
xnor U12125 (N_12125,N_11871,N_11614);
nor U12126 (N_12126,N_11663,N_11934);
xnor U12127 (N_12127,N_11128,N_11291);
nand U12128 (N_12128,N_11214,N_11520);
and U12129 (N_12129,N_11120,N_11952);
and U12130 (N_12130,N_11043,N_11852);
and U12131 (N_12131,N_11412,N_11992);
or U12132 (N_12132,N_11330,N_11806);
nor U12133 (N_12133,N_11512,N_11116);
or U12134 (N_12134,N_11584,N_11204);
or U12135 (N_12135,N_11127,N_11581);
or U12136 (N_12136,N_11795,N_11494);
and U12137 (N_12137,N_11596,N_11487);
nor U12138 (N_12138,N_11514,N_11536);
xnor U12139 (N_12139,N_11949,N_11951);
nor U12140 (N_12140,N_11689,N_11156);
nand U12141 (N_12141,N_11259,N_11775);
nand U12142 (N_12142,N_11991,N_11533);
and U12143 (N_12143,N_11877,N_11732);
or U12144 (N_12144,N_11167,N_11179);
nand U12145 (N_12145,N_11542,N_11048);
nor U12146 (N_12146,N_11263,N_11704);
xnor U12147 (N_12147,N_11861,N_11959);
and U12148 (N_12148,N_11176,N_11900);
nand U12149 (N_12149,N_11130,N_11844);
nor U12150 (N_12150,N_11578,N_11217);
nand U12151 (N_12151,N_11771,N_11436);
nand U12152 (N_12152,N_11995,N_11102);
xnor U12153 (N_12153,N_11895,N_11376);
nor U12154 (N_12154,N_11531,N_11506);
nor U12155 (N_12155,N_11654,N_11858);
or U12156 (N_12156,N_11621,N_11620);
nor U12157 (N_12157,N_11975,N_11173);
xnor U12158 (N_12158,N_11281,N_11209);
nand U12159 (N_12159,N_11212,N_11862);
nor U12160 (N_12160,N_11242,N_11629);
nor U12161 (N_12161,N_11273,N_11087);
xor U12162 (N_12162,N_11500,N_11423);
or U12163 (N_12163,N_11318,N_11668);
xor U12164 (N_12164,N_11316,N_11722);
xor U12165 (N_12165,N_11363,N_11425);
nand U12166 (N_12166,N_11392,N_11968);
nand U12167 (N_12167,N_11278,N_11875);
or U12168 (N_12168,N_11296,N_11053);
or U12169 (N_12169,N_11312,N_11577);
nand U12170 (N_12170,N_11997,N_11637);
and U12171 (N_12171,N_11563,N_11152);
and U12172 (N_12172,N_11652,N_11402);
and U12173 (N_12173,N_11582,N_11007);
or U12174 (N_12174,N_11019,N_11583);
nor U12175 (N_12175,N_11640,N_11626);
or U12176 (N_12176,N_11041,N_11322);
nand U12177 (N_12177,N_11225,N_11115);
and U12178 (N_12178,N_11674,N_11797);
or U12179 (N_12179,N_11780,N_11237);
and U12180 (N_12180,N_11504,N_11365);
and U12181 (N_12181,N_11104,N_11409);
or U12182 (N_12182,N_11397,N_11264);
or U12183 (N_12183,N_11791,N_11993);
xor U12184 (N_12184,N_11326,N_11143);
xnor U12185 (N_12185,N_11381,N_11659);
xnor U12186 (N_12186,N_11280,N_11427);
nor U12187 (N_12187,N_11810,N_11618);
nor U12188 (N_12188,N_11989,N_11117);
nor U12189 (N_12189,N_11725,N_11250);
xor U12190 (N_12190,N_11111,N_11857);
nor U12191 (N_12191,N_11586,N_11557);
or U12192 (N_12192,N_11687,N_11611);
and U12193 (N_12193,N_11293,N_11125);
nor U12194 (N_12194,N_11624,N_11825);
xor U12195 (N_12195,N_11607,N_11794);
or U12196 (N_12196,N_11313,N_11118);
xor U12197 (N_12197,N_11416,N_11085);
and U12198 (N_12198,N_11486,N_11545);
xnor U12199 (N_12199,N_11391,N_11966);
and U12200 (N_12200,N_11961,N_11484);
nand U12201 (N_12201,N_11170,N_11932);
nor U12202 (N_12202,N_11140,N_11133);
xor U12203 (N_12203,N_11319,N_11601);
nand U12204 (N_12204,N_11440,N_11605);
and U12205 (N_12205,N_11905,N_11306);
nand U12206 (N_12206,N_11297,N_11792);
nor U12207 (N_12207,N_11081,N_11693);
nor U12208 (N_12208,N_11508,N_11767);
and U12209 (N_12209,N_11892,N_11244);
nand U12210 (N_12210,N_11914,N_11004);
and U12211 (N_12211,N_11163,N_11332);
nand U12212 (N_12212,N_11101,N_11200);
nor U12213 (N_12213,N_11817,N_11371);
xor U12214 (N_12214,N_11956,N_11031);
xnor U12215 (N_12215,N_11551,N_11255);
or U12216 (N_12216,N_11713,N_11707);
or U12217 (N_12217,N_11216,N_11705);
or U12218 (N_12218,N_11369,N_11869);
xor U12219 (N_12219,N_11191,N_11856);
nand U12220 (N_12220,N_11566,N_11307);
nand U12221 (N_12221,N_11454,N_11277);
nor U12222 (N_12222,N_11833,N_11336);
xor U12223 (N_12223,N_11253,N_11028);
or U12224 (N_12224,N_11887,N_11701);
or U12225 (N_12225,N_11061,N_11597);
nand U12226 (N_12226,N_11820,N_11121);
or U12227 (N_12227,N_11062,N_11522);
or U12228 (N_12228,N_11226,N_11631);
nand U12229 (N_12229,N_11576,N_11235);
nand U12230 (N_12230,N_11422,N_11465);
and U12231 (N_12231,N_11915,N_11234);
nor U12232 (N_12232,N_11863,N_11612);
nand U12233 (N_12233,N_11954,N_11119);
and U12234 (N_12234,N_11351,N_11841);
xor U12235 (N_12235,N_11496,N_11924);
nand U12236 (N_12236,N_11408,N_11113);
and U12237 (N_12237,N_11060,N_11681);
xnor U12238 (N_12238,N_11739,N_11148);
and U12239 (N_12239,N_11906,N_11548);
and U12240 (N_12240,N_11978,N_11883);
xnor U12241 (N_12241,N_11590,N_11922);
xor U12242 (N_12242,N_11194,N_11638);
or U12243 (N_12243,N_11516,N_11498);
nor U12244 (N_12244,N_11515,N_11196);
or U12245 (N_12245,N_11401,N_11393);
and U12246 (N_12246,N_11579,N_11642);
nor U12247 (N_12247,N_11013,N_11671);
nor U12248 (N_12248,N_11926,N_11823);
nor U12249 (N_12249,N_11415,N_11902);
or U12250 (N_12250,N_11463,N_11132);
nor U12251 (N_12251,N_11752,N_11036);
and U12252 (N_12252,N_11539,N_11723);
or U12253 (N_12253,N_11149,N_11161);
xor U12254 (N_12254,N_11809,N_11289);
xor U12255 (N_12255,N_11067,N_11650);
or U12256 (N_12256,N_11604,N_11505);
or U12257 (N_12257,N_11719,N_11799);
xor U12258 (N_12258,N_11044,N_11122);
nand U12259 (N_12259,N_11846,N_11199);
nor U12260 (N_12260,N_11692,N_11758);
or U12261 (N_12261,N_11965,N_11763);
and U12262 (N_12262,N_11231,N_11364);
and U12263 (N_12263,N_11449,N_11488);
nor U12264 (N_12264,N_11447,N_11571);
or U12265 (N_12265,N_11808,N_11315);
nor U12266 (N_12266,N_11697,N_11768);
nor U12267 (N_12267,N_11647,N_11881);
nor U12268 (N_12268,N_11930,N_11016);
nor U12269 (N_12269,N_11439,N_11192);
xor U12270 (N_12270,N_11543,N_11201);
xnor U12271 (N_12271,N_11348,N_11183);
or U12272 (N_12272,N_11368,N_11145);
and U12273 (N_12273,N_11055,N_11451);
xor U12274 (N_12274,N_11347,N_11977);
nand U12275 (N_12275,N_11655,N_11783);
or U12276 (N_12276,N_11038,N_11793);
xor U12277 (N_12277,N_11314,N_11050);
and U12278 (N_12278,N_11916,N_11680);
nor U12279 (N_12279,N_11948,N_11181);
xnor U12280 (N_12280,N_11248,N_11165);
nand U12281 (N_12281,N_11124,N_11673);
and U12282 (N_12282,N_11838,N_11839);
nand U12283 (N_12283,N_11374,N_11193);
and U12284 (N_12284,N_11925,N_11550);
and U12285 (N_12285,N_11106,N_11011);
xnor U12286 (N_12286,N_11093,N_11058);
or U12287 (N_12287,N_11517,N_11899);
nand U12288 (N_12288,N_11185,N_11386);
or U12289 (N_12289,N_11262,N_11528);
or U12290 (N_12290,N_11008,N_11051);
and U12291 (N_12291,N_11643,N_11646);
xor U12292 (N_12292,N_11420,N_11999);
nand U12293 (N_12293,N_11068,N_11559);
nand U12294 (N_12294,N_11931,N_11822);
nor U12295 (N_12295,N_11269,N_11112);
xor U12296 (N_12296,N_11166,N_11299);
nand U12297 (N_12297,N_11240,N_11395);
xor U12298 (N_12298,N_11510,N_11661);
or U12299 (N_12299,N_11241,N_11354);
and U12300 (N_12300,N_11000,N_11828);
xnor U12301 (N_12301,N_11202,N_11032);
and U12302 (N_12302,N_11341,N_11721);
nor U12303 (N_12303,N_11970,N_11383);
nand U12304 (N_12304,N_11069,N_11325);
nand U12305 (N_12305,N_11407,N_11920);
nand U12306 (N_12306,N_11230,N_11766);
nor U12307 (N_12307,N_11755,N_11399);
and U12308 (N_12308,N_11359,N_11186);
or U12309 (N_12309,N_11479,N_11309);
and U12310 (N_12310,N_11885,N_11893);
and U12311 (N_12311,N_11888,N_11355);
or U12312 (N_12312,N_11110,N_11047);
nand U12313 (N_12313,N_11947,N_11855);
and U12314 (N_12314,N_11746,N_11246);
and U12315 (N_12315,N_11083,N_11818);
nor U12316 (N_12316,N_11633,N_11287);
nand U12317 (N_12317,N_11985,N_11350);
nor U12318 (N_12318,N_11022,N_11649);
nor U12319 (N_12319,N_11834,N_11349);
nor U12320 (N_12320,N_11981,N_11426);
and U12321 (N_12321,N_11261,N_11215);
nor U12322 (N_12322,N_11518,N_11513);
or U12323 (N_12323,N_11731,N_11600);
nand U12324 (N_12324,N_11410,N_11743);
nand U12325 (N_12325,N_11434,N_11435);
nand U12326 (N_12326,N_11238,N_11664);
xnor U12327 (N_12327,N_11957,N_11442);
xor U12328 (N_12328,N_11323,N_11034);
and U12329 (N_12329,N_11837,N_11076);
nor U12330 (N_12330,N_11608,N_11720);
nand U12331 (N_12331,N_11080,N_11045);
or U12332 (N_12332,N_11591,N_11819);
nand U12333 (N_12333,N_11310,N_11352);
nor U12334 (N_12334,N_11572,N_11236);
and U12335 (N_12335,N_11891,N_11568);
and U12336 (N_12336,N_11471,N_11461);
nor U12337 (N_12337,N_11836,N_11702);
nor U12338 (N_12338,N_11162,N_11311);
xor U12339 (N_12339,N_11346,N_11475);
and U12340 (N_12340,N_11218,N_11321);
or U12341 (N_12341,N_11800,N_11411);
nand U12342 (N_12342,N_11065,N_11703);
xnor U12343 (N_12343,N_11049,N_11589);
or U12344 (N_12344,N_11552,N_11645);
xnor U12345 (N_12345,N_11786,N_11005);
xor U12346 (N_12346,N_11843,N_11738);
nor U12347 (N_12347,N_11431,N_11367);
nand U12348 (N_12348,N_11727,N_11188);
nand U12349 (N_12349,N_11252,N_11599);
nand U12350 (N_12350,N_11779,N_11708);
nor U12351 (N_12351,N_11091,N_11001);
nand U12352 (N_12352,N_11878,N_11762);
and U12353 (N_12353,N_11963,N_11403);
nor U12354 (N_12354,N_11908,N_11464);
nor U12355 (N_12355,N_11988,N_11082);
and U12356 (N_12356,N_11329,N_11561);
nor U12357 (N_12357,N_11950,N_11150);
nand U12358 (N_12358,N_11042,N_11481);
nand U12359 (N_12359,N_11448,N_11501);
or U12360 (N_12360,N_11615,N_11781);
nand U12361 (N_12361,N_11294,N_11135);
nor U12362 (N_12362,N_11711,N_11361);
nor U12363 (N_12363,N_11283,N_11443);
nand U12364 (N_12364,N_11832,N_11353);
or U12365 (N_12365,N_11728,N_11864);
nor U12366 (N_12366,N_11164,N_11327);
and U12367 (N_12367,N_11414,N_11360);
nand U12368 (N_12368,N_11847,N_11056);
xnor U12369 (N_12369,N_11700,N_11627);
and U12370 (N_12370,N_11413,N_11630);
nor U12371 (N_12371,N_11089,N_11239);
xnor U12372 (N_12372,N_11983,N_11724);
nand U12373 (N_12373,N_11910,N_11010);
xor U12374 (N_12374,N_11077,N_11994);
and U12375 (N_12375,N_11757,N_11021);
and U12376 (N_12376,N_11971,N_11628);
or U12377 (N_12377,N_11593,N_11622);
nand U12378 (N_12378,N_11798,N_11222);
nor U12379 (N_12379,N_11644,N_11560);
nor U12380 (N_12380,N_11251,N_11195);
nand U12381 (N_12381,N_11097,N_11258);
or U12382 (N_12382,N_11666,N_11718);
nor U12383 (N_12383,N_11595,N_11938);
or U12384 (N_12384,N_11754,N_11670);
nor U12385 (N_12385,N_11715,N_11580);
nand U12386 (N_12386,N_11866,N_11063);
nor U12387 (N_12387,N_11333,N_11473);
and U12388 (N_12388,N_11398,N_11874);
nand U12389 (N_12389,N_11598,N_11656);
xor U12390 (N_12390,N_11662,N_11182);
or U12391 (N_12391,N_11676,N_11641);
nand U12392 (N_12392,N_11492,N_11477);
xnor U12393 (N_12393,N_11074,N_11964);
nand U12394 (N_12394,N_11174,N_11564);
or U12395 (N_12395,N_11027,N_11429);
and U12396 (N_12396,N_11245,N_11814);
nand U12397 (N_12397,N_11417,N_11868);
nor U12398 (N_12398,N_11220,N_11495);
xor U12399 (N_12399,N_11851,N_11460);
nand U12400 (N_12400,N_11737,N_11017);
and U12401 (N_12401,N_11927,N_11602);
xnor U12402 (N_12402,N_11865,N_11079);
xnor U12403 (N_12403,N_11980,N_11770);
and U12404 (N_12404,N_11002,N_11158);
or U12405 (N_12405,N_11357,N_11382);
xnor U12406 (N_12406,N_11733,N_11458);
nand U12407 (N_12407,N_11675,N_11476);
xor U12408 (N_12408,N_11678,N_11690);
and U12409 (N_12409,N_11485,N_11750);
xnor U12410 (N_12410,N_11030,N_11208);
xnor U12411 (N_12411,N_11606,N_11086);
and U12412 (N_12412,N_11884,N_11984);
and U12413 (N_12413,N_11131,N_11276);
nor U12414 (N_12414,N_11573,N_11632);
nand U12415 (N_12415,N_11073,N_11691);
or U12416 (N_12416,N_11558,N_11334);
nand U12417 (N_12417,N_11567,N_11870);
xnor U12418 (N_12418,N_11223,N_11099);
nand U12419 (N_12419,N_11592,N_11901);
or U12420 (N_12420,N_11249,N_11816);
nor U12421 (N_12421,N_11206,N_11356);
and U12422 (N_12422,N_11788,N_11811);
nand U12423 (N_12423,N_11390,N_11812);
or U12424 (N_12424,N_11740,N_11136);
xor U12425 (N_12425,N_11677,N_11271);
or U12426 (N_12426,N_11617,N_11441);
nand U12427 (N_12427,N_11912,N_11040);
nor U12428 (N_12428,N_11928,N_11509);
xor U12429 (N_12429,N_11636,N_11913);
xnor U12430 (N_12430,N_11109,N_11039);
or U12431 (N_12431,N_11585,N_11284);
nand U12432 (N_12432,N_11694,N_11213);
and U12433 (N_12433,N_11343,N_11525);
xor U12434 (N_12434,N_11790,N_11491);
nand U12435 (N_12435,N_11379,N_11247);
and U12436 (N_12436,N_11177,N_11378);
and U12437 (N_12437,N_11243,N_11660);
or U12438 (N_12438,N_11438,N_11502);
nand U12439 (N_12439,N_11546,N_11153);
or U12440 (N_12440,N_11867,N_11698);
nor U12441 (N_12441,N_11972,N_11565);
or U12442 (N_12442,N_11574,N_11544);
xor U12443 (N_12443,N_11210,N_11541);
nand U12444 (N_12444,N_11377,N_11778);
or U12445 (N_12445,N_11679,N_11274);
and U12446 (N_12446,N_11126,N_11519);
or U12447 (N_12447,N_11026,N_11172);
xnor U12448 (N_12448,N_11753,N_11462);
nand U12449 (N_12449,N_11396,N_11078);
xor U12450 (N_12450,N_11178,N_11996);
or U12451 (N_12451,N_11105,N_11897);
or U12452 (N_12452,N_11424,N_11096);
or U12453 (N_12453,N_11180,N_11796);
or U12454 (N_12454,N_11942,N_11388);
or U12455 (N_12455,N_11939,N_11765);
or U12456 (N_12456,N_11918,N_11540);
nor U12457 (N_12457,N_11455,N_11470);
nor U12458 (N_12458,N_11072,N_11482);
or U12459 (N_12459,N_11159,N_11735);
xnor U12460 (N_12460,N_11923,N_11946);
nor U12461 (N_12461,N_11538,N_11639);
xor U12462 (N_12462,N_11890,N_11103);
nor U12463 (N_12463,N_11987,N_11830);
xnor U12464 (N_12464,N_11478,N_11882);
and U12465 (N_12465,N_11095,N_11842);
xor U12466 (N_12466,N_11155,N_11729);
xor U12467 (N_12467,N_11684,N_11267);
or U12468 (N_12468,N_11634,N_11328);
nor U12469 (N_12469,N_11958,N_11682);
and U12470 (N_12470,N_11233,N_11052);
xor U12471 (N_12471,N_11092,N_11683);
nand U12472 (N_12472,N_11672,N_11827);
nor U12473 (N_12473,N_11187,N_11903);
and U12474 (N_12474,N_11445,N_11787);
nand U12475 (N_12475,N_11756,N_11457);
nand U12476 (N_12476,N_11990,N_11015);
nand U12477 (N_12477,N_11845,N_11523);
or U12478 (N_12478,N_11726,N_11651);
or U12479 (N_12479,N_11511,N_11169);
xnor U12480 (N_12480,N_11657,N_11717);
or U12481 (N_12481,N_11035,N_11962);
nor U12482 (N_12482,N_11033,N_11982);
nand U12483 (N_12483,N_11282,N_11300);
or U12484 (N_12484,N_11748,N_11860);
xnor U12485 (N_12485,N_11406,N_11784);
or U12486 (N_12486,N_11037,N_11751);
and U12487 (N_12487,N_11257,N_11419);
nor U12488 (N_12488,N_11499,N_11909);
nand U12489 (N_12489,N_11123,N_11807);
nor U12490 (N_12490,N_11292,N_11160);
nor U12491 (N_12491,N_11298,N_11696);
nand U12492 (N_12492,N_11937,N_11279);
nor U12493 (N_12493,N_11260,N_11175);
nand U12494 (N_12494,N_11911,N_11821);
xor U12495 (N_12495,N_11474,N_11879);
nand U12496 (N_12496,N_11452,N_11387);
nor U12497 (N_12497,N_11446,N_11094);
xnor U12498 (N_12498,N_11108,N_11941);
nand U12499 (N_12499,N_11141,N_11904);
or U12500 (N_12500,N_11589,N_11209);
nand U12501 (N_12501,N_11671,N_11515);
or U12502 (N_12502,N_11055,N_11962);
or U12503 (N_12503,N_11959,N_11713);
nor U12504 (N_12504,N_11009,N_11776);
nand U12505 (N_12505,N_11216,N_11967);
nor U12506 (N_12506,N_11437,N_11379);
nor U12507 (N_12507,N_11881,N_11014);
and U12508 (N_12508,N_11027,N_11116);
and U12509 (N_12509,N_11471,N_11295);
or U12510 (N_12510,N_11875,N_11381);
and U12511 (N_12511,N_11001,N_11193);
and U12512 (N_12512,N_11009,N_11108);
and U12513 (N_12513,N_11218,N_11358);
and U12514 (N_12514,N_11714,N_11286);
or U12515 (N_12515,N_11959,N_11829);
nand U12516 (N_12516,N_11583,N_11298);
nor U12517 (N_12517,N_11244,N_11901);
and U12518 (N_12518,N_11217,N_11521);
nand U12519 (N_12519,N_11663,N_11064);
nand U12520 (N_12520,N_11576,N_11920);
xor U12521 (N_12521,N_11875,N_11449);
xnor U12522 (N_12522,N_11112,N_11267);
and U12523 (N_12523,N_11392,N_11550);
xor U12524 (N_12524,N_11250,N_11359);
nand U12525 (N_12525,N_11903,N_11746);
nand U12526 (N_12526,N_11875,N_11467);
and U12527 (N_12527,N_11526,N_11019);
nor U12528 (N_12528,N_11934,N_11831);
nor U12529 (N_12529,N_11987,N_11203);
and U12530 (N_12530,N_11535,N_11688);
nand U12531 (N_12531,N_11238,N_11584);
nor U12532 (N_12532,N_11849,N_11964);
nor U12533 (N_12533,N_11955,N_11561);
or U12534 (N_12534,N_11931,N_11543);
nand U12535 (N_12535,N_11578,N_11939);
nor U12536 (N_12536,N_11908,N_11050);
xor U12537 (N_12537,N_11041,N_11639);
xor U12538 (N_12538,N_11825,N_11961);
nand U12539 (N_12539,N_11231,N_11541);
or U12540 (N_12540,N_11462,N_11876);
or U12541 (N_12541,N_11433,N_11840);
nand U12542 (N_12542,N_11989,N_11540);
or U12543 (N_12543,N_11325,N_11042);
xnor U12544 (N_12544,N_11153,N_11742);
nand U12545 (N_12545,N_11910,N_11603);
nand U12546 (N_12546,N_11816,N_11180);
and U12547 (N_12547,N_11784,N_11658);
nand U12548 (N_12548,N_11019,N_11817);
nand U12549 (N_12549,N_11861,N_11381);
nor U12550 (N_12550,N_11041,N_11272);
xnor U12551 (N_12551,N_11682,N_11257);
and U12552 (N_12552,N_11287,N_11297);
xor U12553 (N_12553,N_11223,N_11402);
xnor U12554 (N_12554,N_11826,N_11117);
or U12555 (N_12555,N_11119,N_11023);
nor U12556 (N_12556,N_11438,N_11201);
or U12557 (N_12557,N_11919,N_11191);
nand U12558 (N_12558,N_11230,N_11583);
nand U12559 (N_12559,N_11563,N_11252);
xnor U12560 (N_12560,N_11814,N_11610);
xnor U12561 (N_12561,N_11537,N_11106);
or U12562 (N_12562,N_11777,N_11873);
nor U12563 (N_12563,N_11747,N_11960);
and U12564 (N_12564,N_11906,N_11763);
or U12565 (N_12565,N_11121,N_11778);
and U12566 (N_12566,N_11083,N_11446);
xor U12567 (N_12567,N_11663,N_11943);
nor U12568 (N_12568,N_11980,N_11181);
and U12569 (N_12569,N_11864,N_11794);
and U12570 (N_12570,N_11409,N_11788);
or U12571 (N_12571,N_11547,N_11029);
or U12572 (N_12572,N_11035,N_11392);
xor U12573 (N_12573,N_11216,N_11400);
xor U12574 (N_12574,N_11748,N_11295);
nor U12575 (N_12575,N_11021,N_11847);
nand U12576 (N_12576,N_11063,N_11154);
and U12577 (N_12577,N_11354,N_11551);
xnor U12578 (N_12578,N_11575,N_11249);
xnor U12579 (N_12579,N_11165,N_11296);
and U12580 (N_12580,N_11435,N_11088);
and U12581 (N_12581,N_11424,N_11150);
nor U12582 (N_12582,N_11184,N_11508);
xor U12583 (N_12583,N_11377,N_11611);
and U12584 (N_12584,N_11968,N_11213);
nor U12585 (N_12585,N_11863,N_11446);
nor U12586 (N_12586,N_11616,N_11250);
nor U12587 (N_12587,N_11771,N_11390);
nand U12588 (N_12588,N_11407,N_11902);
xor U12589 (N_12589,N_11001,N_11588);
xor U12590 (N_12590,N_11274,N_11644);
and U12591 (N_12591,N_11737,N_11008);
xor U12592 (N_12592,N_11466,N_11145);
nor U12593 (N_12593,N_11348,N_11001);
nand U12594 (N_12594,N_11590,N_11111);
nor U12595 (N_12595,N_11151,N_11289);
and U12596 (N_12596,N_11646,N_11089);
or U12597 (N_12597,N_11233,N_11803);
nor U12598 (N_12598,N_11316,N_11680);
and U12599 (N_12599,N_11246,N_11308);
and U12600 (N_12600,N_11071,N_11045);
and U12601 (N_12601,N_11165,N_11014);
and U12602 (N_12602,N_11901,N_11490);
xnor U12603 (N_12603,N_11303,N_11807);
xnor U12604 (N_12604,N_11726,N_11746);
nor U12605 (N_12605,N_11119,N_11789);
or U12606 (N_12606,N_11273,N_11135);
nor U12607 (N_12607,N_11582,N_11700);
or U12608 (N_12608,N_11926,N_11964);
nand U12609 (N_12609,N_11166,N_11228);
nor U12610 (N_12610,N_11098,N_11080);
or U12611 (N_12611,N_11102,N_11754);
nor U12612 (N_12612,N_11511,N_11078);
xnor U12613 (N_12613,N_11068,N_11561);
nor U12614 (N_12614,N_11399,N_11373);
and U12615 (N_12615,N_11271,N_11181);
xor U12616 (N_12616,N_11897,N_11748);
xor U12617 (N_12617,N_11135,N_11895);
xor U12618 (N_12618,N_11698,N_11003);
or U12619 (N_12619,N_11749,N_11036);
nor U12620 (N_12620,N_11298,N_11454);
nand U12621 (N_12621,N_11548,N_11335);
and U12622 (N_12622,N_11115,N_11594);
nand U12623 (N_12623,N_11362,N_11449);
nand U12624 (N_12624,N_11610,N_11739);
and U12625 (N_12625,N_11275,N_11324);
nor U12626 (N_12626,N_11958,N_11770);
xor U12627 (N_12627,N_11342,N_11156);
or U12628 (N_12628,N_11145,N_11816);
xnor U12629 (N_12629,N_11994,N_11767);
or U12630 (N_12630,N_11233,N_11734);
or U12631 (N_12631,N_11419,N_11564);
nand U12632 (N_12632,N_11750,N_11598);
nand U12633 (N_12633,N_11363,N_11903);
xnor U12634 (N_12634,N_11882,N_11174);
nor U12635 (N_12635,N_11801,N_11788);
nor U12636 (N_12636,N_11883,N_11651);
nand U12637 (N_12637,N_11780,N_11707);
nor U12638 (N_12638,N_11373,N_11344);
or U12639 (N_12639,N_11732,N_11304);
nand U12640 (N_12640,N_11660,N_11525);
nor U12641 (N_12641,N_11526,N_11539);
nand U12642 (N_12642,N_11486,N_11352);
or U12643 (N_12643,N_11557,N_11909);
and U12644 (N_12644,N_11172,N_11110);
or U12645 (N_12645,N_11210,N_11836);
nand U12646 (N_12646,N_11474,N_11495);
xor U12647 (N_12647,N_11014,N_11300);
or U12648 (N_12648,N_11741,N_11130);
and U12649 (N_12649,N_11910,N_11295);
nand U12650 (N_12650,N_11603,N_11752);
nand U12651 (N_12651,N_11938,N_11479);
nand U12652 (N_12652,N_11748,N_11928);
or U12653 (N_12653,N_11978,N_11528);
nor U12654 (N_12654,N_11265,N_11432);
or U12655 (N_12655,N_11368,N_11545);
or U12656 (N_12656,N_11966,N_11572);
or U12657 (N_12657,N_11228,N_11894);
or U12658 (N_12658,N_11896,N_11636);
nand U12659 (N_12659,N_11445,N_11017);
and U12660 (N_12660,N_11573,N_11500);
and U12661 (N_12661,N_11012,N_11978);
nand U12662 (N_12662,N_11253,N_11569);
xnor U12663 (N_12663,N_11550,N_11339);
and U12664 (N_12664,N_11777,N_11648);
xnor U12665 (N_12665,N_11562,N_11616);
nor U12666 (N_12666,N_11941,N_11899);
or U12667 (N_12667,N_11277,N_11249);
nor U12668 (N_12668,N_11562,N_11736);
xor U12669 (N_12669,N_11042,N_11377);
or U12670 (N_12670,N_11582,N_11765);
nor U12671 (N_12671,N_11715,N_11855);
nand U12672 (N_12672,N_11063,N_11445);
xnor U12673 (N_12673,N_11304,N_11193);
or U12674 (N_12674,N_11264,N_11175);
xnor U12675 (N_12675,N_11316,N_11643);
xor U12676 (N_12676,N_11473,N_11556);
nand U12677 (N_12677,N_11568,N_11707);
nor U12678 (N_12678,N_11014,N_11833);
or U12679 (N_12679,N_11280,N_11749);
xor U12680 (N_12680,N_11661,N_11380);
or U12681 (N_12681,N_11201,N_11272);
nor U12682 (N_12682,N_11379,N_11694);
nand U12683 (N_12683,N_11127,N_11407);
or U12684 (N_12684,N_11550,N_11682);
xor U12685 (N_12685,N_11632,N_11106);
xnor U12686 (N_12686,N_11952,N_11868);
nand U12687 (N_12687,N_11987,N_11523);
nand U12688 (N_12688,N_11173,N_11086);
xnor U12689 (N_12689,N_11035,N_11048);
or U12690 (N_12690,N_11511,N_11845);
nand U12691 (N_12691,N_11956,N_11424);
nand U12692 (N_12692,N_11021,N_11108);
or U12693 (N_12693,N_11269,N_11811);
or U12694 (N_12694,N_11878,N_11051);
and U12695 (N_12695,N_11165,N_11034);
nand U12696 (N_12696,N_11730,N_11627);
or U12697 (N_12697,N_11791,N_11606);
and U12698 (N_12698,N_11357,N_11444);
nor U12699 (N_12699,N_11321,N_11609);
nor U12700 (N_12700,N_11201,N_11252);
or U12701 (N_12701,N_11207,N_11226);
and U12702 (N_12702,N_11308,N_11456);
nor U12703 (N_12703,N_11321,N_11887);
xor U12704 (N_12704,N_11123,N_11359);
nand U12705 (N_12705,N_11651,N_11732);
nor U12706 (N_12706,N_11053,N_11566);
nor U12707 (N_12707,N_11346,N_11271);
nor U12708 (N_12708,N_11623,N_11194);
nand U12709 (N_12709,N_11145,N_11603);
or U12710 (N_12710,N_11869,N_11934);
nand U12711 (N_12711,N_11731,N_11779);
and U12712 (N_12712,N_11732,N_11085);
nor U12713 (N_12713,N_11253,N_11282);
nand U12714 (N_12714,N_11637,N_11153);
nor U12715 (N_12715,N_11332,N_11572);
nand U12716 (N_12716,N_11464,N_11980);
or U12717 (N_12717,N_11001,N_11051);
nand U12718 (N_12718,N_11150,N_11616);
and U12719 (N_12719,N_11025,N_11955);
and U12720 (N_12720,N_11134,N_11658);
nor U12721 (N_12721,N_11242,N_11402);
nand U12722 (N_12722,N_11767,N_11024);
nand U12723 (N_12723,N_11412,N_11984);
or U12724 (N_12724,N_11917,N_11536);
xnor U12725 (N_12725,N_11919,N_11365);
nor U12726 (N_12726,N_11288,N_11817);
nor U12727 (N_12727,N_11336,N_11923);
nand U12728 (N_12728,N_11495,N_11650);
or U12729 (N_12729,N_11283,N_11121);
xnor U12730 (N_12730,N_11433,N_11438);
or U12731 (N_12731,N_11875,N_11644);
xnor U12732 (N_12732,N_11360,N_11618);
nor U12733 (N_12733,N_11488,N_11936);
or U12734 (N_12734,N_11302,N_11090);
or U12735 (N_12735,N_11123,N_11948);
and U12736 (N_12736,N_11307,N_11519);
nor U12737 (N_12737,N_11089,N_11779);
nor U12738 (N_12738,N_11627,N_11458);
nor U12739 (N_12739,N_11703,N_11051);
nor U12740 (N_12740,N_11385,N_11168);
nand U12741 (N_12741,N_11071,N_11596);
xor U12742 (N_12742,N_11845,N_11242);
nand U12743 (N_12743,N_11327,N_11990);
nor U12744 (N_12744,N_11151,N_11858);
xnor U12745 (N_12745,N_11684,N_11054);
nand U12746 (N_12746,N_11348,N_11674);
and U12747 (N_12747,N_11683,N_11271);
and U12748 (N_12748,N_11592,N_11707);
and U12749 (N_12749,N_11112,N_11786);
and U12750 (N_12750,N_11154,N_11281);
or U12751 (N_12751,N_11753,N_11212);
and U12752 (N_12752,N_11651,N_11404);
nand U12753 (N_12753,N_11192,N_11335);
nor U12754 (N_12754,N_11575,N_11459);
nand U12755 (N_12755,N_11577,N_11036);
or U12756 (N_12756,N_11142,N_11243);
nand U12757 (N_12757,N_11507,N_11203);
xnor U12758 (N_12758,N_11956,N_11885);
or U12759 (N_12759,N_11844,N_11780);
xor U12760 (N_12760,N_11009,N_11085);
or U12761 (N_12761,N_11745,N_11278);
and U12762 (N_12762,N_11651,N_11467);
or U12763 (N_12763,N_11441,N_11711);
nor U12764 (N_12764,N_11082,N_11227);
and U12765 (N_12765,N_11734,N_11410);
nor U12766 (N_12766,N_11725,N_11325);
or U12767 (N_12767,N_11181,N_11508);
or U12768 (N_12768,N_11718,N_11655);
nand U12769 (N_12769,N_11173,N_11871);
or U12770 (N_12770,N_11480,N_11532);
xor U12771 (N_12771,N_11664,N_11960);
or U12772 (N_12772,N_11668,N_11160);
nand U12773 (N_12773,N_11809,N_11738);
xor U12774 (N_12774,N_11881,N_11038);
or U12775 (N_12775,N_11959,N_11988);
nor U12776 (N_12776,N_11276,N_11649);
nand U12777 (N_12777,N_11396,N_11189);
xor U12778 (N_12778,N_11177,N_11893);
nor U12779 (N_12779,N_11401,N_11840);
or U12780 (N_12780,N_11773,N_11851);
nand U12781 (N_12781,N_11950,N_11019);
xnor U12782 (N_12782,N_11328,N_11411);
nor U12783 (N_12783,N_11340,N_11445);
nor U12784 (N_12784,N_11089,N_11269);
or U12785 (N_12785,N_11015,N_11437);
nand U12786 (N_12786,N_11441,N_11677);
or U12787 (N_12787,N_11367,N_11329);
nand U12788 (N_12788,N_11838,N_11361);
nand U12789 (N_12789,N_11442,N_11239);
nor U12790 (N_12790,N_11220,N_11101);
or U12791 (N_12791,N_11141,N_11784);
xnor U12792 (N_12792,N_11896,N_11557);
nand U12793 (N_12793,N_11529,N_11251);
nand U12794 (N_12794,N_11124,N_11316);
xnor U12795 (N_12795,N_11172,N_11589);
nand U12796 (N_12796,N_11308,N_11883);
nor U12797 (N_12797,N_11710,N_11513);
and U12798 (N_12798,N_11786,N_11622);
nand U12799 (N_12799,N_11105,N_11204);
nor U12800 (N_12800,N_11413,N_11079);
and U12801 (N_12801,N_11257,N_11623);
xor U12802 (N_12802,N_11698,N_11759);
xnor U12803 (N_12803,N_11632,N_11767);
nor U12804 (N_12804,N_11341,N_11660);
xnor U12805 (N_12805,N_11749,N_11901);
nor U12806 (N_12806,N_11526,N_11157);
nor U12807 (N_12807,N_11864,N_11950);
nor U12808 (N_12808,N_11155,N_11683);
and U12809 (N_12809,N_11229,N_11211);
and U12810 (N_12810,N_11068,N_11452);
or U12811 (N_12811,N_11347,N_11564);
and U12812 (N_12812,N_11451,N_11617);
nand U12813 (N_12813,N_11372,N_11841);
or U12814 (N_12814,N_11600,N_11116);
nor U12815 (N_12815,N_11965,N_11844);
xnor U12816 (N_12816,N_11037,N_11560);
or U12817 (N_12817,N_11042,N_11302);
nor U12818 (N_12818,N_11185,N_11346);
nand U12819 (N_12819,N_11628,N_11146);
and U12820 (N_12820,N_11276,N_11514);
nand U12821 (N_12821,N_11953,N_11167);
or U12822 (N_12822,N_11324,N_11339);
or U12823 (N_12823,N_11201,N_11870);
xnor U12824 (N_12824,N_11221,N_11966);
and U12825 (N_12825,N_11560,N_11144);
xnor U12826 (N_12826,N_11239,N_11599);
nand U12827 (N_12827,N_11930,N_11452);
and U12828 (N_12828,N_11940,N_11046);
nand U12829 (N_12829,N_11645,N_11017);
and U12830 (N_12830,N_11393,N_11556);
xor U12831 (N_12831,N_11243,N_11575);
nor U12832 (N_12832,N_11578,N_11337);
xor U12833 (N_12833,N_11957,N_11998);
and U12834 (N_12834,N_11806,N_11979);
nor U12835 (N_12835,N_11413,N_11317);
nand U12836 (N_12836,N_11342,N_11648);
and U12837 (N_12837,N_11695,N_11892);
xor U12838 (N_12838,N_11370,N_11980);
nor U12839 (N_12839,N_11816,N_11875);
xnor U12840 (N_12840,N_11357,N_11784);
xor U12841 (N_12841,N_11725,N_11780);
and U12842 (N_12842,N_11222,N_11891);
nor U12843 (N_12843,N_11091,N_11507);
nand U12844 (N_12844,N_11408,N_11443);
xnor U12845 (N_12845,N_11731,N_11906);
xor U12846 (N_12846,N_11353,N_11383);
or U12847 (N_12847,N_11150,N_11401);
and U12848 (N_12848,N_11285,N_11069);
or U12849 (N_12849,N_11626,N_11586);
and U12850 (N_12850,N_11142,N_11203);
nor U12851 (N_12851,N_11398,N_11013);
or U12852 (N_12852,N_11707,N_11284);
nor U12853 (N_12853,N_11668,N_11535);
nor U12854 (N_12854,N_11611,N_11640);
nor U12855 (N_12855,N_11717,N_11400);
or U12856 (N_12856,N_11463,N_11976);
nand U12857 (N_12857,N_11648,N_11136);
or U12858 (N_12858,N_11127,N_11496);
or U12859 (N_12859,N_11862,N_11180);
or U12860 (N_12860,N_11216,N_11077);
nand U12861 (N_12861,N_11546,N_11251);
or U12862 (N_12862,N_11654,N_11241);
or U12863 (N_12863,N_11533,N_11388);
nor U12864 (N_12864,N_11001,N_11412);
nand U12865 (N_12865,N_11695,N_11547);
and U12866 (N_12866,N_11303,N_11126);
nand U12867 (N_12867,N_11835,N_11174);
xnor U12868 (N_12868,N_11815,N_11775);
xor U12869 (N_12869,N_11668,N_11717);
and U12870 (N_12870,N_11771,N_11156);
nand U12871 (N_12871,N_11445,N_11979);
or U12872 (N_12872,N_11424,N_11250);
nor U12873 (N_12873,N_11130,N_11718);
xnor U12874 (N_12874,N_11222,N_11452);
or U12875 (N_12875,N_11641,N_11749);
nand U12876 (N_12876,N_11100,N_11752);
or U12877 (N_12877,N_11463,N_11149);
nor U12878 (N_12878,N_11212,N_11262);
nand U12879 (N_12879,N_11087,N_11567);
nand U12880 (N_12880,N_11192,N_11788);
and U12881 (N_12881,N_11343,N_11635);
nor U12882 (N_12882,N_11071,N_11635);
nand U12883 (N_12883,N_11946,N_11882);
nor U12884 (N_12884,N_11581,N_11160);
nand U12885 (N_12885,N_11736,N_11846);
xor U12886 (N_12886,N_11681,N_11647);
and U12887 (N_12887,N_11116,N_11551);
or U12888 (N_12888,N_11045,N_11942);
xor U12889 (N_12889,N_11796,N_11930);
and U12890 (N_12890,N_11936,N_11685);
nor U12891 (N_12891,N_11454,N_11265);
or U12892 (N_12892,N_11770,N_11714);
xnor U12893 (N_12893,N_11464,N_11817);
xnor U12894 (N_12894,N_11091,N_11931);
xnor U12895 (N_12895,N_11649,N_11244);
nand U12896 (N_12896,N_11650,N_11055);
nand U12897 (N_12897,N_11275,N_11496);
xnor U12898 (N_12898,N_11510,N_11208);
and U12899 (N_12899,N_11155,N_11668);
nand U12900 (N_12900,N_11131,N_11810);
nor U12901 (N_12901,N_11246,N_11544);
or U12902 (N_12902,N_11643,N_11833);
nand U12903 (N_12903,N_11310,N_11995);
nand U12904 (N_12904,N_11427,N_11972);
nor U12905 (N_12905,N_11576,N_11296);
nor U12906 (N_12906,N_11210,N_11348);
xnor U12907 (N_12907,N_11742,N_11052);
nand U12908 (N_12908,N_11847,N_11427);
and U12909 (N_12909,N_11764,N_11894);
xnor U12910 (N_12910,N_11793,N_11582);
nand U12911 (N_12911,N_11946,N_11610);
and U12912 (N_12912,N_11621,N_11231);
xnor U12913 (N_12913,N_11090,N_11718);
nand U12914 (N_12914,N_11275,N_11629);
and U12915 (N_12915,N_11753,N_11660);
xnor U12916 (N_12916,N_11158,N_11721);
nand U12917 (N_12917,N_11507,N_11208);
nor U12918 (N_12918,N_11450,N_11026);
xor U12919 (N_12919,N_11527,N_11304);
or U12920 (N_12920,N_11387,N_11896);
xor U12921 (N_12921,N_11821,N_11336);
nor U12922 (N_12922,N_11584,N_11477);
and U12923 (N_12923,N_11608,N_11446);
nor U12924 (N_12924,N_11136,N_11182);
or U12925 (N_12925,N_11464,N_11326);
and U12926 (N_12926,N_11367,N_11358);
xnor U12927 (N_12927,N_11812,N_11077);
xnor U12928 (N_12928,N_11676,N_11842);
xor U12929 (N_12929,N_11465,N_11050);
nor U12930 (N_12930,N_11646,N_11212);
or U12931 (N_12931,N_11594,N_11815);
or U12932 (N_12932,N_11075,N_11864);
nor U12933 (N_12933,N_11895,N_11203);
nor U12934 (N_12934,N_11295,N_11643);
xor U12935 (N_12935,N_11708,N_11285);
nand U12936 (N_12936,N_11069,N_11459);
nor U12937 (N_12937,N_11430,N_11760);
or U12938 (N_12938,N_11914,N_11390);
nand U12939 (N_12939,N_11612,N_11282);
nand U12940 (N_12940,N_11581,N_11111);
xor U12941 (N_12941,N_11989,N_11017);
and U12942 (N_12942,N_11989,N_11807);
or U12943 (N_12943,N_11506,N_11391);
nand U12944 (N_12944,N_11983,N_11125);
or U12945 (N_12945,N_11973,N_11204);
nand U12946 (N_12946,N_11535,N_11654);
xnor U12947 (N_12947,N_11736,N_11959);
or U12948 (N_12948,N_11857,N_11104);
xnor U12949 (N_12949,N_11316,N_11017);
nor U12950 (N_12950,N_11295,N_11511);
or U12951 (N_12951,N_11668,N_11250);
nand U12952 (N_12952,N_11027,N_11082);
and U12953 (N_12953,N_11700,N_11354);
nor U12954 (N_12954,N_11139,N_11195);
nor U12955 (N_12955,N_11731,N_11189);
nand U12956 (N_12956,N_11959,N_11433);
or U12957 (N_12957,N_11647,N_11418);
and U12958 (N_12958,N_11896,N_11806);
or U12959 (N_12959,N_11734,N_11505);
xor U12960 (N_12960,N_11879,N_11825);
or U12961 (N_12961,N_11011,N_11891);
xor U12962 (N_12962,N_11078,N_11225);
xnor U12963 (N_12963,N_11825,N_11188);
or U12964 (N_12964,N_11241,N_11912);
nand U12965 (N_12965,N_11995,N_11984);
and U12966 (N_12966,N_11950,N_11430);
or U12967 (N_12967,N_11405,N_11104);
nand U12968 (N_12968,N_11497,N_11072);
xor U12969 (N_12969,N_11541,N_11697);
xnor U12970 (N_12970,N_11561,N_11906);
nor U12971 (N_12971,N_11702,N_11721);
nor U12972 (N_12972,N_11424,N_11610);
and U12973 (N_12973,N_11491,N_11531);
and U12974 (N_12974,N_11320,N_11893);
xor U12975 (N_12975,N_11337,N_11328);
nand U12976 (N_12976,N_11288,N_11969);
nor U12977 (N_12977,N_11962,N_11301);
xnor U12978 (N_12978,N_11381,N_11185);
and U12979 (N_12979,N_11061,N_11612);
and U12980 (N_12980,N_11261,N_11766);
nand U12981 (N_12981,N_11976,N_11642);
nand U12982 (N_12982,N_11942,N_11435);
and U12983 (N_12983,N_11588,N_11684);
nor U12984 (N_12984,N_11788,N_11967);
nand U12985 (N_12985,N_11818,N_11932);
or U12986 (N_12986,N_11713,N_11198);
nand U12987 (N_12987,N_11678,N_11395);
and U12988 (N_12988,N_11850,N_11778);
and U12989 (N_12989,N_11771,N_11317);
or U12990 (N_12990,N_11610,N_11975);
xnor U12991 (N_12991,N_11441,N_11248);
or U12992 (N_12992,N_11963,N_11624);
or U12993 (N_12993,N_11392,N_11983);
xor U12994 (N_12994,N_11431,N_11467);
nand U12995 (N_12995,N_11596,N_11208);
and U12996 (N_12996,N_11603,N_11295);
and U12997 (N_12997,N_11377,N_11886);
nand U12998 (N_12998,N_11562,N_11288);
nor U12999 (N_12999,N_11270,N_11207);
nand U13000 (N_13000,N_12570,N_12996);
or U13001 (N_13001,N_12291,N_12511);
nand U13002 (N_13002,N_12114,N_12587);
and U13003 (N_13003,N_12762,N_12653);
xor U13004 (N_13004,N_12021,N_12728);
xor U13005 (N_13005,N_12068,N_12669);
nor U13006 (N_13006,N_12843,N_12520);
nor U13007 (N_13007,N_12585,N_12834);
xor U13008 (N_13008,N_12503,N_12253);
nor U13009 (N_13009,N_12213,N_12255);
nand U13010 (N_13010,N_12647,N_12527);
or U13011 (N_13011,N_12613,N_12096);
or U13012 (N_13012,N_12284,N_12407);
nand U13013 (N_13013,N_12897,N_12808);
or U13014 (N_13014,N_12107,N_12494);
nand U13015 (N_13015,N_12868,N_12374);
nor U13016 (N_13016,N_12203,N_12964);
xor U13017 (N_13017,N_12058,N_12634);
nand U13018 (N_13018,N_12844,N_12989);
or U13019 (N_13019,N_12973,N_12557);
and U13020 (N_13020,N_12912,N_12629);
nor U13021 (N_13021,N_12856,N_12947);
or U13022 (N_13022,N_12162,N_12283);
nand U13023 (N_13023,N_12375,N_12645);
xor U13024 (N_13024,N_12098,N_12157);
xor U13025 (N_13025,N_12811,N_12339);
nand U13026 (N_13026,N_12313,N_12217);
xnor U13027 (N_13027,N_12774,N_12396);
or U13028 (N_13028,N_12499,N_12441);
nand U13029 (N_13029,N_12818,N_12332);
or U13030 (N_13030,N_12477,N_12931);
nor U13031 (N_13031,N_12467,N_12508);
and U13032 (N_13032,N_12362,N_12517);
and U13033 (N_13033,N_12817,N_12803);
nand U13034 (N_13034,N_12319,N_12836);
xnor U13035 (N_13035,N_12016,N_12501);
and U13036 (N_13036,N_12541,N_12397);
xor U13037 (N_13037,N_12698,N_12143);
xnor U13038 (N_13038,N_12750,N_12936);
and U13039 (N_13039,N_12672,N_12083);
xor U13040 (N_13040,N_12516,N_12558);
and U13041 (N_13041,N_12932,N_12318);
nor U13042 (N_13042,N_12500,N_12040);
or U13043 (N_13043,N_12982,N_12150);
xnor U13044 (N_13044,N_12457,N_12333);
xnor U13045 (N_13045,N_12350,N_12458);
nor U13046 (N_13046,N_12109,N_12713);
nand U13047 (N_13047,N_12343,N_12617);
nor U13048 (N_13048,N_12166,N_12665);
and U13049 (N_13049,N_12430,N_12799);
or U13050 (N_13050,N_12925,N_12418);
nand U13051 (N_13051,N_12227,N_12814);
nor U13052 (N_13052,N_12215,N_12905);
or U13053 (N_13053,N_12990,N_12384);
nor U13054 (N_13054,N_12195,N_12697);
xnor U13055 (N_13055,N_12102,N_12340);
xor U13056 (N_13056,N_12294,N_12743);
xor U13057 (N_13057,N_12572,N_12346);
or U13058 (N_13058,N_12940,N_12254);
xnor U13059 (N_13059,N_12059,N_12046);
and U13060 (N_13060,N_12067,N_12325);
nand U13061 (N_13061,N_12639,N_12322);
nor U13062 (N_13062,N_12405,N_12413);
nand U13063 (N_13063,N_12012,N_12184);
xor U13064 (N_13064,N_12221,N_12079);
nand U13065 (N_13065,N_12116,N_12507);
xnor U13066 (N_13066,N_12180,N_12171);
nand U13067 (N_13067,N_12474,N_12419);
nand U13068 (N_13068,N_12773,N_12351);
or U13069 (N_13069,N_12509,N_12937);
or U13070 (N_13070,N_12190,N_12770);
xor U13071 (N_13071,N_12382,N_12226);
nand U13072 (N_13072,N_12565,N_12798);
xnor U13073 (N_13073,N_12013,N_12666);
xor U13074 (N_13074,N_12555,N_12801);
nor U13075 (N_13075,N_12251,N_12686);
xor U13076 (N_13076,N_12906,N_12780);
xor U13077 (N_13077,N_12510,N_12470);
nand U13078 (N_13078,N_12719,N_12212);
and U13079 (N_13079,N_12584,N_12734);
and U13080 (N_13080,N_12658,N_12688);
xnor U13081 (N_13081,N_12775,N_12939);
nand U13082 (N_13082,N_12514,N_12469);
xnor U13083 (N_13083,N_12691,N_12409);
nand U13084 (N_13084,N_12546,N_12327);
nand U13085 (N_13085,N_12700,N_12614);
nor U13086 (N_13086,N_12204,N_12824);
and U13087 (N_13087,N_12442,N_12471);
xnor U13088 (N_13088,N_12263,N_12256);
nand U13089 (N_13089,N_12378,N_12001);
xor U13090 (N_13090,N_12276,N_12929);
or U13091 (N_13091,N_12337,N_12249);
nor U13092 (N_13092,N_12523,N_12224);
nand U13093 (N_13093,N_12790,N_12135);
xnor U13094 (N_13094,N_12596,N_12417);
and U13095 (N_13095,N_12659,N_12085);
xnor U13096 (N_13096,N_12571,N_12926);
and U13097 (N_13097,N_12784,N_12475);
or U13098 (N_13098,N_12705,N_12815);
xor U13099 (N_13099,N_12176,N_12125);
xnor U13100 (N_13100,N_12307,N_12336);
nor U13101 (N_13101,N_12359,N_12954);
nor U13102 (N_13102,N_12353,N_12090);
xnor U13103 (N_13103,N_12295,N_12866);
or U13104 (N_13104,N_12859,N_12789);
and U13105 (N_13105,N_12449,N_12450);
nor U13106 (N_13106,N_12308,N_12826);
xnor U13107 (N_13107,N_12694,N_12317);
and U13108 (N_13108,N_12388,N_12802);
and U13109 (N_13109,N_12660,N_12064);
nand U13110 (N_13110,N_12074,N_12497);
and U13111 (N_13111,N_12118,N_12676);
xnor U13112 (N_13112,N_12273,N_12505);
nor U13113 (N_13113,N_12537,N_12881);
nor U13114 (N_13114,N_12345,N_12722);
nor U13115 (N_13115,N_12515,N_12717);
xor U13116 (N_13116,N_12875,N_12163);
nand U13117 (N_13117,N_12731,N_12039);
and U13118 (N_13118,N_12197,N_12385);
nor U13119 (N_13119,N_12795,N_12214);
xor U13120 (N_13120,N_12753,N_12895);
nor U13121 (N_13121,N_12105,N_12211);
or U13122 (N_13122,N_12923,N_12946);
xor U13123 (N_13123,N_12618,N_12243);
nor U13124 (N_13124,N_12987,N_12855);
nand U13125 (N_13125,N_12806,N_12431);
xor U13126 (N_13126,N_12029,N_12193);
and U13127 (N_13127,N_12194,N_12447);
and U13128 (N_13128,N_12955,N_12683);
or U13129 (N_13129,N_12225,N_12573);
nand U13130 (N_13130,N_12230,N_12741);
nor U13131 (N_13131,N_12463,N_12680);
and U13132 (N_13132,N_12594,N_12246);
or U13133 (N_13133,N_12348,N_12275);
and U13134 (N_13134,N_12129,N_12662);
and U13135 (N_13135,N_12257,N_12455);
and U13136 (N_13136,N_12192,N_12592);
nand U13137 (N_13137,N_12637,N_12465);
or U13138 (N_13138,N_12828,N_12266);
nor U13139 (N_13139,N_12055,N_12742);
nand U13140 (N_13140,N_12380,N_12078);
or U13141 (N_13141,N_12354,N_12739);
and U13142 (N_13142,N_12299,N_12286);
xnor U13143 (N_13143,N_12562,N_12586);
nor U13144 (N_13144,N_12402,N_12981);
or U13145 (N_13145,N_12916,N_12406);
xnor U13146 (N_13146,N_12858,N_12347);
and U13147 (N_13147,N_12481,N_12525);
or U13148 (N_13148,N_12498,N_12485);
and U13149 (N_13149,N_12646,N_12974);
nor U13150 (N_13150,N_12518,N_12149);
xnor U13151 (N_13151,N_12771,N_12349);
nand U13152 (N_13152,N_12324,N_12264);
or U13153 (N_13153,N_12321,N_12306);
nor U13154 (N_13154,N_12595,N_12600);
nor U13155 (N_13155,N_12651,N_12123);
and U13156 (N_13156,N_12502,N_12769);
or U13157 (N_13157,N_12599,N_12445);
nor U13158 (N_13158,N_12994,N_12311);
nand U13159 (N_13159,N_12182,N_12785);
nor U13160 (N_13160,N_12876,N_12809);
or U13161 (N_13161,N_12603,N_12052);
or U13162 (N_13162,N_12464,N_12673);
nand U13163 (N_13163,N_12484,N_12297);
xor U13164 (N_13164,N_12708,N_12443);
and U13165 (N_13165,N_12038,N_12604);
and U13166 (N_13166,N_12577,N_12159);
nor U13167 (N_13167,N_12652,N_12877);
and U13168 (N_13168,N_12127,N_12301);
and U13169 (N_13169,N_12018,N_12490);
nor U13170 (N_13170,N_12810,N_12144);
nor U13171 (N_13171,N_12696,N_12941);
or U13172 (N_13172,N_12715,N_12179);
xor U13173 (N_13173,N_12681,N_12846);
xnor U13174 (N_13174,N_12272,N_12909);
nor U13175 (N_13175,N_12609,N_12986);
and U13176 (N_13176,N_12482,N_12426);
xnor U13177 (N_13177,N_12066,N_12328);
nor U13178 (N_13178,N_12737,N_12712);
and U13179 (N_13179,N_12980,N_12838);
nand U13180 (N_13180,N_12433,N_12685);
xnor U13181 (N_13181,N_12099,N_12796);
nand U13182 (N_13182,N_12383,N_12667);
xnor U13183 (N_13183,N_12574,N_12285);
or U13184 (N_13184,N_12977,N_12261);
or U13185 (N_13185,N_12034,N_12232);
xnor U13186 (N_13186,N_12216,N_12030);
xnor U13187 (N_13187,N_12593,N_12804);
nand U13188 (N_13188,N_12746,N_12128);
nand U13189 (N_13189,N_12281,N_12335);
and U13190 (N_13190,N_12424,N_12521);
nand U13191 (N_13191,N_12528,N_12080);
xnor U13192 (N_13192,N_12334,N_12398);
or U13193 (N_13193,N_12854,N_12188);
xor U13194 (N_13194,N_12205,N_12893);
or U13195 (N_13195,N_12120,N_12917);
nor U13196 (N_13196,N_12124,N_12438);
nand U13197 (N_13197,N_12690,N_12002);
and U13198 (N_13198,N_12744,N_12037);
or U13199 (N_13199,N_12111,N_12958);
xor U13200 (N_13200,N_12053,N_12057);
and U13201 (N_13201,N_12601,N_12401);
nor U13202 (N_13202,N_12569,N_12265);
xnor U13203 (N_13203,N_12807,N_12891);
nand U13204 (N_13204,N_12131,N_12874);
and U13205 (N_13205,N_12506,N_12394);
nand U13206 (N_13206,N_12693,N_12414);
and U13207 (N_13207,N_12865,N_12644);
and U13208 (N_13208,N_12429,N_12260);
nand U13209 (N_13209,N_12439,N_12165);
xnor U13210 (N_13210,N_12456,N_12371);
nor U13211 (N_13211,N_12671,N_12864);
xor U13212 (N_13212,N_12091,N_12183);
nand U13213 (N_13213,N_12886,N_12145);
and U13214 (N_13214,N_12615,N_12075);
or U13215 (N_13215,N_12692,N_12970);
nor U13216 (N_13216,N_12702,N_12787);
nand U13217 (N_13217,N_12041,N_12269);
and U13218 (N_13218,N_12472,N_12062);
nor U13219 (N_13219,N_12797,N_12331);
nand U13220 (N_13220,N_12461,N_12271);
and U13221 (N_13221,N_12373,N_12077);
or U13222 (N_13222,N_12309,N_12952);
or U13223 (N_13223,N_12675,N_12218);
and U13224 (N_13224,N_12329,N_12048);
or U13225 (N_13225,N_12556,N_12655);
xor U13226 (N_13226,N_12454,N_12137);
xnor U13227 (N_13227,N_12519,N_12017);
xor U13228 (N_13228,N_12612,N_12819);
and U13229 (N_13229,N_12065,N_12201);
xor U13230 (N_13230,N_12045,N_12303);
or U13231 (N_13231,N_12704,N_12151);
xor U13232 (N_13232,N_12544,N_12154);
and U13233 (N_13233,N_12907,N_12852);
or U13234 (N_13234,N_12718,N_12765);
nor U13235 (N_13235,N_12567,N_12878);
or U13236 (N_13236,N_12033,N_12689);
xor U13237 (N_13237,N_12342,N_12626);
xnor U13238 (N_13238,N_12156,N_12060);
nor U13239 (N_13239,N_12606,N_12316);
xor U13240 (N_13240,N_12983,N_12219);
or U13241 (N_13241,N_12736,N_12582);
or U13242 (N_13242,N_12579,N_12435);
xor U13243 (N_13243,N_12976,N_12238);
nor U13244 (N_13244,N_12022,N_12234);
nor U13245 (N_13245,N_12270,N_12492);
nor U13246 (N_13246,N_12842,N_12978);
xor U13247 (N_13247,N_12024,N_12493);
nand U13248 (N_13248,N_12522,N_12504);
nor U13249 (N_13249,N_12436,N_12312);
nand U13250 (N_13250,N_12568,N_12229);
and U13251 (N_13251,N_12813,N_12816);
nand U13252 (N_13252,N_12108,N_12870);
nand U13253 (N_13253,N_12512,N_12368);
nor U13254 (N_13254,N_12185,N_12140);
and U13255 (N_13255,N_12551,N_12539);
nor U13256 (N_13256,N_12478,N_12235);
nand U13257 (N_13257,N_12250,N_12622);
or U13258 (N_13258,N_12241,N_12513);
nor U13259 (N_13259,N_12141,N_12158);
or U13260 (N_13260,N_12302,N_12921);
nand U13261 (N_13261,N_12126,N_12489);
or U13262 (N_13262,N_12869,N_12277);
nor U13263 (N_13263,N_12026,N_12290);
and U13264 (N_13264,N_12061,N_12621);
and U13265 (N_13265,N_12751,N_12670);
nand U13266 (N_13266,N_12699,N_12892);
nor U13267 (N_13267,N_12081,N_12729);
and U13268 (N_13268,N_12186,N_12563);
nor U13269 (N_13269,N_12187,N_12304);
nand U13270 (N_13270,N_12636,N_12259);
or U13271 (N_13271,N_12360,N_12935);
or U13272 (N_13272,N_12355,N_12677);
and U13273 (N_13273,N_12679,N_12831);
nand U13274 (N_13274,N_12829,N_12850);
and U13275 (N_13275,N_12293,N_12000);
nor U13276 (N_13276,N_12781,N_12625);
nor U13277 (N_13277,N_12928,N_12920);
nand U13278 (N_13278,N_12155,N_12133);
or U13279 (N_13279,N_12548,N_12641);
nand U13280 (N_13280,N_12530,N_12997);
xor U13281 (N_13281,N_12369,N_12460);
nand U13282 (N_13282,N_12879,N_12386);
or U13283 (N_13283,N_12027,N_12998);
and U13284 (N_13284,N_12487,N_12404);
xor U13285 (N_13285,N_12962,N_12341);
or U13286 (N_13286,N_12242,N_12389);
xor U13287 (N_13287,N_12300,N_12451);
or U13288 (N_13288,N_12376,N_12411);
nor U13289 (N_13289,N_12791,N_12757);
or U13290 (N_13290,N_12610,N_12993);
nand U13291 (N_13291,N_12305,N_12915);
nor U13292 (N_13292,N_12483,N_12209);
nor U13293 (N_13293,N_12545,N_12961);
nand U13294 (N_13294,N_12589,N_12486);
nand U13295 (N_13295,N_12934,N_12930);
nor U13296 (N_13296,N_12848,N_12367);
nand U13297 (N_13297,N_12086,N_12153);
xor U13298 (N_13298,N_12160,N_12009);
xnor U13299 (N_13299,N_12248,N_12540);
nor U13300 (N_13300,N_12616,N_12082);
nor U13301 (N_13301,N_12132,N_12536);
nor U13302 (N_13302,N_12758,N_12421);
xnor U13303 (N_13303,N_12198,N_12550);
nand U13304 (N_13304,N_12890,N_12245);
and U13305 (N_13305,N_12377,N_12338);
or U13306 (N_13306,N_12535,N_12172);
xor U13307 (N_13307,N_12995,N_12358);
or U13308 (N_13308,N_12752,N_12788);
xor U13309 (N_13309,N_12278,N_12533);
or U13310 (N_13310,N_12361,N_12170);
xnor U13311 (N_13311,N_12965,N_12709);
or U13312 (N_13312,N_12792,N_12168);
nand U13313 (N_13313,N_12944,N_12624);
nand U13314 (N_13314,N_12656,N_12553);
nor U13315 (N_13315,N_12089,N_12725);
or U13316 (N_13316,N_12006,N_12820);
xor U13317 (N_13317,N_12244,N_12237);
and U13318 (N_13318,N_12889,N_12674);
nor U13319 (N_13319,N_12400,N_12607);
nor U13320 (N_13320,N_12833,N_12069);
and U13321 (N_13321,N_12867,N_12236);
nand U13322 (N_13322,N_12044,N_12650);
nand U13323 (N_13323,N_12764,N_12444);
nand U13324 (N_13324,N_12730,N_12035);
or U13325 (N_13325,N_12914,N_12768);
nor U13326 (N_13326,N_12957,N_12608);
and U13327 (N_13327,N_12142,N_12072);
nor U13328 (N_13328,N_12543,N_12760);
nand U13329 (N_13329,N_12560,N_12630);
xnor U13330 (N_13330,N_12476,N_12365);
nor U13331 (N_13331,N_12779,N_12605);
nor U13332 (N_13332,N_12191,N_12206);
or U13333 (N_13333,N_12279,N_12363);
nor U13334 (N_13334,N_12706,N_12590);
nand U13335 (N_13335,N_12851,N_12588);
nor U13336 (N_13336,N_12177,N_12972);
nor U13337 (N_13337,N_12231,N_12181);
nand U13338 (N_13338,N_12748,N_12196);
and U13339 (N_13339,N_12975,N_12761);
and U13340 (N_13340,N_12938,N_12529);
nand U13341 (N_13341,N_12822,N_12777);
or U13342 (N_13342,N_12036,N_12434);
nor U13343 (N_13343,N_12364,N_12979);
or U13344 (N_13344,N_12247,N_12152);
nand U13345 (N_13345,N_12884,N_12448);
xnor U13346 (N_13346,N_12724,N_12664);
nand U13347 (N_13347,N_12745,N_12580);
or U13348 (N_13348,N_12922,N_12711);
nand U13349 (N_13349,N_12678,N_12025);
nor U13350 (N_13350,N_12805,N_12392);
nand U13351 (N_13351,N_12684,N_12948);
and U13352 (N_13352,N_12391,N_12416);
xor U13353 (N_13353,N_12619,N_12583);
nor U13354 (N_13354,N_12871,N_12552);
and U13355 (N_13355,N_12960,N_12648);
or U13356 (N_13356,N_12880,N_12554);
xnor U13357 (N_13357,N_12898,N_12425);
or U13358 (N_13358,N_12959,N_12110);
nand U13359 (N_13359,N_12491,N_12575);
xnor U13360 (N_13360,N_12468,N_12668);
nand U13361 (N_13361,N_12410,N_12070);
or U13362 (N_13362,N_12913,N_12412);
nand U13363 (N_13363,N_12032,N_12296);
xnor U13364 (N_13364,N_12106,N_12985);
nor U13365 (N_13365,N_12175,N_12902);
xor U13366 (N_13366,N_12314,N_12632);
xnor U13367 (N_13367,N_12904,N_12657);
nand U13368 (N_13368,N_12682,N_12462);
and U13369 (N_13369,N_12357,N_12597);
xnor U13370 (N_13370,N_12031,N_12428);
nor U13371 (N_13371,N_12095,N_12274);
nand U13372 (N_13372,N_12547,N_12950);
nor U13373 (N_13373,N_12703,N_12687);
xnor U13374 (N_13374,N_12390,N_12863);
and U13375 (N_13375,N_12559,N_12427);
nor U13376 (N_13376,N_12210,N_12113);
or U13377 (N_13377,N_12759,N_12049);
and U13378 (N_13378,N_12763,N_12812);
nand U13379 (N_13379,N_12130,N_12740);
and U13380 (N_13380,N_12782,N_12051);
and U13381 (N_13381,N_12956,N_12716);
nand U13382 (N_13382,N_12860,N_12918);
xnor U13383 (N_13383,N_12161,N_12887);
nand U13384 (N_13384,N_12872,N_12097);
nand U13385 (N_13385,N_12654,N_12847);
or U13386 (N_13386,N_12087,N_12991);
nand U13387 (N_13387,N_12169,N_12043);
nor U13388 (N_13388,N_12623,N_12310);
nand U13389 (N_13389,N_12849,N_12640);
nor U13390 (N_13390,N_12092,N_12823);
and U13391 (N_13391,N_12873,N_12453);
xnor U13392 (N_13392,N_12800,N_12208);
nand U13393 (N_13393,N_12945,N_12240);
xor U13394 (N_13394,N_12627,N_12054);
nand U13395 (N_13395,N_12258,N_12220);
nor U13396 (N_13396,N_12942,N_12119);
nand U13397 (N_13397,N_12015,N_12289);
and U13398 (N_13398,N_12073,N_12786);
and U13399 (N_13399,N_12422,N_12825);
and U13400 (N_13400,N_12199,N_12888);
nand U13401 (N_13401,N_12933,N_12984);
nor U13402 (N_13402,N_12628,N_12840);
or U13403 (N_13403,N_12381,N_12200);
xor U13404 (N_13404,N_12901,N_12710);
xnor U13405 (N_13405,N_12766,N_12727);
and U13406 (N_13406,N_12134,N_12927);
or U13407 (N_13407,N_12794,N_12581);
or U13408 (N_13408,N_12011,N_12479);
nand U13409 (N_13409,N_12720,N_12830);
or U13410 (N_13410,N_12835,N_12738);
and U13411 (N_13411,N_12366,N_12268);
or U13412 (N_13412,N_12862,N_12028);
nor U13413 (N_13413,N_12020,N_12056);
xor U13414 (N_13414,N_12415,N_12999);
and U13415 (N_13415,N_12591,N_12003);
or U13416 (N_13416,N_12004,N_12735);
nand U13417 (N_13417,N_12047,N_12370);
and U13418 (N_13418,N_12459,N_12178);
nor U13419 (N_13419,N_12222,N_12233);
xnor U13420 (N_13420,N_12146,N_12164);
and U13421 (N_13421,N_12023,N_12971);
or U13422 (N_13422,N_12423,N_12910);
and U13423 (N_13423,N_12420,N_12701);
nor U13424 (N_13424,N_12620,N_12841);
and U13425 (N_13425,N_12756,N_12282);
nor U13426 (N_13426,N_12919,N_12298);
nor U13427 (N_13427,N_12578,N_12943);
and U13428 (N_13428,N_12267,N_12532);
and U13429 (N_13429,N_12951,N_12496);
nor U13430 (N_13430,N_12292,N_12372);
nand U13431 (N_13431,N_12598,N_12440);
xnor U13432 (N_13432,N_12063,N_12772);
and U13433 (N_13433,N_12323,N_12076);
and U13434 (N_13434,N_12894,N_12963);
or U13435 (N_13435,N_12949,N_12122);
or U13436 (N_13436,N_12320,N_12395);
xnor U13437 (N_13437,N_12908,N_12403);
nor U13438 (N_13438,N_12988,N_12531);
nand U13439 (N_13439,N_12561,N_12538);
xnor U13440 (N_13440,N_12602,N_12262);
xnor U13441 (N_13441,N_12857,N_12139);
xor U13442 (N_13442,N_12393,N_12007);
or U13443 (N_13443,N_12189,N_12723);
nor U13444 (N_13444,N_12352,N_12534);
xor U13445 (N_13445,N_12642,N_12911);
xor U13446 (N_13446,N_12138,N_12326);
or U13447 (N_13447,N_12387,N_12721);
or U13448 (N_13448,N_12754,N_12549);
or U13449 (N_13449,N_12287,N_12084);
xnor U13450 (N_13450,N_12631,N_12526);
nor U13451 (N_13451,N_12638,N_12953);
nor U13452 (N_13452,N_12473,N_12408);
xnor U13453 (N_13453,N_12432,N_12564);
nor U13454 (N_13454,N_12399,N_12695);
xor U13455 (N_13455,N_12566,N_12117);
and U13456 (N_13456,N_12755,N_12732);
or U13457 (N_13457,N_12207,N_12280);
nor U13458 (N_13458,N_12480,N_12356);
xor U13459 (N_13459,N_12853,N_12966);
xor U13460 (N_13460,N_12252,N_12778);
and U13461 (N_13461,N_12147,N_12707);
nor U13462 (N_13462,N_12832,N_12733);
and U13463 (N_13463,N_12749,N_12005);
or U13464 (N_13464,N_12845,N_12542);
and U13465 (N_13465,N_12315,N_12992);
nor U13466 (N_13466,N_12896,N_12969);
xor U13467 (N_13467,N_12094,N_12783);
or U13468 (N_13468,N_12330,N_12202);
nor U13469 (N_13469,N_12767,N_12611);
nor U13470 (N_13470,N_12173,N_12167);
nor U13471 (N_13471,N_12288,N_12223);
or U13472 (N_13472,N_12101,N_12344);
xor U13473 (N_13473,N_12228,N_12714);
or U13474 (N_13474,N_12633,N_12882);
xor U13475 (N_13475,N_12649,N_12466);
xor U13476 (N_13476,N_12924,N_12239);
or U13477 (N_13477,N_12121,N_12014);
xnor U13478 (N_13478,N_12821,N_12839);
xnor U13479 (N_13479,N_12071,N_12663);
xor U13480 (N_13480,N_12661,N_12576);
and U13481 (N_13481,N_12136,N_12635);
or U13482 (N_13482,N_12643,N_12827);
or U13483 (N_13483,N_12010,N_12899);
nand U13484 (N_13484,N_12883,N_12967);
xor U13485 (N_13485,N_12793,N_12488);
and U13486 (N_13486,N_12008,N_12042);
xnor U13487 (N_13487,N_12903,N_12452);
xor U13488 (N_13488,N_12174,N_12050);
xor U13489 (N_13489,N_12437,N_12861);
nand U13490 (N_13490,N_12837,N_12100);
and U13491 (N_13491,N_12019,N_12900);
nand U13492 (N_13492,N_12093,N_12776);
nand U13493 (N_13493,N_12379,N_12885);
or U13494 (N_13494,N_12747,N_12088);
nand U13495 (N_13495,N_12446,N_12104);
nor U13496 (N_13496,N_12524,N_12112);
and U13497 (N_13497,N_12148,N_12103);
and U13498 (N_13498,N_12115,N_12495);
or U13499 (N_13499,N_12726,N_12968);
and U13500 (N_13500,N_12025,N_12922);
nand U13501 (N_13501,N_12597,N_12903);
or U13502 (N_13502,N_12557,N_12988);
and U13503 (N_13503,N_12004,N_12415);
and U13504 (N_13504,N_12590,N_12013);
and U13505 (N_13505,N_12122,N_12397);
xor U13506 (N_13506,N_12474,N_12976);
or U13507 (N_13507,N_12267,N_12865);
nor U13508 (N_13508,N_12843,N_12108);
xnor U13509 (N_13509,N_12541,N_12385);
xnor U13510 (N_13510,N_12097,N_12315);
nor U13511 (N_13511,N_12629,N_12340);
or U13512 (N_13512,N_12166,N_12251);
nand U13513 (N_13513,N_12818,N_12959);
and U13514 (N_13514,N_12983,N_12629);
or U13515 (N_13515,N_12644,N_12825);
xnor U13516 (N_13516,N_12528,N_12950);
nor U13517 (N_13517,N_12411,N_12699);
or U13518 (N_13518,N_12532,N_12557);
or U13519 (N_13519,N_12947,N_12006);
xor U13520 (N_13520,N_12899,N_12074);
or U13521 (N_13521,N_12077,N_12432);
and U13522 (N_13522,N_12392,N_12293);
nand U13523 (N_13523,N_12515,N_12317);
nand U13524 (N_13524,N_12892,N_12431);
or U13525 (N_13525,N_12868,N_12844);
nor U13526 (N_13526,N_12682,N_12822);
nand U13527 (N_13527,N_12917,N_12430);
xnor U13528 (N_13528,N_12993,N_12312);
and U13529 (N_13529,N_12424,N_12358);
and U13530 (N_13530,N_12438,N_12262);
nor U13531 (N_13531,N_12182,N_12358);
and U13532 (N_13532,N_12333,N_12572);
xnor U13533 (N_13533,N_12252,N_12624);
nor U13534 (N_13534,N_12933,N_12165);
and U13535 (N_13535,N_12711,N_12205);
nand U13536 (N_13536,N_12497,N_12122);
xor U13537 (N_13537,N_12576,N_12991);
nand U13538 (N_13538,N_12044,N_12580);
nand U13539 (N_13539,N_12779,N_12707);
xnor U13540 (N_13540,N_12353,N_12501);
nor U13541 (N_13541,N_12567,N_12352);
nand U13542 (N_13542,N_12129,N_12146);
or U13543 (N_13543,N_12273,N_12500);
or U13544 (N_13544,N_12188,N_12829);
nor U13545 (N_13545,N_12003,N_12601);
and U13546 (N_13546,N_12005,N_12819);
nand U13547 (N_13547,N_12900,N_12683);
nor U13548 (N_13548,N_12800,N_12981);
or U13549 (N_13549,N_12016,N_12724);
and U13550 (N_13550,N_12435,N_12895);
and U13551 (N_13551,N_12042,N_12364);
xor U13552 (N_13552,N_12053,N_12596);
nor U13553 (N_13553,N_12569,N_12628);
nor U13554 (N_13554,N_12937,N_12444);
nand U13555 (N_13555,N_12367,N_12435);
nand U13556 (N_13556,N_12763,N_12271);
xor U13557 (N_13557,N_12228,N_12836);
nand U13558 (N_13558,N_12176,N_12845);
nand U13559 (N_13559,N_12833,N_12307);
and U13560 (N_13560,N_12721,N_12101);
xor U13561 (N_13561,N_12505,N_12594);
nor U13562 (N_13562,N_12472,N_12438);
nor U13563 (N_13563,N_12374,N_12024);
and U13564 (N_13564,N_12331,N_12729);
nand U13565 (N_13565,N_12032,N_12412);
nand U13566 (N_13566,N_12041,N_12633);
nor U13567 (N_13567,N_12887,N_12853);
or U13568 (N_13568,N_12982,N_12958);
nor U13569 (N_13569,N_12677,N_12090);
nor U13570 (N_13570,N_12307,N_12233);
nand U13571 (N_13571,N_12219,N_12949);
and U13572 (N_13572,N_12906,N_12764);
nor U13573 (N_13573,N_12848,N_12461);
xnor U13574 (N_13574,N_12589,N_12715);
nand U13575 (N_13575,N_12876,N_12325);
or U13576 (N_13576,N_12864,N_12432);
or U13577 (N_13577,N_12965,N_12619);
or U13578 (N_13578,N_12284,N_12918);
and U13579 (N_13579,N_12193,N_12468);
or U13580 (N_13580,N_12883,N_12374);
and U13581 (N_13581,N_12558,N_12813);
nand U13582 (N_13582,N_12769,N_12036);
or U13583 (N_13583,N_12139,N_12764);
nor U13584 (N_13584,N_12736,N_12964);
nor U13585 (N_13585,N_12513,N_12224);
nor U13586 (N_13586,N_12814,N_12337);
nor U13587 (N_13587,N_12239,N_12000);
nor U13588 (N_13588,N_12919,N_12263);
xnor U13589 (N_13589,N_12454,N_12297);
or U13590 (N_13590,N_12012,N_12617);
nor U13591 (N_13591,N_12930,N_12845);
nand U13592 (N_13592,N_12050,N_12782);
xor U13593 (N_13593,N_12022,N_12489);
nor U13594 (N_13594,N_12048,N_12238);
or U13595 (N_13595,N_12312,N_12523);
nand U13596 (N_13596,N_12704,N_12689);
nor U13597 (N_13597,N_12729,N_12501);
xor U13598 (N_13598,N_12270,N_12917);
xor U13599 (N_13599,N_12011,N_12950);
nand U13600 (N_13600,N_12810,N_12988);
nand U13601 (N_13601,N_12070,N_12237);
nor U13602 (N_13602,N_12395,N_12246);
xor U13603 (N_13603,N_12974,N_12997);
nor U13604 (N_13604,N_12762,N_12827);
xor U13605 (N_13605,N_12592,N_12981);
nor U13606 (N_13606,N_12389,N_12598);
nor U13607 (N_13607,N_12509,N_12541);
and U13608 (N_13608,N_12128,N_12938);
nor U13609 (N_13609,N_12615,N_12262);
or U13610 (N_13610,N_12873,N_12189);
nand U13611 (N_13611,N_12578,N_12529);
and U13612 (N_13612,N_12892,N_12549);
or U13613 (N_13613,N_12593,N_12183);
nor U13614 (N_13614,N_12112,N_12527);
nor U13615 (N_13615,N_12555,N_12056);
and U13616 (N_13616,N_12481,N_12609);
nor U13617 (N_13617,N_12449,N_12416);
nor U13618 (N_13618,N_12610,N_12333);
nor U13619 (N_13619,N_12299,N_12707);
and U13620 (N_13620,N_12004,N_12939);
or U13621 (N_13621,N_12330,N_12744);
or U13622 (N_13622,N_12657,N_12512);
xnor U13623 (N_13623,N_12688,N_12617);
xnor U13624 (N_13624,N_12261,N_12281);
xor U13625 (N_13625,N_12542,N_12608);
nor U13626 (N_13626,N_12782,N_12989);
or U13627 (N_13627,N_12497,N_12704);
nand U13628 (N_13628,N_12653,N_12925);
xnor U13629 (N_13629,N_12048,N_12726);
nand U13630 (N_13630,N_12691,N_12180);
nor U13631 (N_13631,N_12105,N_12444);
or U13632 (N_13632,N_12271,N_12899);
and U13633 (N_13633,N_12179,N_12518);
nor U13634 (N_13634,N_12613,N_12366);
xor U13635 (N_13635,N_12051,N_12461);
xor U13636 (N_13636,N_12602,N_12725);
and U13637 (N_13637,N_12186,N_12416);
or U13638 (N_13638,N_12568,N_12514);
xnor U13639 (N_13639,N_12673,N_12991);
xor U13640 (N_13640,N_12634,N_12356);
nor U13641 (N_13641,N_12316,N_12782);
and U13642 (N_13642,N_12152,N_12404);
and U13643 (N_13643,N_12949,N_12739);
xor U13644 (N_13644,N_12243,N_12917);
or U13645 (N_13645,N_12566,N_12561);
nor U13646 (N_13646,N_12473,N_12245);
and U13647 (N_13647,N_12265,N_12031);
nand U13648 (N_13648,N_12032,N_12186);
and U13649 (N_13649,N_12109,N_12909);
nand U13650 (N_13650,N_12490,N_12827);
and U13651 (N_13651,N_12886,N_12419);
and U13652 (N_13652,N_12174,N_12992);
and U13653 (N_13653,N_12851,N_12734);
nand U13654 (N_13654,N_12171,N_12373);
nor U13655 (N_13655,N_12581,N_12906);
or U13656 (N_13656,N_12879,N_12969);
nor U13657 (N_13657,N_12519,N_12640);
nand U13658 (N_13658,N_12708,N_12815);
nor U13659 (N_13659,N_12382,N_12722);
nand U13660 (N_13660,N_12475,N_12093);
or U13661 (N_13661,N_12219,N_12769);
or U13662 (N_13662,N_12005,N_12790);
nand U13663 (N_13663,N_12874,N_12704);
nand U13664 (N_13664,N_12774,N_12717);
xnor U13665 (N_13665,N_12394,N_12189);
xnor U13666 (N_13666,N_12706,N_12870);
or U13667 (N_13667,N_12090,N_12658);
or U13668 (N_13668,N_12640,N_12448);
nor U13669 (N_13669,N_12159,N_12395);
xnor U13670 (N_13670,N_12003,N_12039);
nor U13671 (N_13671,N_12278,N_12552);
and U13672 (N_13672,N_12178,N_12676);
nand U13673 (N_13673,N_12392,N_12568);
or U13674 (N_13674,N_12370,N_12507);
nand U13675 (N_13675,N_12324,N_12962);
and U13676 (N_13676,N_12527,N_12077);
nand U13677 (N_13677,N_12180,N_12495);
nor U13678 (N_13678,N_12415,N_12773);
nand U13679 (N_13679,N_12362,N_12857);
and U13680 (N_13680,N_12991,N_12879);
and U13681 (N_13681,N_12834,N_12517);
nor U13682 (N_13682,N_12225,N_12749);
and U13683 (N_13683,N_12706,N_12052);
nor U13684 (N_13684,N_12667,N_12410);
nand U13685 (N_13685,N_12668,N_12900);
and U13686 (N_13686,N_12551,N_12519);
nor U13687 (N_13687,N_12641,N_12046);
xnor U13688 (N_13688,N_12717,N_12972);
nor U13689 (N_13689,N_12616,N_12791);
nor U13690 (N_13690,N_12416,N_12641);
nor U13691 (N_13691,N_12927,N_12207);
and U13692 (N_13692,N_12677,N_12582);
xor U13693 (N_13693,N_12108,N_12728);
nand U13694 (N_13694,N_12799,N_12113);
nor U13695 (N_13695,N_12572,N_12175);
nor U13696 (N_13696,N_12793,N_12624);
nor U13697 (N_13697,N_12074,N_12925);
and U13698 (N_13698,N_12551,N_12901);
or U13699 (N_13699,N_12761,N_12967);
xnor U13700 (N_13700,N_12743,N_12604);
xnor U13701 (N_13701,N_12993,N_12733);
nand U13702 (N_13702,N_12827,N_12842);
xor U13703 (N_13703,N_12173,N_12060);
nand U13704 (N_13704,N_12828,N_12676);
and U13705 (N_13705,N_12853,N_12996);
nor U13706 (N_13706,N_12926,N_12073);
nand U13707 (N_13707,N_12991,N_12599);
xor U13708 (N_13708,N_12950,N_12902);
nor U13709 (N_13709,N_12268,N_12010);
nor U13710 (N_13710,N_12353,N_12147);
nor U13711 (N_13711,N_12067,N_12021);
or U13712 (N_13712,N_12776,N_12575);
and U13713 (N_13713,N_12390,N_12524);
or U13714 (N_13714,N_12320,N_12293);
or U13715 (N_13715,N_12210,N_12411);
nand U13716 (N_13716,N_12166,N_12800);
nand U13717 (N_13717,N_12368,N_12020);
xor U13718 (N_13718,N_12732,N_12852);
xnor U13719 (N_13719,N_12904,N_12959);
and U13720 (N_13720,N_12220,N_12898);
nand U13721 (N_13721,N_12847,N_12299);
or U13722 (N_13722,N_12635,N_12126);
or U13723 (N_13723,N_12536,N_12052);
or U13724 (N_13724,N_12477,N_12958);
nor U13725 (N_13725,N_12090,N_12967);
or U13726 (N_13726,N_12748,N_12526);
or U13727 (N_13727,N_12023,N_12371);
xnor U13728 (N_13728,N_12549,N_12436);
and U13729 (N_13729,N_12127,N_12718);
nand U13730 (N_13730,N_12181,N_12153);
and U13731 (N_13731,N_12422,N_12750);
xnor U13732 (N_13732,N_12408,N_12761);
nand U13733 (N_13733,N_12994,N_12638);
and U13734 (N_13734,N_12072,N_12804);
or U13735 (N_13735,N_12544,N_12667);
nand U13736 (N_13736,N_12656,N_12326);
xor U13737 (N_13737,N_12012,N_12022);
xor U13738 (N_13738,N_12511,N_12648);
nor U13739 (N_13739,N_12569,N_12458);
or U13740 (N_13740,N_12097,N_12091);
nand U13741 (N_13741,N_12877,N_12899);
xnor U13742 (N_13742,N_12675,N_12516);
xnor U13743 (N_13743,N_12925,N_12353);
and U13744 (N_13744,N_12996,N_12433);
nand U13745 (N_13745,N_12047,N_12674);
and U13746 (N_13746,N_12285,N_12661);
nor U13747 (N_13747,N_12016,N_12665);
nand U13748 (N_13748,N_12022,N_12026);
nor U13749 (N_13749,N_12102,N_12599);
nand U13750 (N_13750,N_12744,N_12775);
or U13751 (N_13751,N_12016,N_12352);
nor U13752 (N_13752,N_12750,N_12090);
xnor U13753 (N_13753,N_12677,N_12514);
xor U13754 (N_13754,N_12296,N_12352);
xor U13755 (N_13755,N_12924,N_12152);
or U13756 (N_13756,N_12839,N_12969);
and U13757 (N_13757,N_12217,N_12933);
and U13758 (N_13758,N_12917,N_12226);
and U13759 (N_13759,N_12942,N_12523);
nor U13760 (N_13760,N_12891,N_12014);
and U13761 (N_13761,N_12314,N_12304);
nand U13762 (N_13762,N_12154,N_12506);
nand U13763 (N_13763,N_12596,N_12681);
and U13764 (N_13764,N_12320,N_12279);
or U13765 (N_13765,N_12350,N_12180);
or U13766 (N_13766,N_12128,N_12035);
and U13767 (N_13767,N_12206,N_12264);
and U13768 (N_13768,N_12081,N_12170);
nand U13769 (N_13769,N_12825,N_12538);
and U13770 (N_13770,N_12380,N_12351);
and U13771 (N_13771,N_12044,N_12321);
or U13772 (N_13772,N_12350,N_12678);
xor U13773 (N_13773,N_12010,N_12008);
and U13774 (N_13774,N_12000,N_12095);
and U13775 (N_13775,N_12423,N_12298);
and U13776 (N_13776,N_12774,N_12378);
nor U13777 (N_13777,N_12261,N_12642);
xor U13778 (N_13778,N_12612,N_12542);
and U13779 (N_13779,N_12236,N_12339);
nor U13780 (N_13780,N_12797,N_12973);
and U13781 (N_13781,N_12597,N_12630);
or U13782 (N_13782,N_12858,N_12667);
nand U13783 (N_13783,N_12957,N_12264);
and U13784 (N_13784,N_12354,N_12869);
and U13785 (N_13785,N_12208,N_12674);
and U13786 (N_13786,N_12048,N_12937);
nand U13787 (N_13787,N_12151,N_12169);
and U13788 (N_13788,N_12368,N_12395);
nor U13789 (N_13789,N_12312,N_12644);
or U13790 (N_13790,N_12334,N_12417);
and U13791 (N_13791,N_12289,N_12437);
and U13792 (N_13792,N_12888,N_12599);
or U13793 (N_13793,N_12930,N_12735);
or U13794 (N_13794,N_12858,N_12311);
or U13795 (N_13795,N_12729,N_12849);
or U13796 (N_13796,N_12862,N_12233);
xor U13797 (N_13797,N_12334,N_12444);
xor U13798 (N_13798,N_12901,N_12366);
xor U13799 (N_13799,N_12773,N_12296);
nor U13800 (N_13800,N_12335,N_12326);
and U13801 (N_13801,N_12306,N_12042);
nor U13802 (N_13802,N_12206,N_12019);
nor U13803 (N_13803,N_12895,N_12521);
nor U13804 (N_13804,N_12161,N_12348);
and U13805 (N_13805,N_12192,N_12024);
and U13806 (N_13806,N_12889,N_12763);
nand U13807 (N_13807,N_12559,N_12012);
or U13808 (N_13808,N_12281,N_12085);
nand U13809 (N_13809,N_12929,N_12335);
nor U13810 (N_13810,N_12641,N_12189);
nor U13811 (N_13811,N_12486,N_12459);
nand U13812 (N_13812,N_12454,N_12740);
nor U13813 (N_13813,N_12998,N_12312);
and U13814 (N_13814,N_12836,N_12531);
xnor U13815 (N_13815,N_12044,N_12916);
and U13816 (N_13816,N_12071,N_12389);
or U13817 (N_13817,N_12282,N_12468);
or U13818 (N_13818,N_12840,N_12563);
nand U13819 (N_13819,N_12502,N_12102);
nand U13820 (N_13820,N_12341,N_12963);
nand U13821 (N_13821,N_12109,N_12048);
and U13822 (N_13822,N_12291,N_12730);
nand U13823 (N_13823,N_12642,N_12365);
nand U13824 (N_13824,N_12534,N_12870);
nand U13825 (N_13825,N_12757,N_12712);
xnor U13826 (N_13826,N_12529,N_12982);
or U13827 (N_13827,N_12317,N_12350);
nor U13828 (N_13828,N_12847,N_12352);
xnor U13829 (N_13829,N_12208,N_12333);
nor U13830 (N_13830,N_12568,N_12705);
xor U13831 (N_13831,N_12784,N_12864);
or U13832 (N_13832,N_12736,N_12908);
xnor U13833 (N_13833,N_12322,N_12826);
nand U13834 (N_13834,N_12869,N_12049);
nor U13835 (N_13835,N_12212,N_12103);
or U13836 (N_13836,N_12533,N_12664);
nor U13837 (N_13837,N_12340,N_12106);
nor U13838 (N_13838,N_12160,N_12784);
and U13839 (N_13839,N_12256,N_12190);
or U13840 (N_13840,N_12283,N_12926);
xnor U13841 (N_13841,N_12433,N_12543);
and U13842 (N_13842,N_12672,N_12912);
nor U13843 (N_13843,N_12657,N_12477);
or U13844 (N_13844,N_12690,N_12802);
xor U13845 (N_13845,N_12296,N_12668);
and U13846 (N_13846,N_12971,N_12609);
xnor U13847 (N_13847,N_12882,N_12286);
or U13848 (N_13848,N_12247,N_12873);
nand U13849 (N_13849,N_12564,N_12450);
nand U13850 (N_13850,N_12649,N_12142);
and U13851 (N_13851,N_12127,N_12035);
nand U13852 (N_13852,N_12731,N_12256);
xor U13853 (N_13853,N_12365,N_12378);
nand U13854 (N_13854,N_12973,N_12930);
xor U13855 (N_13855,N_12272,N_12454);
xnor U13856 (N_13856,N_12649,N_12008);
nand U13857 (N_13857,N_12547,N_12982);
nand U13858 (N_13858,N_12501,N_12055);
and U13859 (N_13859,N_12698,N_12342);
nand U13860 (N_13860,N_12246,N_12286);
and U13861 (N_13861,N_12042,N_12399);
nand U13862 (N_13862,N_12672,N_12777);
xor U13863 (N_13863,N_12334,N_12018);
nand U13864 (N_13864,N_12408,N_12452);
or U13865 (N_13865,N_12057,N_12112);
and U13866 (N_13866,N_12448,N_12036);
xnor U13867 (N_13867,N_12761,N_12629);
or U13868 (N_13868,N_12650,N_12274);
nand U13869 (N_13869,N_12798,N_12196);
and U13870 (N_13870,N_12717,N_12679);
nor U13871 (N_13871,N_12849,N_12456);
nand U13872 (N_13872,N_12958,N_12938);
and U13873 (N_13873,N_12636,N_12717);
nand U13874 (N_13874,N_12845,N_12722);
nor U13875 (N_13875,N_12856,N_12976);
or U13876 (N_13876,N_12718,N_12705);
or U13877 (N_13877,N_12612,N_12732);
or U13878 (N_13878,N_12026,N_12078);
nand U13879 (N_13879,N_12511,N_12783);
and U13880 (N_13880,N_12135,N_12150);
and U13881 (N_13881,N_12281,N_12715);
nand U13882 (N_13882,N_12992,N_12329);
or U13883 (N_13883,N_12063,N_12191);
nor U13884 (N_13884,N_12351,N_12718);
or U13885 (N_13885,N_12543,N_12002);
nand U13886 (N_13886,N_12459,N_12549);
xor U13887 (N_13887,N_12024,N_12049);
and U13888 (N_13888,N_12309,N_12184);
nand U13889 (N_13889,N_12525,N_12944);
nor U13890 (N_13890,N_12063,N_12102);
xor U13891 (N_13891,N_12545,N_12699);
or U13892 (N_13892,N_12741,N_12477);
nor U13893 (N_13893,N_12763,N_12957);
and U13894 (N_13894,N_12579,N_12069);
xnor U13895 (N_13895,N_12909,N_12373);
xnor U13896 (N_13896,N_12180,N_12857);
nand U13897 (N_13897,N_12011,N_12433);
xor U13898 (N_13898,N_12799,N_12198);
or U13899 (N_13899,N_12689,N_12974);
xnor U13900 (N_13900,N_12887,N_12342);
nor U13901 (N_13901,N_12988,N_12328);
or U13902 (N_13902,N_12184,N_12162);
nand U13903 (N_13903,N_12484,N_12821);
or U13904 (N_13904,N_12074,N_12042);
or U13905 (N_13905,N_12979,N_12234);
nor U13906 (N_13906,N_12476,N_12659);
and U13907 (N_13907,N_12809,N_12302);
and U13908 (N_13908,N_12750,N_12879);
or U13909 (N_13909,N_12143,N_12609);
nor U13910 (N_13910,N_12074,N_12082);
nor U13911 (N_13911,N_12930,N_12647);
nand U13912 (N_13912,N_12362,N_12334);
xor U13913 (N_13913,N_12512,N_12958);
xnor U13914 (N_13914,N_12716,N_12570);
and U13915 (N_13915,N_12845,N_12929);
and U13916 (N_13916,N_12188,N_12572);
or U13917 (N_13917,N_12522,N_12523);
and U13918 (N_13918,N_12693,N_12691);
nor U13919 (N_13919,N_12199,N_12478);
and U13920 (N_13920,N_12836,N_12308);
and U13921 (N_13921,N_12491,N_12118);
and U13922 (N_13922,N_12699,N_12554);
nor U13923 (N_13923,N_12277,N_12601);
xor U13924 (N_13924,N_12864,N_12198);
xor U13925 (N_13925,N_12752,N_12793);
xor U13926 (N_13926,N_12608,N_12717);
xnor U13927 (N_13927,N_12738,N_12702);
or U13928 (N_13928,N_12618,N_12769);
xor U13929 (N_13929,N_12993,N_12617);
or U13930 (N_13930,N_12781,N_12400);
nor U13931 (N_13931,N_12703,N_12644);
nor U13932 (N_13932,N_12550,N_12649);
and U13933 (N_13933,N_12505,N_12891);
xor U13934 (N_13934,N_12989,N_12269);
xor U13935 (N_13935,N_12286,N_12111);
or U13936 (N_13936,N_12506,N_12194);
xnor U13937 (N_13937,N_12236,N_12357);
xor U13938 (N_13938,N_12633,N_12497);
nor U13939 (N_13939,N_12807,N_12379);
nor U13940 (N_13940,N_12907,N_12462);
and U13941 (N_13941,N_12382,N_12054);
or U13942 (N_13942,N_12917,N_12265);
nor U13943 (N_13943,N_12985,N_12986);
xor U13944 (N_13944,N_12487,N_12398);
nor U13945 (N_13945,N_12213,N_12184);
and U13946 (N_13946,N_12030,N_12010);
nand U13947 (N_13947,N_12982,N_12132);
or U13948 (N_13948,N_12448,N_12922);
and U13949 (N_13949,N_12827,N_12136);
and U13950 (N_13950,N_12906,N_12078);
xnor U13951 (N_13951,N_12955,N_12446);
or U13952 (N_13952,N_12581,N_12260);
nand U13953 (N_13953,N_12270,N_12252);
or U13954 (N_13954,N_12068,N_12425);
nor U13955 (N_13955,N_12642,N_12959);
nor U13956 (N_13956,N_12166,N_12640);
and U13957 (N_13957,N_12291,N_12600);
xnor U13958 (N_13958,N_12300,N_12182);
nand U13959 (N_13959,N_12047,N_12552);
xor U13960 (N_13960,N_12889,N_12325);
nand U13961 (N_13961,N_12947,N_12249);
nand U13962 (N_13962,N_12512,N_12520);
and U13963 (N_13963,N_12628,N_12572);
and U13964 (N_13964,N_12557,N_12519);
and U13965 (N_13965,N_12384,N_12243);
or U13966 (N_13966,N_12154,N_12565);
nor U13967 (N_13967,N_12234,N_12759);
xor U13968 (N_13968,N_12466,N_12011);
nand U13969 (N_13969,N_12199,N_12732);
nor U13970 (N_13970,N_12817,N_12953);
or U13971 (N_13971,N_12355,N_12306);
xnor U13972 (N_13972,N_12925,N_12765);
nor U13973 (N_13973,N_12795,N_12187);
nand U13974 (N_13974,N_12195,N_12980);
nor U13975 (N_13975,N_12334,N_12491);
nor U13976 (N_13976,N_12197,N_12046);
xor U13977 (N_13977,N_12546,N_12445);
or U13978 (N_13978,N_12738,N_12509);
nand U13979 (N_13979,N_12308,N_12513);
xnor U13980 (N_13980,N_12006,N_12374);
or U13981 (N_13981,N_12818,N_12531);
nand U13982 (N_13982,N_12781,N_12640);
xor U13983 (N_13983,N_12255,N_12782);
xor U13984 (N_13984,N_12380,N_12591);
nand U13985 (N_13985,N_12877,N_12890);
or U13986 (N_13986,N_12938,N_12239);
xnor U13987 (N_13987,N_12101,N_12131);
nand U13988 (N_13988,N_12121,N_12911);
and U13989 (N_13989,N_12755,N_12447);
or U13990 (N_13990,N_12811,N_12477);
nor U13991 (N_13991,N_12814,N_12535);
xor U13992 (N_13992,N_12651,N_12348);
xnor U13993 (N_13993,N_12739,N_12964);
and U13994 (N_13994,N_12249,N_12520);
nor U13995 (N_13995,N_12622,N_12978);
xnor U13996 (N_13996,N_12149,N_12339);
nand U13997 (N_13997,N_12192,N_12528);
or U13998 (N_13998,N_12514,N_12563);
xnor U13999 (N_13999,N_12898,N_12502);
or U14000 (N_14000,N_13700,N_13112);
nand U14001 (N_14001,N_13558,N_13770);
xnor U14002 (N_14002,N_13133,N_13439);
or U14003 (N_14003,N_13247,N_13016);
or U14004 (N_14004,N_13529,N_13861);
xnor U14005 (N_14005,N_13073,N_13410);
or U14006 (N_14006,N_13272,N_13198);
nor U14007 (N_14007,N_13052,N_13603);
nand U14008 (N_14008,N_13682,N_13689);
or U14009 (N_14009,N_13932,N_13291);
or U14010 (N_14010,N_13680,N_13701);
nor U14011 (N_14011,N_13955,N_13222);
nor U14012 (N_14012,N_13438,N_13948);
or U14013 (N_14013,N_13616,N_13165);
or U14014 (N_14014,N_13171,N_13132);
nand U14015 (N_14015,N_13725,N_13578);
and U14016 (N_14016,N_13402,N_13371);
nand U14017 (N_14017,N_13140,N_13684);
or U14018 (N_14018,N_13671,N_13117);
xnor U14019 (N_14019,N_13376,N_13562);
nor U14020 (N_14020,N_13254,N_13460);
xnor U14021 (N_14021,N_13798,N_13512);
nand U14022 (N_14022,N_13323,N_13006);
nor U14023 (N_14023,N_13642,N_13647);
or U14024 (N_14024,N_13366,N_13385);
nand U14025 (N_14025,N_13063,N_13361);
xnor U14026 (N_14026,N_13098,N_13940);
and U14027 (N_14027,N_13625,N_13226);
nand U14028 (N_14028,N_13949,N_13008);
nand U14029 (N_14029,N_13049,N_13885);
and U14030 (N_14030,N_13736,N_13193);
xnor U14031 (N_14031,N_13277,N_13930);
or U14032 (N_14032,N_13836,N_13213);
nand U14033 (N_14033,N_13629,N_13546);
nand U14034 (N_14034,N_13174,N_13741);
nand U14035 (N_14035,N_13234,N_13574);
nor U14036 (N_14036,N_13261,N_13034);
and U14037 (N_14037,N_13168,N_13211);
nor U14038 (N_14038,N_13941,N_13173);
nand U14039 (N_14039,N_13145,N_13243);
nand U14040 (N_14040,N_13424,N_13362);
or U14041 (N_14041,N_13594,N_13199);
or U14042 (N_14042,N_13888,N_13744);
and U14043 (N_14043,N_13271,N_13720);
xor U14044 (N_14044,N_13509,N_13002);
nand U14045 (N_14045,N_13815,N_13242);
nor U14046 (N_14046,N_13550,N_13635);
xor U14047 (N_14047,N_13347,N_13292);
and U14048 (N_14048,N_13055,N_13980);
nor U14049 (N_14049,N_13417,N_13936);
and U14050 (N_14050,N_13917,N_13586);
nor U14051 (N_14051,N_13910,N_13833);
nand U14052 (N_14052,N_13392,N_13022);
and U14053 (N_14053,N_13054,N_13229);
nand U14054 (N_14054,N_13609,N_13928);
xnor U14055 (N_14055,N_13982,N_13020);
nand U14056 (N_14056,N_13709,N_13080);
and U14057 (N_14057,N_13528,N_13040);
nor U14058 (N_14058,N_13494,N_13737);
nor U14059 (N_14059,N_13164,N_13547);
xnor U14060 (N_14060,N_13202,N_13563);
xnor U14061 (N_14061,N_13100,N_13543);
xor U14062 (N_14062,N_13263,N_13752);
and U14063 (N_14063,N_13809,N_13458);
nand U14064 (N_14064,N_13905,N_13381);
and U14065 (N_14065,N_13337,N_13889);
xnor U14066 (N_14066,N_13190,N_13697);
and U14067 (N_14067,N_13095,N_13985);
nand U14068 (N_14068,N_13568,N_13601);
or U14069 (N_14069,N_13026,N_13903);
nor U14070 (N_14070,N_13677,N_13379);
or U14071 (N_14071,N_13688,N_13517);
or U14072 (N_14072,N_13446,N_13459);
and U14073 (N_14073,N_13303,N_13879);
nor U14074 (N_14074,N_13904,N_13351);
nor U14075 (N_14075,N_13967,N_13175);
and U14076 (N_14076,N_13289,N_13778);
or U14077 (N_14077,N_13750,N_13456);
and U14078 (N_14078,N_13056,N_13108);
nor U14079 (N_14079,N_13753,N_13728);
nor U14080 (N_14080,N_13602,N_13825);
or U14081 (N_14081,N_13078,N_13826);
and U14082 (N_14082,N_13397,N_13530);
and U14083 (N_14083,N_13152,N_13768);
nand U14084 (N_14084,N_13411,N_13294);
nor U14085 (N_14085,N_13676,N_13617);
nor U14086 (N_14086,N_13404,N_13577);
nor U14087 (N_14087,N_13669,N_13201);
nor U14088 (N_14088,N_13626,N_13837);
xnor U14089 (N_14089,N_13564,N_13510);
or U14090 (N_14090,N_13071,N_13760);
or U14091 (N_14091,N_13899,N_13307);
nor U14092 (N_14092,N_13114,N_13604);
nand U14093 (N_14093,N_13575,N_13331);
nor U14094 (N_14094,N_13349,N_13862);
nor U14095 (N_14095,N_13824,N_13285);
nor U14096 (N_14096,N_13644,N_13342);
or U14097 (N_14097,N_13161,N_13495);
and U14098 (N_14098,N_13631,N_13805);
nand U14099 (N_14099,N_13085,N_13516);
xnor U14100 (N_14100,N_13138,N_13110);
nand U14101 (N_14101,N_13645,N_13525);
nand U14102 (N_14102,N_13148,N_13027);
or U14103 (N_14103,N_13396,N_13665);
nor U14104 (N_14104,N_13388,N_13829);
nand U14105 (N_14105,N_13075,N_13533);
nand U14106 (N_14106,N_13441,N_13074);
and U14107 (N_14107,N_13999,N_13156);
nor U14108 (N_14108,N_13311,N_13442);
or U14109 (N_14109,N_13194,N_13527);
nor U14110 (N_14110,N_13365,N_13325);
xor U14111 (N_14111,N_13238,N_13790);
nor U14112 (N_14112,N_13421,N_13913);
or U14113 (N_14113,N_13419,N_13327);
and U14114 (N_14114,N_13092,N_13561);
and U14115 (N_14115,N_13178,N_13176);
xnor U14116 (N_14116,N_13687,N_13210);
nand U14117 (N_14117,N_13158,N_13852);
xor U14118 (N_14118,N_13989,N_13184);
or U14119 (N_14119,N_13032,N_13641);
and U14120 (N_14120,N_13759,N_13692);
xnor U14121 (N_14121,N_13393,N_13583);
xor U14122 (N_14122,N_13659,N_13183);
xor U14123 (N_14123,N_13290,N_13960);
nor U14124 (N_14124,N_13192,N_13990);
nand U14125 (N_14125,N_13849,N_13037);
or U14126 (N_14126,N_13299,N_13070);
nand U14127 (N_14127,N_13490,N_13857);
nor U14128 (N_14128,N_13549,N_13358);
or U14129 (N_14129,N_13363,N_13621);
and U14130 (N_14130,N_13186,N_13881);
nand U14131 (N_14131,N_13934,N_13783);
or U14132 (N_14132,N_13036,N_13988);
xor U14133 (N_14133,N_13129,N_13666);
xnor U14134 (N_14134,N_13422,N_13735);
or U14135 (N_14135,N_13104,N_13703);
and U14136 (N_14136,N_13639,N_13251);
and U14137 (N_14137,N_13506,N_13432);
and U14138 (N_14138,N_13801,N_13762);
xnor U14139 (N_14139,N_13970,N_13172);
nand U14140 (N_14140,N_13592,N_13423);
nand U14141 (N_14141,N_13465,N_13144);
xnor U14142 (N_14142,N_13330,N_13137);
nand U14143 (N_14143,N_13806,N_13281);
xor U14144 (N_14144,N_13360,N_13312);
xor U14145 (N_14145,N_13004,N_13792);
xnor U14146 (N_14146,N_13452,N_13570);
and U14147 (N_14147,N_13695,N_13011);
nand U14148 (N_14148,N_13386,N_13814);
and U14149 (N_14149,N_13819,N_13914);
nand U14150 (N_14150,N_13035,N_13526);
and U14151 (N_14151,N_13891,N_13590);
or U14152 (N_14152,N_13916,N_13122);
and U14153 (N_14153,N_13265,N_13038);
or U14154 (N_14154,N_13429,N_13010);
or U14155 (N_14155,N_13364,N_13808);
and U14156 (N_14156,N_13420,N_13799);
nor U14157 (N_14157,N_13922,N_13043);
and U14158 (N_14158,N_13179,N_13116);
nand U14159 (N_14159,N_13953,N_13355);
and U14160 (N_14160,N_13968,N_13180);
xnor U14161 (N_14161,N_13064,N_13042);
or U14162 (N_14162,N_13650,N_13557);
xor U14163 (N_14163,N_13431,N_13217);
nor U14164 (N_14164,N_13683,N_13607);
nand U14165 (N_14165,N_13821,N_13001);
xnor U14166 (N_14166,N_13727,N_13489);
xor U14167 (N_14167,N_13542,N_13295);
xor U14168 (N_14168,N_13636,N_13375);
or U14169 (N_14169,N_13784,N_13227);
xnor U14170 (N_14170,N_13651,N_13538);
nand U14171 (N_14171,N_13069,N_13264);
xnor U14172 (N_14172,N_13951,N_13482);
and U14173 (N_14173,N_13785,N_13216);
and U14174 (N_14174,N_13139,N_13864);
nor U14175 (N_14175,N_13492,N_13103);
nor U14176 (N_14176,N_13499,N_13167);
nor U14177 (N_14177,N_13304,N_13196);
nor U14178 (N_14178,N_13153,N_13126);
xnor U14179 (N_14179,N_13445,N_13933);
or U14180 (N_14180,N_13209,N_13044);
and U14181 (N_14181,N_13915,N_13339);
nand U14182 (N_14182,N_13028,N_13079);
xnor U14183 (N_14183,N_13537,N_13923);
and U14184 (N_14184,N_13845,N_13493);
xnor U14185 (N_14185,N_13867,N_13003);
nand U14186 (N_14186,N_13444,N_13455);
nor U14187 (N_14187,N_13344,N_13434);
and U14188 (N_14188,N_13812,N_13518);
or U14189 (N_14189,N_13280,N_13698);
nand U14190 (N_14190,N_13128,N_13314);
nor U14191 (N_14191,N_13977,N_13605);
nor U14192 (N_14192,N_13566,N_13478);
xor U14193 (N_14193,N_13508,N_13062);
nand U14194 (N_14194,N_13552,N_13912);
xor U14195 (N_14195,N_13719,N_13502);
or U14196 (N_14196,N_13253,N_13433);
nor U14197 (N_14197,N_13597,N_13739);
nor U14198 (N_14198,N_13320,N_13598);
nand U14199 (N_14199,N_13863,N_13302);
and U14200 (N_14200,N_13974,N_13279);
nand U14201 (N_14201,N_13992,N_13149);
nand U14202 (N_14202,N_13556,N_13484);
or U14203 (N_14203,N_13769,N_13795);
nand U14204 (N_14204,N_13130,N_13803);
and U14205 (N_14205,N_13485,N_13147);
xor U14206 (N_14206,N_13013,N_13997);
nand U14207 (N_14207,N_13157,N_13730);
and U14208 (N_14208,N_13704,N_13944);
nor U14209 (N_14209,N_13163,N_13487);
xnor U14210 (N_14210,N_13774,N_13865);
and U14211 (N_14211,N_13731,N_13582);
and U14212 (N_14212,N_13966,N_13531);
xnor U14213 (N_14213,N_13426,N_13077);
and U14214 (N_14214,N_13443,N_13696);
nand U14215 (N_14215,N_13775,N_13749);
or U14216 (N_14216,N_13593,N_13800);
nand U14217 (N_14217,N_13875,N_13614);
xor U14218 (N_14218,N_13779,N_13699);
or U14219 (N_14219,N_13535,N_13816);
nand U14220 (N_14220,N_13995,N_13324);
nand U14221 (N_14221,N_13082,N_13335);
xor U14222 (N_14222,N_13757,N_13322);
nor U14223 (N_14223,N_13898,N_13882);
and U14224 (N_14224,N_13802,N_13634);
xnor U14225 (N_14225,N_13878,N_13576);
or U14226 (N_14226,N_13747,N_13571);
nand U14227 (N_14227,N_13789,N_13370);
xnor U14228 (N_14228,N_13893,N_13346);
nand U14229 (N_14229,N_13019,N_13679);
and U14230 (N_14230,N_13522,N_13232);
or U14231 (N_14231,N_13150,N_13024);
and U14232 (N_14232,N_13476,N_13464);
nand U14233 (N_14233,N_13722,N_13657);
or U14234 (N_14234,N_13600,N_13200);
and U14235 (N_14235,N_13328,N_13931);
nor U14236 (N_14236,N_13670,N_13258);
nor U14237 (N_14237,N_13207,N_13113);
nand U14238 (N_14238,N_13500,N_13610);
and U14239 (N_14239,N_13479,N_13664);
nor U14240 (N_14240,N_13937,N_13154);
nor U14241 (N_14241,N_13050,N_13230);
nand U14242 (N_14242,N_13978,N_13548);
or U14243 (N_14243,N_13579,N_13282);
nor U14244 (N_14244,N_13950,N_13545);
xnor U14245 (N_14245,N_13662,N_13830);
xnor U14246 (N_14246,N_13214,N_13694);
or U14247 (N_14247,N_13846,N_13096);
and U14248 (N_14248,N_13613,N_13276);
and U14249 (N_14249,N_13619,N_13461);
xor U14250 (N_14250,N_13565,N_13345);
or U14251 (N_14251,N_13855,N_13884);
nor U14252 (N_14252,N_13283,N_13266);
nor U14253 (N_14253,N_13847,N_13319);
and U14254 (N_14254,N_13856,N_13733);
and U14255 (N_14255,N_13394,N_13854);
xnor U14256 (N_14256,N_13298,N_13972);
nand U14257 (N_14257,N_13109,N_13555);
and U14258 (N_14258,N_13668,N_13707);
or U14259 (N_14259,N_13356,N_13716);
and U14260 (N_14260,N_13726,N_13656);
xnor U14261 (N_14261,N_13943,N_13804);
xnor U14262 (N_14262,N_13851,N_13581);
and U14263 (N_14263,N_13615,N_13191);
nand U14264 (N_14264,N_13329,N_13678);
xnor U14265 (N_14265,N_13909,N_13823);
or U14266 (N_14266,N_13467,N_13497);
or U14267 (N_14267,N_13275,N_13880);
and U14268 (N_14268,N_13751,N_13900);
xor U14269 (N_14269,N_13136,N_13208);
nand U14270 (N_14270,N_13127,N_13892);
or U14271 (N_14271,N_13296,N_13724);
nor U14272 (N_14272,N_13952,N_13890);
nand U14273 (N_14273,N_13119,N_13352);
nor U14274 (N_14274,N_13667,N_13300);
or U14275 (N_14275,N_13973,N_13297);
nor U14276 (N_14276,N_13195,N_13551);
xnor U14277 (N_14277,N_13633,N_13541);
nor U14278 (N_14278,N_13712,N_13767);
nor U14279 (N_14279,N_13734,N_13118);
nor U14280 (N_14280,N_13181,N_13067);
nor U14281 (N_14281,N_13732,N_13742);
nor U14282 (N_14282,N_13975,N_13378);
xor U14283 (N_14283,N_13462,N_13929);
and U14284 (N_14284,N_13486,N_13206);
nand U14285 (N_14285,N_13348,N_13691);
or U14286 (N_14286,N_13764,N_13853);
and U14287 (N_14287,N_13637,N_13964);
and U14288 (N_14288,N_13418,N_13483);
and U14289 (N_14289,N_13448,N_13959);
nand U14290 (N_14290,N_13313,N_13146);
nand U14291 (N_14291,N_13938,N_13763);
nor U14292 (N_14292,N_13817,N_13134);
or U14293 (N_14293,N_13559,N_13661);
and U14294 (N_14294,N_13231,N_13969);
or U14295 (N_14295,N_13869,N_13796);
nor U14296 (N_14296,N_13873,N_13256);
or U14297 (N_14297,N_13205,N_13447);
nand U14298 (N_14298,N_13850,N_13954);
nor U14299 (N_14299,N_13084,N_13189);
nand U14300 (N_14300,N_13389,N_13906);
and U14301 (N_14301,N_13491,N_13620);
or U14302 (N_14302,N_13534,N_13408);
nor U14303 (N_14303,N_13239,N_13368);
nand U14304 (N_14304,N_13791,N_13235);
and U14305 (N_14305,N_13017,N_13984);
xnor U14306 (N_14306,N_13539,N_13336);
or U14307 (N_14307,N_13811,N_13093);
nand U14308 (N_14308,N_13761,N_13310);
nand U14309 (N_14309,N_13515,N_13588);
and U14310 (N_14310,N_13781,N_13965);
or U14311 (N_14311,N_13987,N_13745);
nand U14312 (N_14312,N_13723,N_13437);
nand U14313 (N_14313,N_13470,N_13454);
xnor U14314 (N_14314,N_13640,N_13685);
nor U14315 (N_14315,N_13939,N_13106);
and U14316 (N_14316,N_13244,N_13436);
and U14317 (N_14317,N_13513,N_13755);
nor U14318 (N_14318,N_13204,N_13057);
and U14319 (N_14319,N_13942,N_13794);
nor U14320 (N_14320,N_13252,N_13115);
nand U14321 (N_14321,N_13041,N_13007);
or U14322 (N_14322,N_13409,N_13618);
nor U14323 (N_14323,N_13776,N_13608);
xor U14324 (N_14324,N_13628,N_13377);
xnor U14325 (N_14325,N_13160,N_13868);
xor U14326 (N_14326,N_13961,N_13390);
and U14327 (N_14327,N_13591,N_13046);
nor U14328 (N_14328,N_13714,N_13463);
and U14329 (N_14329,N_13838,N_13693);
nand U14330 (N_14330,N_13068,N_13511);
nor U14331 (N_14331,N_13935,N_13589);
or U14332 (N_14332,N_13507,N_13469);
or U14333 (N_14333,N_13842,N_13877);
nor U14334 (N_14334,N_13874,N_13627);
xnor U14335 (N_14335,N_13983,N_13993);
or U14336 (N_14336,N_13729,N_13269);
nor U14337 (N_14337,N_13083,N_13748);
nand U14338 (N_14338,N_13267,N_13706);
and U14339 (N_14339,N_13876,N_13758);
nor U14340 (N_14340,N_13369,N_13690);
or U14341 (N_14341,N_13412,N_13717);
and U14342 (N_14342,N_13498,N_13273);
or U14343 (N_14343,N_13503,N_13756);
nand U14344 (N_14344,N_13318,N_13653);
nor U14345 (N_14345,N_13123,N_13274);
and U14346 (N_14346,N_13257,N_13284);
nand U14347 (N_14347,N_13249,N_13713);
or U14348 (N_14348,N_13357,N_13124);
or U14349 (N_14349,N_13143,N_13612);
xor U14350 (N_14350,N_13520,N_13449);
nor U14351 (N_14351,N_13228,N_13976);
nor U14352 (N_14352,N_13766,N_13341);
or U14353 (N_14353,N_13772,N_13262);
and U14354 (N_14354,N_13840,N_13648);
nand U14355 (N_14355,N_13587,N_13185);
nor U14356 (N_14356,N_13260,N_13524);
and U14357 (N_14357,N_13957,N_13025);
and U14358 (N_14358,N_13309,N_13606);
xnor U14359 (N_14359,N_13946,N_13278);
nor U14360 (N_14360,N_13215,N_13250);
nand U14361 (N_14361,N_13481,N_13643);
and U14362 (N_14362,N_13415,N_13746);
nor U14363 (N_14363,N_13673,N_13018);
or U14364 (N_14364,N_13771,N_13780);
or U14365 (N_14365,N_13155,N_13197);
xnor U14366 (N_14366,N_13848,N_13872);
or U14367 (N_14367,N_13918,N_13947);
or U14368 (N_14368,N_13945,N_13121);
nor U14369 (N_14369,N_13921,N_13457);
nand U14370 (N_14370,N_13340,N_13622);
and U14371 (N_14371,N_13416,N_13708);
nor U14372 (N_14372,N_13089,N_13962);
xor U14373 (N_14373,N_13956,N_13996);
nor U14374 (N_14374,N_13523,N_13859);
xnor U14375 (N_14375,N_13400,N_13111);
xnor U14376 (N_14376,N_13675,N_13187);
nor U14377 (N_14377,N_13182,N_13505);
or U14378 (N_14378,N_13886,N_13797);
nand U14379 (N_14379,N_13480,N_13086);
nor U14380 (N_14380,N_13632,N_13532);
or U14381 (N_14381,N_13553,N_13177);
and U14382 (N_14382,N_13401,N_13718);
and U14383 (N_14383,N_13354,N_13536);
xor U14384 (N_14384,N_13087,N_13504);
nor U14385 (N_14385,N_13924,N_13000);
nand U14386 (N_14386,N_13715,N_13223);
nor U14387 (N_14387,N_13301,N_13573);
nor U14388 (N_14388,N_13427,N_13501);
or U14389 (N_14389,N_13286,N_13896);
xnor U14390 (N_14390,N_13475,N_13827);
and U14391 (N_14391,N_13496,N_13142);
xor U14392 (N_14392,N_13107,N_13958);
xnor U14393 (N_14393,N_13765,N_13488);
nand U14394 (N_14394,N_13151,N_13188);
or U14395 (N_14395,N_13674,N_13981);
nor U14396 (N_14396,N_13374,N_13843);
and U14397 (N_14397,N_13754,N_13926);
xnor U14398 (N_14398,N_13560,N_13860);
nand U14399 (N_14399,N_13646,N_13908);
nand U14400 (N_14400,N_13813,N_13822);
and U14401 (N_14401,N_13514,N_13031);
and U14402 (N_14402,N_13450,N_13088);
nand U14403 (N_14403,N_13051,N_13061);
xnor U14404 (N_14404,N_13245,N_13711);
or U14405 (N_14405,N_13787,N_13986);
xnor U14406 (N_14406,N_13584,N_13477);
nor U14407 (N_14407,N_13435,N_13065);
nand U14408 (N_14408,N_13248,N_13383);
xnor U14409 (N_14409,N_13023,N_13072);
xor U14410 (N_14410,N_13220,N_13246);
and U14411 (N_14411,N_13911,N_13094);
nand U14412 (N_14412,N_13858,N_13554);
and U14413 (N_14413,N_13326,N_13241);
or U14414 (N_14414,N_13332,N_13162);
nor U14415 (N_14415,N_13818,N_13721);
and U14416 (N_14416,N_13793,N_13039);
and U14417 (N_14417,N_13569,N_13540);
or U14418 (N_14418,N_13472,N_13414);
nor U14419 (N_14419,N_13466,N_13403);
xor U14420 (N_14420,N_13630,N_13212);
nand U14421 (N_14421,N_13810,N_13090);
nand U14422 (N_14422,N_13407,N_13372);
xor U14423 (N_14423,N_13471,N_13773);
and U14424 (N_14424,N_13743,N_13315);
nor U14425 (N_14425,N_13474,N_13097);
xor U14426 (N_14426,N_13473,N_13963);
nand U14427 (N_14427,N_13658,N_13270);
nor U14428 (N_14428,N_13870,N_13014);
nand U14429 (N_14429,N_13125,N_13373);
or U14430 (N_14430,N_13353,N_13045);
xor U14431 (N_14431,N_13159,N_13901);
nor U14432 (N_14432,N_13091,N_13521);
nand U14433 (N_14433,N_13585,N_13135);
nor U14434 (N_14434,N_13702,N_13406);
and U14435 (N_14435,N_13705,N_13306);
xnor U14436 (N_14436,N_13048,N_13897);
nor U14437 (N_14437,N_13623,N_13219);
nor U14438 (N_14438,N_13820,N_13102);
or U14439 (N_14439,N_13287,N_13203);
nand U14440 (N_14440,N_13076,N_13686);
xnor U14441 (N_14441,N_13887,N_13580);
nor U14442 (N_14442,N_13994,N_13567);
or U14443 (N_14443,N_13468,N_13652);
or U14444 (N_14444,N_13308,N_13255);
nand U14445 (N_14445,N_13105,N_13059);
nand U14446 (N_14446,N_13920,N_13405);
nand U14447 (N_14447,N_13807,N_13738);
nor U14448 (N_14448,N_13380,N_13399);
or U14449 (N_14449,N_13572,N_13894);
and U14450 (N_14450,N_13828,N_13015);
nor U14451 (N_14451,N_13991,N_13060);
nand U14452 (N_14452,N_13288,N_13866);
nand U14453 (N_14453,N_13343,N_13233);
nor U14454 (N_14454,N_13971,N_13544);
nand U14455 (N_14455,N_13321,N_13871);
or U14456 (N_14456,N_13218,N_13047);
and U14457 (N_14457,N_13009,N_13638);
nand U14458 (N_14458,N_13259,N_13021);
and U14459 (N_14459,N_13236,N_13654);
or U14460 (N_14460,N_13305,N_13120);
xnor U14461 (N_14461,N_13831,N_13788);
nor U14462 (N_14462,N_13649,N_13005);
nand U14463 (N_14463,N_13367,N_13012);
xnor U14464 (N_14464,N_13066,N_13169);
xnor U14465 (N_14465,N_13835,N_13334);
and U14466 (N_14466,N_13053,N_13663);
nor U14467 (N_14467,N_13237,N_13672);
nand U14468 (N_14468,N_13919,N_13029);
and U14469 (N_14469,N_13841,N_13710);
and U14470 (N_14470,N_13240,N_13333);
xnor U14471 (N_14471,N_13786,N_13681);
xnor U14472 (N_14472,N_13316,N_13225);
xor U14473 (N_14473,N_13268,N_13081);
and U14474 (N_14474,N_13998,N_13033);
or U14475 (N_14475,N_13660,N_13611);
nor U14476 (N_14476,N_13839,N_13782);
or U14477 (N_14477,N_13141,N_13131);
xor U14478 (N_14478,N_13387,N_13883);
nand U14479 (N_14479,N_13451,N_13391);
or U14480 (N_14480,N_13359,N_13979);
or U14481 (N_14481,N_13338,N_13101);
or U14482 (N_14482,N_13596,N_13430);
and U14483 (N_14483,N_13834,N_13398);
nand U14484 (N_14484,N_13832,N_13224);
xnor U14485 (N_14485,N_13395,N_13293);
xor U14486 (N_14486,N_13382,N_13740);
nor U14487 (N_14487,N_13907,N_13902);
and U14488 (N_14488,N_13599,N_13413);
or U14489 (N_14489,N_13927,N_13519);
or U14490 (N_14490,N_13624,N_13777);
and U14491 (N_14491,N_13170,N_13166);
xor U14492 (N_14492,N_13595,N_13317);
nand U14493 (N_14493,N_13453,N_13428);
nor U14494 (N_14494,N_13384,N_13440);
or U14495 (N_14495,N_13925,N_13221);
nor U14496 (N_14496,N_13844,N_13099);
xnor U14497 (N_14497,N_13425,N_13655);
xnor U14498 (N_14498,N_13030,N_13895);
and U14499 (N_14499,N_13058,N_13350);
xnor U14500 (N_14500,N_13664,N_13432);
and U14501 (N_14501,N_13387,N_13785);
or U14502 (N_14502,N_13245,N_13976);
and U14503 (N_14503,N_13146,N_13750);
or U14504 (N_14504,N_13748,N_13901);
nand U14505 (N_14505,N_13621,N_13058);
nand U14506 (N_14506,N_13568,N_13979);
nand U14507 (N_14507,N_13442,N_13097);
or U14508 (N_14508,N_13238,N_13815);
nand U14509 (N_14509,N_13884,N_13106);
xor U14510 (N_14510,N_13247,N_13335);
xor U14511 (N_14511,N_13523,N_13790);
nor U14512 (N_14512,N_13063,N_13652);
xnor U14513 (N_14513,N_13187,N_13377);
and U14514 (N_14514,N_13087,N_13131);
nor U14515 (N_14515,N_13479,N_13965);
and U14516 (N_14516,N_13179,N_13306);
nand U14517 (N_14517,N_13173,N_13032);
nand U14518 (N_14518,N_13203,N_13396);
or U14519 (N_14519,N_13820,N_13286);
or U14520 (N_14520,N_13635,N_13058);
nand U14521 (N_14521,N_13999,N_13388);
xor U14522 (N_14522,N_13760,N_13797);
and U14523 (N_14523,N_13739,N_13544);
or U14524 (N_14524,N_13487,N_13258);
or U14525 (N_14525,N_13145,N_13741);
nand U14526 (N_14526,N_13708,N_13182);
nand U14527 (N_14527,N_13412,N_13470);
nand U14528 (N_14528,N_13774,N_13684);
or U14529 (N_14529,N_13742,N_13891);
nor U14530 (N_14530,N_13644,N_13782);
nor U14531 (N_14531,N_13669,N_13694);
or U14532 (N_14532,N_13321,N_13012);
nor U14533 (N_14533,N_13440,N_13762);
nand U14534 (N_14534,N_13762,N_13121);
nand U14535 (N_14535,N_13624,N_13394);
nand U14536 (N_14536,N_13236,N_13083);
and U14537 (N_14537,N_13280,N_13978);
xor U14538 (N_14538,N_13544,N_13987);
and U14539 (N_14539,N_13749,N_13576);
xor U14540 (N_14540,N_13605,N_13951);
or U14541 (N_14541,N_13111,N_13041);
nor U14542 (N_14542,N_13611,N_13436);
and U14543 (N_14543,N_13449,N_13685);
and U14544 (N_14544,N_13107,N_13979);
and U14545 (N_14545,N_13600,N_13380);
and U14546 (N_14546,N_13075,N_13435);
or U14547 (N_14547,N_13394,N_13519);
nand U14548 (N_14548,N_13926,N_13078);
nand U14549 (N_14549,N_13196,N_13451);
nor U14550 (N_14550,N_13586,N_13894);
or U14551 (N_14551,N_13469,N_13836);
and U14552 (N_14552,N_13295,N_13164);
nor U14553 (N_14553,N_13565,N_13939);
nand U14554 (N_14554,N_13734,N_13566);
nand U14555 (N_14555,N_13300,N_13855);
nor U14556 (N_14556,N_13352,N_13764);
or U14557 (N_14557,N_13771,N_13525);
and U14558 (N_14558,N_13901,N_13655);
nand U14559 (N_14559,N_13356,N_13577);
or U14560 (N_14560,N_13619,N_13928);
nand U14561 (N_14561,N_13071,N_13647);
and U14562 (N_14562,N_13335,N_13938);
nor U14563 (N_14563,N_13482,N_13333);
nand U14564 (N_14564,N_13865,N_13172);
nand U14565 (N_14565,N_13330,N_13036);
nand U14566 (N_14566,N_13344,N_13851);
and U14567 (N_14567,N_13287,N_13942);
xor U14568 (N_14568,N_13632,N_13406);
and U14569 (N_14569,N_13546,N_13784);
nand U14570 (N_14570,N_13438,N_13248);
and U14571 (N_14571,N_13516,N_13989);
nand U14572 (N_14572,N_13161,N_13609);
or U14573 (N_14573,N_13297,N_13593);
nor U14574 (N_14574,N_13379,N_13628);
nand U14575 (N_14575,N_13799,N_13227);
nor U14576 (N_14576,N_13293,N_13004);
and U14577 (N_14577,N_13179,N_13332);
xor U14578 (N_14578,N_13216,N_13204);
nor U14579 (N_14579,N_13714,N_13198);
nor U14580 (N_14580,N_13144,N_13471);
or U14581 (N_14581,N_13002,N_13700);
and U14582 (N_14582,N_13581,N_13983);
nor U14583 (N_14583,N_13803,N_13358);
nor U14584 (N_14584,N_13470,N_13512);
nand U14585 (N_14585,N_13351,N_13300);
xor U14586 (N_14586,N_13828,N_13349);
nor U14587 (N_14587,N_13209,N_13728);
or U14588 (N_14588,N_13555,N_13115);
and U14589 (N_14589,N_13515,N_13602);
nand U14590 (N_14590,N_13474,N_13901);
nor U14591 (N_14591,N_13446,N_13835);
and U14592 (N_14592,N_13101,N_13311);
nor U14593 (N_14593,N_13490,N_13335);
xnor U14594 (N_14594,N_13951,N_13905);
xnor U14595 (N_14595,N_13882,N_13112);
or U14596 (N_14596,N_13495,N_13301);
xnor U14597 (N_14597,N_13948,N_13898);
xnor U14598 (N_14598,N_13798,N_13421);
nor U14599 (N_14599,N_13083,N_13736);
nand U14600 (N_14600,N_13509,N_13890);
and U14601 (N_14601,N_13433,N_13423);
xnor U14602 (N_14602,N_13891,N_13799);
nand U14603 (N_14603,N_13500,N_13276);
nand U14604 (N_14604,N_13297,N_13073);
or U14605 (N_14605,N_13405,N_13798);
nor U14606 (N_14606,N_13434,N_13512);
or U14607 (N_14607,N_13974,N_13847);
xor U14608 (N_14608,N_13718,N_13961);
xnor U14609 (N_14609,N_13199,N_13566);
and U14610 (N_14610,N_13523,N_13688);
or U14611 (N_14611,N_13309,N_13787);
or U14612 (N_14612,N_13400,N_13645);
nor U14613 (N_14613,N_13705,N_13564);
nor U14614 (N_14614,N_13975,N_13060);
and U14615 (N_14615,N_13842,N_13782);
nor U14616 (N_14616,N_13215,N_13908);
or U14617 (N_14617,N_13608,N_13768);
nor U14618 (N_14618,N_13736,N_13085);
and U14619 (N_14619,N_13101,N_13728);
nor U14620 (N_14620,N_13565,N_13722);
and U14621 (N_14621,N_13378,N_13569);
or U14622 (N_14622,N_13150,N_13772);
nand U14623 (N_14623,N_13617,N_13863);
nand U14624 (N_14624,N_13453,N_13841);
nand U14625 (N_14625,N_13309,N_13462);
nand U14626 (N_14626,N_13987,N_13033);
or U14627 (N_14627,N_13947,N_13014);
nand U14628 (N_14628,N_13641,N_13225);
nand U14629 (N_14629,N_13547,N_13630);
nor U14630 (N_14630,N_13109,N_13644);
nor U14631 (N_14631,N_13682,N_13747);
and U14632 (N_14632,N_13409,N_13628);
and U14633 (N_14633,N_13412,N_13908);
nor U14634 (N_14634,N_13873,N_13527);
nor U14635 (N_14635,N_13246,N_13422);
and U14636 (N_14636,N_13940,N_13515);
and U14637 (N_14637,N_13684,N_13604);
nor U14638 (N_14638,N_13504,N_13010);
xor U14639 (N_14639,N_13082,N_13962);
nand U14640 (N_14640,N_13369,N_13802);
xor U14641 (N_14641,N_13068,N_13512);
nand U14642 (N_14642,N_13685,N_13056);
or U14643 (N_14643,N_13947,N_13098);
and U14644 (N_14644,N_13689,N_13886);
and U14645 (N_14645,N_13801,N_13667);
xnor U14646 (N_14646,N_13930,N_13897);
and U14647 (N_14647,N_13281,N_13666);
xor U14648 (N_14648,N_13942,N_13606);
and U14649 (N_14649,N_13062,N_13652);
xor U14650 (N_14650,N_13841,N_13725);
xor U14651 (N_14651,N_13757,N_13635);
or U14652 (N_14652,N_13842,N_13241);
or U14653 (N_14653,N_13650,N_13604);
nor U14654 (N_14654,N_13203,N_13636);
nand U14655 (N_14655,N_13562,N_13982);
xnor U14656 (N_14656,N_13626,N_13436);
nand U14657 (N_14657,N_13092,N_13693);
nor U14658 (N_14658,N_13824,N_13632);
nand U14659 (N_14659,N_13179,N_13866);
nand U14660 (N_14660,N_13072,N_13120);
and U14661 (N_14661,N_13120,N_13838);
xnor U14662 (N_14662,N_13899,N_13500);
and U14663 (N_14663,N_13940,N_13599);
xnor U14664 (N_14664,N_13205,N_13711);
xor U14665 (N_14665,N_13240,N_13320);
xor U14666 (N_14666,N_13344,N_13027);
or U14667 (N_14667,N_13609,N_13573);
or U14668 (N_14668,N_13798,N_13126);
or U14669 (N_14669,N_13972,N_13498);
or U14670 (N_14670,N_13278,N_13976);
nand U14671 (N_14671,N_13589,N_13568);
and U14672 (N_14672,N_13614,N_13236);
xor U14673 (N_14673,N_13247,N_13356);
or U14674 (N_14674,N_13973,N_13866);
xor U14675 (N_14675,N_13988,N_13985);
nor U14676 (N_14676,N_13830,N_13156);
xor U14677 (N_14677,N_13512,N_13404);
and U14678 (N_14678,N_13424,N_13911);
nor U14679 (N_14679,N_13710,N_13422);
and U14680 (N_14680,N_13204,N_13809);
xnor U14681 (N_14681,N_13387,N_13255);
nand U14682 (N_14682,N_13845,N_13639);
xnor U14683 (N_14683,N_13250,N_13980);
nor U14684 (N_14684,N_13414,N_13152);
and U14685 (N_14685,N_13395,N_13157);
nor U14686 (N_14686,N_13679,N_13075);
or U14687 (N_14687,N_13911,N_13489);
and U14688 (N_14688,N_13778,N_13689);
xor U14689 (N_14689,N_13897,N_13506);
or U14690 (N_14690,N_13238,N_13176);
or U14691 (N_14691,N_13062,N_13626);
nor U14692 (N_14692,N_13495,N_13878);
or U14693 (N_14693,N_13824,N_13212);
and U14694 (N_14694,N_13091,N_13962);
nand U14695 (N_14695,N_13206,N_13741);
or U14696 (N_14696,N_13108,N_13168);
nand U14697 (N_14697,N_13264,N_13734);
nor U14698 (N_14698,N_13090,N_13742);
nor U14699 (N_14699,N_13434,N_13115);
xor U14700 (N_14700,N_13388,N_13816);
nand U14701 (N_14701,N_13322,N_13959);
nand U14702 (N_14702,N_13499,N_13555);
nand U14703 (N_14703,N_13455,N_13253);
or U14704 (N_14704,N_13347,N_13980);
xnor U14705 (N_14705,N_13001,N_13236);
nand U14706 (N_14706,N_13806,N_13950);
xnor U14707 (N_14707,N_13577,N_13664);
nand U14708 (N_14708,N_13562,N_13439);
nor U14709 (N_14709,N_13109,N_13220);
or U14710 (N_14710,N_13427,N_13198);
xor U14711 (N_14711,N_13323,N_13531);
and U14712 (N_14712,N_13859,N_13773);
nor U14713 (N_14713,N_13294,N_13899);
xnor U14714 (N_14714,N_13689,N_13224);
xnor U14715 (N_14715,N_13419,N_13017);
and U14716 (N_14716,N_13516,N_13035);
nor U14717 (N_14717,N_13678,N_13502);
xnor U14718 (N_14718,N_13604,N_13265);
xnor U14719 (N_14719,N_13565,N_13424);
xnor U14720 (N_14720,N_13413,N_13188);
xnor U14721 (N_14721,N_13620,N_13737);
nor U14722 (N_14722,N_13798,N_13325);
and U14723 (N_14723,N_13304,N_13980);
xor U14724 (N_14724,N_13372,N_13108);
xnor U14725 (N_14725,N_13890,N_13562);
nand U14726 (N_14726,N_13875,N_13769);
nor U14727 (N_14727,N_13427,N_13967);
and U14728 (N_14728,N_13486,N_13161);
nand U14729 (N_14729,N_13645,N_13720);
or U14730 (N_14730,N_13800,N_13113);
nand U14731 (N_14731,N_13510,N_13490);
xor U14732 (N_14732,N_13934,N_13111);
nand U14733 (N_14733,N_13353,N_13142);
xor U14734 (N_14734,N_13459,N_13029);
or U14735 (N_14735,N_13708,N_13061);
or U14736 (N_14736,N_13972,N_13282);
xnor U14737 (N_14737,N_13596,N_13842);
nor U14738 (N_14738,N_13463,N_13922);
nand U14739 (N_14739,N_13456,N_13061);
nand U14740 (N_14740,N_13302,N_13378);
nand U14741 (N_14741,N_13385,N_13514);
nand U14742 (N_14742,N_13737,N_13880);
nand U14743 (N_14743,N_13816,N_13278);
xor U14744 (N_14744,N_13215,N_13178);
or U14745 (N_14745,N_13824,N_13054);
nor U14746 (N_14746,N_13645,N_13403);
and U14747 (N_14747,N_13455,N_13237);
or U14748 (N_14748,N_13570,N_13492);
and U14749 (N_14749,N_13882,N_13336);
and U14750 (N_14750,N_13737,N_13366);
and U14751 (N_14751,N_13863,N_13020);
xnor U14752 (N_14752,N_13824,N_13898);
xnor U14753 (N_14753,N_13011,N_13122);
nor U14754 (N_14754,N_13280,N_13856);
or U14755 (N_14755,N_13615,N_13618);
or U14756 (N_14756,N_13903,N_13759);
and U14757 (N_14757,N_13642,N_13204);
and U14758 (N_14758,N_13011,N_13231);
and U14759 (N_14759,N_13996,N_13975);
and U14760 (N_14760,N_13784,N_13512);
xnor U14761 (N_14761,N_13157,N_13401);
xnor U14762 (N_14762,N_13390,N_13746);
nor U14763 (N_14763,N_13030,N_13380);
nand U14764 (N_14764,N_13105,N_13869);
xor U14765 (N_14765,N_13185,N_13363);
or U14766 (N_14766,N_13799,N_13560);
nor U14767 (N_14767,N_13710,N_13677);
nand U14768 (N_14768,N_13633,N_13832);
nand U14769 (N_14769,N_13045,N_13950);
xnor U14770 (N_14770,N_13652,N_13834);
or U14771 (N_14771,N_13878,N_13885);
and U14772 (N_14772,N_13006,N_13963);
xor U14773 (N_14773,N_13810,N_13638);
xnor U14774 (N_14774,N_13994,N_13194);
or U14775 (N_14775,N_13533,N_13653);
nor U14776 (N_14776,N_13122,N_13417);
nor U14777 (N_14777,N_13201,N_13724);
xnor U14778 (N_14778,N_13397,N_13154);
xor U14779 (N_14779,N_13414,N_13042);
nor U14780 (N_14780,N_13338,N_13448);
or U14781 (N_14781,N_13189,N_13059);
xnor U14782 (N_14782,N_13135,N_13253);
or U14783 (N_14783,N_13928,N_13152);
xnor U14784 (N_14784,N_13284,N_13348);
or U14785 (N_14785,N_13920,N_13143);
nor U14786 (N_14786,N_13949,N_13805);
and U14787 (N_14787,N_13587,N_13260);
xnor U14788 (N_14788,N_13020,N_13560);
or U14789 (N_14789,N_13258,N_13278);
xnor U14790 (N_14790,N_13287,N_13752);
and U14791 (N_14791,N_13110,N_13849);
and U14792 (N_14792,N_13722,N_13367);
nor U14793 (N_14793,N_13960,N_13896);
or U14794 (N_14794,N_13921,N_13774);
nand U14795 (N_14795,N_13128,N_13037);
nand U14796 (N_14796,N_13000,N_13274);
nor U14797 (N_14797,N_13707,N_13601);
xnor U14798 (N_14798,N_13639,N_13713);
xnor U14799 (N_14799,N_13105,N_13465);
and U14800 (N_14800,N_13713,N_13283);
and U14801 (N_14801,N_13878,N_13877);
and U14802 (N_14802,N_13611,N_13320);
nand U14803 (N_14803,N_13076,N_13096);
and U14804 (N_14804,N_13785,N_13119);
nor U14805 (N_14805,N_13626,N_13991);
and U14806 (N_14806,N_13841,N_13022);
xnor U14807 (N_14807,N_13400,N_13613);
nor U14808 (N_14808,N_13367,N_13099);
or U14809 (N_14809,N_13510,N_13651);
xor U14810 (N_14810,N_13626,N_13940);
xor U14811 (N_14811,N_13707,N_13016);
nand U14812 (N_14812,N_13329,N_13443);
or U14813 (N_14813,N_13068,N_13240);
nand U14814 (N_14814,N_13835,N_13570);
or U14815 (N_14815,N_13164,N_13106);
nand U14816 (N_14816,N_13762,N_13313);
nand U14817 (N_14817,N_13653,N_13448);
and U14818 (N_14818,N_13433,N_13895);
and U14819 (N_14819,N_13513,N_13600);
nand U14820 (N_14820,N_13096,N_13941);
or U14821 (N_14821,N_13467,N_13552);
nand U14822 (N_14822,N_13116,N_13259);
and U14823 (N_14823,N_13154,N_13186);
nand U14824 (N_14824,N_13865,N_13410);
or U14825 (N_14825,N_13660,N_13542);
and U14826 (N_14826,N_13440,N_13394);
xnor U14827 (N_14827,N_13933,N_13467);
nand U14828 (N_14828,N_13875,N_13752);
and U14829 (N_14829,N_13427,N_13696);
nor U14830 (N_14830,N_13565,N_13098);
and U14831 (N_14831,N_13214,N_13612);
and U14832 (N_14832,N_13559,N_13418);
or U14833 (N_14833,N_13355,N_13548);
xnor U14834 (N_14834,N_13649,N_13348);
nor U14835 (N_14835,N_13390,N_13853);
nand U14836 (N_14836,N_13038,N_13197);
xor U14837 (N_14837,N_13221,N_13099);
and U14838 (N_14838,N_13382,N_13892);
xor U14839 (N_14839,N_13217,N_13821);
and U14840 (N_14840,N_13303,N_13389);
and U14841 (N_14841,N_13207,N_13352);
nand U14842 (N_14842,N_13975,N_13183);
xnor U14843 (N_14843,N_13429,N_13277);
xnor U14844 (N_14844,N_13917,N_13531);
nor U14845 (N_14845,N_13055,N_13589);
nor U14846 (N_14846,N_13677,N_13197);
or U14847 (N_14847,N_13509,N_13613);
and U14848 (N_14848,N_13695,N_13116);
xor U14849 (N_14849,N_13851,N_13930);
or U14850 (N_14850,N_13388,N_13680);
and U14851 (N_14851,N_13914,N_13842);
or U14852 (N_14852,N_13537,N_13989);
nand U14853 (N_14853,N_13370,N_13953);
xnor U14854 (N_14854,N_13437,N_13756);
and U14855 (N_14855,N_13123,N_13773);
or U14856 (N_14856,N_13427,N_13802);
nor U14857 (N_14857,N_13173,N_13188);
and U14858 (N_14858,N_13146,N_13097);
or U14859 (N_14859,N_13777,N_13883);
xnor U14860 (N_14860,N_13345,N_13967);
nand U14861 (N_14861,N_13421,N_13229);
or U14862 (N_14862,N_13493,N_13366);
xnor U14863 (N_14863,N_13249,N_13091);
nand U14864 (N_14864,N_13807,N_13535);
nand U14865 (N_14865,N_13031,N_13601);
nor U14866 (N_14866,N_13405,N_13346);
nor U14867 (N_14867,N_13854,N_13782);
nor U14868 (N_14868,N_13593,N_13480);
nand U14869 (N_14869,N_13334,N_13385);
or U14870 (N_14870,N_13223,N_13741);
and U14871 (N_14871,N_13741,N_13332);
nor U14872 (N_14872,N_13523,N_13296);
nor U14873 (N_14873,N_13125,N_13703);
nand U14874 (N_14874,N_13797,N_13465);
nand U14875 (N_14875,N_13661,N_13411);
xnor U14876 (N_14876,N_13439,N_13410);
or U14877 (N_14877,N_13557,N_13360);
or U14878 (N_14878,N_13296,N_13030);
or U14879 (N_14879,N_13824,N_13286);
and U14880 (N_14880,N_13674,N_13978);
nor U14881 (N_14881,N_13000,N_13964);
nand U14882 (N_14882,N_13860,N_13648);
or U14883 (N_14883,N_13726,N_13288);
or U14884 (N_14884,N_13141,N_13372);
xnor U14885 (N_14885,N_13538,N_13576);
and U14886 (N_14886,N_13170,N_13520);
nor U14887 (N_14887,N_13933,N_13998);
xnor U14888 (N_14888,N_13444,N_13727);
xor U14889 (N_14889,N_13905,N_13825);
xor U14890 (N_14890,N_13369,N_13692);
and U14891 (N_14891,N_13947,N_13566);
nor U14892 (N_14892,N_13984,N_13264);
nand U14893 (N_14893,N_13701,N_13977);
or U14894 (N_14894,N_13990,N_13344);
xnor U14895 (N_14895,N_13171,N_13002);
and U14896 (N_14896,N_13836,N_13584);
nand U14897 (N_14897,N_13360,N_13335);
nor U14898 (N_14898,N_13274,N_13656);
xor U14899 (N_14899,N_13484,N_13794);
nand U14900 (N_14900,N_13548,N_13950);
nor U14901 (N_14901,N_13621,N_13489);
nor U14902 (N_14902,N_13560,N_13062);
or U14903 (N_14903,N_13731,N_13136);
and U14904 (N_14904,N_13236,N_13141);
nor U14905 (N_14905,N_13975,N_13105);
or U14906 (N_14906,N_13030,N_13567);
or U14907 (N_14907,N_13451,N_13689);
xnor U14908 (N_14908,N_13226,N_13535);
or U14909 (N_14909,N_13432,N_13850);
nand U14910 (N_14910,N_13834,N_13305);
nor U14911 (N_14911,N_13332,N_13166);
nor U14912 (N_14912,N_13282,N_13090);
nor U14913 (N_14913,N_13109,N_13955);
nor U14914 (N_14914,N_13267,N_13503);
nand U14915 (N_14915,N_13716,N_13482);
nand U14916 (N_14916,N_13071,N_13043);
xor U14917 (N_14917,N_13026,N_13448);
or U14918 (N_14918,N_13548,N_13336);
and U14919 (N_14919,N_13166,N_13872);
and U14920 (N_14920,N_13356,N_13384);
or U14921 (N_14921,N_13839,N_13188);
nor U14922 (N_14922,N_13333,N_13190);
and U14923 (N_14923,N_13982,N_13376);
and U14924 (N_14924,N_13529,N_13078);
xor U14925 (N_14925,N_13951,N_13234);
nand U14926 (N_14926,N_13585,N_13347);
and U14927 (N_14927,N_13944,N_13857);
nor U14928 (N_14928,N_13822,N_13381);
nand U14929 (N_14929,N_13442,N_13284);
nor U14930 (N_14930,N_13649,N_13910);
or U14931 (N_14931,N_13026,N_13886);
xor U14932 (N_14932,N_13583,N_13210);
and U14933 (N_14933,N_13558,N_13286);
and U14934 (N_14934,N_13723,N_13457);
nor U14935 (N_14935,N_13993,N_13793);
and U14936 (N_14936,N_13177,N_13758);
nand U14937 (N_14937,N_13885,N_13521);
and U14938 (N_14938,N_13380,N_13325);
or U14939 (N_14939,N_13995,N_13537);
or U14940 (N_14940,N_13684,N_13995);
nor U14941 (N_14941,N_13088,N_13226);
nand U14942 (N_14942,N_13120,N_13414);
xnor U14943 (N_14943,N_13757,N_13344);
xor U14944 (N_14944,N_13395,N_13394);
nand U14945 (N_14945,N_13464,N_13241);
or U14946 (N_14946,N_13329,N_13396);
and U14947 (N_14947,N_13130,N_13631);
nor U14948 (N_14948,N_13704,N_13120);
and U14949 (N_14949,N_13006,N_13155);
nor U14950 (N_14950,N_13445,N_13541);
xnor U14951 (N_14951,N_13360,N_13251);
and U14952 (N_14952,N_13137,N_13134);
or U14953 (N_14953,N_13960,N_13973);
xnor U14954 (N_14954,N_13903,N_13563);
nand U14955 (N_14955,N_13493,N_13084);
nor U14956 (N_14956,N_13431,N_13053);
nor U14957 (N_14957,N_13843,N_13251);
xnor U14958 (N_14958,N_13565,N_13415);
nand U14959 (N_14959,N_13952,N_13749);
nor U14960 (N_14960,N_13156,N_13122);
xor U14961 (N_14961,N_13458,N_13253);
xnor U14962 (N_14962,N_13962,N_13598);
or U14963 (N_14963,N_13203,N_13667);
or U14964 (N_14964,N_13039,N_13994);
nand U14965 (N_14965,N_13201,N_13605);
xor U14966 (N_14966,N_13852,N_13990);
xnor U14967 (N_14967,N_13808,N_13807);
and U14968 (N_14968,N_13106,N_13761);
or U14969 (N_14969,N_13591,N_13538);
nand U14970 (N_14970,N_13988,N_13537);
and U14971 (N_14971,N_13548,N_13224);
nand U14972 (N_14972,N_13411,N_13816);
nand U14973 (N_14973,N_13416,N_13402);
nor U14974 (N_14974,N_13775,N_13022);
or U14975 (N_14975,N_13282,N_13738);
xnor U14976 (N_14976,N_13808,N_13153);
nand U14977 (N_14977,N_13652,N_13700);
and U14978 (N_14978,N_13564,N_13897);
and U14979 (N_14979,N_13915,N_13508);
nor U14980 (N_14980,N_13956,N_13984);
nor U14981 (N_14981,N_13742,N_13388);
xor U14982 (N_14982,N_13192,N_13217);
nand U14983 (N_14983,N_13197,N_13221);
xnor U14984 (N_14984,N_13064,N_13339);
and U14985 (N_14985,N_13670,N_13531);
nor U14986 (N_14986,N_13662,N_13123);
xnor U14987 (N_14987,N_13227,N_13436);
xnor U14988 (N_14988,N_13753,N_13071);
or U14989 (N_14989,N_13900,N_13211);
and U14990 (N_14990,N_13351,N_13276);
and U14991 (N_14991,N_13981,N_13102);
nor U14992 (N_14992,N_13875,N_13906);
and U14993 (N_14993,N_13635,N_13414);
and U14994 (N_14994,N_13211,N_13183);
and U14995 (N_14995,N_13747,N_13637);
xor U14996 (N_14996,N_13606,N_13385);
nand U14997 (N_14997,N_13789,N_13466);
nand U14998 (N_14998,N_13337,N_13897);
nor U14999 (N_14999,N_13925,N_13397);
or UO_0 (O_0,N_14707,N_14350);
xor UO_1 (O_1,N_14750,N_14600);
or UO_2 (O_2,N_14845,N_14433);
and UO_3 (O_3,N_14537,N_14729);
or UO_4 (O_4,N_14688,N_14692);
and UO_5 (O_5,N_14812,N_14076);
xor UO_6 (O_6,N_14749,N_14360);
nand UO_7 (O_7,N_14969,N_14910);
and UO_8 (O_8,N_14569,N_14813);
or UO_9 (O_9,N_14514,N_14663);
nand UO_10 (O_10,N_14238,N_14856);
and UO_11 (O_11,N_14735,N_14627);
xor UO_12 (O_12,N_14353,N_14030);
and UO_13 (O_13,N_14681,N_14649);
and UO_14 (O_14,N_14033,N_14876);
or UO_15 (O_15,N_14023,N_14134);
nor UO_16 (O_16,N_14348,N_14595);
nand UO_17 (O_17,N_14039,N_14215);
nand UO_18 (O_18,N_14788,N_14272);
or UO_19 (O_19,N_14046,N_14316);
nor UO_20 (O_20,N_14066,N_14269);
xor UO_21 (O_21,N_14024,N_14650);
or UO_22 (O_22,N_14993,N_14555);
xnor UO_23 (O_23,N_14774,N_14962);
xnor UO_24 (O_24,N_14295,N_14485);
or UO_25 (O_25,N_14769,N_14805);
xor UO_26 (O_26,N_14539,N_14850);
or UO_27 (O_27,N_14223,N_14868);
or UO_28 (O_28,N_14286,N_14331);
nor UO_29 (O_29,N_14712,N_14773);
and UO_30 (O_30,N_14109,N_14966);
and UO_31 (O_31,N_14148,N_14888);
xor UO_32 (O_32,N_14414,N_14654);
xnor UO_33 (O_33,N_14800,N_14280);
xnor UO_34 (O_34,N_14072,N_14963);
and UO_35 (O_35,N_14018,N_14077);
nor UO_36 (O_36,N_14621,N_14402);
or UO_37 (O_37,N_14975,N_14709);
nand UO_38 (O_38,N_14323,N_14655);
nand UO_39 (O_39,N_14113,N_14541);
nor UO_40 (O_40,N_14190,N_14778);
xor UO_41 (O_41,N_14670,N_14921);
or UO_42 (O_42,N_14300,N_14154);
xnor UO_43 (O_43,N_14596,N_14391);
nand UO_44 (O_44,N_14535,N_14886);
and UO_45 (O_45,N_14951,N_14898);
and UO_46 (O_46,N_14617,N_14753);
nand UO_47 (O_47,N_14846,N_14081);
or UO_48 (O_48,N_14458,N_14719);
nand UO_49 (O_49,N_14837,N_14984);
nor UO_50 (O_50,N_14647,N_14313);
nor UO_51 (O_51,N_14150,N_14147);
xnor UO_52 (O_52,N_14254,N_14032);
or UO_53 (O_53,N_14720,N_14802);
nor UO_54 (O_54,N_14151,N_14542);
or UO_55 (O_55,N_14387,N_14330);
and UO_56 (O_56,N_14156,N_14820);
and UO_57 (O_57,N_14763,N_14970);
nor UO_58 (O_58,N_14227,N_14204);
nor UO_59 (O_59,N_14472,N_14594);
nor UO_60 (O_60,N_14806,N_14599);
or UO_61 (O_61,N_14543,N_14138);
or UO_62 (O_62,N_14765,N_14088);
and UO_63 (O_63,N_14576,N_14112);
nor UO_64 (O_64,N_14176,N_14628);
or UO_65 (O_65,N_14416,N_14995);
or UO_66 (O_66,N_14834,N_14724);
nand UO_67 (O_67,N_14142,N_14009);
nand UO_68 (O_68,N_14690,N_14613);
nor UO_69 (O_69,N_14905,N_14397);
nor UO_70 (O_70,N_14140,N_14137);
or UO_71 (O_71,N_14925,N_14955);
or UO_72 (O_72,N_14352,N_14698);
or UO_73 (O_73,N_14872,N_14120);
nand UO_74 (O_74,N_14551,N_14478);
and UO_75 (O_75,N_14849,N_14567);
and UO_76 (O_76,N_14207,N_14721);
nand UO_77 (O_77,N_14145,N_14693);
or UO_78 (O_78,N_14909,N_14470);
or UO_79 (O_79,N_14431,N_14540);
or UO_80 (O_80,N_14530,N_14480);
xor UO_81 (O_81,N_14916,N_14987);
or UO_82 (O_82,N_14495,N_14327);
nor UO_83 (O_83,N_14632,N_14025);
nand UO_84 (O_84,N_14271,N_14777);
nand UO_85 (O_85,N_14240,N_14261);
and UO_86 (O_86,N_14011,N_14284);
nor UO_87 (O_87,N_14074,N_14489);
nand UO_88 (O_88,N_14922,N_14063);
nor UO_89 (O_89,N_14653,N_14465);
nor UO_90 (O_90,N_14205,N_14345);
and UO_91 (O_91,N_14793,N_14099);
and UO_92 (O_92,N_14186,N_14673);
and UO_93 (O_93,N_14061,N_14015);
and UO_94 (O_94,N_14528,N_14000);
nor UO_95 (O_95,N_14708,N_14052);
and UO_96 (O_96,N_14325,N_14432);
xnor UO_97 (O_97,N_14016,N_14761);
xor UO_98 (O_98,N_14726,N_14732);
nand UO_99 (O_99,N_14441,N_14890);
and UO_100 (O_100,N_14652,N_14319);
and UO_101 (O_101,N_14166,N_14310);
or UO_102 (O_102,N_14342,N_14349);
nand UO_103 (O_103,N_14376,N_14976);
nor UO_104 (O_104,N_14162,N_14079);
xnor UO_105 (O_105,N_14340,N_14210);
or UO_106 (O_106,N_14122,N_14427);
xor UO_107 (O_107,N_14356,N_14827);
or UO_108 (O_108,N_14633,N_14188);
and UO_109 (O_109,N_14742,N_14206);
nor UO_110 (O_110,N_14225,N_14260);
or UO_111 (O_111,N_14320,N_14045);
and UO_112 (O_112,N_14752,N_14466);
or UO_113 (O_113,N_14087,N_14386);
nor UO_114 (O_114,N_14611,N_14826);
nand UO_115 (O_115,N_14798,N_14727);
or UO_116 (O_116,N_14958,N_14956);
xnor UO_117 (O_117,N_14497,N_14307);
nand UO_118 (O_118,N_14588,N_14919);
xor UO_119 (O_119,N_14844,N_14091);
or UO_120 (O_120,N_14494,N_14343);
nand UO_121 (O_121,N_14629,N_14440);
nor UO_122 (O_122,N_14401,N_14159);
xor UO_123 (O_123,N_14518,N_14899);
xor UO_124 (O_124,N_14559,N_14579);
xor UO_125 (O_125,N_14104,N_14980);
nor UO_126 (O_126,N_14776,N_14604);
or UO_127 (O_127,N_14854,N_14593);
or UO_128 (O_128,N_14141,N_14029);
nor UO_129 (O_129,N_14398,N_14682);
nand UO_130 (O_130,N_14094,N_14783);
nor UO_131 (O_131,N_14680,N_14370);
and UO_132 (O_132,N_14329,N_14863);
nand UO_133 (O_133,N_14430,N_14843);
nor UO_134 (O_134,N_14454,N_14500);
or UO_135 (O_135,N_14483,N_14298);
or UO_136 (O_136,N_14879,N_14312);
nand UO_137 (O_137,N_14672,N_14108);
nor UO_138 (O_138,N_14838,N_14287);
nand UO_139 (O_139,N_14195,N_14381);
and UO_140 (O_140,N_14417,N_14625);
xnor UO_141 (O_141,N_14201,N_14125);
or UO_142 (O_142,N_14920,N_14338);
xor UO_143 (O_143,N_14887,N_14563);
or UO_144 (O_144,N_14981,N_14823);
and UO_145 (O_145,N_14321,N_14092);
nand UO_146 (O_146,N_14998,N_14198);
nand UO_147 (O_147,N_14219,N_14368);
and UO_148 (O_148,N_14436,N_14407);
and UO_149 (O_149,N_14311,N_14160);
nand UO_150 (O_150,N_14175,N_14279);
xnor UO_151 (O_151,N_14564,N_14169);
or UO_152 (O_152,N_14772,N_14220);
nor UO_153 (O_153,N_14102,N_14477);
nand UO_154 (O_154,N_14795,N_14382);
or UO_155 (O_155,N_14249,N_14013);
nand UO_156 (O_156,N_14933,N_14722);
nand UO_157 (O_157,N_14770,N_14133);
nor UO_158 (O_158,N_14245,N_14276);
xor UO_159 (O_159,N_14505,N_14118);
or UO_160 (O_160,N_14967,N_14359);
or UO_161 (O_161,N_14532,N_14103);
and UO_162 (O_162,N_14943,N_14114);
nor UO_163 (O_163,N_14105,N_14895);
or UO_164 (O_164,N_14244,N_14467);
or UO_165 (O_165,N_14631,N_14048);
nand UO_166 (O_166,N_14246,N_14193);
nand UO_167 (O_167,N_14351,N_14004);
nand UO_168 (O_168,N_14582,N_14334);
or UO_169 (O_169,N_14498,N_14506);
nand UO_170 (O_170,N_14581,N_14393);
or UO_171 (O_171,N_14314,N_14425);
xnor UO_172 (O_172,N_14136,N_14525);
xnor UO_173 (O_173,N_14828,N_14347);
nor UO_174 (O_174,N_14283,N_14728);
xor UO_175 (O_175,N_14930,N_14366);
or UO_176 (O_176,N_14258,N_14107);
nor UO_177 (O_177,N_14230,N_14253);
xor UO_178 (O_178,N_14678,N_14715);
nor UO_179 (O_179,N_14301,N_14549);
nor UO_180 (O_180,N_14664,N_14865);
nor UO_181 (O_181,N_14903,N_14622);
nor UO_182 (O_182,N_14167,N_14035);
and UO_183 (O_183,N_14282,N_14578);
nand UO_184 (O_184,N_14126,N_14262);
nor UO_185 (O_185,N_14404,N_14453);
or UO_186 (O_186,N_14346,N_14626);
xor UO_187 (O_187,N_14168,N_14096);
nand UO_188 (O_188,N_14158,N_14413);
nand UO_189 (O_189,N_14866,N_14143);
xor UO_190 (O_190,N_14211,N_14934);
and UO_191 (O_191,N_14270,N_14135);
nor UO_192 (O_192,N_14019,N_14713);
nand UO_193 (O_193,N_14180,N_14818);
xnor UO_194 (O_194,N_14651,N_14026);
xnor UO_195 (O_195,N_14624,N_14194);
xor UO_196 (O_196,N_14247,N_14869);
xor UO_197 (O_197,N_14531,N_14871);
and UO_198 (O_198,N_14557,N_14212);
or UO_199 (O_199,N_14702,N_14835);
and UO_200 (O_200,N_14476,N_14442);
or UO_201 (O_201,N_14444,N_14725);
nor UO_202 (O_202,N_14322,N_14510);
or UO_203 (O_203,N_14296,N_14131);
and UO_204 (O_204,N_14764,N_14511);
nand UO_205 (O_205,N_14691,N_14926);
or UO_206 (O_206,N_14419,N_14801);
and UO_207 (O_207,N_14751,N_14685);
and UO_208 (O_208,N_14208,N_14568);
and UO_209 (O_209,N_14289,N_14915);
nand UO_210 (O_210,N_14251,N_14332);
and UO_211 (O_211,N_14878,N_14789);
xor UO_212 (O_212,N_14181,N_14139);
nor UO_213 (O_213,N_14456,N_14947);
xor UO_214 (O_214,N_14928,N_14936);
nand UO_215 (O_215,N_14517,N_14297);
nand UO_216 (O_216,N_14504,N_14710);
and UO_217 (O_217,N_14609,N_14833);
and UO_218 (O_218,N_14191,N_14931);
nand UO_219 (O_219,N_14723,N_14526);
and UO_220 (O_220,N_14968,N_14819);
and UO_221 (O_221,N_14304,N_14659);
xnor UO_222 (O_222,N_14946,N_14512);
xor UO_223 (O_223,N_14683,N_14572);
nor UO_224 (O_224,N_14460,N_14080);
nor UO_225 (O_225,N_14775,N_14335);
and UO_226 (O_226,N_14097,N_14503);
xnor UO_227 (O_227,N_14027,N_14084);
and UO_228 (O_228,N_14830,N_14734);
nor UO_229 (O_229,N_14950,N_14640);
xor UO_230 (O_230,N_14577,N_14235);
xor UO_231 (O_231,N_14157,N_14389);
nand UO_232 (O_232,N_14999,N_14612);
nor UO_233 (O_233,N_14883,N_14447);
nor UO_234 (O_234,N_14420,N_14885);
xor UO_235 (O_235,N_14941,N_14248);
and UO_236 (O_236,N_14014,N_14214);
nor UO_237 (O_237,N_14893,N_14877);
nor UO_238 (O_238,N_14446,N_14001);
xnor UO_239 (O_239,N_14994,N_14974);
and UO_240 (O_240,N_14400,N_14779);
or UO_241 (O_241,N_14859,N_14508);
xor UO_242 (O_242,N_14816,N_14686);
nor UO_243 (O_243,N_14667,N_14803);
nor UO_244 (O_244,N_14439,N_14303);
nand UO_245 (O_245,N_14855,N_14443);
nand UO_246 (O_246,N_14049,N_14583);
and UO_247 (O_247,N_14768,N_14513);
and UO_248 (O_248,N_14379,N_14597);
or UO_249 (O_249,N_14315,N_14605);
nand UO_250 (O_250,N_14042,N_14545);
or UO_251 (O_251,N_14797,N_14882);
and UO_252 (O_252,N_14203,N_14115);
or UO_253 (O_253,N_14089,N_14556);
and UO_254 (O_254,N_14471,N_14550);
xor UO_255 (O_255,N_14744,N_14022);
nand UO_256 (O_256,N_14435,N_14365);
and UO_257 (O_257,N_14964,N_14068);
nand UO_258 (O_258,N_14252,N_14308);
and UO_259 (O_259,N_14945,N_14491);
or UO_260 (O_260,N_14700,N_14957);
nor UO_261 (O_261,N_14705,N_14418);
nand UO_262 (O_262,N_14699,N_14533);
or UO_263 (O_263,N_14357,N_14601);
xnor UO_264 (O_264,N_14747,N_14236);
and UO_265 (O_265,N_14374,N_14638);
nand UO_266 (O_266,N_14237,N_14410);
or UO_267 (O_267,N_14731,N_14992);
xnor UO_268 (O_268,N_14684,N_14677);
and UO_269 (O_269,N_14170,N_14012);
and UO_270 (O_270,N_14179,N_14810);
xnor UO_271 (O_271,N_14986,N_14644);
or UO_272 (O_272,N_14554,N_14274);
nor UO_273 (O_273,N_14369,N_14294);
and UO_274 (O_274,N_14977,N_14646);
nor UO_275 (O_275,N_14474,N_14257);
nand UO_276 (O_276,N_14917,N_14047);
and UO_277 (O_277,N_14982,N_14570);
xor UO_278 (O_278,N_14390,N_14598);
nand UO_279 (O_279,N_14161,N_14703);
nor UO_280 (O_280,N_14372,N_14266);
nor UO_281 (O_281,N_14486,N_14146);
or UO_282 (O_282,N_14536,N_14488);
nor UO_283 (O_283,N_14317,N_14522);
and UO_284 (O_284,N_14501,N_14095);
nand UO_285 (O_285,N_14658,N_14694);
xor UO_286 (O_286,N_14464,N_14060);
nand UO_287 (O_287,N_14527,N_14200);
xnor UO_288 (O_288,N_14949,N_14794);
xor UO_289 (O_289,N_14232,N_14424);
nor UO_290 (O_290,N_14880,N_14648);
nor UO_291 (O_291,N_14028,N_14187);
xnor UO_292 (O_292,N_14755,N_14911);
nor UO_293 (O_293,N_14552,N_14451);
and UO_294 (O_294,N_14469,N_14121);
nor UO_295 (O_295,N_14538,N_14737);
nand UO_296 (O_296,N_14071,N_14100);
nand UO_297 (O_297,N_14429,N_14054);
xor UO_298 (O_298,N_14894,N_14717);
xor UO_299 (O_299,N_14757,N_14050);
nor UO_300 (O_300,N_14056,N_14935);
xor UO_301 (O_301,N_14116,N_14098);
nor UO_302 (O_302,N_14623,N_14005);
or UO_303 (O_303,N_14267,N_14086);
or UO_304 (O_304,N_14634,N_14502);
or UO_305 (O_305,N_14814,N_14473);
xnor UO_306 (O_306,N_14620,N_14383);
and UO_307 (O_307,N_14106,N_14889);
xnor UO_308 (O_308,N_14288,N_14457);
or UO_309 (O_309,N_14388,N_14078);
nand UO_310 (O_310,N_14990,N_14636);
xnor UO_311 (O_311,N_14479,N_14580);
nor UO_312 (O_312,N_14746,N_14197);
and UO_313 (O_313,N_14041,N_14165);
and UO_314 (O_314,N_14482,N_14129);
xnor UO_315 (O_315,N_14585,N_14881);
and UO_316 (O_316,N_14913,N_14006);
nor UO_317 (O_317,N_14864,N_14792);
nor UO_318 (O_318,N_14831,N_14277);
or UO_319 (O_319,N_14704,N_14224);
nor UO_320 (O_320,N_14127,N_14733);
nand UO_321 (O_321,N_14155,N_14676);
xor UO_322 (O_322,N_14534,N_14637);
nand UO_323 (O_323,N_14496,N_14822);
nor UO_324 (O_324,N_14020,N_14739);
or UO_325 (O_325,N_14101,N_14767);
nand UO_326 (O_326,N_14562,N_14445);
or UO_327 (O_327,N_14616,N_14674);
nor UO_328 (O_328,N_14697,N_14668);
or UO_329 (O_329,N_14642,N_14748);
or UO_330 (O_330,N_14860,N_14031);
or UO_331 (O_331,N_14111,N_14468);
nor UO_332 (O_332,N_14250,N_14043);
xor UO_333 (O_333,N_14278,N_14972);
or UO_334 (O_334,N_14265,N_14602);
or UO_335 (O_335,N_14759,N_14932);
and UO_336 (O_336,N_14988,N_14592);
or UO_337 (O_337,N_14051,N_14953);
or UO_338 (O_338,N_14036,N_14874);
xor UO_339 (O_339,N_14069,N_14840);
nor UO_340 (O_340,N_14259,N_14177);
xor UO_341 (O_341,N_14085,N_14809);
nand UO_342 (O_342,N_14918,N_14487);
xnor UO_343 (O_343,N_14523,N_14363);
nand UO_344 (O_344,N_14128,N_14093);
or UO_345 (O_345,N_14558,N_14607);
or UO_346 (O_346,N_14875,N_14784);
nor UO_347 (O_347,N_14660,N_14754);
nor UO_348 (O_348,N_14461,N_14228);
nand UO_349 (O_349,N_14293,N_14804);
nor UO_350 (O_350,N_14217,N_14218);
and UO_351 (O_351,N_14643,N_14153);
or UO_352 (O_352,N_14689,N_14870);
nor UO_353 (O_353,N_14841,N_14760);
nand UO_354 (O_354,N_14184,N_14825);
nor UO_355 (O_355,N_14229,N_14507);
xnor UO_356 (O_356,N_14944,N_14861);
xor UO_357 (O_357,N_14687,N_14178);
and UO_358 (O_358,N_14891,N_14971);
xor UO_359 (O_359,N_14923,N_14952);
nand UO_360 (O_360,N_14738,N_14399);
xnor UO_361 (O_361,N_14324,N_14242);
xnor UO_362 (O_362,N_14927,N_14010);
nor UO_363 (O_363,N_14213,N_14671);
nor UO_364 (O_364,N_14481,N_14392);
nand UO_365 (O_365,N_14853,N_14371);
and UO_366 (O_366,N_14124,N_14450);
nand UO_367 (O_367,N_14897,N_14939);
nand UO_368 (O_368,N_14657,N_14589);
nand UO_369 (O_369,N_14786,N_14339);
and UO_370 (O_370,N_14997,N_14665);
nor UO_371 (O_371,N_14173,N_14736);
or UO_372 (O_372,N_14358,N_14756);
nand UO_373 (O_373,N_14333,N_14566);
nor UO_374 (O_374,N_14979,N_14422);
or UO_375 (O_375,N_14233,N_14851);
or UO_376 (O_376,N_14038,N_14591);
and UO_377 (O_377,N_14183,N_14209);
or UO_378 (O_378,N_14438,N_14529);
and UO_379 (O_379,N_14571,N_14256);
nor UO_380 (O_380,N_14202,N_14790);
nand UO_381 (O_381,N_14847,N_14395);
nor UO_382 (O_382,N_14908,N_14985);
xor UO_383 (O_383,N_14515,N_14618);
and UO_384 (O_384,N_14065,N_14002);
nand UO_385 (O_385,N_14394,N_14003);
nor UO_386 (O_386,N_14884,N_14415);
or UO_387 (O_387,N_14044,N_14901);
xnor UO_388 (O_388,N_14055,N_14264);
xor UO_389 (O_389,N_14608,N_14403);
or UO_390 (O_390,N_14836,N_14546);
or UO_391 (O_391,N_14318,N_14808);
xnor UO_392 (O_392,N_14656,N_14679);
or UO_393 (O_393,N_14408,N_14163);
nand UO_394 (O_394,N_14701,N_14852);
and UO_395 (O_395,N_14791,N_14706);
xnor UO_396 (O_396,N_14412,N_14714);
or UO_397 (O_397,N_14058,N_14263);
and UO_398 (O_398,N_14017,N_14938);
nor UO_399 (O_399,N_14615,N_14275);
xor UO_400 (O_400,N_14377,N_14815);
xor UO_401 (O_401,N_14575,N_14299);
and UO_402 (O_402,N_14164,N_14355);
xnor UO_403 (O_403,N_14606,N_14639);
or UO_404 (O_404,N_14306,N_14520);
nor UO_405 (O_405,N_14149,N_14516);
or UO_406 (O_406,N_14904,N_14452);
nor UO_407 (O_407,N_14172,N_14302);
nor UO_408 (O_408,N_14455,N_14716);
xor UO_409 (O_409,N_14243,N_14123);
nor UO_410 (O_410,N_14959,N_14226);
nand UO_411 (O_411,N_14059,N_14584);
nand UO_412 (O_412,N_14573,N_14428);
nor UO_413 (O_413,N_14780,N_14221);
or UO_414 (O_414,N_14799,N_14782);
nor UO_415 (O_415,N_14216,N_14586);
or UO_416 (O_416,N_14380,N_14130);
and UO_417 (O_417,N_14900,N_14189);
xor UO_418 (O_418,N_14222,N_14367);
xnor UO_419 (O_419,N_14057,N_14336);
or UO_420 (O_420,N_14948,N_14423);
xnor UO_421 (O_421,N_14940,N_14560);
xnor UO_422 (O_422,N_14796,N_14290);
xor UO_423 (O_423,N_14070,N_14305);
nand UO_424 (O_424,N_14448,N_14519);
xnor UO_425 (O_425,N_14090,N_14848);
nand UO_426 (O_426,N_14973,N_14082);
nor UO_427 (O_427,N_14929,N_14341);
nor UO_428 (O_428,N_14661,N_14730);
nor UO_429 (O_429,N_14405,N_14766);
nor UO_430 (O_430,N_14040,N_14490);
or UO_431 (O_431,N_14745,N_14034);
xnor UO_432 (O_432,N_14185,N_14544);
nand UO_433 (O_433,N_14174,N_14037);
xor UO_434 (O_434,N_14378,N_14493);
nor UO_435 (O_435,N_14337,N_14914);
nand UO_436 (O_436,N_14053,N_14811);
xnor UO_437 (O_437,N_14696,N_14384);
xor UO_438 (O_438,N_14965,N_14459);
and UO_439 (O_439,N_14561,N_14907);
and UO_440 (O_440,N_14857,N_14326);
nand UO_441 (O_441,N_14906,N_14364);
nor UO_442 (O_442,N_14695,N_14182);
and UO_443 (O_443,N_14492,N_14421);
xor UO_444 (O_444,N_14449,N_14375);
or UO_445 (O_445,N_14743,N_14630);
xnor UO_446 (O_446,N_14064,N_14762);
nand UO_447 (O_447,N_14829,N_14821);
nor UO_448 (O_448,N_14021,N_14824);
or UO_449 (O_449,N_14565,N_14989);
or UO_450 (O_450,N_14110,N_14832);
nand UO_451 (O_451,N_14171,N_14902);
xor UO_452 (O_452,N_14385,N_14409);
xnor UO_453 (O_453,N_14574,N_14067);
or UO_454 (O_454,N_14281,N_14771);
nand UO_455 (O_455,N_14132,N_14231);
nand UO_456 (O_456,N_14807,N_14666);
and UO_457 (O_457,N_14521,N_14268);
nor UO_458 (O_458,N_14741,N_14344);
nand UO_459 (O_459,N_14484,N_14411);
nor UO_460 (O_460,N_14960,N_14273);
and UO_461 (O_461,N_14373,N_14475);
xor UO_462 (O_462,N_14961,N_14285);
and UO_463 (O_463,N_14309,N_14144);
xnor UO_464 (O_464,N_14437,N_14610);
and UO_465 (O_465,N_14007,N_14152);
and UO_466 (O_466,N_14912,N_14787);
nand UO_467 (O_467,N_14645,N_14509);
and UO_468 (O_468,N_14292,N_14553);
xor UO_469 (O_469,N_14758,N_14083);
nand UO_470 (O_470,N_14937,N_14396);
or UO_471 (O_471,N_14117,N_14196);
xor UO_472 (O_472,N_14842,N_14675);
nor UO_473 (O_473,N_14075,N_14635);
nor UO_474 (O_474,N_14619,N_14858);
or UO_475 (O_475,N_14354,N_14192);
nor UO_476 (O_476,N_14996,N_14867);
and UO_477 (O_477,N_14669,N_14839);
nor UO_478 (O_478,N_14978,N_14062);
xnor UO_479 (O_479,N_14817,N_14361);
and UO_480 (O_480,N_14896,N_14718);
xor UO_481 (O_481,N_14073,N_14983);
and UO_482 (O_482,N_14641,N_14547);
nor UO_483 (O_483,N_14662,N_14524);
and UO_484 (O_484,N_14862,N_14740);
xnor UO_485 (O_485,N_14954,N_14942);
and UO_486 (O_486,N_14499,N_14781);
nand UO_487 (O_487,N_14434,N_14587);
or UO_488 (O_488,N_14991,N_14119);
or UO_489 (O_489,N_14463,N_14614);
and UO_490 (O_490,N_14785,N_14924);
or UO_491 (O_491,N_14241,N_14426);
xnor UO_492 (O_492,N_14873,N_14328);
nor UO_493 (O_493,N_14291,N_14234);
and UO_494 (O_494,N_14462,N_14199);
or UO_495 (O_495,N_14548,N_14362);
nor UO_496 (O_496,N_14711,N_14892);
or UO_497 (O_497,N_14008,N_14406);
and UO_498 (O_498,N_14590,N_14239);
xor UO_499 (O_499,N_14255,N_14603);
nor UO_500 (O_500,N_14848,N_14058);
nor UO_501 (O_501,N_14730,N_14871);
and UO_502 (O_502,N_14565,N_14510);
and UO_503 (O_503,N_14626,N_14241);
xor UO_504 (O_504,N_14275,N_14908);
nor UO_505 (O_505,N_14590,N_14930);
nand UO_506 (O_506,N_14735,N_14612);
xnor UO_507 (O_507,N_14873,N_14676);
nor UO_508 (O_508,N_14006,N_14834);
or UO_509 (O_509,N_14399,N_14229);
nor UO_510 (O_510,N_14333,N_14437);
or UO_511 (O_511,N_14815,N_14249);
nand UO_512 (O_512,N_14328,N_14841);
nand UO_513 (O_513,N_14844,N_14085);
and UO_514 (O_514,N_14032,N_14193);
nor UO_515 (O_515,N_14150,N_14851);
nor UO_516 (O_516,N_14931,N_14798);
nor UO_517 (O_517,N_14268,N_14736);
nand UO_518 (O_518,N_14959,N_14704);
or UO_519 (O_519,N_14500,N_14094);
and UO_520 (O_520,N_14394,N_14573);
nand UO_521 (O_521,N_14043,N_14637);
nand UO_522 (O_522,N_14071,N_14927);
or UO_523 (O_523,N_14009,N_14950);
nand UO_524 (O_524,N_14618,N_14233);
and UO_525 (O_525,N_14931,N_14479);
and UO_526 (O_526,N_14540,N_14918);
and UO_527 (O_527,N_14520,N_14413);
nor UO_528 (O_528,N_14639,N_14592);
xor UO_529 (O_529,N_14713,N_14397);
or UO_530 (O_530,N_14034,N_14284);
xnor UO_531 (O_531,N_14339,N_14637);
xnor UO_532 (O_532,N_14764,N_14790);
nor UO_533 (O_533,N_14028,N_14427);
or UO_534 (O_534,N_14514,N_14706);
or UO_535 (O_535,N_14701,N_14567);
or UO_536 (O_536,N_14566,N_14976);
or UO_537 (O_537,N_14566,N_14314);
nand UO_538 (O_538,N_14680,N_14492);
or UO_539 (O_539,N_14935,N_14479);
nand UO_540 (O_540,N_14139,N_14035);
or UO_541 (O_541,N_14871,N_14793);
or UO_542 (O_542,N_14738,N_14964);
xnor UO_543 (O_543,N_14391,N_14697);
nand UO_544 (O_544,N_14738,N_14463);
nand UO_545 (O_545,N_14725,N_14898);
and UO_546 (O_546,N_14683,N_14534);
nand UO_547 (O_547,N_14121,N_14354);
nor UO_548 (O_548,N_14774,N_14666);
and UO_549 (O_549,N_14536,N_14857);
or UO_550 (O_550,N_14502,N_14796);
and UO_551 (O_551,N_14687,N_14221);
nand UO_552 (O_552,N_14412,N_14434);
and UO_553 (O_553,N_14541,N_14206);
nand UO_554 (O_554,N_14147,N_14399);
and UO_555 (O_555,N_14152,N_14798);
nor UO_556 (O_556,N_14835,N_14943);
nor UO_557 (O_557,N_14269,N_14866);
or UO_558 (O_558,N_14464,N_14067);
or UO_559 (O_559,N_14481,N_14364);
nor UO_560 (O_560,N_14861,N_14381);
xor UO_561 (O_561,N_14176,N_14599);
nor UO_562 (O_562,N_14540,N_14462);
xnor UO_563 (O_563,N_14153,N_14430);
or UO_564 (O_564,N_14861,N_14800);
nor UO_565 (O_565,N_14483,N_14435);
xnor UO_566 (O_566,N_14892,N_14664);
or UO_567 (O_567,N_14834,N_14034);
xor UO_568 (O_568,N_14950,N_14515);
and UO_569 (O_569,N_14543,N_14515);
or UO_570 (O_570,N_14767,N_14179);
or UO_571 (O_571,N_14676,N_14636);
xnor UO_572 (O_572,N_14528,N_14493);
or UO_573 (O_573,N_14518,N_14202);
and UO_574 (O_574,N_14612,N_14207);
nand UO_575 (O_575,N_14353,N_14829);
and UO_576 (O_576,N_14412,N_14052);
nand UO_577 (O_577,N_14118,N_14168);
nand UO_578 (O_578,N_14550,N_14845);
xor UO_579 (O_579,N_14650,N_14705);
nand UO_580 (O_580,N_14999,N_14734);
or UO_581 (O_581,N_14879,N_14356);
nor UO_582 (O_582,N_14398,N_14008);
and UO_583 (O_583,N_14893,N_14808);
xnor UO_584 (O_584,N_14201,N_14087);
nor UO_585 (O_585,N_14385,N_14750);
nor UO_586 (O_586,N_14102,N_14238);
or UO_587 (O_587,N_14013,N_14170);
nor UO_588 (O_588,N_14012,N_14758);
or UO_589 (O_589,N_14516,N_14771);
and UO_590 (O_590,N_14934,N_14071);
xnor UO_591 (O_591,N_14961,N_14637);
nor UO_592 (O_592,N_14318,N_14195);
xnor UO_593 (O_593,N_14455,N_14446);
and UO_594 (O_594,N_14754,N_14561);
and UO_595 (O_595,N_14938,N_14911);
nor UO_596 (O_596,N_14773,N_14084);
and UO_597 (O_597,N_14593,N_14620);
nand UO_598 (O_598,N_14677,N_14744);
xnor UO_599 (O_599,N_14899,N_14877);
nand UO_600 (O_600,N_14291,N_14576);
nor UO_601 (O_601,N_14294,N_14402);
xor UO_602 (O_602,N_14205,N_14279);
xnor UO_603 (O_603,N_14554,N_14894);
nand UO_604 (O_604,N_14476,N_14952);
nand UO_605 (O_605,N_14330,N_14930);
and UO_606 (O_606,N_14345,N_14203);
nand UO_607 (O_607,N_14206,N_14486);
xnor UO_608 (O_608,N_14170,N_14239);
xnor UO_609 (O_609,N_14930,N_14430);
nor UO_610 (O_610,N_14465,N_14412);
nor UO_611 (O_611,N_14667,N_14523);
nand UO_612 (O_612,N_14711,N_14386);
nand UO_613 (O_613,N_14657,N_14317);
or UO_614 (O_614,N_14602,N_14697);
xnor UO_615 (O_615,N_14826,N_14190);
nand UO_616 (O_616,N_14262,N_14979);
nor UO_617 (O_617,N_14953,N_14693);
xor UO_618 (O_618,N_14331,N_14667);
or UO_619 (O_619,N_14997,N_14253);
nor UO_620 (O_620,N_14175,N_14209);
nor UO_621 (O_621,N_14935,N_14579);
nand UO_622 (O_622,N_14369,N_14923);
and UO_623 (O_623,N_14398,N_14511);
or UO_624 (O_624,N_14489,N_14742);
or UO_625 (O_625,N_14085,N_14838);
and UO_626 (O_626,N_14112,N_14343);
xor UO_627 (O_627,N_14730,N_14344);
nand UO_628 (O_628,N_14896,N_14315);
and UO_629 (O_629,N_14400,N_14116);
nand UO_630 (O_630,N_14220,N_14482);
or UO_631 (O_631,N_14701,N_14681);
nor UO_632 (O_632,N_14894,N_14212);
xnor UO_633 (O_633,N_14813,N_14462);
nor UO_634 (O_634,N_14861,N_14076);
xor UO_635 (O_635,N_14198,N_14010);
or UO_636 (O_636,N_14077,N_14017);
nor UO_637 (O_637,N_14107,N_14537);
nand UO_638 (O_638,N_14027,N_14579);
nand UO_639 (O_639,N_14712,N_14246);
and UO_640 (O_640,N_14313,N_14798);
or UO_641 (O_641,N_14844,N_14534);
nor UO_642 (O_642,N_14153,N_14025);
or UO_643 (O_643,N_14169,N_14798);
xnor UO_644 (O_644,N_14758,N_14543);
and UO_645 (O_645,N_14050,N_14395);
or UO_646 (O_646,N_14905,N_14636);
and UO_647 (O_647,N_14119,N_14686);
nand UO_648 (O_648,N_14911,N_14003);
nand UO_649 (O_649,N_14643,N_14323);
nor UO_650 (O_650,N_14655,N_14420);
xor UO_651 (O_651,N_14307,N_14765);
and UO_652 (O_652,N_14461,N_14752);
xor UO_653 (O_653,N_14759,N_14221);
xnor UO_654 (O_654,N_14618,N_14401);
nand UO_655 (O_655,N_14044,N_14515);
xor UO_656 (O_656,N_14563,N_14128);
xnor UO_657 (O_657,N_14937,N_14576);
or UO_658 (O_658,N_14291,N_14513);
or UO_659 (O_659,N_14611,N_14707);
nor UO_660 (O_660,N_14121,N_14730);
nor UO_661 (O_661,N_14751,N_14478);
or UO_662 (O_662,N_14957,N_14807);
and UO_663 (O_663,N_14077,N_14627);
or UO_664 (O_664,N_14834,N_14945);
nand UO_665 (O_665,N_14244,N_14601);
and UO_666 (O_666,N_14796,N_14511);
or UO_667 (O_667,N_14512,N_14971);
and UO_668 (O_668,N_14300,N_14428);
nand UO_669 (O_669,N_14218,N_14975);
or UO_670 (O_670,N_14359,N_14749);
nor UO_671 (O_671,N_14043,N_14505);
xor UO_672 (O_672,N_14094,N_14415);
xnor UO_673 (O_673,N_14037,N_14432);
and UO_674 (O_674,N_14274,N_14349);
nand UO_675 (O_675,N_14316,N_14445);
xnor UO_676 (O_676,N_14553,N_14615);
nand UO_677 (O_677,N_14563,N_14421);
or UO_678 (O_678,N_14883,N_14006);
or UO_679 (O_679,N_14817,N_14014);
nor UO_680 (O_680,N_14631,N_14766);
nor UO_681 (O_681,N_14062,N_14479);
xor UO_682 (O_682,N_14415,N_14998);
or UO_683 (O_683,N_14639,N_14504);
nor UO_684 (O_684,N_14748,N_14328);
nand UO_685 (O_685,N_14998,N_14576);
nor UO_686 (O_686,N_14498,N_14143);
or UO_687 (O_687,N_14562,N_14764);
and UO_688 (O_688,N_14882,N_14131);
nor UO_689 (O_689,N_14593,N_14139);
nand UO_690 (O_690,N_14807,N_14971);
xor UO_691 (O_691,N_14642,N_14984);
xor UO_692 (O_692,N_14435,N_14878);
or UO_693 (O_693,N_14654,N_14652);
or UO_694 (O_694,N_14370,N_14471);
and UO_695 (O_695,N_14311,N_14526);
xor UO_696 (O_696,N_14918,N_14191);
nor UO_697 (O_697,N_14438,N_14123);
and UO_698 (O_698,N_14583,N_14481);
xor UO_699 (O_699,N_14634,N_14224);
nor UO_700 (O_700,N_14419,N_14830);
nor UO_701 (O_701,N_14373,N_14634);
nand UO_702 (O_702,N_14514,N_14819);
nand UO_703 (O_703,N_14628,N_14902);
xor UO_704 (O_704,N_14484,N_14933);
or UO_705 (O_705,N_14815,N_14059);
nand UO_706 (O_706,N_14949,N_14349);
or UO_707 (O_707,N_14405,N_14947);
nor UO_708 (O_708,N_14553,N_14180);
nor UO_709 (O_709,N_14163,N_14470);
xor UO_710 (O_710,N_14908,N_14339);
nand UO_711 (O_711,N_14216,N_14027);
and UO_712 (O_712,N_14201,N_14154);
or UO_713 (O_713,N_14533,N_14665);
nand UO_714 (O_714,N_14714,N_14967);
nand UO_715 (O_715,N_14730,N_14200);
and UO_716 (O_716,N_14624,N_14648);
nand UO_717 (O_717,N_14441,N_14471);
nor UO_718 (O_718,N_14313,N_14899);
xnor UO_719 (O_719,N_14447,N_14693);
xnor UO_720 (O_720,N_14543,N_14133);
nand UO_721 (O_721,N_14140,N_14980);
nor UO_722 (O_722,N_14361,N_14769);
xor UO_723 (O_723,N_14317,N_14282);
and UO_724 (O_724,N_14348,N_14764);
nand UO_725 (O_725,N_14540,N_14140);
and UO_726 (O_726,N_14425,N_14233);
nand UO_727 (O_727,N_14444,N_14757);
and UO_728 (O_728,N_14946,N_14546);
and UO_729 (O_729,N_14181,N_14642);
or UO_730 (O_730,N_14859,N_14885);
nand UO_731 (O_731,N_14899,N_14953);
nand UO_732 (O_732,N_14903,N_14886);
and UO_733 (O_733,N_14579,N_14090);
nor UO_734 (O_734,N_14614,N_14314);
nand UO_735 (O_735,N_14046,N_14277);
nand UO_736 (O_736,N_14714,N_14110);
nor UO_737 (O_737,N_14987,N_14549);
xor UO_738 (O_738,N_14430,N_14768);
nand UO_739 (O_739,N_14008,N_14000);
nand UO_740 (O_740,N_14612,N_14905);
and UO_741 (O_741,N_14907,N_14043);
or UO_742 (O_742,N_14600,N_14605);
and UO_743 (O_743,N_14169,N_14795);
and UO_744 (O_744,N_14472,N_14815);
or UO_745 (O_745,N_14200,N_14984);
or UO_746 (O_746,N_14922,N_14645);
nor UO_747 (O_747,N_14412,N_14692);
nand UO_748 (O_748,N_14326,N_14482);
and UO_749 (O_749,N_14951,N_14263);
or UO_750 (O_750,N_14793,N_14887);
nand UO_751 (O_751,N_14639,N_14097);
nand UO_752 (O_752,N_14746,N_14806);
nand UO_753 (O_753,N_14260,N_14808);
and UO_754 (O_754,N_14754,N_14251);
and UO_755 (O_755,N_14975,N_14420);
nand UO_756 (O_756,N_14356,N_14073);
xor UO_757 (O_757,N_14482,N_14313);
and UO_758 (O_758,N_14379,N_14517);
xor UO_759 (O_759,N_14968,N_14182);
xnor UO_760 (O_760,N_14438,N_14259);
nor UO_761 (O_761,N_14884,N_14947);
and UO_762 (O_762,N_14193,N_14713);
and UO_763 (O_763,N_14105,N_14248);
xor UO_764 (O_764,N_14220,N_14078);
or UO_765 (O_765,N_14926,N_14228);
nand UO_766 (O_766,N_14992,N_14024);
and UO_767 (O_767,N_14372,N_14165);
nand UO_768 (O_768,N_14639,N_14022);
xnor UO_769 (O_769,N_14519,N_14851);
and UO_770 (O_770,N_14628,N_14748);
nor UO_771 (O_771,N_14685,N_14957);
or UO_772 (O_772,N_14554,N_14057);
nor UO_773 (O_773,N_14639,N_14621);
xor UO_774 (O_774,N_14174,N_14689);
nor UO_775 (O_775,N_14123,N_14598);
xnor UO_776 (O_776,N_14524,N_14604);
or UO_777 (O_777,N_14635,N_14567);
or UO_778 (O_778,N_14399,N_14267);
nand UO_779 (O_779,N_14131,N_14579);
nand UO_780 (O_780,N_14272,N_14185);
and UO_781 (O_781,N_14701,N_14052);
xnor UO_782 (O_782,N_14293,N_14474);
xnor UO_783 (O_783,N_14395,N_14445);
xnor UO_784 (O_784,N_14454,N_14741);
xor UO_785 (O_785,N_14404,N_14390);
nand UO_786 (O_786,N_14561,N_14166);
or UO_787 (O_787,N_14499,N_14658);
nor UO_788 (O_788,N_14252,N_14646);
and UO_789 (O_789,N_14527,N_14155);
nand UO_790 (O_790,N_14549,N_14684);
nor UO_791 (O_791,N_14496,N_14600);
and UO_792 (O_792,N_14771,N_14156);
or UO_793 (O_793,N_14081,N_14107);
or UO_794 (O_794,N_14211,N_14154);
and UO_795 (O_795,N_14545,N_14600);
or UO_796 (O_796,N_14397,N_14927);
or UO_797 (O_797,N_14948,N_14420);
xnor UO_798 (O_798,N_14523,N_14142);
and UO_799 (O_799,N_14782,N_14151);
and UO_800 (O_800,N_14976,N_14782);
nor UO_801 (O_801,N_14406,N_14637);
nor UO_802 (O_802,N_14393,N_14514);
and UO_803 (O_803,N_14808,N_14629);
and UO_804 (O_804,N_14569,N_14768);
and UO_805 (O_805,N_14377,N_14708);
and UO_806 (O_806,N_14280,N_14186);
nand UO_807 (O_807,N_14414,N_14946);
or UO_808 (O_808,N_14700,N_14607);
nor UO_809 (O_809,N_14293,N_14900);
nor UO_810 (O_810,N_14546,N_14272);
xor UO_811 (O_811,N_14918,N_14859);
xnor UO_812 (O_812,N_14252,N_14427);
or UO_813 (O_813,N_14466,N_14799);
xor UO_814 (O_814,N_14466,N_14227);
xor UO_815 (O_815,N_14171,N_14424);
nor UO_816 (O_816,N_14950,N_14590);
and UO_817 (O_817,N_14032,N_14084);
xor UO_818 (O_818,N_14744,N_14762);
nand UO_819 (O_819,N_14814,N_14390);
nand UO_820 (O_820,N_14214,N_14898);
and UO_821 (O_821,N_14628,N_14804);
nand UO_822 (O_822,N_14043,N_14453);
nand UO_823 (O_823,N_14973,N_14818);
xnor UO_824 (O_824,N_14212,N_14746);
and UO_825 (O_825,N_14971,N_14882);
xnor UO_826 (O_826,N_14179,N_14385);
or UO_827 (O_827,N_14125,N_14625);
xor UO_828 (O_828,N_14575,N_14774);
or UO_829 (O_829,N_14344,N_14500);
xor UO_830 (O_830,N_14489,N_14454);
and UO_831 (O_831,N_14902,N_14919);
xnor UO_832 (O_832,N_14210,N_14306);
xor UO_833 (O_833,N_14073,N_14636);
and UO_834 (O_834,N_14786,N_14751);
xor UO_835 (O_835,N_14280,N_14705);
nand UO_836 (O_836,N_14779,N_14545);
or UO_837 (O_837,N_14535,N_14178);
nand UO_838 (O_838,N_14697,N_14761);
nor UO_839 (O_839,N_14017,N_14267);
xnor UO_840 (O_840,N_14345,N_14686);
or UO_841 (O_841,N_14046,N_14756);
nor UO_842 (O_842,N_14651,N_14685);
and UO_843 (O_843,N_14073,N_14858);
nand UO_844 (O_844,N_14768,N_14720);
nand UO_845 (O_845,N_14234,N_14059);
nand UO_846 (O_846,N_14768,N_14341);
xor UO_847 (O_847,N_14663,N_14395);
xnor UO_848 (O_848,N_14868,N_14577);
or UO_849 (O_849,N_14509,N_14559);
and UO_850 (O_850,N_14392,N_14704);
xnor UO_851 (O_851,N_14186,N_14281);
nand UO_852 (O_852,N_14380,N_14532);
xor UO_853 (O_853,N_14166,N_14262);
nand UO_854 (O_854,N_14539,N_14155);
or UO_855 (O_855,N_14717,N_14481);
nand UO_856 (O_856,N_14026,N_14520);
xor UO_857 (O_857,N_14248,N_14426);
xnor UO_858 (O_858,N_14256,N_14082);
nor UO_859 (O_859,N_14721,N_14715);
xor UO_860 (O_860,N_14405,N_14193);
and UO_861 (O_861,N_14477,N_14527);
and UO_862 (O_862,N_14720,N_14029);
nor UO_863 (O_863,N_14692,N_14452);
and UO_864 (O_864,N_14328,N_14699);
nor UO_865 (O_865,N_14375,N_14764);
nand UO_866 (O_866,N_14531,N_14325);
or UO_867 (O_867,N_14415,N_14847);
xnor UO_868 (O_868,N_14156,N_14630);
xnor UO_869 (O_869,N_14212,N_14169);
nor UO_870 (O_870,N_14704,N_14393);
xnor UO_871 (O_871,N_14685,N_14749);
nand UO_872 (O_872,N_14129,N_14403);
and UO_873 (O_873,N_14256,N_14421);
nor UO_874 (O_874,N_14694,N_14639);
xnor UO_875 (O_875,N_14000,N_14692);
or UO_876 (O_876,N_14114,N_14413);
xnor UO_877 (O_877,N_14898,N_14217);
xor UO_878 (O_878,N_14471,N_14806);
or UO_879 (O_879,N_14017,N_14658);
or UO_880 (O_880,N_14737,N_14292);
nor UO_881 (O_881,N_14553,N_14409);
nand UO_882 (O_882,N_14452,N_14458);
nand UO_883 (O_883,N_14373,N_14232);
nor UO_884 (O_884,N_14154,N_14336);
or UO_885 (O_885,N_14123,N_14978);
and UO_886 (O_886,N_14997,N_14802);
xnor UO_887 (O_887,N_14852,N_14106);
or UO_888 (O_888,N_14067,N_14969);
and UO_889 (O_889,N_14071,N_14874);
xor UO_890 (O_890,N_14180,N_14346);
and UO_891 (O_891,N_14552,N_14997);
or UO_892 (O_892,N_14566,N_14971);
nand UO_893 (O_893,N_14138,N_14752);
xnor UO_894 (O_894,N_14924,N_14715);
nor UO_895 (O_895,N_14254,N_14361);
and UO_896 (O_896,N_14709,N_14283);
nor UO_897 (O_897,N_14823,N_14033);
xor UO_898 (O_898,N_14990,N_14041);
or UO_899 (O_899,N_14770,N_14663);
and UO_900 (O_900,N_14633,N_14347);
nor UO_901 (O_901,N_14625,N_14065);
and UO_902 (O_902,N_14277,N_14820);
xnor UO_903 (O_903,N_14146,N_14911);
nand UO_904 (O_904,N_14876,N_14976);
nor UO_905 (O_905,N_14064,N_14328);
or UO_906 (O_906,N_14104,N_14818);
nor UO_907 (O_907,N_14489,N_14886);
xor UO_908 (O_908,N_14486,N_14817);
nand UO_909 (O_909,N_14562,N_14274);
and UO_910 (O_910,N_14834,N_14562);
and UO_911 (O_911,N_14769,N_14316);
and UO_912 (O_912,N_14014,N_14737);
nand UO_913 (O_913,N_14465,N_14877);
nand UO_914 (O_914,N_14262,N_14586);
nand UO_915 (O_915,N_14900,N_14807);
or UO_916 (O_916,N_14426,N_14420);
or UO_917 (O_917,N_14396,N_14301);
or UO_918 (O_918,N_14394,N_14477);
nand UO_919 (O_919,N_14485,N_14337);
or UO_920 (O_920,N_14885,N_14671);
and UO_921 (O_921,N_14112,N_14570);
nor UO_922 (O_922,N_14119,N_14854);
nand UO_923 (O_923,N_14353,N_14319);
or UO_924 (O_924,N_14205,N_14897);
xnor UO_925 (O_925,N_14696,N_14148);
and UO_926 (O_926,N_14525,N_14605);
and UO_927 (O_927,N_14353,N_14762);
nor UO_928 (O_928,N_14686,N_14726);
and UO_929 (O_929,N_14707,N_14885);
and UO_930 (O_930,N_14554,N_14272);
nor UO_931 (O_931,N_14119,N_14337);
or UO_932 (O_932,N_14278,N_14476);
or UO_933 (O_933,N_14265,N_14931);
xnor UO_934 (O_934,N_14080,N_14804);
and UO_935 (O_935,N_14605,N_14106);
nor UO_936 (O_936,N_14451,N_14654);
nor UO_937 (O_937,N_14288,N_14644);
or UO_938 (O_938,N_14732,N_14777);
xor UO_939 (O_939,N_14016,N_14669);
and UO_940 (O_940,N_14985,N_14861);
and UO_941 (O_941,N_14687,N_14546);
or UO_942 (O_942,N_14673,N_14097);
and UO_943 (O_943,N_14870,N_14932);
nand UO_944 (O_944,N_14193,N_14111);
nand UO_945 (O_945,N_14688,N_14876);
xor UO_946 (O_946,N_14755,N_14057);
nor UO_947 (O_947,N_14833,N_14058);
nor UO_948 (O_948,N_14179,N_14766);
and UO_949 (O_949,N_14990,N_14560);
xnor UO_950 (O_950,N_14427,N_14223);
xnor UO_951 (O_951,N_14685,N_14735);
nor UO_952 (O_952,N_14247,N_14400);
nand UO_953 (O_953,N_14521,N_14164);
nand UO_954 (O_954,N_14602,N_14357);
xor UO_955 (O_955,N_14055,N_14799);
xor UO_956 (O_956,N_14207,N_14402);
and UO_957 (O_957,N_14659,N_14300);
nor UO_958 (O_958,N_14421,N_14099);
or UO_959 (O_959,N_14463,N_14130);
or UO_960 (O_960,N_14693,N_14731);
and UO_961 (O_961,N_14105,N_14887);
xnor UO_962 (O_962,N_14954,N_14722);
and UO_963 (O_963,N_14513,N_14516);
xnor UO_964 (O_964,N_14452,N_14132);
xor UO_965 (O_965,N_14322,N_14689);
nor UO_966 (O_966,N_14677,N_14906);
nor UO_967 (O_967,N_14076,N_14933);
xnor UO_968 (O_968,N_14397,N_14374);
and UO_969 (O_969,N_14392,N_14911);
and UO_970 (O_970,N_14653,N_14305);
or UO_971 (O_971,N_14318,N_14238);
and UO_972 (O_972,N_14771,N_14806);
nor UO_973 (O_973,N_14087,N_14504);
nand UO_974 (O_974,N_14052,N_14970);
and UO_975 (O_975,N_14308,N_14393);
nand UO_976 (O_976,N_14555,N_14360);
nand UO_977 (O_977,N_14195,N_14135);
or UO_978 (O_978,N_14329,N_14307);
and UO_979 (O_979,N_14860,N_14353);
xor UO_980 (O_980,N_14508,N_14916);
xnor UO_981 (O_981,N_14322,N_14024);
nor UO_982 (O_982,N_14472,N_14403);
xor UO_983 (O_983,N_14709,N_14868);
xnor UO_984 (O_984,N_14974,N_14897);
and UO_985 (O_985,N_14017,N_14699);
nand UO_986 (O_986,N_14070,N_14852);
nand UO_987 (O_987,N_14964,N_14973);
nor UO_988 (O_988,N_14188,N_14663);
nor UO_989 (O_989,N_14296,N_14417);
or UO_990 (O_990,N_14520,N_14586);
nor UO_991 (O_991,N_14467,N_14722);
nand UO_992 (O_992,N_14990,N_14292);
nand UO_993 (O_993,N_14575,N_14723);
or UO_994 (O_994,N_14303,N_14117);
xor UO_995 (O_995,N_14647,N_14061);
nor UO_996 (O_996,N_14083,N_14975);
and UO_997 (O_997,N_14370,N_14583);
or UO_998 (O_998,N_14831,N_14794);
and UO_999 (O_999,N_14578,N_14711);
nand UO_1000 (O_1000,N_14657,N_14798);
and UO_1001 (O_1001,N_14629,N_14111);
xor UO_1002 (O_1002,N_14236,N_14290);
nor UO_1003 (O_1003,N_14960,N_14937);
xor UO_1004 (O_1004,N_14393,N_14459);
nor UO_1005 (O_1005,N_14549,N_14572);
nand UO_1006 (O_1006,N_14293,N_14417);
and UO_1007 (O_1007,N_14292,N_14385);
xnor UO_1008 (O_1008,N_14710,N_14790);
nand UO_1009 (O_1009,N_14401,N_14000);
nor UO_1010 (O_1010,N_14815,N_14903);
or UO_1011 (O_1011,N_14648,N_14878);
nand UO_1012 (O_1012,N_14238,N_14234);
nor UO_1013 (O_1013,N_14645,N_14025);
nand UO_1014 (O_1014,N_14556,N_14756);
xor UO_1015 (O_1015,N_14740,N_14313);
or UO_1016 (O_1016,N_14242,N_14899);
nor UO_1017 (O_1017,N_14740,N_14412);
nor UO_1018 (O_1018,N_14352,N_14773);
nor UO_1019 (O_1019,N_14302,N_14669);
or UO_1020 (O_1020,N_14516,N_14028);
nor UO_1021 (O_1021,N_14489,N_14636);
xnor UO_1022 (O_1022,N_14084,N_14544);
and UO_1023 (O_1023,N_14103,N_14041);
or UO_1024 (O_1024,N_14609,N_14183);
nand UO_1025 (O_1025,N_14395,N_14088);
xnor UO_1026 (O_1026,N_14802,N_14429);
and UO_1027 (O_1027,N_14069,N_14496);
xor UO_1028 (O_1028,N_14514,N_14321);
or UO_1029 (O_1029,N_14296,N_14040);
and UO_1030 (O_1030,N_14249,N_14069);
and UO_1031 (O_1031,N_14326,N_14124);
xnor UO_1032 (O_1032,N_14306,N_14456);
xor UO_1033 (O_1033,N_14243,N_14832);
and UO_1034 (O_1034,N_14458,N_14934);
nand UO_1035 (O_1035,N_14465,N_14444);
xor UO_1036 (O_1036,N_14584,N_14555);
and UO_1037 (O_1037,N_14300,N_14408);
nand UO_1038 (O_1038,N_14045,N_14634);
nand UO_1039 (O_1039,N_14958,N_14439);
or UO_1040 (O_1040,N_14290,N_14985);
or UO_1041 (O_1041,N_14635,N_14054);
xnor UO_1042 (O_1042,N_14008,N_14481);
and UO_1043 (O_1043,N_14840,N_14581);
or UO_1044 (O_1044,N_14571,N_14446);
xnor UO_1045 (O_1045,N_14585,N_14896);
nor UO_1046 (O_1046,N_14132,N_14914);
and UO_1047 (O_1047,N_14600,N_14040);
nor UO_1048 (O_1048,N_14047,N_14572);
and UO_1049 (O_1049,N_14127,N_14543);
xor UO_1050 (O_1050,N_14459,N_14050);
xor UO_1051 (O_1051,N_14224,N_14454);
and UO_1052 (O_1052,N_14723,N_14324);
or UO_1053 (O_1053,N_14737,N_14062);
nand UO_1054 (O_1054,N_14605,N_14880);
nand UO_1055 (O_1055,N_14473,N_14518);
nand UO_1056 (O_1056,N_14940,N_14133);
and UO_1057 (O_1057,N_14256,N_14027);
xnor UO_1058 (O_1058,N_14314,N_14024);
xor UO_1059 (O_1059,N_14213,N_14320);
nor UO_1060 (O_1060,N_14759,N_14271);
xnor UO_1061 (O_1061,N_14265,N_14788);
nor UO_1062 (O_1062,N_14616,N_14713);
and UO_1063 (O_1063,N_14073,N_14543);
nand UO_1064 (O_1064,N_14683,N_14294);
nor UO_1065 (O_1065,N_14064,N_14856);
nand UO_1066 (O_1066,N_14090,N_14222);
nor UO_1067 (O_1067,N_14089,N_14653);
and UO_1068 (O_1068,N_14102,N_14248);
nand UO_1069 (O_1069,N_14268,N_14509);
nor UO_1070 (O_1070,N_14959,N_14000);
xor UO_1071 (O_1071,N_14707,N_14307);
and UO_1072 (O_1072,N_14912,N_14158);
or UO_1073 (O_1073,N_14020,N_14841);
or UO_1074 (O_1074,N_14689,N_14519);
nand UO_1075 (O_1075,N_14450,N_14333);
or UO_1076 (O_1076,N_14190,N_14069);
and UO_1077 (O_1077,N_14164,N_14182);
and UO_1078 (O_1078,N_14876,N_14566);
xor UO_1079 (O_1079,N_14928,N_14663);
nand UO_1080 (O_1080,N_14325,N_14043);
and UO_1081 (O_1081,N_14435,N_14228);
nand UO_1082 (O_1082,N_14348,N_14743);
xor UO_1083 (O_1083,N_14190,N_14182);
and UO_1084 (O_1084,N_14415,N_14908);
or UO_1085 (O_1085,N_14129,N_14611);
nand UO_1086 (O_1086,N_14566,N_14934);
and UO_1087 (O_1087,N_14079,N_14334);
and UO_1088 (O_1088,N_14258,N_14025);
nand UO_1089 (O_1089,N_14331,N_14677);
nor UO_1090 (O_1090,N_14410,N_14088);
and UO_1091 (O_1091,N_14374,N_14608);
nand UO_1092 (O_1092,N_14572,N_14725);
nand UO_1093 (O_1093,N_14925,N_14891);
and UO_1094 (O_1094,N_14963,N_14677);
xnor UO_1095 (O_1095,N_14370,N_14485);
nor UO_1096 (O_1096,N_14519,N_14473);
nor UO_1097 (O_1097,N_14025,N_14328);
and UO_1098 (O_1098,N_14208,N_14091);
nand UO_1099 (O_1099,N_14709,N_14944);
or UO_1100 (O_1100,N_14662,N_14555);
xor UO_1101 (O_1101,N_14637,N_14725);
nor UO_1102 (O_1102,N_14762,N_14477);
xor UO_1103 (O_1103,N_14209,N_14438);
nand UO_1104 (O_1104,N_14413,N_14637);
or UO_1105 (O_1105,N_14355,N_14601);
nand UO_1106 (O_1106,N_14457,N_14106);
or UO_1107 (O_1107,N_14479,N_14400);
xor UO_1108 (O_1108,N_14304,N_14534);
or UO_1109 (O_1109,N_14743,N_14071);
xor UO_1110 (O_1110,N_14658,N_14407);
or UO_1111 (O_1111,N_14665,N_14617);
nand UO_1112 (O_1112,N_14127,N_14871);
nor UO_1113 (O_1113,N_14364,N_14356);
xor UO_1114 (O_1114,N_14408,N_14600);
nor UO_1115 (O_1115,N_14042,N_14207);
xor UO_1116 (O_1116,N_14386,N_14677);
nor UO_1117 (O_1117,N_14024,N_14849);
and UO_1118 (O_1118,N_14712,N_14531);
or UO_1119 (O_1119,N_14511,N_14539);
nand UO_1120 (O_1120,N_14919,N_14041);
nand UO_1121 (O_1121,N_14493,N_14471);
nand UO_1122 (O_1122,N_14278,N_14721);
nand UO_1123 (O_1123,N_14581,N_14087);
xor UO_1124 (O_1124,N_14144,N_14405);
nor UO_1125 (O_1125,N_14846,N_14315);
and UO_1126 (O_1126,N_14051,N_14700);
nand UO_1127 (O_1127,N_14771,N_14951);
or UO_1128 (O_1128,N_14596,N_14778);
or UO_1129 (O_1129,N_14544,N_14153);
and UO_1130 (O_1130,N_14234,N_14334);
nand UO_1131 (O_1131,N_14231,N_14058);
nor UO_1132 (O_1132,N_14332,N_14126);
and UO_1133 (O_1133,N_14206,N_14720);
xor UO_1134 (O_1134,N_14527,N_14019);
nand UO_1135 (O_1135,N_14088,N_14906);
nor UO_1136 (O_1136,N_14122,N_14156);
nand UO_1137 (O_1137,N_14223,N_14888);
or UO_1138 (O_1138,N_14505,N_14519);
and UO_1139 (O_1139,N_14938,N_14419);
or UO_1140 (O_1140,N_14650,N_14841);
nor UO_1141 (O_1141,N_14003,N_14719);
or UO_1142 (O_1142,N_14223,N_14984);
nor UO_1143 (O_1143,N_14871,N_14704);
or UO_1144 (O_1144,N_14493,N_14796);
and UO_1145 (O_1145,N_14812,N_14071);
nor UO_1146 (O_1146,N_14668,N_14842);
nand UO_1147 (O_1147,N_14943,N_14581);
xor UO_1148 (O_1148,N_14870,N_14010);
xor UO_1149 (O_1149,N_14518,N_14261);
xnor UO_1150 (O_1150,N_14435,N_14727);
or UO_1151 (O_1151,N_14606,N_14330);
or UO_1152 (O_1152,N_14638,N_14342);
or UO_1153 (O_1153,N_14636,N_14643);
nand UO_1154 (O_1154,N_14596,N_14510);
or UO_1155 (O_1155,N_14553,N_14273);
nand UO_1156 (O_1156,N_14605,N_14133);
nor UO_1157 (O_1157,N_14871,N_14110);
nor UO_1158 (O_1158,N_14339,N_14565);
nor UO_1159 (O_1159,N_14735,N_14967);
xor UO_1160 (O_1160,N_14345,N_14661);
xor UO_1161 (O_1161,N_14198,N_14544);
nand UO_1162 (O_1162,N_14840,N_14794);
xnor UO_1163 (O_1163,N_14080,N_14886);
xor UO_1164 (O_1164,N_14434,N_14300);
and UO_1165 (O_1165,N_14544,N_14471);
and UO_1166 (O_1166,N_14501,N_14795);
or UO_1167 (O_1167,N_14765,N_14112);
xor UO_1168 (O_1168,N_14620,N_14344);
nand UO_1169 (O_1169,N_14793,N_14925);
xnor UO_1170 (O_1170,N_14280,N_14706);
or UO_1171 (O_1171,N_14298,N_14774);
xor UO_1172 (O_1172,N_14437,N_14521);
and UO_1173 (O_1173,N_14844,N_14338);
nor UO_1174 (O_1174,N_14735,N_14942);
or UO_1175 (O_1175,N_14862,N_14115);
nand UO_1176 (O_1176,N_14077,N_14638);
and UO_1177 (O_1177,N_14727,N_14362);
and UO_1178 (O_1178,N_14590,N_14025);
or UO_1179 (O_1179,N_14450,N_14097);
nor UO_1180 (O_1180,N_14938,N_14429);
nand UO_1181 (O_1181,N_14282,N_14680);
nor UO_1182 (O_1182,N_14013,N_14685);
or UO_1183 (O_1183,N_14692,N_14546);
and UO_1184 (O_1184,N_14874,N_14009);
and UO_1185 (O_1185,N_14331,N_14597);
and UO_1186 (O_1186,N_14786,N_14424);
xor UO_1187 (O_1187,N_14558,N_14089);
nor UO_1188 (O_1188,N_14533,N_14001);
nand UO_1189 (O_1189,N_14712,N_14071);
nand UO_1190 (O_1190,N_14573,N_14833);
xor UO_1191 (O_1191,N_14251,N_14375);
xor UO_1192 (O_1192,N_14251,N_14118);
and UO_1193 (O_1193,N_14897,N_14598);
nand UO_1194 (O_1194,N_14720,N_14686);
nand UO_1195 (O_1195,N_14193,N_14574);
or UO_1196 (O_1196,N_14991,N_14177);
nand UO_1197 (O_1197,N_14523,N_14861);
xor UO_1198 (O_1198,N_14947,N_14188);
nor UO_1199 (O_1199,N_14931,N_14715);
nand UO_1200 (O_1200,N_14138,N_14301);
and UO_1201 (O_1201,N_14245,N_14596);
nand UO_1202 (O_1202,N_14537,N_14297);
and UO_1203 (O_1203,N_14190,N_14640);
nand UO_1204 (O_1204,N_14479,N_14374);
nand UO_1205 (O_1205,N_14816,N_14491);
xor UO_1206 (O_1206,N_14543,N_14548);
nor UO_1207 (O_1207,N_14436,N_14034);
xor UO_1208 (O_1208,N_14890,N_14052);
and UO_1209 (O_1209,N_14077,N_14218);
nand UO_1210 (O_1210,N_14895,N_14062);
nand UO_1211 (O_1211,N_14119,N_14445);
nand UO_1212 (O_1212,N_14117,N_14724);
and UO_1213 (O_1213,N_14391,N_14233);
or UO_1214 (O_1214,N_14529,N_14778);
xor UO_1215 (O_1215,N_14368,N_14325);
nand UO_1216 (O_1216,N_14972,N_14420);
or UO_1217 (O_1217,N_14255,N_14864);
nand UO_1218 (O_1218,N_14377,N_14960);
nand UO_1219 (O_1219,N_14030,N_14587);
and UO_1220 (O_1220,N_14646,N_14111);
nor UO_1221 (O_1221,N_14498,N_14172);
and UO_1222 (O_1222,N_14965,N_14056);
nor UO_1223 (O_1223,N_14677,N_14801);
or UO_1224 (O_1224,N_14351,N_14501);
or UO_1225 (O_1225,N_14295,N_14841);
xnor UO_1226 (O_1226,N_14393,N_14487);
nor UO_1227 (O_1227,N_14456,N_14147);
nor UO_1228 (O_1228,N_14950,N_14610);
and UO_1229 (O_1229,N_14443,N_14420);
nand UO_1230 (O_1230,N_14296,N_14393);
and UO_1231 (O_1231,N_14576,N_14474);
xor UO_1232 (O_1232,N_14076,N_14104);
xor UO_1233 (O_1233,N_14987,N_14002);
xor UO_1234 (O_1234,N_14654,N_14939);
xor UO_1235 (O_1235,N_14112,N_14044);
xor UO_1236 (O_1236,N_14176,N_14248);
nor UO_1237 (O_1237,N_14388,N_14224);
and UO_1238 (O_1238,N_14384,N_14916);
and UO_1239 (O_1239,N_14293,N_14720);
nand UO_1240 (O_1240,N_14213,N_14702);
nor UO_1241 (O_1241,N_14698,N_14526);
or UO_1242 (O_1242,N_14169,N_14072);
or UO_1243 (O_1243,N_14395,N_14839);
and UO_1244 (O_1244,N_14329,N_14848);
xnor UO_1245 (O_1245,N_14074,N_14578);
xnor UO_1246 (O_1246,N_14565,N_14367);
nor UO_1247 (O_1247,N_14441,N_14889);
nand UO_1248 (O_1248,N_14207,N_14381);
or UO_1249 (O_1249,N_14152,N_14912);
and UO_1250 (O_1250,N_14999,N_14751);
or UO_1251 (O_1251,N_14444,N_14675);
or UO_1252 (O_1252,N_14607,N_14655);
and UO_1253 (O_1253,N_14357,N_14089);
or UO_1254 (O_1254,N_14425,N_14501);
and UO_1255 (O_1255,N_14970,N_14458);
or UO_1256 (O_1256,N_14115,N_14189);
nor UO_1257 (O_1257,N_14880,N_14422);
and UO_1258 (O_1258,N_14279,N_14482);
nor UO_1259 (O_1259,N_14246,N_14880);
and UO_1260 (O_1260,N_14235,N_14033);
or UO_1261 (O_1261,N_14690,N_14878);
nand UO_1262 (O_1262,N_14771,N_14501);
or UO_1263 (O_1263,N_14720,N_14169);
and UO_1264 (O_1264,N_14960,N_14654);
nor UO_1265 (O_1265,N_14954,N_14431);
or UO_1266 (O_1266,N_14041,N_14525);
nand UO_1267 (O_1267,N_14583,N_14294);
and UO_1268 (O_1268,N_14302,N_14820);
or UO_1269 (O_1269,N_14492,N_14255);
nor UO_1270 (O_1270,N_14891,N_14348);
nor UO_1271 (O_1271,N_14229,N_14391);
and UO_1272 (O_1272,N_14501,N_14390);
nor UO_1273 (O_1273,N_14688,N_14434);
nor UO_1274 (O_1274,N_14701,N_14054);
xnor UO_1275 (O_1275,N_14876,N_14831);
xnor UO_1276 (O_1276,N_14587,N_14590);
xor UO_1277 (O_1277,N_14850,N_14593);
nor UO_1278 (O_1278,N_14377,N_14154);
nor UO_1279 (O_1279,N_14425,N_14034);
nor UO_1280 (O_1280,N_14376,N_14938);
nand UO_1281 (O_1281,N_14150,N_14689);
and UO_1282 (O_1282,N_14901,N_14709);
or UO_1283 (O_1283,N_14559,N_14823);
and UO_1284 (O_1284,N_14499,N_14180);
and UO_1285 (O_1285,N_14674,N_14427);
nand UO_1286 (O_1286,N_14271,N_14895);
nor UO_1287 (O_1287,N_14013,N_14230);
and UO_1288 (O_1288,N_14041,N_14032);
nand UO_1289 (O_1289,N_14299,N_14259);
and UO_1290 (O_1290,N_14152,N_14842);
nor UO_1291 (O_1291,N_14027,N_14383);
or UO_1292 (O_1292,N_14458,N_14640);
nor UO_1293 (O_1293,N_14236,N_14132);
or UO_1294 (O_1294,N_14158,N_14636);
nor UO_1295 (O_1295,N_14452,N_14000);
and UO_1296 (O_1296,N_14735,N_14283);
nand UO_1297 (O_1297,N_14020,N_14021);
nand UO_1298 (O_1298,N_14462,N_14636);
or UO_1299 (O_1299,N_14352,N_14992);
and UO_1300 (O_1300,N_14623,N_14140);
nand UO_1301 (O_1301,N_14291,N_14659);
or UO_1302 (O_1302,N_14831,N_14941);
xnor UO_1303 (O_1303,N_14174,N_14990);
nor UO_1304 (O_1304,N_14117,N_14384);
xor UO_1305 (O_1305,N_14821,N_14658);
and UO_1306 (O_1306,N_14595,N_14212);
nor UO_1307 (O_1307,N_14703,N_14939);
and UO_1308 (O_1308,N_14397,N_14915);
nor UO_1309 (O_1309,N_14796,N_14844);
and UO_1310 (O_1310,N_14904,N_14588);
nor UO_1311 (O_1311,N_14141,N_14383);
nor UO_1312 (O_1312,N_14561,N_14839);
nor UO_1313 (O_1313,N_14406,N_14431);
xor UO_1314 (O_1314,N_14599,N_14494);
or UO_1315 (O_1315,N_14317,N_14272);
xor UO_1316 (O_1316,N_14780,N_14209);
nor UO_1317 (O_1317,N_14736,N_14518);
and UO_1318 (O_1318,N_14019,N_14035);
nor UO_1319 (O_1319,N_14082,N_14321);
and UO_1320 (O_1320,N_14525,N_14176);
or UO_1321 (O_1321,N_14180,N_14697);
or UO_1322 (O_1322,N_14458,N_14463);
nor UO_1323 (O_1323,N_14467,N_14569);
or UO_1324 (O_1324,N_14286,N_14983);
xnor UO_1325 (O_1325,N_14586,N_14574);
xnor UO_1326 (O_1326,N_14274,N_14532);
xnor UO_1327 (O_1327,N_14638,N_14741);
nor UO_1328 (O_1328,N_14220,N_14288);
nand UO_1329 (O_1329,N_14513,N_14602);
xnor UO_1330 (O_1330,N_14235,N_14322);
or UO_1331 (O_1331,N_14892,N_14543);
or UO_1332 (O_1332,N_14133,N_14834);
nand UO_1333 (O_1333,N_14628,N_14909);
and UO_1334 (O_1334,N_14293,N_14975);
xor UO_1335 (O_1335,N_14812,N_14092);
xor UO_1336 (O_1336,N_14545,N_14110);
and UO_1337 (O_1337,N_14663,N_14955);
nand UO_1338 (O_1338,N_14511,N_14802);
and UO_1339 (O_1339,N_14277,N_14430);
nand UO_1340 (O_1340,N_14496,N_14644);
nor UO_1341 (O_1341,N_14573,N_14230);
nand UO_1342 (O_1342,N_14720,N_14280);
xor UO_1343 (O_1343,N_14125,N_14180);
and UO_1344 (O_1344,N_14650,N_14451);
nand UO_1345 (O_1345,N_14383,N_14733);
nor UO_1346 (O_1346,N_14520,N_14606);
nand UO_1347 (O_1347,N_14087,N_14110);
nand UO_1348 (O_1348,N_14881,N_14738);
and UO_1349 (O_1349,N_14141,N_14453);
nor UO_1350 (O_1350,N_14706,N_14545);
or UO_1351 (O_1351,N_14418,N_14316);
nor UO_1352 (O_1352,N_14245,N_14339);
and UO_1353 (O_1353,N_14736,N_14166);
nor UO_1354 (O_1354,N_14915,N_14362);
xnor UO_1355 (O_1355,N_14397,N_14089);
or UO_1356 (O_1356,N_14806,N_14938);
or UO_1357 (O_1357,N_14818,N_14802);
nor UO_1358 (O_1358,N_14824,N_14498);
nand UO_1359 (O_1359,N_14652,N_14985);
nand UO_1360 (O_1360,N_14254,N_14989);
or UO_1361 (O_1361,N_14076,N_14855);
or UO_1362 (O_1362,N_14545,N_14036);
or UO_1363 (O_1363,N_14293,N_14132);
or UO_1364 (O_1364,N_14940,N_14272);
or UO_1365 (O_1365,N_14685,N_14850);
nor UO_1366 (O_1366,N_14115,N_14238);
nor UO_1367 (O_1367,N_14250,N_14707);
xnor UO_1368 (O_1368,N_14586,N_14558);
xnor UO_1369 (O_1369,N_14635,N_14265);
xor UO_1370 (O_1370,N_14599,N_14326);
nand UO_1371 (O_1371,N_14786,N_14760);
nand UO_1372 (O_1372,N_14665,N_14935);
and UO_1373 (O_1373,N_14214,N_14259);
and UO_1374 (O_1374,N_14839,N_14797);
and UO_1375 (O_1375,N_14069,N_14707);
nor UO_1376 (O_1376,N_14608,N_14143);
and UO_1377 (O_1377,N_14643,N_14929);
xor UO_1378 (O_1378,N_14093,N_14144);
and UO_1379 (O_1379,N_14171,N_14318);
and UO_1380 (O_1380,N_14443,N_14291);
and UO_1381 (O_1381,N_14764,N_14558);
and UO_1382 (O_1382,N_14257,N_14848);
and UO_1383 (O_1383,N_14231,N_14263);
nand UO_1384 (O_1384,N_14034,N_14484);
xnor UO_1385 (O_1385,N_14694,N_14042);
xnor UO_1386 (O_1386,N_14237,N_14029);
nor UO_1387 (O_1387,N_14425,N_14303);
and UO_1388 (O_1388,N_14494,N_14193);
xnor UO_1389 (O_1389,N_14585,N_14364);
and UO_1390 (O_1390,N_14757,N_14980);
or UO_1391 (O_1391,N_14006,N_14263);
xnor UO_1392 (O_1392,N_14688,N_14804);
xor UO_1393 (O_1393,N_14785,N_14983);
xor UO_1394 (O_1394,N_14235,N_14777);
nand UO_1395 (O_1395,N_14022,N_14467);
nor UO_1396 (O_1396,N_14923,N_14382);
or UO_1397 (O_1397,N_14234,N_14451);
xor UO_1398 (O_1398,N_14803,N_14273);
nor UO_1399 (O_1399,N_14948,N_14215);
or UO_1400 (O_1400,N_14613,N_14615);
nor UO_1401 (O_1401,N_14811,N_14295);
and UO_1402 (O_1402,N_14292,N_14298);
nor UO_1403 (O_1403,N_14053,N_14220);
or UO_1404 (O_1404,N_14568,N_14696);
and UO_1405 (O_1405,N_14671,N_14553);
or UO_1406 (O_1406,N_14692,N_14977);
nand UO_1407 (O_1407,N_14279,N_14427);
and UO_1408 (O_1408,N_14670,N_14980);
nand UO_1409 (O_1409,N_14847,N_14016);
xnor UO_1410 (O_1410,N_14278,N_14648);
or UO_1411 (O_1411,N_14665,N_14041);
nand UO_1412 (O_1412,N_14836,N_14762);
xor UO_1413 (O_1413,N_14360,N_14056);
xnor UO_1414 (O_1414,N_14879,N_14894);
and UO_1415 (O_1415,N_14064,N_14760);
nor UO_1416 (O_1416,N_14211,N_14523);
xor UO_1417 (O_1417,N_14072,N_14533);
xnor UO_1418 (O_1418,N_14663,N_14925);
nor UO_1419 (O_1419,N_14931,N_14378);
nor UO_1420 (O_1420,N_14406,N_14759);
and UO_1421 (O_1421,N_14839,N_14485);
nand UO_1422 (O_1422,N_14166,N_14861);
and UO_1423 (O_1423,N_14842,N_14627);
or UO_1424 (O_1424,N_14765,N_14733);
or UO_1425 (O_1425,N_14177,N_14191);
nand UO_1426 (O_1426,N_14723,N_14152);
and UO_1427 (O_1427,N_14920,N_14701);
or UO_1428 (O_1428,N_14529,N_14909);
nand UO_1429 (O_1429,N_14657,N_14190);
nor UO_1430 (O_1430,N_14471,N_14047);
nor UO_1431 (O_1431,N_14520,N_14142);
xnor UO_1432 (O_1432,N_14432,N_14798);
nand UO_1433 (O_1433,N_14602,N_14773);
and UO_1434 (O_1434,N_14117,N_14810);
and UO_1435 (O_1435,N_14166,N_14445);
xor UO_1436 (O_1436,N_14720,N_14104);
nor UO_1437 (O_1437,N_14790,N_14638);
or UO_1438 (O_1438,N_14236,N_14972);
xnor UO_1439 (O_1439,N_14351,N_14673);
and UO_1440 (O_1440,N_14910,N_14773);
or UO_1441 (O_1441,N_14686,N_14234);
nand UO_1442 (O_1442,N_14554,N_14482);
nor UO_1443 (O_1443,N_14678,N_14777);
xnor UO_1444 (O_1444,N_14090,N_14710);
and UO_1445 (O_1445,N_14481,N_14117);
and UO_1446 (O_1446,N_14654,N_14560);
nand UO_1447 (O_1447,N_14956,N_14626);
and UO_1448 (O_1448,N_14593,N_14488);
nand UO_1449 (O_1449,N_14383,N_14098);
nand UO_1450 (O_1450,N_14762,N_14561);
and UO_1451 (O_1451,N_14505,N_14467);
or UO_1452 (O_1452,N_14371,N_14013);
xnor UO_1453 (O_1453,N_14322,N_14388);
nand UO_1454 (O_1454,N_14022,N_14237);
and UO_1455 (O_1455,N_14689,N_14497);
and UO_1456 (O_1456,N_14631,N_14922);
nand UO_1457 (O_1457,N_14825,N_14937);
or UO_1458 (O_1458,N_14467,N_14261);
nand UO_1459 (O_1459,N_14825,N_14698);
or UO_1460 (O_1460,N_14308,N_14753);
nand UO_1461 (O_1461,N_14730,N_14589);
and UO_1462 (O_1462,N_14657,N_14632);
xnor UO_1463 (O_1463,N_14377,N_14886);
nor UO_1464 (O_1464,N_14697,N_14832);
or UO_1465 (O_1465,N_14251,N_14128);
xor UO_1466 (O_1466,N_14704,N_14772);
xnor UO_1467 (O_1467,N_14810,N_14349);
nor UO_1468 (O_1468,N_14366,N_14617);
or UO_1469 (O_1469,N_14913,N_14296);
nor UO_1470 (O_1470,N_14261,N_14291);
or UO_1471 (O_1471,N_14286,N_14183);
nor UO_1472 (O_1472,N_14150,N_14854);
and UO_1473 (O_1473,N_14848,N_14865);
nand UO_1474 (O_1474,N_14241,N_14200);
nand UO_1475 (O_1475,N_14020,N_14948);
xnor UO_1476 (O_1476,N_14774,N_14822);
xor UO_1477 (O_1477,N_14417,N_14537);
xor UO_1478 (O_1478,N_14950,N_14744);
and UO_1479 (O_1479,N_14263,N_14887);
nand UO_1480 (O_1480,N_14967,N_14845);
or UO_1481 (O_1481,N_14189,N_14623);
and UO_1482 (O_1482,N_14602,N_14543);
nand UO_1483 (O_1483,N_14352,N_14517);
or UO_1484 (O_1484,N_14746,N_14978);
nor UO_1485 (O_1485,N_14886,N_14851);
xnor UO_1486 (O_1486,N_14691,N_14211);
and UO_1487 (O_1487,N_14094,N_14770);
nand UO_1488 (O_1488,N_14453,N_14765);
xor UO_1489 (O_1489,N_14331,N_14400);
and UO_1490 (O_1490,N_14695,N_14843);
nand UO_1491 (O_1491,N_14925,N_14349);
xor UO_1492 (O_1492,N_14453,N_14158);
xnor UO_1493 (O_1493,N_14677,N_14413);
or UO_1494 (O_1494,N_14614,N_14628);
and UO_1495 (O_1495,N_14656,N_14253);
or UO_1496 (O_1496,N_14212,N_14315);
xnor UO_1497 (O_1497,N_14221,N_14800);
or UO_1498 (O_1498,N_14571,N_14012);
and UO_1499 (O_1499,N_14632,N_14863);
nand UO_1500 (O_1500,N_14890,N_14717);
or UO_1501 (O_1501,N_14512,N_14596);
xnor UO_1502 (O_1502,N_14544,N_14831);
xnor UO_1503 (O_1503,N_14798,N_14713);
nand UO_1504 (O_1504,N_14545,N_14626);
or UO_1505 (O_1505,N_14195,N_14011);
or UO_1506 (O_1506,N_14263,N_14189);
or UO_1507 (O_1507,N_14653,N_14002);
and UO_1508 (O_1508,N_14069,N_14752);
and UO_1509 (O_1509,N_14798,N_14146);
nand UO_1510 (O_1510,N_14736,N_14657);
xnor UO_1511 (O_1511,N_14899,N_14764);
xor UO_1512 (O_1512,N_14411,N_14508);
and UO_1513 (O_1513,N_14723,N_14807);
nor UO_1514 (O_1514,N_14599,N_14545);
or UO_1515 (O_1515,N_14007,N_14834);
xor UO_1516 (O_1516,N_14883,N_14498);
nor UO_1517 (O_1517,N_14089,N_14031);
nand UO_1518 (O_1518,N_14697,N_14895);
or UO_1519 (O_1519,N_14463,N_14117);
xnor UO_1520 (O_1520,N_14938,N_14271);
nand UO_1521 (O_1521,N_14109,N_14715);
nor UO_1522 (O_1522,N_14918,N_14503);
and UO_1523 (O_1523,N_14449,N_14802);
nor UO_1524 (O_1524,N_14252,N_14138);
xnor UO_1525 (O_1525,N_14130,N_14828);
nand UO_1526 (O_1526,N_14837,N_14589);
or UO_1527 (O_1527,N_14376,N_14255);
or UO_1528 (O_1528,N_14053,N_14694);
and UO_1529 (O_1529,N_14657,N_14064);
and UO_1530 (O_1530,N_14943,N_14075);
nor UO_1531 (O_1531,N_14414,N_14715);
nor UO_1532 (O_1532,N_14616,N_14775);
nor UO_1533 (O_1533,N_14233,N_14444);
nor UO_1534 (O_1534,N_14722,N_14113);
nor UO_1535 (O_1535,N_14958,N_14087);
or UO_1536 (O_1536,N_14260,N_14888);
and UO_1537 (O_1537,N_14457,N_14283);
nand UO_1538 (O_1538,N_14738,N_14089);
nand UO_1539 (O_1539,N_14555,N_14980);
or UO_1540 (O_1540,N_14877,N_14616);
xor UO_1541 (O_1541,N_14276,N_14787);
xnor UO_1542 (O_1542,N_14791,N_14002);
nand UO_1543 (O_1543,N_14471,N_14574);
or UO_1544 (O_1544,N_14820,N_14765);
nand UO_1545 (O_1545,N_14492,N_14849);
xnor UO_1546 (O_1546,N_14950,N_14455);
and UO_1547 (O_1547,N_14529,N_14267);
nor UO_1548 (O_1548,N_14015,N_14309);
nand UO_1549 (O_1549,N_14331,N_14021);
xnor UO_1550 (O_1550,N_14426,N_14799);
nor UO_1551 (O_1551,N_14131,N_14955);
nor UO_1552 (O_1552,N_14910,N_14261);
and UO_1553 (O_1553,N_14579,N_14281);
nor UO_1554 (O_1554,N_14891,N_14369);
or UO_1555 (O_1555,N_14412,N_14397);
or UO_1556 (O_1556,N_14493,N_14461);
nor UO_1557 (O_1557,N_14310,N_14164);
and UO_1558 (O_1558,N_14444,N_14018);
nand UO_1559 (O_1559,N_14730,N_14300);
and UO_1560 (O_1560,N_14920,N_14856);
xnor UO_1561 (O_1561,N_14318,N_14236);
nor UO_1562 (O_1562,N_14301,N_14482);
xnor UO_1563 (O_1563,N_14521,N_14927);
xor UO_1564 (O_1564,N_14747,N_14928);
and UO_1565 (O_1565,N_14104,N_14742);
xnor UO_1566 (O_1566,N_14811,N_14837);
xnor UO_1567 (O_1567,N_14583,N_14111);
xor UO_1568 (O_1568,N_14050,N_14544);
and UO_1569 (O_1569,N_14080,N_14862);
nand UO_1570 (O_1570,N_14062,N_14441);
nor UO_1571 (O_1571,N_14774,N_14622);
or UO_1572 (O_1572,N_14690,N_14749);
or UO_1573 (O_1573,N_14811,N_14197);
xor UO_1574 (O_1574,N_14545,N_14471);
nand UO_1575 (O_1575,N_14152,N_14374);
nor UO_1576 (O_1576,N_14818,N_14820);
xnor UO_1577 (O_1577,N_14943,N_14870);
and UO_1578 (O_1578,N_14281,N_14934);
or UO_1579 (O_1579,N_14057,N_14199);
xor UO_1580 (O_1580,N_14408,N_14071);
and UO_1581 (O_1581,N_14634,N_14005);
nor UO_1582 (O_1582,N_14409,N_14618);
or UO_1583 (O_1583,N_14044,N_14385);
or UO_1584 (O_1584,N_14910,N_14937);
nor UO_1585 (O_1585,N_14609,N_14055);
or UO_1586 (O_1586,N_14675,N_14322);
and UO_1587 (O_1587,N_14180,N_14751);
xor UO_1588 (O_1588,N_14491,N_14548);
and UO_1589 (O_1589,N_14133,N_14522);
or UO_1590 (O_1590,N_14763,N_14053);
xnor UO_1591 (O_1591,N_14229,N_14175);
xnor UO_1592 (O_1592,N_14186,N_14745);
xor UO_1593 (O_1593,N_14158,N_14916);
or UO_1594 (O_1594,N_14593,N_14361);
nor UO_1595 (O_1595,N_14093,N_14781);
or UO_1596 (O_1596,N_14683,N_14263);
and UO_1597 (O_1597,N_14988,N_14963);
and UO_1598 (O_1598,N_14392,N_14159);
and UO_1599 (O_1599,N_14768,N_14417);
or UO_1600 (O_1600,N_14324,N_14979);
xor UO_1601 (O_1601,N_14281,N_14018);
or UO_1602 (O_1602,N_14408,N_14526);
or UO_1603 (O_1603,N_14428,N_14399);
xnor UO_1604 (O_1604,N_14293,N_14151);
xnor UO_1605 (O_1605,N_14934,N_14709);
and UO_1606 (O_1606,N_14220,N_14708);
nor UO_1607 (O_1607,N_14671,N_14392);
nand UO_1608 (O_1608,N_14743,N_14666);
and UO_1609 (O_1609,N_14671,N_14415);
or UO_1610 (O_1610,N_14176,N_14047);
or UO_1611 (O_1611,N_14564,N_14952);
nor UO_1612 (O_1612,N_14295,N_14244);
and UO_1613 (O_1613,N_14049,N_14089);
nor UO_1614 (O_1614,N_14743,N_14316);
or UO_1615 (O_1615,N_14971,N_14806);
nand UO_1616 (O_1616,N_14396,N_14496);
nor UO_1617 (O_1617,N_14200,N_14457);
xor UO_1618 (O_1618,N_14030,N_14854);
xnor UO_1619 (O_1619,N_14346,N_14197);
and UO_1620 (O_1620,N_14276,N_14966);
xnor UO_1621 (O_1621,N_14437,N_14331);
and UO_1622 (O_1622,N_14026,N_14174);
or UO_1623 (O_1623,N_14594,N_14116);
nand UO_1624 (O_1624,N_14414,N_14693);
or UO_1625 (O_1625,N_14251,N_14232);
or UO_1626 (O_1626,N_14449,N_14768);
or UO_1627 (O_1627,N_14047,N_14326);
xnor UO_1628 (O_1628,N_14071,N_14055);
nand UO_1629 (O_1629,N_14092,N_14950);
or UO_1630 (O_1630,N_14046,N_14614);
or UO_1631 (O_1631,N_14688,N_14614);
and UO_1632 (O_1632,N_14138,N_14764);
and UO_1633 (O_1633,N_14650,N_14470);
nand UO_1634 (O_1634,N_14937,N_14676);
nor UO_1635 (O_1635,N_14964,N_14373);
and UO_1636 (O_1636,N_14032,N_14219);
and UO_1637 (O_1637,N_14836,N_14764);
or UO_1638 (O_1638,N_14639,N_14823);
nor UO_1639 (O_1639,N_14482,N_14404);
nor UO_1640 (O_1640,N_14661,N_14547);
and UO_1641 (O_1641,N_14278,N_14083);
nand UO_1642 (O_1642,N_14733,N_14717);
and UO_1643 (O_1643,N_14896,N_14860);
and UO_1644 (O_1644,N_14556,N_14389);
or UO_1645 (O_1645,N_14360,N_14240);
nand UO_1646 (O_1646,N_14299,N_14264);
nor UO_1647 (O_1647,N_14694,N_14499);
nand UO_1648 (O_1648,N_14685,N_14345);
xnor UO_1649 (O_1649,N_14075,N_14370);
nand UO_1650 (O_1650,N_14047,N_14667);
xnor UO_1651 (O_1651,N_14928,N_14315);
or UO_1652 (O_1652,N_14253,N_14335);
and UO_1653 (O_1653,N_14343,N_14875);
nand UO_1654 (O_1654,N_14183,N_14109);
nand UO_1655 (O_1655,N_14178,N_14817);
nand UO_1656 (O_1656,N_14914,N_14629);
and UO_1657 (O_1657,N_14351,N_14755);
or UO_1658 (O_1658,N_14897,N_14913);
nand UO_1659 (O_1659,N_14346,N_14044);
and UO_1660 (O_1660,N_14736,N_14664);
nand UO_1661 (O_1661,N_14391,N_14975);
nand UO_1662 (O_1662,N_14915,N_14080);
nor UO_1663 (O_1663,N_14042,N_14408);
and UO_1664 (O_1664,N_14881,N_14545);
nand UO_1665 (O_1665,N_14364,N_14993);
and UO_1666 (O_1666,N_14985,N_14482);
nand UO_1667 (O_1667,N_14528,N_14112);
nand UO_1668 (O_1668,N_14261,N_14607);
nand UO_1669 (O_1669,N_14385,N_14694);
nor UO_1670 (O_1670,N_14876,N_14505);
nand UO_1671 (O_1671,N_14527,N_14898);
nor UO_1672 (O_1672,N_14788,N_14604);
or UO_1673 (O_1673,N_14197,N_14768);
and UO_1674 (O_1674,N_14310,N_14427);
xor UO_1675 (O_1675,N_14112,N_14158);
and UO_1676 (O_1676,N_14234,N_14770);
and UO_1677 (O_1677,N_14895,N_14641);
nor UO_1678 (O_1678,N_14269,N_14123);
nor UO_1679 (O_1679,N_14976,N_14441);
xor UO_1680 (O_1680,N_14627,N_14816);
xnor UO_1681 (O_1681,N_14813,N_14559);
or UO_1682 (O_1682,N_14590,N_14899);
xor UO_1683 (O_1683,N_14453,N_14566);
xor UO_1684 (O_1684,N_14556,N_14381);
or UO_1685 (O_1685,N_14253,N_14436);
and UO_1686 (O_1686,N_14245,N_14924);
nand UO_1687 (O_1687,N_14681,N_14820);
or UO_1688 (O_1688,N_14764,N_14166);
nand UO_1689 (O_1689,N_14538,N_14811);
or UO_1690 (O_1690,N_14277,N_14142);
and UO_1691 (O_1691,N_14496,N_14857);
nor UO_1692 (O_1692,N_14286,N_14838);
nand UO_1693 (O_1693,N_14149,N_14294);
nand UO_1694 (O_1694,N_14309,N_14479);
nand UO_1695 (O_1695,N_14701,N_14774);
or UO_1696 (O_1696,N_14120,N_14469);
xor UO_1697 (O_1697,N_14681,N_14760);
nand UO_1698 (O_1698,N_14061,N_14325);
or UO_1699 (O_1699,N_14721,N_14713);
and UO_1700 (O_1700,N_14657,N_14618);
or UO_1701 (O_1701,N_14196,N_14035);
nand UO_1702 (O_1702,N_14378,N_14304);
or UO_1703 (O_1703,N_14252,N_14925);
or UO_1704 (O_1704,N_14493,N_14090);
nor UO_1705 (O_1705,N_14452,N_14419);
xor UO_1706 (O_1706,N_14904,N_14591);
nor UO_1707 (O_1707,N_14171,N_14550);
or UO_1708 (O_1708,N_14095,N_14164);
and UO_1709 (O_1709,N_14695,N_14474);
and UO_1710 (O_1710,N_14859,N_14908);
and UO_1711 (O_1711,N_14597,N_14811);
and UO_1712 (O_1712,N_14536,N_14020);
and UO_1713 (O_1713,N_14829,N_14285);
or UO_1714 (O_1714,N_14487,N_14628);
or UO_1715 (O_1715,N_14277,N_14707);
nor UO_1716 (O_1716,N_14843,N_14634);
nand UO_1717 (O_1717,N_14090,N_14746);
nand UO_1718 (O_1718,N_14509,N_14807);
xnor UO_1719 (O_1719,N_14162,N_14308);
or UO_1720 (O_1720,N_14518,N_14650);
nor UO_1721 (O_1721,N_14962,N_14097);
and UO_1722 (O_1722,N_14968,N_14427);
xor UO_1723 (O_1723,N_14153,N_14183);
and UO_1724 (O_1724,N_14348,N_14411);
nor UO_1725 (O_1725,N_14347,N_14823);
nor UO_1726 (O_1726,N_14705,N_14282);
nand UO_1727 (O_1727,N_14559,N_14860);
nand UO_1728 (O_1728,N_14653,N_14334);
nand UO_1729 (O_1729,N_14462,N_14818);
and UO_1730 (O_1730,N_14831,N_14699);
nor UO_1731 (O_1731,N_14580,N_14304);
and UO_1732 (O_1732,N_14708,N_14208);
nor UO_1733 (O_1733,N_14613,N_14753);
nand UO_1734 (O_1734,N_14368,N_14704);
nor UO_1735 (O_1735,N_14173,N_14440);
nand UO_1736 (O_1736,N_14567,N_14405);
and UO_1737 (O_1737,N_14909,N_14031);
xor UO_1738 (O_1738,N_14256,N_14978);
xnor UO_1739 (O_1739,N_14826,N_14065);
and UO_1740 (O_1740,N_14570,N_14271);
nand UO_1741 (O_1741,N_14284,N_14986);
nand UO_1742 (O_1742,N_14114,N_14659);
xor UO_1743 (O_1743,N_14019,N_14285);
nand UO_1744 (O_1744,N_14308,N_14860);
nand UO_1745 (O_1745,N_14493,N_14574);
xor UO_1746 (O_1746,N_14389,N_14778);
or UO_1747 (O_1747,N_14096,N_14494);
nand UO_1748 (O_1748,N_14901,N_14484);
nor UO_1749 (O_1749,N_14661,N_14816);
or UO_1750 (O_1750,N_14610,N_14306);
or UO_1751 (O_1751,N_14618,N_14403);
nor UO_1752 (O_1752,N_14455,N_14896);
nand UO_1753 (O_1753,N_14747,N_14406);
or UO_1754 (O_1754,N_14171,N_14695);
xor UO_1755 (O_1755,N_14321,N_14988);
xnor UO_1756 (O_1756,N_14410,N_14165);
nor UO_1757 (O_1757,N_14049,N_14429);
xor UO_1758 (O_1758,N_14107,N_14881);
or UO_1759 (O_1759,N_14568,N_14221);
or UO_1760 (O_1760,N_14209,N_14354);
or UO_1761 (O_1761,N_14684,N_14431);
xor UO_1762 (O_1762,N_14470,N_14641);
and UO_1763 (O_1763,N_14412,N_14010);
nand UO_1764 (O_1764,N_14425,N_14077);
nand UO_1765 (O_1765,N_14087,N_14307);
nor UO_1766 (O_1766,N_14198,N_14235);
nor UO_1767 (O_1767,N_14127,N_14861);
xor UO_1768 (O_1768,N_14184,N_14319);
nor UO_1769 (O_1769,N_14729,N_14843);
nor UO_1770 (O_1770,N_14782,N_14408);
nor UO_1771 (O_1771,N_14917,N_14138);
or UO_1772 (O_1772,N_14644,N_14919);
xnor UO_1773 (O_1773,N_14774,N_14179);
or UO_1774 (O_1774,N_14307,N_14604);
or UO_1775 (O_1775,N_14577,N_14012);
and UO_1776 (O_1776,N_14389,N_14054);
nor UO_1777 (O_1777,N_14628,N_14406);
nor UO_1778 (O_1778,N_14680,N_14375);
and UO_1779 (O_1779,N_14748,N_14468);
or UO_1780 (O_1780,N_14293,N_14982);
xor UO_1781 (O_1781,N_14169,N_14578);
or UO_1782 (O_1782,N_14628,N_14701);
xnor UO_1783 (O_1783,N_14530,N_14159);
nand UO_1784 (O_1784,N_14554,N_14935);
and UO_1785 (O_1785,N_14990,N_14211);
or UO_1786 (O_1786,N_14575,N_14847);
or UO_1787 (O_1787,N_14406,N_14504);
xnor UO_1788 (O_1788,N_14168,N_14128);
xor UO_1789 (O_1789,N_14344,N_14925);
nand UO_1790 (O_1790,N_14936,N_14786);
xnor UO_1791 (O_1791,N_14582,N_14247);
and UO_1792 (O_1792,N_14696,N_14112);
nand UO_1793 (O_1793,N_14494,N_14750);
nand UO_1794 (O_1794,N_14451,N_14562);
and UO_1795 (O_1795,N_14595,N_14796);
nor UO_1796 (O_1796,N_14513,N_14700);
nand UO_1797 (O_1797,N_14970,N_14337);
and UO_1798 (O_1798,N_14869,N_14446);
or UO_1799 (O_1799,N_14172,N_14686);
nand UO_1800 (O_1800,N_14147,N_14205);
or UO_1801 (O_1801,N_14209,N_14808);
xnor UO_1802 (O_1802,N_14620,N_14590);
nand UO_1803 (O_1803,N_14229,N_14329);
or UO_1804 (O_1804,N_14889,N_14133);
and UO_1805 (O_1805,N_14478,N_14151);
nor UO_1806 (O_1806,N_14018,N_14978);
nor UO_1807 (O_1807,N_14027,N_14237);
xor UO_1808 (O_1808,N_14152,N_14810);
nand UO_1809 (O_1809,N_14170,N_14227);
and UO_1810 (O_1810,N_14380,N_14681);
nand UO_1811 (O_1811,N_14662,N_14629);
xor UO_1812 (O_1812,N_14832,N_14769);
or UO_1813 (O_1813,N_14988,N_14110);
or UO_1814 (O_1814,N_14892,N_14062);
or UO_1815 (O_1815,N_14905,N_14844);
nor UO_1816 (O_1816,N_14517,N_14670);
nor UO_1817 (O_1817,N_14178,N_14852);
and UO_1818 (O_1818,N_14847,N_14727);
or UO_1819 (O_1819,N_14426,N_14197);
nor UO_1820 (O_1820,N_14797,N_14001);
and UO_1821 (O_1821,N_14671,N_14254);
and UO_1822 (O_1822,N_14836,N_14976);
and UO_1823 (O_1823,N_14454,N_14939);
and UO_1824 (O_1824,N_14931,N_14920);
xnor UO_1825 (O_1825,N_14548,N_14600);
xor UO_1826 (O_1826,N_14330,N_14639);
or UO_1827 (O_1827,N_14404,N_14031);
nor UO_1828 (O_1828,N_14357,N_14536);
xor UO_1829 (O_1829,N_14692,N_14478);
xnor UO_1830 (O_1830,N_14595,N_14517);
nor UO_1831 (O_1831,N_14943,N_14903);
and UO_1832 (O_1832,N_14618,N_14156);
or UO_1833 (O_1833,N_14500,N_14873);
nand UO_1834 (O_1834,N_14442,N_14053);
xor UO_1835 (O_1835,N_14599,N_14617);
nor UO_1836 (O_1836,N_14306,N_14518);
xor UO_1837 (O_1837,N_14921,N_14067);
nor UO_1838 (O_1838,N_14246,N_14716);
nand UO_1839 (O_1839,N_14254,N_14093);
or UO_1840 (O_1840,N_14712,N_14548);
xnor UO_1841 (O_1841,N_14313,N_14418);
xnor UO_1842 (O_1842,N_14238,N_14070);
xnor UO_1843 (O_1843,N_14547,N_14825);
nand UO_1844 (O_1844,N_14385,N_14850);
or UO_1845 (O_1845,N_14279,N_14066);
and UO_1846 (O_1846,N_14903,N_14843);
or UO_1847 (O_1847,N_14836,N_14477);
nand UO_1848 (O_1848,N_14930,N_14206);
nor UO_1849 (O_1849,N_14743,N_14897);
or UO_1850 (O_1850,N_14577,N_14839);
nor UO_1851 (O_1851,N_14370,N_14645);
xnor UO_1852 (O_1852,N_14774,N_14078);
nand UO_1853 (O_1853,N_14084,N_14419);
or UO_1854 (O_1854,N_14578,N_14278);
xnor UO_1855 (O_1855,N_14611,N_14270);
xnor UO_1856 (O_1856,N_14860,N_14563);
and UO_1857 (O_1857,N_14653,N_14323);
nor UO_1858 (O_1858,N_14314,N_14916);
nor UO_1859 (O_1859,N_14087,N_14638);
or UO_1860 (O_1860,N_14123,N_14858);
or UO_1861 (O_1861,N_14994,N_14768);
and UO_1862 (O_1862,N_14156,N_14997);
and UO_1863 (O_1863,N_14181,N_14076);
or UO_1864 (O_1864,N_14382,N_14895);
xnor UO_1865 (O_1865,N_14203,N_14768);
and UO_1866 (O_1866,N_14482,N_14821);
nor UO_1867 (O_1867,N_14122,N_14101);
nor UO_1868 (O_1868,N_14357,N_14311);
xnor UO_1869 (O_1869,N_14814,N_14951);
and UO_1870 (O_1870,N_14962,N_14901);
and UO_1871 (O_1871,N_14677,N_14068);
nand UO_1872 (O_1872,N_14749,N_14529);
nor UO_1873 (O_1873,N_14054,N_14528);
nor UO_1874 (O_1874,N_14125,N_14535);
or UO_1875 (O_1875,N_14641,N_14030);
nor UO_1876 (O_1876,N_14585,N_14307);
and UO_1877 (O_1877,N_14991,N_14755);
nand UO_1878 (O_1878,N_14700,N_14407);
xor UO_1879 (O_1879,N_14116,N_14159);
nand UO_1880 (O_1880,N_14397,N_14810);
nor UO_1881 (O_1881,N_14521,N_14928);
or UO_1882 (O_1882,N_14421,N_14302);
or UO_1883 (O_1883,N_14153,N_14214);
or UO_1884 (O_1884,N_14441,N_14007);
nor UO_1885 (O_1885,N_14964,N_14273);
xor UO_1886 (O_1886,N_14769,N_14694);
nor UO_1887 (O_1887,N_14030,N_14994);
nor UO_1888 (O_1888,N_14678,N_14366);
nand UO_1889 (O_1889,N_14796,N_14180);
nor UO_1890 (O_1890,N_14164,N_14231);
xor UO_1891 (O_1891,N_14553,N_14382);
or UO_1892 (O_1892,N_14856,N_14196);
and UO_1893 (O_1893,N_14829,N_14035);
xor UO_1894 (O_1894,N_14277,N_14800);
xor UO_1895 (O_1895,N_14762,N_14600);
xnor UO_1896 (O_1896,N_14285,N_14477);
and UO_1897 (O_1897,N_14372,N_14335);
nand UO_1898 (O_1898,N_14247,N_14099);
xor UO_1899 (O_1899,N_14475,N_14686);
or UO_1900 (O_1900,N_14405,N_14149);
nor UO_1901 (O_1901,N_14821,N_14418);
xnor UO_1902 (O_1902,N_14011,N_14030);
and UO_1903 (O_1903,N_14396,N_14369);
nand UO_1904 (O_1904,N_14111,N_14804);
and UO_1905 (O_1905,N_14867,N_14960);
nand UO_1906 (O_1906,N_14617,N_14512);
and UO_1907 (O_1907,N_14745,N_14649);
nand UO_1908 (O_1908,N_14508,N_14552);
nor UO_1909 (O_1909,N_14077,N_14304);
nand UO_1910 (O_1910,N_14740,N_14397);
or UO_1911 (O_1911,N_14595,N_14574);
nand UO_1912 (O_1912,N_14895,N_14579);
nor UO_1913 (O_1913,N_14723,N_14562);
xnor UO_1914 (O_1914,N_14462,N_14982);
or UO_1915 (O_1915,N_14387,N_14077);
or UO_1916 (O_1916,N_14198,N_14707);
nor UO_1917 (O_1917,N_14478,N_14674);
nand UO_1918 (O_1918,N_14709,N_14144);
and UO_1919 (O_1919,N_14580,N_14513);
nand UO_1920 (O_1920,N_14071,N_14004);
and UO_1921 (O_1921,N_14684,N_14151);
and UO_1922 (O_1922,N_14927,N_14049);
and UO_1923 (O_1923,N_14995,N_14314);
nand UO_1924 (O_1924,N_14095,N_14144);
and UO_1925 (O_1925,N_14402,N_14359);
nand UO_1926 (O_1926,N_14921,N_14813);
and UO_1927 (O_1927,N_14427,N_14403);
nor UO_1928 (O_1928,N_14201,N_14502);
and UO_1929 (O_1929,N_14230,N_14198);
or UO_1930 (O_1930,N_14941,N_14315);
or UO_1931 (O_1931,N_14935,N_14975);
nand UO_1932 (O_1932,N_14652,N_14180);
and UO_1933 (O_1933,N_14149,N_14186);
nor UO_1934 (O_1934,N_14275,N_14676);
nor UO_1935 (O_1935,N_14513,N_14693);
xnor UO_1936 (O_1936,N_14573,N_14931);
nand UO_1937 (O_1937,N_14911,N_14543);
and UO_1938 (O_1938,N_14286,N_14006);
and UO_1939 (O_1939,N_14409,N_14430);
nor UO_1940 (O_1940,N_14632,N_14172);
xnor UO_1941 (O_1941,N_14148,N_14470);
nor UO_1942 (O_1942,N_14110,N_14505);
nand UO_1943 (O_1943,N_14433,N_14391);
nand UO_1944 (O_1944,N_14712,N_14309);
nand UO_1945 (O_1945,N_14995,N_14601);
nor UO_1946 (O_1946,N_14920,N_14649);
and UO_1947 (O_1947,N_14068,N_14534);
nand UO_1948 (O_1948,N_14308,N_14893);
xnor UO_1949 (O_1949,N_14861,N_14919);
nand UO_1950 (O_1950,N_14946,N_14159);
or UO_1951 (O_1951,N_14128,N_14056);
nor UO_1952 (O_1952,N_14869,N_14110);
nand UO_1953 (O_1953,N_14498,N_14373);
nand UO_1954 (O_1954,N_14297,N_14224);
and UO_1955 (O_1955,N_14361,N_14999);
xor UO_1956 (O_1956,N_14350,N_14513);
or UO_1957 (O_1957,N_14323,N_14563);
nor UO_1958 (O_1958,N_14949,N_14659);
and UO_1959 (O_1959,N_14163,N_14558);
xnor UO_1960 (O_1960,N_14494,N_14835);
and UO_1961 (O_1961,N_14368,N_14904);
or UO_1962 (O_1962,N_14879,N_14901);
xor UO_1963 (O_1963,N_14803,N_14139);
nor UO_1964 (O_1964,N_14427,N_14910);
nor UO_1965 (O_1965,N_14349,N_14063);
or UO_1966 (O_1966,N_14119,N_14265);
or UO_1967 (O_1967,N_14812,N_14636);
and UO_1968 (O_1968,N_14598,N_14794);
or UO_1969 (O_1969,N_14503,N_14168);
nand UO_1970 (O_1970,N_14886,N_14713);
or UO_1971 (O_1971,N_14764,N_14054);
nor UO_1972 (O_1972,N_14214,N_14160);
xor UO_1973 (O_1973,N_14455,N_14813);
nor UO_1974 (O_1974,N_14914,N_14806);
and UO_1975 (O_1975,N_14859,N_14694);
or UO_1976 (O_1976,N_14305,N_14374);
and UO_1977 (O_1977,N_14580,N_14727);
or UO_1978 (O_1978,N_14341,N_14645);
nor UO_1979 (O_1979,N_14127,N_14946);
nand UO_1980 (O_1980,N_14226,N_14169);
xnor UO_1981 (O_1981,N_14604,N_14415);
and UO_1982 (O_1982,N_14902,N_14630);
or UO_1983 (O_1983,N_14233,N_14038);
or UO_1984 (O_1984,N_14233,N_14562);
nor UO_1985 (O_1985,N_14988,N_14995);
or UO_1986 (O_1986,N_14822,N_14305);
and UO_1987 (O_1987,N_14986,N_14501);
nor UO_1988 (O_1988,N_14484,N_14576);
nand UO_1989 (O_1989,N_14240,N_14030);
or UO_1990 (O_1990,N_14406,N_14039);
and UO_1991 (O_1991,N_14195,N_14432);
xnor UO_1992 (O_1992,N_14730,N_14233);
nor UO_1993 (O_1993,N_14533,N_14914);
nor UO_1994 (O_1994,N_14114,N_14903);
xnor UO_1995 (O_1995,N_14666,N_14467);
and UO_1996 (O_1996,N_14008,N_14158);
xor UO_1997 (O_1997,N_14449,N_14418);
nand UO_1998 (O_1998,N_14659,N_14190);
or UO_1999 (O_1999,N_14877,N_14257);
endmodule