module basic_1000_10000_1500_100_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_747,In_930);
or U1 (N_1,In_482,In_91);
nand U2 (N_2,In_759,In_289);
nand U3 (N_3,In_235,In_379);
or U4 (N_4,In_674,In_226);
xnor U5 (N_5,In_439,In_621);
or U6 (N_6,In_384,In_590);
and U7 (N_7,In_151,In_497);
and U8 (N_8,In_98,In_523);
and U9 (N_9,In_274,In_798);
xor U10 (N_10,In_34,In_706);
and U11 (N_11,In_503,In_432);
and U12 (N_12,In_312,In_317);
nor U13 (N_13,In_69,In_137);
xnor U14 (N_14,In_173,In_760);
and U15 (N_15,In_501,In_1);
and U16 (N_16,In_638,In_500);
xnor U17 (N_17,In_163,In_766);
nand U18 (N_18,In_936,In_722);
nor U19 (N_19,In_829,In_389);
nor U20 (N_20,In_825,In_239);
and U21 (N_21,In_918,In_333);
nor U22 (N_22,In_189,In_701);
nor U23 (N_23,In_716,In_277);
nand U24 (N_24,In_818,In_492);
xnor U25 (N_25,In_461,In_190);
or U26 (N_26,In_487,In_550);
or U27 (N_27,In_38,In_229);
nand U28 (N_28,In_643,In_376);
nand U29 (N_29,In_102,In_49);
nand U30 (N_30,In_132,In_0);
or U31 (N_31,In_107,In_982);
and U32 (N_32,In_844,In_115);
or U33 (N_33,In_17,In_308);
xor U34 (N_34,In_567,In_542);
xor U35 (N_35,In_426,In_950);
nand U36 (N_36,In_291,In_271);
and U37 (N_37,In_207,In_3);
nand U38 (N_38,In_357,In_11);
or U39 (N_39,In_519,In_719);
xnor U40 (N_40,In_361,In_336);
nand U41 (N_41,In_404,In_203);
or U42 (N_42,In_632,In_608);
nand U43 (N_43,In_339,In_170);
xnor U44 (N_44,In_961,In_453);
or U45 (N_45,In_616,In_718);
and U46 (N_46,In_983,In_954);
nand U47 (N_47,In_628,In_721);
nor U48 (N_48,In_378,In_438);
xnor U49 (N_49,In_865,In_594);
nand U50 (N_50,In_963,In_978);
nand U51 (N_51,In_228,In_543);
and U52 (N_52,In_39,In_45);
xnor U53 (N_53,In_211,In_295);
or U54 (N_54,In_247,In_757);
nor U55 (N_55,In_222,In_843);
xnor U56 (N_56,In_690,In_462);
xor U57 (N_57,In_960,In_609);
xnor U58 (N_58,In_198,In_79);
nand U59 (N_59,In_791,In_645);
xnor U60 (N_60,In_21,In_510);
or U61 (N_61,In_612,In_631);
and U62 (N_62,In_78,In_332);
nor U63 (N_63,In_301,In_576);
nor U64 (N_64,In_342,In_705);
xnor U65 (N_65,In_552,In_19);
nor U66 (N_66,In_955,In_823);
xnor U67 (N_67,In_329,In_991);
xnor U68 (N_68,In_304,In_363);
xor U69 (N_69,In_553,In_831);
or U70 (N_70,In_633,In_6);
xnor U71 (N_71,In_33,In_598);
nand U72 (N_72,In_67,In_602);
xnor U73 (N_73,In_422,In_24);
or U74 (N_74,In_143,In_580);
or U75 (N_75,In_514,In_935);
or U76 (N_76,In_990,In_273);
xor U77 (N_77,In_777,In_95);
nor U78 (N_78,In_650,In_181);
nor U79 (N_79,In_356,In_997);
xor U80 (N_80,In_14,In_377);
or U81 (N_81,In_571,In_99);
and U82 (N_82,In_54,In_655);
xnor U83 (N_83,In_326,In_726);
or U84 (N_84,In_898,In_415);
nand U85 (N_85,In_10,In_666);
or U86 (N_86,In_212,In_707);
nand U87 (N_87,In_662,In_306);
or U88 (N_88,In_617,In_485);
or U89 (N_89,In_168,In_434);
nor U90 (N_90,In_278,In_601);
nand U91 (N_91,In_296,In_535);
xor U92 (N_92,In_223,In_187);
xnor U93 (N_93,In_160,In_157);
and U94 (N_94,In_150,In_261);
and U95 (N_95,In_962,In_735);
nand U96 (N_96,In_870,In_806);
or U97 (N_97,In_688,In_209);
nand U98 (N_98,In_814,In_347);
xnor U99 (N_99,In_206,In_520);
nand U100 (N_100,In_345,N_84);
or U101 (N_101,In_886,In_358);
xnor U102 (N_102,In_551,In_882);
and U103 (N_103,In_921,In_913);
nor U104 (N_104,In_344,In_298);
or U105 (N_105,In_391,In_816);
or U106 (N_106,In_942,In_850);
nand U107 (N_107,In_527,In_600);
and U108 (N_108,In_660,In_425);
or U109 (N_109,In_125,In_511);
nand U110 (N_110,In_193,In_723);
and U111 (N_111,In_665,In_986);
nor U112 (N_112,In_903,In_614);
nor U113 (N_113,In_381,N_65);
xor U114 (N_114,In_984,N_93);
nand U115 (N_115,In_945,In_155);
nand U116 (N_116,N_13,In_815);
nand U117 (N_117,In_675,In_324);
and U118 (N_118,N_22,In_569);
nor U119 (N_119,In_50,In_568);
nand U120 (N_120,In_664,In_283);
xor U121 (N_121,In_753,In_836);
or U122 (N_122,N_67,In_540);
or U123 (N_123,In_869,In_738);
nor U124 (N_124,In_549,N_76);
nor U125 (N_125,In_889,In_796);
nor U126 (N_126,In_44,In_595);
nand U127 (N_127,In_491,N_43);
xnor U128 (N_128,In_490,In_746);
nor U129 (N_129,In_443,N_42);
or U130 (N_130,In_775,In_242);
xnor U131 (N_131,In_479,In_793);
nand U132 (N_132,In_530,In_225);
nand U133 (N_133,In_219,N_66);
and U134 (N_134,In_498,In_284);
nand U135 (N_135,In_546,In_998);
nor U136 (N_136,In_974,In_373);
or U137 (N_137,In_365,In_262);
and U138 (N_138,N_37,In_813);
and U139 (N_139,In_893,In_641);
xnor U140 (N_140,N_47,In_504);
xor U141 (N_141,N_98,In_895);
nor U142 (N_142,In_258,In_183);
xnor U143 (N_143,In_362,In_27);
nand U144 (N_144,In_383,In_682);
and U145 (N_145,In_449,In_169);
nand U146 (N_146,In_156,In_400);
and U147 (N_147,N_16,In_750);
nand U148 (N_148,In_88,In_172);
and U149 (N_149,In_894,In_253);
nor U150 (N_150,In_934,In_162);
and U151 (N_151,In_695,In_756);
and U152 (N_152,In_647,In_360);
and U153 (N_153,In_709,In_622);
and U154 (N_154,In_944,In_354);
or U155 (N_155,In_459,In_605);
nor U156 (N_156,In_60,In_84);
or U157 (N_157,In_184,In_513);
and U158 (N_158,In_596,In_409);
or U159 (N_159,In_769,In_348);
or U160 (N_160,In_976,In_956);
xor U161 (N_161,N_44,In_496);
xnor U162 (N_162,In_74,In_30);
xnor U163 (N_163,In_845,In_532);
nand U164 (N_164,In_732,In_15);
xor U165 (N_165,N_2,In_794);
xnor U166 (N_166,N_25,In_764);
nor U167 (N_167,In_557,In_968);
xnor U168 (N_168,In_204,In_186);
and U169 (N_169,In_781,In_4);
nand U170 (N_170,In_120,In_82);
or U171 (N_171,In_464,In_855);
nand U172 (N_172,In_499,In_452);
and U173 (N_173,In_320,In_281);
and U174 (N_174,In_70,N_89);
nor U175 (N_175,In_398,In_819);
nand U176 (N_176,In_86,In_474);
and U177 (N_177,N_7,In_779);
xor U178 (N_178,In_947,In_288);
or U179 (N_179,N_96,In_681);
or U180 (N_180,In_672,In_202);
and U181 (N_181,In_122,In_197);
xnor U182 (N_182,In_280,In_915);
xnor U183 (N_183,In_85,In_914);
nand U184 (N_184,In_531,In_221);
nor U185 (N_185,N_95,In_311);
and U186 (N_186,In_587,In_299);
nand U187 (N_187,In_801,In_410);
or U188 (N_188,In_118,In_581);
xnor U189 (N_189,In_224,In_165);
or U190 (N_190,N_46,In_965);
and U191 (N_191,In_724,In_953);
xnor U192 (N_192,In_573,In_538);
and U193 (N_193,In_254,In_985);
or U194 (N_194,In_57,N_39);
nand U195 (N_195,N_33,In_250);
xnor U196 (N_196,In_698,In_987);
nand U197 (N_197,In_751,In_249);
nand U198 (N_198,In_637,In_938);
or U199 (N_199,In_536,In_846);
nor U200 (N_200,N_115,N_130);
nand U201 (N_201,In_677,In_401);
nand U202 (N_202,N_199,N_108);
nand U203 (N_203,In_372,In_548);
and U204 (N_204,In_959,In_444);
xor U205 (N_205,In_577,N_159);
or U206 (N_206,In_396,In_830);
xnor U207 (N_207,In_23,N_128);
and U208 (N_208,N_171,In_524);
nand U209 (N_209,In_729,In_25);
nand U210 (N_210,In_795,In_68);
or U211 (N_211,In_136,In_896);
nor U212 (N_212,In_649,In_179);
nor U213 (N_213,In_941,In_268);
nor U214 (N_214,In_309,N_78);
nor U215 (N_215,In_335,In_191);
nand U216 (N_216,In_463,In_591);
nor U217 (N_217,N_32,N_196);
and U218 (N_218,N_155,In_436);
xor U219 (N_219,N_85,N_101);
or U220 (N_220,N_58,In_743);
nor U221 (N_221,In_266,In_267);
nor U222 (N_222,In_104,In_822);
or U223 (N_223,In_419,N_88);
or U224 (N_224,In_782,In_758);
or U225 (N_225,In_592,In_270);
xnor U226 (N_226,In_584,In_678);
or U227 (N_227,In_12,In_403);
xor U228 (N_228,N_168,N_11);
nand U229 (N_229,In_127,In_353);
nand U230 (N_230,In_390,In_644);
and U231 (N_231,In_697,In_977);
and U232 (N_232,In_939,In_314);
and U233 (N_233,In_467,In_445);
nand U234 (N_234,In_113,In_87);
and U235 (N_235,In_138,In_611);
and U236 (N_236,In_486,In_528);
xnor U237 (N_237,N_127,In_32);
nor U238 (N_238,In_374,In_251);
xor U239 (N_239,In_689,In_768);
nor U240 (N_240,In_465,N_17);
or U241 (N_241,In_734,In_773);
or U242 (N_242,N_174,In_651);
or U243 (N_243,N_18,N_197);
nor U244 (N_244,N_74,In_979);
nand U245 (N_245,In_446,In_243);
and U246 (N_246,In_663,N_4);
nand U247 (N_247,In_785,N_102);
xnor U248 (N_248,In_94,In_367);
and U249 (N_249,N_122,In_740);
nand U250 (N_250,In_371,In_744);
or U251 (N_251,In_506,In_177);
and U252 (N_252,In_386,In_881);
or U253 (N_253,In_355,In_20);
nand U254 (N_254,In_153,N_79);
nor U255 (N_255,N_179,In_593);
xnor U256 (N_256,N_1,In_880);
xor U257 (N_257,In_282,In_720);
or U258 (N_258,In_946,In_106);
xor U259 (N_259,In_255,N_82);
nand U260 (N_260,In_803,In_131);
and U261 (N_261,In_708,In_62);
nor U262 (N_262,In_233,N_48);
nand U263 (N_263,In_123,In_399);
xor U264 (N_264,N_104,In_725);
nor U265 (N_265,In_244,In_625);
nand U266 (N_266,In_269,In_161);
and U267 (N_267,N_38,In_780);
or U268 (N_268,In_413,In_405);
or U269 (N_269,In_788,In_275);
nor U270 (N_270,In_185,In_901);
nor U271 (N_271,In_739,In_421);
nand U272 (N_272,In_879,N_170);
and U273 (N_273,In_578,N_87);
or U274 (N_274,N_20,In_97);
xor U275 (N_275,N_12,In_676);
and U276 (N_276,N_73,In_630);
and U277 (N_277,In_101,In_860);
nor U278 (N_278,In_512,In_388);
and U279 (N_279,N_41,In_827);
nand U280 (N_280,In_926,In_770);
xor U281 (N_281,In_900,In_703);
xor U282 (N_282,In_731,In_92);
or U283 (N_283,In_303,In_736);
nand U284 (N_284,In_749,In_811);
or U285 (N_285,In_554,In_240);
xor U286 (N_286,In_810,In_76);
or U287 (N_287,N_77,N_35);
nor U288 (N_288,In_236,N_176);
or U289 (N_289,In_826,N_119);
nor U290 (N_290,N_172,In_516);
nand U291 (N_291,N_116,In_652);
nor U292 (N_292,In_544,In_47);
and U293 (N_293,In_103,In_321);
nor U294 (N_294,In_375,In_741);
and U295 (N_295,In_395,In_263);
xnor U296 (N_296,N_175,N_49);
nor U297 (N_297,In_792,In_64);
or U298 (N_298,In_981,In_146);
or U299 (N_299,In_521,In_313);
nor U300 (N_300,N_211,N_36);
xnor U301 (N_301,N_270,N_235);
xnor U302 (N_302,N_54,In_192);
nor U303 (N_303,In_975,In_351);
or U304 (N_304,In_322,In_996);
nor U305 (N_305,In_964,N_83);
xor U306 (N_306,N_253,N_293);
xnor U307 (N_307,In_610,In_340);
or U308 (N_308,In_925,In_636);
nand U309 (N_309,N_154,In_126);
nor U310 (N_310,In_646,N_152);
and U311 (N_311,In_394,N_185);
nor U312 (N_312,N_265,In_680);
xnor U313 (N_313,In_878,In_623);
nand U314 (N_314,In_875,In_885);
nor U315 (N_315,In_809,In_48);
and U316 (N_316,In_564,In_642);
nor U317 (N_317,In_290,In_863);
nor U318 (N_318,In_835,N_21);
xor U319 (N_319,In_116,In_951);
nor U320 (N_320,In_256,N_0);
nand U321 (N_321,In_684,In_285);
and U322 (N_322,N_19,In_957);
or U323 (N_323,In_5,N_278);
nor U324 (N_324,N_145,In_22);
nand U325 (N_325,In_928,In_216);
and U326 (N_326,N_286,In_839);
nand U327 (N_327,In_158,N_255);
nand U328 (N_328,N_169,N_257);
nor U329 (N_329,In_999,N_231);
and U330 (N_330,In_784,In_346);
nor U331 (N_331,In_145,N_214);
nor U332 (N_332,In_7,In_370);
xor U333 (N_333,N_147,In_517);
nand U334 (N_334,In_754,N_269);
nor U335 (N_335,In_349,In_494);
nand U336 (N_336,In_8,In_89);
or U337 (N_337,In_26,N_206);
nor U338 (N_338,In_402,In_110);
nand U339 (N_339,N_258,In_245);
nor U340 (N_340,In_112,N_292);
and U341 (N_341,In_683,In_534);
nand U342 (N_342,In_518,N_166);
and U343 (N_343,In_884,In_460);
nand U344 (N_344,In_331,In_142);
nor U345 (N_345,In_43,In_588);
and U346 (N_346,N_121,In_667);
nor U347 (N_347,In_966,N_259);
nor U348 (N_348,In_994,In_539);
or U349 (N_349,In_417,N_281);
nand U350 (N_350,In_315,In_488);
and U351 (N_351,In_176,In_714);
and U352 (N_352,In_265,N_229);
or U353 (N_353,N_266,In_297);
and U354 (N_354,In_472,In_995);
nand U355 (N_355,In_330,In_635);
or U356 (N_356,In_967,N_51);
nor U357 (N_357,In_727,N_202);
nand U358 (N_358,N_131,In_687);
and U359 (N_359,N_236,In_752);
or U360 (N_360,N_183,N_162);
xnor U361 (N_361,N_124,In_385);
nand U362 (N_362,In_820,N_224);
and U363 (N_363,In_180,N_220);
nor U364 (N_364,In_178,In_134);
nor U365 (N_365,N_72,N_62);
xnor U366 (N_366,In_515,N_28);
xor U367 (N_367,In_495,In_406);
and U368 (N_368,N_272,In_717);
xor U369 (N_369,N_29,N_285);
and U370 (N_370,In_767,In_748);
nor U371 (N_371,N_97,In_72);
nor U372 (N_372,In_246,In_469);
xor U373 (N_373,In_624,In_279);
or U374 (N_374,In_71,In_489);
nor U375 (N_375,In_93,In_971);
nor U376 (N_376,In_407,N_10);
nor U377 (N_377,In_917,In_570);
or U378 (N_378,N_227,In_509);
or U379 (N_379,N_153,In_343);
nand U380 (N_380,N_252,In_42);
or U381 (N_381,In_607,In_90);
nor U382 (N_382,N_191,N_164);
and U383 (N_383,In_615,In_9);
nor U384 (N_384,N_50,N_297);
or U385 (N_385,In_359,In_973);
nor U386 (N_386,N_243,In_582);
nor U387 (N_387,In_411,In_606);
xor U388 (N_388,N_157,N_56);
or U389 (N_389,N_280,N_118);
nand U390 (N_390,In_905,In_73);
and U391 (N_391,N_27,N_52);
and U392 (N_392,In_877,In_380);
or U393 (N_393,In_537,In_484);
nor U394 (N_394,In_883,N_218);
xor U395 (N_395,N_125,N_284);
xor U396 (N_396,N_230,In_970);
nor U397 (N_397,In_114,In_774);
and U398 (N_398,N_298,In_435);
nand U399 (N_399,N_143,In_937);
xnor U400 (N_400,N_358,In_307);
xor U401 (N_401,In_972,In_148);
nand U402 (N_402,In_730,In_437);
nor U403 (N_403,In_199,N_261);
and U404 (N_404,In_59,N_329);
and U405 (N_405,N_212,In_338);
nor U406 (N_406,In_352,In_58);
and U407 (N_407,In_694,N_290);
xor U408 (N_408,In_989,N_26);
nor U409 (N_409,N_379,N_239);
xnor U410 (N_410,N_111,N_385);
xor U411 (N_411,N_15,In_585);
nor U412 (N_412,In_393,N_342);
nor U413 (N_413,In_100,In_711);
and U414 (N_414,In_824,N_354);
nand U415 (N_415,In_857,In_685);
xor U416 (N_416,In_217,N_198);
xnor U417 (N_417,N_393,N_369);
nand U418 (N_418,In_919,N_264);
xnor U419 (N_419,N_283,In_305);
or U420 (N_420,N_362,In_526);
xor U421 (N_421,In_135,In_61);
or U422 (N_422,In_414,In_629);
xor U423 (N_423,In_201,In_525);
xor U424 (N_424,N_40,In_627);
xor U425 (N_425,In_657,In_949);
or U426 (N_426,In_715,In_28);
xnor U427 (N_427,In_856,In_679);
nor U428 (N_428,N_317,In_533);
and U429 (N_429,In_670,N_263);
nand U430 (N_430,N_161,In_252);
nand U431 (N_431,N_207,N_373);
xor U432 (N_432,N_129,In_63);
or U433 (N_433,In_442,N_333);
and U434 (N_434,In_626,N_318);
or U435 (N_435,In_864,N_312);
nand U436 (N_436,In_911,In_565);
nand U437 (N_437,In_907,N_319);
nor U438 (N_438,In_428,N_346);
and U439 (N_439,N_117,In_272);
nor U440 (N_440,In_412,In_130);
nor U441 (N_441,N_142,In_46);
nor U442 (N_442,N_363,In_128);
nand U443 (N_443,In_728,N_330);
and U444 (N_444,N_374,N_303);
and U445 (N_445,In_851,In_904);
or U446 (N_446,In_833,In_659);
xor U447 (N_447,N_248,In_174);
nand U448 (N_448,In_171,N_344);
nand U449 (N_449,N_233,N_364);
nor U450 (N_450,N_387,In_859);
or U451 (N_451,N_282,N_361);
nand U452 (N_452,In_583,N_337);
nor U453 (N_453,In_556,N_240);
or U454 (N_454,N_357,N_69);
and U455 (N_455,In_81,In_572);
nand U456 (N_456,In_144,In_508);
nand U457 (N_457,N_120,N_194);
nand U458 (N_458,N_57,N_5);
xor U459 (N_459,In_891,N_332);
xnor U460 (N_460,In_238,N_215);
xor U461 (N_461,N_192,In_105);
xnor U462 (N_462,In_948,In_188);
or U463 (N_463,In_868,N_241);
and U464 (N_464,N_9,N_322);
nand U465 (N_465,In_364,N_226);
nor U466 (N_466,In_772,N_313);
and U467 (N_467,In_789,In_408);
xor U468 (N_468,In_931,N_70);
xnor U469 (N_469,In_451,In_575);
nand U470 (N_470,N_349,In_502);
or U471 (N_471,N_160,In_597);
nor U472 (N_472,N_398,In_673);
or U473 (N_473,In_765,In_755);
nor U474 (N_474,In_586,In_807);
and U475 (N_475,In_507,In_619);
nor U476 (N_476,N_156,N_203);
nor U477 (N_477,N_113,N_291);
or U478 (N_478,N_378,In_952);
xnor U479 (N_479,In_195,In_866);
nand U480 (N_480,N_351,In_933);
xor U481 (N_481,N_389,In_771);
nor U482 (N_482,N_109,In_154);
and U483 (N_483,In_111,In_832);
or U484 (N_484,In_147,N_80);
xor U485 (N_485,N_68,N_237);
and U486 (N_486,In_80,In_887);
or U487 (N_487,In_117,In_328);
and U488 (N_488,In_13,N_277);
and U489 (N_489,N_34,In_319);
or U490 (N_490,N_133,N_186);
or U491 (N_491,In_232,N_139);
and U492 (N_492,N_201,In_108);
xor U493 (N_493,In_121,In_51);
nand U494 (N_494,In_561,In_558);
nor U495 (N_495,N_340,N_267);
xnor U496 (N_496,In_762,In_215);
or U497 (N_497,N_365,N_132);
xnor U498 (N_498,In_294,In_862);
and U499 (N_499,In_861,N_238);
nor U500 (N_500,In_547,N_181);
nor U501 (N_501,In_52,In_668);
and U502 (N_502,In_906,N_195);
nor U503 (N_503,N_447,In_119);
xnor U504 (N_504,In_327,N_189);
nor U505 (N_505,In_293,N_489);
nor U506 (N_506,In_218,In_416);
nor U507 (N_507,N_419,In_702);
or U508 (N_508,In_529,N_225);
xnor U509 (N_509,In_292,In_841);
nand U510 (N_510,N_327,In_713);
nor U511 (N_511,In_423,N_494);
and U512 (N_512,N_417,In_969);
or U513 (N_513,In_654,N_216);
nor U514 (N_514,N_222,N_366);
and U515 (N_515,In_992,N_436);
or U516 (N_516,N_367,N_484);
or U517 (N_517,N_310,In_802);
nand U518 (N_518,In_213,In_924);
or U519 (N_519,N_427,N_454);
or U520 (N_520,N_453,N_432);
xnor U521 (N_521,N_30,N_23);
and U522 (N_522,N_409,In_257);
and U523 (N_523,N_53,N_420);
nand U524 (N_524,In_234,N_204);
and U525 (N_525,N_136,N_193);
and U526 (N_526,In_276,In_175);
or U527 (N_527,N_444,N_244);
or U528 (N_528,In_763,In_686);
nor U529 (N_529,N_311,In_778);
and U530 (N_530,N_356,N_221);
nand U531 (N_531,In_661,In_541);
nor U532 (N_532,In_696,In_671);
nor U533 (N_533,N_219,N_479);
or U534 (N_534,N_422,In_194);
nand U535 (N_535,N_343,N_251);
or U536 (N_536,N_141,N_302);
nor U537 (N_537,N_403,N_167);
and U538 (N_538,In_337,In_812);
nand U539 (N_539,In_231,In_366);
or U540 (N_540,N_396,N_348);
nor U541 (N_541,In_574,In_958);
xnor U542 (N_542,In_808,N_469);
and U543 (N_543,In_302,N_429);
xor U544 (N_544,N_324,N_81);
xnor U545 (N_545,In_910,In_478);
nand U546 (N_546,N_91,N_71);
or U547 (N_547,N_341,N_99);
or U548 (N_548,N_246,In_842);
or U549 (N_549,In_653,N_213);
nand U550 (N_550,In_699,In_787);
nor U551 (N_551,N_45,N_480);
and U552 (N_552,In_522,In_560);
nor U553 (N_553,In_505,N_471);
nand U554 (N_554,N_497,N_180);
xnor U555 (N_555,N_323,In_873);
and U556 (N_556,N_123,N_209);
or U557 (N_557,N_135,N_232);
nand U558 (N_558,N_86,N_331);
or U559 (N_559,N_483,In_888);
or U560 (N_560,In_83,In_458);
nor U561 (N_561,In_56,In_237);
or U562 (N_562,In_922,In_35);
and U563 (N_563,In_139,N_405);
nand U564 (N_564,N_382,N_462);
nor U565 (N_565,In_943,In_733);
xor U566 (N_566,N_413,N_178);
nor U567 (N_567,In_369,In_420);
nand U568 (N_568,In_797,In_493);
nor U569 (N_569,In_710,N_138);
xnor U570 (N_570,In_545,N_493);
nand U571 (N_571,N_6,In_424);
xnor U572 (N_572,In_848,N_182);
or U573 (N_573,In_429,N_187);
or U574 (N_574,In_620,In_700);
nor U575 (N_575,In_704,In_310);
or U576 (N_576,N_63,In_2);
nor U577 (N_577,In_634,N_390);
or U578 (N_578,N_472,N_395);
and U579 (N_579,In_241,In_37);
nand U580 (N_580,N_360,N_146);
nor U581 (N_581,N_328,N_465);
xor U582 (N_582,In_562,In_927);
nor U583 (N_583,In_325,N_450);
nand U584 (N_584,N_217,In_455);
and U585 (N_585,N_485,In_427);
and U586 (N_586,In_761,N_210);
or U587 (N_587,In_450,N_279);
nor U588 (N_588,N_406,In_164);
and U589 (N_589,N_384,In_109);
or U590 (N_590,In_656,In_742);
nor U591 (N_591,N_24,N_359);
xor U592 (N_592,In_563,N_440);
nor U593 (N_593,N_92,In_599);
xnor U594 (N_594,N_350,N_260);
xor U595 (N_595,In_316,In_471);
nand U596 (N_596,In_899,N_437);
nor U597 (N_597,N_418,N_490);
nand U598 (N_598,N_473,N_60);
nand U599 (N_599,N_307,N_449);
and U600 (N_600,N_445,N_151);
nand U601 (N_601,In_804,In_433);
nand U602 (N_602,N_468,N_520);
or U603 (N_603,In_470,N_534);
xnor U604 (N_604,In_200,N_150);
and U605 (N_605,N_394,N_140);
or U606 (N_606,N_308,In_640);
xor U607 (N_607,N_540,In_259);
nand U608 (N_608,N_64,N_495);
or U609 (N_609,N_527,N_158);
nand U610 (N_610,N_321,N_515);
and U611 (N_611,N_335,N_8);
nor U612 (N_612,N_412,In_786);
and U613 (N_613,N_407,In_940);
and U614 (N_614,N_134,N_564);
and U615 (N_615,In_858,In_923);
and U616 (N_616,N_434,In_849);
xor U617 (N_617,N_190,In_932);
xnor U618 (N_618,In_75,N_250);
nand U619 (N_619,N_397,N_173);
nand U620 (N_620,N_539,N_459);
nor U621 (N_621,N_315,In_392);
or U622 (N_622,In_712,In_847);
and U623 (N_623,In_334,N_438);
or U624 (N_624,N_441,N_506);
nor U625 (N_625,N_326,N_585);
nand U626 (N_626,N_163,In_920);
nand U627 (N_627,N_325,N_103);
nand U628 (N_628,N_205,N_568);
nand U629 (N_629,In_648,In_140);
and U630 (N_630,N_458,In_431);
or U631 (N_631,N_383,N_275);
xor U632 (N_632,In_834,In_988);
nor U633 (N_633,In_318,N_505);
xnor U634 (N_634,N_100,In_397);
nor U635 (N_635,In_890,In_872);
and U636 (N_636,N_481,N_509);
nor U637 (N_637,N_455,In_691);
nor U638 (N_638,N_500,N_518);
nor U639 (N_639,In_876,N_595);
or U640 (N_640,In_776,In_53);
nand U641 (N_641,In_993,In_480);
or U642 (N_642,N_482,N_487);
nand U643 (N_643,N_496,N_561);
xnor U644 (N_644,N_59,In_817);
nand U645 (N_645,N_256,N_289);
nand U646 (N_646,N_376,N_542);
or U647 (N_647,In_618,N_460);
nand U648 (N_648,In_65,In_783);
nand U649 (N_649,N_268,In_182);
xor U650 (N_650,N_347,In_166);
and U651 (N_651,N_535,N_296);
xnor U652 (N_652,In_350,N_305);
and U653 (N_653,N_531,N_563);
xor U654 (N_654,N_591,In_799);
or U655 (N_655,N_421,In_853);
or U656 (N_656,N_245,In_828);
nor U657 (N_657,N_106,N_557);
or U658 (N_658,N_569,In_133);
xnor U659 (N_659,N_314,N_584);
nand U660 (N_660,N_476,N_491);
or U661 (N_661,N_3,N_549);
xor U662 (N_662,In_867,In_248);
nand U663 (N_663,In_897,N_488);
and U664 (N_664,N_400,In_96);
xnor U665 (N_665,N_426,N_565);
and U666 (N_666,N_503,N_165);
or U667 (N_667,N_587,In_323);
nor U668 (N_668,In_167,In_430);
xnor U669 (N_669,In_287,N_149);
and U670 (N_670,N_309,In_902);
nor U671 (N_671,N_528,N_208);
nor U672 (N_672,In_16,In_210);
xnor U673 (N_673,N_94,In_264);
or U674 (N_674,N_271,In_613);
xnor U675 (N_675,N_404,N_474);
and U676 (N_676,N_448,N_596);
and U677 (N_677,N_583,In_214);
nand U678 (N_678,N_401,N_75);
nand U679 (N_679,N_414,In_141);
xor U680 (N_680,In_579,In_18);
and U681 (N_681,In_227,N_274);
nor U682 (N_682,N_288,N_112);
and U683 (N_683,In_205,N_590);
and U684 (N_684,N_467,N_299);
or U685 (N_685,N_456,N_31);
xor U686 (N_686,N_592,In_41);
and U687 (N_687,N_188,N_273);
and U688 (N_688,N_352,In_382);
and U689 (N_689,N_566,In_208);
xor U690 (N_690,N_184,N_439);
xor U691 (N_691,N_525,N_548);
nor U692 (N_692,N_381,In_892);
xnor U693 (N_693,N_533,In_566);
xor U694 (N_694,N_554,N_523);
nor U695 (N_695,N_295,N_200);
nor U696 (N_696,N_416,N_599);
and U697 (N_697,N_538,N_570);
or U698 (N_698,In_466,In_980);
or U699 (N_699,N_550,N_276);
and U700 (N_700,In_418,N_499);
or U701 (N_701,N_696,N_679);
nand U702 (N_702,In_230,In_929);
nor U703 (N_703,N_391,In_805);
and U704 (N_704,N_643,N_148);
and U705 (N_705,N_573,N_144);
nor U706 (N_706,N_639,N_368);
and U707 (N_707,N_606,In_916);
nor U708 (N_708,N_567,N_619);
or U709 (N_709,N_647,N_674);
or U710 (N_710,N_610,N_555);
or U711 (N_711,In_871,N_234);
or U712 (N_712,N_632,N_611);
or U713 (N_713,N_262,N_524);
nand U714 (N_714,N_688,In_368);
or U715 (N_715,N_501,N_578);
and U716 (N_716,N_380,N_682);
nor U717 (N_717,N_510,N_301);
or U718 (N_718,N_553,N_636);
nor U719 (N_719,N_625,N_177);
and U720 (N_720,N_242,N_580);
nor U721 (N_721,N_442,N_593);
or U722 (N_722,N_470,N_623);
xor U723 (N_723,N_695,In_77);
nand U724 (N_724,N_624,N_223);
or U725 (N_725,In_456,In_737);
nand U726 (N_726,N_620,N_613);
or U727 (N_727,In_476,N_601);
nor U728 (N_728,N_486,N_651);
nor U729 (N_729,N_399,N_642);
nor U730 (N_730,N_320,N_228);
or U731 (N_731,N_693,N_655);
or U732 (N_732,N_114,N_677);
xnor U733 (N_733,N_532,N_616);
and U734 (N_734,N_452,In_483);
xor U735 (N_735,N_14,N_517);
nand U736 (N_736,N_552,In_639);
and U737 (N_737,N_294,N_556);
nand U738 (N_738,N_603,N_635);
nand U739 (N_739,In_838,In_693);
nor U740 (N_740,N_423,N_594);
nand U741 (N_741,In_66,In_692);
and U742 (N_742,N_589,N_402);
xor U743 (N_743,N_526,In_473);
nand U744 (N_744,N_687,N_663);
nor U745 (N_745,N_574,N_504);
nand U746 (N_746,N_345,N_254);
and U747 (N_747,N_466,N_435);
and U748 (N_748,In_124,N_615);
or U749 (N_749,N_464,N_637);
or U750 (N_750,N_477,N_628);
and U751 (N_751,N_650,N_137);
nand U752 (N_752,In_800,N_680);
nand U753 (N_753,N_670,N_475);
or U754 (N_754,N_662,N_110);
nand U755 (N_755,In_448,In_29);
xnor U756 (N_756,In_31,N_547);
nand U757 (N_757,N_660,N_551);
or U758 (N_758,N_249,N_664);
nand U759 (N_759,In_477,N_698);
nor U760 (N_760,N_576,N_247);
and U761 (N_761,In_658,N_446);
xnor U762 (N_762,N_575,In_286);
xor U763 (N_763,N_644,N_622);
nand U764 (N_764,N_652,N_463);
xor U765 (N_765,N_654,N_649);
nor U766 (N_766,N_353,N_306);
or U767 (N_767,N_388,N_640);
xnor U768 (N_768,N_507,N_377);
or U769 (N_769,N_571,N_681);
xnor U770 (N_770,N_697,N_641);
or U771 (N_771,N_638,N_582);
xor U772 (N_772,N_577,N_656);
and U773 (N_773,N_689,N_408);
nor U774 (N_774,N_586,In_475);
xnor U775 (N_775,N_692,N_90);
or U776 (N_776,N_699,In_152);
and U777 (N_777,N_672,N_673);
xor U778 (N_778,N_598,N_657);
nor U779 (N_779,N_617,N_375);
nor U780 (N_780,N_107,N_433);
xnor U781 (N_781,N_411,In_555);
and U782 (N_782,N_300,N_424);
nand U783 (N_783,In_457,N_630);
xnor U784 (N_784,N_653,N_648);
nor U785 (N_785,N_629,N_634);
xor U786 (N_786,In_36,N_355);
xor U787 (N_787,In_854,N_543);
and U788 (N_788,N_336,In_603);
or U789 (N_789,In_196,In_745);
nor U790 (N_790,N_621,N_597);
nand U791 (N_791,N_686,N_645);
and U792 (N_792,N_492,In_260);
nor U793 (N_793,N_658,N_631);
or U794 (N_794,N_536,N_287);
nor U795 (N_795,N_684,In_874);
or U796 (N_796,In_220,In_447);
xor U797 (N_797,N_428,N_316);
xor U798 (N_798,N_371,In_559);
nand U799 (N_799,N_608,N_443);
nand U800 (N_800,N_667,N_754);
and U801 (N_801,In_468,N_430);
xnor U802 (N_802,In_341,In_454);
xnor U803 (N_803,N_633,N_668);
or U804 (N_804,N_781,N_786);
nor U805 (N_805,N_715,N_704);
or U806 (N_806,N_709,In_604);
xnor U807 (N_807,N_773,N_609);
nand U808 (N_808,N_694,In_387);
nor U809 (N_809,N_304,N_775);
xnor U810 (N_810,N_415,N_55);
nand U811 (N_811,N_743,N_738);
and U812 (N_812,N_334,N_706);
xnor U813 (N_813,N_744,N_605);
and U814 (N_814,N_798,N_579);
and U815 (N_815,N_782,N_370);
or U816 (N_816,N_126,In_159);
and U817 (N_817,N_607,N_748);
and U818 (N_818,In_441,N_457);
xor U819 (N_819,N_666,N_339);
and U820 (N_820,N_750,N_546);
nand U821 (N_821,In_40,N_516);
and U822 (N_822,N_514,N_522);
or U823 (N_823,In_912,N_762);
xor U824 (N_824,In_149,N_386);
or U825 (N_825,N_779,N_778);
nor U826 (N_826,N_730,N_410);
nor U827 (N_827,In_821,N_105);
or U828 (N_828,N_747,N_739);
xor U829 (N_829,N_724,N_760);
nor U830 (N_830,N_767,N_716);
nor U831 (N_831,N_713,N_794);
xnor U832 (N_832,N_752,N_646);
nand U833 (N_833,N_755,N_338);
nand U834 (N_834,N_707,N_759);
xor U835 (N_835,N_431,N_751);
or U836 (N_836,N_771,N_671);
or U837 (N_837,N_612,N_498);
xor U838 (N_838,N_702,In_481);
nand U839 (N_839,N_511,N_61);
or U840 (N_840,N_729,N_478);
nor U841 (N_841,N_558,N_799);
nand U842 (N_842,N_392,N_451);
or U843 (N_843,N_659,N_519);
nor U844 (N_844,N_722,N_600);
nand U845 (N_845,N_736,N_718);
xor U846 (N_846,N_756,N_726);
xor U847 (N_847,N_602,N_737);
nor U848 (N_848,N_772,N_753);
nor U849 (N_849,N_720,N_793);
nand U850 (N_850,N_774,N_691);
nand U851 (N_851,N_626,In_790);
xor U852 (N_852,N_797,N_559);
and U853 (N_853,N_581,N_719);
xnor U854 (N_854,N_502,N_717);
and U855 (N_855,N_769,N_776);
and U856 (N_856,N_795,N_758);
or U857 (N_857,N_711,N_796);
xor U858 (N_858,N_545,N_705);
xnor U859 (N_859,N_734,N_461);
nand U860 (N_860,N_676,N_768);
nor U861 (N_861,N_683,N_731);
and U862 (N_862,In_300,N_770);
nand U863 (N_863,N_665,N_669);
nor U864 (N_864,N_746,N_588);
and U865 (N_865,N_513,N_560);
and U866 (N_866,N_740,N_791);
xor U867 (N_867,N_788,N_765);
or U868 (N_868,N_690,In_669);
nand U869 (N_869,N_685,In_589);
nand U870 (N_870,In_840,N_530);
xor U871 (N_871,In_909,N_512);
xnor U872 (N_872,In_852,N_562);
and U873 (N_873,N_425,In_440);
nand U874 (N_874,In_55,N_792);
and U875 (N_875,N_712,N_763);
nor U876 (N_876,N_710,N_708);
nor U877 (N_877,N_604,N_618);
or U878 (N_878,N_780,N_537);
nand U879 (N_879,N_508,N_741);
xor U880 (N_880,N_541,N_735);
or U881 (N_881,N_790,N_728);
and U882 (N_882,N_675,N_745);
xnor U883 (N_883,N_785,N_529);
or U884 (N_884,N_727,N_761);
or U885 (N_885,In_837,N_661);
or U886 (N_886,N_714,N_766);
and U887 (N_887,N_627,N_733);
nor U888 (N_888,In_129,N_732);
nand U889 (N_889,N_723,N_721);
nor U890 (N_890,N_372,N_703);
xor U891 (N_891,N_614,N_544);
or U892 (N_892,N_725,N_700);
or U893 (N_893,N_749,N_678);
nand U894 (N_894,N_521,In_908);
xnor U895 (N_895,N_784,N_701);
nand U896 (N_896,N_789,N_572);
nand U897 (N_897,N_742,N_783);
or U898 (N_898,N_787,N_764);
nor U899 (N_899,N_757,N_777);
nor U900 (N_900,N_880,N_806);
or U901 (N_901,N_805,N_835);
xor U902 (N_902,N_807,N_837);
nand U903 (N_903,N_882,N_866);
and U904 (N_904,N_895,N_808);
nand U905 (N_905,N_879,N_862);
and U906 (N_906,N_846,N_830);
nor U907 (N_907,N_871,N_874);
xnor U908 (N_908,N_825,N_824);
and U909 (N_909,N_899,N_864);
nand U910 (N_910,N_881,N_849);
and U911 (N_911,N_811,N_813);
nor U912 (N_912,N_861,N_851);
nand U913 (N_913,N_833,N_840);
xnor U914 (N_914,N_836,N_868);
nor U915 (N_915,N_883,N_845);
xnor U916 (N_916,N_823,N_892);
nor U917 (N_917,N_832,N_886);
nand U918 (N_918,N_810,N_856);
or U919 (N_919,N_884,N_848);
xor U920 (N_920,N_863,N_827);
nand U921 (N_921,N_817,N_819);
nor U922 (N_922,N_821,N_828);
xor U923 (N_923,N_852,N_869);
or U924 (N_924,N_838,N_815);
xor U925 (N_925,N_855,N_812);
xor U926 (N_926,N_844,N_872);
and U927 (N_927,N_818,N_896);
nand U928 (N_928,N_850,N_822);
and U929 (N_929,N_870,N_878);
nand U930 (N_930,N_857,N_814);
nor U931 (N_931,N_809,N_877);
and U932 (N_932,N_893,N_831);
nand U933 (N_933,N_826,N_804);
nor U934 (N_934,N_803,N_834);
nand U935 (N_935,N_843,N_887);
and U936 (N_936,N_820,N_829);
nor U937 (N_937,N_898,N_842);
xor U938 (N_938,N_894,N_891);
or U939 (N_939,N_839,N_867);
xor U940 (N_940,N_875,N_853);
and U941 (N_941,N_876,N_873);
nand U942 (N_942,N_858,N_841);
and U943 (N_943,N_865,N_801);
xnor U944 (N_944,N_847,N_890);
nand U945 (N_945,N_885,N_860);
xnor U946 (N_946,N_897,N_859);
nand U947 (N_947,N_800,N_802);
and U948 (N_948,N_888,N_816);
nand U949 (N_949,N_854,N_889);
or U950 (N_950,N_896,N_861);
or U951 (N_951,N_825,N_843);
nand U952 (N_952,N_841,N_801);
and U953 (N_953,N_818,N_817);
or U954 (N_954,N_800,N_822);
nor U955 (N_955,N_837,N_812);
nand U956 (N_956,N_809,N_859);
nand U957 (N_957,N_887,N_877);
and U958 (N_958,N_840,N_867);
xor U959 (N_959,N_807,N_856);
nor U960 (N_960,N_831,N_867);
xor U961 (N_961,N_863,N_870);
xor U962 (N_962,N_845,N_813);
xnor U963 (N_963,N_893,N_825);
or U964 (N_964,N_853,N_871);
or U965 (N_965,N_825,N_804);
or U966 (N_966,N_872,N_882);
xnor U967 (N_967,N_883,N_852);
xnor U968 (N_968,N_849,N_813);
and U969 (N_969,N_898,N_801);
and U970 (N_970,N_821,N_858);
nand U971 (N_971,N_849,N_844);
xnor U972 (N_972,N_857,N_875);
or U973 (N_973,N_817,N_850);
xnor U974 (N_974,N_846,N_811);
nand U975 (N_975,N_875,N_804);
xnor U976 (N_976,N_856,N_875);
and U977 (N_977,N_867,N_803);
or U978 (N_978,N_866,N_883);
xnor U979 (N_979,N_878,N_804);
xnor U980 (N_980,N_868,N_847);
nand U981 (N_981,N_898,N_812);
and U982 (N_982,N_805,N_822);
nand U983 (N_983,N_834,N_898);
or U984 (N_984,N_866,N_858);
nor U985 (N_985,N_811,N_848);
and U986 (N_986,N_864,N_831);
nor U987 (N_987,N_802,N_877);
xor U988 (N_988,N_868,N_894);
or U989 (N_989,N_836,N_809);
and U990 (N_990,N_804,N_885);
xnor U991 (N_991,N_864,N_841);
nand U992 (N_992,N_857,N_854);
xnor U993 (N_993,N_879,N_816);
nor U994 (N_994,N_850,N_851);
or U995 (N_995,N_845,N_804);
and U996 (N_996,N_823,N_830);
xnor U997 (N_997,N_886,N_842);
xnor U998 (N_998,N_806,N_826);
or U999 (N_999,N_853,N_860);
nor U1000 (N_1000,N_901,N_932);
xor U1001 (N_1001,N_918,N_929);
nand U1002 (N_1002,N_900,N_926);
xnor U1003 (N_1003,N_987,N_956);
nor U1004 (N_1004,N_965,N_974);
xor U1005 (N_1005,N_917,N_997);
and U1006 (N_1006,N_938,N_933);
or U1007 (N_1007,N_950,N_923);
or U1008 (N_1008,N_966,N_924);
or U1009 (N_1009,N_925,N_916);
or U1010 (N_1010,N_991,N_998);
or U1011 (N_1011,N_921,N_903);
or U1012 (N_1012,N_905,N_967);
nand U1013 (N_1013,N_931,N_981);
xnor U1014 (N_1014,N_960,N_961);
nor U1015 (N_1015,N_953,N_978);
nand U1016 (N_1016,N_976,N_927);
xnor U1017 (N_1017,N_944,N_928);
xor U1018 (N_1018,N_910,N_964);
nor U1019 (N_1019,N_954,N_971);
and U1020 (N_1020,N_947,N_937);
or U1021 (N_1021,N_955,N_904);
nor U1022 (N_1022,N_969,N_982);
nand U1023 (N_1023,N_946,N_984);
nand U1024 (N_1024,N_940,N_996);
nand U1025 (N_1025,N_963,N_951);
and U1026 (N_1026,N_922,N_906);
nor U1027 (N_1027,N_945,N_973);
or U1028 (N_1028,N_994,N_999);
or U1029 (N_1029,N_989,N_913);
nand U1030 (N_1030,N_942,N_914);
nand U1031 (N_1031,N_907,N_975);
xnor U1032 (N_1032,N_972,N_968);
or U1033 (N_1033,N_970,N_957);
and U1034 (N_1034,N_988,N_930);
nor U1035 (N_1035,N_990,N_908);
xor U1036 (N_1036,N_902,N_985);
and U1037 (N_1037,N_915,N_936);
and U1038 (N_1038,N_911,N_919);
xnor U1039 (N_1039,N_992,N_952);
nor U1040 (N_1040,N_935,N_959);
nor U1041 (N_1041,N_939,N_909);
and U1042 (N_1042,N_958,N_949);
nor U1043 (N_1043,N_993,N_943);
or U1044 (N_1044,N_948,N_962);
and U1045 (N_1045,N_980,N_983);
or U1046 (N_1046,N_941,N_979);
xnor U1047 (N_1047,N_934,N_912);
nand U1048 (N_1048,N_986,N_977);
nand U1049 (N_1049,N_995,N_920);
xor U1050 (N_1050,N_900,N_962);
and U1051 (N_1051,N_906,N_910);
or U1052 (N_1052,N_937,N_961);
nor U1053 (N_1053,N_904,N_929);
nor U1054 (N_1054,N_990,N_940);
nand U1055 (N_1055,N_973,N_996);
or U1056 (N_1056,N_980,N_987);
nand U1057 (N_1057,N_965,N_982);
nand U1058 (N_1058,N_964,N_984);
and U1059 (N_1059,N_979,N_932);
and U1060 (N_1060,N_918,N_974);
nor U1061 (N_1061,N_979,N_951);
nand U1062 (N_1062,N_952,N_926);
nor U1063 (N_1063,N_935,N_951);
or U1064 (N_1064,N_986,N_954);
xnor U1065 (N_1065,N_910,N_975);
and U1066 (N_1066,N_999,N_950);
xor U1067 (N_1067,N_997,N_945);
and U1068 (N_1068,N_964,N_911);
or U1069 (N_1069,N_903,N_926);
nand U1070 (N_1070,N_904,N_949);
nor U1071 (N_1071,N_946,N_916);
nand U1072 (N_1072,N_910,N_926);
xor U1073 (N_1073,N_967,N_973);
and U1074 (N_1074,N_916,N_938);
or U1075 (N_1075,N_921,N_982);
xor U1076 (N_1076,N_958,N_953);
and U1077 (N_1077,N_910,N_936);
nand U1078 (N_1078,N_935,N_985);
nor U1079 (N_1079,N_938,N_978);
or U1080 (N_1080,N_903,N_925);
nand U1081 (N_1081,N_988,N_990);
nand U1082 (N_1082,N_997,N_948);
or U1083 (N_1083,N_927,N_978);
and U1084 (N_1084,N_936,N_920);
nand U1085 (N_1085,N_925,N_941);
and U1086 (N_1086,N_969,N_933);
xnor U1087 (N_1087,N_921,N_925);
nor U1088 (N_1088,N_945,N_901);
nand U1089 (N_1089,N_950,N_976);
nor U1090 (N_1090,N_942,N_982);
nand U1091 (N_1091,N_968,N_938);
and U1092 (N_1092,N_972,N_941);
xnor U1093 (N_1093,N_993,N_978);
nand U1094 (N_1094,N_990,N_903);
xor U1095 (N_1095,N_900,N_930);
xor U1096 (N_1096,N_911,N_977);
xnor U1097 (N_1097,N_975,N_955);
or U1098 (N_1098,N_986,N_912);
xnor U1099 (N_1099,N_926,N_928);
nor U1100 (N_1100,N_1066,N_1028);
nand U1101 (N_1101,N_1092,N_1091);
xor U1102 (N_1102,N_1036,N_1096);
or U1103 (N_1103,N_1018,N_1088);
xnor U1104 (N_1104,N_1086,N_1049);
xor U1105 (N_1105,N_1027,N_1097);
and U1106 (N_1106,N_1043,N_1022);
nand U1107 (N_1107,N_1065,N_1077);
nand U1108 (N_1108,N_1014,N_1073);
nor U1109 (N_1109,N_1057,N_1008);
and U1110 (N_1110,N_1024,N_1039);
nor U1111 (N_1111,N_1023,N_1087);
or U1112 (N_1112,N_1081,N_1055);
and U1113 (N_1113,N_1054,N_1029);
xor U1114 (N_1114,N_1053,N_1079);
or U1115 (N_1115,N_1031,N_1009);
nand U1116 (N_1116,N_1042,N_1015);
and U1117 (N_1117,N_1032,N_1021);
or U1118 (N_1118,N_1095,N_1068);
or U1119 (N_1119,N_1004,N_1016);
nor U1120 (N_1120,N_1084,N_1030);
xor U1121 (N_1121,N_1076,N_1074);
or U1122 (N_1122,N_1085,N_1063);
nor U1123 (N_1123,N_1026,N_1011);
or U1124 (N_1124,N_1038,N_1040);
and U1125 (N_1125,N_1093,N_1045);
xor U1126 (N_1126,N_1047,N_1098);
nor U1127 (N_1127,N_1025,N_1099);
xnor U1128 (N_1128,N_1046,N_1037);
xor U1129 (N_1129,N_1078,N_1060);
nand U1130 (N_1130,N_1019,N_1048);
nand U1131 (N_1131,N_1094,N_1082);
nor U1132 (N_1132,N_1071,N_1061);
or U1133 (N_1133,N_1090,N_1064);
and U1134 (N_1134,N_1089,N_1035);
or U1135 (N_1135,N_1000,N_1070);
xnor U1136 (N_1136,N_1052,N_1033);
xor U1137 (N_1137,N_1083,N_1059);
and U1138 (N_1138,N_1012,N_1001);
and U1139 (N_1139,N_1003,N_1075);
xor U1140 (N_1140,N_1058,N_1069);
nor U1141 (N_1141,N_1002,N_1010);
nor U1142 (N_1142,N_1067,N_1056);
xor U1143 (N_1143,N_1051,N_1013);
and U1144 (N_1144,N_1006,N_1005);
nor U1145 (N_1145,N_1007,N_1044);
and U1146 (N_1146,N_1072,N_1017);
xnor U1147 (N_1147,N_1020,N_1050);
xnor U1148 (N_1148,N_1041,N_1062);
nor U1149 (N_1149,N_1034,N_1080);
nand U1150 (N_1150,N_1031,N_1025);
and U1151 (N_1151,N_1036,N_1021);
nand U1152 (N_1152,N_1085,N_1042);
nand U1153 (N_1153,N_1088,N_1057);
nor U1154 (N_1154,N_1059,N_1056);
and U1155 (N_1155,N_1008,N_1062);
or U1156 (N_1156,N_1028,N_1090);
or U1157 (N_1157,N_1055,N_1027);
or U1158 (N_1158,N_1095,N_1024);
nor U1159 (N_1159,N_1005,N_1041);
or U1160 (N_1160,N_1005,N_1080);
nor U1161 (N_1161,N_1075,N_1019);
nand U1162 (N_1162,N_1051,N_1097);
or U1163 (N_1163,N_1039,N_1086);
or U1164 (N_1164,N_1094,N_1062);
xnor U1165 (N_1165,N_1026,N_1027);
or U1166 (N_1166,N_1080,N_1000);
nor U1167 (N_1167,N_1026,N_1005);
or U1168 (N_1168,N_1050,N_1026);
or U1169 (N_1169,N_1022,N_1067);
or U1170 (N_1170,N_1055,N_1038);
and U1171 (N_1171,N_1013,N_1004);
or U1172 (N_1172,N_1071,N_1075);
nor U1173 (N_1173,N_1071,N_1055);
xnor U1174 (N_1174,N_1002,N_1099);
or U1175 (N_1175,N_1010,N_1067);
xnor U1176 (N_1176,N_1052,N_1005);
nand U1177 (N_1177,N_1031,N_1029);
or U1178 (N_1178,N_1078,N_1048);
and U1179 (N_1179,N_1026,N_1022);
nor U1180 (N_1180,N_1013,N_1000);
and U1181 (N_1181,N_1068,N_1089);
nand U1182 (N_1182,N_1094,N_1099);
nand U1183 (N_1183,N_1034,N_1037);
xor U1184 (N_1184,N_1097,N_1087);
and U1185 (N_1185,N_1091,N_1045);
xnor U1186 (N_1186,N_1065,N_1011);
nor U1187 (N_1187,N_1059,N_1098);
and U1188 (N_1188,N_1018,N_1059);
and U1189 (N_1189,N_1089,N_1047);
nand U1190 (N_1190,N_1037,N_1014);
nand U1191 (N_1191,N_1036,N_1087);
nand U1192 (N_1192,N_1027,N_1005);
nand U1193 (N_1193,N_1046,N_1090);
xor U1194 (N_1194,N_1007,N_1075);
and U1195 (N_1195,N_1071,N_1078);
and U1196 (N_1196,N_1001,N_1074);
xor U1197 (N_1197,N_1073,N_1068);
nand U1198 (N_1198,N_1036,N_1007);
xor U1199 (N_1199,N_1044,N_1063);
or U1200 (N_1200,N_1174,N_1194);
nand U1201 (N_1201,N_1157,N_1100);
xnor U1202 (N_1202,N_1152,N_1189);
nor U1203 (N_1203,N_1166,N_1135);
nor U1204 (N_1204,N_1120,N_1140);
nor U1205 (N_1205,N_1198,N_1164);
nand U1206 (N_1206,N_1149,N_1102);
nor U1207 (N_1207,N_1114,N_1162);
xnor U1208 (N_1208,N_1179,N_1186);
xor U1209 (N_1209,N_1172,N_1143);
nand U1210 (N_1210,N_1191,N_1103);
or U1211 (N_1211,N_1178,N_1144);
nand U1212 (N_1212,N_1126,N_1109);
and U1213 (N_1213,N_1124,N_1115);
nand U1214 (N_1214,N_1111,N_1136);
or U1215 (N_1215,N_1190,N_1130);
nor U1216 (N_1216,N_1110,N_1112);
nor U1217 (N_1217,N_1145,N_1197);
xor U1218 (N_1218,N_1138,N_1129);
nor U1219 (N_1219,N_1141,N_1139);
or U1220 (N_1220,N_1105,N_1133);
nand U1221 (N_1221,N_1163,N_1137);
or U1222 (N_1222,N_1151,N_1131);
nand U1223 (N_1223,N_1193,N_1187);
nor U1224 (N_1224,N_1176,N_1155);
and U1225 (N_1225,N_1175,N_1159);
or U1226 (N_1226,N_1183,N_1168);
and U1227 (N_1227,N_1113,N_1148);
and U1228 (N_1228,N_1107,N_1142);
nand U1229 (N_1229,N_1118,N_1160);
nor U1230 (N_1230,N_1173,N_1127);
nor U1231 (N_1231,N_1158,N_1156);
nor U1232 (N_1232,N_1161,N_1154);
nand U1233 (N_1233,N_1165,N_1147);
nor U1234 (N_1234,N_1106,N_1119);
and U1235 (N_1235,N_1184,N_1181);
nor U1236 (N_1236,N_1153,N_1180);
nand U1237 (N_1237,N_1150,N_1108);
nor U1238 (N_1238,N_1171,N_1104);
xor U1239 (N_1239,N_1123,N_1121);
or U1240 (N_1240,N_1167,N_1132);
nand U1241 (N_1241,N_1122,N_1169);
nor U1242 (N_1242,N_1188,N_1125);
or U1243 (N_1243,N_1185,N_1177);
or U1244 (N_1244,N_1146,N_1116);
nand U1245 (N_1245,N_1128,N_1192);
xor U1246 (N_1246,N_1182,N_1101);
and U1247 (N_1247,N_1195,N_1170);
nand U1248 (N_1248,N_1196,N_1199);
nor U1249 (N_1249,N_1117,N_1134);
or U1250 (N_1250,N_1169,N_1158);
and U1251 (N_1251,N_1167,N_1116);
xor U1252 (N_1252,N_1137,N_1196);
nand U1253 (N_1253,N_1157,N_1122);
nand U1254 (N_1254,N_1141,N_1161);
nand U1255 (N_1255,N_1175,N_1140);
and U1256 (N_1256,N_1149,N_1138);
nor U1257 (N_1257,N_1142,N_1140);
xnor U1258 (N_1258,N_1172,N_1170);
or U1259 (N_1259,N_1138,N_1104);
and U1260 (N_1260,N_1171,N_1176);
xor U1261 (N_1261,N_1164,N_1135);
nand U1262 (N_1262,N_1165,N_1122);
xor U1263 (N_1263,N_1131,N_1130);
nor U1264 (N_1264,N_1143,N_1162);
and U1265 (N_1265,N_1110,N_1157);
xnor U1266 (N_1266,N_1108,N_1143);
or U1267 (N_1267,N_1193,N_1103);
or U1268 (N_1268,N_1162,N_1178);
xor U1269 (N_1269,N_1157,N_1102);
nor U1270 (N_1270,N_1102,N_1147);
or U1271 (N_1271,N_1113,N_1157);
and U1272 (N_1272,N_1165,N_1105);
nand U1273 (N_1273,N_1159,N_1111);
nand U1274 (N_1274,N_1139,N_1140);
xnor U1275 (N_1275,N_1161,N_1152);
nand U1276 (N_1276,N_1194,N_1187);
nor U1277 (N_1277,N_1199,N_1116);
nand U1278 (N_1278,N_1167,N_1119);
nor U1279 (N_1279,N_1125,N_1192);
nand U1280 (N_1280,N_1101,N_1129);
nand U1281 (N_1281,N_1110,N_1162);
xnor U1282 (N_1282,N_1197,N_1199);
xor U1283 (N_1283,N_1140,N_1147);
and U1284 (N_1284,N_1146,N_1120);
nand U1285 (N_1285,N_1150,N_1189);
xor U1286 (N_1286,N_1137,N_1195);
nor U1287 (N_1287,N_1100,N_1144);
or U1288 (N_1288,N_1103,N_1170);
and U1289 (N_1289,N_1151,N_1129);
xnor U1290 (N_1290,N_1122,N_1146);
xnor U1291 (N_1291,N_1128,N_1154);
nor U1292 (N_1292,N_1143,N_1127);
or U1293 (N_1293,N_1116,N_1150);
nand U1294 (N_1294,N_1176,N_1119);
nand U1295 (N_1295,N_1115,N_1196);
or U1296 (N_1296,N_1138,N_1195);
nand U1297 (N_1297,N_1141,N_1153);
or U1298 (N_1298,N_1144,N_1111);
nor U1299 (N_1299,N_1109,N_1139);
xnor U1300 (N_1300,N_1208,N_1250);
nor U1301 (N_1301,N_1223,N_1226);
nor U1302 (N_1302,N_1272,N_1246);
nand U1303 (N_1303,N_1260,N_1299);
nand U1304 (N_1304,N_1229,N_1241);
or U1305 (N_1305,N_1247,N_1206);
xor U1306 (N_1306,N_1218,N_1245);
or U1307 (N_1307,N_1254,N_1283);
nand U1308 (N_1308,N_1274,N_1234);
nor U1309 (N_1309,N_1291,N_1267);
nand U1310 (N_1310,N_1284,N_1243);
or U1311 (N_1311,N_1235,N_1232);
or U1312 (N_1312,N_1293,N_1236);
and U1313 (N_1313,N_1201,N_1237);
xor U1314 (N_1314,N_1200,N_1242);
nand U1315 (N_1315,N_1249,N_1212);
xor U1316 (N_1316,N_1204,N_1202);
xor U1317 (N_1317,N_1266,N_1248);
nor U1318 (N_1318,N_1231,N_1285);
nand U1319 (N_1319,N_1259,N_1230);
or U1320 (N_1320,N_1262,N_1282);
or U1321 (N_1321,N_1275,N_1251);
xnor U1322 (N_1322,N_1228,N_1215);
or U1323 (N_1323,N_1256,N_1258);
nor U1324 (N_1324,N_1255,N_1219);
or U1325 (N_1325,N_1289,N_1278);
or U1326 (N_1326,N_1225,N_1286);
xnor U1327 (N_1327,N_1280,N_1216);
and U1328 (N_1328,N_1224,N_1244);
nand U1329 (N_1329,N_1205,N_1214);
and U1330 (N_1330,N_1287,N_1210);
nor U1331 (N_1331,N_1261,N_1222);
nor U1332 (N_1332,N_1269,N_1279);
or U1333 (N_1333,N_1297,N_1227);
nand U1334 (N_1334,N_1257,N_1264);
nor U1335 (N_1335,N_1298,N_1288);
and U1336 (N_1336,N_1217,N_1220);
xnor U1337 (N_1337,N_1292,N_1203);
and U1338 (N_1338,N_1239,N_1273);
xor U1339 (N_1339,N_1240,N_1281);
nor U1340 (N_1340,N_1238,N_1221);
xor U1341 (N_1341,N_1268,N_1207);
nand U1342 (N_1342,N_1271,N_1263);
or U1343 (N_1343,N_1211,N_1252);
nor U1344 (N_1344,N_1296,N_1295);
xor U1345 (N_1345,N_1277,N_1294);
nand U1346 (N_1346,N_1270,N_1209);
nor U1347 (N_1347,N_1233,N_1265);
or U1348 (N_1348,N_1276,N_1213);
or U1349 (N_1349,N_1253,N_1290);
nor U1350 (N_1350,N_1217,N_1246);
xnor U1351 (N_1351,N_1223,N_1280);
nor U1352 (N_1352,N_1218,N_1283);
or U1353 (N_1353,N_1257,N_1202);
nand U1354 (N_1354,N_1223,N_1298);
nand U1355 (N_1355,N_1277,N_1214);
or U1356 (N_1356,N_1287,N_1232);
or U1357 (N_1357,N_1236,N_1251);
nor U1358 (N_1358,N_1266,N_1202);
or U1359 (N_1359,N_1224,N_1274);
xor U1360 (N_1360,N_1293,N_1254);
nor U1361 (N_1361,N_1277,N_1212);
and U1362 (N_1362,N_1270,N_1243);
nor U1363 (N_1363,N_1227,N_1210);
xnor U1364 (N_1364,N_1280,N_1259);
and U1365 (N_1365,N_1222,N_1234);
nor U1366 (N_1366,N_1240,N_1269);
and U1367 (N_1367,N_1203,N_1257);
nand U1368 (N_1368,N_1271,N_1225);
or U1369 (N_1369,N_1227,N_1241);
nor U1370 (N_1370,N_1241,N_1256);
nand U1371 (N_1371,N_1212,N_1260);
nor U1372 (N_1372,N_1263,N_1253);
xnor U1373 (N_1373,N_1292,N_1240);
nand U1374 (N_1374,N_1268,N_1236);
nand U1375 (N_1375,N_1225,N_1259);
nor U1376 (N_1376,N_1208,N_1218);
nor U1377 (N_1377,N_1278,N_1281);
and U1378 (N_1378,N_1266,N_1293);
xnor U1379 (N_1379,N_1249,N_1243);
and U1380 (N_1380,N_1200,N_1247);
nor U1381 (N_1381,N_1293,N_1287);
or U1382 (N_1382,N_1284,N_1279);
xnor U1383 (N_1383,N_1222,N_1297);
nor U1384 (N_1384,N_1276,N_1226);
nor U1385 (N_1385,N_1219,N_1294);
xnor U1386 (N_1386,N_1239,N_1221);
nor U1387 (N_1387,N_1235,N_1277);
xor U1388 (N_1388,N_1233,N_1290);
xor U1389 (N_1389,N_1293,N_1289);
and U1390 (N_1390,N_1234,N_1265);
and U1391 (N_1391,N_1218,N_1299);
nor U1392 (N_1392,N_1206,N_1210);
xor U1393 (N_1393,N_1256,N_1233);
nor U1394 (N_1394,N_1229,N_1263);
nor U1395 (N_1395,N_1217,N_1242);
nor U1396 (N_1396,N_1234,N_1221);
nor U1397 (N_1397,N_1265,N_1227);
nand U1398 (N_1398,N_1222,N_1218);
nor U1399 (N_1399,N_1240,N_1267);
and U1400 (N_1400,N_1313,N_1394);
nand U1401 (N_1401,N_1373,N_1380);
nand U1402 (N_1402,N_1379,N_1397);
xnor U1403 (N_1403,N_1372,N_1354);
and U1404 (N_1404,N_1305,N_1392);
xnor U1405 (N_1405,N_1355,N_1361);
or U1406 (N_1406,N_1382,N_1393);
nor U1407 (N_1407,N_1317,N_1328);
or U1408 (N_1408,N_1367,N_1368);
nand U1409 (N_1409,N_1330,N_1311);
nand U1410 (N_1410,N_1395,N_1365);
and U1411 (N_1411,N_1364,N_1337);
nand U1412 (N_1412,N_1327,N_1346);
and U1413 (N_1413,N_1362,N_1352);
or U1414 (N_1414,N_1345,N_1391);
nand U1415 (N_1415,N_1360,N_1310);
nand U1416 (N_1416,N_1307,N_1343);
and U1417 (N_1417,N_1363,N_1374);
nor U1418 (N_1418,N_1390,N_1325);
or U1419 (N_1419,N_1319,N_1399);
and U1420 (N_1420,N_1335,N_1353);
xor U1421 (N_1421,N_1369,N_1385);
nand U1422 (N_1422,N_1387,N_1302);
and U1423 (N_1423,N_1314,N_1331);
xnor U1424 (N_1424,N_1304,N_1383);
xnor U1425 (N_1425,N_1357,N_1301);
and U1426 (N_1426,N_1347,N_1309);
or U1427 (N_1427,N_1303,N_1332);
or U1428 (N_1428,N_1315,N_1329);
nand U1429 (N_1429,N_1378,N_1375);
nor U1430 (N_1430,N_1312,N_1308);
or U1431 (N_1431,N_1388,N_1333);
xnor U1432 (N_1432,N_1340,N_1370);
and U1433 (N_1433,N_1389,N_1341);
nand U1434 (N_1434,N_1316,N_1338);
nand U1435 (N_1435,N_1336,N_1358);
or U1436 (N_1436,N_1356,N_1396);
nor U1437 (N_1437,N_1306,N_1344);
nor U1438 (N_1438,N_1351,N_1348);
and U1439 (N_1439,N_1366,N_1377);
nand U1440 (N_1440,N_1376,N_1318);
nor U1441 (N_1441,N_1350,N_1386);
and U1442 (N_1442,N_1381,N_1371);
and U1443 (N_1443,N_1384,N_1349);
and U1444 (N_1444,N_1323,N_1322);
and U1445 (N_1445,N_1324,N_1398);
nor U1446 (N_1446,N_1321,N_1342);
or U1447 (N_1447,N_1320,N_1334);
nand U1448 (N_1448,N_1359,N_1326);
and U1449 (N_1449,N_1300,N_1339);
nor U1450 (N_1450,N_1326,N_1301);
xnor U1451 (N_1451,N_1312,N_1364);
xor U1452 (N_1452,N_1334,N_1397);
nor U1453 (N_1453,N_1325,N_1356);
nand U1454 (N_1454,N_1364,N_1366);
xnor U1455 (N_1455,N_1312,N_1341);
or U1456 (N_1456,N_1376,N_1351);
xnor U1457 (N_1457,N_1380,N_1322);
nor U1458 (N_1458,N_1347,N_1313);
nor U1459 (N_1459,N_1314,N_1305);
xnor U1460 (N_1460,N_1373,N_1337);
xor U1461 (N_1461,N_1347,N_1383);
or U1462 (N_1462,N_1347,N_1360);
nor U1463 (N_1463,N_1317,N_1383);
xor U1464 (N_1464,N_1365,N_1314);
xnor U1465 (N_1465,N_1339,N_1381);
nand U1466 (N_1466,N_1394,N_1380);
nor U1467 (N_1467,N_1332,N_1346);
nand U1468 (N_1468,N_1355,N_1372);
xnor U1469 (N_1469,N_1343,N_1315);
xor U1470 (N_1470,N_1311,N_1372);
xor U1471 (N_1471,N_1335,N_1330);
xor U1472 (N_1472,N_1306,N_1379);
nand U1473 (N_1473,N_1340,N_1355);
or U1474 (N_1474,N_1376,N_1374);
or U1475 (N_1475,N_1399,N_1393);
and U1476 (N_1476,N_1394,N_1372);
nand U1477 (N_1477,N_1357,N_1343);
nor U1478 (N_1478,N_1310,N_1362);
and U1479 (N_1479,N_1389,N_1305);
nand U1480 (N_1480,N_1367,N_1347);
nand U1481 (N_1481,N_1385,N_1335);
or U1482 (N_1482,N_1301,N_1364);
nor U1483 (N_1483,N_1355,N_1382);
and U1484 (N_1484,N_1324,N_1392);
xnor U1485 (N_1485,N_1356,N_1312);
xnor U1486 (N_1486,N_1379,N_1323);
nand U1487 (N_1487,N_1384,N_1360);
nand U1488 (N_1488,N_1391,N_1373);
xnor U1489 (N_1489,N_1371,N_1333);
and U1490 (N_1490,N_1368,N_1363);
xnor U1491 (N_1491,N_1379,N_1380);
nand U1492 (N_1492,N_1350,N_1370);
and U1493 (N_1493,N_1389,N_1332);
nor U1494 (N_1494,N_1383,N_1346);
nor U1495 (N_1495,N_1373,N_1388);
nor U1496 (N_1496,N_1330,N_1379);
and U1497 (N_1497,N_1319,N_1310);
and U1498 (N_1498,N_1320,N_1352);
or U1499 (N_1499,N_1320,N_1332);
or U1500 (N_1500,N_1450,N_1449);
nand U1501 (N_1501,N_1468,N_1480);
or U1502 (N_1502,N_1431,N_1476);
or U1503 (N_1503,N_1473,N_1484);
or U1504 (N_1504,N_1443,N_1490);
xor U1505 (N_1505,N_1463,N_1456);
nor U1506 (N_1506,N_1413,N_1414);
nor U1507 (N_1507,N_1416,N_1423);
or U1508 (N_1508,N_1433,N_1441);
xnor U1509 (N_1509,N_1471,N_1429);
nor U1510 (N_1510,N_1467,N_1486);
xor U1511 (N_1511,N_1428,N_1422);
xnor U1512 (N_1512,N_1474,N_1410);
nor U1513 (N_1513,N_1405,N_1407);
nand U1514 (N_1514,N_1430,N_1406);
nand U1515 (N_1515,N_1465,N_1472);
xnor U1516 (N_1516,N_1454,N_1427);
nor U1517 (N_1517,N_1448,N_1451);
nand U1518 (N_1518,N_1447,N_1493);
nand U1519 (N_1519,N_1477,N_1419);
nor U1520 (N_1520,N_1408,N_1415);
or U1521 (N_1521,N_1446,N_1432);
and U1522 (N_1522,N_1488,N_1496);
nand U1523 (N_1523,N_1403,N_1479);
nand U1524 (N_1524,N_1444,N_1495);
xnor U1525 (N_1525,N_1499,N_1402);
or U1526 (N_1526,N_1475,N_1460);
nor U1527 (N_1527,N_1436,N_1492);
or U1528 (N_1528,N_1485,N_1455);
nand U1529 (N_1529,N_1401,N_1421);
nand U1530 (N_1530,N_1453,N_1478);
nor U1531 (N_1531,N_1466,N_1418);
or U1532 (N_1532,N_1498,N_1487);
xor U1533 (N_1533,N_1482,N_1458);
or U1534 (N_1534,N_1469,N_1400);
nand U1535 (N_1535,N_1457,N_1434);
nand U1536 (N_1536,N_1470,N_1424);
and U1537 (N_1537,N_1464,N_1445);
nand U1538 (N_1538,N_1411,N_1437);
and U1539 (N_1539,N_1494,N_1439);
xnor U1540 (N_1540,N_1489,N_1481);
nand U1541 (N_1541,N_1497,N_1452);
and U1542 (N_1542,N_1459,N_1404);
xor U1543 (N_1543,N_1438,N_1461);
nand U1544 (N_1544,N_1417,N_1420);
xnor U1545 (N_1545,N_1426,N_1435);
xor U1546 (N_1546,N_1462,N_1440);
nor U1547 (N_1547,N_1409,N_1483);
nand U1548 (N_1548,N_1491,N_1442);
and U1549 (N_1549,N_1412,N_1425);
xnor U1550 (N_1550,N_1464,N_1417);
nor U1551 (N_1551,N_1451,N_1439);
and U1552 (N_1552,N_1416,N_1425);
or U1553 (N_1553,N_1450,N_1423);
and U1554 (N_1554,N_1439,N_1409);
xnor U1555 (N_1555,N_1412,N_1478);
nor U1556 (N_1556,N_1473,N_1411);
or U1557 (N_1557,N_1447,N_1401);
nand U1558 (N_1558,N_1489,N_1448);
or U1559 (N_1559,N_1410,N_1495);
or U1560 (N_1560,N_1467,N_1499);
xor U1561 (N_1561,N_1437,N_1485);
xnor U1562 (N_1562,N_1461,N_1493);
or U1563 (N_1563,N_1490,N_1460);
xor U1564 (N_1564,N_1497,N_1476);
xnor U1565 (N_1565,N_1498,N_1422);
nand U1566 (N_1566,N_1477,N_1437);
nor U1567 (N_1567,N_1435,N_1406);
xnor U1568 (N_1568,N_1490,N_1488);
xor U1569 (N_1569,N_1405,N_1447);
or U1570 (N_1570,N_1449,N_1421);
xnor U1571 (N_1571,N_1468,N_1453);
and U1572 (N_1572,N_1425,N_1449);
xnor U1573 (N_1573,N_1413,N_1420);
and U1574 (N_1574,N_1406,N_1439);
nor U1575 (N_1575,N_1479,N_1400);
xnor U1576 (N_1576,N_1479,N_1486);
or U1577 (N_1577,N_1494,N_1430);
and U1578 (N_1578,N_1446,N_1474);
nor U1579 (N_1579,N_1441,N_1450);
or U1580 (N_1580,N_1499,N_1492);
nor U1581 (N_1581,N_1432,N_1492);
nand U1582 (N_1582,N_1452,N_1482);
nand U1583 (N_1583,N_1406,N_1494);
or U1584 (N_1584,N_1423,N_1431);
and U1585 (N_1585,N_1478,N_1483);
nand U1586 (N_1586,N_1480,N_1409);
nand U1587 (N_1587,N_1493,N_1406);
or U1588 (N_1588,N_1402,N_1413);
or U1589 (N_1589,N_1401,N_1407);
or U1590 (N_1590,N_1464,N_1454);
nand U1591 (N_1591,N_1424,N_1432);
and U1592 (N_1592,N_1477,N_1424);
and U1593 (N_1593,N_1410,N_1424);
nand U1594 (N_1594,N_1454,N_1447);
nand U1595 (N_1595,N_1495,N_1422);
xor U1596 (N_1596,N_1488,N_1450);
or U1597 (N_1597,N_1463,N_1442);
nand U1598 (N_1598,N_1485,N_1482);
xnor U1599 (N_1599,N_1404,N_1447);
nor U1600 (N_1600,N_1596,N_1576);
nor U1601 (N_1601,N_1552,N_1547);
and U1602 (N_1602,N_1575,N_1554);
xnor U1603 (N_1603,N_1539,N_1520);
xor U1604 (N_1604,N_1500,N_1546);
nor U1605 (N_1605,N_1569,N_1589);
nor U1606 (N_1606,N_1579,N_1507);
nor U1607 (N_1607,N_1526,N_1581);
or U1608 (N_1608,N_1551,N_1592);
nand U1609 (N_1609,N_1591,N_1541);
and U1610 (N_1610,N_1513,N_1540);
nor U1611 (N_1611,N_1511,N_1522);
xnor U1612 (N_1612,N_1586,N_1515);
xnor U1613 (N_1613,N_1524,N_1523);
xor U1614 (N_1614,N_1510,N_1594);
xor U1615 (N_1615,N_1543,N_1544);
or U1616 (N_1616,N_1557,N_1536);
nor U1617 (N_1617,N_1514,N_1574);
nor U1618 (N_1618,N_1585,N_1504);
nor U1619 (N_1619,N_1567,N_1508);
nand U1620 (N_1620,N_1517,N_1590);
xor U1621 (N_1621,N_1593,N_1503);
and U1622 (N_1622,N_1519,N_1528);
nor U1623 (N_1623,N_1545,N_1568);
and U1624 (N_1624,N_1599,N_1560);
and U1625 (N_1625,N_1559,N_1565);
nor U1626 (N_1626,N_1577,N_1584);
xnor U1627 (N_1627,N_1570,N_1512);
xor U1628 (N_1628,N_1597,N_1538);
and U1629 (N_1629,N_1558,N_1525);
nor U1630 (N_1630,N_1502,N_1566);
and U1631 (N_1631,N_1527,N_1587);
and U1632 (N_1632,N_1532,N_1542);
and U1633 (N_1633,N_1573,N_1583);
or U1634 (N_1634,N_1555,N_1506);
nor U1635 (N_1635,N_1531,N_1516);
or U1636 (N_1636,N_1505,N_1535);
xnor U1637 (N_1637,N_1529,N_1578);
nand U1638 (N_1638,N_1549,N_1580);
xnor U1639 (N_1639,N_1563,N_1582);
xor U1640 (N_1640,N_1562,N_1534);
xor U1641 (N_1641,N_1595,N_1501);
xnor U1642 (N_1642,N_1533,N_1561);
and U1643 (N_1643,N_1588,N_1521);
xor U1644 (N_1644,N_1518,N_1550);
or U1645 (N_1645,N_1548,N_1556);
nand U1646 (N_1646,N_1571,N_1530);
xor U1647 (N_1647,N_1537,N_1509);
xor U1648 (N_1648,N_1572,N_1564);
nand U1649 (N_1649,N_1598,N_1553);
nand U1650 (N_1650,N_1543,N_1516);
nand U1651 (N_1651,N_1556,N_1538);
nor U1652 (N_1652,N_1560,N_1576);
nand U1653 (N_1653,N_1558,N_1554);
xor U1654 (N_1654,N_1505,N_1538);
nor U1655 (N_1655,N_1517,N_1516);
or U1656 (N_1656,N_1552,N_1568);
nand U1657 (N_1657,N_1570,N_1547);
and U1658 (N_1658,N_1528,N_1585);
xor U1659 (N_1659,N_1533,N_1502);
or U1660 (N_1660,N_1506,N_1522);
nand U1661 (N_1661,N_1558,N_1505);
nand U1662 (N_1662,N_1570,N_1591);
or U1663 (N_1663,N_1520,N_1564);
or U1664 (N_1664,N_1528,N_1552);
and U1665 (N_1665,N_1523,N_1581);
or U1666 (N_1666,N_1507,N_1565);
nand U1667 (N_1667,N_1558,N_1545);
nand U1668 (N_1668,N_1556,N_1587);
xnor U1669 (N_1669,N_1503,N_1568);
xor U1670 (N_1670,N_1577,N_1520);
and U1671 (N_1671,N_1545,N_1541);
nand U1672 (N_1672,N_1585,N_1537);
xnor U1673 (N_1673,N_1541,N_1525);
nand U1674 (N_1674,N_1554,N_1525);
nand U1675 (N_1675,N_1521,N_1590);
or U1676 (N_1676,N_1538,N_1555);
nand U1677 (N_1677,N_1512,N_1598);
xor U1678 (N_1678,N_1536,N_1553);
and U1679 (N_1679,N_1513,N_1516);
nand U1680 (N_1680,N_1589,N_1543);
nor U1681 (N_1681,N_1544,N_1500);
nand U1682 (N_1682,N_1582,N_1583);
or U1683 (N_1683,N_1566,N_1550);
nand U1684 (N_1684,N_1538,N_1504);
nor U1685 (N_1685,N_1529,N_1586);
nor U1686 (N_1686,N_1517,N_1537);
nor U1687 (N_1687,N_1553,N_1580);
nand U1688 (N_1688,N_1584,N_1533);
and U1689 (N_1689,N_1573,N_1507);
xnor U1690 (N_1690,N_1502,N_1572);
nor U1691 (N_1691,N_1597,N_1581);
and U1692 (N_1692,N_1561,N_1505);
xor U1693 (N_1693,N_1535,N_1567);
and U1694 (N_1694,N_1576,N_1537);
nand U1695 (N_1695,N_1582,N_1543);
nand U1696 (N_1696,N_1543,N_1560);
nor U1697 (N_1697,N_1578,N_1581);
xor U1698 (N_1698,N_1586,N_1507);
nand U1699 (N_1699,N_1594,N_1541);
nor U1700 (N_1700,N_1698,N_1650);
or U1701 (N_1701,N_1667,N_1664);
and U1702 (N_1702,N_1668,N_1646);
nand U1703 (N_1703,N_1620,N_1622);
xnor U1704 (N_1704,N_1687,N_1681);
or U1705 (N_1705,N_1606,N_1691);
nor U1706 (N_1706,N_1651,N_1605);
nor U1707 (N_1707,N_1641,N_1654);
or U1708 (N_1708,N_1662,N_1675);
nor U1709 (N_1709,N_1657,N_1665);
or U1710 (N_1710,N_1655,N_1670);
and U1711 (N_1711,N_1640,N_1623);
and U1712 (N_1712,N_1659,N_1683);
and U1713 (N_1713,N_1621,N_1608);
nand U1714 (N_1714,N_1626,N_1678);
nand U1715 (N_1715,N_1642,N_1603);
or U1716 (N_1716,N_1688,N_1663);
or U1717 (N_1717,N_1671,N_1633);
nor U1718 (N_1718,N_1649,N_1638);
xor U1719 (N_1719,N_1631,N_1653);
xnor U1720 (N_1720,N_1679,N_1636);
or U1721 (N_1721,N_1682,N_1611);
and U1722 (N_1722,N_1694,N_1616);
or U1723 (N_1723,N_1697,N_1666);
and U1724 (N_1724,N_1684,N_1689);
nand U1725 (N_1725,N_1673,N_1685);
or U1726 (N_1726,N_1604,N_1674);
xor U1727 (N_1727,N_1602,N_1669);
or U1728 (N_1728,N_1639,N_1613);
nand U1729 (N_1729,N_1692,N_1634);
xnor U1730 (N_1730,N_1635,N_1658);
and U1731 (N_1731,N_1628,N_1647);
or U1732 (N_1732,N_1629,N_1612);
xnor U1733 (N_1733,N_1615,N_1661);
nand U1734 (N_1734,N_1644,N_1695);
or U1735 (N_1735,N_1643,N_1618);
or U1736 (N_1736,N_1686,N_1610);
nor U1737 (N_1737,N_1676,N_1648);
nand U1738 (N_1738,N_1652,N_1609);
xor U1739 (N_1739,N_1677,N_1624);
nand U1740 (N_1740,N_1672,N_1619);
nand U1741 (N_1741,N_1600,N_1632);
nand U1742 (N_1742,N_1696,N_1614);
nor U1743 (N_1743,N_1699,N_1680);
nor U1744 (N_1744,N_1660,N_1617);
nand U1745 (N_1745,N_1690,N_1645);
and U1746 (N_1746,N_1627,N_1601);
xor U1747 (N_1747,N_1625,N_1630);
xor U1748 (N_1748,N_1607,N_1656);
and U1749 (N_1749,N_1637,N_1693);
xnor U1750 (N_1750,N_1647,N_1699);
or U1751 (N_1751,N_1697,N_1644);
nor U1752 (N_1752,N_1617,N_1662);
or U1753 (N_1753,N_1679,N_1600);
nand U1754 (N_1754,N_1691,N_1647);
xnor U1755 (N_1755,N_1689,N_1616);
nand U1756 (N_1756,N_1645,N_1600);
and U1757 (N_1757,N_1673,N_1645);
nand U1758 (N_1758,N_1690,N_1695);
or U1759 (N_1759,N_1693,N_1619);
nand U1760 (N_1760,N_1665,N_1661);
nand U1761 (N_1761,N_1619,N_1625);
nand U1762 (N_1762,N_1678,N_1690);
nor U1763 (N_1763,N_1677,N_1627);
nand U1764 (N_1764,N_1685,N_1663);
xnor U1765 (N_1765,N_1655,N_1605);
and U1766 (N_1766,N_1687,N_1600);
and U1767 (N_1767,N_1697,N_1686);
xor U1768 (N_1768,N_1627,N_1637);
xnor U1769 (N_1769,N_1605,N_1691);
nand U1770 (N_1770,N_1639,N_1616);
or U1771 (N_1771,N_1625,N_1688);
xnor U1772 (N_1772,N_1623,N_1624);
or U1773 (N_1773,N_1661,N_1641);
nand U1774 (N_1774,N_1638,N_1615);
nand U1775 (N_1775,N_1676,N_1632);
nand U1776 (N_1776,N_1652,N_1616);
nor U1777 (N_1777,N_1650,N_1658);
nor U1778 (N_1778,N_1606,N_1617);
and U1779 (N_1779,N_1657,N_1660);
or U1780 (N_1780,N_1687,N_1669);
nand U1781 (N_1781,N_1647,N_1629);
and U1782 (N_1782,N_1641,N_1650);
and U1783 (N_1783,N_1672,N_1697);
nor U1784 (N_1784,N_1635,N_1630);
nand U1785 (N_1785,N_1654,N_1648);
nor U1786 (N_1786,N_1679,N_1603);
or U1787 (N_1787,N_1685,N_1622);
nor U1788 (N_1788,N_1665,N_1618);
xor U1789 (N_1789,N_1661,N_1699);
or U1790 (N_1790,N_1625,N_1609);
nand U1791 (N_1791,N_1699,N_1692);
or U1792 (N_1792,N_1604,N_1671);
nand U1793 (N_1793,N_1638,N_1605);
and U1794 (N_1794,N_1663,N_1628);
xor U1795 (N_1795,N_1691,N_1636);
nor U1796 (N_1796,N_1698,N_1689);
nor U1797 (N_1797,N_1673,N_1669);
nand U1798 (N_1798,N_1673,N_1661);
xnor U1799 (N_1799,N_1694,N_1651);
nor U1800 (N_1800,N_1702,N_1762);
xnor U1801 (N_1801,N_1748,N_1749);
xnor U1802 (N_1802,N_1744,N_1743);
nor U1803 (N_1803,N_1774,N_1769);
nor U1804 (N_1804,N_1721,N_1764);
and U1805 (N_1805,N_1719,N_1772);
nor U1806 (N_1806,N_1728,N_1741);
nor U1807 (N_1807,N_1757,N_1722);
nor U1808 (N_1808,N_1779,N_1782);
nor U1809 (N_1809,N_1738,N_1715);
nand U1810 (N_1810,N_1766,N_1730);
or U1811 (N_1811,N_1704,N_1780);
nand U1812 (N_1812,N_1793,N_1759);
nand U1813 (N_1813,N_1754,N_1787);
nand U1814 (N_1814,N_1765,N_1739);
xnor U1815 (N_1815,N_1768,N_1703);
nor U1816 (N_1816,N_1709,N_1770);
nor U1817 (N_1817,N_1712,N_1714);
and U1818 (N_1818,N_1725,N_1735);
or U1819 (N_1819,N_1700,N_1750);
nor U1820 (N_1820,N_1734,N_1751);
nor U1821 (N_1821,N_1752,N_1777);
and U1822 (N_1822,N_1797,N_1789);
xor U1823 (N_1823,N_1760,N_1740);
and U1824 (N_1824,N_1708,N_1746);
and U1825 (N_1825,N_1724,N_1742);
xor U1826 (N_1826,N_1745,N_1737);
nor U1827 (N_1827,N_1732,N_1753);
and U1828 (N_1828,N_1710,N_1771);
xnor U1829 (N_1829,N_1776,N_1729);
or U1830 (N_1830,N_1773,N_1726);
or U1831 (N_1831,N_1747,N_1720);
and U1832 (N_1832,N_1755,N_1775);
and U1833 (N_1833,N_1786,N_1783);
nand U1834 (N_1834,N_1788,N_1701);
or U1835 (N_1835,N_1718,N_1713);
nor U1836 (N_1836,N_1756,N_1727);
and U1837 (N_1837,N_1761,N_1781);
xnor U1838 (N_1838,N_1717,N_1763);
or U1839 (N_1839,N_1706,N_1733);
or U1840 (N_1840,N_1723,N_1799);
xnor U1841 (N_1841,N_1795,N_1711);
nand U1842 (N_1842,N_1792,N_1778);
and U1843 (N_1843,N_1784,N_1791);
or U1844 (N_1844,N_1767,N_1758);
and U1845 (N_1845,N_1705,N_1796);
or U1846 (N_1846,N_1707,N_1798);
or U1847 (N_1847,N_1716,N_1736);
nand U1848 (N_1848,N_1731,N_1785);
and U1849 (N_1849,N_1790,N_1794);
nand U1850 (N_1850,N_1764,N_1799);
xnor U1851 (N_1851,N_1795,N_1710);
or U1852 (N_1852,N_1759,N_1712);
xnor U1853 (N_1853,N_1727,N_1750);
or U1854 (N_1854,N_1774,N_1767);
nand U1855 (N_1855,N_1728,N_1765);
nand U1856 (N_1856,N_1781,N_1711);
xor U1857 (N_1857,N_1700,N_1707);
and U1858 (N_1858,N_1788,N_1731);
or U1859 (N_1859,N_1763,N_1747);
nor U1860 (N_1860,N_1728,N_1789);
nand U1861 (N_1861,N_1713,N_1781);
and U1862 (N_1862,N_1770,N_1792);
or U1863 (N_1863,N_1704,N_1759);
or U1864 (N_1864,N_1739,N_1751);
or U1865 (N_1865,N_1712,N_1743);
nand U1866 (N_1866,N_1734,N_1732);
nand U1867 (N_1867,N_1759,N_1763);
nand U1868 (N_1868,N_1767,N_1787);
and U1869 (N_1869,N_1755,N_1758);
or U1870 (N_1870,N_1790,N_1709);
or U1871 (N_1871,N_1745,N_1775);
nand U1872 (N_1872,N_1748,N_1779);
nor U1873 (N_1873,N_1720,N_1778);
or U1874 (N_1874,N_1715,N_1731);
xnor U1875 (N_1875,N_1726,N_1779);
and U1876 (N_1876,N_1713,N_1716);
nor U1877 (N_1877,N_1752,N_1723);
xnor U1878 (N_1878,N_1704,N_1711);
or U1879 (N_1879,N_1741,N_1761);
xor U1880 (N_1880,N_1751,N_1798);
xor U1881 (N_1881,N_1713,N_1755);
and U1882 (N_1882,N_1701,N_1725);
and U1883 (N_1883,N_1715,N_1763);
nor U1884 (N_1884,N_1798,N_1794);
and U1885 (N_1885,N_1733,N_1743);
xnor U1886 (N_1886,N_1706,N_1742);
xor U1887 (N_1887,N_1763,N_1746);
nor U1888 (N_1888,N_1711,N_1762);
nand U1889 (N_1889,N_1795,N_1718);
xnor U1890 (N_1890,N_1746,N_1747);
nand U1891 (N_1891,N_1701,N_1791);
and U1892 (N_1892,N_1768,N_1713);
nand U1893 (N_1893,N_1762,N_1740);
nor U1894 (N_1894,N_1761,N_1715);
and U1895 (N_1895,N_1737,N_1788);
nand U1896 (N_1896,N_1758,N_1751);
xor U1897 (N_1897,N_1784,N_1746);
xnor U1898 (N_1898,N_1704,N_1716);
or U1899 (N_1899,N_1711,N_1739);
nand U1900 (N_1900,N_1890,N_1802);
or U1901 (N_1901,N_1876,N_1834);
and U1902 (N_1902,N_1891,N_1848);
and U1903 (N_1903,N_1897,N_1888);
xor U1904 (N_1904,N_1878,N_1889);
xnor U1905 (N_1905,N_1807,N_1844);
and U1906 (N_1906,N_1813,N_1814);
or U1907 (N_1907,N_1870,N_1879);
or U1908 (N_1908,N_1837,N_1832);
or U1909 (N_1909,N_1875,N_1886);
nor U1910 (N_1910,N_1882,N_1872);
or U1911 (N_1911,N_1821,N_1885);
or U1912 (N_1912,N_1853,N_1812);
and U1913 (N_1913,N_1852,N_1858);
or U1914 (N_1914,N_1839,N_1893);
and U1915 (N_1915,N_1895,N_1880);
nor U1916 (N_1916,N_1887,N_1871);
nor U1917 (N_1917,N_1836,N_1846);
xor U1918 (N_1918,N_1830,N_1864);
nand U1919 (N_1919,N_1896,N_1829);
xnor U1920 (N_1920,N_1809,N_1883);
xnor U1921 (N_1921,N_1847,N_1845);
nor U1922 (N_1922,N_1842,N_1861);
xor U1923 (N_1923,N_1850,N_1803);
xnor U1924 (N_1924,N_1867,N_1801);
or U1925 (N_1925,N_1856,N_1819);
and U1926 (N_1926,N_1818,N_1815);
nand U1927 (N_1927,N_1825,N_1873);
or U1928 (N_1928,N_1810,N_1884);
nor U1929 (N_1929,N_1851,N_1800);
xor U1930 (N_1930,N_1805,N_1831);
nand U1931 (N_1931,N_1817,N_1874);
nand U1932 (N_1932,N_1826,N_1804);
or U1933 (N_1933,N_1863,N_1854);
or U1934 (N_1934,N_1841,N_1835);
xor U1935 (N_1935,N_1868,N_1849);
nor U1936 (N_1936,N_1865,N_1898);
nor U1937 (N_1937,N_1824,N_1894);
or U1938 (N_1938,N_1811,N_1827);
and U1939 (N_1939,N_1899,N_1840);
and U1940 (N_1940,N_1820,N_1869);
or U1941 (N_1941,N_1833,N_1843);
nor U1942 (N_1942,N_1857,N_1808);
nor U1943 (N_1943,N_1823,N_1822);
xnor U1944 (N_1944,N_1860,N_1816);
and U1945 (N_1945,N_1806,N_1866);
nor U1946 (N_1946,N_1859,N_1855);
nor U1947 (N_1947,N_1877,N_1828);
or U1948 (N_1948,N_1838,N_1862);
or U1949 (N_1949,N_1881,N_1892);
nor U1950 (N_1950,N_1881,N_1845);
xnor U1951 (N_1951,N_1809,N_1852);
xnor U1952 (N_1952,N_1890,N_1848);
xnor U1953 (N_1953,N_1813,N_1841);
and U1954 (N_1954,N_1820,N_1813);
xnor U1955 (N_1955,N_1850,N_1848);
xor U1956 (N_1956,N_1819,N_1896);
and U1957 (N_1957,N_1871,N_1888);
nand U1958 (N_1958,N_1898,N_1818);
and U1959 (N_1959,N_1820,N_1893);
nand U1960 (N_1960,N_1802,N_1808);
xnor U1961 (N_1961,N_1874,N_1825);
nor U1962 (N_1962,N_1814,N_1810);
and U1963 (N_1963,N_1850,N_1815);
nor U1964 (N_1964,N_1897,N_1874);
nor U1965 (N_1965,N_1897,N_1831);
xnor U1966 (N_1966,N_1870,N_1848);
nor U1967 (N_1967,N_1863,N_1879);
xnor U1968 (N_1968,N_1813,N_1821);
or U1969 (N_1969,N_1800,N_1865);
or U1970 (N_1970,N_1844,N_1859);
or U1971 (N_1971,N_1881,N_1844);
xor U1972 (N_1972,N_1819,N_1863);
nor U1973 (N_1973,N_1865,N_1820);
xnor U1974 (N_1974,N_1861,N_1898);
nor U1975 (N_1975,N_1821,N_1888);
xnor U1976 (N_1976,N_1856,N_1826);
and U1977 (N_1977,N_1833,N_1880);
xor U1978 (N_1978,N_1895,N_1805);
nor U1979 (N_1979,N_1892,N_1857);
xor U1980 (N_1980,N_1877,N_1811);
and U1981 (N_1981,N_1803,N_1852);
and U1982 (N_1982,N_1833,N_1865);
xor U1983 (N_1983,N_1807,N_1867);
nor U1984 (N_1984,N_1879,N_1855);
nor U1985 (N_1985,N_1843,N_1847);
xnor U1986 (N_1986,N_1807,N_1837);
nand U1987 (N_1987,N_1840,N_1817);
xor U1988 (N_1988,N_1808,N_1848);
nand U1989 (N_1989,N_1881,N_1816);
nor U1990 (N_1990,N_1892,N_1852);
and U1991 (N_1991,N_1812,N_1808);
or U1992 (N_1992,N_1801,N_1829);
and U1993 (N_1993,N_1840,N_1804);
nor U1994 (N_1994,N_1825,N_1896);
nor U1995 (N_1995,N_1835,N_1877);
nor U1996 (N_1996,N_1821,N_1822);
and U1997 (N_1997,N_1837,N_1835);
nor U1998 (N_1998,N_1897,N_1807);
nor U1999 (N_1999,N_1814,N_1804);
nand U2000 (N_2000,N_1953,N_1922);
nand U2001 (N_2001,N_1982,N_1916);
or U2002 (N_2002,N_1912,N_1959);
and U2003 (N_2003,N_1937,N_1971);
or U2004 (N_2004,N_1929,N_1907);
or U2005 (N_2005,N_1933,N_1964);
and U2006 (N_2006,N_1990,N_1936);
nand U2007 (N_2007,N_1958,N_1960);
nand U2008 (N_2008,N_1921,N_1915);
nand U2009 (N_2009,N_1952,N_1995);
nand U2010 (N_2010,N_1902,N_1954);
or U2011 (N_2011,N_1926,N_1981);
and U2012 (N_2012,N_1980,N_1955);
nand U2013 (N_2013,N_1943,N_1908);
or U2014 (N_2014,N_1904,N_1913);
nand U2015 (N_2015,N_1901,N_1925);
and U2016 (N_2016,N_1932,N_1944);
and U2017 (N_2017,N_1987,N_1985);
or U2018 (N_2018,N_1919,N_1984);
nor U2019 (N_2019,N_1930,N_1951);
or U2020 (N_2020,N_1947,N_1975);
nand U2021 (N_2021,N_1965,N_1993);
nand U2022 (N_2022,N_1920,N_1957);
nor U2023 (N_2023,N_1978,N_1988);
xnor U2024 (N_2024,N_1923,N_1974);
xor U2025 (N_2025,N_1994,N_1956);
xnor U2026 (N_2026,N_1934,N_1961);
nor U2027 (N_2027,N_1950,N_1977);
xnor U2028 (N_2028,N_1948,N_1939);
xnor U2029 (N_2029,N_1998,N_1979);
and U2030 (N_2030,N_1927,N_1928);
nor U2031 (N_2031,N_1949,N_1962);
and U2032 (N_2032,N_1996,N_1983);
and U2033 (N_2033,N_1918,N_1963);
xor U2034 (N_2034,N_1900,N_1911);
xnor U2035 (N_2035,N_1940,N_1970);
or U2036 (N_2036,N_1986,N_1969);
or U2037 (N_2037,N_1910,N_1905);
xor U2038 (N_2038,N_1935,N_1909);
and U2039 (N_2039,N_1989,N_1914);
or U2040 (N_2040,N_1972,N_1942);
nor U2041 (N_2041,N_1941,N_1991);
and U2042 (N_2042,N_1997,N_1992);
nor U2043 (N_2043,N_1945,N_1967);
or U2044 (N_2044,N_1924,N_1946);
and U2045 (N_2045,N_1931,N_1917);
xnor U2046 (N_2046,N_1999,N_1903);
or U2047 (N_2047,N_1973,N_1938);
or U2048 (N_2048,N_1968,N_1906);
nand U2049 (N_2049,N_1976,N_1966);
and U2050 (N_2050,N_1941,N_1908);
nand U2051 (N_2051,N_1963,N_1951);
nor U2052 (N_2052,N_1901,N_1907);
or U2053 (N_2053,N_1972,N_1911);
xnor U2054 (N_2054,N_1936,N_1974);
or U2055 (N_2055,N_1951,N_1957);
xnor U2056 (N_2056,N_1980,N_1909);
and U2057 (N_2057,N_1968,N_1953);
nor U2058 (N_2058,N_1941,N_1954);
and U2059 (N_2059,N_1992,N_1923);
nor U2060 (N_2060,N_1996,N_1912);
xnor U2061 (N_2061,N_1930,N_1998);
nand U2062 (N_2062,N_1969,N_1922);
or U2063 (N_2063,N_1961,N_1921);
nor U2064 (N_2064,N_1954,N_1918);
xnor U2065 (N_2065,N_1927,N_1976);
xor U2066 (N_2066,N_1974,N_1934);
nor U2067 (N_2067,N_1908,N_1928);
and U2068 (N_2068,N_1932,N_1938);
xnor U2069 (N_2069,N_1909,N_1996);
nand U2070 (N_2070,N_1997,N_1999);
or U2071 (N_2071,N_1999,N_1966);
nor U2072 (N_2072,N_1987,N_1982);
or U2073 (N_2073,N_1922,N_1995);
or U2074 (N_2074,N_1912,N_1990);
and U2075 (N_2075,N_1922,N_1986);
xor U2076 (N_2076,N_1998,N_1952);
or U2077 (N_2077,N_1918,N_1996);
nand U2078 (N_2078,N_1934,N_1946);
nor U2079 (N_2079,N_1955,N_1984);
xnor U2080 (N_2080,N_1986,N_1974);
and U2081 (N_2081,N_1988,N_1997);
nor U2082 (N_2082,N_1943,N_1900);
nand U2083 (N_2083,N_1991,N_1925);
or U2084 (N_2084,N_1939,N_1923);
and U2085 (N_2085,N_1971,N_1976);
xnor U2086 (N_2086,N_1928,N_1992);
or U2087 (N_2087,N_1908,N_1999);
xnor U2088 (N_2088,N_1939,N_1910);
xor U2089 (N_2089,N_1962,N_1943);
and U2090 (N_2090,N_1953,N_1937);
xnor U2091 (N_2091,N_1917,N_1936);
xor U2092 (N_2092,N_1964,N_1958);
nand U2093 (N_2093,N_1980,N_1979);
nor U2094 (N_2094,N_1904,N_1959);
nand U2095 (N_2095,N_1942,N_1941);
and U2096 (N_2096,N_1937,N_1903);
and U2097 (N_2097,N_1914,N_1908);
xor U2098 (N_2098,N_1968,N_1949);
nor U2099 (N_2099,N_1932,N_1924);
and U2100 (N_2100,N_2032,N_2021);
xor U2101 (N_2101,N_2093,N_2059);
and U2102 (N_2102,N_2017,N_2038);
nor U2103 (N_2103,N_2031,N_2062);
and U2104 (N_2104,N_2068,N_2092);
nor U2105 (N_2105,N_2004,N_2066);
and U2106 (N_2106,N_2053,N_2088);
nor U2107 (N_2107,N_2078,N_2033);
and U2108 (N_2108,N_2075,N_2011);
nor U2109 (N_2109,N_2094,N_2001);
or U2110 (N_2110,N_2065,N_2002);
nor U2111 (N_2111,N_2003,N_2030);
nor U2112 (N_2112,N_2085,N_2025);
or U2113 (N_2113,N_2014,N_2063);
and U2114 (N_2114,N_2056,N_2047);
xnor U2115 (N_2115,N_2079,N_2041);
nand U2116 (N_2116,N_2044,N_2042);
or U2117 (N_2117,N_2070,N_2034);
nand U2118 (N_2118,N_2029,N_2067);
and U2119 (N_2119,N_2005,N_2027);
and U2120 (N_2120,N_2028,N_2097);
nand U2121 (N_2121,N_2087,N_2071);
or U2122 (N_2122,N_2051,N_2072);
and U2123 (N_2123,N_2008,N_2074);
nand U2124 (N_2124,N_2081,N_2023);
nor U2125 (N_2125,N_2077,N_2082);
or U2126 (N_2126,N_2012,N_2060);
and U2127 (N_2127,N_2098,N_2040);
xor U2128 (N_2128,N_2010,N_2058);
xor U2129 (N_2129,N_2064,N_2009);
xor U2130 (N_2130,N_2006,N_2019);
nand U2131 (N_2131,N_2073,N_2035);
xnor U2132 (N_2132,N_2057,N_2050);
nand U2133 (N_2133,N_2022,N_2061);
nor U2134 (N_2134,N_2076,N_2052);
nor U2135 (N_2135,N_2080,N_2043);
nor U2136 (N_2136,N_2086,N_2083);
nand U2137 (N_2137,N_2096,N_2069);
and U2138 (N_2138,N_2007,N_2045);
and U2139 (N_2139,N_2024,N_2018);
xnor U2140 (N_2140,N_2036,N_2095);
nand U2141 (N_2141,N_2049,N_2013);
nand U2142 (N_2142,N_2090,N_2039);
or U2143 (N_2143,N_2089,N_2048);
xor U2144 (N_2144,N_2016,N_2020);
nor U2145 (N_2145,N_2026,N_2037);
nand U2146 (N_2146,N_2015,N_2000);
and U2147 (N_2147,N_2055,N_2054);
nand U2148 (N_2148,N_2084,N_2091);
xor U2149 (N_2149,N_2099,N_2046);
xnor U2150 (N_2150,N_2038,N_2090);
or U2151 (N_2151,N_2042,N_2011);
nand U2152 (N_2152,N_2071,N_2096);
nand U2153 (N_2153,N_2010,N_2056);
or U2154 (N_2154,N_2023,N_2069);
and U2155 (N_2155,N_2042,N_2068);
nor U2156 (N_2156,N_2021,N_2002);
or U2157 (N_2157,N_2091,N_2066);
and U2158 (N_2158,N_2052,N_2014);
nor U2159 (N_2159,N_2054,N_2028);
and U2160 (N_2160,N_2088,N_2021);
and U2161 (N_2161,N_2002,N_2096);
nand U2162 (N_2162,N_2058,N_2047);
nor U2163 (N_2163,N_2036,N_2076);
nand U2164 (N_2164,N_2075,N_2042);
nand U2165 (N_2165,N_2040,N_2061);
nor U2166 (N_2166,N_2002,N_2066);
or U2167 (N_2167,N_2085,N_2097);
or U2168 (N_2168,N_2081,N_2085);
nand U2169 (N_2169,N_2062,N_2036);
and U2170 (N_2170,N_2086,N_2017);
xor U2171 (N_2171,N_2073,N_2017);
nand U2172 (N_2172,N_2080,N_2048);
xor U2173 (N_2173,N_2091,N_2065);
nor U2174 (N_2174,N_2016,N_2000);
nand U2175 (N_2175,N_2086,N_2002);
nand U2176 (N_2176,N_2018,N_2093);
nor U2177 (N_2177,N_2082,N_2002);
nand U2178 (N_2178,N_2048,N_2036);
xor U2179 (N_2179,N_2023,N_2053);
xnor U2180 (N_2180,N_2072,N_2050);
nor U2181 (N_2181,N_2049,N_2043);
and U2182 (N_2182,N_2055,N_2091);
and U2183 (N_2183,N_2050,N_2084);
xnor U2184 (N_2184,N_2037,N_2068);
nand U2185 (N_2185,N_2055,N_2019);
nor U2186 (N_2186,N_2061,N_2009);
nor U2187 (N_2187,N_2030,N_2091);
nor U2188 (N_2188,N_2007,N_2087);
or U2189 (N_2189,N_2089,N_2009);
xor U2190 (N_2190,N_2095,N_2061);
xnor U2191 (N_2191,N_2077,N_2006);
or U2192 (N_2192,N_2040,N_2074);
xor U2193 (N_2193,N_2032,N_2082);
xor U2194 (N_2194,N_2045,N_2072);
nand U2195 (N_2195,N_2073,N_2052);
or U2196 (N_2196,N_2019,N_2075);
or U2197 (N_2197,N_2023,N_2082);
and U2198 (N_2198,N_2091,N_2039);
nand U2199 (N_2199,N_2001,N_2085);
nor U2200 (N_2200,N_2176,N_2103);
or U2201 (N_2201,N_2139,N_2149);
xor U2202 (N_2202,N_2152,N_2191);
nor U2203 (N_2203,N_2123,N_2146);
nor U2204 (N_2204,N_2117,N_2189);
xor U2205 (N_2205,N_2151,N_2153);
nand U2206 (N_2206,N_2195,N_2122);
nor U2207 (N_2207,N_2168,N_2194);
nor U2208 (N_2208,N_2101,N_2179);
nor U2209 (N_2209,N_2170,N_2129);
nand U2210 (N_2210,N_2142,N_2119);
nor U2211 (N_2211,N_2130,N_2133);
nor U2212 (N_2212,N_2184,N_2120);
xnor U2213 (N_2213,N_2127,N_2169);
or U2214 (N_2214,N_2166,N_2187);
and U2215 (N_2215,N_2134,N_2199);
or U2216 (N_2216,N_2155,N_2107);
nand U2217 (N_2217,N_2156,N_2147);
and U2218 (N_2218,N_2128,N_2197);
nand U2219 (N_2219,N_2118,N_2125);
and U2220 (N_2220,N_2150,N_2100);
and U2221 (N_2221,N_2173,N_2108);
and U2222 (N_2222,N_2190,N_2165);
xor U2223 (N_2223,N_2177,N_2132);
nor U2224 (N_2224,N_2102,N_2154);
nor U2225 (N_2225,N_2121,N_2126);
nor U2226 (N_2226,N_2115,N_2140);
and U2227 (N_2227,N_2110,N_2136);
and U2228 (N_2228,N_2180,N_2159);
or U2229 (N_2229,N_2158,N_2178);
xor U2230 (N_2230,N_2171,N_2131);
nand U2231 (N_2231,N_2193,N_2112);
xnor U2232 (N_2232,N_2172,N_2160);
or U2233 (N_2233,N_2196,N_2167);
nand U2234 (N_2234,N_2148,N_2192);
nor U2235 (N_2235,N_2174,N_2137);
nand U2236 (N_2236,N_2114,N_2188);
nor U2237 (N_2237,N_2106,N_2113);
nor U2238 (N_2238,N_2185,N_2141);
nand U2239 (N_2239,N_2138,N_2163);
or U2240 (N_2240,N_2181,N_2161);
xor U2241 (N_2241,N_2143,N_2116);
or U2242 (N_2242,N_2104,N_2111);
nand U2243 (N_2243,N_2175,N_2183);
or U2244 (N_2244,N_2198,N_2145);
or U2245 (N_2245,N_2144,N_2109);
and U2246 (N_2246,N_2164,N_2105);
nor U2247 (N_2247,N_2135,N_2157);
nand U2248 (N_2248,N_2186,N_2182);
xor U2249 (N_2249,N_2162,N_2124);
xor U2250 (N_2250,N_2124,N_2176);
xor U2251 (N_2251,N_2106,N_2140);
and U2252 (N_2252,N_2137,N_2188);
or U2253 (N_2253,N_2148,N_2100);
xnor U2254 (N_2254,N_2159,N_2151);
nor U2255 (N_2255,N_2189,N_2183);
xnor U2256 (N_2256,N_2162,N_2114);
nor U2257 (N_2257,N_2119,N_2184);
or U2258 (N_2258,N_2128,N_2182);
xnor U2259 (N_2259,N_2156,N_2168);
and U2260 (N_2260,N_2182,N_2115);
xor U2261 (N_2261,N_2142,N_2141);
nand U2262 (N_2262,N_2185,N_2136);
nand U2263 (N_2263,N_2118,N_2119);
xnor U2264 (N_2264,N_2195,N_2159);
nor U2265 (N_2265,N_2105,N_2144);
or U2266 (N_2266,N_2146,N_2101);
nand U2267 (N_2267,N_2125,N_2148);
or U2268 (N_2268,N_2125,N_2111);
or U2269 (N_2269,N_2149,N_2130);
or U2270 (N_2270,N_2126,N_2139);
xor U2271 (N_2271,N_2161,N_2166);
or U2272 (N_2272,N_2124,N_2148);
and U2273 (N_2273,N_2133,N_2148);
or U2274 (N_2274,N_2102,N_2110);
xnor U2275 (N_2275,N_2176,N_2137);
nor U2276 (N_2276,N_2158,N_2167);
and U2277 (N_2277,N_2125,N_2186);
nor U2278 (N_2278,N_2102,N_2166);
nor U2279 (N_2279,N_2168,N_2177);
nand U2280 (N_2280,N_2198,N_2180);
xnor U2281 (N_2281,N_2192,N_2119);
nor U2282 (N_2282,N_2124,N_2138);
nor U2283 (N_2283,N_2124,N_2131);
nand U2284 (N_2284,N_2171,N_2143);
and U2285 (N_2285,N_2100,N_2160);
and U2286 (N_2286,N_2127,N_2168);
xor U2287 (N_2287,N_2139,N_2147);
or U2288 (N_2288,N_2197,N_2133);
xnor U2289 (N_2289,N_2140,N_2189);
xnor U2290 (N_2290,N_2189,N_2157);
xnor U2291 (N_2291,N_2111,N_2129);
xnor U2292 (N_2292,N_2186,N_2165);
nor U2293 (N_2293,N_2151,N_2118);
nor U2294 (N_2294,N_2176,N_2199);
nor U2295 (N_2295,N_2156,N_2115);
or U2296 (N_2296,N_2193,N_2192);
nand U2297 (N_2297,N_2170,N_2109);
or U2298 (N_2298,N_2149,N_2185);
xor U2299 (N_2299,N_2120,N_2106);
xnor U2300 (N_2300,N_2244,N_2258);
nor U2301 (N_2301,N_2221,N_2202);
and U2302 (N_2302,N_2286,N_2245);
xnor U2303 (N_2303,N_2228,N_2238);
or U2304 (N_2304,N_2211,N_2247);
or U2305 (N_2305,N_2250,N_2257);
nor U2306 (N_2306,N_2227,N_2223);
or U2307 (N_2307,N_2290,N_2275);
xor U2308 (N_2308,N_2295,N_2246);
nor U2309 (N_2309,N_2253,N_2287);
and U2310 (N_2310,N_2251,N_2285);
xor U2311 (N_2311,N_2273,N_2237);
or U2312 (N_2312,N_2281,N_2270);
nor U2313 (N_2313,N_2222,N_2239);
or U2314 (N_2314,N_2259,N_2242);
or U2315 (N_2315,N_2214,N_2299);
or U2316 (N_2316,N_2274,N_2289);
nor U2317 (N_2317,N_2224,N_2208);
xor U2318 (N_2318,N_2230,N_2240);
nand U2319 (N_2319,N_2241,N_2262);
nor U2320 (N_2320,N_2296,N_2200);
nand U2321 (N_2321,N_2283,N_2206);
xnor U2322 (N_2322,N_2267,N_2272);
and U2323 (N_2323,N_2218,N_2280);
and U2324 (N_2324,N_2201,N_2215);
or U2325 (N_2325,N_2288,N_2209);
and U2326 (N_2326,N_2266,N_2232);
nand U2327 (N_2327,N_2271,N_2292);
or U2328 (N_2328,N_2212,N_2264);
or U2329 (N_2329,N_2203,N_2229);
or U2330 (N_2330,N_2210,N_2260);
and U2331 (N_2331,N_2265,N_2231);
xnor U2332 (N_2332,N_2219,N_2226);
nand U2333 (N_2333,N_2236,N_2207);
nor U2334 (N_2334,N_2233,N_2256);
xnor U2335 (N_2335,N_2254,N_2248);
xor U2336 (N_2336,N_2235,N_2205);
nor U2337 (N_2337,N_2282,N_2243);
nand U2338 (N_2338,N_2234,N_2293);
and U2339 (N_2339,N_2291,N_2217);
xor U2340 (N_2340,N_2276,N_2263);
or U2341 (N_2341,N_2216,N_2204);
and U2342 (N_2342,N_2249,N_2268);
xnor U2343 (N_2343,N_2261,N_2213);
nand U2344 (N_2344,N_2297,N_2298);
or U2345 (N_2345,N_2269,N_2284);
xor U2346 (N_2346,N_2252,N_2279);
nand U2347 (N_2347,N_2277,N_2225);
xor U2348 (N_2348,N_2294,N_2255);
and U2349 (N_2349,N_2278,N_2220);
xor U2350 (N_2350,N_2288,N_2219);
nor U2351 (N_2351,N_2213,N_2284);
nand U2352 (N_2352,N_2228,N_2294);
or U2353 (N_2353,N_2236,N_2230);
xnor U2354 (N_2354,N_2227,N_2243);
nor U2355 (N_2355,N_2258,N_2288);
nand U2356 (N_2356,N_2271,N_2277);
and U2357 (N_2357,N_2214,N_2208);
or U2358 (N_2358,N_2286,N_2228);
xor U2359 (N_2359,N_2240,N_2219);
or U2360 (N_2360,N_2248,N_2279);
or U2361 (N_2361,N_2271,N_2211);
or U2362 (N_2362,N_2273,N_2247);
or U2363 (N_2363,N_2270,N_2232);
and U2364 (N_2364,N_2259,N_2244);
and U2365 (N_2365,N_2249,N_2217);
nand U2366 (N_2366,N_2234,N_2209);
and U2367 (N_2367,N_2210,N_2296);
or U2368 (N_2368,N_2274,N_2213);
nor U2369 (N_2369,N_2222,N_2291);
or U2370 (N_2370,N_2212,N_2263);
nand U2371 (N_2371,N_2233,N_2232);
nand U2372 (N_2372,N_2260,N_2224);
or U2373 (N_2373,N_2284,N_2280);
or U2374 (N_2374,N_2225,N_2254);
nor U2375 (N_2375,N_2272,N_2201);
or U2376 (N_2376,N_2231,N_2229);
or U2377 (N_2377,N_2227,N_2244);
nand U2378 (N_2378,N_2229,N_2282);
or U2379 (N_2379,N_2228,N_2216);
nand U2380 (N_2380,N_2279,N_2250);
nor U2381 (N_2381,N_2230,N_2237);
xor U2382 (N_2382,N_2215,N_2214);
or U2383 (N_2383,N_2270,N_2259);
nand U2384 (N_2384,N_2268,N_2235);
xor U2385 (N_2385,N_2284,N_2271);
or U2386 (N_2386,N_2277,N_2275);
and U2387 (N_2387,N_2295,N_2244);
nand U2388 (N_2388,N_2203,N_2285);
xor U2389 (N_2389,N_2289,N_2210);
or U2390 (N_2390,N_2209,N_2284);
and U2391 (N_2391,N_2220,N_2272);
nand U2392 (N_2392,N_2254,N_2217);
nand U2393 (N_2393,N_2217,N_2219);
or U2394 (N_2394,N_2294,N_2245);
xnor U2395 (N_2395,N_2272,N_2286);
or U2396 (N_2396,N_2248,N_2200);
xnor U2397 (N_2397,N_2204,N_2268);
or U2398 (N_2398,N_2263,N_2288);
xor U2399 (N_2399,N_2261,N_2274);
nor U2400 (N_2400,N_2329,N_2369);
and U2401 (N_2401,N_2303,N_2358);
nand U2402 (N_2402,N_2399,N_2380);
xnor U2403 (N_2403,N_2379,N_2327);
nor U2404 (N_2404,N_2368,N_2345);
or U2405 (N_2405,N_2313,N_2364);
or U2406 (N_2406,N_2307,N_2316);
or U2407 (N_2407,N_2384,N_2397);
nor U2408 (N_2408,N_2301,N_2339);
nand U2409 (N_2409,N_2374,N_2365);
or U2410 (N_2410,N_2360,N_2342);
xnor U2411 (N_2411,N_2341,N_2322);
nand U2412 (N_2412,N_2347,N_2387);
or U2413 (N_2413,N_2393,N_2340);
nor U2414 (N_2414,N_2398,N_2337);
nand U2415 (N_2415,N_2315,N_2336);
and U2416 (N_2416,N_2382,N_2376);
or U2417 (N_2417,N_2330,N_2312);
xnor U2418 (N_2418,N_2324,N_2305);
and U2419 (N_2419,N_2356,N_2353);
and U2420 (N_2420,N_2325,N_2359);
and U2421 (N_2421,N_2388,N_2395);
nand U2422 (N_2422,N_2386,N_2318);
nor U2423 (N_2423,N_2300,N_2378);
or U2424 (N_2424,N_2302,N_2354);
nor U2425 (N_2425,N_2333,N_2343);
and U2426 (N_2426,N_2396,N_2331);
or U2427 (N_2427,N_2381,N_2335);
nand U2428 (N_2428,N_2314,N_2366);
and U2429 (N_2429,N_2308,N_2319);
nand U2430 (N_2430,N_2317,N_2311);
and U2431 (N_2431,N_2309,N_2372);
or U2432 (N_2432,N_2392,N_2362);
xnor U2433 (N_2433,N_2328,N_2352);
and U2434 (N_2434,N_2350,N_2383);
and U2435 (N_2435,N_2363,N_2349);
xor U2436 (N_2436,N_2348,N_2346);
and U2437 (N_2437,N_2389,N_2370);
xnor U2438 (N_2438,N_2390,N_2323);
nand U2439 (N_2439,N_2320,N_2357);
and U2440 (N_2440,N_2310,N_2344);
and U2441 (N_2441,N_2304,N_2391);
nand U2442 (N_2442,N_2385,N_2351);
xor U2443 (N_2443,N_2338,N_2332);
nor U2444 (N_2444,N_2334,N_2306);
nor U2445 (N_2445,N_2355,N_2375);
xnor U2446 (N_2446,N_2321,N_2373);
nand U2447 (N_2447,N_2361,N_2367);
xnor U2448 (N_2448,N_2326,N_2377);
or U2449 (N_2449,N_2394,N_2371);
xnor U2450 (N_2450,N_2328,N_2372);
and U2451 (N_2451,N_2322,N_2301);
nor U2452 (N_2452,N_2330,N_2307);
nand U2453 (N_2453,N_2338,N_2371);
nand U2454 (N_2454,N_2373,N_2338);
nor U2455 (N_2455,N_2378,N_2374);
and U2456 (N_2456,N_2389,N_2397);
nand U2457 (N_2457,N_2398,N_2396);
nor U2458 (N_2458,N_2398,N_2316);
and U2459 (N_2459,N_2315,N_2351);
or U2460 (N_2460,N_2380,N_2352);
xnor U2461 (N_2461,N_2362,N_2346);
and U2462 (N_2462,N_2325,N_2321);
xor U2463 (N_2463,N_2378,N_2377);
nand U2464 (N_2464,N_2310,N_2373);
or U2465 (N_2465,N_2353,N_2306);
nor U2466 (N_2466,N_2393,N_2343);
nand U2467 (N_2467,N_2311,N_2366);
xnor U2468 (N_2468,N_2380,N_2366);
or U2469 (N_2469,N_2300,N_2389);
xnor U2470 (N_2470,N_2390,N_2392);
xor U2471 (N_2471,N_2370,N_2393);
xnor U2472 (N_2472,N_2365,N_2321);
and U2473 (N_2473,N_2324,N_2370);
nor U2474 (N_2474,N_2387,N_2307);
or U2475 (N_2475,N_2324,N_2398);
nor U2476 (N_2476,N_2342,N_2302);
nand U2477 (N_2477,N_2378,N_2304);
and U2478 (N_2478,N_2350,N_2396);
nand U2479 (N_2479,N_2336,N_2330);
nand U2480 (N_2480,N_2383,N_2391);
nor U2481 (N_2481,N_2345,N_2364);
nand U2482 (N_2482,N_2362,N_2324);
nand U2483 (N_2483,N_2341,N_2308);
nor U2484 (N_2484,N_2322,N_2328);
nor U2485 (N_2485,N_2399,N_2302);
and U2486 (N_2486,N_2359,N_2334);
and U2487 (N_2487,N_2389,N_2321);
and U2488 (N_2488,N_2369,N_2309);
nand U2489 (N_2489,N_2316,N_2326);
and U2490 (N_2490,N_2381,N_2325);
nand U2491 (N_2491,N_2339,N_2358);
nand U2492 (N_2492,N_2331,N_2364);
nand U2493 (N_2493,N_2313,N_2388);
or U2494 (N_2494,N_2326,N_2300);
nand U2495 (N_2495,N_2392,N_2308);
and U2496 (N_2496,N_2317,N_2310);
nand U2497 (N_2497,N_2307,N_2372);
xnor U2498 (N_2498,N_2329,N_2382);
xor U2499 (N_2499,N_2302,N_2303);
nand U2500 (N_2500,N_2414,N_2493);
nand U2501 (N_2501,N_2451,N_2489);
nand U2502 (N_2502,N_2450,N_2448);
or U2503 (N_2503,N_2444,N_2485);
nor U2504 (N_2504,N_2492,N_2496);
nor U2505 (N_2505,N_2484,N_2436);
or U2506 (N_2506,N_2438,N_2467);
nor U2507 (N_2507,N_2473,N_2410);
xor U2508 (N_2508,N_2432,N_2446);
or U2509 (N_2509,N_2400,N_2461);
nand U2510 (N_2510,N_2417,N_2482);
xnor U2511 (N_2511,N_2404,N_2402);
nand U2512 (N_2512,N_2457,N_2477);
xnor U2513 (N_2513,N_2491,N_2463);
nand U2514 (N_2514,N_2474,N_2415);
xor U2515 (N_2515,N_2453,N_2434);
nand U2516 (N_2516,N_2406,N_2460);
and U2517 (N_2517,N_2431,N_2418);
xnor U2518 (N_2518,N_2483,N_2405);
and U2519 (N_2519,N_2426,N_2464);
nand U2520 (N_2520,N_2428,N_2425);
nand U2521 (N_2521,N_2490,N_2433);
xor U2522 (N_2522,N_2455,N_2435);
and U2523 (N_2523,N_2494,N_2440);
and U2524 (N_2524,N_2470,N_2447);
nand U2525 (N_2525,N_2462,N_2480);
or U2526 (N_2526,N_2421,N_2495);
nor U2527 (N_2527,N_2443,N_2413);
and U2528 (N_2528,N_2499,N_2469);
nand U2529 (N_2529,N_2407,N_2481);
nand U2530 (N_2530,N_2459,N_2456);
nand U2531 (N_2531,N_2449,N_2437);
nand U2532 (N_2532,N_2479,N_2430);
xnor U2533 (N_2533,N_2424,N_2486);
nand U2534 (N_2534,N_2478,N_2487);
or U2535 (N_2535,N_2420,N_2416);
xor U2536 (N_2536,N_2442,N_2476);
and U2537 (N_2537,N_2497,N_2409);
xor U2538 (N_2538,N_2466,N_2471);
nor U2539 (N_2539,N_2475,N_2439);
or U2540 (N_2540,N_2419,N_2408);
xor U2541 (N_2541,N_2411,N_2429);
or U2542 (N_2542,N_2498,N_2445);
xor U2543 (N_2543,N_2427,N_2472);
xnor U2544 (N_2544,N_2488,N_2423);
xnor U2545 (N_2545,N_2468,N_2454);
and U2546 (N_2546,N_2465,N_2441);
xnor U2547 (N_2547,N_2403,N_2422);
and U2548 (N_2548,N_2412,N_2458);
and U2549 (N_2549,N_2452,N_2401);
and U2550 (N_2550,N_2479,N_2431);
nor U2551 (N_2551,N_2426,N_2492);
and U2552 (N_2552,N_2423,N_2460);
nand U2553 (N_2553,N_2462,N_2425);
nor U2554 (N_2554,N_2454,N_2407);
nand U2555 (N_2555,N_2493,N_2443);
xnor U2556 (N_2556,N_2413,N_2460);
nand U2557 (N_2557,N_2465,N_2463);
nor U2558 (N_2558,N_2405,N_2442);
nor U2559 (N_2559,N_2463,N_2475);
nand U2560 (N_2560,N_2463,N_2400);
or U2561 (N_2561,N_2412,N_2424);
xor U2562 (N_2562,N_2432,N_2481);
nand U2563 (N_2563,N_2400,N_2424);
nor U2564 (N_2564,N_2437,N_2468);
and U2565 (N_2565,N_2409,N_2445);
xnor U2566 (N_2566,N_2483,N_2429);
and U2567 (N_2567,N_2493,N_2412);
xnor U2568 (N_2568,N_2458,N_2465);
xor U2569 (N_2569,N_2433,N_2497);
nor U2570 (N_2570,N_2413,N_2418);
or U2571 (N_2571,N_2453,N_2417);
or U2572 (N_2572,N_2478,N_2470);
and U2573 (N_2573,N_2410,N_2418);
nand U2574 (N_2574,N_2469,N_2466);
or U2575 (N_2575,N_2429,N_2461);
nand U2576 (N_2576,N_2470,N_2441);
and U2577 (N_2577,N_2495,N_2447);
xnor U2578 (N_2578,N_2430,N_2465);
xnor U2579 (N_2579,N_2499,N_2484);
or U2580 (N_2580,N_2480,N_2449);
and U2581 (N_2581,N_2486,N_2460);
nand U2582 (N_2582,N_2414,N_2416);
nand U2583 (N_2583,N_2487,N_2495);
xnor U2584 (N_2584,N_2462,N_2486);
or U2585 (N_2585,N_2491,N_2476);
or U2586 (N_2586,N_2489,N_2492);
xnor U2587 (N_2587,N_2476,N_2468);
or U2588 (N_2588,N_2431,N_2466);
xor U2589 (N_2589,N_2482,N_2420);
nand U2590 (N_2590,N_2481,N_2449);
xor U2591 (N_2591,N_2415,N_2423);
xor U2592 (N_2592,N_2427,N_2413);
nand U2593 (N_2593,N_2487,N_2427);
nand U2594 (N_2594,N_2411,N_2474);
or U2595 (N_2595,N_2488,N_2478);
or U2596 (N_2596,N_2469,N_2462);
nor U2597 (N_2597,N_2444,N_2430);
xnor U2598 (N_2598,N_2420,N_2432);
and U2599 (N_2599,N_2442,N_2431);
nand U2600 (N_2600,N_2526,N_2536);
or U2601 (N_2601,N_2525,N_2542);
xnor U2602 (N_2602,N_2566,N_2510);
or U2603 (N_2603,N_2593,N_2559);
nor U2604 (N_2604,N_2550,N_2595);
or U2605 (N_2605,N_2544,N_2569);
nand U2606 (N_2606,N_2583,N_2531);
nand U2607 (N_2607,N_2557,N_2578);
xor U2608 (N_2608,N_2560,N_2534);
nand U2609 (N_2609,N_2565,N_2570);
and U2610 (N_2610,N_2543,N_2574);
or U2611 (N_2611,N_2521,N_2573);
or U2612 (N_2612,N_2571,N_2585);
and U2613 (N_2613,N_2532,N_2556);
xor U2614 (N_2614,N_2572,N_2512);
xor U2615 (N_2615,N_2515,N_2505);
and U2616 (N_2616,N_2501,N_2540);
nor U2617 (N_2617,N_2568,N_2586);
nor U2618 (N_2618,N_2517,N_2598);
or U2619 (N_2619,N_2529,N_2592);
or U2620 (N_2620,N_2551,N_2514);
or U2621 (N_2621,N_2504,N_2558);
and U2622 (N_2622,N_2513,N_2554);
or U2623 (N_2623,N_2528,N_2527);
xor U2624 (N_2624,N_2508,N_2503);
or U2625 (N_2625,N_2575,N_2577);
and U2626 (N_2626,N_2530,N_2576);
nand U2627 (N_2627,N_2507,N_2594);
nand U2628 (N_2628,N_2590,N_2502);
and U2629 (N_2629,N_2509,N_2549);
or U2630 (N_2630,N_2516,N_2541);
or U2631 (N_2631,N_2555,N_2519);
xnor U2632 (N_2632,N_2587,N_2547);
xor U2633 (N_2633,N_2581,N_2537);
nand U2634 (N_2634,N_2582,N_2539);
nand U2635 (N_2635,N_2546,N_2596);
xor U2636 (N_2636,N_2548,N_2562);
xnor U2637 (N_2637,N_2561,N_2563);
nor U2638 (N_2638,N_2591,N_2580);
nand U2639 (N_2639,N_2506,N_2500);
xor U2640 (N_2640,N_2535,N_2584);
and U2641 (N_2641,N_2533,N_2567);
or U2642 (N_2642,N_2524,N_2597);
or U2643 (N_2643,N_2538,N_2522);
xor U2644 (N_2644,N_2599,N_2588);
or U2645 (N_2645,N_2523,N_2545);
and U2646 (N_2646,N_2589,N_2553);
and U2647 (N_2647,N_2520,N_2564);
or U2648 (N_2648,N_2518,N_2552);
nor U2649 (N_2649,N_2511,N_2579);
nand U2650 (N_2650,N_2566,N_2588);
nor U2651 (N_2651,N_2503,N_2558);
nor U2652 (N_2652,N_2536,N_2577);
and U2653 (N_2653,N_2534,N_2515);
and U2654 (N_2654,N_2577,N_2544);
and U2655 (N_2655,N_2563,N_2549);
or U2656 (N_2656,N_2507,N_2561);
or U2657 (N_2657,N_2581,N_2533);
nor U2658 (N_2658,N_2548,N_2513);
nor U2659 (N_2659,N_2504,N_2557);
and U2660 (N_2660,N_2529,N_2591);
xnor U2661 (N_2661,N_2530,N_2582);
nand U2662 (N_2662,N_2539,N_2551);
xor U2663 (N_2663,N_2517,N_2508);
nor U2664 (N_2664,N_2547,N_2556);
nand U2665 (N_2665,N_2509,N_2534);
nor U2666 (N_2666,N_2537,N_2508);
nand U2667 (N_2667,N_2546,N_2537);
nand U2668 (N_2668,N_2564,N_2505);
nor U2669 (N_2669,N_2521,N_2500);
nor U2670 (N_2670,N_2525,N_2554);
nand U2671 (N_2671,N_2571,N_2520);
nand U2672 (N_2672,N_2574,N_2565);
and U2673 (N_2673,N_2500,N_2585);
and U2674 (N_2674,N_2514,N_2584);
or U2675 (N_2675,N_2552,N_2547);
nand U2676 (N_2676,N_2579,N_2516);
nand U2677 (N_2677,N_2506,N_2524);
xor U2678 (N_2678,N_2599,N_2511);
nor U2679 (N_2679,N_2524,N_2563);
xnor U2680 (N_2680,N_2578,N_2522);
and U2681 (N_2681,N_2533,N_2561);
nor U2682 (N_2682,N_2578,N_2565);
or U2683 (N_2683,N_2575,N_2566);
nor U2684 (N_2684,N_2516,N_2501);
nor U2685 (N_2685,N_2559,N_2561);
xnor U2686 (N_2686,N_2597,N_2575);
nor U2687 (N_2687,N_2521,N_2502);
nand U2688 (N_2688,N_2537,N_2554);
or U2689 (N_2689,N_2581,N_2526);
nor U2690 (N_2690,N_2591,N_2598);
or U2691 (N_2691,N_2538,N_2571);
xor U2692 (N_2692,N_2555,N_2508);
or U2693 (N_2693,N_2548,N_2540);
and U2694 (N_2694,N_2560,N_2550);
xnor U2695 (N_2695,N_2525,N_2515);
nor U2696 (N_2696,N_2549,N_2528);
nor U2697 (N_2697,N_2564,N_2559);
xnor U2698 (N_2698,N_2595,N_2546);
nand U2699 (N_2699,N_2507,N_2540);
nor U2700 (N_2700,N_2667,N_2619);
nor U2701 (N_2701,N_2639,N_2626);
and U2702 (N_2702,N_2649,N_2607);
xnor U2703 (N_2703,N_2652,N_2615);
nor U2704 (N_2704,N_2664,N_2629);
nor U2705 (N_2705,N_2681,N_2697);
nand U2706 (N_2706,N_2687,N_2631);
xnor U2707 (N_2707,N_2668,N_2658);
and U2708 (N_2708,N_2647,N_2684);
or U2709 (N_2709,N_2654,N_2601);
and U2710 (N_2710,N_2611,N_2641);
nor U2711 (N_2711,N_2699,N_2644);
nor U2712 (N_2712,N_2640,N_2600);
and U2713 (N_2713,N_2692,N_2624);
nor U2714 (N_2714,N_2653,N_2636);
nor U2715 (N_2715,N_2674,N_2650);
and U2716 (N_2716,N_2665,N_2645);
xnor U2717 (N_2717,N_2620,N_2691);
nand U2718 (N_2718,N_2693,N_2623);
nor U2719 (N_2719,N_2646,N_2695);
xor U2720 (N_2720,N_2686,N_2632);
xor U2721 (N_2721,N_2633,N_2659);
xnor U2722 (N_2722,N_2696,N_2672);
xnor U2723 (N_2723,N_2662,N_2606);
nand U2724 (N_2724,N_2630,N_2679);
nor U2725 (N_2725,N_2618,N_2613);
or U2726 (N_2726,N_2694,N_2643);
nand U2727 (N_2727,N_2671,N_2660);
or U2728 (N_2728,N_2682,N_2698);
nand U2729 (N_2729,N_2602,N_2617);
xnor U2730 (N_2730,N_2635,N_2680);
nand U2731 (N_2731,N_2609,N_2638);
xor U2732 (N_2732,N_2614,N_2637);
or U2733 (N_2733,N_2675,N_2612);
and U2734 (N_2734,N_2628,N_2677);
and U2735 (N_2735,N_2616,N_2634);
or U2736 (N_2736,N_2678,N_2604);
or U2737 (N_2737,N_2648,N_2683);
and U2738 (N_2738,N_2670,N_2685);
nand U2739 (N_2739,N_2688,N_2608);
and U2740 (N_2740,N_2642,N_2690);
nor U2741 (N_2741,N_2651,N_2655);
xnor U2742 (N_2742,N_2656,N_2676);
and U2743 (N_2743,N_2673,N_2669);
xor U2744 (N_2744,N_2621,N_2627);
and U2745 (N_2745,N_2622,N_2663);
xnor U2746 (N_2746,N_2661,N_2605);
xor U2747 (N_2747,N_2657,N_2603);
nand U2748 (N_2748,N_2610,N_2666);
nor U2749 (N_2749,N_2625,N_2689);
xor U2750 (N_2750,N_2602,N_2673);
or U2751 (N_2751,N_2642,N_2698);
xnor U2752 (N_2752,N_2649,N_2674);
xnor U2753 (N_2753,N_2626,N_2660);
xnor U2754 (N_2754,N_2628,N_2652);
nor U2755 (N_2755,N_2684,N_2691);
xor U2756 (N_2756,N_2601,N_2688);
nor U2757 (N_2757,N_2609,N_2669);
or U2758 (N_2758,N_2659,N_2684);
xnor U2759 (N_2759,N_2643,N_2681);
nand U2760 (N_2760,N_2655,N_2663);
xor U2761 (N_2761,N_2641,N_2660);
nand U2762 (N_2762,N_2685,N_2620);
xor U2763 (N_2763,N_2608,N_2698);
or U2764 (N_2764,N_2645,N_2699);
and U2765 (N_2765,N_2657,N_2679);
nand U2766 (N_2766,N_2646,N_2612);
nand U2767 (N_2767,N_2628,N_2679);
xor U2768 (N_2768,N_2673,N_2620);
and U2769 (N_2769,N_2654,N_2681);
nand U2770 (N_2770,N_2662,N_2654);
nor U2771 (N_2771,N_2645,N_2601);
nand U2772 (N_2772,N_2631,N_2667);
or U2773 (N_2773,N_2683,N_2659);
nand U2774 (N_2774,N_2671,N_2620);
nor U2775 (N_2775,N_2610,N_2693);
nor U2776 (N_2776,N_2675,N_2635);
and U2777 (N_2777,N_2649,N_2634);
xor U2778 (N_2778,N_2635,N_2661);
and U2779 (N_2779,N_2684,N_2624);
nor U2780 (N_2780,N_2677,N_2652);
nand U2781 (N_2781,N_2647,N_2657);
and U2782 (N_2782,N_2682,N_2699);
or U2783 (N_2783,N_2687,N_2677);
nor U2784 (N_2784,N_2684,N_2688);
nor U2785 (N_2785,N_2698,N_2639);
nor U2786 (N_2786,N_2605,N_2639);
or U2787 (N_2787,N_2608,N_2638);
or U2788 (N_2788,N_2678,N_2628);
nand U2789 (N_2789,N_2639,N_2664);
xnor U2790 (N_2790,N_2681,N_2621);
xnor U2791 (N_2791,N_2618,N_2657);
and U2792 (N_2792,N_2637,N_2694);
nor U2793 (N_2793,N_2679,N_2683);
or U2794 (N_2794,N_2673,N_2608);
nor U2795 (N_2795,N_2668,N_2620);
and U2796 (N_2796,N_2654,N_2659);
and U2797 (N_2797,N_2620,N_2649);
xor U2798 (N_2798,N_2636,N_2606);
nand U2799 (N_2799,N_2698,N_2693);
nor U2800 (N_2800,N_2782,N_2719);
and U2801 (N_2801,N_2781,N_2712);
or U2802 (N_2802,N_2730,N_2706);
and U2803 (N_2803,N_2727,N_2756);
or U2804 (N_2804,N_2731,N_2724);
nor U2805 (N_2805,N_2745,N_2784);
xor U2806 (N_2806,N_2790,N_2737);
and U2807 (N_2807,N_2762,N_2794);
or U2808 (N_2808,N_2700,N_2789);
or U2809 (N_2809,N_2760,N_2726);
nor U2810 (N_2810,N_2735,N_2715);
and U2811 (N_2811,N_2744,N_2702);
xnor U2812 (N_2812,N_2777,N_2716);
nand U2813 (N_2813,N_2798,N_2732);
or U2814 (N_2814,N_2766,N_2775);
nor U2815 (N_2815,N_2711,N_2793);
and U2816 (N_2816,N_2739,N_2768);
nor U2817 (N_2817,N_2718,N_2701);
or U2818 (N_2818,N_2796,N_2738);
and U2819 (N_2819,N_2780,N_2758);
and U2820 (N_2820,N_2786,N_2795);
and U2821 (N_2821,N_2788,N_2787);
nand U2822 (N_2822,N_2753,N_2703);
and U2823 (N_2823,N_2722,N_2748);
nor U2824 (N_2824,N_2710,N_2792);
nand U2825 (N_2825,N_2723,N_2774);
or U2826 (N_2826,N_2799,N_2763);
and U2827 (N_2827,N_2704,N_2765);
nor U2828 (N_2828,N_2720,N_2714);
nor U2829 (N_2829,N_2708,N_2733);
or U2830 (N_2830,N_2769,N_2742);
nand U2831 (N_2831,N_2725,N_2771);
nand U2832 (N_2832,N_2783,N_2755);
and U2833 (N_2833,N_2751,N_2707);
and U2834 (N_2834,N_2728,N_2736);
nor U2835 (N_2835,N_2750,N_2717);
nor U2836 (N_2836,N_2749,N_2773);
and U2837 (N_2837,N_2778,N_2752);
and U2838 (N_2838,N_2767,N_2721);
nor U2839 (N_2839,N_2709,N_2791);
and U2840 (N_2840,N_2759,N_2797);
nand U2841 (N_2841,N_2743,N_2776);
nor U2842 (N_2842,N_2740,N_2734);
nand U2843 (N_2843,N_2770,N_2772);
or U2844 (N_2844,N_2785,N_2754);
nor U2845 (N_2845,N_2705,N_2713);
nand U2846 (N_2846,N_2779,N_2761);
nor U2847 (N_2847,N_2757,N_2741);
and U2848 (N_2848,N_2746,N_2729);
xor U2849 (N_2849,N_2747,N_2764);
nand U2850 (N_2850,N_2705,N_2747);
nor U2851 (N_2851,N_2718,N_2770);
nor U2852 (N_2852,N_2713,N_2711);
or U2853 (N_2853,N_2743,N_2730);
nand U2854 (N_2854,N_2703,N_2726);
nor U2855 (N_2855,N_2799,N_2724);
and U2856 (N_2856,N_2765,N_2787);
xor U2857 (N_2857,N_2721,N_2709);
or U2858 (N_2858,N_2767,N_2712);
nor U2859 (N_2859,N_2784,N_2767);
or U2860 (N_2860,N_2735,N_2718);
nor U2861 (N_2861,N_2797,N_2773);
or U2862 (N_2862,N_2710,N_2744);
xor U2863 (N_2863,N_2782,N_2715);
and U2864 (N_2864,N_2744,N_2711);
nor U2865 (N_2865,N_2717,N_2748);
nand U2866 (N_2866,N_2707,N_2786);
and U2867 (N_2867,N_2756,N_2752);
xnor U2868 (N_2868,N_2725,N_2774);
nand U2869 (N_2869,N_2745,N_2780);
or U2870 (N_2870,N_2743,N_2799);
and U2871 (N_2871,N_2798,N_2740);
or U2872 (N_2872,N_2704,N_2762);
and U2873 (N_2873,N_2752,N_2784);
or U2874 (N_2874,N_2707,N_2749);
nand U2875 (N_2875,N_2747,N_2787);
and U2876 (N_2876,N_2769,N_2723);
nor U2877 (N_2877,N_2729,N_2701);
or U2878 (N_2878,N_2713,N_2735);
or U2879 (N_2879,N_2760,N_2707);
and U2880 (N_2880,N_2715,N_2703);
nand U2881 (N_2881,N_2730,N_2722);
nor U2882 (N_2882,N_2795,N_2774);
or U2883 (N_2883,N_2792,N_2796);
and U2884 (N_2884,N_2709,N_2788);
xnor U2885 (N_2885,N_2783,N_2752);
nand U2886 (N_2886,N_2729,N_2713);
or U2887 (N_2887,N_2707,N_2729);
or U2888 (N_2888,N_2761,N_2784);
and U2889 (N_2889,N_2749,N_2735);
xnor U2890 (N_2890,N_2711,N_2756);
or U2891 (N_2891,N_2785,N_2720);
xor U2892 (N_2892,N_2736,N_2749);
nor U2893 (N_2893,N_2712,N_2760);
nand U2894 (N_2894,N_2789,N_2768);
nor U2895 (N_2895,N_2703,N_2717);
xor U2896 (N_2896,N_2706,N_2729);
or U2897 (N_2897,N_2786,N_2790);
nand U2898 (N_2898,N_2724,N_2797);
and U2899 (N_2899,N_2766,N_2701);
or U2900 (N_2900,N_2824,N_2874);
and U2901 (N_2901,N_2837,N_2846);
xor U2902 (N_2902,N_2892,N_2879);
nand U2903 (N_2903,N_2881,N_2855);
nor U2904 (N_2904,N_2834,N_2840);
nand U2905 (N_2905,N_2872,N_2864);
and U2906 (N_2906,N_2889,N_2868);
and U2907 (N_2907,N_2876,N_2826);
nor U2908 (N_2908,N_2807,N_2829);
nor U2909 (N_2909,N_2818,N_2812);
nand U2910 (N_2910,N_2827,N_2811);
xor U2911 (N_2911,N_2894,N_2899);
xnor U2912 (N_2912,N_2852,N_2884);
nand U2913 (N_2913,N_2803,N_2820);
nand U2914 (N_2914,N_2853,N_2817);
xnor U2915 (N_2915,N_2861,N_2804);
or U2916 (N_2916,N_2886,N_2869);
nor U2917 (N_2917,N_2823,N_2828);
and U2918 (N_2918,N_2841,N_2810);
nor U2919 (N_2919,N_2887,N_2814);
xnor U2920 (N_2920,N_2821,N_2833);
nand U2921 (N_2921,N_2893,N_2862);
nand U2922 (N_2922,N_2805,N_2860);
or U2923 (N_2923,N_2867,N_2842);
nand U2924 (N_2924,N_2815,N_2865);
xor U2925 (N_2925,N_2858,N_2843);
or U2926 (N_2926,N_2830,N_2801);
or U2927 (N_2927,N_2898,N_2848);
nand U2928 (N_2928,N_2870,N_2822);
and U2929 (N_2929,N_2835,N_2854);
nand U2930 (N_2930,N_2806,N_2825);
and U2931 (N_2931,N_2890,N_2885);
nand U2932 (N_2932,N_2897,N_2850);
nor U2933 (N_2933,N_2866,N_2819);
nand U2934 (N_2934,N_2863,N_2802);
nor U2935 (N_2935,N_2888,N_2896);
xnor U2936 (N_2936,N_2878,N_2808);
or U2937 (N_2937,N_2883,N_2831);
or U2938 (N_2938,N_2895,N_2832);
nor U2939 (N_2939,N_2838,N_2816);
or U2940 (N_2940,N_2845,N_2800);
xor U2941 (N_2941,N_2839,N_2844);
or U2942 (N_2942,N_2836,N_2859);
xnor U2943 (N_2943,N_2857,N_2891);
and U2944 (N_2944,N_2849,N_2875);
and U2945 (N_2945,N_2877,N_2873);
or U2946 (N_2946,N_2847,N_2856);
and U2947 (N_2947,N_2880,N_2813);
xor U2948 (N_2948,N_2851,N_2882);
and U2949 (N_2949,N_2809,N_2871);
nor U2950 (N_2950,N_2899,N_2823);
or U2951 (N_2951,N_2894,N_2890);
or U2952 (N_2952,N_2859,N_2864);
nand U2953 (N_2953,N_2833,N_2825);
or U2954 (N_2954,N_2855,N_2828);
nand U2955 (N_2955,N_2809,N_2810);
nor U2956 (N_2956,N_2892,N_2891);
and U2957 (N_2957,N_2811,N_2801);
nand U2958 (N_2958,N_2858,N_2876);
or U2959 (N_2959,N_2837,N_2860);
nand U2960 (N_2960,N_2855,N_2836);
or U2961 (N_2961,N_2888,N_2878);
xnor U2962 (N_2962,N_2894,N_2821);
and U2963 (N_2963,N_2890,N_2865);
nand U2964 (N_2964,N_2846,N_2838);
and U2965 (N_2965,N_2874,N_2870);
and U2966 (N_2966,N_2891,N_2885);
nor U2967 (N_2967,N_2879,N_2852);
nor U2968 (N_2968,N_2814,N_2882);
nand U2969 (N_2969,N_2840,N_2865);
and U2970 (N_2970,N_2821,N_2876);
nor U2971 (N_2971,N_2806,N_2805);
nand U2972 (N_2972,N_2896,N_2805);
nand U2973 (N_2973,N_2840,N_2831);
nor U2974 (N_2974,N_2817,N_2818);
xor U2975 (N_2975,N_2867,N_2872);
nand U2976 (N_2976,N_2871,N_2881);
and U2977 (N_2977,N_2841,N_2814);
nor U2978 (N_2978,N_2806,N_2824);
nand U2979 (N_2979,N_2822,N_2840);
xor U2980 (N_2980,N_2890,N_2827);
nand U2981 (N_2981,N_2899,N_2830);
and U2982 (N_2982,N_2800,N_2838);
or U2983 (N_2983,N_2850,N_2813);
and U2984 (N_2984,N_2831,N_2882);
or U2985 (N_2985,N_2857,N_2881);
nor U2986 (N_2986,N_2884,N_2837);
and U2987 (N_2987,N_2823,N_2873);
xor U2988 (N_2988,N_2884,N_2839);
nand U2989 (N_2989,N_2861,N_2825);
and U2990 (N_2990,N_2838,N_2889);
nand U2991 (N_2991,N_2894,N_2867);
xnor U2992 (N_2992,N_2897,N_2887);
or U2993 (N_2993,N_2877,N_2849);
nand U2994 (N_2994,N_2885,N_2860);
and U2995 (N_2995,N_2886,N_2829);
and U2996 (N_2996,N_2873,N_2884);
and U2997 (N_2997,N_2876,N_2804);
nor U2998 (N_2998,N_2826,N_2867);
nor U2999 (N_2999,N_2836,N_2834);
xnor U3000 (N_3000,N_2960,N_2991);
and U3001 (N_3001,N_2989,N_2909);
nor U3002 (N_3002,N_2918,N_2969);
nor U3003 (N_3003,N_2975,N_2906);
and U3004 (N_3004,N_2964,N_2919);
and U3005 (N_3005,N_2924,N_2993);
and U3006 (N_3006,N_2914,N_2911);
and U3007 (N_3007,N_2998,N_2913);
nor U3008 (N_3008,N_2979,N_2940);
xor U3009 (N_3009,N_2937,N_2957);
xor U3010 (N_3010,N_2954,N_2970);
xnor U3011 (N_3011,N_2965,N_2936);
nand U3012 (N_3012,N_2944,N_2902);
nand U3013 (N_3013,N_2955,N_2903);
xor U3014 (N_3014,N_2928,N_2927);
xor U3015 (N_3015,N_2976,N_2981);
xor U3016 (N_3016,N_2932,N_2967);
and U3017 (N_3017,N_2982,N_2922);
nand U3018 (N_3018,N_2997,N_2904);
nand U3019 (N_3019,N_2956,N_2930);
xnor U3020 (N_3020,N_2963,N_2987);
xor U3021 (N_3021,N_2941,N_2916);
nor U3022 (N_3022,N_2945,N_2961);
nor U3023 (N_3023,N_2947,N_2905);
or U3024 (N_3024,N_2910,N_2948);
nand U3025 (N_3025,N_2929,N_2939);
nor U3026 (N_3026,N_2953,N_2950);
and U3027 (N_3027,N_2952,N_2920);
and U3028 (N_3028,N_2934,N_2925);
or U3029 (N_3029,N_2966,N_2951);
or U3030 (N_3030,N_2977,N_2959);
and U3031 (N_3031,N_2921,N_2943);
and U3032 (N_3032,N_2994,N_2908);
nor U3033 (N_3033,N_2971,N_2915);
and U3034 (N_3034,N_2995,N_2958);
and U3035 (N_3035,N_2984,N_2935);
and U3036 (N_3036,N_2972,N_2938);
or U3037 (N_3037,N_2968,N_2985);
nand U3038 (N_3038,N_2912,N_2907);
nor U3039 (N_3039,N_2901,N_2946);
xnor U3040 (N_3040,N_2974,N_2942);
or U3041 (N_3041,N_2962,N_2988);
and U3042 (N_3042,N_2923,N_2992);
nor U3043 (N_3043,N_2917,N_2931);
xor U3044 (N_3044,N_2986,N_2980);
nand U3045 (N_3045,N_2999,N_2926);
or U3046 (N_3046,N_2973,N_2990);
nor U3047 (N_3047,N_2949,N_2983);
or U3048 (N_3048,N_2996,N_2978);
nand U3049 (N_3049,N_2900,N_2933);
nor U3050 (N_3050,N_2957,N_2955);
nand U3051 (N_3051,N_2948,N_2903);
or U3052 (N_3052,N_2948,N_2933);
nor U3053 (N_3053,N_2954,N_2936);
xor U3054 (N_3054,N_2977,N_2978);
xor U3055 (N_3055,N_2971,N_2962);
xor U3056 (N_3056,N_2975,N_2981);
xnor U3057 (N_3057,N_2990,N_2923);
xnor U3058 (N_3058,N_2973,N_2923);
or U3059 (N_3059,N_2967,N_2942);
nand U3060 (N_3060,N_2986,N_2958);
and U3061 (N_3061,N_2927,N_2920);
or U3062 (N_3062,N_2904,N_2921);
nor U3063 (N_3063,N_2949,N_2974);
xnor U3064 (N_3064,N_2970,N_2913);
nand U3065 (N_3065,N_2900,N_2913);
nor U3066 (N_3066,N_2902,N_2931);
xnor U3067 (N_3067,N_2919,N_2985);
nor U3068 (N_3068,N_2939,N_2915);
xnor U3069 (N_3069,N_2998,N_2936);
or U3070 (N_3070,N_2992,N_2920);
nand U3071 (N_3071,N_2939,N_2928);
or U3072 (N_3072,N_2919,N_2917);
nor U3073 (N_3073,N_2923,N_2905);
nor U3074 (N_3074,N_2964,N_2953);
xor U3075 (N_3075,N_2951,N_2958);
nor U3076 (N_3076,N_2964,N_2944);
or U3077 (N_3077,N_2986,N_2942);
or U3078 (N_3078,N_2933,N_2911);
and U3079 (N_3079,N_2905,N_2989);
nand U3080 (N_3080,N_2977,N_2994);
or U3081 (N_3081,N_2944,N_2965);
xnor U3082 (N_3082,N_2990,N_2993);
and U3083 (N_3083,N_2969,N_2939);
nor U3084 (N_3084,N_2967,N_2930);
nor U3085 (N_3085,N_2907,N_2945);
or U3086 (N_3086,N_2938,N_2983);
or U3087 (N_3087,N_2963,N_2960);
xnor U3088 (N_3088,N_2925,N_2947);
nor U3089 (N_3089,N_2910,N_2932);
xnor U3090 (N_3090,N_2986,N_2944);
xnor U3091 (N_3091,N_2946,N_2934);
or U3092 (N_3092,N_2972,N_2904);
xor U3093 (N_3093,N_2989,N_2903);
or U3094 (N_3094,N_2938,N_2921);
nand U3095 (N_3095,N_2932,N_2930);
xor U3096 (N_3096,N_2951,N_2911);
xor U3097 (N_3097,N_2978,N_2970);
or U3098 (N_3098,N_2929,N_2949);
nor U3099 (N_3099,N_2906,N_2951);
nor U3100 (N_3100,N_3084,N_3042);
nor U3101 (N_3101,N_3023,N_3097);
xor U3102 (N_3102,N_3028,N_3096);
nand U3103 (N_3103,N_3046,N_3006);
and U3104 (N_3104,N_3082,N_3019);
nor U3105 (N_3105,N_3098,N_3031);
or U3106 (N_3106,N_3061,N_3037);
and U3107 (N_3107,N_3045,N_3015);
and U3108 (N_3108,N_3029,N_3020);
nor U3109 (N_3109,N_3086,N_3052);
nand U3110 (N_3110,N_3074,N_3094);
or U3111 (N_3111,N_3051,N_3000);
nor U3112 (N_3112,N_3007,N_3071);
xnor U3113 (N_3113,N_3036,N_3053);
nor U3114 (N_3114,N_3022,N_3054);
nor U3115 (N_3115,N_3058,N_3057);
xor U3116 (N_3116,N_3091,N_3002);
nand U3117 (N_3117,N_3089,N_3034);
xnor U3118 (N_3118,N_3055,N_3050);
xnor U3119 (N_3119,N_3008,N_3044);
or U3120 (N_3120,N_3069,N_3012);
nor U3121 (N_3121,N_3027,N_3014);
or U3122 (N_3122,N_3041,N_3067);
and U3123 (N_3123,N_3077,N_3026);
or U3124 (N_3124,N_3072,N_3049);
or U3125 (N_3125,N_3030,N_3017);
or U3126 (N_3126,N_3085,N_3001);
nor U3127 (N_3127,N_3075,N_3081);
or U3128 (N_3128,N_3059,N_3073);
or U3129 (N_3129,N_3047,N_3099);
nand U3130 (N_3130,N_3080,N_3021);
xor U3131 (N_3131,N_3018,N_3032);
nor U3132 (N_3132,N_3076,N_3038);
or U3133 (N_3133,N_3090,N_3092);
nor U3134 (N_3134,N_3065,N_3009);
and U3135 (N_3135,N_3016,N_3003);
nand U3136 (N_3136,N_3068,N_3011);
or U3137 (N_3137,N_3033,N_3048);
or U3138 (N_3138,N_3024,N_3088);
and U3139 (N_3139,N_3040,N_3060);
nand U3140 (N_3140,N_3043,N_3064);
nand U3141 (N_3141,N_3035,N_3079);
nand U3142 (N_3142,N_3070,N_3005);
or U3143 (N_3143,N_3025,N_3083);
and U3144 (N_3144,N_3095,N_3010);
or U3145 (N_3145,N_3093,N_3087);
nor U3146 (N_3146,N_3039,N_3013);
nor U3147 (N_3147,N_3062,N_3066);
xor U3148 (N_3148,N_3004,N_3063);
nor U3149 (N_3149,N_3056,N_3078);
nor U3150 (N_3150,N_3008,N_3050);
or U3151 (N_3151,N_3070,N_3067);
or U3152 (N_3152,N_3089,N_3096);
or U3153 (N_3153,N_3070,N_3016);
nand U3154 (N_3154,N_3006,N_3022);
nor U3155 (N_3155,N_3096,N_3023);
xor U3156 (N_3156,N_3092,N_3096);
nand U3157 (N_3157,N_3028,N_3019);
xnor U3158 (N_3158,N_3091,N_3026);
and U3159 (N_3159,N_3006,N_3094);
xor U3160 (N_3160,N_3056,N_3009);
nand U3161 (N_3161,N_3026,N_3040);
and U3162 (N_3162,N_3007,N_3030);
or U3163 (N_3163,N_3018,N_3089);
xor U3164 (N_3164,N_3007,N_3047);
nand U3165 (N_3165,N_3039,N_3070);
xnor U3166 (N_3166,N_3087,N_3040);
nand U3167 (N_3167,N_3026,N_3035);
nor U3168 (N_3168,N_3097,N_3070);
xor U3169 (N_3169,N_3040,N_3002);
nand U3170 (N_3170,N_3000,N_3097);
nor U3171 (N_3171,N_3033,N_3084);
nand U3172 (N_3172,N_3068,N_3036);
or U3173 (N_3173,N_3079,N_3046);
xnor U3174 (N_3174,N_3099,N_3008);
xnor U3175 (N_3175,N_3098,N_3021);
nand U3176 (N_3176,N_3005,N_3069);
nand U3177 (N_3177,N_3099,N_3076);
and U3178 (N_3178,N_3055,N_3023);
or U3179 (N_3179,N_3065,N_3023);
or U3180 (N_3180,N_3084,N_3011);
nand U3181 (N_3181,N_3009,N_3005);
or U3182 (N_3182,N_3091,N_3011);
and U3183 (N_3183,N_3042,N_3026);
nand U3184 (N_3184,N_3010,N_3024);
xor U3185 (N_3185,N_3083,N_3055);
nor U3186 (N_3186,N_3023,N_3078);
or U3187 (N_3187,N_3082,N_3099);
xnor U3188 (N_3188,N_3065,N_3081);
nand U3189 (N_3189,N_3005,N_3058);
xnor U3190 (N_3190,N_3094,N_3036);
nand U3191 (N_3191,N_3080,N_3024);
xnor U3192 (N_3192,N_3017,N_3090);
and U3193 (N_3193,N_3025,N_3026);
nor U3194 (N_3194,N_3037,N_3030);
nand U3195 (N_3195,N_3024,N_3070);
or U3196 (N_3196,N_3023,N_3057);
nand U3197 (N_3197,N_3093,N_3083);
and U3198 (N_3198,N_3089,N_3008);
nor U3199 (N_3199,N_3059,N_3035);
xnor U3200 (N_3200,N_3139,N_3119);
nand U3201 (N_3201,N_3177,N_3197);
and U3202 (N_3202,N_3154,N_3179);
or U3203 (N_3203,N_3151,N_3109);
nand U3204 (N_3204,N_3130,N_3162);
or U3205 (N_3205,N_3182,N_3153);
xor U3206 (N_3206,N_3126,N_3189);
xor U3207 (N_3207,N_3196,N_3137);
nor U3208 (N_3208,N_3180,N_3136);
and U3209 (N_3209,N_3188,N_3129);
nand U3210 (N_3210,N_3105,N_3199);
and U3211 (N_3211,N_3140,N_3143);
nor U3212 (N_3212,N_3163,N_3186);
nor U3213 (N_3213,N_3131,N_3144);
xnor U3214 (N_3214,N_3133,N_3114);
nand U3215 (N_3215,N_3155,N_3138);
and U3216 (N_3216,N_3148,N_3127);
or U3217 (N_3217,N_3106,N_3135);
or U3218 (N_3218,N_3159,N_3193);
nor U3219 (N_3219,N_3147,N_3132);
and U3220 (N_3220,N_3146,N_3108);
xnor U3221 (N_3221,N_3101,N_3125);
nor U3222 (N_3222,N_3187,N_3116);
xnor U3223 (N_3223,N_3158,N_3107);
nor U3224 (N_3224,N_3183,N_3103);
or U3225 (N_3225,N_3166,N_3110);
and U3226 (N_3226,N_3102,N_3117);
xnor U3227 (N_3227,N_3142,N_3141);
nand U3228 (N_3228,N_3168,N_3149);
nand U3229 (N_3229,N_3157,N_3128);
and U3230 (N_3230,N_3181,N_3118);
xnor U3231 (N_3231,N_3160,N_3190);
or U3232 (N_3232,N_3122,N_3191);
nand U3233 (N_3233,N_3134,N_3174);
nand U3234 (N_3234,N_3173,N_3115);
nand U3235 (N_3235,N_3112,N_3185);
nand U3236 (N_3236,N_3164,N_3124);
nor U3237 (N_3237,N_3100,N_3169);
or U3238 (N_3238,N_3113,N_3104);
and U3239 (N_3239,N_3192,N_3195);
xor U3240 (N_3240,N_3170,N_3123);
and U3241 (N_3241,N_3120,N_3150);
or U3242 (N_3242,N_3156,N_3172);
xnor U3243 (N_3243,N_3152,N_3176);
and U3244 (N_3244,N_3184,N_3161);
nor U3245 (N_3245,N_3145,N_3167);
xnor U3246 (N_3246,N_3121,N_3111);
or U3247 (N_3247,N_3178,N_3194);
or U3248 (N_3248,N_3165,N_3175);
xor U3249 (N_3249,N_3198,N_3171);
and U3250 (N_3250,N_3181,N_3195);
xor U3251 (N_3251,N_3181,N_3157);
and U3252 (N_3252,N_3137,N_3119);
or U3253 (N_3253,N_3128,N_3141);
or U3254 (N_3254,N_3108,N_3107);
xor U3255 (N_3255,N_3104,N_3129);
nor U3256 (N_3256,N_3172,N_3143);
xor U3257 (N_3257,N_3108,N_3118);
xor U3258 (N_3258,N_3161,N_3155);
and U3259 (N_3259,N_3116,N_3119);
nor U3260 (N_3260,N_3165,N_3135);
or U3261 (N_3261,N_3188,N_3124);
nor U3262 (N_3262,N_3172,N_3114);
xor U3263 (N_3263,N_3172,N_3159);
nand U3264 (N_3264,N_3115,N_3177);
nand U3265 (N_3265,N_3180,N_3141);
xor U3266 (N_3266,N_3183,N_3191);
nor U3267 (N_3267,N_3178,N_3100);
and U3268 (N_3268,N_3123,N_3142);
or U3269 (N_3269,N_3111,N_3153);
or U3270 (N_3270,N_3136,N_3124);
nor U3271 (N_3271,N_3167,N_3186);
xnor U3272 (N_3272,N_3160,N_3165);
or U3273 (N_3273,N_3114,N_3120);
nand U3274 (N_3274,N_3103,N_3138);
or U3275 (N_3275,N_3120,N_3195);
nor U3276 (N_3276,N_3154,N_3177);
or U3277 (N_3277,N_3187,N_3111);
and U3278 (N_3278,N_3152,N_3105);
xnor U3279 (N_3279,N_3113,N_3141);
nor U3280 (N_3280,N_3148,N_3109);
xor U3281 (N_3281,N_3196,N_3151);
xnor U3282 (N_3282,N_3160,N_3115);
or U3283 (N_3283,N_3115,N_3134);
nor U3284 (N_3284,N_3179,N_3158);
or U3285 (N_3285,N_3161,N_3153);
or U3286 (N_3286,N_3138,N_3184);
nand U3287 (N_3287,N_3161,N_3158);
and U3288 (N_3288,N_3104,N_3131);
and U3289 (N_3289,N_3173,N_3178);
nor U3290 (N_3290,N_3141,N_3139);
nor U3291 (N_3291,N_3144,N_3147);
xnor U3292 (N_3292,N_3103,N_3190);
xor U3293 (N_3293,N_3195,N_3169);
nor U3294 (N_3294,N_3150,N_3135);
nand U3295 (N_3295,N_3111,N_3192);
xnor U3296 (N_3296,N_3167,N_3102);
and U3297 (N_3297,N_3178,N_3131);
nor U3298 (N_3298,N_3107,N_3114);
and U3299 (N_3299,N_3158,N_3156);
or U3300 (N_3300,N_3284,N_3275);
nand U3301 (N_3301,N_3215,N_3212);
nand U3302 (N_3302,N_3290,N_3231);
or U3303 (N_3303,N_3260,N_3240);
or U3304 (N_3304,N_3201,N_3253);
xor U3305 (N_3305,N_3247,N_3205);
nor U3306 (N_3306,N_3210,N_3269);
nand U3307 (N_3307,N_3286,N_3298);
nor U3308 (N_3308,N_3296,N_3211);
and U3309 (N_3309,N_3288,N_3230);
nand U3310 (N_3310,N_3226,N_3244);
and U3311 (N_3311,N_3243,N_3202);
xor U3312 (N_3312,N_3209,N_3213);
nor U3313 (N_3313,N_3217,N_3266);
nor U3314 (N_3314,N_3251,N_3270);
or U3315 (N_3315,N_3225,N_3252);
nand U3316 (N_3316,N_3206,N_3220);
nor U3317 (N_3317,N_3249,N_3254);
and U3318 (N_3318,N_3291,N_3256);
and U3319 (N_3319,N_3241,N_3246);
nand U3320 (N_3320,N_3236,N_3214);
or U3321 (N_3321,N_3297,N_3263);
nor U3322 (N_3322,N_3200,N_3228);
nand U3323 (N_3323,N_3282,N_3279);
xnor U3324 (N_3324,N_3283,N_3278);
and U3325 (N_3325,N_3219,N_3287);
and U3326 (N_3326,N_3229,N_3271);
xor U3327 (N_3327,N_3273,N_3221);
xnor U3328 (N_3328,N_3259,N_3280);
xor U3329 (N_3329,N_3203,N_3295);
or U3330 (N_3330,N_3267,N_3264);
nor U3331 (N_3331,N_3222,N_3258);
and U3332 (N_3332,N_3242,N_3232);
xnor U3333 (N_3333,N_3218,N_3257);
nor U3334 (N_3334,N_3265,N_3238);
xnor U3335 (N_3335,N_3234,N_3281);
and U3336 (N_3336,N_3233,N_3227);
nand U3337 (N_3337,N_3276,N_3285);
xnor U3338 (N_3338,N_3299,N_3255);
nand U3339 (N_3339,N_3245,N_3289);
and U3340 (N_3340,N_3250,N_3292);
nand U3341 (N_3341,N_3237,N_3268);
nand U3342 (N_3342,N_3294,N_3262);
or U3343 (N_3343,N_3293,N_3235);
xnor U3344 (N_3344,N_3239,N_3277);
xnor U3345 (N_3345,N_3248,N_3224);
and U3346 (N_3346,N_3207,N_3223);
nor U3347 (N_3347,N_3204,N_3208);
and U3348 (N_3348,N_3272,N_3216);
or U3349 (N_3349,N_3261,N_3274);
or U3350 (N_3350,N_3291,N_3213);
or U3351 (N_3351,N_3297,N_3235);
and U3352 (N_3352,N_3276,N_3237);
nand U3353 (N_3353,N_3238,N_3297);
xnor U3354 (N_3354,N_3229,N_3213);
nor U3355 (N_3355,N_3297,N_3279);
nand U3356 (N_3356,N_3206,N_3237);
and U3357 (N_3357,N_3218,N_3252);
nand U3358 (N_3358,N_3218,N_3248);
or U3359 (N_3359,N_3240,N_3218);
nor U3360 (N_3360,N_3297,N_3275);
and U3361 (N_3361,N_3265,N_3259);
or U3362 (N_3362,N_3213,N_3226);
nand U3363 (N_3363,N_3296,N_3247);
nor U3364 (N_3364,N_3223,N_3200);
and U3365 (N_3365,N_3212,N_3232);
nand U3366 (N_3366,N_3231,N_3238);
xnor U3367 (N_3367,N_3201,N_3246);
nor U3368 (N_3368,N_3255,N_3206);
xnor U3369 (N_3369,N_3234,N_3253);
and U3370 (N_3370,N_3246,N_3252);
nand U3371 (N_3371,N_3205,N_3216);
or U3372 (N_3372,N_3273,N_3262);
or U3373 (N_3373,N_3270,N_3275);
or U3374 (N_3374,N_3294,N_3295);
nor U3375 (N_3375,N_3289,N_3217);
xnor U3376 (N_3376,N_3246,N_3205);
and U3377 (N_3377,N_3211,N_3267);
xor U3378 (N_3378,N_3238,N_3216);
nor U3379 (N_3379,N_3297,N_3269);
xnor U3380 (N_3380,N_3276,N_3234);
xor U3381 (N_3381,N_3251,N_3235);
nor U3382 (N_3382,N_3265,N_3244);
nand U3383 (N_3383,N_3277,N_3215);
nand U3384 (N_3384,N_3223,N_3271);
xor U3385 (N_3385,N_3218,N_3256);
nand U3386 (N_3386,N_3223,N_3293);
and U3387 (N_3387,N_3291,N_3270);
nor U3388 (N_3388,N_3250,N_3259);
nand U3389 (N_3389,N_3285,N_3280);
nand U3390 (N_3390,N_3206,N_3269);
or U3391 (N_3391,N_3283,N_3277);
or U3392 (N_3392,N_3258,N_3240);
xor U3393 (N_3393,N_3236,N_3258);
nor U3394 (N_3394,N_3227,N_3285);
and U3395 (N_3395,N_3283,N_3220);
nor U3396 (N_3396,N_3242,N_3281);
nor U3397 (N_3397,N_3205,N_3208);
xnor U3398 (N_3398,N_3277,N_3286);
and U3399 (N_3399,N_3280,N_3232);
xnor U3400 (N_3400,N_3340,N_3381);
nand U3401 (N_3401,N_3310,N_3376);
nor U3402 (N_3402,N_3334,N_3354);
nand U3403 (N_3403,N_3391,N_3336);
nand U3404 (N_3404,N_3327,N_3352);
nor U3405 (N_3405,N_3312,N_3314);
nor U3406 (N_3406,N_3321,N_3362);
nand U3407 (N_3407,N_3366,N_3389);
xnor U3408 (N_3408,N_3387,N_3360);
xnor U3409 (N_3409,N_3329,N_3322);
xnor U3410 (N_3410,N_3398,N_3399);
xnor U3411 (N_3411,N_3350,N_3332);
or U3412 (N_3412,N_3374,N_3323);
xnor U3413 (N_3413,N_3317,N_3370);
nand U3414 (N_3414,N_3377,N_3363);
nor U3415 (N_3415,N_3313,N_3379);
xor U3416 (N_3416,N_3395,N_3320);
and U3417 (N_3417,N_3302,N_3339);
xnor U3418 (N_3418,N_3305,N_3393);
and U3419 (N_3419,N_3356,N_3392);
or U3420 (N_3420,N_3369,N_3300);
or U3421 (N_3421,N_3342,N_3396);
and U3422 (N_3422,N_3361,N_3337);
nand U3423 (N_3423,N_3375,N_3344);
and U3424 (N_3424,N_3315,N_3357);
nand U3425 (N_3425,N_3368,N_3303);
or U3426 (N_3426,N_3378,N_3383);
nand U3427 (N_3427,N_3319,N_3346);
or U3428 (N_3428,N_3372,N_3338);
nor U3429 (N_3429,N_3390,N_3307);
or U3430 (N_3430,N_3385,N_3325);
nand U3431 (N_3431,N_3380,N_3351);
nor U3432 (N_3432,N_3324,N_3382);
nand U3433 (N_3433,N_3306,N_3347);
and U3434 (N_3434,N_3364,N_3397);
xnor U3435 (N_3435,N_3328,N_3348);
and U3436 (N_3436,N_3343,N_3333);
or U3437 (N_3437,N_3330,N_3359);
or U3438 (N_3438,N_3345,N_3349);
xor U3439 (N_3439,N_3394,N_3365);
or U3440 (N_3440,N_3373,N_3371);
nor U3441 (N_3441,N_3367,N_3358);
or U3442 (N_3442,N_3388,N_3304);
or U3443 (N_3443,N_3318,N_3384);
and U3444 (N_3444,N_3309,N_3308);
and U3445 (N_3445,N_3331,N_3311);
or U3446 (N_3446,N_3326,N_3335);
nor U3447 (N_3447,N_3353,N_3386);
nand U3448 (N_3448,N_3341,N_3301);
nor U3449 (N_3449,N_3355,N_3316);
and U3450 (N_3450,N_3301,N_3322);
xor U3451 (N_3451,N_3388,N_3308);
xor U3452 (N_3452,N_3397,N_3389);
and U3453 (N_3453,N_3383,N_3335);
and U3454 (N_3454,N_3383,N_3389);
and U3455 (N_3455,N_3396,N_3353);
xor U3456 (N_3456,N_3311,N_3390);
xnor U3457 (N_3457,N_3393,N_3328);
xor U3458 (N_3458,N_3386,N_3385);
nor U3459 (N_3459,N_3325,N_3366);
nor U3460 (N_3460,N_3352,N_3302);
nand U3461 (N_3461,N_3352,N_3334);
nand U3462 (N_3462,N_3374,N_3304);
or U3463 (N_3463,N_3310,N_3351);
and U3464 (N_3464,N_3319,N_3355);
xor U3465 (N_3465,N_3392,N_3374);
nand U3466 (N_3466,N_3346,N_3358);
xor U3467 (N_3467,N_3381,N_3376);
nor U3468 (N_3468,N_3363,N_3379);
or U3469 (N_3469,N_3349,N_3319);
or U3470 (N_3470,N_3372,N_3374);
nand U3471 (N_3471,N_3334,N_3346);
nor U3472 (N_3472,N_3366,N_3324);
and U3473 (N_3473,N_3340,N_3398);
and U3474 (N_3474,N_3356,N_3329);
nand U3475 (N_3475,N_3335,N_3348);
or U3476 (N_3476,N_3341,N_3383);
or U3477 (N_3477,N_3316,N_3324);
nand U3478 (N_3478,N_3342,N_3312);
or U3479 (N_3479,N_3327,N_3396);
nor U3480 (N_3480,N_3319,N_3373);
nor U3481 (N_3481,N_3396,N_3343);
and U3482 (N_3482,N_3327,N_3360);
nand U3483 (N_3483,N_3381,N_3358);
and U3484 (N_3484,N_3372,N_3336);
and U3485 (N_3485,N_3382,N_3388);
nor U3486 (N_3486,N_3306,N_3378);
or U3487 (N_3487,N_3313,N_3312);
nand U3488 (N_3488,N_3374,N_3396);
and U3489 (N_3489,N_3300,N_3325);
nor U3490 (N_3490,N_3314,N_3372);
nor U3491 (N_3491,N_3329,N_3330);
and U3492 (N_3492,N_3351,N_3329);
or U3493 (N_3493,N_3385,N_3347);
xor U3494 (N_3494,N_3361,N_3307);
and U3495 (N_3495,N_3312,N_3306);
or U3496 (N_3496,N_3323,N_3358);
xnor U3497 (N_3497,N_3382,N_3327);
nor U3498 (N_3498,N_3350,N_3368);
or U3499 (N_3499,N_3375,N_3359);
xnor U3500 (N_3500,N_3482,N_3431);
or U3501 (N_3501,N_3432,N_3491);
nand U3502 (N_3502,N_3485,N_3423);
or U3503 (N_3503,N_3414,N_3455);
nor U3504 (N_3504,N_3407,N_3463);
nor U3505 (N_3505,N_3418,N_3498);
and U3506 (N_3506,N_3492,N_3420);
and U3507 (N_3507,N_3474,N_3450);
nor U3508 (N_3508,N_3472,N_3490);
nor U3509 (N_3509,N_3409,N_3480);
xor U3510 (N_3510,N_3475,N_3478);
nand U3511 (N_3511,N_3456,N_3433);
nor U3512 (N_3512,N_3443,N_3413);
or U3513 (N_3513,N_3403,N_3457);
or U3514 (N_3514,N_3435,N_3438);
or U3515 (N_3515,N_3496,N_3417);
xor U3516 (N_3516,N_3430,N_3429);
and U3517 (N_3517,N_3400,N_3404);
and U3518 (N_3518,N_3424,N_3405);
and U3519 (N_3519,N_3461,N_3427);
nand U3520 (N_3520,N_3499,N_3448);
xnor U3521 (N_3521,N_3415,N_3444);
or U3522 (N_3522,N_3488,N_3477);
nor U3523 (N_3523,N_3416,N_3419);
xor U3524 (N_3524,N_3483,N_3410);
xnor U3525 (N_3525,N_3487,N_3402);
xor U3526 (N_3526,N_3425,N_3436);
and U3527 (N_3527,N_3412,N_3493);
and U3528 (N_3528,N_3401,N_3447);
or U3529 (N_3529,N_3462,N_3446);
and U3530 (N_3530,N_3466,N_3445);
nor U3531 (N_3531,N_3426,N_3434);
xnor U3532 (N_3532,N_3408,N_3460);
xor U3533 (N_3533,N_3476,N_3428);
or U3534 (N_3534,N_3468,N_3484);
nand U3535 (N_3535,N_3471,N_3440);
and U3536 (N_3536,N_3479,N_3467);
or U3537 (N_3537,N_3459,N_3441);
nand U3538 (N_3538,N_3451,N_3470);
nor U3539 (N_3539,N_3464,N_3411);
nor U3540 (N_3540,N_3406,N_3452);
and U3541 (N_3541,N_3422,N_3469);
or U3542 (N_3542,N_3495,N_3442);
xor U3543 (N_3543,N_3437,N_3473);
nand U3544 (N_3544,N_3465,N_3486);
xor U3545 (N_3545,N_3489,N_3494);
and U3546 (N_3546,N_3497,N_3449);
or U3547 (N_3547,N_3458,N_3421);
or U3548 (N_3548,N_3439,N_3454);
nand U3549 (N_3549,N_3453,N_3481);
and U3550 (N_3550,N_3447,N_3445);
xnor U3551 (N_3551,N_3466,N_3448);
and U3552 (N_3552,N_3485,N_3414);
nor U3553 (N_3553,N_3478,N_3400);
xnor U3554 (N_3554,N_3423,N_3441);
nor U3555 (N_3555,N_3463,N_3489);
nand U3556 (N_3556,N_3489,N_3485);
or U3557 (N_3557,N_3413,N_3416);
xor U3558 (N_3558,N_3419,N_3453);
nor U3559 (N_3559,N_3416,N_3408);
xnor U3560 (N_3560,N_3418,N_3497);
nand U3561 (N_3561,N_3459,N_3476);
and U3562 (N_3562,N_3432,N_3462);
and U3563 (N_3563,N_3442,N_3458);
nor U3564 (N_3564,N_3407,N_3423);
xor U3565 (N_3565,N_3440,N_3422);
nand U3566 (N_3566,N_3402,N_3415);
nand U3567 (N_3567,N_3418,N_3493);
xor U3568 (N_3568,N_3445,N_3460);
and U3569 (N_3569,N_3450,N_3409);
and U3570 (N_3570,N_3452,N_3473);
nand U3571 (N_3571,N_3424,N_3461);
xor U3572 (N_3572,N_3487,N_3417);
or U3573 (N_3573,N_3490,N_3454);
xnor U3574 (N_3574,N_3484,N_3462);
xnor U3575 (N_3575,N_3415,N_3496);
or U3576 (N_3576,N_3407,N_3479);
or U3577 (N_3577,N_3449,N_3474);
nand U3578 (N_3578,N_3429,N_3454);
or U3579 (N_3579,N_3452,N_3421);
xor U3580 (N_3580,N_3499,N_3486);
xnor U3581 (N_3581,N_3446,N_3473);
or U3582 (N_3582,N_3412,N_3425);
nor U3583 (N_3583,N_3487,N_3449);
xor U3584 (N_3584,N_3449,N_3414);
and U3585 (N_3585,N_3409,N_3489);
nand U3586 (N_3586,N_3448,N_3479);
xnor U3587 (N_3587,N_3494,N_3407);
or U3588 (N_3588,N_3444,N_3400);
xor U3589 (N_3589,N_3484,N_3457);
and U3590 (N_3590,N_3418,N_3425);
nand U3591 (N_3591,N_3405,N_3457);
nor U3592 (N_3592,N_3409,N_3435);
xor U3593 (N_3593,N_3463,N_3413);
or U3594 (N_3594,N_3478,N_3465);
nand U3595 (N_3595,N_3492,N_3453);
nand U3596 (N_3596,N_3489,N_3478);
nand U3597 (N_3597,N_3441,N_3406);
xnor U3598 (N_3598,N_3473,N_3444);
nor U3599 (N_3599,N_3459,N_3491);
or U3600 (N_3600,N_3558,N_3502);
nand U3601 (N_3601,N_3547,N_3580);
xnor U3602 (N_3602,N_3576,N_3574);
nor U3603 (N_3603,N_3567,N_3533);
and U3604 (N_3604,N_3554,N_3553);
nor U3605 (N_3605,N_3516,N_3599);
and U3606 (N_3606,N_3579,N_3506);
and U3607 (N_3607,N_3556,N_3501);
nor U3608 (N_3608,N_3577,N_3584);
nor U3609 (N_3609,N_3587,N_3524);
xor U3610 (N_3610,N_3589,N_3583);
or U3611 (N_3611,N_3526,N_3591);
nor U3612 (N_3612,N_3529,N_3595);
nand U3613 (N_3613,N_3540,N_3545);
nor U3614 (N_3614,N_3590,N_3517);
nand U3615 (N_3615,N_3534,N_3566);
xnor U3616 (N_3616,N_3531,N_3571);
nand U3617 (N_3617,N_3518,N_3512);
or U3618 (N_3618,N_3542,N_3565);
or U3619 (N_3619,N_3544,N_3570);
nand U3620 (N_3620,N_3575,N_3532);
nand U3621 (N_3621,N_3562,N_3559);
and U3622 (N_3622,N_3581,N_3519);
and U3623 (N_3623,N_3539,N_3586);
nand U3624 (N_3624,N_3557,N_3594);
nand U3625 (N_3625,N_3546,N_3543);
nor U3626 (N_3626,N_3598,N_3568);
and U3627 (N_3627,N_3552,N_3573);
xor U3628 (N_3628,N_3505,N_3508);
nor U3629 (N_3629,N_3514,N_3593);
nand U3630 (N_3630,N_3507,N_3548);
and U3631 (N_3631,N_3541,N_3527);
nor U3632 (N_3632,N_3538,N_3509);
nand U3633 (N_3633,N_3504,N_3561);
xor U3634 (N_3634,N_3569,N_3525);
nand U3635 (N_3635,N_3592,N_3537);
nand U3636 (N_3636,N_3596,N_3530);
and U3637 (N_3637,N_3503,N_3535);
xor U3638 (N_3638,N_3536,N_3578);
and U3639 (N_3639,N_3582,N_3551);
xor U3640 (N_3640,N_3550,N_3521);
or U3641 (N_3641,N_3528,N_3572);
nor U3642 (N_3642,N_3560,N_3510);
or U3643 (N_3643,N_3555,N_3549);
xnor U3644 (N_3644,N_3515,N_3585);
nor U3645 (N_3645,N_3588,N_3511);
xnor U3646 (N_3646,N_3522,N_3597);
and U3647 (N_3647,N_3520,N_3500);
or U3648 (N_3648,N_3513,N_3563);
or U3649 (N_3649,N_3564,N_3523);
xor U3650 (N_3650,N_3500,N_3574);
nand U3651 (N_3651,N_3598,N_3510);
or U3652 (N_3652,N_3560,N_3570);
and U3653 (N_3653,N_3573,N_3594);
or U3654 (N_3654,N_3576,N_3578);
nand U3655 (N_3655,N_3589,N_3506);
and U3656 (N_3656,N_3576,N_3580);
and U3657 (N_3657,N_3556,N_3566);
and U3658 (N_3658,N_3504,N_3510);
nor U3659 (N_3659,N_3513,N_3562);
nand U3660 (N_3660,N_3583,N_3524);
and U3661 (N_3661,N_3561,N_3553);
and U3662 (N_3662,N_3591,N_3515);
nand U3663 (N_3663,N_3590,N_3581);
or U3664 (N_3664,N_3510,N_3518);
xnor U3665 (N_3665,N_3571,N_3563);
nor U3666 (N_3666,N_3552,N_3563);
nor U3667 (N_3667,N_3569,N_3519);
nand U3668 (N_3668,N_3597,N_3555);
xor U3669 (N_3669,N_3584,N_3549);
xor U3670 (N_3670,N_3566,N_3517);
nand U3671 (N_3671,N_3591,N_3582);
nand U3672 (N_3672,N_3585,N_3545);
nand U3673 (N_3673,N_3549,N_3547);
nand U3674 (N_3674,N_3514,N_3575);
nand U3675 (N_3675,N_3554,N_3527);
and U3676 (N_3676,N_3533,N_3517);
xor U3677 (N_3677,N_3526,N_3525);
xor U3678 (N_3678,N_3534,N_3545);
nor U3679 (N_3679,N_3573,N_3506);
nor U3680 (N_3680,N_3502,N_3541);
and U3681 (N_3681,N_3554,N_3591);
and U3682 (N_3682,N_3509,N_3512);
or U3683 (N_3683,N_3551,N_3548);
and U3684 (N_3684,N_3555,N_3530);
xor U3685 (N_3685,N_3521,N_3517);
nand U3686 (N_3686,N_3564,N_3577);
or U3687 (N_3687,N_3559,N_3514);
or U3688 (N_3688,N_3543,N_3571);
and U3689 (N_3689,N_3550,N_3532);
or U3690 (N_3690,N_3512,N_3597);
or U3691 (N_3691,N_3504,N_3520);
nor U3692 (N_3692,N_3510,N_3573);
nand U3693 (N_3693,N_3569,N_3560);
nor U3694 (N_3694,N_3514,N_3513);
nor U3695 (N_3695,N_3594,N_3552);
nand U3696 (N_3696,N_3574,N_3594);
or U3697 (N_3697,N_3500,N_3546);
and U3698 (N_3698,N_3584,N_3551);
or U3699 (N_3699,N_3539,N_3525);
nor U3700 (N_3700,N_3685,N_3667);
and U3701 (N_3701,N_3680,N_3679);
nor U3702 (N_3702,N_3683,N_3663);
nand U3703 (N_3703,N_3643,N_3678);
and U3704 (N_3704,N_3657,N_3675);
or U3705 (N_3705,N_3658,N_3609);
nor U3706 (N_3706,N_3681,N_3631);
nand U3707 (N_3707,N_3648,N_3651);
xnor U3708 (N_3708,N_3655,N_3692);
xor U3709 (N_3709,N_3637,N_3600);
and U3710 (N_3710,N_3694,N_3647);
xnor U3711 (N_3711,N_3671,N_3634);
xor U3712 (N_3712,N_3687,N_3641);
xnor U3713 (N_3713,N_3659,N_3632);
and U3714 (N_3714,N_3620,N_3615);
or U3715 (N_3715,N_3604,N_3640);
and U3716 (N_3716,N_3630,N_3627);
or U3717 (N_3717,N_3665,N_3639);
and U3718 (N_3718,N_3670,N_3603);
or U3719 (N_3719,N_3698,N_3616);
xnor U3720 (N_3720,N_3626,N_3624);
xor U3721 (N_3721,N_3669,N_3662);
or U3722 (N_3722,N_3619,N_3650);
and U3723 (N_3723,N_3686,N_3673);
or U3724 (N_3724,N_3608,N_3625);
nor U3725 (N_3725,N_3606,N_3695);
xnor U3726 (N_3726,N_3633,N_3682);
or U3727 (N_3727,N_3676,N_3644);
nor U3728 (N_3728,N_3652,N_3623);
xor U3729 (N_3729,N_3668,N_3642);
and U3730 (N_3730,N_3607,N_3621);
xnor U3731 (N_3731,N_3635,N_3661);
xor U3732 (N_3732,N_3617,N_3656);
or U3733 (N_3733,N_3645,N_3649);
or U3734 (N_3734,N_3696,N_3614);
and U3735 (N_3735,N_3622,N_3638);
and U3736 (N_3736,N_3697,N_3628);
and U3737 (N_3737,N_3602,N_3612);
nor U3738 (N_3738,N_3684,N_3605);
nor U3739 (N_3739,N_3699,N_3666);
nor U3740 (N_3740,N_3646,N_3688);
nand U3741 (N_3741,N_3654,N_3689);
nor U3742 (N_3742,N_3636,N_3693);
xor U3743 (N_3743,N_3601,N_3610);
or U3744 (N_3744,N_3613,N_3618);
or U3745 (N_3745,N_3690,N_3629);
xnor U3746 (N_3746,N_3660,N_3674);
xor U3747 (N_3747,N_3653,N_3611);
xor U3748 (N_3748,N_3691,N_3664);
or U3749 (N_3749,N_3677,N_3672);
nand U3750 (N_3750,N_3666,N_3689);
nor U3751 (N_3751,N_3615,N_3600);
and U3752 (N_3752,N_3655,N_3678);
and U3753 (N_3753,N_3699,N_3641);
nor U3754 (N_3754,N_3623,N_3627);
nor U3755 (N_3755,N_3608,N_3622);
or U3756 (N_3756,N_3681,N_3666);
nor U3757 (N_3757,N_3621,N_3649);
xnor U3758 (N_3758,N_3619,N_3633);
xor U3759 (N_3759,N_3630,N_3662);
nor U3760 (N_3760,N_3670,N_3698);
or U3761 (N_3761,N_3681,N_3694);
xor U3762 (N_3762,N_3658,N_3630);
nand U3763 (N_3763,N_3648,N_3695);
nand U3764 (N_3764,N_3601,N_3614);
nand U3765 (N_3765,N_3679,N_3699);
xor U3766 (N_3766,N_3672,N_3663);
nor U3767 (N_3767,N_3606,N_3615);
nand U3768 (N_3768,N_3684,N_3630);
nor U3769 (N_3769,N_3641,N_3633);
nand U3770 (N_3770,N_3680,N_3668);
nand U3771 (N_3771,N_3628,N_3669);
and U3772 (N_3772,N_3634,N_3662);
xnor U3773 (N_3773,N_3673,N_3692);
and U3774 (N_3774,N_3632,N_3609);
and U3775 (N_3775,N_3648,N_3681);
or U3776 (N_3776,N_3682,N_3617);
or U3777 (N_3777,N_3693,N_3617);
or U3778 (N_3778,N_3629,N_3603);
nor U3779 (N_3779,N_3688,N_3650);
nand U3780 (N_3780,N_3696,N_3636);
and U3781 (N_3781,N_3603,N_3696);
nand U3782 (N_3782,N_3647,N_3627);
and U3783 (N_3783,N_3648,N_3649);
nor U3784 (N_3784,N_3656,N_3699);
and U3785 (N_3785,N_3607,N_3613);
nor U3786 (N_3786,N_3614,N_3639);
xnor U3787 (N_3787,N_3667,N_3653);
nor U3788 (N_3788,N_3653,N_3698);
or U3789 (N_3789,N_3646,N_3698);
xor U3790 (N_3790,N_3639,N_3652);
or U3791 (N_3791,N_3675,N_3604);
xnor U3792 (N_3792,N_3689,N_3645);
xor U3793 (N_3793,N_3651,N_3602);
or U3794 (N_3794,N_3621,N_3609);
nor U3795 (N_3795,N_3639,N_3606);
nand U3796 (N_3796,N_3607,N_3622);
xor U3797 (N_3797,N_3659,N_3682);
xnor U3798 (N_3798,N_3632,N_3612);
nor U3799 (N_3799,N_3663,N_3626);
nor U3800 (N_3800,N_3712,N_3794);
or U3801 (N_3801,N_3782,N_3755);
nand U3802 (N_3802,N_3790,N_3771);
nor U3803 (N_3803,N_3795,N_3792);
or U3804 (N_3804,N_3723,N_3745);
nor U3805 (N_3805,N_3714,N_3726);
xnor U3806 (N_3806,N_3798,N_3752);
nand U3807 (N_3807,N_3727,N_3718);
nor U3808 (N_3808,N_3767,N_3735);
nor U3809 (N_3809,N_3719,N_3703);
nor U3810 (N_3810,N_3780,N_3743);
or U3811 (N_3811,N_3777,N_3707);
or U3812 (N_3812,N_3737,N_3775);
nand U3813 (N_3813,N_3700,N_3759);
or U3814 (N_3814,N_3710,N_3785);
or U3815 (N_3815,N_3734,N_3770);
nand U3816 (N_3816,N_3709,N_3746);
and U3817 (N_3817,N_3791,N_3722);
or U3818 (N_3818,N_3788,N_3702);
nand U3819 (N_3819,N_3760,N_3784);
xor U3820 (N_3820,N_3774,N_3793);
nor U3821 (N_3821,N_3779,N_3761);
and U3822 (N_3822,N_3732,N_3766);
nor U3823 (N_3823,N_3704,N_3748);
nor U3824 (N_3824,N_3753,N_3750);
nor U3825 (N_3825,N_3736,N_3730);
and U3826 (N_3826,N_3776,N_3721);
or U3827 (N_3827,N_3705,N_3716);
xnor U3828 (N_3828,N_3733,N_3728);
or U3829 (N_3829,N_3720,N_3768);
xnor U3830 (N_3830,N_3783,N_3701);
nor U3831 (N_3831,N_3756,N_3717);
and U3832 (N_3832,N_3731,N_3725);
or U3833 (N_3833,N_3762,N_3772);
xor U3834 (N_3834,N_3754,N_3739);
nand U3835 (N_3835,N_3740,N_3769);
and U3836 (N_3836,N_3741,N_3744);
and U3837 (N_3837,N_3787,N_3724);
xor U3838 (N_3838,N_3764,N_3742);
and U3839 (N_3839,N_3773,N_3749);
nand U3840 (N_3840,N_3789,N_3781);
and U3841 (N_3841,N_3711,N_3799);
nor U3842 (N_3842,N_3765,N_3778);
nand U3843 (N_3843,N_3738,N_3729);
nand U3844 (N_3844,N_3706,N_3751);
nor U3845 (N_3845,N_3758,N_3708);
xnor U3846 (N_3846,N_3757,N_3796);
and U3847 (N_3847,N_3763,N_3797);
or U3848 (N_3848,N_3747,N_3786);
nand U3849 (N_3849,N_3715,N_3713);
and U3850 (N_3850,N_3750,N_3742);
or U3851 (N_3851,N_3743,N_3740);
nor U3852 (N_3852,N_3704,N_3738);
nor U3853 (N_3853,N_3702,N_3750);
nor U3854 (N_3854,N_3751,N_3717);
or U3855 (N_3855,N_3793,N_3781);
nor U3856 (N_3856,N_3796,N_3761);
or U3857 (N_3857,N_3789,N_3718);
or U3858 (N_3858,N_3742,N_3747);
or U3859 (N_3859,N_3760,N_3724);
nor U3860 (N_3860,N_3712,N_3759);
or U3861 (N_3861,N_3710,N_3701);
xnor U3862 (N_3862,N_3737,N_3798);
or U3863 (N_3863,N_3717,N_3765);
xor U3864 (N_3864,N_3756,N_3725);
xor U3865 (N_3865,N_3735,N_3790);
xor U3866 (N_3866,N_3726,N_3790);
or U3867 (N_3867,N_3764,N_3780);
nand U3868 (N_3868,N_3762,N_3700);
nand U3869 (N_3869,N_3709,N_3779);
xnor U3870 (N_3870,N_3733,N_3725);
nand U3871 (N_3871,N_3752,N_3712);
and U3872 (N_3872,N_3728,N_3795);
nand U3873 (N_3873,N_3724,N_3740);
and U3874 (N_3874,N_3735,N_3775);
and U3875 (N_3875,N_3778,N_3702);
and U3876 (N_3876,N_3734,N_3761);
nand U3877 (N_3877,N_3727,N_3732);
xor U3878 (N_3878,N_3771,N_3714);
nor U3879 (N_3879,N_3741,N_3704);
nand U3880 (N_3880,N_3776,N_3743);
or U3881 (N_3881,N_3776,N_3796);
and U3882 (N_3882,N_3724,N_3766);
xnor U3883 (N_3883,N_3728,N_3704);
nand U3884 (N_3884,N_3766,N_3730);
or U3885 (N_3885,N_3712,N_3708);
xnor U3886 (N_3886,N_3725,N_3742);
xnor U3887 (N_3887,N_3706,N_3765);
or U3888 (N_3888,N_3764,N_3708);
nor U3889 (N_3889,N_3758,N_3715);
and U3890 (N_3890,N_3728,N_3762);
or U3891 (N_3891,N_3727,N_3799);
nor U3892 (N_3892,N_3769,N_3758);
nor U3893 (N_3893,N_3796,N_3743);
xor U3894 (N_3894,N_3792,N_3784);
nor U3895 (N_3895,N_3795,N_3758);
or U3896 (N_3896,N_3772,N_3707);
xnor U3897 (N_3897,N_3729,N_3753);
xnor U3898 (N_3898,N_3721,N_3732);
nor U3899 (N_3899,N_3709,N_3752);
and U3900 (N_3900,N_3831,N_3893);
and U3901 (N_3901,N_3822,N_3850);
and U3902 (N_3902,N_3827,N_3862);
or U3903 (N_3903,N_3878,N_3876);
nor U3904 (N_3904,N_3818,N_3875);
nor U3905 (N_3905,N_3865,N_3814);
xor U3906 (N_3906,N_3881,N_3846);
nor U3907 (N_3907,N_3834,N_3842);
and U3908 (N_3908,N_3877,N_3803);
and U3909 (N_3909,N_3837,N_3815);
nor U3910 (N_3910,N_3861,N_3869);
nor U3911 (N_3911,N_3858,N_3894);
nor U3912 (N_3912,N_3883,N_3891);
nor U3913 (N_3913,N_3809,N_3885);
nor U3914 (N_3914,N_3899,N_3804);
and U3915 (N_3915,N_3808,N_3802);
xor U3916 (N_3916,N_3816,N_3855);
nor U3917 (N_3917,N_3845,N_3800);
nor U3918 (N_3918,N_3867,N_3879);
or U3919 (N_3919,N_3897,N_3833);
or U3920 (N_3920,N_3811,N_3856);
nor U3921 (N_3921,N_3825,N_3860);
xor U3922 (N_3922,N_3848,N_3812);
nor U3923 (N_3923,N_3854,N_3880);
and U3924 (N_3924,N_3896,N_3820);
nand U3925 (N_3925,N_3828,N_3843);
and U3926 (N_3926,N_3806,N_3886);
or U3927 (N_3927,N_3840,N_3898);
nor U3928 (N_3928,N_3817,N_3838);
and U3929 (N_3929,N_3813,N_3863);
and U3930 (N_3930,N_3868,N_3871);
xnor U3931 (N_3931,N_3853,N_3810);
nor U3932 (N_3932,N_3873,N_3821);
nand U3933 (N_3933,N_3801,N_3857);
or U3934 (N_3934,N_3849,N_3852);
or U3935 (N_3935,N_3870,N_3805);
and U3936 (N_3936,N_3819,N_3884);
and U3937 (N_3937,N_3889,N_3826);
nand U3938 (N_3938,N_3830,N_3807);
nand U3939 (N_3939,N_3882,N_3864);
nand U3940 (N_3940,N_3835,N_3874);
or U3941 (N_3941,N_3847,N_3841);
or U3942 (N_3942,N_3887,N_3832);
nor U3943 (N_3943,N_3888,N_3824);
or U3944 (N_3944,N_3851,N_3872);
or U3945 (N_3945,N_3823,N_3844);
nor U3946 (N_3946,N_3890,N_3892);
xnor U3947 (N_3947,N_3836,N_3829);
and U3948 (N_3948,N_3859,N_3839);
nand U3949 (N_3949,N_3895,N_3866);
nor U3950 (N_3950,N_3838,N_3845);
nand U3951 (N_3951,N_3814,N_3842);
or U3952 (N_3952,N_3848,N_3899);
and U3953 (N_3953,N_3841,N_3857);
nor U3954 (N_3954,N_3812,N_3824);
or U3955 (N_3955,N_3805,N_3816);
or U3956 (N_3956,N_3866,N_3814);
nand U3957 (N_3957,N_3887,N_3883);
xor U3958 (N_3958,N_3846,N_3852);
xor U3959 (N_3959,N_3887,N_3839);
nand U3960 (N_3960,N_3886,N_3810);
xor U3961 (N_3961,N_3836,N_3870);
nand U3962 (N_3962,N_3866,N_3807);
nor U3963 (N_3963,N_3822,N_3824);
nor U3964 (N_3964,N_3840,N_3865);
and U3965 (N_3965,N_3803,N_3869);
and U3966 (N_3966,N_3830,N_3855);
xnor U3967 (N_3967,N_3814,N_3859);
or U3968 (N_3968,N_3828,N_3801);
nand U3969 (N_3969,N_3810,N_3892);
nand U3970 (N_3970,N_3877,N_3827);
nand U3971 (N_3971,N_3859,N_3806);
xor U3972 (N_3972,N_3823,N_3882);
nor U3973 (N_3973,N_3883,N_3862);
nor U3974 (N_3974,N_3818,N_3809);
or U3975 (N_3975,N_3825,N_3876);
nor U3976 (N_3976,N_3807,N_3822);
nor U3977 (N_3977,N_3801,N_3891);
and U3978 (N_3978,N_3811,N_3837);
nor U3979 (N_3979,N_3849,N_3860);
nor U3980 (N_3980,N_3837,N_3877);
or U3981 (N_3981,N_3830,N_3818);
xnor U3982 (N_3982,N_3805,N_3836);
xnor U3983 (N_3983,N_3887,N_3860);
xnor U3984 (N_3984,N_3863,N_3810);
nor U3985 (N_3985,N_3840,N_3824);
nor U3986 (N_3986,N_3893,N_3865);
xnor U3987 (N_3987,N_3861,N_3835);
nor U3988 (N_3988,N_3877,N_3821);
nand U3989 (N_3989,N_3844,N_3873);
nand U3990 (N_3990,N_3852,N_3803);
and U3991 (N_3991,N_3875,N_3831);
nor U3992 (N_3992,N_3896,N_3874);
xor U3993 (N_3993,N_3826,N_3886);
xnor U3994 (N_3994,N_3800,N_3846);
xnor U3995 (N_3995,N_3854,N_3822);
nand U3996 (N_3996,N_3818,N_3869);
xnor U3997 (N_3997,N_3868,N_3818);
nand U3998 (N_3998,N_3851,N_3810);
and U3999 (N_3999,N_3820,N_3882);
or U4000 (N_4000,N_3986,N_3966);
nand U4001 (N_4001,N_3983,N_3921);
xor U4002 (N_4002,N_3995,N_3938);
nand U4003 (N_4003,N_3965,N_3999);
nand U4004 (N_4004,N_3927,N_3945);
or U4005 (N_4005,N_3982,N_3990);
nor U4006 (N_4006,N_3923,N_3913);
or U4007 (N_4007,N_3933,N_3956);
or U4008 (N_4008,N_3941,N_3903);
or U4009 (N_4009,N_3924,N_3926);
nand U4010 (N_4010,N_3988,N_3939);
nor U4011 (N_4011,N_3958,N_3900);
nand U4012 (N_4012,N_3974,N_3992);
and U4013 (N_4013,N_3915,N_3910);
or U4014 (N_4014,N_3975,N_3959);
nand U4015 (N_4015,N_3979,N_3929);
and U4016 (N_4016,N_3940,N_3914);
and U4017 (N_4017,N_3947,N_3930);
nand U4018 (N_4018,N_3996,N_3993);
and U4019 (N_4019,N_3948,N_3949);
nor U4020 (N_4020,N_3978,N_3953);
or U4021 (N_4021,N_3918,N_3901);
or U4022 (N_4022,N_3904,N_3932);
nor U4023 (N_4023,N_3931,N_3991);
and U4024 (N_4024,N_3920,N_3909);
xor U4025 (N_4025,N_3994,N_3984);
and U4026 (N_4026,N_3954,N_3970);
nor U4027 (N_4027,N_3946,N_3917);
nand U4028 (N_4028,N_3936,N_3980);
or U4029 (N_4029,N_3944,N_3963);
or U4030 (N_4030,N_3950,N_3961);
nor U4031 (N_4031,N_3987,N_3906);
or U4032 (N_4032,N_3942,N_3951);
xnor U4033 (N_4033,N_3968,N_3912);
and U4034 (N_4034,N_3922,N_3935);
and U4035 (N_4035,N_3907,N_3934);
nor U4036 (N_4036,N_3908,N_3955);
nand U4037 (N_4037,N_3967,N_3998);
xnor U4038 (N_4038,N_3989,N_3960);
nor U4039 (N_4039,N_3902,N_3952);
xnor U4040 (N_4040,N_3916,N_3962);
nand U4041 (N_4041,N_3919,N_3911);
and U4042 (N_4042,N_3985,N_3997);
and U4043 (N_4043,N_3976,N_3957);
nor U4044 (N_4044,N_3964,N_3905);
or U4045 (N_4045,N_3981,N_3928);
or U4046 (N_4046,N_3937,N_3973);
nand U4047 (N_4047,N_3972,N_3971);
nand U4048 (N_4048,N_3969,N_3977);
nor U4049 (N_4049,N_3943,N_3925);
or U4050 (N_4050,N_3991,N_3939);
nand U4051 (N_4051,N_3947,N_3918);
or U4052 (N_4052,N_3905,N_3982);
nand U4053 (N_4053,N_3916,N_3967);
nor U4054 (N_4054,N_3983,N_3982);
or U4055 (N_4055,N_3999,N_3944);
nand U4056 (N_4056,N_3999,N_3920);
and U4057 (N_4057,N_3990,N_3920);
and U4058 (N_4058,N_3924,N_3948);
xor U4059 (N_4059,N_3934,N_3966);
nand U4060 (N_4060,N_3968,N_3929);
and U4061 (N_4061,N_3907,N_3944);
nor U4062 (N_4062,N_3969,N_3979);
and U4063 (N_4063,N_3902,N_3945);
or U4064 (N_4064,N_3994,N_3989);
nor U4065 (N_4065,N_3927,N_3914);
nor U4066 (N_4066,N_3963,N_3968);
nand U4067 (N_4067,N_3912,N_3903);
nand U4068 (N_4068,N_3928,N_3965);
nor U4069 (N_4069,N_3990,N_3939);
and U4070 (N_4070,N_3939,N_3960);
nor U4071 (N_4071,N_3943,N_3920);
xnor U4072 (N_4072,N_3968,N_3922);
xnor U4073 (N_4073,N_3944,N_3900);
xor U4074 (N_4074,N_3902,N_3965);
or U4075 (N_4075,N_3938,N_3907);
nor U4076 (N_4076,N_3980,N_3953);
and U4077 (N_4077,N_3949,N_3959);
xor U4078 (N_4078,N_3993,N_3906);
nand U4079 (N_4079,N_3996,N_3915);
nand U4080 (N_4080,N_3958,N_3963);
nor U4081 (N_4081,N_3952,N_3970);
nand U4082 (N_4082,N_3938,N_3906);
or U4083 (N_4083,N_3909,N_3997);
or U4084 (N_4084,N_3913,N_3944);
xnor U4085 (N_4085,N_3903,N_3989);
nand U4086 (N_4086,N_3994,N_3944);
xor U4087 (N_4087,N_3946,N_3935);
nand U4088 (N_4088,N_3929,N_3909);
nor U4089 (N_4089,N_3981,N_3993);
or U4090 (N_4090,N_3994,N_3909);
nor U4091 (N_4091,N_3923,N_3909);
xnor U4092 (N_4092,N_3901,N_3917);
nor U4093 (N_4093,N_3948,N_3916);
and U4094 (N_4094,N_3940,N_3929);
and U4095 (N_4095,N_3912,N_3901);
xor U4096 (N_4096,N_3929,N_3902);
nor U4097 (N_4097,N_3945,N_3994);
and U4098 (N_4098,N_3904,N_3989);
and U4099 (N_4099,N_3934,N_3981);
nand U4100 (N_4100,N_4005,N_4031);
xnor U4101 (N_4101,N_4030,N_4080);
and U4102 (N_4102,N_4078,N_4083);
xnor U4103 (N_4103,N_4082,N_4054);
nand U4104 (N_4104,N_4048,N_4000);
nand U4105 (N_4105,N_4029,N_4015);
xnor U4106 (N_4106,N_4088,N_4095);
or U4107 (N_4107,N_4017,N_4035);
and U4108 (N_4108,N_4072,N_4009);
and U4109 (N_4109,N_4039,N_4026);
and U4110 (N_4110,N_4075,N_4014);
xnor U4111 (N_4111,N_4069,N_4057);
and U4112 (N_4112,N_4013,N_4033);
nand U4113 (N_4113,N_4018,N_4068);
xnor U4114 (N_4114,N_4047,N_4093);
nand U4115 (N_4115,N_4003,N_4024);
or U4116 (N_4116,N_4043,N_4086);
xnor U4117 (N_4117,N_4051,N_4040);
or U4118 (N_4118,N_4099,N_4049);
and U4119 (N_4119,N_4085,N_4044);
nor U4120 (N_4120,N_4073,N_4037);
nand U4121 (N_4121,N_4089,N_4012);
or U4122 (N_4122,N_4076,N_4045);
nor U4123 (N_4123,N_4041,N_4027);
xor U4124 (N_4124,N_4058,N_4036);
xor U4125 (N_4125,N_4021,N_4008);
xor U4126 (N_4126,N_4087,N_4066);
nand U4127 (N_4127,N_4010,N_4016);
and U4128 (N_4128,N_4067,N_4074);
nor U4129 (N_4129,N_4096,N_4065);
xor U4130 (N_4130,N_4055,N_4052);
and U4131 (N_4131,N_4056,N_4060);
xnor U4132 (N_4132,N_4002,N_4053);
or U4133 (N_4133,N_4090,N_4071);
and U4134 (N_4134,N_4022,N_4064);
nand U4135 (N_4135,N_4025,N_4011);
xnor U4136 (N_4136,N_4092,N_4028);
xnor U4137 (N_4137,N_4050,N_4001);
nor U4138 (N_4138,N_4019,N_4020);
nor U4139 (N_4139,N_4038,N_4077);
nand U4140 (N_4140,N_4070,N_4006);
nand U4141 (N_4141,N_4097,N_4084);
xnor U4142 (N_4142,N_4032,N_4098);
nand U4143 (N_4143,N_4059,N_4007);
or U4144 (N_4144,N_4094,N_4023);
xnor U4145 (N_4145,N_4046,N_4061);
nor U4146 (N_4146,N_4081,N_4062);
xnor U4147 (N_4147,N_4034,N_4004);
xor U4148 (N_4148,N_4079,N_4091);
or U4149 (N_4149,N_4063,N_4042);
and U4150 (N_4150,N_4050,N_4058);
nand U4151 (N_4151,N_4051,N_4062);
nand U4152 (N_4152,N_4043,N_4009);
nand U4153 (N_4153,N_4017,N_4096);
nor U4154 (N_4154,N_4024,N_4011);
or U4155 (N_4155,N_4076,N_4009);
or U4156 (N_4156,N_4028,N_4032);
and U4157 (N_4157,N_4007,N_4051);
nor U4158 (N_4158,N_4031,N_4017);
nor U4159 (N_4159,N_4003,N_4011);
nand U4160 (N_4160,N_4038,N_4013);
and U4161 (N_4161,N_4042,N_4083);
nand U4162 (N_4162,N_4035,N_4037);
nand U4163 (N_4163,N_4004,N_4069);
xor U4164 (N_4164,N_4018,N_4002);
and U4165 (N_4165,N_4055,N_4080);
xnor U4166 (N_4166,N_4078,N_4010);
and U4167 (N_4167,N_4090,N_4096);
and U4168 (N_4168,N_4055,N_4019);
nand U4169 (N_4169,N_4057,N_4021);
and U4170 (N_4170,N_4004,N_4051);
xnor U4171 (N_4171,N_4020,N_4074);
nand U4172 (N_4172,N_4074,N_4030);
xor U4173 (N_4173,N_4064,N_4002);
nor U4174 (N_4174,N_4042,N_4039);
and U4175 (N_4175,N_4086,N_4015);
nand U4176 (N_4176,N_4025,N_4061);
xor U4177 (N_4177,N_4038,N_4035);
nor U4178 (N_4178,N_4071,N_4065);
nor U4179 (N_4179,N_4040,N_4085);
nor U4180 (N_4180,N_4018,N_4053);
and U4181 (N_4181,N_4034,N_4077);
nand U4182 (N_4182,N_4067,N_4071);
nand U4183 (N_4183,N_4005,N_4067);
and U4184 (N_4184,N_4062,N_4025);
and U4185 (N_4185,N_4091,N_4096);
xor U4186 (N_4186,N_4032,N_4017);
or U4187 (N_4187,N_4082,N_4027);
nand U4188 (N_4188,N_4082,N_4067);
and U4189 (N_4189,N_4074,N_4076);
nor U4190 (N_4190,N_4055,N_4000);
and U4191 (N_4191,N_4030,N_4032);
nor U4192 (N_4192,N_4097,N_4059);
nor U4193 (N_4193,N_4077,N_4000);
xnor U4194 (N_4194,N_4024,N_4057);
nor U4195 (N_4195,N_4062,N_4015);
xor U4196 (N_4196,N_4093,N_4022);
xor U4197 (N_4197,N_4088,N_4087);
xor U4198 (N_4198,N_4080,N_4041);
and U4199 (N_4199,N_4077,N_4009);
and U4200 (N_4200,N_4103,N_4179);
nand U4201 (N_4201,N_4107,N_4133);
and U4202 (N_4202,N_4169,N_4161);
and U4203 (N_4203,N_4122,N_4194);
nand U4204 (N_4204,N_4130,N_4191);
nor U4205 (N_4205,N_4146,N_4125);
nor U4206 (N_4206,N_4104,N_4168);
or U4207 (N_4207,N_4147,N_4105);
nor U4208 (N_4208,N_4118,N_4190);
nand U4209 (N_4209,N_4123,N_4158);
nand U4210 (N_4210,N_4184,N_4143);
nand U4211 (N_4211,N_4198,N_4135);
xnor U4212 (N_4212,N_4185,N_4154);
xnor U4213 (N_4213,N_4129,N_4121);
nand U4214 (N_4214,N_4116,N_4138);
nor U4215 (N_4215,N_4100,N_4127);
xnor U4216 (N_4216,N_4112,N_4176);
xnor U4217 (N_4217,N_4163,N_4150);
and U4218 (N_4218,N_4132,N_4145);
and U4219 (N_4219,N_4165,N_4126);
or U4220 (N_4220,N_4114,N_4196);
nor U4221 (N_4221,N_4111,N_4110);
nand U4222 (N_4222,N_4128,N_4120);
and U4223 (N_4223,N_4136,N_4144);
xnor U4224 (N_4224,N_4164,N_4181);
nand U4225 (N_4225,N_4137,N_4152);
xor U4226 (N_4226,N_4109,N_4160);
and U4227 (N_4227,N_4173,N_4124);
or U4228 (N_4228,N_4119,N_4195);
nor U4229 (N_4229,N_4140,N_4186);
and U4230 (N_4230,N_4167,N_4102);
or U4231 (N_4231,N_4180,N_4166);
and U4232 (N_4232,N_4157,N_4178);
or U4233 (N_4233,N_4156,N_4101);
nand U4234 (N_4234,N_4131,N_4188);
xnor U4235 (N_4235,N_4199,N_4189);
xnor U4236 (N_4236,N_4149,N_4108);
nor U4237 (N_4237,N_4187,N_4197);
xor U4238 (N_4238,N_4106,N_4171);
nand U4239 (N_4239,N_4175,N_4155);
or U4240 (N_4240,N_4162,N_4153);
and U4241 (N_4241,N_4183,N_4115);
nand U4242 (N_4242,N_4141,N_4177);
and U4243 (N_4243,N_4113,N_4192);
nand U4244 (N_4244,N_4193,N_4170);
nor U4245 (N_4245,N_4151,N_4139);
or U4246 (N_4246,N_4159,N_4174);
nand U4247 (N_4247,N_4148,N_4142);
and U4248 (N_4248,N_4182,N_4117);
nor U4249 (N_4249,N_4134,N_4172);
and U4250 (N_4250,N_4126,N_4110);
or U4251 (N_4251,N_4119,N_4155);
nand U4252 (N_4252,N_4182,N_4131);
nand U4253 (N_4253,N_4128,N_4183);
xor U4254 (N_4254,N_4181,N_4115);
or U4255 (N_4255,N_4126,N_4114);
xnor U4256 (N_4256,N_4129,N_4137);
nand U4257 (N_4257,N_4177,N_4127);
nor U4258 (N_4258,N_4167,N_4161);
or U4259 (N_4259,N_4196,N_4192);
or U4260 (N_4260,N_4185,N_4194);
or U4261 (N_4261,N_4175,N_4125);
nand U4262 (N_4262,N_4115,N_4193);
nor U4263 (N_4263,N_4192,N_4141);
xor U4264 (N_4264,N_4177,N_4170);
and U4265 (N_4265,N_4145,N_4179);
or U4266 (N_4266,N_4174,N_4129);
xor U4267 (N_4267,N_4149,N_4113);
xor U4268 (N_4268,N_4107,N_4167);
xor U4269 (N_4269,N_4177,N_4153);
nand U4270 (N_4270,N_4165,N_4174);
or U4271 (N_4271,N_4143,N_4154);
xnor U4272 (N_4272,N_4177,N_4130);
nand U4273 (N_4273,N_4198,N_4161);
nor U4274 (N_4274,N_4145,N_4184);
or U4275 (N_4275,N_4135,N_4151);
xor U4276 (N_4276,N_4141,N_4153);
and U4277 (N_4277,N_4132,N_4163);
nand U4278 (N_4278,N_4189,N_4197);
nand U4279 (N_4279,N_4133,N_4115);
xnor U4280 (N_4280,N_4162,N_4113);
nor U4281 (N_4281,N_4190,N_4181);
and U4282 (N_4282,N_4129,N_4194);
or U4283 (N_4283,N_4170,N_4187);
xor U4284 (N_4284,N_4152,N_4167);
nor U4285 (N_4285,N_4162,N_4182);
xor U4286 (N_4286,N_4130,N_4152);
nor U4287 (N_4287,N_4157,N_4167);
nor U4288 (N_4288,N_4127,N_4139);
or U4289 (N_4289,N_4160,N_4105);
nand U4290 (N_4290,N_4134,N_4109);
and U4291 (N_4291,N_4132,N_4104);
nand U4292 (N_4292,N_4169,N_4186);
xor U4293 (N_4293,N_4127,N_4194);
nand U4294 (N_4294,N_4169,N_4115);
nor U4295 (N_4295,N_4121,N_4183);
nor U4296 (N_4296,N_4155,N_4144);
nand U4297 (N_4297,N_4179,N_4104);
nor U4298 (N_4298,N_4168,N_4159);
xor U4299 (N_4299,N_4156,N_4102);
nor U4300 (N_4300,N_4292,N_4210);
or U4301 (N_4301,N_4212,N_4218);
or U4302 (N_4302,N_4236,N_4233);
and U4303 (N_4303,N_4260,N_4201);
and U4304 (N_4304,N_4223,N_4208);
or U4305 (N_4305,N_4246,N_4207);
xnor U4306 (N_4306,N_4248,N_4272);
and U4307 (N_4307,N_4221,N_4261);
nand U4308 (N_4308,N_4295,N_4269);
and U4309 (N_4309,N_4251,N_4265);
nor U4310 (N_4310,N_4284,N_4226);
and U4311 (N_4311,N_4296,N_4200);
nor U4312 (N_4312,N_4298,N_4242);
xnor U4313 (N_4313,N_4277,N_4270);
and U4314 (N_4314,N_4254,N_4288);
xor U4315 (N_4315,N_4234,N_4282);
and U4316 (N_4316,N_4204,N_4243);
and U4317 (N_4317,N_4262,N_4287);
nor U4318 (N_4318,N_4253,N_4294);
or U4319 (N_4319,N_4273,N_4241);
xor U4320 (N_4320,N_4203,N_4299);
and U4321 (N_4321,N_4216,N_4297);
nand U4322 (N_4322,N_4258,N_4228);
and U4323 (N_4323,N_4263,N_4214);
nor U4324 (N_4324,N_4283,N_4281);
xnor U4325 (N_4325,N_4259,N_4245);
nand U4326 (N_4326,N_4229,N_4264);
or U4327 (N_4327,N_4250,N_4202);
and U4328 (N_4328,N_4222,N_4211);
nor U4329 (N_4329,N_4285,N_4225);
nand U4330 (N_4330,N_4240,N_4231);
or U4331 (N_4331,N_4268,N_4266);
nor U4332 (N_4332,N_4235,N_4252);
or U4333 (N_4333,N_4232,N_4255);
or U4334 (N_4334,N_4293,N_4230);
or U4335 (N_4335,N_4206,N_4205);
nor U4336 (N_4336,N_4279,N_4276);
nand U4337 (N_4337,N_4215,N_4239);
or U4338 (N_4338,N_4220,N_4249);
nand U4339 (N_4339,N_4244,N_4289);
or U4340 (N_4340,N_4271,N_4209);
and U4341 (N_4341,N_4257,N_4227);
or U4342 (N_4342,N_4286,N_4278);
nor U4343 (N_4343,N_4224,N_4238);
nand U4344 (N_4344,N_4267,N_4274);
xor U4345 (N_4345,N_4217,N_4213);
or U4346 (N_4346,N_4256,N_4275);
xnor U4347 (N_4347,N_4247,N_4280);
nor U4348 (N_4348,N_4237,N_4291);
nand U4349 (N_4349,N_4290,N_4219);
and U4350 (N_4350,N_4271,N_4267);
and U4351 (N_4351,N_4250,N_4278);
xnor U4352 (N_4352,N_4285,N_4287);
nand U4353 (N_4353,N_4284,N_4251);
and U4354 (N_4354,N_4244,N_4256);
xor U4355 (N_4355,N_4225,N_4286);
or U4356 (N_4356,N_4217,N_4282);
xor U4357 (N_4357,N_4279,N_4273);
nor U4358 (N_4358,N_4253,N_4254);
xnor U4359 (N_4359,N_4270,N_4298);
xnor U4360 (N_4360,N_4204,N_4241);
nand U4361 (N_4361,N_4229,N_4280);
xnor U4362 (N_4362,N_4298,N_4246);
nor U4363 (N_4363,N_4263,N_4265);
xor U4364 (N_4364,N_4202,N_4225);
or U4365 (N_4365,N_4291,N_4211);
and U4366 (N_4366,N_4214,N_4202);
nor U4367 (N_4367,N_4203,N_4211);
or U4368 (N_4368,N_4282,N_4218);
or U4369 (N_4369,N_4234,N_4200);
xor U4370 (N_4370,N_4279,N_4292);
and U4371 (N_4371,N_4236,N_4293);
and U4372 (N_4372,N_4289,N_4208);
nand U4373 (N_4373,N_4207,N_4211);
and U4374 (N_4374,N_4287,N_4295);
xor U4375 (N_4375,N_4250,N_4219);
nor U4376 (N_4376,N_4227,N_4204);
nand U4377 (N_4377,N_4290,N_4238);
or U4378 (N_4378,N_4260,N_4228);
xnor U4379 (N_4379,N_4269,N_4224);
nand U4380 (N_4380,N_4227,N_4203);
and U4381 (N_4381,N_4236,N_4284);
xnor U4382 (N_4382,N_4280,N_4203);
nand U4383 (N_4383,N_4260,N_4278);
xor U4384 (N_4384,N_4231,N_4216);
nor U4385 (N_4385,N_4220,N_4269);
nor U4386 (N_4386,N_4271,N_4228);
or U4387 (N_4387,N_4226,N_4263);
or U4388 (N_4388,N_4265,N_4231);
nand U4389 (N_4389,N_4284,N_4254);
and U4390 (N_4390,N_4296,N_4294);
nand U4391 (N_4391,N_4243,N_4276);
or U4392 (N_4392,N_4233,N_4281);
or U4393 (N_4393,N_4237,N_4295);
nand U4394 (N_4394,N_4255,N_4219);
or U4395 (N_4395,N_4282,N_4276);
nor U4396 (N_4396,N_4288,N_4296);
xor U4397 (N_4397,N_4207,N_4283);
nand U4398 (N_4398,N_4272,N_4232);
nor U4399 (N_4399,N_4270,N_4287);
or U4400 (N_4400,N_4368,N_4314);
nand U4401 (N_4401,N_4301,N_4327);
and U4402 (N_4402,N_4325,N_4382);
or U4403 (N_4403,N_4311,N_4387);
nor U4404 (N_4404,N_4338,N_4397);
nand U4405 (N_4405,N_4320,N_4391);
xnor U4406 (N_4406,N_4303,N_4329);
and U4407 (N_4407,N_4335,N_4394);
xnor U4408 (N_4408,N_4376,N_4362);
xor U4409 (N_4409,N_4356,N_4318);
and U4410 (N_4410,N_4332,N_4324);
nor U4411 (N_4411,N_4313,N_4399);
nand U4412 (N_4412,N_4305,N_4331);
nor U4413 (N_4413,N_4352,N_4380);
xnor U4414 (N_4414,N_4349,N_4328);
nor U4415 (N_4415,N_4348,N_4340);
nand U4416 (N_4416,N_4389,N_4393);
nor U4417 (N_4417,N_4341,N_4396);
or U4418 (N_4418,N_4386,N_4321);
or U4419 (N_4419,N_4359,N_4373);
nor U4420 (N_4420,N_4343,N_4361);
nor U4421 (N_4421,N_4322,N_4315);
xor U4422 (N_4422,N_4358,N_4388);
xnor U4423 (N_4423,N_4308,N_4304);
or U4424 (N_4424,N_4367,N_4385);
nand U4425 (N_4425,N_4354,N_4383);
xnor U4426 (N_4426,N_4323,N_4379);
xnor U4427 (N_4427,N_4330,N_4317);
and U4428 (N_4428,N_4370,N_4363);
nor U4429 (N_4429,N_4319,N_4344);
or U4430 (N_4430,N_4339,N_4381);
or U4431 (N_4431,N_4395,N_4398);
nand U4432 (N_4432,N_4374,N_4347);
xor U4433 (N_4433,N_4364,N_4337);
nand U4434 (N_4434,N_4372,N_4355);
or U4435 (N_4435,N_4357,N_4366);
or U4436 (N_4436,N_4316,N_4351);
or U4437 (N_4437,N_4378,N_4336);
nand U4438 (N_4438,N_4300,N_4353);
xnor U4439 (N_4439,N_4345,N_4334);
nor U4440 (N_4440,N_4384,N_4309);
nor U4441 (N_4441,N_4306,N_4342);
and U4442 (N_4442,N_4369,N_4326);
xor U4443 (N_4443,N_4371,N_4360);
and U4444 (N_4444,N_4312,N_4375);
nand U4445 (N_4445,N_4377,N_4365);
or U4446 (N_4446,N_4350,N_4392);
or U4447 (N_4447,N_4310,N_4307);
xor U4448 (N_4448,N_4333,N_4302);
xnor U4449 (N_4449,N_4390,N_4346);
and U4450 (N_4450,N_4356,N_4383);
and U4451 (N_4451,N_4335,N_4355);
nor U4452 (N_4452,N_4354,N_4353);
or U4453 (N_4453,N_4356,N_4320);
or U4454 (N_4454,N_4367,N_4318);
nor U4455 (N_4455,N_4358,N_4329);
or U4456 (N_4456,N_4308,N_4364);
nand U4457 (N_4457,N_4368,N_4331);
and U4458 (N_4458,N_4307,N_4322);
or U4459 (N_4459,N_4367,N_4357);
xnor U4460 (N_4460,N_4304,N_4320);
nor U4461 (N_4461,N_4394,N_4349);
nor U4462 (N_4462,N_4304,N_4374);
and U4463 (N_4463,N_4393,N_4352);
nor U4464 (N_4464,N_4389,N_4306);
nand U4465 (N_4465,N_4315,N_4346);
nor U4466 (N_4466,N_4315,N_4328);
nand U4467 (N_4467,N_4311,N_4394);
or U4468 (N_4468,N_4381,N_4397);
xor U4469 (N_4469,N_4303,N_4359);
nor U4470 (N_4470,N_4305,N_4377);
or U4471 (N_4471,N_4361,N_4369);
and U4472 (N_4472,N_4398,N_4370);
nor U4473 (N_4473,N_4359,N_4327);
or U4474 (N_4474,N_4349,N_4336);
xor U4475 (N_4475,N_4304,N_4397);
nor U4476 (N_4476,N_4396,N_4306);
or U4477 (N_4477,N_4390,N_4374);
nand U4478 (N_4478,N_4370,N_4329);
xnor U4479 (N_4479,N_4309,N_4317);
nand U4480 (N_4480,N_4361,N_4394);
nand U4481 (N_4481,N_4302,N_4349);
nor U4482 (N_4482,N_4306,N_4339);
nand U4483 (N_4483,N_4347,N_4353);
or U4484 (N_4484,N_4364,N_4370);
and U4485 (N_4485,N_4304,N_4314);
nor U4486 (N_4486,N_4308,N_4374);
nor U4487 (N_4487,N_4372,N_4398);
or U4488 (N_4488,N_4339,N_4328);
and U4489 (N_4489,N_4352,N_4355);
or U4490 (N_4490,N_4303,N_4317);
or U4491 (N_4491,N_4385,N_4357);
or U4492 (N_4492,N_4395,N_4302);
nor U4493 (N_4493,N_4368,N_4339);
xnor U4494 (N_4494,N_4362,N_4380);
xnor U4495 (N_4495,N_4314,N_4391);
xnor U4496 (N_4496,N_4321,N_4318);
xnor U4497 (N_4497,N_4384,N_4371);
xor U4498 (N_4498,N_4382,N_4338);
and U4499 (N_4499,N_4356,N_4373);
nor U4500 (N_4500,N_4484,N_4479);
nand U4501 (N_4501,N_4451,N_4472);
and U4502 (N_4502,N_4415,N_4439);
nand U4503 (N_4503,N_4475,N_4447);
nand U4504 (N_4504,N_4490,N_4488);
xnor U4505 (N_4505,N_4403,N_4455);
nand U4506 (N_4506,N_4492,N_4464);
and U4507 (N_4507,N_4431,N_4453);
nand U4508 (N_4508,N_4494,N_4471);
nand U4509 (N_4509,N_4468,N_4449);
nand U4510 (N_4510,N_4427,N_4441);
xor U4511 (N_4511,N_4485,N_4409);
nor U4512 (N_4512,N_4426,N_4493);
and U4513 (N_4513,N_4466,N_4470);
nor U4514 (N_4514,N_4477,N_4436);
nor U4515 (N_4515,N_4498,N_4499);
nand U4516 (N_4516,N_4440,N_4419);
nand U4517 (N_4517,N_4423,N_4486);
or U4518 (N_4518,N_4474,N_4465);
nor U4519 (N_4519,N_4401,N_4489);
or U4520 (N_4520,N_4448,N_4462);
xor U4521 (N_4521,N_4428,N_4432);
and U4522 (N_4522,N_4481,N_4483);
xor U4523 (N_4523,N_4458,N_4445);
and U4524 (N_4524,N_4480,N_4411);
or U4525 (N_4525,N_4429,N_4405);
nor U4526 (N_4526,N_4482,N_4418);
or U4527 (N_4527,N_4421,N_4438);
and U4528 (N_4528,N_4495,N_4469);
xnor U4529 (N_4529,N_4491,N_4460);
nand U4530 (N_4530,N_4412,N_4446);
nand U4531 (N_4531,N_4414,N_4463);
or U4532 (N_4532,N_4422,N_4457);
nand U4533 (N_4533,N_4476,N_4400);
nor U4534 (N_4534,N_4487,N_4443);
nand U4535 (N_4535,N_4424,N_4473);
nor U4536 (N_4536,N_4410,N_4406);
nor U4537 (N_4537,N_4433,N_4452);
xnor U4538 (N_4538,N_4408,N_4454);
xor U4539 (N_4539,N_4478,N_4496);
or U4540 (N_4540,N_4413,N_4425);
xnor U4541 (N_4541,N_4416,N_4444);
and U4542 (N_4542,N_4407,N_4456);
xnor U4543 (N_4543,N_4434,N_4417);
or U4544 (N_4544,N_4404,N_4450);
xor U4545 (N_4545,N_4497,N_4402);
or U4546 (N_4546,N_4442,N_4437);
xor U4547 (N_4547,N_4420,N_4430);
and U4548 (N_4548,N_4467,N_4461);
xnor U4549 (N_4549,N_4435,N_4459);
xor U4550 (N_4550,N_4401,N_4415);
xor U4551 (N_4551,N_4458,N_4418);
or U4552 (N_4552,N_4409,N_4446);
or U4553 (N_4553,N_4479,N_4439);
nand U4554 (N_4554,N_4409,N_4451);
nor U4555 (N_4555,N_4435,N_4416);
or U4556 (N_4556,N_4463,N_4440);
nand U4557 (N_4557,N_4436,N_4465);
or U4558 (N_4558,N_4487,N_4488);
nand U4559 (N_4559,N_4499,N_4460);
nand U4560 (N_4560,N_4419,N_4406);
or U4561 (N_4561,N_4491,N_4478);
nand U4562 (N_4562,N_4481,N_4447);
nor U4563 (N_4563,N_4442,N_4448);
nand U4564 (N_4564,N_4485,N_4448);
nor U4565 (N_4565,N_4459,N_4444);
and U4566 (N_4566,N_4430,N_4483);
and U4567 (N_4567,N_4400,N_4491);
xor U4568 (N_4568,N_4454,N_4402);
nor U4569 (N_4569,N_4473,N_4466);
nand U4570 (N_4570,N_4415,N_4419);
xor U4571 (N_4571,N_4492,N_4407);
or U4572 (N_4572,N_4452,N_4439);
xor U4573 (N_4573,N_4403,N_4482);
and U4574 (N_4574,N_4499,N_4471);
xnor U4575 (N_4575,N_4490,N_4412);
xor U4576 (N_4576,N_4425,N_4490);
nor U4577 (N_4577,N_4417,N_4488);
xor U4578 (N_4578,N_4408,N_4400);
nor U4579 (N_4579,N_4443,N_4451);
and U4580 (N_4580,N_4467,N_4485);
nor U4581 (N_4581,N_4433,N_4435);
xor U4582 (N_4582,N_4473,N_4432);
and U4583 (N_4583,N_4490,N_4496);
and U4584 (N_4584,N_4494,N_4424);
nand U4585 (N_4585,N_4432,N_4497);
nand U4586 (N_4586,N_4437,N_4422);
xnor U4587 (N_4587,N_4487,N_4484);
nand U4588 (N_4588,N_4489,N_4498);
and U4589 (N_4589,N_4462,N_4498);
and U4590 (N_4590,N_4473,N_4429);
and U4591 (N_4591,N_4488,N_4443);
or U4592 (N_4592,N_4463,N_4408);
nand U4593 (N_4593,N_4482,N_4453);
xnor U4594 (N_4594,N_4471,N_4444);
xor U4595 (N_4595,N_4433,N_4466);
and U4596 (N_4596,N_4491,N_4408);
or U4597 (N_4597,N_4428,N_4493);
nand U4598 (N_4598,N_4463,N_4491);
or U4599 (N_4599,N_4492,N_4456);
xnor U4600 (N_4600,N_4581,N_4579);
or U4601 (N_4601,N_4573,N_4517);
and U4602 (N_4602,N_4525,N_4587);
or U4603 (N_4603,N_4531,N_4553);
and U4604 (N_4604,N_4535,N_4541);
or U4605 (N_4605,N_4500,N_4582);
or U4606 (N_4606,N_4536,N_4518);
xnor U4607 (N_4607,N_4542,N_4556);
or U4608 (N_4608,N_4598,N_4578);
xnor U4609 (N_4609,N_4569,N_4585);
nand U4610 (N_4610,N_4508,N_4543);
xnor U4611 (N_4611,N_4515,N_4549);
or U4612 (N_4612,N_4564,N_4562);
and U4613 (N_4613,N_4575,N_4552);
nand U4614 (N_4614,N_4540,N_4557);
xor U4615 (N_4615,N_4572,N_4513);
nor U4616 (N_4616,N_4593,N_4561);
nand U4617 (N_4617,N_4589,N_4588);
nand U4618 (N_4618,N_4584,N_4506);
and U4619 (N_4619,N_4574,N_4546);
xnor U4620 (N_4620,N_4591,N_4566);
xor U4621 (N_4621,N_4519,N_4505);
nor U4622 (N_4622,N_4567,N_4512);
nor U4623 (N_4623,N_4528,N_4597);
xor U4624 (N_4624,N_4510,N_4570);
nand U4625 (N_4625,N_4547,N_4560);
xnor U4626 (N_4626,N_4555,N_4568);
or U4627 (N_4627,N_4559,N_4521);
or U4628 (N_4628,N_4599,N_4580);
nor U4629 (N_4629,N_4533,N_4595);
nor U4630 (N_4630,N_4522,N_4550);
xnor U4631 (N_4631,N_4503,N_4594);
nor U4632 (N_4632,N_4534,N_4526);
xnor U4633 (N_4633,N_4523,N_4509);
and U4634 (N_4634,N_4545,N_4596);
xor U4635 (N_4635,N_4544,N_4576);
xor U4636 (N_4636,N_4592,N_4502);
and U4637 (N_4637,N_4507,N_4551);
and U4638 (N_4638,N_4558,N_4548);
nand U4639 (N_4639,N_4563,N_4537);
or U4640 (N_4640,N_4554,N_4516);
and U4641 (N_4641,N_4524,N_4577);
and U4642 (N_4642,N_4539,N_4520);
xnor U4643 (N_4643,N_4571,N_4583);
and U4644 (N_4644,N_4511,N_4504);
nor U4645 (N_4645,N_4501,N_4586);
or U4646 (N_4646,N_4590,N_4529);
and U4647 (N_4647,N_4565,N_4532);
nor U4648 (N_4648,N_4538,N_4530);
nand U4649 (N_4649,N_4527,N_4514);
nor U4650 (N_4650,N_4592,N_4575);
and U4651 (N_4651,N_4539,N_4568);
and U4652 (N_4652,N_4510,N_4529);
and U4653 (N_4653,N_4531,N_4525);
nand U4654 (N_4654,N_4546,N_4576);
and U4655 (N_4655,N_4558,N_4531);
xnor U4656 (N_4656,N_4526,N_4523);
nand U4657 (N_4657,N_4516,N_4507);
and U4658 (N_4658,N_4526,N_4539);
or U4659 (N_4659,N_4563,N_4574);
nand U4660 (N_4660,N_4554,N_4587);
or U4661 (N_4661,N_4501,N_4522);
nor U4662 (N_4662,N_4590,N_4557);
nor U4663 (N_4663,N_4587,N_4593);
nor U4664 (N_4664,N_4573,N_4570);
xnor U4665 (N_4665,N_4560,N_4519);
or U4666 (N_4666,N_4527,N_4568);
xor U4667 (N_4667,N_4539,N_4565);
xor U4668 (N_4668,N_4561,N_4518);
or U4669 (N_4669,N_4536,N_4554);
xor U4670 (N_4670,N_4536,N_4575);
nor U4671 (N_4671,N_4566,N_4584);
xor U4672 (N_4672,N_4580,N_4571);
nand U4673 (N_4673,N_4503,N_4599);
nor U4674 (N_4674,N_4574,N_4529);
or U4675 (N_4675,N_4538,N_4583);
and U4676 (N_4676,N_4540,N_4570);
nand U4677 (N_4677,N_4522,N_4540);
nor U4678 (N_4678,N_4516,N_4536);
or U4679 (N_4679,N_4540,N_4577);
nor U4680 (N_4680,N_4564,N_4592);
xor U4681 (N_4681,N_4523,N_4539);
and U4682 (N_4682,N_4549,N_4588);
nand U4683 (N_4683,N_4580,N_4538);
and U4684 (N_4684,N_4527,N_4511);
nand U4685 (N_4685,N_4541,N_4558);
or U4686 (N_4686,N_4553,N_4514);
nand U4687 (N_4687,N_4544,N_4594);
nand U4688 (N_4688,N_4564,N_4529);
or U4689 (N_4689,N_4525,N_4576);
or U4690 (N_4690,N_4510,N_4501);
xor U4691 (N_4691,N_4577,N_4569);
xor U4692 (N_4692,N_4548,N_4595);
nor U4693 (N_4693,N_4586,N_4525);
or U4694 (N_4694,N_4538,N_4599);
xnor U4695 (N_4695,N_4560,N_4589);
nand U4696 (N_4696,N_4522,N_4586);
nor U4697 (N_4697,N_4549,N_4586);
or U4698 (N_4698,N_4538,N_4568);
or U4699 (N_4699,N_4565,N_4524);
nand U4700 (N_4700,N_4624,N_4682);
xnor U4701 (N_4701,N_4671,N_4684);
or U4702 (N_4702,N_4689,N_4664);
xnor U4703 (N_4703,N_4652,N_4635);
or U4704 (N_4704,N_4687,N_4677);
xnor U4705 (N_4705,N_4606,N_4608);
nor U4706 (N_4706,N_4618,N_4640);
nor U4707 (N_4707,N_4633,N_4655);
xnor U4708 (N_4708,N_4601,N_4648);
and U4709 (N_4709,N_4627,N_4673);
nor U4710 (N_4710,N_4649,N_4676);
or U4711 (N_4711,N_4637,N_4607);
nor U4712 (N_4712,N_4678,N_4629);
nor U4713 (N_4713,N_4628,N_4642);
nand U4714 (N_4714,N_4656,N_4644);
nor U4715 (N_4715,N_4612,N_4668);
and U4716 (N_4716,N_4679,N_4638);
or U4717 (N_4717,N_4603,N_4681);
xnor U4718 (N_4718,N_4670,N_4696);
and U4719 (N_4719,N_4672,N_4699);
nand U4720 (N_4720,N_4695,N_4625);
xnor U4721 (N_4721,N_4643,N_4667);
nor U4722 (N_4722,N_4659,N_4663);
xor U4723 (N_4723,N_4657,N_4630);
nor U4724 (N_4724,N_4661,N_4680);
nand U4725 (N_4725,N_4675,N_4662);
nor U4726 (N_4726,N_4639,N_4604);
and U4727 (N_4727,N_4688,N_4613);
and U4728 (N_4728,N_4686,N_4611);
xor U4729 (N_4729,N_4653,N_4691);
and U4730 (N_4730,N_4622,N_4623);
or U4731 (N_4731,N_4626,N_4654);
or U4732 (N_4732,N_4647,N_4698);
nor U4733 (N_4733,N_4660,N_4692);
or U4734 (N_4734,N_4600,N_4634);
and U4735 (N_4735,N_4669,N_4645);
nand U4736 (N_4736,N_4614,N_4641);
nor U4737 (N_4737,N_4621,N_4685);
xor U4738 (N_4738,N_4619,N_4651);
xor U4739 (N_4739,N_4694,N_4615);
or U4740 (N_4740,N_4674,N_4650);
xnor U4741 (N_4741,N_4690,N_4631);
xor U4742 (N_4742,N_4616,N_4693);
nor U4743 (N_4743,N_4610,N_4632);
or U4744 (N_4744,N_4697,N_4617);
xor U4745 (N_4745,N_4620,N_4605);
xnor U4746 (N_4746,N_4683,N_4658);
and U4747 (N_4747,N_4646,N_4602);
nand U4748 (N_4748,N_4665,N_4666);
and U4749 (N_4749,N_4609,N_4636);
and U4750 (N_4750,N_4642,N_4651);
nor U4751 (N_4751,N_4603,N_4653);
or U4752 (N_4752,N_4689,N_4665);
and U4753 (N_4753,N_4642,N_4647);
nand U4754 (N_4754,N_4631,N_4620);
nand U4755 (N_4755,N_4630,N_4642);
or U4756 (N_4756,N_4687,N_4650);
nor U4757 (N_4757,N_4672,N_4652);
xnor U4758 (N_4758,N_4664,N_4615);
nor U4759 (N_4759,N_4680,N_4671);
nor U4760 (N_4760,N_4663,N_4680);
xnor U4761 (N_4761,N_4665,N_4641);
nand U4762 (N_4762,N_4665,N_4656);
or U4763 (N_4763,N_4671,N_4652);
xor U4764 (N_4764,N_4645,N_4639);
and U4765 (N_4765,N_4698,N_4674);
or U4766 (N_4766,N_4639,N_4653);
or U4767 (N_4767,N_4689,N_4610);
nor U4768 (N_4768,N_4699,N_4634);
or U4769 (N_4769,N_4617,N_4698);
or U4770 (N_4770,N_4602,N_4615);
nand U4771 (N_4771,N_4609,N_4689);
nor U4772 (N_4772,N_4629,N_4686);
nand U4773 (N_4773,N_4696,N_4675);
nor U4774 (N_4774,N_4640,N_4654);
and U4775 (N_4775,N_4664,N_4674);
nor U4776 (N_4776,N_4616,N_4678);
xor U4777 (N_4777,N_4687,N_4662);
nor U4778 (N_4778,N_4671,N_4618);
nand U4779 (N_4779,N_4619,N_4627);
xor U4780 (N_4780,N_4658,N_4679);
nor U4781 (N_4781,N_4603,N_4650);
xnor U4782 (N_4782,N_4680,N_4690);
xnor U4783 (N_4783,N_4610,N_4658);
xnor U4784 (N_4784,N_4632,N_4654);
xor U4785 (N_4785,N_4642,N_4679);
xor U4786 (N_4786,N_4679,N_4625);
nand U4787 (N_4787,N_4696,N_4639);
xnor U4788 (N_4788,N_4647,N_4673);
nand U4789 (N_4789,N_4626,N_4646);
and U4790 (N_4790,N_4699,N_4651);
or U4791 (N_4791,N_4617,N_4677);
and U4792 (N_4792,N_4695,N_4637);
or U4793 (N_4793,N_4642,N_4653);
nor U4794 (N_4794,N_4673,N_4684);
or U4795 (N_4795,N_4625,N_4612);
or U4796 (N_4796,N_4632,N_4643);
nand U4797 (N_4797,N_4624,N_4633);
and U4798 (N_4798,N_4690,N_4627);
xor U4799 (N_4799,N_4671,N_4638);
xnor U4800 (N_4800,N_4762,N_4766);
nor U4801 (N_4801,N_4749,N_4733);
xor U4802 (N_4802,N_4750,N_4759);
nor U4803 (N_4803,N_4702,N_4710);
and U4804 (N_4804,N_4752,N_4707);
nand U4805 (N_4805,N_4793,N_4700);
or U4806 (N_4806,N_4796,N_4753);
and U4807 (N_4807,N_4774,N_4747);
xnor U4808 (N_4808,N_4716,N_4737);
nand U4809 (N_4809,N_4731,N_4756);
and U4810 (N_4810,N_4730,N_4776);
xnor U4811 (N_4811,N_4771,N_4738);
nor U4812 (N_4812,N_4721,N_4719);
nor U4813 (N_4813,N_4703,N_4792);
or U4814 (N_4814,N_4798,N_4727);
or U4815 (N_4815,N_4763,N_4795);
nor U4816 (N_4816,N_4781,N_4757);
and U4817 (N_4817,N_4787,N_4754);
xor U4818 (N_4818,N_4728,N_4726);
nor U4819 (N_4819,N_4736,N_4785);
or U4820 (N_4820,N_4718,N_4797);
nor U4821 (N_4821,N_4723,N_4709);
and U4822 (N_4822,N_4745,N_4777);
and U4823 (N_4823,N_4715,N_4765);
or U4824 (N_4824,N_4742,N_4729);
and U4825 (N_4825,N_4712,N_4734);
nor U4826 (N_4826,N_4770,N_4780);
nand U4827 (N_4827,N_4751,N_4741);
xnor U4828 (N_4828,N_4739,N_4768);
or U4829 (N_4829,N_4720,N_4782);
nor U4830 (N_4830,N_4794,N_4708);
xor U4831 (N_4831,N_4732,N_4713);
and U4832 (N_4832,N_4778,N_4786);
xor U4833 (N_4833,N_4748,N_4724);
or U4834 (N_4834,N_4784,N_4744);
and U4835 (N_4835,N_4779,N_4725);
nand U4836 (N_4836,N_4717,N_4722);
nand U4837 (N_4837,N_4764,N_4775);
xor U4838 (N_4838,N_4743,N_4714);
nor U4839 (N_4839,N_4791,N_4711);
nor U4840 (N_4840,N_4704,N_4760);
or U4841 (N_4841,N_4767,N_4746);
or U4842 (N_4842,N_4706,N_4788);
or U4843 (N_4843,N_4761,N_4758);
nor U4844 (N_4844,N_4701,N_4799);
or U4845 (N_4845,N_4783,N_4772);
and U4846 (N_4846,N_4705,N_4740);
nor U4847 (N_4847,N_4789,N_4769);
or U4848 (N_4848,N_4773,N_4755);
and U4849 (N_4849,N_4735,N_4790);
xnor U4850 (N_4850,N_4794,N_4757);
xnor U4851 (N_4851,N_4729,N_4773);
nand U4852 (N_4852,N_4759,N_4795);
nor U4853 (N_4853,N_4782,N_4735);
nand U4854 (N_4854,N_4736,N_4745);
nand U4855 (N_4855,N_4741,N_4716);
and U4856 (N_4856,N_4773,N_4754);
xnor U4857 (N_4857,N_4735,N_4759);
and U4858 (N_4858,N_4755,N_4718);
and U4859 (N_4859,N_4762,N_4775);
or U4860 (N_4860,N_4796,N_4744);
nor U4861 (N_4861,N_4727,N_4760);
nand U4862 (N_4862,N_4767,N_4786);
xnor U4863 (N_4863,N_4739,N_4726);
or U4864 (N_4864,N_4772,N_4793);
nand U4865 (N_4865,N_4727,N_4792);
or U4866 (N_4866,N_4793,N_4754);
nand U4867 (N_4867,N_4798,N_4760);
and U4868 (N_4868,N_4742,N_4782);
nand U4869 (N_4869,N_4719,N_4716);
nor U4870 (N_4870,N_4746,N_4785);
and U4871 (N_4871,N_4714,N_4751);
nand U4872 (N_4872,N_4717,N_4791);
nor U4873 (N_4873,N_4746,N_4773);
and U4874 (N_4874,N_4750,N_4725);
xor U4875 (N_4875,N_4767,N_4730);
nor U4876 (N_4876,N_4732,N_4755);
nor U4877 (N_4877,N_4744,N_4793);
or U4878 (N_4878,N_4798,N_4713);
nand U4879 (N_4879,N_4754,N_4771);
nand U4880 (N_4880,N_4743,N_4779);
or U4881 (N_4881,N_4716,N_4747);
or U4882 (N_4882,N_4792,N_4714);
nand U4883 (N_4883,N_4760,N_4796);
nand U4884 (N_4884,N_4727,N_4794);
and U4885 (N_4885,N_4799,N_4781);
nor U4886 (N_4886,N_4797,N_4713);
nand U4887 (N_4887,N_4732,N_4794);
xor U4888 (N_4888,N_4729,N_4706);
or U4889 (N_4889,N_4786,N_4723);
or U4890 (N_4890,N_4768,N_4780);
or U4891 (N_4891,N_4799,N_4774);
nor U4892 (N_4892,N_4766,N_4779);
and U4893 (N_4893,N_4792,N_4763);
and U4894 (N_4894,N_4720,N_4716);
or U4895 (N_4895,N_4719,N_4731);
nor U4896 (N_4896,N_4728,N_4770);
nor U4897 (N_4897,N_4716,N_4791);
and U4898 (N_4898,N_4702,N_4780);
xnor U4899 (N_4899,N_4769,N_4795);
xnor U4900 (N_4900,N_4840,N_4888);
xor U4901 (N_4901,N_4804,N_4864);
or U4902 (N_4902,N_4805,N_4865);
xor U4903 (N_4903,N_4829,N_4849);
nor U4904 (N_4904,N_4893,N_4841);
and U4905 (N_4905,N_4813,N_4842);
nor U4906 (N_4906,N_4837,N_4818);
or U4907 (N_4907,N_4800,N_4846);
or U4908 (N_4908,N_4814,N_4808);
and U4909 (N_4909,N_4873,N_4897);
nor U4910 (N_4910,N_4826,N_4882);
or U4911 (N_4911,N_4831,N_4879);
or U4912 (N_4912,N_4871,N_4896);
and U4913 (N_4913,N_4880,N_4861);
and U4914 (N_4914,N_4847,N_4899);
and U4915 (N_4915,N_4848,N_4884);
xnor U4916 (N_4916,N_4843,N_4824);
or U4917 (N_4917,N_4830,N_4870);
xnor U4918 (N_4918,N_4890,N_4892);
nor U4919 (N_4919,N_4869,N_4875);
and U4920 (N_4920,N_4801,N_4838);
or U4921 (N_4921,N_4860,N_4876);
nor U4922 (N_4922,N_4859,N_4817);
nand U4923 (N_4923,N_4878,N_4881);
nand U4924 (N_4924,N_4816,N_4812);
xnor U4925 (N_4925,N_4874,N_4809);
nor U4926 (N_4926,N_4839,N_4885);
and U4927 (N_4927,N_4827,N_4853);
xor U4928 (N_4928,N_4891,N_4807);
or U4929 (N_4929,N_4836,N_4866);
or U4930 (N_4930,N_4820,N_4811);
xnor U4931 (N_4931,N_4886,N_4889);
and U4932 (N_4932,N_4823,N_4858);
or U4933 (N_4933,N_4803,N_4851);
nand U4934 (N_4934,N_4825,N_4822);
nand U4935 (N_4935,N_4821,N_4855);
nand U4936 (N_4936,N_4835,N_4898);
and U4937 (N_4937,N_4856,N_4852);
nand U4938 (N_4938,N_4867,N_4834);
nand U4939 (N_4939,N_4877,N_4862);
or U4940 (N_4940,N_4883,N_4844);
or U4941 (N_4941,N_4868,N_4895);
and U4942 (N_4942,N_4872,N_4894);
and U4943 (N_4943,N_4815,N_4887);
nor U4944 (N_4944,N_4828,N_4857);
nor U4945 (N_4945,N_4806,N_4863);
and U4946 (N_4946,N_4850,N_4854);
or U4947 (N_4947,N_4819,N_4832);
and U4948 (N_4948,N_4833,N_4802);
xor U4949 (N_4949,N_4845,N_4810);
or U4950 (N_4950,N_4876,N_4802);
xnor U4951 (N_4951,N_4863,N_4825);
nand U4952 (N_4952,N_4867,N_4820);
nor U4953 (N_4953,N_4873,N_4840);
nor U4954 (N_4954,N_4816,N_4837);
and U4955 (N_4955,N_4826,N_4866);
or U4956 (N_4956,N_4867,N_4886);
nand U4957 (N_4957,N_4830,N_4848);
or U4958 (N_4958,N_4820,N_4876);
or U4959 (N_4959,N_4846,N_4869);
nand U4960 (N_4960,N_4858,N_4872);
and U4961 (N_4961,N_4869,N_4882);
nand U4962 (N_4962,N_4835,N_4895);
xor U4963 (N_4963,N_4888,N_4886);
xor U4964 (N_4964,N_4841,N_4803);
or U4965 (N_4965,N_4857,N_4812);
xnor U4966 (N_4966,N_4885,N_4815);
nor U4967 (N_4967,N_4856,N_4815);
nand U4968 (N_4968,N_4870,N_4833);
and U4969 (N_4969,N_4889,N_4854);
nand U4970 (N_4970,N_4895,N_4882);
nand U4971 (N_4971,N_4858,N_4827);
or U4972 (N_4972,N_4832,N_4812);
nand U4973 (N_4973,N_4880,N_4876);
nand U4974 (N_4974,N_4817,N_4825);
nor U4975 (N_4975,N_4893,N_4882);
and U4976 (N_4976,N_4820,N_4890);
nor U4977 (N_4977,N_4811,N_4882);
and U4978 (N_4978,N_4836,N_4805);
or U4979 (N_4979,N_4877,N_4872);
and U4980 (N_4980,N_4803,N_4868);
and U4981 (N_4981,N_4823,N_4894);
and U4982 (N_4982,N_4802,N_4819);
and U4983 (N_4983,N_4849,N_4863);
nor U4984 (N_4984,N_4827,N_4816);
or U4985 (N_4985,N_4853,N_4868);
nor U4986 (N_4986,N_4852,N_4807);
xnor U4987 (N_4987,N_4808,N_4894);
nor U4988 (N_4988,N_4811,N_4891);
xnor U4989 (N_4989,N_4840,N_4825);
xnor U4990 (N_4990,N_4886,N_4843);
xor U4991 (N_4991,N_4895,N_4864);
nor U4992 (N_4992,N_4834,N_4891);
nor U4993 (N_4993,N_4859,N_4882);
nor U4994 (N_4994,N_4865,N_4835);
and U4995 (N_4995,N_4841,N_4882);
xor U4996 (N_4996,N_4879,N_4865);
and U4997 (N_4997,N_4881,N_4857);
nand U4998 (N_4998,N_4873,N_4841);
xor U4999 (N_4999,N_4884,N_4809);
and U5000 (N_5000,N_4931,N_4970);
and U5001 (N_5001,N_4999,N_4975);
nor U5002 (N_5002,N_4966,N_4945);
xor U5003 (N_5003,N_4994,N_4983);
and U5004 (N_5004,N_4910,N_4992);
nand U5005 (N_5005,N_4958,N_4996);
and U5006 (N_5006,N_4932,N_4965);
xnor U5007 (N_5007,N_4969,N_4972);
nor U5008 (N_5008,N_4933,N_4959);
and U5009 (N_5009,N_4955,N_4985);
nand U5010 (N_5010,N_4976,N_4963);
nor U5011 (N_5011,N_4989,N_4977);
and U5012 (N_5012,N_4938,N_4913);
or U5013 (N_5013,N_4902,N_4939);
xor U5014 (N_5014,N_4952,N_4928);
or U5015 (N_5015,N_4988,N_4949);
xor U5016 (N_5016,N_4917,N_4914);
nand U5017 (N_5017,N_4923,N_4919);
or U5018 (N_5018,N_4986,N_4922);
and U5019 (N_5019,N_4995,N_4912);
and U5020 (N_5020,N_4968,N_4906);
and U5021 (N_5021,N_4901,N_4903);
nand U5022 (N_5022,N_4964,N_4991);
xnor U5023 (N_5023,N_4926,N_4984);
xnor U5024 (N_5024,N_4918,N_4971);
or U5025 (N_5025,N_4925,N_4947);
xor U5026 (N_5026,N_4920,N_4907);
and U5027 (N_5027,N_4993,N_4909);
xnor U5028 (N_5028,N_4905,N_4944);
nand U5029 (N_5029,N_4997,N_4921);
and U5030 (N_5030,N_4911,N_4973);
xor U5031 (N_5031,N_4908,N_4904);
xor U5032 (N_5032,N_4946,N_4967);
and U5033 (N_5033,N_4962,N_4951);
or U5034 (N_5034,N_4974,N_4934);
or U5035 (N_5035,N_4915,N_4940);
or U5036 (N_5036,N_4987,N_4980);
nor U5037 (N_5037,N_4998,N_4957);
nand U5038 (N_5038,N_4982,N_4930);
and U5039 (N_5039,N_4954,N_4929);
nor U5040 (N_5040,N_4953,N_4937);
and U5041 (N_5041,N_4927,N_4979);
nor U5042 (N_5042,N_4956,N_4942);
nor U5043 (N_5043,N_4924,N_4935);
or U5044 (N_5044,N_4990,N_4948);
nor U5045 (N_5045,N_4941,N_4900);
nand U5046 (N_5046,N_4981,N_4936);
or U5047 (N_5047,N_4950,N_4916);
and U5048 (N_5048,N_4961,N_4943);
nor U5049 (N_5049,N_4978,N_4960);
or U5050 (N_5050,N_4986,N_4961);
nand U5051 (N_5051,N_4933,N_4950);
nand U5052 (N_5052,N_4921,N_4902);
and U5053 (N_5053,N_4932,N_4954);
nor U5054 (N_5054,N_4979,N_4992);
or U5055 (N_5055,N_4950,N_4939);
and U5056 (N_5056,N_4984,N_4925);
nand U5057 (N_5057,N_4955,N_4975);
and U5058 (N_5058,N_4943,N_4902);
nand U5059 (N_5059,N_4920,N_4980);
nand U5060 (N_5060,N_4998,N_4939);
or U5061 (N_5061,N_4947,N_4915);
xnor U5062 (N_5062,N_4941,N_4999);
xnor U5063 (N_5063,N_4976,N_4946);
nor U5064 (N_5064,N_4915,N_4921);
nand U5065 (N_5065,N_4969,N_4965);
nand U5066 (N_5066,N_4948,N_4962);
xor U5067 (N_5067,N_4966,N_4919);
and U5068 (N_5068,N_4978,N_4996);
and U5069 (N_5069,N_4966,N_4928);
nor U5070 (N_5070,N_4929,N_4983);
and U5071 (N_5071,N_4987,N_4974);
nor U5072 (N_5072,N_4955,N_4996);
xor U5073 (N_5073,N_4919,N_4978);
and U5074 (N_5074,N_4925,N_4992);
nor U5075 (N_5075,N_4924,N_4988);
and U5076 (N_5076,N_4987,N_4972);
or U5077 (N_5077,N_4916,N_4930);
xnor U5078 (N_5078,N_4951,N_4958);
or U5079 (N_5079,N_4905,N_4902);
or U5080 (N_5080,N_4984,N_4966);
xnor U5081 (N_5081,N_4942,N_4935);
and U5082 (N_5082,N_4905,N_4926);
nand U5083 (N_5083,N_4916,N_4992);
and U5084 (N_5084,N_4943,N_4956);
and U5085 (N_5085,N_4919,N_4903);
nand U5086 (N_5086,N_4984,N_4956);
and U5087 (N_5087,N_4920,N_4975);
nor U5088 (N_5088,N_4942,N_4905);
xor U5089 (N_5089,N_4932,N_4918);
xnor U5090 (N_5090,N_4951,N_4996);
nand U5091 (N_5091,N_4994,N_4966);
and U5092 (N_5092,N_4919,N_4902);
nand U5093 (N_5093,N_4963,N_4968);
xor U5094 (N_5094,N_4939,N_4983);
xnor U5095 (N_5095,N_4934,N_4978);
nand U5096 (N_5096,N_4977,N_4992);
and U5097 (N_5097,N_4949,N_4978);
nor U5098 (N_5098,N_4953,N_4947);
and U5099 (N_5099,N_4969,N_4961);
or U5100 (N_5100,N_5028,N_5065);
and U5101 (N_5101,N_5085,N_5052);
or U5102 (N_5102,N_5054,N_5095);
nand U5103 (N_5103,N_5006,N_5036);
nand U5104 (N_5104,N_5041,N_5045);
nor U5105 (N_5105,N_5059,N_5007);
nor U5106 (N_5106,N_5030,N_5068);
and U5107 (N_5107,N_5099,N_5023);
and U5108 (N_5108,N_5042,N_5035);
nand U5109 (N_5109,N_5015,N_5079);
nand U5110 (N_5110,N_5005,N_5093);
nor U5111 (N_5111,N_5062,N_5090);
nor U5112 (N_5112,N_5047,N_5040);
xnor U5113 (N_5113,N_5025,N_5021);
nor U5114 (N_5114,N_5001,N_5067);
nand U5115 (N_5115,N_5038,N_5027);
or U5116 (N_5116,N_5000,N_5034);
nor U5117 (N_5117,N_5071,N_5044);
nand U5118 (N_5118,N_5058,N_5018);
nand U5119 (N_5119,N_5072,N_5063);
and U5120 (N_5120,N_5024,N_5020);
and U5121 (N_5121,N_5009,N_5048);
nor U5122 (N_5122,N_5026,N_5051);
nand U5123 (N_5123,N_5012,N_5037);
nand U5124 (N_5124,N_5011,N_5076);
and U5125 (N_5125,N_5078,N_5003);
and U5126 (N_5126,N_5086,N_5089);
and U5127 (N_5127,N_5080,N_5096);
or U5128 (N_5128,N_5049,N_5031);
or U5129 (N_5129,N_5013,N_5097);
and U5130 (N_5130,N_5017,N_5060);
xor U5131 (N_5131,N_5056,N_5014);
xnor U5132 (N_5132,N_5091,N_5084);
xor U5133 (N_5133,N_5077,N_5088);
or U5134 (N_5134,N_5019,N_5055);
nand U5135 (N_5135,N_5075,N_5046);
xnor U5136 (N_5136,N_5004,N_5069);
xnor U5137 (N_5137,N_5033,N_5073);
and U5138 (N_5138,N_5032,N_5083);
nor U5139 (N_5139,N_5082,N_5022);
or U5140 (N_5140,N_5039,N_5081);
nand U5141 (N_5141,N_5050,N_5094);
nor U5142 (N_5142,N_5002,N_5043);
nand U5143 (N_5143,N_5029,N_5074);
or U5144 (N_5144,N_5010,N_5057);
nor U5145 (N_5145,N_5008,N_5098);
nor U5146 (N_5146,N_5064,N_5066);
and U5147 (N_5147,N_5087,N_5053);
nand U5148 (N_5148,N_5061,N_5016);
xnor U5149 (N_5149,N_5092,N_5070);
xnor U5150 (N_5150,N_5018,N_5066);
xor U5151 (N_5151,N_5068,N_5090);
nand U5152 (N_5152,N_5032,N_5031);
nand U5153 (N_5153,N_5022,N_5099);
xor U5154 (N_5154,N_5099,N_5089);
nand U5155 (N_5155,N_5098,N_5060);
nand U5156 (N_5156,N_5004,N_5029);
xnor U5157 (N_5157,N_5043,N_5088);
nor U5158 (N_5158,N_5077,N_5050);
nand U5159 (N_5159,N_5091,N_5043);
and U5160 (N_5160,N_5056,N_5091);
nor U5161 (N_5161,N_5086,N_5073);
nand U5162 (N_5162,N_5029,N_5013);
nand U5163 (N_5163,N_5085,N_5066);
xor U5164 (N_5164,N_5073,N_5042);
or U5165 (N_5165,N_5018,N_5091);
or U5166 (N_5166,N_5044,N_5094);
or U5167 (N_5167,N_5061,N_5081);
nand U5168 (N_5168,N_5093,N_5033);
nand U5169 (N_5169,N_5044,N_5028);
or U5170 (N_5170,N_5095,N_5055);
nand U5171 (N_5171,N_5081,N_5076);
nand U5172 (N_5172,N_5091,N_5058);
xor U5173 (N_5173,N_5040,N_5073);
xnor U5174 (N_5174,N_5046,N_5030);
xor U5175 (N_5175,N_5061,N_5022);
nor U5176 (N_5176,N_5012,N_5061);
xnor U5177 (N_5177,N_5024,N_5073);
and U5178 (N_5178,N_5060,N_5089);
nor U5179 (N_5179,N_5009,N_5073);
or U5180 (N_5180,N_5034,N_5018);
and U5181 (N_5181,N_5048,N_5089);
xor U5182 (N_5182,N_5083,N_5023);
or U5183 (N_5183,N_5080,N_5032);
nand U5184 (N_5184,N_5080,N_5068);
and U5185 (N_5185,N_5005,N_5047);
nand U5186 (N_5186,N_5098,N_5055);
nor U5187 (N_5187,N_5013,N_5033);
nor U5188 (N_5188,N_5062,N_5094);
nand U5189 (N_5189,N_5031,N_5062);
or U5190 (N_5190,N_5009,N_5041);
and U5191 (N_5191,N_5064,N_5035);
and U5192 (N_5192,N_5017,N_5077);
and U5193 (N_5193,N_5010,N_5066);
and U5194 (N_5194,N_5034,N_5096);
nor U5195 (N_5195,N_5038,N_5054);
xnor U5196 (N_5196,N_5092,N_5034);
xor U5197 (N_5197,N_5072,N_5045);
xnor U5198 (N_5198,N_5019,N_5012);
or U5199 (N_5199,N_5062,N_5084);
or U5200 (N_5200,N_5125,N_5173);
nor U5201 (N_5201,N_5186,N_5190);
xnor U5202 (N_5202,N_5110,N_5137);
nor U5203 (N_5203,N_5165,N_5181);
xor U5204 (N_5204,N_5164,N_5116);
or U5205 (N_5205,N_5168,N_5152);
and U5206 (N_5206,N_5189,N_5148);
xnor U5207 (N_5207,N_5182,N_5143);
nor U5208 (N_5208,N_5149,N_5160);
nor U5209 (N_5209,N_5145,N_5153);
nand U5210 (N_5210,N_5156,N_5107);
or U5211 (N_5211,N_5169,N_5151);
nand U5212 (N_5212,N_5159,N_5140);
xor U5213 (N_5213,N_5150,N_5119);
nor U5214 (N_5214,N_5141,N_5105);
xor U5215 (N_5215,N_5198,N_5127);
and U5216 (N_5216,N_5108,N_5100);
nor U5217 (N_5217,N_5128,N_5162);
or U5218 (N_5218,N_5183,N_5179);
xor U5219 (N_5219,N_5113,N_5187);
xor U5220 (N_5220,N_5139,N_5120);
or U5221 (N_5221,N_5178,N_5154);
nor U5222 (N_5222,N_5136,N_5191);
and U5223 (N_5223,N_5196,N_5163);
nand U5224 (N_5224,N_5170,N_5129);
or U5225 (N_5225,N_5114,N_5122);
and U5226 (N_5226,N_5177,N_5132);
or U5227 (N_5227,N_5197,N_5176);
nand U5228 (N_5228,N_5185,N_5171);
and U5229 (N_5229,N_5104,N_5193);
or U5230 (N_5230,N_5199,N_5123);
and U5231 (N_5231,N_5188,N_5133);
or U5232 (N_5232,N_5155,N_5130);
and U5233 (N_5233,N_5157,N_5134);
or U5234 (N_5234,N_5172,N_5106);
or U5235 (N_5235,N_5142,N_5112);
nor U5236 (N_5236,N_5109,N_5102);
xnor U5237 (N_5237,N_5118,N_5126);
xor U5238 (N_5238,N_5180,N_5124);
and U5239 (N_5239,N_5144,N_5167);
nand U5240 (N_5240,N_5174,N_5117);
and U5241 (N_5241,N_5175,N_5161);
and U5242 (N_5242,N_5103,N_5147);
and U5243 (N_5243,N_5111,N_5192);
or U5244 (N_5244,N_5131,N_5195);
and U5245 (N_5245,N_5166,N_5115);
or U5246 (N_5246,N_5135,N_5194);
nand U5247 (N_5247,N_5121,N_5138);
and U5248 (N_5248,N_5101,N_5184);
nor U5249 (N_5249,N_5158,N_5146);
nand U5250 (N_5250,N_5191,N_5164);
xnor U5251 (N_5251,N_5146,N_5121);
or U5252 (N_5252,N_5114,N_5193);
nand U5253 (N_5253,N_5138,N_5165);
and U5254 (N_5254,N_5155,N_5136);
xnor U5255 (N_5255,N_5129,N_5199);
xor U5256 (N_5256,N_5150,N_5111);
and U5257 (N_5257,N_5136,N_5119);
and U5258 (N_5258,N_5176,N_5133);
or U5259 (N_5259,N_5177,N_5122);
nor U5260 (N_5260,N_5101,N_5147);
or U5261 (N_5261,N_5180,N_5154);
nand U5262 (N_5262,N_5171,N_5174);
or U5263 (N_5263,N_5179,N_5109);
xnor U5264 (N_5264,N_5133,N_5178);
nand U5265 (N_5265,N_5197,N_5181);
or U5266 (N_5266,N_5158,N_5182);
xor U5267 (N_5267,N_5112,N_5189);
or U5268 (N_5268,N_5193,N_5124);
xor U5269 (N_5269,N_5193,N_5187);
nor U5270 (N_5270,N_5167,N_5183);
nor U5271 (N_5271,N_5148,N_5135);
and U5272 (N_5272,N_5153,N_5169);
and U5273 (N_5273,N_5166,N_5157);
or U5274 (N_5274,N_5181,N_5121);
nand U5275 (N_5275,N_5137,N_5128);
or U5276 (N_5276,N_5182,N_5175);
xnor U5277 (N_5277,N_5143,N_5159);
nand U5278 (N_5278,N_5112,N_5182);
or U5279 (N_5279,N_5138,N_5151);
and U5280 (N_5280,N_5152,N_5125);
or U5281 (N_5281,N_5164,N_5199);
xnor U5282 (N_5282,N_5176,N_5175);
nor U5283 (N_5283,N_5110,N_5103);
and U5284 (N_5284,N_5137,N_5194);
nand U5285 (N_5285,N_5183,N_5121);
nor U5286 (N_5286,N_5152,N_5167);
xnor U5287 (N_5287,N_5151,N_5176);
and U5288 (N_5288,N_5167,N_5190);
or U5289 (N_5289,N_5173,N_5121);
and U5290 (N_5290,N_5111,N_5117);
xnor U5291 (N_5291,N_5178,N_5140);
and U5292 (N_5292,N_5111,N_5102);
or U5293 (N_5293,N_5108,N_5180);
nand U5294 (N_5294,N_5181,N_5145);
or U5295 (N_5295,N_5109,N_5189);
and U5296 (N_5296,N_5187,N_5102);
xnor U5297 (N_5297,N_5146,N_5185);
xor U5298 (N_5298,N_5115,N_5169);
nand U5299 (N_5299,N_5133,N_5100);
and U5300 (N_5300,N_5263,N_5232);
nand U5301 (N_5301,N_5242,N_5211);
nand U5302 (N_5302,N_5249,N_5285);
or U5303 (N_5303,N_5216,N_5246);
nor U5304 (N_5304,N_5255,N_5258);
nand U5305 (N_5305,N_5239,N_5229);
and U5306 (N_5306,N_5218,N_5243);
or U5307 (N_5307,N_5270,N_5299);
or U5308 (N_5308,N_5212,N_5228);
or U5309 (N_5309,N_5259,N_5262);
or U5310 (N_5310,N_5296,N_5226);
or U5311 (N_5311,N_5222,N_5268);
xnor U5312 (N_5312,N_5292,N_5235);
or U5313 (N_5313,N_5207,N_5209);
or U5314 (N_5314,N_5294,N_5273);
nand U5315 (N_5315,N_5254,N_5298);
xnor U5316 (N_5316,N_5286,N_5213);
xor U5317 (N_5317,N_5274,N_5247);
or U5318 (N_5318,N_5215,N_5267);
xor U5319 (N_5319,N_5275,N_5225);
or U5320 (N_5320,N_5223,N_5276);
or U5321 (N_5321,N_5265,N_5236);
and U5322 (N_5322,N_5205,N_5260);
or U5323 (N_5323,N_5264,N_5250);
nand U5324 (N_5324,N_5269,N_5200);
nand U5325 (N_5325,N_5290,N_5234);
xnor U5326 (N_5326,N_5224,N_5214);
xnor U5327 (N_5327,N_5253,N_5245);
or U5328 (N_5328,N_5277,N_5256);
nor U5329 (N_5329,N_5271,N_5241);
nor U5330 (N_5330,N_5272,N_5201);
or U5331 (N_5331,N_5231,N_5293);
or U5332 (N_5332,N_5233,N_5281);
nand U5333 (N_5333,N_5221,N_5284);
xor U5334 (N_5334,N_5238,N_5278);
nor U5335 (N_5335,N_5251,N_5210);
xor U5336 (N_5336,N_5288,N_5206);
or U5337 (N_5337,N_5227,N_5204);
or U5338 (N_5338,N_5219,N_5230);
nand U5339 (N_5339,N_5282,N_5248);
nand U5340 (N_5340,N_5280,N_5297);
nand U5341 (N_5341,N_5287,N_5295);
and U5342 (N_5342,N_5217,N_5220);
nand U5343 (N_5343,N_5283,N_5240);
xor U5344 (N_5344,N_5261,N_5203);
nand U5345 (N_5345,N_5202,N_5291);
or U5346 (N_5346,N_5252,N_5208);
or U5347 (N_5347,N_5266,N_5244);
xnor U5348 (N_5348,N_5257,N_5237);
xor U5349 (N_5349,N_5289,N_5279);
xnor U5350 (N_5350,N_5256,N_5269);
or U5351 (N_5351,N_5299,N_5244);
nor U5352 (N_5352,N_5275,N_5252);
nor U5353 (N_5353,N_5235,N_5293);
or U5354 (N_5354,N_5282,N_5221);
xor U5355 (N_5355,N_5256,N_5234);
and U5356 (N_5356,N_5282,N_5289);
and U5357 (N_5357,N_5274,N_5281);
nor U5358 (N_5358,N_5205,N_5257);
and U5359 (N_5359,N_5202,N_5229);
xor U5360 (N_5360,N_5213,N_5212);
xnor U5361 (N_5361,N_5225,N_5210);
nor U5362 (N_5362,N_5285,N_5220);
xor U5363 (N_5363,N_5214,N_5256);
xnor U5364 (N_5364,N_5215,N_5277);
nor U5365 (N_5365,N_5266,N_5292);
nand U5366 (N_5366,N_5240,N_5251);
and U5367 (N_5367,N_5221,N_5256);
or U5368 (N_5368,N_5244,N_5227);
nand U5369 (N_5369,N_5281,N_5222);
nand U5370 (N_5370,N_5202,N_5285);
nor U5371 (N_5371,N_5269,N_5219);
or U5372 (N_5372,N_5274,N_5262);
nand U5373 (N_5373,N_5268,N_5261);
nor U5374 (N_5374,N_5218,N_5291);
or U5375 (N_5375,N_5296,N_5238);
or U5376 (N_5376,N_5230,N_5235);
and U5377 (N_5377,N_5204,N_5269);
and U5378 (N_5378,N_5252,N_5277);
xor U5379 (N_5379,N_5214,N_5282);
nor U5380 (N_5380,N_5293,N_5219);
nor U5381 (N_5381,N_5295,N_5224);
nand U5382 (N_5382,N_5288,N_5289);
and U5383 (N_5383,N_5225,N_5212);
or U5384 (N_5384,N_5246,N_5225);
nor U5385 (N_5385,N_5207,N_5228);
nand U5386 (N_5386,N_5260,N_5208);
nand U5387 (N_5387,N_5271,N_5257);
and U5388 (N_5388,N_5203,N_5281);
and U5389 (N_5389,N_5290,N_5276);
nor U5390 (N_5390,N_5293,N_5258);
nand U5391 (N_5391,N_5273,N_5252);
and U5392 (N_5392,N_5262,N_5208);
or U5393 (N_5393,N_5256,N_5223);
or U5394 (N_5394,N_5252,N_5289);
nor U5395 (N_5395,N_5212,N_5230);
nand U5396 (N_5396,N_5276,N_5247);
nor U5397 (N_5397,N_5244,N_5221);
nor U5398 (N_5398,N_5290,N_5210);
nor U5399 (N_5399,N_5243,N_5276);
and U5400 (N_5400,N_5389,N_5387);
nand U5401 (N_5401,N_5329,N_5364);
nand U5402 (N_5402,N_5340,N_5362);
or U5403 (N_5403,N_5302,N_5331);
xor U5404 (N_5404,N_5324,N_5306);
nor U5405 (N_5405,N_5383,N_5353);
nor U5406 (N_5406,N_5328,N_5349);
xnor U5407 (N_5407,N_5357,N_5337);
nor U5408 (N_5408,N_5333,N_5380);
nand U5409 (N_5409,N_5373,N_5393);
xor U5410 (N_5410,N_5348,N_5317);
xor U5411 (N_5411,N_5338,N_5304);
nor U5412 (N_5412,N_5351,N_5361);
nand U5413 (N_5413,N_5311,N_5371);
xnor U5414 (N_5414,N_5335,N_5355);
nor U5415 (N_5415,N_5326,N_5359);
or U5416 (N_5416,N_5346,N_5307);
and U5417 (N_5417,N_5342,N_5379);
or U5418 (N_5418,N_5367,N_5374);
xor U5419 (N_5419,N_5396,N_5310);
nor U5420 (N_5420,N_5345,N_5386);
or U5421 (N_5421,N_5382,N_5366);
nor U5422 (N_5422,N_5391,N_5316);
nor U5423 (N_5423,N_5365,N_5341);
nand U5424 (N_5424,N_5318,N_5325);
and U5425 (N_5425,N_5399,N_5301);
nand U5426 (N_5426,N_5336,N_5381);
nor U5427 (N_5427,N_5323,N_5384);
and U5428 (N_5428,N_5397,N_5352);
xor U5429 (N_5429,N_5305,N_5388);
nand U5430 (N_5430,N_5363,N_5358);
and U5431 (N_5431,N_5344,N_5360);
xor U5432 (N_5432,N_5370,N_5343);
or U5433 (N_5433,N_5375,N_5308);
nor U5434 (N_5434,N_5394,N_5369);
nand U5435 (N_5435,N_5315,N_5372);
nor U5436 (N_5436,N_5350,N_5303);
nand U5437 (N_5437,N_5327,N_5321);
xor U5438 (N_5438,N_5330,N_5300);
and U5439 (N_5439,N_5385,N_5377);
xor U5440 (N_5440,N_5322,N_5395);
and U5441 (N_5441,N_5313,N_5356);
xnor U5442 (N_5442,N_5354,N_5376);
nor U5443 (N_5443,N_5390,N_5314);
nor U5444 (N_5444,N_5309,N_5378);
or U5445 (N_5445,N_5398,N_5320);
nor U5446 (N_5446,N_5347,N_5339);
nor U5447 (N_5447,N_5392,N_5332);
nor U5448 (N_5448,N_5312,N_5368);
nand U5449 (N_5449,N_5319,N_5334);
or U5450 (N_5450,N_5330,N_5309);
nand U5451 (N_5451,N_5308,N_5324);
or U5452 (N_5452,N_5356,N_5399);
xnor U5453 (N_5453,N_5352,N_5310);
and U5454 (N_5454,N_5371,N_5338);
and U5455 (N_5455,N_5362,N_5325);
and U5456 (N_5456,N_5348,N_5391);
and U5457 (N_5457,N_5390,N_5307);
nor U5458 (N_5458,N_5392,N_5329);
xor U5459 (N_5459,N_5374,N_5359);
and U5460 (N_5460,N_5325,N_5305);
and U5461 (N_5461,N_5392,N_5365);
nor U5462 (N_5462,N_5395,N_5318);
xor U5463 (N_5463,N_5350,N_5325);
nand U5464 (N_5464,N_5353,N_5306);
or U5465 (N_5465,N_5300,N_5321);
or U5466 (N_5466,N_5374,N_5391);
xnor U5467 (N_5467,N_5328,N_5363);
or U5468 (N_5468,N_5392,N_5320);
or U5469 (N_5469,N_5338,N_5382);
nand U5470 (N_5470,N_5340,N_5343);
and U5471 (N_5471,N_5365,N_5324);
xnor U5472 (N_5472,N_5300,N_5390);
xor U5473 (N_5473,N_5390,N_5397);
xnor U5474 (N_5474,N_5300,N_5302);
or U5475 (N_5475,N_5323,N_5361);
nor U5476 (N_5476,N_5333,N_5323);
nand U5477 (N_5477,N_5309,N_5312);
nand U5478 (N_5478,N_5376,N_5383);
xor U5479 (N_5479,N_5319,N_5357);
or U5480 (N_5480,N_5305,N_5384);
and U5481 (N_5481,N_5394,N_5362);
xnor U5482 (N_5482,N_5354,N_5395);
and U5483 (N_5483,N_5305,N_5304);
or U5484 (N_5484,N_5387,N_5300);
nor U5485 (N_5485,N_5395,N_5368);
or U5486 (N_5486,N_5365,N_5337);
nand U5487 (N_5487,N_5323,N_5313);
nor U5488 (N_5488,N_5380,N_5353);
or U5489 (N_5489,N_5358,N_5338);
xor U5490 (N_5490,N_5399,N_5387);
nor U5491 (N_5491,N_5382,N_5349);
nand U5492 (N_5492,N_5353,N_5371);
and U5493 (N_5493,N_5352,N_5329);
xor U5494 (N_5494,N_5376,N_5364);
nand U5495 (N_5495,N_5373,N_5307);
and U5496 (N_5496,N_5393,N_5359);
nor U5497 (N_5497,N_5323,N_5325);
or U5498 (N_5498,N_5317,N_5382);
nor U5499 (N_5499,N_5303,N_5342);
nor U5500 (N_5500,N_5423,N_5440);
xor U5501 (N_5501,N_5467,N_5483);
xor U5502 (N_5502,N_5438,N_5452);
nor U5503 (N_5503,N_5471,N_5484);
or U5504 (N_5504,N_5458,N_5410);
nand U5505 (N_5505,N_5439,N_5492);
nor U5506 (N_5506,N_5480,N_5441);
nor U5507 (N_5507,N_5427,N_5488);
and U5508 (N_5508,N_5418,N_5494);
nand U5509 (N_5509,N_5422,N_5463);
nor U5510 (N_5510,N_5413,N_5434);
nor U5511 (N_5511,N_5495,N_5404);
or U5512 (N_5512,N_5490,N_5470);
and U5513 (N_5513,N_5474,N_5421);
xor U5514 (N_5514,N_5496,N_5444);
xnor U5515 (N_5515,N_5460,N_5411);
xnor U5516 (N_5516,N_5435,N_5402);
nor U5517 (N_5517,N_5445,N_5476);
nand U5518 (N_5518,N_5407,N_5455);
or U5519 (N_5519,N_5447,N_5469);
xnor U5520 (N_5520,N_5428,N_5465);
nand U5521 (N_5521,N_5481,N_5478);
and U5522 (N_5522,N_5457,N_5405);
xor U5523 (N_5523,N_5412,N_5482);
and U5524 (N_5524,N_5437,N_5449);
or U5525 (N_5525,N_5420,N_5448);
nor U5526 (N_5526,N_5400,N_5491);
nand U5527 (N_5527,N_5450,N_5406);
nand U5528 (N_5528,N_5433,N_5453);
nand U5529 (N_5529,N_5426,N_5485);
and U5530 (N_5530,N_5454,N_5416);
and U5531 (N_5531,N_5446,N_5489);
and U5532 (N_5532,N_5443,N_5464);
and U5533 (N_5533,N_5430,N_5409);
nor U5534 (N_5534,N_5415,N_5472);
or U5535 (N_5535,N_5493,N_5459);
and U5536 (N_5536,N_5408,N_5451);
nand U5537 (N_5537,N_5477,N_5431);
and U5538 (N_5538,N_5461,N_5429);
and U5539 (N_5539,N_5479,N_5486);
xnor U5540 (N_5540,N_5497,N_5403);
nor U5541 (N_5541,N_5499,N_5419);
and U5542 (N_5542,N_5473,N_5425);
nor U5543 (N_5543,N_5466,N_5475);
and U5544 (N_5544,N_5442,N_5498);
or U5545 (N_5545,N_5462,N_5414);
and U5546 (N_5546,N_5436,N_5401);
or U5547 (N_5547,N_5424,N_5417);
xor U5548 (N_5548,N_5487,N_5468);
xor U5549 (N_5549,N_5456,N_5432);
xnor U5550 (N_5550,N_5445,N_5477);
and U5551 (N_5551,N_5460,N_5447);
nor U5552 (N_5552,N_5467,N_5477);
nor U5553 (N_5553,N_5422,N_5452);
xnor U5554 (N_5554,N_5466,N_5400);
and U5555 (N_5555,N_5439,N_5442);
nand U5556 (N_5556,N_5468,N_5434);
nand U5557 (N_5557,N_5492,N_5431);
or U5558 (N_5558,N_5486,N_5440);
and U5559 (N_5559,N_5455,N_5453);
xnor U5560 (N_5560,N_5423,N_5421);
nor U5561 (N_5561,N_5404,N_5420);
xor U5562 (N_5562,N_5420,N_5443);
and U5563 (N_5563,N_5427,N_5432);
or U5564 (N_5564,N_5464,N_5472);
and U5565 (N_5565,N_5492,N_5406);
or U5566 (N_5566,N_5495,N_5480);
xnor U5567 (N_5567,N_5405,N_5420);
nor U5568 (N_5568,N_5480,N_5494);
and U5569 (N_5569,N_5429,N_5421);
and U5570 (N_5570,N_5414,N_5475);
and U5571 (N_5571,N_5437,N_5492);
and U5572 (N_5572,N_5403,N_5435);
or U5573 (N_5573,N_5457,N_5473);
nand U5574 (N_5574,N_5411,N_5463);
and U5575 (N_5575,N_5474,N_5497);
xor U5576 (N_5576,N_5429,N_5416);
and U5577 (N_5577,N_5498,N_5405);
nand U5578 (N_5578,N_5468,N_5485);
or U5579 (N_5579,N_5446,N_5481);
nand U5580 (N_5580,N_5427,N_5430);
nor U5581 (N_5581,N_5462,N_5472);
xnor U5582 (N_5582,N_5431,N_5476);
xnor U5583 (N_5583,N_5486,N_5498);
and U5584 (N_5584,N_5475,N_5490);
nor U5585 (N_5585,N_5428,N_5483);
nand U5586 (N_5586,N_5466,N_5477);
or U5587 (N_5587,N_5442,N_5424);
and U5588 (N_5588,N_5428,N_5438);
nand U5589 (N_5589,N_5454,N_5427);
xor U5590 (N_5590,N_5416,N_5442);
xnor U5591 (N_5591,N_5443,N_5423);
and U5592 (N_5592,N_5481,N_5453);
xor U5593 (N_5593,N_5455,N_5491);
nor U5594 (N_5594,N_5423,N_5412);
nor U5595 (N_5595,N_5426,N_5422);
nor U5596 (N_5596,N_5464,N_5496);
or U5597 (N_5597,N_5483,N_5474);
and U5598 (N_5598,N_5485,N_5492);
xor U5599 (N_5599,N_5440,N_5456);
and U5600 (N_5600,N_5589,N_5586);
nand U5601 (N_5601,N_5587,N_5503);
and U5602 (N_5602,N_5571,N_5561);
nor U5603 (N_5603,N_5551,N_5511);
nor U5604 (N_5604,N_5599,N_5550);
or U5605 (N_5605,N_5565,N_5575);
and U5606 (N_5606,N_5516,N_5553);
nand U5607 (N_5607,N_5596,N_5583);
nor U5608 (N_5608,N_5549,N_5527);
xor U5609 (N_5609,N_5534,N_5513);
xor U5610 (N_5610,N_5570,N_5555);
and U5611 (N_5611,N_5563,N_5522);
and U5612 (N_5612,N_5593,N_5548);
or U5613 (N_5613,N_5509,N_5542);
nor U5614 (N_5614,N_5526,N_5582);
or U5615 (N_5615,N_5559,N_5543);
and U5616 (N_5616,N_5584,N_5564);
xnor U5617 (N_5617,N_5541,N_5512);
nor U5618 (N_5618,N_5537,N_5544);
and U5619 (N_5619,N_5525,N_5528);
and U5620 (N_5620,N_5580,N_5501);
nand U5621 (N_5621,N_5560,N_5535);
xor U5622 (N_5622,N_5576,N_5556);
xor U5623 (N_5623,N_5500,N_5507);
and U5624 (N_5624,N_5569,N_5594);
nor U5625 (N_5625,N_5574,N_5505);
nor U5626 (N_5626,N_5538,N_5590);
or U5627 (N_5627,N_5572,N_5521);
nor U5628 (N_5628,N_5539,N_5519);
or U5629 (N_5629,N_5523,N_5531);
and U5630 (N_5630,N_5573,N_5545);
nand U5631 (N_5631,N_5529,N_5567);
xor U5632 (N_5632,N_5585,N_5536);
nor U5633 (N_5633,N_5524,N_5568);
nand U5634 (N_5634,N_5577,N_5562);
nor U5635 (N_5635,N_5515,N_5554);
nand U5636 (N_5636,N_5581,N_5557);
and U5637 (N_5637,N_5598,N_5504);
xnor U5638 (N_5638,N_5532,N_5578);
nand U5639 (N_5639,N_5558,N_5502);
or U5640 (N_5640,N_5591,N_5533);
nand U5641 (N_5641,N_5566,N_5547);
nor U5642 (N_5642,N_5592,N_5546);
nand U5643 (N_5643,N_5588,N_5520);
xnor U5644 (N_5644,N_5508,N_5597);
xnor U5645 (N_5645,N_5510,N_5518);
nor U5646 (N_5646,N_5517,N_5506);
and U5647 (N_5647,N_5514,N_5530);
nand U5648 (N_5648,N_5552,N_5540);
and U5649 (N_5649,N_5595,N_5579);
xnor U5650 (N_5650,N_5532,N_5503);
nor U5651 (N_5651,N_5504,N_5594);
nand U5652 (N_5652,N_5570,N_5513);
and U5653 (N_5653,N_5516,N_5554);
nand U5654 (N_5654,N_5529,N_5517);
nor U5655 (N_5655,N_5568,N_5503);
and U5656 (N_5656,N_5512,N_5577);
xnor U5657 (N_5657,N_5562,N_5586);
or U5658 (N_5658,N_5523,N_5589);
or U5659 (N_5659,N_5531,N_5534);
nor U5660 (N_5660,N_5513,N_5559);
nand U5661 (N_5661,N_5579,N_5572);
or U5662 (N_5662,N_5526,N_5585);
or U5663 (N_5663,N_5574,N_5542);
or U5664 (N_5664,N_5524,N_5506);
and U5665 (N_5665,N_5590,N_5552);
nand U5666 (N_5666,N_5575,N_5510);
xor U5667 (N_5667,N_5536,N_5533);
and U5668 (N_5668,N_5591,N_5585);
nor U5669 (N_5669,N_5535,N_5540);
and U5670 (N_5670,N_5549,N_5568);
nand U5671 (N_5671,N_5513,N_5535);
and U5672 (N_5672,N_5529,N_5574);
nor U5673 (N_5673,N_5559,N_5532);
nand U5674 (N_5674,N_5581,N_5597);
nor U5675 (N_5675,N_5507,N_5552);
nand U5676 (N_5676,N_5509,N_5501);
nand U5677 (N_5677,N_5506,N_5547);
or U5678 (N_5678,N_5516,N_5575);
nor U5679 (N_5679,N_5574,N_5593);
or U5680 (N_5680,N_5507,N_5504);
or U5681 (N_5681,N_5560,N_5516);
xnor U5682 (N_5682,N_5512,N_5537);
nand U5683 (N_5683,N_5511,N_5596);
xor U5684 (N_5684,N_5537,N_5594);
xor U5685 (N_5685,N_5544,N_5570);
nor U5686 (N_5686,N_5511,N_5520);
or U5687 (N_5687,N_5576,N_5551);
nand U5688 (N_5688,N_5572,N_5570);
nand U5689 (N_5689,N_5585,N_5555);
and U5690 (N_5690,N_5561,N_5528);
nor U5691 (N_5691,N_5539,N_5581);
nand U5692 (N_5692,N_5598,N_5517);
and U5693 (N_5693,N_5534,N_5566);
xor U5694 (N_5694,N_5587,N_5595);
xor U5695 (N_5695,N_5533,N_5584);
nor U5696 (N_5696,N_5595,N_5545);
xnor U5697 (N_5697,N_5516,N_5538);
nand U5698 (N_5698,N_5540,N_5584);
nand U5699 (N_5699,N_5552,N_5564);
or U5700 (N_5700,N_5618,N_5623);
and U5701 (N_5701,N_5692,N_5612);
nand U5702 (N_5702,N_5657,N_5636);
nand U5703 (N_5703,N_5676,N_5699);
xnor U5704 (N_5704,N_5640,N_5606);
nand U5705 (N_5705,N_5689,N_5629);
xnor U5706 (N_5706,N_5695,N_5675);
nor U5707 (N_5707,N_5674,N_5617);
nor U5708 (N_5708,N_5631,N_5652);
xnor U5709 (N_5709,N_5698,N_5609);
nand U5710 (N_5710,N_5682,N_5684);
or U5711 (N_5711,N_5634,N_5637);
xor U5712 (N_5712,N_5645,N_5690);
nand U5713 (N_5713,N_5646,N_5608);
or U5714 (N_5714,N_5626,N_5613);
nor U5715 (N_5715,N_5648,N_5678);
or U5716 (N_5716,N_5696,N_5615);
or U5717 (N_5717,N_5641,N_5662);
xnor U5718 (N_5718,N_5672,N_5654);
nor U5719 (N_5719,N_5611,N_5625);
xnor U5720 (N_5720,N_5603,N_5664);
xor U5721 (N_5721,N_5668,N_5681);
nand U5722 (N_5722,N_5663,N_5604);
xnor U5723 (N_5723,N_5644,N_5688);
xor U5724 (N_5724,N_5628,N_5694);
or U5725 (N_5725,N_5658,N_5660);
and U5726 (N_5726,N_5677,N_5622);
or U5727 (N_5727,N_5642,N_5627);
nand U5728 (N_5728,N_5614,N_5616);
or U5729 (N_5729,N_5638,N_5633);
nor U5730 (N_5730,N_5602,N_5630);
or U5731 (N_5731,N_5685,N_5621);
or U5732 (N_5732,N_5673,N_5635);
nor U5733 (N_5733,N_5686,N_5643);
nand U5734 (N_5734,N_5649,N_5651);
nor U5735 (N_5735,N_5632,N_5691);
or U5736 (N_5736,N_5661,N_5610);
or U5737 (N_5737,N_5679,N_5669);
and U5738 (N_5738,N_5620,N_5656);
xnor U5739 (N_5739,N_5601,N_5653);
nor U5740 (N_5740,N_5650,N_5666);
or U5741 (N_5741,N_5687,N_5639);
nor U5742 (N_5742,N_5665,N_5605);
nand U5743 (N_5743,N_5671,N_5693);
and U5744 (N_5744,N_5670,N_5619);
xnor U5745 (N_5745,N_5655,N_5683);
nor U5746 (N_5746,N_5659,N_5600);
or U5747 (N_5747,N_5667,N_5647);
xor U5748 (N_5748,N_5697,N_5607);
nand U5749 (N_5749,N_5680,N_5624);
and U5750 (N_5750,N_5637,N_5633);
nand U5751 (N_5751,N_5685,N_5637);
nand U5752 (N_5752,N_5634,N_5608);
and U5753 (N_5753,N_5626,N_5681);
nand U5754 (N_5754,N_5649,N_5658);
and U5755 (N_5755,N_5661,N_5658);
nand U5756 (N_5756,N_5618,N_5698);
nor U5757 (N_5757,N_5682,N_5612);
xnor U5758 (N_5758,N_5629,N_5601);
nand U5759 (N_5759,N_5617,N_5612);
xnor U5760 (N_5760,N_5698,N_5603);
and U5761 (N_5761,N_5692,N_5631);
or U5762 (N_5762,N_5613,N_5684);
and U5763 (N_5763,N_5636,N_5678);
and U5764 (N_5764,N_5674,N_5695);
or U5765 (N_5765,N_5696,N_5677);
xor U5766 (N_5766,N_5669,N_5657);
xor U5767 (N_5767,N_5653,N_5683);
and U5768 (N_5768,N_5681,N_5698);
or U5769 (N_5769,N_5628,N_5630);
xor U5770 (N_5770,N_5690,N_5608);
nor U5771 (N_5771,N_5615,N_5664);
nor U5772 (N_5772,N_5687,N_5669);
nor U5773 (N_5773,N_5606,N_5614);
nor U5774 (N_5774,N_5640,N_5674);
nor U5775 (N_5775,N_5605,N_5680);
xnor U5776 (N_5776,N_5684,N_5639);
nand U5777 (N_5777,N_5604,N_5623);
and U5778 (N_5778,N_5603,N_5622);
or U5779 (N_5779,N_5691,N_5636);
and U5780 (N_5780,N_5623,N_5642);
nand U5781 (N_5781,N_5698,N_5628);
or U5782 (N_5782,N_5625,N_5696);
and U5783 (N_5783,N_5670,N_5660);
xnor U5784 (N_5784,N_5676,N_5683);
nand U5785 (N_5785,N_5609,N_5693);
xor U5786 (N_5786,N_5616,N_5691);
and U5787 (N_5787,N_5699,N_5612);
nand U5788 (N_5788,N_5673,N_5617);
nand U5789 (N_5789,N_5603,N_5608);
nand U5790 (N_5790,N_5655,N_5631);
xor U5791 (N_5791,N_5643,N_5618);
nor U5792 (N_5792,N_5630,N_5647);
or U5793 (N_5793,N_5645,N_5668);
xnor U5794 (N_5794,N_5680,N_5633);
and U5795 (N_5795,N_5601,N_5628);
or U5796 (N_5796,N_5638,N_5676);
or U5797 (N_5797,N_5633,N_5614);
xor U5798 (N_5798,N_5652,N_5657);
nand U5799 (N_5799,N_5660,N_5662);
xor U5800 (N_5800,N_5700,N_5726);
nand U5801 (N_5801,N_5716,N_5729);
nor U5802 (N_5802,N_5754,N_5746);
xor U5803 (N_5803,N_5772,N_5723);
nor U5804 (N_5804,N_5705,N_5702);
and U5805 (N_5805,N_5712,N_5718);
xnor U5806 (N_5806,N_5794,N_5736);
nand U5807 (N_5807,N_5785,N_5721);
nor U5808 (N_5808,N_5713,N_5766);
nand U5809 (N_5809,N_5776,N_5792);
nor U5810 (N_5810,N_5780,N_5722);
and U5811 (N_5811,N_5737,N_5757);
or U5812 (N_5812,N_5724,N_5782);
and U5813 (N_5813,N_5743,N_5745);
nand U5814 (N_5814,N_5706,N_5731);
nand U5815 (N_5815,N_5799,N_5768);
or U5816 (N_5816,N_5742,N_5787);
or U5817 (N_5817,N_5781,N_5751);
and U5818 (N_5818,N_5786,N_5771);
and U5819 (N_5819,N_5725,N_5703);
nand U5820 (N_5820,N_5733,N_5773);
and U5821 (N_5821,N_5797,N_5789);
xor U5822 (N_5822,N_5748,N_5753);
or U5823 (N_5823,N_5719,N_5777);
nand U5824 (N_5824,N_5788,N_5714);
and U5825 (N_5825,N_5717,N_5784);
xor U5826 (N_5826,N_5738,N_5756);
and U5827 (N_5827,N_5730,N_5755);
or U5828 (N_5828,N_5798,N_5727);
or U5829 (N_5829,N_5759,N_5732);
nand U5830 (N_5830,N_5708,N_5711);
or U5831 (N_5831,N_5779,N_5762);
xnor U5832 (N_5832,N_5704,N_5761);
nand U5833 (N_5833,N_5752,N_5790);
nand U5834 (N_5834,N_5778,N_5774);
nor U5835 (N_5835,N_5765,N_5728);
xnor U5836 (N_5836,N_5739,N_5707);
nor U5837 (N_5837,N_5710,N_5796);
or U5838 (N_5838,N_5770,N_5741);
xnor U5839 (N_5839,N_5735,N_5734);
xor U5840 (N_5840,N_5769,N_5783);
or U5841 (N_5841,N_5709,N_5747);
and U5842 (N_5842,N_5744,N_5764);
nand U5843 (N_5843,N_5750,N_5763);
xnor U5844 (N_5844,N_5715,N_5760);
nand U5845 (N_5845,N_5758,N_5740);
nor U5846 (N_5846,N_5701,N_5767);
xnor U5847 (N_5847,N_5720,N_5791);
nand U5848 (N_5848,N_5749,N_5795);
or U5849 (N_5849,N_5793,N_5775);
and U5850 (N_5850,N_5742,N_5736);
nor U5851 (N_5851,N_5762,N_5712);
and U5852 (N_5852,N_5795,N_5731);
nand U5853 (N_5853,N_5743,N_5761);
nor U5854 (N_5854,N_5701,N_5745);
or U5855 (N_5855,N_5765,N_5774);
nor U5856 (N_5856,N_5722,N_5724);
and U5857 (N_5857,N_5783,N_5702);
nor U5858 (N_5858,N_5783,N_5740);
xor U5859 (N_5859,N_5750,N_5772);
nor U5860 (N_5860,N_5795,N_5746);
and U5861 (N_5861,N_5713,N_5725);
or U5862 (N_5862,N_5730,N_5769);
and U5863 (N_5863,N_5774,N_5794);
nand U5864 (N_5864,N_5781,N_5721);
nand U5865 (N_5865,N_5702,N_5794);
or U5866 (N_5866,N_5792,N_5745);
and U5867 (N_5867,N_5748,N_5787);
xnor U5868 (N_5868,N_5706,N_5716);
or U5869 (N_5869,N_5725,N_5795);
xnor U5870 (N_5870,N_5705,N_5723);
or U5871 (N_5871,N_5799,N_5772);
nand U5872 (N_5872,N_5757,N_5759);
nand U5873 (N_5873,N_5753,N_5719);
xnor U5874 (N_5874,N_5754,N_5724);
and U5875 (N_5875,N_5725,N_5773);
and U5876 (N_5876,N_5781,N_5717);
nand U5877 (N_5877,N_5724,N_5742);
or U5878 (N_5878,N_5767,N_5737);
nand U5879 (N_5879,N_5745,N_5766);
and U5880 (N_5880,N_5754,N_5740);
xnor U5881 (N_5881,N_5700,N_5799);
and U5882 (N_5882,N_5799,N_5732);
nor U5883 (N_5883,N_5794,N_5716);
xnor U5884 (N_5884,N_5761,N_5783);
nand U5885 (N_5885,N_5719,N_5756);
nand U5886 (N_5886,N_5713,N_5745);
nand U5887 (N_5887,N_5789,N_5710);
nor U5888 (N_5888,N_5733,N_5790);
nand U5889 (N_5889,N_5755,N_5780);
and U5890 (N_5890,N_5766,N_5799);
or U5891 (N_5891,N_5741,N_5703);
nand U5892 (N_5892,N_5783,N_5781);
nor U5893 (N_5893,N_5747,N_5713);
and U5894 (N_5894,N_5780,N_5735);
or U5895 (N_5895,N_5713,N_5789);
nor U5896 (N_5896,N_5708,N_5700);
nand U5897 (N_5897,N_5790,N_5714);
and U5898 (N_5898,N_5774,N_5759);
nand U5899 (N_5899,N_5710,N_5786);
nand U5900 (N_5900,N_5818,N_5826);
or U5901 (N_5901,N_5875,N_5829);
or U5902 (N_5902,N_5834,N_5827);
xor U5903 (N_5903,N_5858,N_5882);
nor U5904 (N_5904,N_5808,N_5844);
nor U5905 (N_5905,N_5821,N_5864);
nand U5906 (N_5906,N_5868,N_5837);
and U5907 (N_5907,N_5862,N_5895);
and U5908 (N_5908,N_5867,N_5846);
or U5909 (N_5909,N_5878,N_5804);
and U5910 (N_5910,N_5886,N_5812);
or U5911 (N_5911,N_5891,N_5876);
xor U5912 (N_5912,N_5887,N_5888);
nor U5913 (N_5913,N_5849,N_5847);
and U5914 (N_5914,N_5881,N_5838);
nand U5915 (N_5915,N_5832,N_5850);
xnor U5916 (N_5916,N_5820,N_5872);
xor U5917 (N_5917,N_5817,N_5885);
and U5918 (N_5918,N_5815,N_5880);
or U5919 (N_5919,N_5830,N_5800);
nor U5920 (N_5920,N_5842,N_5898);
and U5921 (N_5921,N_5874,N_5836);
xor U5922 (N_5922,N_5893,N_5890);
or U5923 (N_5923,N_5845,N_5828);
and U5924 (N_5924,N_5823,N_5816);
xnor U5925 (N_5925,N_5831,N_5883);
nor U5926 (N_5926,N_5896,N_5855);
nor U5927 (N_5927,N_5889,N_5839);
nand U5928 (N_5928,N_5869,N_5840);
and U5929 (N_5929,N_5835,N_5801);
xor U5930 (N_5930,N_5859,N_5825);
nand U5931 (N_5931,N_5810,N_5813);
nor U5932 (N_5932,N_5806,N_5852);
and U5933 (N_5933,N_5870,N_5877);
and U5934 (N_5934,N_5809,N_5841);
nor U5935 (N_5935,N_5848,N_5803);
and U5936 (N_5936,N_5860,N_5856);
nor U5937 (N_5937,N_5894,N_5805);
nand U5938 (N_5938,N_5814,N_5853);
xor U5939 (N_5939,N_5863,N_5865);
xor U5940 (N_5940,N_5899,N_5879);
and U5941 (N_5941,N_5811,N_5857);
or U5942 (N_5942,N_5824,N_5884);
nand U5943 (N_5943,N_5802,N_5892);
xnor U5944 (N_5944,N_5873,N_5861);
and U5945 (N_5945,N_5897,N_5833);
or U5946 (N_5946,N_5819,N_5807);
or U5947 (N_5947,N_5871,N_5822);
nand U5948 (N_5948,N_5866,N_5843);
nor U5949 (N_5949,N_5854,N_5851);
or U5950 (N_5950,N_5837,N_5897);
xnor U5951 (N_5951,N_5834,N_5826);
xor U5952 (N_5952,N_5895,N_5875);
and U5953 (N_5953,N_5874,N_5855);
xor U5954 (N_5954,N_5813,N_5825);
or U5955 (N_5955,N_5804,N_5819);
and U5956 (N_5956,N_5878,N_5855);
xnor U5957 (N_5957,N_5846,N_5871);
nand U5958 (N_5958,N_5804,N_5837);
and U5959 (N_5959,N_5865,N_5804);
xor U5960 (N_5960,N_5863,N_5892);
xnor U5961 (N_5961,N_5880,N_5865);
or U5962 (N_5962,N_5861,N_5851);
xnor U5963 (N_5963,N_5869,N_5873);
xnor U5964 (N_5964,N_5891,N_5862);
nor U5965 (N_5965,N_5864,N_5811);
nand U5966 (N_5966,N_5864,N_5840);
and U5967 (N_5967,N_5890,N_5824);
or U5968 (N_5968,N_5842,N_5859);
nor U5969 (N_5969,N_5847,N_5897);
nand U5970 (N_5970,N_5888,N_5841);
nor U5971 (N_5971,N_5846,N_5810);
nand U5972 (N_5972,N_5889,N_5801);
and U5973 (N_5973,N_5820,N_5805);
nor U5974 (N_5974,N_5811,N_5892);
nor U5975 (N_5975,N_5857,N_5831);
xor U5976 (N_5976,N_5807,N_5800);
xnor U5977 (N_5977,N_5859,N_5834);
xnor U5978 (N_5978,N_5899,N_5817);
xor U5979 (N_5979,N_5858,N_5854);
nand U5980 (N_5980,N_5868,N_5879);
xor U5981 (N_5981,N_5882,N_5842);
and U5982 (N_5982,N_5877,N_5862);
or U5983 (N_5983,N_5841,N_5858);
nand U5984 (N_5984,N_5840,N_5810);
xor U5985 (N_5985,N_5831,N_5806);
xnor U5986 (N_5986,N_5895,N_5866);
nand U5987 (N_5987,N_5810,N_5868);
and U5988 (N_5988,N_5898,N_5829);
xnor U5989 (N_5989,N_5870,N_5885);
nand U5990 (N_5990,N_5855,N_5815);
nand U5991 (N_5991,N_5843,N_5857);
nor U5992 (N_5992,N_5821,N_5845);
and U5993 (N_5993,N_5865,N_5810);
and U5994 (N_5994,N_5867,N_5813);
nand U5995 (N_5995,N_5847,N_5896);
and U5996 (N_5996,N_5833,N_5808);
nand U5997 (N_5997,N_5894,N_5895);
or U5998 (N_5998,N_5857,N_5859);
and U5999 (N_5999,N_5821,N_5835);
or U6000 (N_6000,N_5944,N_5999);
nor U6001 (N_6001,N_5925,N_5998);
and U6002 (N_6002,N_5911,N_5910);
nor U6003 (N_6003,N_5954,N_5937);
or U6004 (N_6004,N_5950,N_5966);
nand U6005 (N_6005,N_5956,N_5986);
or U6006 (N_6006,N_5917,N_5949);
xor U6007 (N_6007,N_5970,N_5931);
nor U6008 (N_6008,N_5982,N_5947);
or U6009 (N_6009,N_5934,N_5920);
and U6010 (N_6010,N_5997,N_5918);
nand U6011 (N_6011,N_5984,N_5940);
nor U6012 (N_6012,N_5973,N_5935);
and U6013 (N_6013,N_5968,N_5967);
nand U6014 (N_6014,N_5916,N_5914);
xor U6015 (N_6015,N_5957,N_5938);
nor U6016 (N_6016,N_5933,N_5905);
nand U6017 (N_6017,N_5928,N_5969);
and U6018 (N_6018,N_5955,N_5921);
xor U6019 (N_6019,N_5962,N_5902);
and U6020 (N_6020,N_5953,N_5923);
xor U6021 (N_6021,N_5965,N_5961);
xor U6022 (N_6022,N_5988,N_5939);
nand U6023 (N_6023,N_5919,N_5912);
or U6024 (N_6024,N_5908,N_5951);
xnor U6025 (N_6025,N_5959,N_5994);
and U6026 (N_6026,N_5991,N_5929);
or U6027 (N_6027,N_5915,N_5909);
or U6028 (N_6028,N_5936,N_5977);
or U6029 (N_6029,N_5989,N_5941);
or U6030 (N_6030,N_5903,N_5926);
nand U6031 (N_6031,N_5992,N_5907);
or U6032 (N_6032,N_5942,N_5996);
and U6033 (N_6033,N_5971,N_5943);
and U6034 (N_6034,N_5904,N_5980);
xnor U6035 (N_6035,N_5985,N_5976);
xor U6036 (N_6036,N_5995,N_5974);
xor U6037 (N_6037,N_5958,N_5930);
and U6038 (N_6038,N_5946,N_5963);
xnor U6039 (N_6039,N_5948,N_5927);
or U6040 (N_6040,N_5960,N_5932);
xnor U6041 (N_6041,N_5983,N_5990);
nand U6042 (N_6042,N_5964,N_5952);
xnor U6043 (N_6043,N_5906,N_5978);
or U6044 (N_6044,N_5922,N_5924);
nand U6045 (N_6045,N_5913,N_5972);
xor U6046 (N_6046,N_5975,N_5987);
or U6047 (N_6047,N_5981,N_5979);
xnor U6048 (N_6048,N_5901,N_5945);
nand U6049 (N_6049,N_5993,N_5900);
nand U6050 (N_6050,N_5966,N_5939);
nor U6051 (N_6051,N_5938,N_5933);
nand U6052 (N_6052,N_5998,N_5966);
and U6053 (N_6053,N_5975,N_5946);
and U6054 (N_6054,N_5915,N_5914);
or U6055 (N_6055,N_5968,N_5935);
or U6056 (N_6056,N_5992,N_5972);
or U6057 (N_6057,N_5950,N_5925);
and U6058 (N_6058,N_5951,N_5996);
nand U6059 (N_6059,N_5981,N_5936);
nor U6060 (N_6060,N_5970,N_5937);
nor U6061 (N_6061,N_5962,N_5982);
xor U6062 (N_6062,N_5941,N_5966);
or U6063 (N_6063,N_5919,N_5928);
xor U6064 (N_6064,N_5983,N_5909);
or U6065 (N_6065,N_5949,N_5923);
nor U6066 (N_6066,N_5918,N_5916);
xnor U6067 (N_6067,N_5924,N_5903);
nand U6068 (N_6068,N_5931,N_5926);
nand U6069 (N_6069,N_5959,N_5938);
and U6070 (N_6070,N_5900,N_5962);
or U6071 (N_6071,N_5910,N_5990);
and U6072 (N_6072,N_5986,N_5999);
nor U6073 (N_6073,N_5975,N_5993);
and U6074 (N_6074,N_5923,N_5978);
and U6075 (N_6075,N_5909,N_5997);
nand U6076 (N_6076,N_5953,N_5927);
nand U6077 (N_6077,N_5991,N_5925);
xor U6078 (N_6078,N_5966,N_5977);
xor U6079 (N_6079,N_5988,N_5913);
xor U6080 (N_6080,N_5985,N_5935);
nor U6081 (N_6081,N_5924,N_5968);
nor U6082 (N_6082,N_5947,N_5905);
or U6083 (N_6083,N_5942,N_5979);
and U6084 (N_6084,N_5982,N_5905);
xnor U6085 (N_6085,N_5942,N_5986);
nand U6086 (N_6086,N_5974,N_5911);
xor U6087 (N_6087,N_5963,N_5970);
or U6088 (N_6088,N_5957,N_5968);
or U6089 (N_6089,N_5950,N_5916);
or U6090 (N_6090,N_5922,N_5920);
or U6091 (N_6091,N_5973,N_5979);
xnor U6092 (N_6092,N_5937,N_5959);
or U6093 (N_6093,N_5984,N_5935);
xnor U6094 (N_6094,N_5937,N_5938);
nor U6095 (N_6095,N_5954,N_5922);
or U6096 (N_6096,N_5965,N_5908);
or U6097 (N_6097,N_5940,N_5927);
and U6098 (N_6098,N_5923,N_5921);
xor U6099 (N_6099,N_5965,N_5956);
nand U6100 (N_6100,N_6053,N_6079);
nor U6101 (N_6101,N_6008,N_6036);
xnor U6102 (N_6102,N_6063,N_6033);
xnor U6103 (N_6103,N_6074,N_6092);
and U6104 (N_6104,N_6059,N_6041);
xor U6105 (N_6105,N_6093,N_6001);
nand U6106 (N_6106,N_6046,N_6034);
and U6107 (N_6107,N_6009,N_6006);
nor U6108 (N_6108,N_6018,N_6027);
and U6109 (N_6109,N_6091,N_6057);
nand U6110 (N_6110,N_6032,N_6013);
or U6111 (N_6111,N_6024,N_6003);
xor U6112 (N_6112,N_6068,N_6081);
nor U6113 (N_6113,N_6031,N_6066);
xnor U6114 (N_6114,N_6049,N_6060);
or U6115 (N_6115,N_6095,N_6025);
and U6116 (N_6116,N_6012,N_6082);
or U6117 (N_6117,N_6071,N_6010);
and U6118 (N_6118,N_6039,N_6050);
and U6119 (N_6119,N_6097,N_6083);
or U6120 (N_6120,N_6069,N_6077);
or U6121 (N_6121,N_6043,N_6085);
xor U6122 (N_6122,N_6017,N_6087);
nand U6123 (N_6123,N_6099,N_6056);
or U6124 (N_6124,N_6045,N_6086);
nor U6125 (N_6125,N_6048,N_6040);
and U6126 (N_6126,N_6002,N_6023);
or U6127 (N_6127,N_6028,N_6042);
nand U6128 (N_6128,N_6065,N_6052);
nor U6129 (N_6129,N_6073,N_6089);
xnor U6130 (N_6130,N_6070,N_6038);
nand U6131 (N_6131,N_6088,N_6047);
or U6132 (N_6132,N_6007,N_6072);
xor U6133 (N_6133,N_6000,N_6011);
nor U6134 (N_6134,N_6076,N_6005);
xnor U6135 (N_6135,N_6096,N_6015);
nand U6136 (N_6136,N_6062,N_6030);
nand U6137 (N_6137,N_6098,N_6020);
xor U6138 (N_6138,N_6084,N_6094);
or U6139 (N_6139,N_6058,N_6080);
nand U6140 (N_6140,N_6019,N_6067);
nor U6141 (N_6141,N_6044,N_6064);
nand U6142 (N_6142,N_6075,N_6051);
nand U6143 (N_6143,N_6021,N_6022);
nand U6144 (N_6144,N_6016,N_6014);
or U6145 (N_6145,N_6035,N_6029);
xnor U6146 (N_6146,N_6037,N_6078);
nor U6147 (N_6147,N_6061,N_6026);
and U6148 (N_6148,N_6054,N_6055);
nand U6149 (N_6149,N_6090,N_6004);
nor U6150 (N_6150,N_6048,N_6095);
or U6151 (N_6151,N_6075,N_6020);
xnor U6152 (N_6152,N_6066,N_6099);
and U6153 (N_6153,N_6034,N_6050);
nand U6154 (N_6154,N_6005,N_6018);
or U6155 (N_6155,N_6057,N_6060);
xor U6156 (N_6156,N_6021,N_6086);
xor U6157 (N_6157,N_6078,N_6054);
nand U6158 (N_6158,N_6077,N_6088);
xnor U6159 (N_6159,N_6070,N_6043);
xnor U6160 (N_6160,N_6092,N_6080);
xor U6161 (N_6161,N_6084,N_6070);
nand U6162 (N_6162,N_6045,N_6017);
xnor U6163 (N_6163,N_6057,N_6014);
nor U6164 (N_6164,N_6059,N_6005);
nor U6165 (N_6165,N_6063,N_6091);
xor U6166 (N_6166,N_6004,N_6098);
xor U6167 (N_6167,N_6071,N_6000);
or U6168 (N_6168,N_6075,N_6030);
nor U6169 (N_6169,N_6071,N_6093);
and U6170 (N_6170,N_6012,N_6070);
nand U6171 (N_6171,N_6009,N_6098);
nor U6172 (N_6172,N_6086,N_6083);
and U6173 (N_6173,N_6018,N_6015);
nor U6174 (N_6174,N_6040,N_6078);
or U6175 (N_6175,N_6073,N_6096);
or U6176 (N_6176,N_6004,N_6006);
and U6177 (N_6177,N_6050,N_6018);
nand U6178 (N_6178,N_6016,N_6090);
nor U6179 (N_6179,N_6044,N_6004);
and U6180 (N_6180,N_6048,N_6006);
and U6181 (N_6181,N_6080,N_6089);
and U6182 (N_6182,N_6050,N_6082);
xnor U6183 (N_6183,N_6059,N_6019);
and U6184 (N_6184,N_6031,N_6041);
nand U6185 (N_6185,N_6051,N_6049);
and U6186 (N_6186,N_6047,N_6037);
and U6187 (N_6187,N_6003,N_6055);
or U6188 (N_6188,N_6062,N_6020);
nand U6189 (N_6189,N_6035,N_6016);
nand U6190 (N_6190,N_6084,N_6092);
nand U6191 (N_6191,N_6006,N_6076);
nand U6192 (N_6192,N_6065,N_6037);
or U6193 (N_6193,N_6008,N_6090);
and U6194 (N_6194,N_6007,N_6020);
nand U6195 (N_6195,N_6099,N_6036);
nand U6196 (N_6196,N_6051,N_6002);
xnor U6197 (N_6197,N_6051,N_6091);
nand U6198 (N_6198,N_6003,N_6050);
and U6199 (N_6199,N_6074,N_6008);
or U6200 (N_6200,N_6130,N_6124);
nand U6201 (N_6201,N_6143,N_6168);
xor U6202 (N_6202,N_6183,N_6157);
or U6203 (N_6203,N_6131,N_6159);
nor U6204 (N_6204,N_6151,N_6165);
and U6205 (N_6205,N_6198,N_6113);
xnor U6206 (N_6206,N_6188,N_6136);
or U6207 (N_6207,N_6181,N_6109);
nor U6208 (N_6208,N_6197,N_6179);
nand U6209 (N_6209,N_6135,N_6175);
nand U6210 (N_6210,N_6133,N_6166);
nor U6211 (N_6211,N_6108,N_6184);
nor U6212 (N_6212,N_6123,N_6173);
xor U6213 (N_6213,N_6101,N_6112);
xor U6214 (N_6214,N_6120,N_6107);
and U6215 (N_6215,N_6164,N_6150);
and U6216 (N_6216,N_6161,N_6119);
and U6217 (N_6217,N_6155,N_6189);
xnor U6218 (N_6218,N_6193,N_6138);
and U6219 (N_6219,N_6180,N_6187);
xor U6220 (N_6220,N_6167,N_6154);
nand U6221 (N_6221,N_6185,N_6176);
nand U6222 (N_6222,N_6139,N_6192);
nand U6223 (N_6223,N_6127,N_6115);
and U6224 (N_6224,N_6141,N_6178);
and U6225 (N_6225,N_6140,N_6114);
nor U6226 (N_6226,N_6177,N_6195);
nand U6227 (N_6227,N_6100,N_6102);
or U6228 (N_6228,N_6134,N_6172);
or U6229 (N_6229,N_6149,N_6170);
or U6230 (N_6230,N_6162,N_6194);
nor U6231 (N_6231,N_6129,N_6116);
nand U6232 (N_6232,N_6182,N_6186);
nor U6233 (N_6233,N_6153,N_6147);
or U6234 (N_6234,N_6110,N_6117);
nor U6235 (N_6235,N_6171,N_6174);
nand U6236 (N_6236,N_6144,N_6191);
nor U6237 (N_6237,N_6132,N_6169);
nor U6238 (N_6238,N_6152,N_6158);
xor U6239 (N_6239,N_6111,N_6105);
nand U6240 (N_6240,N_6125,N_6142);
nor U6241 (N_6241,N_6156,N_6137);
xor U6242 (N_6242,N_6104,N_6160);
or U6243 (N_6243,N_6121,N_6190);
and U6244 (N_6244,N_6126,N_6163);
xnor U6245 (N_6245,N_6122,N_6148);
or U6246 (N_6246,N_6199,N_6103);
nor U6247 (N_6247,N_6128,N_6118);
or U6248 (N_6248,N_6146,N_6196);
and U6249 (N_6249,N_6145,N_6106);
xnor U6250 (N_6250,N_6197,N_6142);
or U6251 (N_6251,N_6161,N_6153);
or U6252 (N_6252,N_6186,N_6101);
nor U6253 (N_6253,N_6111,N_6120);
or U6254 (N_6254,N_6118,N_6135);
and U6255 (N_6255,N_6188,N_6122);
xor U6256 (N_6256,N_6163,N_6174);
and U6257 (N_6257,N_6161,N_6122);
and U6258 (N_6258,N_6191,N_6116);
and U6259 (N_6259,N_6193,N_6126);
or U6260 (N_6260,N_6180,N_6135);
or U6261 (N_6261,N_6132,N_6125);
xor U6262 (N_6262,N_6160,N_6113);
xor U6263 (N_6263,N_6197,N_6187);
and U6264 (N_6264,N_6150,N_6195);
xor U6265 (N_6265,N_6196,N_6114);
or U6266 (N_6266,N_6188,N_6148);
or U6267 (N_6267,N_6171,N_6140);
or U6268 (N_6268,N_6146,N_6153);
or U6269 (N_6269,N_6170,N_6156);
nand U6270 (N_6270,N_6180,N_6131);
or U6271 (N_6271,N_6110,N_6181);
xnor U6272 (N_6272,N_6196,N_6123);
xnor U6273 (N_6273,N_6101,N_6169);
nor U6274 (N_6274,N_6158,N_6159);
or U6275 (N_6275,N_6185,N_6145);
or U6276 (N_6276,N_6157,N_6178);
nor U6277 (N_6277,N_6116,N_6110);
or U6278 (N_6278,N_6132,N_6129);
xnor U6279 (N_6279,N_6132,N_6126);
nor U6280 (N_6280,N_6147,N_6196);
xor U6281 (N_6281,N_6102,N_6137);
xnor U6282 (N_6282,N_6184,N_6149);
nand U6283 (N_6283,N_6145,N_6143);
nand U6284 (N_6284,N_6121,N_6111);
and U6285 (N_6285,N_6152,N_6124);
xor U6286 (N_6286,N_6165,N_6174);
nor U6287 (N_6287,N_6165,N_6121);
xnor U6288 (N_6288,N_6135,N_6121);
and U6289 (N_6289,N_6168,N_6188);
xor U6290 (N_6290,N_6184,N_6130);
and U6291 (N_6291,N_6182,N_6198);
nand U6292 (N_6292,N_6137,N_6157);
or U6293 (N_6293,N_6142,N_6169);
or U6294 (N_6294,N_6171,N_6186);
nor U6295 (N_6295,N_6157,N_6193);
and U6296 (N_6296,N_6130,N_6185);
nor U6297 (N_6297,N_6137,N_6190);
and U6298 (N_6298,N_6141,N_6114);
nor U6299 (N_6299,N_6124,N_6107);
xor U6300 (N_6300,N_6269,N_6299);
or U6301 (N_6301,N_6205,N_6277);
and U6302 (N_6302,N_6294,N_6268);
nand U6303 (N_6303,N_6263,N_6260);
or U6304 (N_6304,N_6286,N_6261);
and U6305 (N_6305,N_6221,N_6288);
and U6306 (N_6306,N_6287,N_6264);
and U6307 (N_6307,N_6280,N_6236);
nor U6308 (N_6308,N_6275,N_6231);
xnor U6309 (N_6309,N_6239,N_6214);
nand U6310 (N_6310,N_6291,N_6265);
xor U6311 (N_6311,N_6241,N_6203);
nand U6312 (N_6312,N_6272,N_6242);
and U6313 (N_6313,N_6215,N_6250);
or U6314 (N_6314,N_6212,N_6200);
and U6315 (N_6315,N_6222,N_6283);
xnor U6316 (N_6316,N_6237,N_6229);
or U6317 (N_6317,N_6225,N_6248);
xnor U6318 (N_6318,N_6249,N_6274);
or U6319 (N_6319,N_6211,N_6298);
and U6320 (N_6320,N_6273,N_6233);
and U6321 (N_6321,N_6276,N_6297);
nand U6322 (N_6322,N_6246,N_6234);
or U6323 (N_6323,N_6257,N_6208);
nor U6324 (N_6324,N_6207,N_6278);
and U6325 (N_6325,N_6279,N_6293);
nor U6326 (N_6326,N_6271,N_6245);
nor U6327 (N_6327,N_6251,N_6282);
nand U6328 (N_6328,N_6267,N_6210);
xnor U6329 (N_6329,N_6284,N_6219);
nor U6330 (N_6330,N_6226,N_6266);
xnor U6331 (N_6331,N_6204,N_6254);
nor U6332 (N_6332,N_6289,N_6258);
nor U6333 (N_6333,N_6228,N_6220);
nor U6334 (N_6334,N_6255,N_6270);
nand U6335 (N_6335,N_6230,N_6259);
or U6336 (N_6336,N_6216,N_6296);
or U6337 (N_6337,N_6252,N_6238);
and U6338 (N_6338,N_6256,N_6253);
nand U6339 (N_6339,N_6290,N_6281);
and U6340 (N_6340,N_6244,N_6227);
nand U6341 (N_6341,N_6240,N_6202);
and U6342 (N_6342,N_6206,N_6235);
xor U6343 (N_6343,N_6243,N_6223);
xnor U6344 (N_6344,N_6285,N_6209);
nor U6345 (N_6345,N_6292,N_6247);
xnor U6346 (N_6346,N_6201,N_6295);
nor U6347 (N_6347,N_6218,N_6224);
nand U6348 (N_6348,N_6217,N_6213);
or U6349 (N_6349,N_6262,N_6232);
xnor U6350 (N_6350,N_6237,N_6277);
nand U6351 (N_6351,N_6242,N_6280);
nor U6352 (N_6352,N_6201,N_6293);
xor U6353 (N_6353,N_6260,N_6257);
or U6354 (N_6354,N_6246,N_6211);
xor U6355 (N_6355,N_6276,N_6263);
and U6356 (N_6356,N_6289,N_6226);
nor U6357 (N_6357,N_6290,N_6248);
nand U6358 (N_6358,N_6210,N_6278);
or U6359 (N_6359,N_6297,N_6241);
xnor U6360 (N_6360,N_6200,N_6225);
nor U6361 (N_6361,N_6247,N_6254);
xor U6362 (N_6362,N_6246,N_6278);
or U6363 (N_6363,N_6240,N_6282);
nor U6364 (N_6364,N_6276,N_6288);
nor U6365 (N_6365,N_6223,N_6287);
nor U6366 (N_6366,N_6246,N_6251);
xor U6367 (N_6367,N_6227,N_6249);
or U6368 (N_6368,N_6291,N_6276);
nand U6369 (N_6369,N_6270,N_6237);
xor U6370 (N_6370,N_6276,N_6277);
or U6371 (N_6371,N_6293,N_6266);
xnor U6372 (N_6372,N_6252,N_6242);
and U6373 (N_6373,N_6292,N_6289);
and U6374 (N_6374,N_6234,N_6272);
nor U6375 (N_6375,N_6297,N_6245);
or U6376 (N_6376,N_6258,N_6230);
or U6377 (N_6377,N_6232,N_6282);
xnor U6378 (N_6378,N_6247,N_6207);
xnor U6379 (N_6379,N_6235,N_6283);
nor U6380 (N_6380,N_6224,N_6292);
xnor U6381 (N_6381,N_6221,N_6261);
nor U6382 (N_6382,N_6219,N_6241);
or U6383 (N_6383,N_6256,N_6238);
or U6384 (N_6384,N_6273,N_6256);
or U6385 (N_6385,N_6249,N_6218);
nor U6386 (N_6386,N_6229,N_6278);
nand U6387 (N_6387,N_6208,N_6279);
and U6388 (N_6388,N_6216,N_6266);
xor U6389 (N_6389,N_6255,N_6232);
xor U6390 (N_6390,N_6250,N_6238);
or U6391 (N_6391,N_6288,N_6220);
nor U6392 (N_6392,N_6271,N_6229);
xnor U6393 (N_6393,N_6208,N_6274);
nor U6394 (N_6394,N_6243,N_6206);
xor U6395 (N_6395,N_6284,N_6242);
or U6396 (N_6396,N_6249,N_6230);
xor U6397 (N_6397,N_6201,N_6262);
and U6398 (N_6398,N_6278,N_6208);
or U6399 (N_6399,N_6281,N_6286);
and U6400 (N_6400,N_6383,N_6357);
and U6401 (N_6401,N_6342,N_6372);
and U6402 (N_6402,N_6325,N_6390);
nand U6403 (N_6403,N_6341,N_6380);
or U6404 (N_6404,N_6387,N_6334);
nand U6405 (N_6405,N_6310,N_6358);
xor U6406 (N_6406,N_6305,N_6324);
nand U6407 (N_6407,N_6355,N_6371);
nand U6408 (N_6408,N_6388,N_6395);
and U6409 (N_6409,N_6301,N_6336);
nor U6410 (N_6410,N_6317,N_6314);
nand U6411 (N_6411,N_6396,N_6338);
nor U6412 (N_6412,N_6359,N_6354);
nand U6413 (N_6413,N_6381,N_6377);
or U6414 (N_6414,N_6329,N_6389);
and U6415 (N_6415,N_6374,N_6308);
and U6416 (N_6416,N_6348,N_6315);
and U6417 (N_6417,N_6313,N_6347);
nor U6418 (N_6418,N_6356,N_6382);
or U6419 (N_6419,N_6302,N_6367);
xor U6420 (N_6420,N_6343,N_6340);
nand U6421 (N_6421,N_6370,N_6397);
xor U6422 (N_6422,N_6327,N_6304);
or U6423 (N_6423,N_6332,N_6392);
xor U6424 (N_6424,N_6376,N_6352);
nor U6425 (N_6425,N_6379,N_6399);
xor U6426 (N_6426,N_6300,N_6316);
or U6427 (N_6427,N_6333,N_6394);
nor U6428 (N_6428,N_6386,N_6319);
nand U6429 (N_6429,N_6346,N_6368);
nor U6430 (N_6430,N_6361,N_6309);
nor U6431 (N_6431,N_6323,N_6378);
nand U6432 (N_6432,N_6366,N_6303);
nand U6433 (N_6433,N_6373,N_6339);
or U6434 (N_6434,N_6328,N_6335);
xor U6435 (N_6435,N_6385,N_6345);
nand U6436 (N_6436,N_6330,N_6311);
or U6437 (N_6437,N_6365,N_6318);
nand U6438 (N_6438,N_6363,N_6398);
nand U6439 (N_6439,N_6320,N_6369);
nor U6440 (N_6440,N_6393,N_6331);
and U6441 (N_6441,N_6326,N_6306);
nor U6442 (N_6442,N_6349,N_6344);
or U6443 (N_6443,N_6375,N_6362);
and U6444 (N_6444,N_6312,N_6350);
or U6445 (N_6445,N_6321,N_6351);
and U6446 (N_6446,N_6391,N_6307);
nor U6447 (N_6447,N_6364,N_6337);
and U6448 (N_6448,N_6360,N_6322);
xnor U6449 (N_6449,N_6353,N_6384);
or U6450 (N_6450,N_6323,N_6362);
nand U6451 (N_6451,N_6398,N_6396);
or U6452 (N_6452,N_6325,N_6315);
nor U6453 (N_6453,N_6384,N_6323);
xor U6454 (N_6454,N_6312,N_6331);
and U6455 (N_6455,N_6307,N_6358);
nand U6456 (N_6456,N_6363,N_6360);
nor U6457 (N_6457,N_6367,N_6306);
xnor U6458 (N_6458,N_6345,N_6359);
nand U6459 (N_6459,N_6346,N_6359);
or U6460 (N_6460,N_6308,N_6332);
nand U6461 (N_6461,N_6339,N_6351);
or U6462 (N_6462,N_6305,N_6386);
and U6463 (N_6463,N_6325,N_6341);
nor U6464 (N_6464,N_6312,N_6363);
and U6465 (N_6465,N_6374,N_6348);
and U6466 (N_6466,N_6374,N_6310);
nand U6467 (N_6467,N_6307,N_6352);
nand U6468 (N_6468,N_6344,N_6328);
and U6469 (N_6469,N_6395,N_6386);
nand U6470 (N_6470,N_6358,N_6317);
nand U6471 (N_6471,N_6315,N_6308);
and U6472 (N_6472,N_6305,N_6375);
or U6473 (N_6473,N_6355,N_6377);
or U6474 (N_6474,N_6365,N_6313);
xnor U6475 (N_6475,N_6375,N_6336);
nand U6476 (N_6476,N_6399,N_6350);
or U6477 (N_6477,N_6395,N_6380);
xor U6478 (N_6478,N_6336,N_6378);
nand U6479 (N_6479,N_6320,N_6343);
nand U6480 (N_6480,N_6346,N_6305);
and U6481 (N_6481,N_6371,N_6351);
nand U6482 (N_6482,N_6388,N_6396);
nand U6483 (N_6483,N_6306,N_6342);
xor U6484 (N_6484,N_6387,N_6311);
and U6485 (N_6485,N_6305,N_6358);
nor U6486 (N_6486,N_6312,N_6357);
nand U6487 (N_6487,N_6322,N_6359);
nand U6488 (N_6488,N_6375,N_6330);
and U6489 (N_6489,N_6345,N_6322);
nand U6490 (N_6490,N_6336,N_6314);
or U6491 (N_6491,N_6399,N_6342);
and U6492 (N_6492,N_6336,N_6322);
nand U6493 (N_6493,N_6368,N_6314);
xor U6494 (N_6494,N_6305,N_6314);
xnor U6495 (N_6495,N_6398,N_6359);
xor U6496 (N_6496,N_6392,N_6371);
nand U6497 (N_6497,N_6371,N_6334);
nand U6498 (N_6498,N_6373,N_6310);
and U6499 (N_6499,N_6365,N_6320);
nand U6500 (N_6500,N_6413,N_6429);
or U6501 (N_6501,N_6433,N_6454);
nand U6502 (N_6502,N_6445,N_6421);
and U6503 (N_6503,N_6439,N_6485);
nor U6504 (N_6504,N_6481,N_6463);
or U6505 (N_6505,N_6480,N_6446);
nor U6506 (N_6506,N_6473,N_6467);
and U6507 (N_6507,N_6475,N_6482);
or U6508 (N_6508,N_6428,N_6487);
xor U6509 (N_6509,N_6405,N_6432);
nand U6510 (N_6510,N_6474,N_6401);
or U6511 (N_6511,N_6497,N_6417);
xnor U6512 (N_6512,N_6465,N_6422);
and U6513 (N_6513,N_6420,N_6476);
or U6514 (N_6514,N_6409,N_6494);
and U6515 (N_6515,N_6489,N_6495);
and U6516 (N_6516,N_6450,N_6410);
nand U6517 (N_6517,N_6464,N_6424);
xnor U6518 (N_6518,N_6466,N_6498);
nand U6519 (N_6519,N_6478,N_6451);
and U6520 (N_6520,N_6431,N_6444);
xor U6521 (N_6521,N_6449,N_6436);
or U6522 (N_6522,N_6496,N_6403);
xnor U6523 (N_6523,N_6414,N_6479);
xor U6524 (N_6524,N_6423,N_6408);
nand U6525 (N_6525,N_6483,N_6492);
nor U6526 (N_6526,N_6459,N_6460);
nor U6527 (N_6527,N_6400,N_6461);
or U6528 (N_6528,N_6455,N_6402);
nor U6529 (N_6529,N_6484,N_6430);
or U6530 (N_6530,N_6457,N_6448);
nor U6531 (N_6531,N_6419,N_6404);
and U6532 (N_6532,N_6440,N_6438);
nand U6533 (N_6533,N_6426,N_6488);
nand U6534 (N_6534,N_6499,N_6418);
nor U6535 (N_6535,N_6458,N_6462);
nor U6536 (N_6536,N_6441,N_6407);
and U6537 (N_6537,N_6456,N_6411);
xor U6538 (N_6538,N_6415,N_6472);
nand U6539 (N_6539,N_6412,N_6471);
nand U6540 (N_6540,N_6452,N_6435);
xnor U6541 (N_6541,N_6425,N_6443);
and U6542 (N_6542,N_6470,N_6416);
nand U6543 (N_6543,N_6442,N_6491);
or U6544 (N_6544,N_6437,N_6477);
and U6545 (N_6545,N_6406,N_6490);
and U6546 (N_6546,N_6427,N_6434);
nand U6547 (N_6547,N_6468,N_6469);
and U6548 (N_6548,N_6447,N_6493);
nor U6549 (N_6549,N_6486,N_6453);
xor U6550 (N_6550,N_6493,N_6491);
xnor U6551 (N_6551,N_6484,N_6494);
xnor U6552 (N_6552,N_6445,N_6406);
nor U6553 (N_6553,N_6478,N_6436);
nor U6554 (N_6554,N_6422,N_6431);
nor U6555 (N_6555,N_6456,N_6472);
nand U6556 (N_6556,N_6436,N_6467);
and U6557 (N_6557,N_6407,N_6422);
or U6558 (N_6558,N_6447,N_6414);
or U6559 (N_6559,N_6494,N_6455);
nand U6560 (N_6560,N_6476,N_6439);
nand U6561 (N_6561,N_6494,N_6421);
or U6562 (N_6562,N_6432,N_6487);
xnor U6563 (N_6563,N_6464,N_6462);
nor U6564 (N_6564,N_6475,N_6431);
nor U6565 (N_6565,N_6425,N_6414);
and U6566 (N_6566,N_6415,N_6420);
nor U6567 (N_6567,N_6460,N_6454);
or U6568 (N_6568,N_6475,N_6478);
nand U6569 (N_6569,N_6412,N_6452);
or U6570 (N_6570,N_6428,N_6425);
xnor U6571 (N_6571,N_6426,N_6499);
nand U6572 (N_6572,N_6451,N_6414);
nor U6573 (N_6573,N_6492,N_6479);
xor U6574 (N_6574,N_6449,N_6489);
nor U6575 (N_6575,N_6456,N_6475);
or U6576 (N_6576,N_6421,N_6430);
or U6577 (N_6577,N_6499,N_6492);
nand U6578 (N_6578,N_6483,N_6430);
and U6579 (N_6579,N_6425,N_6432);
nand U6580 (N_6580,N_6422,N_6437);
nand U6581 (N_6581,N_6497,N_6440);
and U6582 (N_6582,N_6460,N_6474);
nand U6583 (N_6583,N_6451,N_6429);
nor U6584 (N_6584,N_6451,N_6448);
nand U6585 (N_6585,N_6422,N_6490);
and U6586 (N_6586,N_6425,N_6486);
xnor U6587 (N_6587,N_6451,N_6485);
and U6588 (N_6588,N_6411,N_6477);
xnor U6589 (N_6589,N_6429,N_6495);
nand U6590 (N_6590,N_6454,N_6446);
nand U6591 (N_6591,N_6412,N_6456);
or U6592 (N_6592,N_6467,N_6453);
and U6593 (N_6593,N_6470,N_6418);
and U6594 (N_6594,N_6444,N_6484);
or U6595 (N_6595,N_6483,N_6476);
or U6596 (N_6596,N_6474,N_6455);
nor U6597 (N_6597,N_6424,N_6471);
nand U6598 (N_6598,N_6412,N_6437);
nand U6599 (N_6599,N_6491,N_6492);
or U6600 (N_6600,N_6594,N_6531);
or U6601 (N_6601,N_6507,N_6590);
nor U6602 (N_6602,N_6540,N_6517);
nand U6603 (N_6603,N_6514,N_6599);
nor U6604 (N_6604,N_6521,N_6587);
or U6605 (N_6605,N_6560,N_6589);
xnor U6606 (N_6606,N_6503,N_6538);
xnor U6607 (N_6607,N_6552,N_6523);
or U6608 (N_6608,N_6570,N_6545);
xor U6609 (N_6609,N_6592,N_6509);
xor U6610 (N_6610,N_6564,N_6568);
or U6611 (N_6611,N_6567,N_6586);
and U6612 (N_6612,N_6544,N_6534);
nand U6613 (N_6613,N_6510,N_6578);
and U6614 (N_6614,N_6550,N_6546);
nor U6615 (N_6615,N_6504,N_6561);
or U6616 (N_6616,N_6576,N_6520);
and U6617 (N_6617,N_6582,N_6522);
and U6618 (N_6618,N_6557,N_6584);
xnor U6619 (N_6619,N_6555,N_6597);
nand U6620 (N_6620,N_6566,N_6593);
nor U6621 (N_6621,N_6542,N_6549);
or U6622 (N_6622,N_6580,N_6554);
nand U6623 (N_6623,N_6506,N_6572);
or U6624 (N_6624,N_6595,N_6562);
and U6625 (N_6625,N_6537,N_6532);
or U6626 (N_6626,N_6543,N_6530);
or U6627 (N_6627,N_6548,N_6518);
and U6628 (N_6628,N_6525,N_6565);
and U6629 (N_6629,N_6571,N_6574);
nand U6630 (N_6630,N_6556,N_6547);
xor U6631 (N_6631,N_6512,N_6598);
nor U6632 (N_6632,N_6511,N_6533);
and U6633 (N_6633,N_6501,N_6539);
nor U6634 (N_6634,N_6558,N_6527);
nand U6635 (N_6635,N_6502,N_6516);
or U6636 (N_6636,N_6596,N_6519);
or U6637 (N_6637,N_6563,N_6575);
xnor U6638 (N_6638,N_6505,N_6513);
xnor U6639 (N_6639,N_6588,N_6529);
xnor U6640 (N_6640,N_6500,N_6508);
nor U6641 (N_6641,N_6579,N_6528);
nand U6642 (N_6642,N_6551,N_6581);
nand U6643 (N_6643,N_6524,N_6585);
xnor U6644 (N_6644,N_6583,N_6526);
xnor U6645 (N_6645,N_6591,N_6569);
or U6646 (N_6646,N_6553,N_6536);
nand U6647 (N_6647,N_6559,N_6573);
or U6648 (N_6648,N_6535,N_6577);
nor U6649 (N_6649,N_6541,N_6515);
and U6650 (N_6650,N_6591,N_6510);
or U6651 (N_6651,N_6577,N_6530);
and U6652 (N_6652,N_6548,N_6563);
or U6653 (N_6653,N_6524,N_6586);
nand U6654 (N_6654,N_6532,N_6507);
and U6655 (N_6655,N_6555,N_6541);
or U6656 (N_6656,N_6565,N_6538);
nor U6657 (N_6657,N_6523,N_6556);
nand U6658 (N_6658,N_6595,N_6557);
nor U6659 (N_6659,N_6533,N_6539);
and U6660 (N_6660,N_6526,N_6520);
or U6661 (N_6661,N_6514,N_6571);
xor U6662 (N_6662,N_6514,N_6503);
nor U6663 (N_6663,N_6543,N_6522);
and U6664 (N_6664,N_6541,N_6563);
and U6665 (N_6665,N_6542,N_6539);
xor U6666 (N_6666,N_6511,N_6503);
or U6667 (N_6667,N_6584,N_6529);
xnor U6668 (N_6668,N_6546,N_6531);
and U6669 (N_6669,N_6514,N_6565);
xor U6670 (N_6670,N_6590,N_6562);
nor U6671 (N_6671,N_6553,N_6506);
xor U6672 (N_6672,N_6597,N_6501);
or U6673 (N_6673,N_6578,N_6538);
nand U6674 (N_6674,N_6560,N_6555);
nand U6675 (N_6675,N_6577,N_6569);
and U6676 (N_6676,N_6564,N_6597);
xnor U6677 (N_6677,N_6564,N_6512);
or U6678 (N_6678,N_6521,N_6527);
xor U6679 (N_6679,N_6517,N_6561);
or U6680 (N_6680,N_6504,N_6534);
nand U6681 (N_6681,N_6587,N_6582);
or U6682 (N_6682,N_6599,N_6521);
or U6683 (N_6683,N_6551,N_6540);
and U6684 (N_6684,N_6532,N_6513);
and U6685 (N_6685,N_6552,N_6546);
and U6686 (N_6686,N_6515,N_6570);
nand U6687 (N_6687,N_6535,N_6576);
or U6688 (N_6688,N_6560,N_6510);
and U6689 (N_6689,N_6525,N_6537);
xnor U6690 (N_6690,N_6517,N_6557);
nor U6691 (N_6691,N_6508,N_6579);
or U6692 (N_6692,N_6547,N_6510);
nor U6693 (N_6693,N_6597,N_6581);
xnor U6694 (N_6694,N_6520,N_6540);
xnor U6695 (N_6695,N_6572,N_6594);
xor U6696 (N_6696,N_6544,N_6584);
xor U6697 (N_6697,N_6592,N_6596);
xnor U6698 (N_6698,N_6567,N_6535);
xor U6699 (N_6699,N_6519,N_6540);
nand U6700 (N_6700,N_6637,N_6640);
xor U6701 (N_6701,N_6642,N_6609);
xnor U6702 (N_6702,N_6632,N_6634);
xor U6703 (N_6703,N_6679,N_6664);
xor U6704 (N_6704,N_6682,N_6680);
and U6705 (N_6705,N_6659,N_6654);
nand U6706 (N_6706,N_6620,N_6687);
and U6707 (N_6707,N_6644,N_6621);
xnor U6708 (N_6708,N_6694,N_6658);
and U6709 (N_6709,N_6618,N_6631);
nand U6710 (N_6710,N_6635,N_6651);
nand U6711 (N_6711,N_6646,N_6643);
or U6712 (N_6712,N_6653,N_6633);
nand U6713 (N_6713,N_6669,N_6602);
and U6714 (N_6714,N_6629,N_6665);
xnor U6715 (N_6715,N_6656,N_6675);
or U6716 (N_6716,N_6625,N_6668);
nand U6717 (N_6717,N_6697,N_6677);
nor U6718 (N_6718,N_6673,N_6652);
nor U6719 (N_6719,N_6648,N_6661);
xnor U6720 (N_6720,N_6696,N_6610);
nand U6721 (N_6721,N_6662,N_6671);
nor U6722 (N_6722,N_6608,N_6627);
and U6723 (N_6723,N_6636,N_6614);
nand U6724 (N_6724,N_6681,N_6623);
and U6725 (N_6725,N_6611,N_6650);
nand U6726 (N_6726,N_6691,N_6641);
nor U6727 (N_6727,N_6606,N_6600);
xnor U6728 (N_6728,N_6624,N_6683);
nand U6729 (N_6729,N_6695,N_6699);
nand U6730 (N_6730,N_6685,N_6622);
xnor U6731 (N_6731,N_6626,N_6674);
xor U6732 (N_6732,N_6647,N_6645);
nand U6733 (N_6733,N_6670,N_6684);
and U6734 (N_6734,N_6667,N_6663);
or U6735 (N_6735,N_6630,N_6660);
nor U6736 (N_6736,N_6666,N_6657);
or U6737 (N_6737,N_6616,N_6612);
nor U6738 (N_6738,N_6605,N_6686);
nor U6739 (N_6739,N_6615,N_6676);
xor U6740 (N_6740,N_6639,N_6604);
and U6741 (N_6741,N_6603,N_6638);
and U6742 (N_6742,N_6649,N_6601);
and U6743 (N_6743,N_6607,N_6672);
xnor U6744 (N_6744,N_6692,N_6613);
nand U6745 (N_6745,N_6698,N_6689);
or U6746 (N_6746,N_6688,N_6655);
and U6747 (N_6747,N_6690,N_6693);
nand U6748 (N_6748,N_6617,N_6628);
nand U6749 (N_6749,N_6678,N_6619);
nor U6750 (N_6750,N_6624,N_6670);
nor U6751 (N_6751,N_6627,N_6680);
and U6752 (N_6752,N_6612,N_6614);
or U6753 (N_6753,N_6673,N_6680);
or U6754 (N_6754,N_6649,N_6633);
or U6755 (N_6755,N_6648,N_6626);
or U6756 (N_6756,N_6666,N_6603);
xor U6757 (N_6757,N_6673,N_6625);
nor U6758 (N_6758,N_6632,N_6684);
nand U6759 (N_6759,N_6697,N_6688);
nand U6760 (N_6760,N_6662,N_6600);
nor U6761 (N_6761,N_6637,N_6634);
xor U6762 (N_6762,N_6650,N_6633);
and U6763 (N_6763,N_6651,N_6657);
and U6764 (N_6764,N_6629,N_6611);
and U6765 (N_6765,N_6670,N_6682);
or U6766 (N_6766,N_6675,N_6669);
nand U6767 (N_6767,N_6690,N_6694);
nand U6768 (N_6768,N_6686,N_6611);
nor U6769 (N_6769,N_6613,N_6667);
or U6770 (N_6770,N_6624,N_6677);
xnor U6771 (N_6771,N_6607,N_6635);
nor U6772 (N_6772,N_6638,N_6628);
nand U6773 (N_6773,N_6675,N_6635);
xor U6774 (N_6774,N_6634,N_6674);
xnor U6775 (N_6775,N_6682,N_6681);
xor U6776 (N_6776,N_6648,N_6652);
xnor U6777 (N_6777,N_6684,N_6642);
and U6778 (N_6778,N_6667,N_6697);
xnor U6779 (N_6779,N_6673,N_6614);
and U6780 (N_6780,N_6696,N_6606);
or U6781 (N_6781,N_6669,N_6617);
xor U6782 (N_6782,N_6699,N_6676);
nor U6783 (N_6783,N_6655,N_6643);
and U6784 (N_6784,N_6610,N_6660);
or U6785 (N_6785,N_6647,N_6678);
nor U6786 (N_6786,N_6634,N_6673);
and U6787 (N_6787,N_6664,N_6651);
xor U6788 (N_6788,N_6697,N_6662);
nand U6789 (N_6789,N_6631,N_6628);
nor U6790 (N_6790,N_6638,N_6611);
nor U6791 (N_6791,N_6609,N_6660);
nand U6792 (N_6792,N_6642,N_6634);
nor U6793 (N_6793,N_6618,N_6655);
xnor U6794 (N_6794,N_6656,N_6624);
or U6795 (N_6795,N_6676,N_6662);
nor U6796 (N_6796,N_6622,N_6628);
nand U6797 (N_6797,N_6692,N_6601);
nand U6798 (N_6798,N_6665,N_6632);
xor U6799 (N_6799,N_6633,N_6673);
nor U6800 (N_6800,N_6755,N_6775);
and U6801 (N_6801,N_6793,N_6725);
xor U6802 (N_6802,N_6744,N_6700);
and U6803 (N_6803,N_6754,N_6706);
nor U6804 (N_6804,N_6746,N_6787);
and U6805 (N_6805,N_6734,N_6719);
nor U6806 (N_6806,N_6759,N_6765);
or U6807 (N_6807,N_6756,N_6799);
nand U6808 (N_6808,N_6729,N_6789);
xnor U6809 (N_6809,N_6797,N_6795);
and U6810 (N_6810,N_6742,N_6739);
or U6811 (N_6811,N_6732,N_6714);
nand U6812 (N_6812,N_6713,N_6772);
xor U6813 (N_6813,N_6781,N_6753);
xnor U6814 (N_6814,N_6758,N_6785);
and U6815 (N_6815,N_6716,N_6743);
xor U6816 (N_6816,N_6777,N_6735);
nand U6817 (N_6817,N_6748,N_6733);
nor U6818 (N_6818,N_6710,N_6702);
xnor U6819 (N_6819,N_6778,N_6701);
nand U6820 (N_6820,N_6774,N_6740);
or U6821 (N_6821,N_6711,N_6731);
xnor U6822 (N_6822,N_6783,N_6730);
nand U6823 (N_6823,N_6715,N_6750);
nor U6824 (N_6824,N_6747,N_6738);
or U6825 (N_6825,N_6771,N_6760);
or U6826 (N_6826,N_6752,N_6727);
xnor U6827 (N_6827,N_6769,N_6770);
or U6828 (N_6828,N_6709,N_6764);
xnor U6829 (N_6829,N_6762,N_6717);
or U6830 (N_6830,N_6728,N_6724);
and U6831 (N_6831,N_6720,N_6788);
nand U6832 (N_6832,N_6712,N_6773);
or U6833 (N_6833,N_6703,N_6768);
or U6834 (N_6834,N_6721,N_6708);
nor U6835 (N_6835,N_6780,N_6790);
nand U6836 (N_6836,N_6761,N_6726);
nor U6837 (N_6837,N_6707,N_6763);
nand U6838 (N_6838,N_6798,N_6767);
and U6839 (N_6839,N_6722,N_6704);
and U6840 (N_6840,N_6745,N_6792);
or U6841 (N_6841,N_6796,N_6784);
nor U6842 (N_6842,N_6749,N_6794);
xnor U6843 (N_6843,N_6766,N_6736);
or U6844 (N_6844,N_6776,N_6782);
xnor U6845 (N_6845,N_6737,N_6757);
nor U6846 (N_6846,N_6779,N_6751);
nand U6847 (N_6847,N_6786,N_6723);
nand U6848 (N_6848,N_6705,N_6791);
nor U6849 (N_6849,N_6741,N_6718);
xnor U6850 (N_6850,N_6776,N_6765);
nor U6851 (N_6851,N_6720,N_6768);
nor U6852 (N_6852,N_6763,N_6765);
and U6853 (N_6853,N_6785,N_6704);
xnor U6854 (N_6854,N_6772,N_6783);
nand U6855 (N_6855,N_6795,N_6720);
xnor U6856 (N_6856,N_6710,N_6790);
xnor U6857 (N_6857,N_6715,N_6749);
nand U6858 (N_6858,N_6768,N_6740);
xor U6859 (N_6859,N_6702,N_6789);
nor U6860 (N_6860,N_6784,N_6751);
or U6861 (N_6861,N_6727,N_6787);
xor U6862 (N_6862,N_6750,N_6775);
nor U6863 (N_6863,N_6785,N_6786);
and U6864 (N_6864,N_6702,N_6772);
or U6865 (N_6865,N_6747,N_6784);
nand U6866 (N_6866,N_6790,N_6702);
and U6867 (N_6867,N_6794,N_6734);
xor U6868 (N_6868,N_6752,N_6763);
or U6869 (N_6869,N_6791,N_6706);
and U6870 (N_6870,N_6709,N_6761);
nand U6871 (N_6871,N_6788,N_6753);
nor U6872 (N_6872,N_6742,N_6774);
or U6873 (N_6873,N_6705,N_6723);
xor U6874 (N_6874,N_6758,N_6745);
or U6875 (N_6875,N_6791,N_6733);
nor U6876 (N_6876,N_6751,N_6754);
and U6877 (N_6877,N_6751,N_6790);
nor U6878 (N_6878,N_6769,N_6705);
xnor U6879 (N_6879,N_6748,N_6791);
or U6880 (N_6880,N_6733,N_6765);
nand U6881 (N_6881,N_6751,N_6702);
or U6882 (N_6882,N_6709,N_6739);
or U6883 (N_6883,N_6789,N_6719);
nand U6884 (N_6884,N_6774,N_6768);
or U6885 (N_6885,N_6730,N_6740);
nor U6886 (N_6886,N_6765,N_6724);
nand U6887 (N_6887,N_6736,N_6763);
and U6888 (N_6888,N_6729,N_6755);
and U6889 (N_6889,N_6711,N_6782);
nor U6890 (N_6890,N_6747,N_6706);
xor U6891 (N_6891,N_6742,N_6799);
nor U6892 (N_6892,N_6707,N_6777);
xor U6893 (N_6893,N_6777,N_6715);
nor U6894 (N_6894,N_6745,N_6788);
and U6895 (N_6895,N_6704,N_6743);
xor U6896 (N_6896,N_6715,N_6799);
or U6897 (N_6897,N_6790,N_6729);
and U6898 (N_6898,N_6781,N_6702);
xor U6899 (N_6899,N_6754,N_6731);
or U6900 (N_6900,N_6847,N_6817);
nor U6901 (N_6901,N_6875,N_6830);
and U6902 (N_6902,N_6889,N_6822);
xor U6903 (N_6903,N_6800,N_6890);
and U6904 (N_6904,N_6801,N_6862);
and U6905 (N_6905,N_6879,N_6885);
nand U6906 (N_6906,N_6892,N_6818);
and U6907 (N_6907,N_6807,N_6894);
or U6908 (N_6908,N_6828,N_6806);
or U6909 (N_6909,N_6821,N_6881);
nand U6910 (N_6910,N_6874,N_6829);
and U6911 (N_6911,N_6831,N_6868);
and U6912 (N_6912,N_6826,N_6886);
xnor U6913 (N_6913,N_6873,N_6814);
or U6914 (N_6914,N_6880,N_6856);
xor U6915 (N_6915,N_6893,N_6871);
and U6916 (N_6916,N_6857,N_6863);
nor U6917 (N_6917,N_6802,N_6809);
and U6918 (N_6918,N_6858,N_6882);
and U6919 (N_6919,N_6860,N_6841);
and U6920 (N_6920,N_6837,N_6876);
and U6921 (N_6921,N_6811,N_6861);
and U6922 (N_6922,N_6854,N_6812);
nand U6923 (N_6923,N_6855,N_6897);
xnor U6924 (N_6924,N_6842,N_6835);
or U6925 (N_6925,N_6899,N_6804);
nand U6926 (N_6926,N_6816,N_6846);
xor U6927 (N_6927,N_6877,N_6859);
or U6928 (N_6928,N_6891,N_6878);
xnor U6929 (N_6929,N_6827,N_6864);
xnor U6930 (N_6930,N_6838,N_6845);
xnor U6931 (N_6931,N_6808,N_6844);
and U6932 (N_6932,N_6883,N_6836);
xnor U6933 (N_6933,N_6834,N_6810);
xor U6934 (N_6934,N_6896,N_6839);
nor U6935 (N_6935,N_6813,N_6870);
nor U6936 (N_6936,N_6803,N_6850);
nor U6937 (N_6937,N_6898,N_6848);
nand U6938 (N_6938,N_6869,N_6852);
xnor U6939 (N_6939,N_6865,N_6888);
xnor U6940 (N_6940,N_6815,N_6895);
or U6941 (N_6941,N_6823,N_6820);
nand U6942 (N_6942,N_6805,N_6851);
xnor U6943 (N_6943,N_6872,N_6825);
xnor U6944 (N_6944,N_6840,N_6843);
and U6945 (N_6945,N_6819,N_6884);
or U6946 (N_6946,N_6853,N_6849);
nor U6947 (N_6947,N_6832,N_6867);
or U6948 (N_6948,N_6824,N_6887);
nor U6949 (N_6949,N_6833,N_6866);
xnor U6950 (N_6950,N_6870,N_6882);
xnor U6951 (N_6951,N_6890,N_6832);
nand U6952 (N_6952,N_6849,N_6858);
nor U6953 (N_6953,N_6809,N_6883);
nor U6954 (N_6954,N_6854,N_6817);
or U6955 (N_6955,N_6809,N_6820);
or U6956 (N_6956,N_6884,N_6891);
xor U6957 (N_6957,N_6832,N_6810);
and U6958 (N_6958,N_6841,N_6868);
nor U6959 (N_6959,N_6856,N_6882);
and U6960 (N_6960,N_6891,N_6846);
xor U6961 (N_6961,N_6843,N_6803);
nor U6962 (N_6962,N_6896,N_6875);
nor U6963 (N_6963,N_6810,N_6888);
nand U6964 (N_6964,N_6857,N_6853);
xnor U6965 (N_6965,N_6890,N_6850);
nand U6966 (N_6966,N_6837,N_6811);
and U6967 (N_6967,N_6894,N_6805);
and U6968 (N_6968,N_6832,N_6877);
nand U6969 (N_6969,N_6811,N_6888);
nor U6970 (N_6970,N_6823,N_6809);
and U6971 (N_6971,N_6898,N_6895);
xor U6972 (N_6972,N_6843,N_6881);
nand U6973 (N_6973,N_6843,N_6812);
xnor U6974 (N_6974,N_6829,N_6824);
and U6975 (N_6975,N_6829,N_6886);
xor U6976 (N_6976,N_6856,N_6893);
nand U6977 (N_6977,N_6899,N_6805);
and U6978 (N_6978,N_6811,N_6831);
nor U6979 (N_6979,N_6802,N_6863);
nor U6980 (N_6980,N_6823,N_6882);
or U6981 (N_6981,N_6802,N_6803);
and U6982 (N_6982,N_6868,N_6812);
or U6983 (N_6983,N_6893,N_6805);
nor U6984 (N_6984,N_6845,N_6818);
xor U6985 (N_6985,N_6806,N_6878);
nor U6986 (N_6986,N_6816,N_6824);
nor U6987 (N_6987,N_6806,N_6805);
xor U6988 (N_6988,N_6824,N_6890);
and U6989 (N_6989,N_6830,N_6896);
nor U6990 (N_6990,N_6882,N_6886);
xnor U6991 (N_6991,N_6802,N_6870);
or U6992 (N_6992,N_6824,N_6879);
or U6993 (N_6993,N_6848,N_6823);
and U6994 (N_6994,N_6801,N_6861);
or U6995 (N_6995,N_6898,N_6812);
nand U6996 (N_6996,N_6887,N_6814);
or U6997 (N_6997,N_6878,N_6841);
nor U6998 (N_6998,N_6829,N_6890);
nor U6999 (N_6999,N_6888,N_6822);
nand U7000 (N_7000,N_6936,N_6902);
nor U7001 (N_7001,N_6953,N_6974);
and U7002 (N_7002,N_6991,N_6919);
nand U7003 (N_7003,N_6926,N_6925);
and U7004 (N_7004,N_6927,N_6978);
xnor U7005 (N_7005,N_6966,N_6999);
or U7006 (N_7006,N_6943,N_6921);
xor U7007 (N_7007,N_6982,N_6907);
nor U7008 (N_7008,N_6923,N_6979);
xor U7009 (N_7009,N_6914,N_6901);
nor U7010 (N_7010,N_6985,N_6964);
xnor U7011 (N_7011,N_6983,N_6946);
xnor U7012 (N_7012,N_6909,N_6935);
xor U7013 (N_7013,N_6910,N_6951);
and U7014 (N_7014,N_6960,N_6992);
xnor U7015 (N_7015,N_6988,N_6931);
xnor U7016 (N_7016,N_6934,N_6958);
or U7017 (N_7017,N_6913,N_6957);
and U7018 (N_7018,N_6916,N_6937);
and U7019 (N_7019,N_6994,N_6917);
or U7020 (N_7020,N_6924,N_6980);
nand U7021 (N_7021,N_6948,N_6963);
nand U7022 (N_7022,N_6969,N_6971);
or U7023 (N_7023,N_6904,N_6947);
nor U7024 (N_7024,N_6911,N_6959);
nand U7025 (N_7025,N_6965,N_6920);
nand U7026 (N_7026,N_6922,N_6950);
nor U7027 (N_7027,N_6976,N_6900);
or U7028 (N_7028,N_6955,N_6952);
or U7029 (N_7029,N_6908,N_6929);
and U7030 (N_7030,N_6990,N_6970);
nand U7031 (N_7031,N_6981,N_6915);
xnor U7032 (N_7032,N_6918,N_6998);
or U7033 (N_7033,N_6996,N_6944);
nand U7034 (N_7034,N_6939,N_6940);
and U7035 (N_7035,N_6962,N_6972);
nor U7036 (N_7036,N_6997,N_6930);
xor U7037 (N_7037,N_6956,N_6928);
nand U7038 (N_7038,N_6932,N_6975);
and U7039 (N_7039,N_6954,N_6905);
xnor U7040 (N_7040,N_6986,N_6973);
nand U7041 (N_7041,N_6912,N_6987);
or U7042 (N_7042,N_6933,N_6949);
xor U7043 (N_7043,N_6995,N_6977);
nor U7044 (N_7044,N_6942,N_6989);
nand U7045 (N_7045,N_6961,N_6906);
xor U7046 (N_7046,N_6968,N_6941);
and U7047 (N_7047,N_6993,N_6903);
and U7048 (N_7048,N_6984,N_6945);
and U7049 (N_7049,N_6967,N_6938);
nor U7050 (N_7050,N_6989,N_6984);
nand U7051 (N_7051,N_6938,N_6913);
or U7052 (N_7052,N_6977,N_6987);
xnor U7053 (N_7053,N_6919,N_6963);
or U7054 (N_7054,N_6957,N_6943);
xnor U7055 (N_7055,N_6976,N_6998);
nor U7056 (N_7056,N_6906,N_6953);
xnor U7057 (N_7057,N_6921,N_6993);
nand U7058 (N_7058,N_6976,N_6913);
nor U7059 (N_7059,N_6992,N_6941);
or U7060 (N_7060,N_6959,N_6918);
and U7061 (N_7061,N_6963,N_6990);
or U7062 (N_7062,N_6900,N_6938);
nand U7063 (N_7063,N_6941,N_6971);
nor U7064 (N_7064,N_6942,N_6903);
nand U7065 (N_7065,N_6937,N_6950);
xnor U7066 (N_7066,N_6911,N_6993);
nor U7067 (N_7067,N_6912,N_6946);
and U7068 (N_7068,N_6966,N_6988);
and U7069 (N_7069,N_6928,N_6999);
nor U7070 (N_7070,N_6916,N_6985);
nand U7071 (N_7071,N_6972,N_6926);
nand U7072 (N_7072,N_6935,N_6944);
and U7073 (N_7073,N_6968,N_6934);
nand U7074 (N_7074,N_6980,N_6937);
nor U7075 (N_7075,N_6955,N_6909);
nor U7076 (N_7076,N_6905,N_6924);
nand U7077 (N_7077,N_6973,N_6992);
or U7078 (N_7078,N_6956,N_6908);
xor U7079 (N_7079,N_6956,N_6997);
and U7080 (N_7080,N_6948,N_6954);
nand U7081 (N_7081,N_6999,N_6959);
and U7082 (N_7082,N_6916,N_6999);
and U7083 (N_7083,N_6947,N_6982);
xor U7084 (N_7084,N_6925,N_6959);
or U7085 (N_7085,N_6931,N_6972);
xnor U7086 (N_7086,N_6949,N_6974);
and U7087 (N_7087,N_6973,N_6957);
xor U7088 (N_7088,N_6931,N_6934);
and U7089 (N_7089,N_6971,N_6953);
nand U7090 (N_7090,N_6918,N_6912);
nand U7091 (N_7091,N_6956,N_6949);
nand U7092 (N_7092,N_6966,N_6962);
nand U7093 (N_7093,N_6914,N_6996);
nand U7094 (N_7094,N_6994,N_6999);
nand U7095 (N_7095,N_6913,N_6919);
and U7096 (N_7096,N_6942,N_6969);
and U7097 (N_7097,N_6945,N_6948);
nor U7098 (N_7098,N_6913,N_6981);
nor U7099 (N_7099,N_6945,N_6962);
xor U7100 (N_7100,N_7035,N_7004);
and U7101 (N_7101,N_7039,N_7001);
xnor U7102 (N_7102,N_7064,N_7014);
nor U7103 (N_7103,N_7029,N_7028);
xnor U7104 (N_7104,N_7078,N_7036);
and U7105 (N_7105,N_7037,N_7056);
xor U7106 (N_7106,N_7043,N_7055);
and U7107 (N_7107,N_7032,N_7025);
and U7108 (N_7108,N_7099,N_7005);
nor U7109 (N_7109,N_7031,N_7017);
nor U7110 (N_7110,N_7093,N_7098);
nor U7111 (N_7111,N_7076,N_7053);
or U7112 (N_7112,N_7050,N_7080);
nand U7113 (N_7113,N_7022,N_7047);
nor U7114 (N_7114,N_7008,N_7075);
nor U7115 (N_7115,N_7010,N_7018);
and U7116 (N_7116,N_7045,N_7069);
or U7117 (N_7117,N_7074,N_7067);
and U7118 (N_7118,N_7003,N_7042);
nor U7119 (N_7119,N_7086,N_7051);
nor U7120 (N_7120,N_7044,N_7012);
xor U7121 (N_7121,N_7068,N_7092);
xor U7122 (N_7122,N_7024,N_7002);
and U7123 (N_7123,N_7020,N_7090);
nand U7124 (N_7124,N_7011,N_7006);
xnor U7125 (N_7125,N_7073,N_7089);
nor U7126 (N_7126,N_7065,N_7041);
or U7127 (N_7127,N_7081,N_7058);
nor U7128 (N_7128,N_7033,N_7009);
and U7129 (N_7129,N_7083,N_7097);
nor U7130 (N_7130,N_7070,N_7057);
nor U7131 (N_7131,N_7054,N_7040);
xnor U7132 (N_7132,N_7013,N_7052);
or U7133 (N_7133,N_7034,N_7071);
xnor U7134 (N_7134,N_7061,N_7096);
or U7135 (N_7135,N_7016,N_7079);
xor U7136 (N_7136,N_7000,N_7019);
or U7137 (N_7137,N_7027,N_7049);
and U7138 (N_7138,N_7038,N_7091);
and U7139 (N_7139,N_7059,N_7095);
nor U7140 (N_7140,N_7007,N_7060);
xnor U7141 (N_7141,N_7066,N_7085);
nor U7142 (N_7142,N_7023,N_7030);
or U7143 (N_7143,N_7077,N_7021);
or U7144 (N_7144,N_7026,N_7048);
or U7145 (N_7145,N_7046,N_7082);
and U7146 (N_7146,N_7063,N_7087);
or U7147 (N_7147,N_7094,N_7088);
nor U7148 (N_7148,N_7062,N_7084);
or U7149 (N_7149,N_7072,N_7015);
nor U7150 (N_7150,N_7012,N_7061);
xnor U7151 (N_7151,N_7045,N_7091);
xnor U7152 (N_7152,N_7069,N_7061);
nor U7153 (N_7153,N_7043,N_7009);
xor U7154 (N_7154,N_7098,N_7004);
nand U7155 (N_7155,N_7059,N_7084);
nand U7156 (N_7156,N_7080,N_7040);
xor U7157 (N_7157,N_7054,N_7019);
xor U7158 (N_7158,N_7005,N_7038);
xor U7159 (N_7159,N_7056,N_7010);
or U7160 (N_7160,N_7074,N_7039);
xnor U7161 (N_7161,N_7097,N_7085);
nor U7162 (N_7162,N_7080,N_7090);
nor U7163 (N_7163,N_7064,N_7063);
or U7164 (N_7164,N_7050,N_7014);
and U7165 (N_7165,N_7058,N_7086);
and U7166 (N_7166,N_7091,N_7065);
and U7167 (N_7167,N_7047,N_7046);
nor U7168 (N_7168,N_7074,N_7046);
or U7169 (N_7169,N_7082,N_7048);
nand U7170 (N_7170,N_7080,N_7057);
and U7171 (N_7171,N_7038,N_7053);
nand U7172 (N_7172,N_7010,N_7036);
nor U7173 (N_7173,N_7093,N_7086);
and U7174 (N_7174,N_7015,N_7074);
nor U7175 (N_7175,N_7087,N_7007);
xor U7176 (N_7176,N_7013,N_7016);
and U7177 (N_7177,N_7069,N_7009);
nor U7178 (N_7178,N_7008,N_7065);
or U7179 (N_7179,N_7094,N_7082);
or U7180 (N_7180,N_7089,N_7052);
or U7181 (N_7181,N_7021,N_7034);
xnor U7182 (N_7182,N_7037,N_7099);
nand U7183 (N_7183,N_7040,N_7004);
nor U7184 (N_7184,N_7073,N_7093);
xor U7185 (N_7185,N_7003,N_7074);
or U7186 (N_7186,N_7097,N_7081);
xor U7187 (N_7187,N_7071,N_7072);
nand U7188 (N_7188,N_7078,N_7097);
nor U7189 (N_7189,N_7018,N_7085);
nand U7190 (N_7190,N_7086,N_7032);
nand U7191 (N_7191,N_7071,N_7044);
and U7192 (N_7192,N_7070,N_7073);
xnor U7193 (N_7193,N_7068,N_7029);
nand U7194 (N_7194,N_7021,N_7092);
xor U7195 (N_7195,N_7066,N_7006);
and U7196 (N_7196,N_7050,N_7078);
nor U7197 (N_7197,N_7016,N_7099);
and U7198 (N_7198,N_7094,N_7076);
xor U7199 (N_7199,N_7096,N_7065);
or U7200 (N_7200,N_7137,N_7169);
and U7201 (N_7201,N_7194,N_7132);
or U7202 (N_7202,N_7157,N_7148);
and U7203 (N_7203,N_7166,N_7183);
or U7204 (N_7204,N_7177,N_7156);
nor U7205 (N_7205,N_7143,N_7184);
nand U7206 (N_7206,N_7149,N_7173);
xnor U7207 (N_7207,N_7117,N_7175);
and U7208 (N_7208,N_7134,N_7159);
or U7209 (N_7209,N_7139,N_7171);
or U7210 (N_7210,N_7112,N_7146);
or U7211 (N_7211,N_7118,N_7103);
xor U7212 (N_7212,N_7123,N_7174);
or U7213 (N_7213,N_7193,N_7119);
nor U7214 (N_7214,N_7172,N_7108);
nor U7215 (N_7215,N_7100,N_7182);
nand U7216 (N_7216,N_7167,N_7135);
xor U7217 (N_7217,N_7114,N_7142);
nand U7218 (N_7218,N_7136,N_7107);
or U7219 (N_7219,N_7187,N_7185);
and U7220 (N_7220,N_7162,N_7198);
nor U7221 (N_7221,N_7105,N_7106);
nand U7222 (N_7222,N_7195,N_7120);
or U7223 (N_7223,N_7168,N_7115);
nor U7224 (N_7224,N_7186,N_7141);
xor U7225 (N_7225,N_7155,N_7192);
and U7226 (N_7226,N_7113,N_7165);
or U7227 (N_7227,N_7178,N_7191);
or U7228 (N_7228,N_7179,N_7180);
nand U7229 (N_7229,N_7121,N_7197);
xnor U7230 (N_7230,N_7170,N_7122);
nor U7231 (N_7231,N_7164,N_7125);
or U7232 (N_7232,N_7127,N_7147);
nand U7233 (N_7233,N_7181,N_7140);
or U7234 (N_7234,N_7153,N_7109);
nand U7235 (N_7235,N_7188,N_7199);
and U7236 (N_7236,N_7128,N_7126);
and U7237 (N_7237,N_7152,N_7129);
nand U7238 (N_7238,N_7110,N_7130);
xnor U7239 (N_7239,N_7160,N_7150);
xnor U7240 (N_7240,N_7131,N_7124);
and U7241 (N_7241,N_7138,N_7145);
nand U7242 (N_7242,N_7158,N_7161);
and U7243 (N_7243,N_7111,N_7104);
nand U7244 (N_7244,N_7163,N_7102);
xor U7245 (N_7245,N_7133,N_7196);
and U7246 (N_7246,N_7154,N_7189);
nor U7247 (N_7247,N_7144,N_7176);
nor U7248 (N_7248,N_7190,N_7151);
xor U7249 (N_7249,N_7101,N_7116);
or U7250 (N_7250,N_7100,N_7124);
xor U7251 (N_7251,N_7118,N_7116);
or U7252 (N_7252,N_7138,N_7190);
and U7253 (N_7253,N_7182,N_7102);
xnor U7254 (N_7254,N_7182,N_7148);
or U7255 (N_7255,N_7174,N_7108);
and U7256 (N_7256,N_7169,N_7127);
nand U7257 (N_7257,N_7186,N_7134);
nor U7258 (N_7258,N_7108,N_7159);
nand U7259 (N_7259,N_7136,N_7175);
nand U7260 (N_7260,N_7167,N_7186);
nand U7261 (N_7261,N_7168,N_7100);
xor U7262 (N_7262,N_7112,N_7106);
or U7263 (N_7263,N_7175,N_7141);
xor U7264 (N_7264,N_7175,N_7106);
or U7265 (N_7265,N_7120,N_7167);
xor U7266 (N_7266,N_7108,N_7130);
nor U7267 (N_7267,N_7186,N_7170);
nor U7268 (N_7268,N_7106,N_7167);
nor U7269 (N_7269,N_7124,N_7144);
or U7270 (N_7270,N_7136,N_7187);
nor U7271 (N_7271,N_7126,N_7110);
nand U7272 (N_7272,N_7179,N_7148);
xor U7273 (N_7273,N_7177,N_7164);
nor U7274 (N_7274,N_7149,N_7199);
nor U7275 (N_7275,N_7191,N_7198);
and U7276 (N_7276,N_7170,N_7103);
nand U7277 (N_7277,N_7128,N_7156);
nor U7278 (N_7278,N_7154,N_7196);
xor U7279 (N_7279,N_7133,N_7109);
xnor U7280 (N_7280,N_7126,N_7115);
nand U7281 (N_7281,N_7192,N_7112);
nor U7282 (N_7282,N_7100,N_7150);
xnor U7283 (N_7283,N_7104,N_7193);
nand U7284 (N_7284,N_7173,N_7108);
nand U7285 (N_7285,N_7193,N_7195);
and U7286 (N_7286,N_7148,N_7118);
nor U7287 (N_7287,N_7116,N_7112);
and U7288 (N_7288,N_7175,N_7142);
nand U7289 (N_7289,N_7162,N_7127);
xnor U7290 (N_7290,N_7147,N_7120);
xor U7291 (N_7291,N_7185,N_7101);
xnor U7292 (N_7292,N_7197,N_7128);
and U7293 (N_7293,N_7124,N_7166);
and U7294 (N_7294,N_7147,N_7151);
nor U7295 (N_7295,N_7190,N_7152);
or U7296 (N_7296,N_7183,N_7104);
and U7297 (N_7297,N_7179,N_7163);
xor U7298 (N_7298,N_7163,N_7152);
and U7299 (N_7299,N_7183,N_7191);
xnor U7300 (N_7300,N_7238,N_7290);
and U7301 (N_7301,N_7273,N_7218);
and U7302 (N_7302,N_7237,N_7266);
nand U7303 (N_7303,N_7228,N_7270);
xor U7304 (N_7304,N_7264,N_7234);
nor U7305 (N_7305,N_7274,N_7253);
nor U7306 (N_7306,N_7254,N_7250);
and U7307 (N_7307,N_7229,N_7241);
nor U7308 (N_7308,N_7246,N_7239);
nand U7309 (N_7309,N_7226,N_7277);
and U7310 (N_7310,N_7262,N_7242);
xnor U7311 (N_7311,N_7208,N_7296);
xor U7312 (N_7312,N_7295,N_7215);
nor U7313 (N_7313,N_7224,N_7235);
xnor U7314 (N_7314,N_7271,N_7269);
nand U7315 (N_7315,N_7275,N_7200);
nand U7316 (N_7316,N_7223,N_7207);
nand U7317 (N_7317,N_7248,N_7217);
nand U7318 (N_7318,N_7272,N_7203);
or U7319 (N_7319,N_7268,N_7287);
nor U7320 (N_7320,N_7256,N_7243);
xnor U7321 (N_7321,N_7214,N_7219);
xor U7322 (N_7322,N_7299,N_7288);
nand U7323 (N_7323,N_7213,N_7282);
or U7324 (N_7324,N_7210,N_7281);
nand U7325 (N_7325,N_7244,N_7258);
or U7326 (N_7326,N_7216,N_7212);
nor U7327 (N_7327,N_7286,N_7204);
or U7328 (N_7328,N_7280,N_7221);
nor U7329 (N_7329,N_7202,N_7261);
and U7330 (N_7330,N_7249,N_7259);
nor U7331 (N_7331,N_7267,N_7201);
nor U7332 (N_7332,N_7245,N_7236);
or U7333 (N_7333,N_7209,N_7220);
and U7334 (N_7334,N_7230,N_7285);
nand U7335 (N_7335,N_7247,N_7205);
and U7336 (N_7336,N_7206,N_7227);
xor U7337 (N_7337,N_7279,N_7251);
nand U7338 (N_7338,N_7252,N_7225);
nor U7339 (N_7339,N_7257,N_7292);
and U7340 (N_7340,N_7265,N_7289);
nand U7341 (N_7341,N_7294,N_7232);
or U7342 (N_7342,N_7297,N_7276);
xnor U7343 (N_7343,N_7260,N_7263);
nor U7344 (N_7344,N_7233,N_7255);
nand U7345 (N_7345,N_7240,N_7278);
or U7346 (N_7346,N_7211,N_7231);
or U7347 (N_7347,N_7293,N_7298);
and U7348 (N_7348,N_7284,N_7222);
and U7349 (N_7349,N_7283,N_7291);
nand U7350 (N_7350,N_7233,N_7225);
nand U7351 (N_7351,N_7265,N_7213);
nand U7352 (N_7352,N_7259,N_7244);
xnor U7353 (N_7353,N_7219,N_7230);
and U7354 (N_7354,N_7219,N_7242);
or U7355 (N_7355,N_7290,N_7253);
xor U7356 (N_7356,N_7273,N_7238);
nand U7357 (N_7357,N_7264,N_7251);
or U7358 (N_7358,N_7213,N_7242);
or U7359 (N_7359,N_7284,N_7225);
xor U7360 (N_7360,N_7241,N_7279);
or U7361 (N_7361,N_7258,N_7230);
xor U7362 (N_7362,N_7243,N_7286);
nand U7363 (N_7363,N_7211,N_7224);
and U7364 (N_7364,N_7271,N_7213);
nand U7365 (N_7365,N_7285,N_7222);
nor U7366 (N_7366,N_7267,N_7210);
xor U7367 (N_7367,N_7216,N_7268);
xnor U7368 (N_7368,N_7256,N_7297);
nor U7369 (N_7369,N_7220,N_7259);
nand U7370 (N_7370,N_7223,N_7288);
xnor U7371 (N_7371,N_7265,N_7211);
or U7372 (N_7372,N_7263,N_7276);
and U7373 (N_7373,N_7240,N_7257);
nor U7374 (N_7374,N_7210,N_7261);
and U7375 (N_7375,N_7208,N_7212);
xnor U7376 (N_7376,N_7269,N_7207);
or U7377 (N_7377,N_7271,N_7237);
or U7378 (N_7378,N_7270,N_7298);
xnor U7379 (N_7379,N_7273,N_7274);
or U7380 (N_7380,N_7250,N_7298);
xnor U7381 (N_7381,N_7272,N_7209);
xor U7382 (N_7382,N_7297,N_7259);
nor U7383 (N_7383,N_7202,N_7235);
and U7384 (N_7384,N_7286,N_7221);
nand U7385 (N_7385,N_7200,N_7216);
and U7386 (N_7386,N_7290,N_7223);
and U7387 (N_7387,N_7261,N_7291);
nand U7388 (N_7388,N_7204,N_7228);
nor U7389 (N_7389,N_7245,N_7239);
and U7390 (N_7390,N_7273,N_7277);
xor U7391 (N_7391,N_7228,N_7254);
or U7392 (N_7392,N_7259,N_7298);
nor U7393 (N_7393,N_7262,N_7241);
nand U7394 (N_7394,N_7212,N_7250);
xnor U7395 (N_7395,N_7246,N_7232);
nand U7396 (N_7396,N_7260,N_7261);
and U7397 (N_7397,N_7278,N_7202);
nor U7398 (N_7398,N_7231,N_7214);
xnor U7399 (N_7399,N_7285,N_7295);
or U7400 (N_7400,N_7317,N_7301);
and U7401 (N_7401,N_7366,N_7340);
xor U7402 (N_7402,N_7342,N_7363);
nor U7403 (N_7403,N_7381,N_7364);
or U7404 (N_7404,N_7356,N_7350);
or U7405 (N_7405,N_7353,N_7390);
nor U7406 (N_7406,N_7307,N_7369);
xnor U7407 (N_7407,N_7338,N_7303);
or U7408 (N_7408,N_7341,N_7377);
or U7409 (N_7409,N_7359,N_7360);
nor U7410 (N_7410,N_7352,N_7371);
nor U7411 (N_7411,N_7302,N_7330);
and U7412 (N_7412,N_7329,N_7361);
xnor U7413 (N_7413,N_7395,N_7374);
nand U7414 (N_7414,N_7368,N_7305);
nand U7415 (N_7415,N_7336,N_7322);
nand U7416 (N_7416,N_7370,N_7345);
or U7417 (N_7417,N_7397,N_7357);
xnor U7418 (N_7418,N_7367,N_7316);
nand U7419 (N_7419,N_7326,N_7324);
nor U7420 (N_7420,N_7319,N_7398);
nand U7421 (N_7421,N_7393,N_7348);
xor U7422 (N_7422,N_7333,N_7378);
nor U7423 (N_7423,N_7313,N_7396);
nand U7424 (N_7424,N_7391,N_7321);
nand U7425 (N_7425,N_7347,N_7300);
nor U7426 (N_7426,N_7388,N_7335);
nand U7427 (N_7427,N_7339,N_7354);
or U7428 (N_7428,N_7355,N_7394);
nand U7429 (N_7429,N_7306,N_7349);
and U7430 (N_7430,N_7323,N_7332);
and U7431 (N_7431,N_7351,N_7383);
or U7432 (N_7432,N_7314,N_7365);
or U7433 (N_7433,N_7318,N_7325);
xnor U7434 (N_7434,N_7386,N_7337);
nor U7435 (N_7435,N_7344,N_7311);
xnor U7436 (N_7436,N_7379,N_7327);
nand U7437 (N_7437,N_7389,N_7372);
and U7438 (N_7438,N_7315,N_7308);
nand U7439 (N_7439,N_7392,N_7343);
xor U7440 (N_7440,N_7309,N_7328);
nor U7441 (N_7441,N_7312,N_7358);
nor U7442 (N_7442,N_7380,N_7375);
nor U7443 (N_7443,N_7320,N_7362);
xnor U7444 (N_7444,N_7385,N_7346);
and U7445 (N_7445,N_7376,N_7373);
nor U7446 (N_7446,N_7334,N_7310);
and U7447 (N_7447,N_7382,N_7384);
or U7448 (N_7448,N_7304,N_7399);
xor U7449 (N_7449,N_7331,N_7387);
or U7450 (N_7450,N_7375,N_7324);
or U7451 (N_7451,N_7330,N_7350);
nor U7452 (N_7452,N_7341,N_7311);
nor U7453 (N_7453,N_7328,N_7333);
nor U7454 (N_7454,N_7392,N_7361);
and U7455 (N_7455,N_7390,N_7340);
xor U7456 (N_7456,N_7398,N_7349);
and U7457 (N_7457,N_7381,N_7390);
nand U7458 (N_7458,N_7391,N_7399);
or U7459 (N_7459,N_7304,N_7397);
nor U7460 (N_7460,N_7310,N_7383);
and U7461 (N_7461,N_7386,N_7378);
or U7462 (N_7462,N_7368,N_7321);
nor U7463 (N_7463,N_7303,N_7359);
nor U7464 (N_7464,N_7360,N_7326);
nor U7465 (N_7465,N_7328,N_7357);
or U7466 (N_7466,N_7327,N_7310);
nor U7467 (N_7467,N_7374,N_7323);
nand U7468 (N_7468,N_7371,N_7350);
or U7469 (N_7469,N_7394,N_7322);
or U7470 (N_7470,N_7361,N_7338);
and U7471 (N_7471,N_7308,N_7370);
and U7472 (N_7472,N_7320,N_7317);
and U7473 (N_7473,N_7363,N_7357);
xor U7474 (N_7474,N_7350,N_7322);
xnor U7475 (N_7475,N_7377,N_7395);
or U7476 (N_7476,N_7335,N_7369);
and U7477 (N_7477,N_7342,N_7382);
or U7478 (N_7478,N_7353,N_7335);
or U7479 (N_7479,N_7388,N_7310);
and U7480 (N_7480,N_7336,N_7385);
and U7481 (N_7481,N_7395,N_7366);
and U7482 (N_7482,N_7356,N_7312);
or U7483 (N_7483,N_7360,N_7303);
or U7484 (N_7484,N_7363,N_7320);
or U7485 (N_7485,N_7396,N_7367);
xor U7486 (N_7486,N_7303,N_7372);
xnor U7487 (N_7487,N_7399,N_7383);
nand U7488 (N_7488,N_7370,N_7304);
xor U7489 (N_7489,N_7329,N_7343);
or U7490 (N_7490,N_7362,N_7336);
and U7491 (N_7491,N_7348,N_7330);
nand U7492 (N_7492,N_7385,N_7398);
or U7493 (N_7493,N_7362,N_7303);
nand U7494 (N_7494,N_7371,N_7337);
nand U7495 (N_7495,N_7334,N_7361);
and U7496 (N_7496,N_7306,N_7376);
nand U7497 (N_7497,N_7329,N_7310);
nor U7498 (N_7498,N_7359,N_7373);
xnor U7499 (N_7499,N_7314,N_7375);
nand U7500 (N_7500,N_7455,N_7444);
and U7501 (N_7501,N_7412,N_7452);
and U7502 (N_7502,N_7484,N_7460);
xnor U7503 (N_7503,N_7401,N_7470);
or U7504 (N_7504,N_7417,N_7447);
nand U7505 (N_7505,N_7402,N_7481);
and U7506 (N_7506,N_7420,N_7410);
nor U7507 (N_7507,N_7445,N_7498);
and U7508 (N_7508,N_7495,N_7450);
and U7509 (N_7509,N_7487,N_7449);
xor U7510 (N_7510,N_7427,N_7482);
or U7511 (N_7511,N_7461,N_7467);
nor U7512 (N_7512,N_7439,N_7476);
or U7513 (N_7513,N_7400,N_7490);
and U7514 (N_7514,N_7413,N_7422);
nand U7515 (N_7515,N_7443,N_7474);
or U7516 (N_7516,N_7463,N_7434);
and U7517 (N_7517,N_7414,N_7441);
or U7518 (N_7518,N_7471,N_7426);
xnor U7519 (N_7519,N_7469,N_7408);
nor U7520 (N_7520,N_7483,N_7462);
nor U7521 (N_7521,N_7451,N_7403);
nand U7522 (N_7522,N_7453,N_7488);
nor U7523 (N_7523,N_7480,N_7423);
xnor U7524 (N_7524,N_7416,N_7466);
nor U7525 (N_7525,N_7475,N_7431);
and U7526 (N_7526,N_7485,N_7468);
or U7527 (N_7527,N_7492,N_7433);
nand U7528 (N_7528,N_7419,N_7440);
and U7529 (N_7529,N_7454,N_7457);
xor U7530 (N_7530,N_7465,N_7429);
and U7531 (N_7531,N_7478,N_7493);
nor U7532 (N_7532,N_7486,N_7424);
nand U7533 (N_7533,N_7407,N_7415);
nand U7534 (N_7534,N_7437,N_7496);
nor U7535 (N_7535,N_7494,N_7491);
xnor U7536 (N_7536,N_7499,N_7473);
xnor U7537 (N_7537,N_7442,N_7438);
xnor U7538 (N_7538,N_7406,N_7497);
nand U7539 (N_7539,N_7428,N_7459);
xnor U7540 (N_7540,N_7418,N_7405);
xor U7541 (N_7541,N_7446,N_7404);
nor U7542 (N_7542,N_7430,N_7456);
or U7543 (N_7543,N_7458,N_7435);
nand U7544 (N_7544,N_7436,N_7477);
and U7545 (N_7545,N_7421,N_7411);
nand U7546 (N_7546,N_7432,N_7409);
or U7547 (N_7547,N_7448,N_7425);
nand U7548 (N_7548,N_7489,N_7479);
xor U7549 (N_7549,N_7472,N_7464);
nand U7550 (N_7550,N_7446,N_7484);
xnor U7551 (N_7551,N_7487,N_7419);
and U7552 (N_7552,N_7464,N_7444);
nand U7553 (N_7553,N_7404,N_7442);
and U7554 (N_7554,N_7415,N_7468);
nand U7555 (N_7555,N_7462,N_7472);
nor U7556 (N_7556,N_7481,N_7423);
nor U7557 (N_7557,N_7402,N_7453);
xor U7558 (N_7558,N_7480,N_7407);
and U7559 (N_7559,N_7424,N_7472);
or U7560 (N_7560,N_7498,N_7444);
xnor U7561 (N_7561,N_7402,N_7464);
nor U7562 (N_7562,N_7445,N_7441);
xnor U7563 (N_7563,N_7419,N_7444);
or U7564 (N_7564,N_7469,N_7424);
nand U7565 (N_7565,N_7436,N_7476);
xor U7566 (N_7566,N_7422,N_7402);
nand U7567 (N_7567,N_7474,N_7432);
and U7568 (N_7568,N_7481,N_7446);
xnor U7569 (N_7569,N_7415,N_7422);
nand U7570 (N_7570,N_7482,N_7433);
nor U7571 (N_7571,N_7429,N_7412);
nor U7572 (N_7572,N_7406,N_7456);
or U7573 (N_7573,N_7494,N_7467);
xnor U7574 (N_7574,N_7423,N_7498);
xor U7575 (N_7575,N_7439,N_7408);
xnor U7576 (N_7576,N_7434,N_7479);
and U7577 (N_7577,N_7450,N_7468);
nand U7578 (N_7578,N_7452,N_7436);
nand U7579 (N_7579,N_7439,N_7471);
and U7580 (N_7580,N_7465,N_7475);
and U7581 (N_7581,N_7469,N_7478);
nand U7582 (N_7582,N_7431,N_7459);
nand U7583 (N_7583,N_7401,N_7400);
and U7584 (N_7584,N_7498,N_7449);
nor U7585 (N_7585,N_7473,N_7455);
nor U7586 (N_7586,N_7462,N_7454);
xor U7587 (N_7587,N_7450,N_7429);
and U7588 (N_7588,N_7430,N_7476);
xnor U7589 (N_7589,N_7424,N_7462);
nor U7590 (N_7590,N_7495,N_7422);
nand U7591 (N_7591,N_7438,N_7420);
xor U7592 (N_7592,N_7486,N_7478);
xnor U7593 (N_7593,N_7486,N_7409);
nor U7594 (N_7594,N_7495,N_7470);
nor U7595 (N_7595,N_7441,N_7402);
and U7596 (N_7596,N_7494,N_7456);
xor U7597 (N_7597,N_7415,N_7452);
nand U7598 (N_7598,N_7419,N_7438);
and U7599 (N_7599,N_7433,N_7478);
nor U7600 (N_7600,N_7501,N_7545);
or U7601 (N_7601,N_7574,N_7576);
nor U7602 (N_7602,N_7573,N_7528);
xnor U7603 (N_7603,N_7555,N_7580);
or U7604 (N_7604,N_7527,N_7548);
xor U7605 (N_7605,N_7549,N_7592);
or U7606 (N_7606,N_7599,N_7591);
or U7607 (N_7607,N_7500,N_7522);
xor U7608 (N_7608,N_7565,N_7561);
or U7609 (N_7609,N_7582,N_7550);
xor U7610 (N_7610,N_7568,N_7532);
nand U7611 (N_7611,N_7577,N_7514);
or U7612 (N_7612,N_7571,N_7579);
xnor U7613 (N_7613,N_7583,N_7556);
and U7614 (N_7614,N_7525,N_7590);
nor U7615 (N_7615,N_7569,N_7533);
nand U7616 (N_7616,N_7524,N_7529);
nor U7617 (N_7617,N_7538,N_7523);
xor U7618 (N_7618,N_7503,N_7530);
xor U7619 (N_7619,N_7560,N_7512);
and U7620 (N_7620,N_7589,N_7507);
and U7621 (N_7621,N_7534,N_7519);
nor U7622 (N_7622,N_7557,N_7513);
nor U7623 (N_7623,N_7578,N_7593);
and U7624 (N_7624,N_7517,N_7510);
xor U7625 (N_7625,N_7515,N_7588);
nand U7626 (N_7626,N_7572,N_7508);
and U7627 (N_7627,N_7520,N_7506);
or U7628 (N_7628,N_7558,N_7543);
and U7629 (N_7629,N_7585,N_7547);
nand U7630 (N_7630,N_7502,N_7567);
xnor U7631 (N_7631,N_7584,N_7544);
nand U7632 (N_7632,N_7505,N_7553);
xnor U7633 (N_7633,N_7563,N_7597);
nand U7634 (N_7634,N_7540,N_7541);
nor U7635 (N_7635,N_7594,N_7581);
nor U7636 (N_7636,N_7554,N_7537);
nor U7637 (N_7637,N_7516,N_7562);
or U7638 (N_7638,N_7559,N_7509);
or U7639 (N_7639,N_7536,N_7552);
and U7640 (N_7640,N_7504,N_7542);
and U7641 (N_7641,N_7564,N_7596);
and U7642 (N_7642,N_7595,N_7521);
nand U7643 (N_7643,N_7598,N_7586);
and U7644 (N_7644,N_7566,N_7575);
nor U7645 (N_7645,N_7587,N_7570);
xor U7646 (N_7646,N_7511,N_7535);
or U7647 (N_7647,N_7531,N_7518);
xnor U7648 (N_7648,N_7539,N_7551);
nand U7649 (N_7649,N_7526,N_7546);
and U7650 (N_7650,N_7516,N_7514);
and U7651 (N_7651,N_7597,N_7576);
and U7652 (N_7652,N_7525,N_7561);
and U7653 (N_7653,N_7548,N_7506);
and U7654 (N_7654,N_7572,N_7502);
or U7655 (N_7655,N_7546,N_7501);
or U7656 (N_7656,N_7500,N_7532);
nor U7657 (N_7657,N_7554,N_7560);
or U7658 (N_7658,N_7592,N_7579);
or U7659 (N_7659,N_7592,N_7557);
and U7660 (N_7660,N_7532,N_7533);
nand U7661 (N_7661,N_7505,N_7554);
nand U7662 (N_7662,N_7504,N_7538);
xnor U7663 (N_7663,N_7553,N_7570);
nor U7664 (N_7664,N_7501,N_7556);
nand U7665 (N_7665,N_7530,N_7524);
or U7666 (N_7666,N_7593,N_7597);
nand U7667 (N_7667,N_7526,N_7571);
nand U7668 (N_7668,N_7539,N_7569);
and U7669 (N_7669,N_7549,N_7583);
nor U7670 (N_7670,N_7519,N_7520);
nor U7671 (N_7671,N_7587,N_7538);
xor U7672 (N_7672,N_7554,N_7596);
nor U7673 (N_7673,N_7512,N_7574);
or U7674 (N_7674,N_7564,N_7549);
xor U7675 (N_7675,N_7593,N_7592);
or U7676 (N_7676,N_7518,N_7598);
nand U7677 (N_7677,N_7544,N_7501);
or U7678 (N_7678,N_7583,N_7534);
nand U7679 (N_7679,N_7500,N_7509);
and U7680 (N_7680,N_7516,N_7504);
nor U7681 (N_7681,N_7569,N_7542);
nand U7682 (N_7682,N_7519,N_7569);
or U7683 (N_7683,N_7574,N_7505);
nor U7684 (N_7684,N_7540,N_7572);
nand U7685 (N_7685,N_7566,N_7595);
xnor U7686 (N_7686,N_7594,N_7579);
and U7687 (N_7687,N_7552,N_7581);
nand U7688 (N_7688,N_7511,N_7579);
or U7689 (N_7689,N_7531,N_7594);
nor U7690 (N_7690,N_7532,N_7524);
or U7691 (N_7691,N_7513,N_7589);
or U7692 (N_7692,N_7575,N_7530);
or U7693 (N_7693,N_7569,N_7501);
nor U7694 (N_7694,N_7576,N_7584);
nand U7695 (N_7695,N_7522,N_7541);
nand U7696 (N_7696,N_7566,N_7538);
nor U7697 (N_7697,N_7589,N_7571);
or U7698 (N_7698,N_7507,N_7546);
or U7699 (N_7699,N_7566,N_7545);
or U7700 (N_7700,N_7689,N_7603);
nand U7701 (N_7701,N_7607,N_7691);
nor U7702 (N_7702,N_7670,N_7602);
xor U7703 (N_7703,N_7652,N_7638);
nand U7704 (N_7704,N_7699,N_7694);
nand U7705 (N_7705,N_7679,N_7614);
and U7706 (N_7706,N_7627,N_7674);
xnor U7707 (N_7707,N_7608,N_7620);
nor U7708 (N_7708,N_7681,N_7676);
or U7709 (N_7709,N_7637,N_7693);
nor U7710 (N_7710,N_7644,N_7671);
nor U7711 (N_7711,N_7660,N_7636);
xor U7712 (N_7712,N_7697,N_7600);
nand U7713 (N_7713,N_7621,N_7605);
nand U7714 (N_7714,N_7624,N_7639);
xor U7715 (N_7715,N_7669,N_7675);
and U7716 (N_7716,N_7649,N_7640);
or U7717 (N_7717,N_7630,N_7686);
and U7718 (N_7718,N_7632,N_7692);
xnor U7719 (N_7719,N_7678,N_7648);
nor U7720 (N_7720,N_7601,N_7612);
and U7721 (N_7721,N_7695,N_7617);
nand U7722 (N_7722,N_7610,N_7604);
xnor U7723 (N_7723,N_7615,N_7667);
nor U7724 (N_7724,N_7655,N_7668);
nand U7725 (N_7725,N_7633,N_7622);
xnor U7726 (N_7726,N_7626,N_7653);
nand U7727 (N_7727,N_7611,N_7651);
or U7728 (N_7728,N_7616,N_7683);
nor U7729 (N_7729,N_7635,N_7663);
xnor U7730 (N_7730,N_7646,N_7677);
nand U7731 (N_7731,N_7665,N_7634);
nand U7732 (N_7732,N_7613,N_7685);
and U7733 (N_7733,N_7698,N_7658);
nand U7734 (N_7734,N_7650,N_7664);
nor U7735 (N_7735,N_7609,N_7645);
nor U7736 (N_7736,N_7631,N_7643);
nand U7737 (N_7737,N_7688,N_7696);
and U7738 (N_7738,N_7642,N_7623);
nand U7739 (N_7739,N_7672,N_7680);
and U7740 (N_7740,N_7656,N_7654);
nor U7741 (N_7741,N_7661,N_7618);
nor U7742 (N_7742,N_7629,N_7659);
xor U7743 (N_7743,N_7666,N_7657);
nand U7744 (N_7744,N_7619,N_7628);
nor U7745 (N_7745,N_7684,N_7647);
or U7746 (N_7746,N_7662,N_7641);
nand U7747 (N_7747,N_7625,N_7682);
xor U7748 (N_7748,N_7687,N_7673);
xnor U7749 (N_7749,N_7606,N_7690);
or U7750 (N_7750,N_7600,N_7667);
nor U7751 (N_7751,N_7685,N_7696);
xnor U7752 (N_7752,N_7618,N_7616);
nor U7753 (N_7753,N_7665,N_7666);
and U7754 (N_7754,N_7627,N_7677);
or U7755 (N_7755,N_7634,N_7620);
nor U7756 (N_7756,N_7646,N_7694);
nor U7757 (N_7757,N_7602,N_7631);
nor U7758 (N_7758,N_7660,N_7686);
xor U7759 (N_7759,N_7681,N_7636);
nand U7760 (N_7760,N_7634,N_7673);
nand U7761 (N_7761,N_7656,N_7634);
nand U7762 (N_7762,N_7688,N_7644);
nand U7763 (N_7763,N_7655,N_7616);
xor U7764 (N_7764,N_7664,N_7634);
nand U7765 (N_7765,N_7683,N_7617);
xor U7766 (N_7766,N_7645,N_7657);
nor U7767 (N_7767,N_7686,N_7645);
nand U7768 (N_7768,N_7687,N_7635);
nor U7769 (N_7769,N_7689,N_7663);
xnor U7770 (N_7770,N_7611,N_7646);
xnor U7771 (N_7771,N_7665,N_7687);
xor U7772 (N_7772,N_7644,N_7664);
or U7773 (N_7773,N_7616,N_7609);
xor U7774 (N_7774,N_7607,N_7612);
xor U7775 (N_7775,N_7685,N_7677);
or U7776 (N_7776,N_7618,N_7615);
nor U7777 (N_7777,N_7677,N_7654);
or U7778 (N_7778,N_7604,N_7612);
and U7779 (N_7779,N_7624,N_7669);
nor U7780 (N_7780,N_7657,N_7617);
xnor U7781 (N_7781,N_7667,N_7617);
nand U7782 (N_7782,N_7620,N_7630);
xor U7783 (N_7783,N_7613,N_7651);
or U7784 (N_7784,N_7674,N_7615);
and U7785 (N_7785,N_7629,N_7619);
nor U7786 (N_7786,N_7608,N_7671);
xnor U7787 (N_7787,N_7666,N_7682);
xnor U7788 (N_7788,N_7695,N_7641);
xnor U7789 (N_7789,N_7687,N_7646);
xnor U7790 (N_7790,N_7644,N_7667);
xnor U7791 (N_7791,N_7612,N_7632);
nor U7792 (N_7792,N_7692,N_7627);
xor U7793 (N_7793,N_7627,N_7668);
or U7794 (N_7794,N_7632,N_7629);
nor U7795 (N_7795,N_7696,N_7690);
nand U7796 (N_7796,N_7638,N_7603);
nand U7797 (N_7797,N_7649,N_7629);
nand U7798 (N_7798,N_7692,N_7658);
nor U7799 (N_7799,N_7653,N_7659);
nand U7800 (N_7800,N_7703,N_7760);
or U7801 (N_7801,N_7717,N_7737);
nor U7802 (N_7802,N_7755,N_7724);
xnor U7803 (N_7803,N_7726,N_7711);
and U7804 (N_7804,N_7767,N_7780);
xnor U7805 (N_7805,N_7746,N_7732);
nand U7806 (N_7806,N_7768,N_7796);
or U7807 (N_7807,N_7781,N_7713);
nand U7808 (N_7808,N_7740,N_7754);
nand U7809 (N_7809,N_7762,N_7734);
and U7810 (N_7810,N_7789,N_7777);
or U7811 (N_7811,N_7775,N_7715);
and U7812 (N_7812,N_7798,N_7778);
nor U7813 (N_7813,N_7774,N_7743);
xnor U7814 (N_7814,N_7779,N_7736);
and U7815 (N_7815,N_7799,N_7741);
xnor U7816 (N_7816,N_7752,N_7757);
nor U7817 (N_7817,N_7719,N_7756);
or U7818 (N_7818,N_7700,N_7764);
or U7819 (N_7819,N_7788,N_7794);
xnor U7820 (N_7820,N_7735,N_7738);
nor U7821 (N_7821,N_7769,N_7776);
and U7822 (N_7822,N_7771,N_7744);
or U7823 (N_7823,N_7716,N_7733);
or U7824 (N_7824,N_7793,N_7772);
or U7825 (N_7825,N_7785,N_7704);
nand U7826 (N_7826,N_7765,N_7723);
xor U7827 (N_7827,N_7795,N_7739);
xor U7828 (N_7828,N_7792,N_7742);
nor U7829 (N_7829,N_7705,N_7725);
xor U7830 (N_7830,N_7731,N_7783);
and U7831 (N_7831,N_7710,N_7728);
xor U7832 (N_7832,N_7787,N_7753);
xnor U7833 (N_7833,N_7718,N_7707);
nor U7834 (N_7834,N_7714,N_7722);
xor U7835 (N_7835,N_7730,N_7750);
nor U7836 (N_7836,N_7763,N_7790);
xor U7837 (N_7837,N_7727,N_7745);
xor U7838 (N_7838,N_7758,N_7751);
nor U7839 (N_7839,N_7702,N_7709);
nand U7840 (N_7840,N_7729,N_7747);
nor U7841 (N_7841,N_7784,N_7759);
and U7842 (N_7842,N_7766,N_7749);
nor U7843 (N_7843,N_7773,N_7748);
xor U7844 (N_7844,N_7701,N_7706);
or U7845 (N_7845,N_7761,N_7782);
or U7846 (N_7846,N_7797,N_7791);
and U7847 (N_7847,N_7770,N_7721);
nor U7848 (N_7848,N_7720,N_7712);
xor U7849 (N_7849,N_7708,N_7786);
nand U7850 (N_7850,N_7780,N_7746);
xnor U7851 (N_7851,N_7701,N_7719);
or U7852 (N_7852,N_7725,N_7726);
nand U7853 (N_7853,N_7786,N_7709);
nor U7854 (N_7854,N_7788,N_7744);
or U7855 (N_7855,N_7704,N_7709);
nand U7856 (N_7856,N_7772,N_7753);
or U7857 (N_7857,N_7775,N_7778);
and U7858 (N_7858,N_7750,N_7745);
nor U7859 (N_7859,N_7749,N_7718);
or U7860 (N_7860,N_7738,N_7792);
nor U7861 (N_7861,N_7728,N_7753);
and U7862 (N_7862,N_7727,N_7704);
nand U7863 (N_7863,N_7770,N_7799);
xor U7864 (N_7864,N_7741,N_7793);
nor U7865 (N_7865,N_7739,N_7725);
and U7866 (N_7866,N_7761,N_7751);
xnor U7867 (N_7867,N_7712,N_7726);
nor U7868 (N_7868,N_7708,N_7790);
or U7869 (N_7869,N_7737,N_7756);
nand U7870 (N_7870,N_7707,N_7725);
nor U7871 (N_7871,N_7774,N_7794);
nand U7872 (N_7872,N_7769,N_7716);
xnor U7873 (N_7873,N_7720,N_7768);
nand U7874 (N_7874,N_7763,N_7744);
nand U7875 (N_7875,N_7713,N_7754);
nand U7876 (N_7876,N_7746,N_7715);
or U7877 (N_7877,N_7718,N_7730);
nand U7878 (N_7878,N_7704,N_7721);
or U7879 (N_7879,N_7747,N_7797);
or U7880 (N_7880,N_7717,N_7775);
nand U7881 (N_7881,N_7738,N_7728);
or U7882 (N_7882,N_7762,N_7758);
nand U7883 (N_7883,N_7712,N_7760);
and U7884 (N_7884,N_7723,N_7747);
nand U7885 (N_7885,N_7716,N_7767);
and U7886 (N_7886,N_7705,N_7772);
nand U7887 (N_7887,N_7707,N_7788);
and U7888 (N_7888,N_7781,N_7747);
xor U7889 (N_7889,N_7758,N_7724);
nand U7890 (N_7890,N_7710,N_7737);
xnor U7891 (N_7891,N_7783,N_7710);
or U7892 (N_7892,N_7708,N_7715);
and U7893 (N_7893,N_7799,N_7765);
or U7894 (N_7894,N_7741,N_7706);
and U7895 (N_7895,N_7751,N_7768);
nand U7896 (N_7896,N_7707,N_7792);
nor U7897 (N_7897,N_7794,N_7767);
xnor U7898 (N_7898,N_7744,N_7707);
and U7899 (N_7899,N_7735,N_7723);
nand U7900 (N_7900,N_7850,N_7843);
nand U7901 (N_7901,N_7823,N_7819);
and U7902 (N_7902,N_7855,N_7835);
nand U7903 (N_7903,N_7879,N_7874);
or U7904 (N_7904,N_7813,N_7889);
xnor U7905 (N_7905,N_7882,N_7804);
nor U7906 (N_7906,N_7801,N_7807);
nor U7907 (N_7907,N_7837,N_7890);
xnor U7908 (N_7908,N_7824,N_7853);
xor U7909 (N_7909,N_7846,N_7836);
nand U7910 (N_7910,N_7832,N_7815);
or U7911 (N_7911,N_7886,N_7854);
and U7912 (N_7912,N_7896,N_7861);
nor U7913 (N_7913,N_7873,N_7869);
xor U7914 (N_7914,N_7857,N_7872);
or U7915 (N_7915,N_7851,N_7885);
xor U7916 (N_7916,N_7898,N_7814);
and U7917 (N_7917,N_7867,N_7820);
and U7918 (N_7918,N_7810,N_7821);
or U7919 (N_7919,N_7870,N_7827);
and U7920 (N_7920,N_7839,N_7860);
or U7921 (N_7921,N_7842,N_7863);
and U7922 (N_7922,N_7871,N_7856);
nor U7923 (N_7923,N_7877,N_7894);
xnor U7924 (N_7924,N_7805,N_7876);
and U7925 (N_7925,N_7822,N_7800);
nor U7926 (N_7926,N_7875,N_7816);
and U7927 (N_7927,N_7868,N_7808);
xor U7928 (N_7928,N_7849,N_7852);
and U7929 (N_7929,N_7859,N_7881);
or U7930 (N_7930,N_7847,N_7840);
and U7931 (N_7931,N_7884,N_7834);
and U7932 (N_7932,N_7812,N_7865);
or U7933 (N_7933,N_7888,N_7893);
nor U7934 (N_7934,N_7817,N_7895);
or U7935 (N_7935,N_7864,N_7845);
nand U7936 (N_7936,N_7887,N_7878);
xor U7937 (N_7937,N_7848,N_7802);
and U7938 (N_7938,N_7803,N_7826);
and U7939 (N_7939,N_7833,N_7811);
nor U7940 (N_7940,N_7866,N_7862);
xnor U7941 (N_7941,N_7830,N_7829);
xor U7942 (N_7942,N_7825,N_7818);
xor U7943 (N_7943,N_7831,N_7838);
nand U7944 (N_7944,N_7899,N_7892);
and U7945 (N_7945,N_7809,N_7844);
xor U7946 (N_7946,N_7880,N_7858);
or U7947 (N_7947,N_7806,N_7897);
or U7948 (N_7948,N_7883,N_7841);
nor U7949 (N_7949,N_7891,N_7828);
and U7950 (N_7950,N_7817,N_7821);
nor U7951 (N_7951,N_7828,N_7805);
or U7952 (N_7952,N_7880,N_7852);
or U7953 (N_7953,N_7887,N_7813);
nor U7954 (N_7954,N_7871,N_7860);
nand U7955 (N_7955,N_7866,N_7817);
or U7956 (N_7956,N_7876,N_7880);
or U7957 (N_7957,N_7868,N_7809);
and U7958 (N_7958,N_7811,N_7874);
nor U7959 (N_7959,N_7832,N_7860);
nand U7960 (N_7960,N_7808,N_7877);
and U7961 (N_7961,N_7893,N_7859);
or U7962 (N_7962,N_7850,N_7871);
xnor U7963 (N_7963,N_7869,N_7887);
nor U7964 (N_7964,N_7808,N_7854);
and U7965 (N_7965,N_7893,N_7802);
or U7966 (N_7966,N_7898,N_7862);
nor U7967 (N_7967,N_7860,N_7896);
or U7968 (N_7968,N_7816,N_7829);
nand U7969 (N_7969,N_7819,N_7816);
or U7970 (N_7970,N_7856,N_7849);
xor U7971 (N_7971,N_7837,N_7820);
and U7972 (N_7972,N_7873,N_7861);
or U7973 (N_7973,N_7821,N_7847);
and U7974 (N_7974,N_7808,N_7881);
nand U7975 (N_7975,N_7884,N_7829);
nand U7976 (N_7976,N_7833,N_7881);
nand U7977 (N_7977,N_7883,N_7848);
nor U7978 (N_7978,N_7818,N_7853);
nand U7979 (N_7979,N_7814,N_7842);
and U7980 (N_7980,N_7834,N_7871);
nor U7981 (N_7981,N_7865,N_7826);
or U7982 (N_7982,N_7821,N_7871);
or U7983 (N_7983,N_7899,N_7895);
xnor U7984 (N_7984,N_7835,N_7850);
and U7985 (N_7985,N_7822,N_7842);
and U7986 (N_7986,N_7867,N_7844);
or U7987 (N_7987,N_7825,N_7855);
nor U7988 (N_7988,N_7817,N_7802);
and U7989 (N_7989,N_7809,N_7885);
nand U7990 (N_7990,N_7833,N_7817);
or U7991 (N_7991,N_7808,N_7827);
nand U7992 (N_7992,N_7807,N_7829);
nor U7993 (N_7993,N_7825,N_7800);
nor U7994 (N_7994,N_7813,N_7848);
xor U7995 (N_7995,N_7881,N_7847);
and U7996 (N_7996,N_7835,N_7874);
and U7997 (N_7997,N_7832,N_7859);
and U7998 (N_7998,N_7846,N_7819);
nand U7999 (N_7999,N_7825,N_7843);
or U8000 (N_8000,N_7984,N_7951);
xor U8001 (N_8001,N_7995,N_7987);
and U8002 (N_8002,N_7961,N_7981);
and U8003 (N_8003,N_7982,N_7923);
and U8004 (N_8004,N_7915,N_7999);
nand U8005 (N_8005,N_7932,N_7996);
xnor U8006 (N_8006,N_7994,N_7957);
and U8007 (N_8007,N_7969,N_7988);
or U8008 (N_8008,N_7983,N_7971);
nand U8009 (N_8009,N_7935,N_7960);
or U8010 (N_8010,N_7955,N_7940);
nor U8011 (N_8011,N_7922,N_7916);
or U8012 (N_8012,N_7975,N_7904);
and U8013 (N_8013,N_7978,N_7934);
and U8014 (N_8014,N_7917,N_7977);
or U8015 (N_8015,N_7964,N_7924);
xor U8016 (N_8016,N_7950,N_7998);
and U8017 (N_8017,N_7930,N_7945);
or U8018 (N_8018,N_7905,N_7985);
or U8019 (N_8019,N_7929,N_7900);
xnor U8020 (N_8020,N_7979,N_7910);
xnor U8021 (N_8021,N_7967,N_7942);
or U8022 (N_8022,N_7933,N_7909);
and U8023 (N_8023,N_7963,N_7954);
nand U8024 (N_8024,N_7901,N_7938);
nor U8025 (N_8025,N_7958,N_7939);
or U8026 (N_8026,N_7913,N_7956);
nand U8027 (N_8027,N_7966,N_7902);
nor U8028 (N_8028,N_7931,N_7919);
nand U8029 (N_8029,N_7944,N_7949);
or U8030 (N_8030,N_7946,N_7903);
nand U8031 (N_8031,N_7928,N_7906);
nor U8032 (N_8032,N_7908,N_7997);
nor U8033 (N_8033,N_7947,N_7918);
nor U8034 (N_8034,N_7948,N_7992);
xnor U8035 (N_8035,N_7986,N_7941);
nand U8036 (N_8036,N_7937,N_7980);
nor U8037 (N_8037,N_7914,N_7926);
xnor U8038 (N_8038,N_7953,N_7952);
xor U8039 (N_8039,N_7920,N_7976);
xor U8040 (N_8040,N_7991,N_7907);
or U8041 (N_8041,N_7936,N_7921);
or U8042 (N_8042,N_7965,N_7973);
and U8043 (N_8043,N_7968,N_7974);
xor U8044 (N_8044,N_7970,N_7925);
nor U8045 (N_8045,N_7912,N_7993);
and U8046 (N_8046,N_7927,N_7962);
xor U8047 (N_8047,N_7959,N_7972);
nor U8048 (N_8048,N_7989,N_7911);
nand U8049 (N_8049,N_7943,N_7990);
or U8050 (N_8050,N_7905,N_7973);
nand U8051 (N_8051,N_7930,N_7947);
or U8052 (N_8052,N_7995,N_7964);
or U8053 (N_8053,N_7969,N_7959);
xnor U8054 (N_8054,N_7990,N_7954);
xor U8055 (N_8055,N_7999,N_7939);
xor U8056 (N_8056,N_7978,N_7969);
xnor U8057 (N_8057,N_7936,N_7979);
and U8058 (N_8058,N_7921,N_7906);
xor U8059 (N_8059,N_7933,N_7995);
nand U8060 (N_8060,N_7944,N_7919);
nor U8061 (N_8061,N_7974,N_7946);
xor U8062 (N_8062,N_7909,N_7953);
nand U8063 (N_8063,N_7937,N_7993);
nor U8064 (N_8064,N_7903,N_7980);
nor U8065 (N_8065,N_7907,N_7938);
nand U8066 (N_8066,N_7982,N_7935);
and U8067 (N_8067,N_7912,N_7937);
nand U8068 (N_8068,N_7998,N_7909);
nand U8069 (N_8069,N_7920,N_7994);
and U8070 (N_8070,N_7914,N_7907);
nand U8071 (N_8071,N_7947,N_7960);
nand U8072 (N_8072,N_7992,N_7940);
and U8073 (N_8073,N_7989,N_7983);
nor U8074 (N_8074,N_7993,N_7932);
and U8075 (N_8075,N_7973,N_7960);
and U8076 (N_8076,N_7990,N_7950);
nor U8077 (N_8077,N_7961,N_7926);
nand U8078 (N_8078,N_7993,N_7967);
nand U8079 (N_8079,N_7956,N_7947);
or U8080 (N_8080,N_7996,N_7981);
nand U8081 (N_8081,N_7969,N_7901);
and U8082 (N_8082,N_7961,N_7904);
xor U8083 (N_8083,N_7982,N_7947);
or U8084 (N_8084,N_7989,N_7994);
or U8085 (N_8085,N_7941,N_7939);
nor U8086 (N_8086,N_7904,N_7994);
nor U8087 (N_8087,N_7988,N_7948);
nor U8088 (N_8088,N_7928,N_7903);
nor U8089 (N_8089,N_7908,N_7943);
nor U8090 (N_8090,N_7995,N_7953);
nand U8091 (N_8091,N_7944,N_7926);
nand U8092 (N_8092,N_7967,N_7963);
nor U8093 (N_8093,N_7903,N_7912);
nor U8094 (N_8094,N_7909,N_7950);
or U8095 (N_8095,N_7955,N_7966);
and U8096 (N_8096,N_7986,N_7927);
nor U8097 (N_8097,N_7945,N_7969);
nor U8098 (N_8098,N_7990,N_7983);
or U8099 (N_8099,N_7979,N_7952);
and U8100 (N_8100,N_8014,N_8024);
or U8101 (N_8101,N_8055,N_8008);
and U8102 (N_8102,N_8079,N_8089);
xnor U8103 (N_8103,N_8078,N_8092);
xnor U8104 (N_8104,N_8074,N_8041);
and U8105 (N_8105,N_8060,N_8042);
nor U8106 (N_8106,N_8009,N_8017);
nand U8107 (N_8107,N_8066,N_8071);
or U8108 (N_8108,N_8002,N_8007);
nor U8109 (N_8109,N_8084,N_8077);
or U8110 (N_8110,N_8062,N_8052);
nor U8111 (N_8111,N_8083,N_8019);
or U8112 (N_8112,N_8094,N_8044);
and U8113 (N_8113,N_8098,N_8049);
and U8114 (N_8114,N_8095,N_8030);
xor U8115 (N_8115,N_8099,N_8093);
nor U8116 (N_8116,N_8018,N_8068);
nand U8117 (N_8117,N_8040,N_8022);
nand U8118 (N_8118,N_8067,N_8065);
and U8119 (N_8119,N_8006,N_8064);
nand U8120 (N_8120,N_8043,N_8063);
xor U8121 (N_8121,N_8028,N_8073);
nor U8122 (N_8122,N_8037,N_8059);
xor U8123 (N_8123,N_8096,N_8003);
or U8124 (N_8124,N_8023,N_8012);
and U8125 (N_8125,N_8004,N_8038);
and U8126 (N_8126,N_8045,N_8082);
nor U8127 (N_8127,N_8031,N_8035);
nand U8128 (N_8128,N_8054,N_8032);
and U8129 (N_8129,N_8046,N_8025);
nand U8130 (N_8130,N_8086,N_8021);
xnor U8131 (N_8131,N_8061,N_8050);
nor U8132 (N_8132,N_8034,N_8001);
nor U8133 (N_8133,N_8051,N_8057);
xor U8134 (N_8134,N_8070,N_8020);
nor U8135 (N_8135,N_8072,N_8005);
and U8136 (N_8136,N_8026,N_8058);
nor U8137 (N_8137,N_8033,N_8013);
nand U8138 (N_8138,N_8027,N_8010);
or U8139 (N_8139,N_8076,N_8069);
nand U8140 (N_8140,N_8048,N_8097);
xor U8141 (N_8141,N_8056,N_8085);
nor U8142 (N_8142,N_8000,N_8080);
xnor U8143 (N_8143,N_8036,N_8081);
or U8144 (N_8144,N_8088,N_8039);
xor U8145 (N_8145,N_8091,N_8053);
xnor U8146 (N_8146,N_8011,N_8075);
and U8147 (N_8147,N_8016,N_8047);
nand U8148 (N_8148,N_8090,N_8015);
nor U8149 (N_8149,N_8087,N_8029);
nand U8150 (N_8150,N_8033,N_8017);
or U8151 (N_8151,N_8008,N_8044);
nand U8152 (N_8152,N_8001,N_8084);
or U8153 (N_8153,N_8073,N_8032);
xor U8154 (N_8154,N_8071,N_8090);
and U8155 (N_8155,N_8049,N_8070);
or U8156 (N_8156,N_8042,N_8067);
xor U8157 (N_8157,N_8049,N_8095);
xnor U8158 (N_8158,N_8087,N_8050);
nand U8159 (N_8159,N_8029,N_8013);
and U8160 (N_8160,N_8007,N_8025);
or U8161 (N_8161,N_8059,N_8091);
and U8162 (N_8162,N_8059,N_8042);
or U8163 (N_8163,N_8088,N_8026);
xor U8164 (N_8164,N_8025,N_8019);
or U8165 (N_8165,N_8056,N_8090);
and U8166 (N_8166,N_8078,N_8093);
xnor U8167 (N_8167,N_8008,N_8084);
nor U8168 (N_8168,N_8058,N_8031);
nor U8169 (N_8169,N_8021,N_8067);
nor U8170 (N_8170,N_8047,N_8042);
nor U8171 (N_8171,N_8048,N_8043);
and U8172 (N_8172,N_8009,N_8025);
nand U8173 (N_8173,N_8056,N_8068);
xor U8174 (N_8174,N_8038,N_8049);
nor U8175 (N_8175,N_8029,N_8005);
nand U8176 (N_8176,N_8009,N_8024);
nor U8177 (N_8177,N_8054,N_8079);
xnor U8178 (N_8178,N_8082,N_8064);
xor U8179 (N_8179,N_8010,N_8082);
or U8180 (N_8180,N_8031,N_8056);
nand U8181 (N_8181,N_8095,N_8077);
or U8182 (N_8182,N_8027,N_8045);
nand U8183 (N_8183,N_8028,N_8020);
or U8184 (N_8184,N_8022,N_8032);
or U8185 (N_8185,N_8013,N_8022);
nand U8186 (N_8186,N_8039,N_8064);
nand U8187 (N_8187,N_8018,N_8067);
nand U8188 (N_8188,N_8081,N_8099);
xor U8189 (N_8189,N_8017,N_8057);
xnor U8190 (N_8190,N_8051,N_8077);
and U8191 (N_8191,N_8070,N_8097);
xor U8192 (N_8192,N_8092,N_8010);
nor U8193 (N_8193,N_8076,N_8072);
nand U8194 (N_8194,N_8049,N_8085);
or U8195 (N_8195,N_8012,N_8003);
or U8196 (N_8196,N_8052,N_8040);
xor U8197 (N_8197,N_8038,N_8028);
and U8198 (N_8198,N_8049,N_8066);
and U8199 (N_8199,N_8079,N_8010);
nor U8200 (N_8200,N_8176,N_8146);
xor U8201 (N_8201,N_8183,N_8150);
nand U8202 (N_8202,N_8194,N_8141);
nor U8203 (N_8203,N_8144,N_8139);
nor U8204 (N_8204,N_8197,N_8182);
or U8205 (N_8205,N_8126,N_8192);
nand U8206 (N_8206,N_8187,N_8105);
and U8207 (N_8207,N_8188,N_8104);
xnor U8208 (N_8208,N_8158,N_8123);
nand U8209 (N_8209,N_8125,N_8112);
xor U8210 (N_8210,N_8173,N_8100);
xnor U8211 (N_8211,N_8122,N_8151);
or U8212 (N_8212,N_8138,N_8175);
xor U8213 (N_8213,N_8142,N_8172);
nand U8214 (N_8214,N_8109,N_8124);
nand U8215 (N_8215,N_8143,N_8190);
and U8216 (N_8216,N_8106,N_8116);
and U8217 (N_8217,N_8119,N_8169);
nor U8218 (N_8218,N_8107,N_8103);
xor U8219 (N_8219,N_8121,N_8185);
or U8220 (N_8220,N_8156,N_8131);
nand U8221 (N_8221,N_8136,N_8181);
nand U8222 (N_8222,N_8117,N_8167);
xor U8223 (N_8223,N_8159,N_8163);
nand U8224 (N_8224,N_8134,N_8184);
and U8225 (N_8225,N_8128,N_8174);
xor U8226 (N_8226,N_8129,N_8199);
nand U8227 (N_8227,N_8154,N_8118);
or U8228 (N_8228,N_8108,N_8157);
nor U8229 (N_8229,N_8102,N_8115);
xor U8230 (N_8230,N_8149,N_8198);
xnor U8231 (N_8231,N_8152,N_8148);
xnor U8232 (N_8232,N_8120,N_8164);
nor U8233 (N_8233,N_8110,N_8196);
or U8234 (N_8234,N_8101,N_8127);
nor U8235 (N_8235,N_8168,N_8114);
or U8236 (N_8236,N_8113,N_8147);
nor U8237 (N_8237,N_8153,N_8135);
nand U8238 (N_8238,N_8160,N_8165);
nand U8239 (N_8239,N_8166,N_8140);
and U8240 (N_8240,N_8133,N_8179);
xnor U8241 (N_8241,N_8186,N_8170);
nand U8242 (N_8242,N_8193,N_8137);
nand U8243 (N_8243,N_8111,N_8130);
and U8244 (N_8244,N_8180,N_8132);
xor U8245 (N_8245,N_8161,N_8145);
nand U8246 (N_8246,N_8155,N_8191);
and U8247 (N_8247,N_8162,N_8178);
xor U8248 (N_8248,N_8177,N_8171);
or U8249 (N_8249,N_8195,N_8189);
nand U8250 (N_8250,N_8124,N_8100);
nor U8251 (N_8251,N_8151,N_8199);
and U8252 (N_8252,N_8186,N_8108);
xnor U8253 (N_8253,N_8140,N_8186);
xor U8254 (N_8254,N_8157,N_8145);
xor U8255 (N_8255,N_8150,N_8105);
xnor U8256 (N_8256,N_8166,N_8133);
nor U8257 (N_8257,N_8186,N_8191);
or U8258 (N_8258,N_8146,N_8122);
and U8259 (N_8259,N_8137,N_8171);
xor U8260 (N_8260,N_8128,N_8150);
xnor U8261 (N_8261,N_8180,N_8149);
or U8262 (N_8262,N_8181,N_8172);
or U8263 (N_8263,N_8149,N_8143);
or U8264 (N_8264,N_8112,N_8174);
nand U8265 (N_8265,N_8150,N_8124);
nand U8266 (N_8266,N_8104,N_8180);
or U8267 (N_8267,N_8195,N_8171);
nand U8268 (N_8268,N_8163,N_8114);
xor U8269 (N_8269,N_8191,N_8165);
xnor U8270 (N_8270,N_8156,N_8114);
and U8271 (N_8271,N_8182,N_8154);
nand U8272 (N_8272,N_8182,N_8157);
nand U8273 (N_8273,N_8122,N_8169);
xnor U8274 (N_8274,N_8155,N_8152);
or U8275 (N_8275,N_8187,N_8184);
nand U8276 (N_8276,N_8127,N_8104);
xnor U8277 (N_8277,N_8151,N_8126);
or U8278 (N_8278,N_8104,N_8184);
and U8279 (N_8279,N_8110,N_8112);
nand U8280 (N_8280,N_8107,N_8187);
xnor U8281 (N_8281,N_8115,N_8148);
or U8282 (N_8282,N_8152,N_8193);
and U8283 (N_8283,N_8144,N_8187);
and U8284 (N_8284,N_8146,N_8152);
nand U8285 (N_8285,N_8185,N_8167);
nand U8286 (N_8286,N_8164,N_8135);
nor U8287 (N_8287,N_8118,N_8171);
nand U8288 (N_8288,N_8120,N_8176);
nor U8289 (N_8289,N_8122,N_8195);
xor U8290 (N_8290,N_8134,N_8144);
and U8291 (N_8291,N_8118,N_8157);
and U8292 (N_8292,N_8161,N_8126);
nor U8293 (N_8293,N_8192,N_8119);
and U8294 (N_8294,N_8115,N_8157);
or U8295 (N_8295,N_8150,N_8193);
nand U8296 (N_8296,N_8122,N_8106);
and U8297 (N_8297,N_8149,N_8158);
nor U8298 (N_8298,N_8107,N_8182);
nor U8299 (N_8299,N_8160,N_8149);
or U8300 (N_8300,N_8256,N_8260);
or U8301 (N_8301,N_8210,N_8275);
xor U8302 (N_8302,N_8270,N_8265);
or U8303 (N_8303,N_8282,N_8208);
and U8304 (N_8304,N_8225,N_8230);
nand U8305 (N_8305,N_8204,N_8262);
nor U8306 (N_8306,N_8207,N_8279);
or U8307 (N_8307,N_8232,N_8287);
nand U8308 (N_8308,N_8242,N_8272);
or U8309 (N_8309,N_8258,N_8257);
and U8310 (N_8310,N_8268,N_8226);
or U8311 (N_8311,N_8290,N_8201);
and U8312 (N_8312,N_8278,N_8292);
or U8313 (N_8313,N_8216,N_8212);
nand U8314 (N_8314,N_8266,N_8296);
or U8315 (N_8315,N_8238,N_8246);
nor U8316 (N_8316,N_8217,N_8222);
xor U8317 (N_8317,N_8248,N_8285);
nand U8318 (N_8318,N_8289,N_8298);
or U8319 (N_8319,N_8293,N_8228);
and U8320 (N_8320,N_8281,N_8218);
nor U8321 (N_8321,N_8202,N_8271);
nor U8322 (N_8322,N_8229,N_8273);
or U8323 (N_8323,N_8243,N_8236);
or U8324 (N_8324,N_8255,N_8252);
nand U8325 (N_8325,N_8263,N_8239);
or U8326 (N_8326,N_8237,N_8245);
and U8327 (N_8327,N_8288,N_8205);
or U8328 (N_8328,N_8284,N_8264);
nor U8329 (N_8329,N_8240,N_8251);
nand U8330 (N_8330,N_8261,N_8291);
nand U8331 (N_8331,N_8277,N_8294);
or U8332 (N_8332,N_8220,N_8241);
or U8333 (N_8333,N_8254,N_8213);
nand U8334 (N_8334,N_8219,N_8249);
nand U8335 (N_8335,N_8247,N_8215);
and U8336 (N_8336,N_8244,N_8269);
nor U8337 (N_8337,N_8214,N_8200);
xor U8338 (N_8338,N_8259,N_8280);
and U8339 (N_8339,N_8253,N_8276);
nor U8340 (N_8340,N_8299,N_8295);
or U8341 (N_8341,N_8274,N_8231);
and U8342 (N_8342,N_8283,N_8209);
nand U8343 (N_8343,N_8206,N_8234);
nand U8344 (N_8344,N_8221,N_8233);
nor U8345 (N_8345,N_8203,N_8250);
and U8346 (N_8346,N_8211,N_8224);
nor U8347 (N_8347,N_8297,N_8267);
or U8348 (N_8348,N_8286,N_8223);
and U8349 (N_8349,N_8227,N_8235);
and U8350 (N_8350,N_8268,N_8280);
or U8351 (N_8351,N_8286,N_8258);
nor U8352 (N_8352,N_8270,N_8283);
nor U8353 (N_8353,N_8277,N_8206);
nand U8354 (N_8354,N_8299,N_8213);
and U8355 (N_8355,N_8286,N_8230);
nor U8356 (N_8356,N_8272,N_8233);
xor U8357 (N_8357,N_8227,N_8236);
nand U8358 (N_8358,N_8288,N_8220);
nand U8359 (N_8359,N_8224,N_8216);
nand U8360 (N_8360,N_8268,N_8295);
or U8361 (N_8361,N_8250,N_8255);
xnor U8362 (N_8362,N_8211,N_8297);
xor U8363 (N_8363,N_8262,N_8299);
xor U8364 (N_8364,N_8208,N_8250);
nor U8365 (N_8365,N_8269,N_8259);
nor U8366 (N_8366,N_8258,N_8223);
xnor U8367 (N_8367,N_8250,N_8239);
nor U8368 (N_8368,N_8295,N_8212);
nor U8369 (N_8369,N_8251,N_8207);
xor U8370 (N_8370,N_8256,N_8224);
or U8371 (N_8371,N_8205,N_8200);
nand U8372 (N_8372,N_8253,N_8251);
nand U8373 (N_8373,N_8284,N_8296);
nor U8374 (N_8374,N_8230,N_8224);
and U8375 (N_8375,N_8290,N_8231);
nand U8376 (N_8376,N_8292,N_8207);
nor U8377 (N_8377,N_8255,N_8284);
nor U8378 (N_8378,N_8270,N_8282);
nor U8379 (N_8379,N_8204,N_8275);
xor U8380 (N_8380,N_8273,N_8235);
or U8381 (N_8381,N_8211,N_8280);
xor U8382 (N_8382,N_8213,N_8241);
nor U8383 (N_8383,N_8261,N_8274);
nand U8384 (N_8384,N_8269,N_8292);
or U8385 (N_8385,N_8202,N_8278);
or U8386 (N_8386,N_8258,N_8259);
xnor U8387 (N_8387,N_8276,N_8234);
nand U8388 (N_8388,N_8214,N_8270);
nand U8389 (N_8389,N_8254,N_8231);
and U8390 (N_8390,N_8292,N_8232);
or U8391 (N_8391,N_8293,N_8246);
xor U8392 (N_8392,N_8232,N_8226);
nor U8393 (N_8393,N_8264,N_8239);
xnor U8394 (N_8394,N_8252,N_8222);
or U8395 (N_8395,N_8205,N_8298);
and U8396 (N_8396,N_8255,N_8296);
or U8397 (N_8397,N_8284,N_8261);
nand U8398 (N_8398,N_8246,N_8242);
and U8399 (N_8399,N_8229,N_8295);
nand U8400 (N_8400,N_8361,N_8344);
or U8401 (N_8401,N_8360,N_8356);
and U8402 (N_8402,N_8366,N_8367);
nand U8403 (N_8403,N_8315,N_8321);
or U8404 (N_8404,N_8300,N_8376);
and U8405 (N_8405,N_8357,N_8341);
and U8406 (N_8406,N_8369,N_8354);
nand U8407 (N_8407,N_8302,N_8373);
nand U8408 (N_8408,N_8333,N_8345);
and U8409 (N_8409,N_8313,N_8337);
xor U8410 (N_8410,N_8370,N_8378);
and U8411 (N_8411,N_8314,N_8355);
nor U8412 (N_8412,N_8359,N_8377);
nand U8413 (N_8413,N_8322,N_8385);
and U8414 (N_8414,N_8349,N_8303);
and U8415 (N_8415,N_8365,N_8346);
or U8416 (N_8416,N_8340,N_8375);
xor U8417 (N_8417,N_8325,N_8393);
and U8418 (N_8418,N_8396,N_8362);
xnor U8419 (N_8419,N_8309,N_8311);
nor U8420 (N_8420,N_8352,N_8331);
xor U8421 (N_8421,N_8374,N_8308);
and U8422 (N_8422,N_8388,N_8343);
nor U8423 (N_8423,N_8364,N_8394);
nand U8424 (N_8424,N_8312,N_8381);
nand U8425 (N_8425,N_8330,N_8327);
xor U8426 (N_8426,N_8324,N_8336);
nor U8427 (N_8427,N_8307,N_8391);
nor U8428 (N_8428,N_8338,N_8323);
nand U8429 (N_8429,N_8363,N_8319);
and U8430 (N_8430,N_8353,N_8329);
nand U8431 (N_8431,N_8348,N_8326);
nor U8432 (N_8432,N_8335,N_8328);
nand U8433 (N_8433,N_8383,N_8358);
or U8434 (N_8434,N_8390,N_8304);
or U8435 (N_8435,N_8395,N_8379);
nor U8436 (N_8436,N_8306,N_8372);
xor U8437 (N_8437,N_8310,N_8318);
nand U8438 (N_8438,N_8380,N_8386);
xor U8439 (N_8439,N_8317,N_8320);
xor U8440 (N_8440,N_8387,N_8392);
xnor U8441 (N_8441,N_8305,N_8301);
xor U8442 (N_8442,N_8339,N_8397);
and U8443 (N_8443,N_8350,N_8382);
xnor U8444 (N_8444,N_8351,N_8368);
nand U8445 (N_8445,N_8342,N_8389);
xor U8446 (N_8446,N_8398,N_8316);
or U8447 (N_8447,N_8384,N_8399);
nor U8448 (N_8448,N_8371,N_8334);
nand U8449 (N_8449,N_8347,N_8332);
and U8450 (N_8450,N_8342,N_8367);
or U8451 (N_8451,N_8335,N_8303);
nand U8452 (N_8452,N_8303,N_8330);
nand U8453 (N_8453,N_8375,N_8334);
and U8454 (N_8454,N_8365,N_8352);
and U8455 (N_8455,N_8320,N_8395);
and U8456 (N_8456,N_8353,N_8390);
or U8457 (N_8457,N_8374,N_8301);
or U8458 (N_8458,N_8330,N_8334);
xnor U8459 (N_8459,N_8337,N_8399);
nor U8460 (N_8460,N_8364,N_8361);
nor U8461 (N_8461,N_8311,N_8321);
and U8462 (N_8462,N_8361,N_8329);
xnor U8463 (N_8463,N_8358,N_8335);
nand U8464 (N_8464,N_8308,N_8388);
or U8465 (N_8465,N_8359,N_8347);
nand U8466 (N_8466,N_8304,N_8351);
nor U8467 (N_8467,N_8353,N_8302);
nand U8468 (N_8468,N_8344,N_8346);
or U8469 (N_8469,N_8315,N_8318);
xnor U8470 (N_8470,N_8372,N_8340);
xnor U8471 (N_8471,N_8312,N_8375);
or U8472 (N_8472,N_8347,N_8397);
or U8473 (N_8473,N_8315,N_8371);
nor U8474 (N_8474,N_8335,N_8321);
nor U8475 (N_8475,N_8327,N_8387);
xor U8476 (N_8476,N_8312,N_8377);
and U8477 (N_8477,N_8357,N_8353);
or U8478 (N_8478,N_8318,N_8332);
xnor U8479 (N_8479,N_8378,N_8360);
or U8480 (N_8480,N_8376,N_8394);
xnor U8481 (N_8481,N_8339,N_8313);
and U8482 (N_8482,N_8368,N_8309);
xnor U8483 (N_8483,N_8354,N_8308);
or U8484 (N_8484,N_8384,N_8387);
or U8485 (N_8485,N_8329,N_8356);
nor U8486 (N_8486,N_8387,N_8314);
or U8487 (N_8487,N_8327,N_8313);
nor U8488 (N_8488,N_8318,N_8312);
and U8489 (N_8489,N_8392,N_8349);
or U8490 (N_8490,N_8390,N_8308);
or U8491 (N_8491,N_8376,N_8381);
xor U8492 (N_8492,N_8394,N_8362);
nand U8493 (N_8493,N_8377,N_8392);
nor U8494 (N_8494,N_8318,N_8328);
or U8495 (N_8495,N_8386,N_8304);
and U8496 (N_8496,N_8330,N_8319);
nand U8497 (N_8497,N_8366,N_8338);
nand U8498 (N_8498,N_8389,N_8307);
or U8499 (N_8499,N_8333,N_8381);
and U8500 (N_8500,N_8455,N_8457);
nor U8501 (N_8501,N_8490,N_8409);
nor U8502 (N_8502,N_8492,N_8414);
xnor U8503 (N_8503,N_8450,N_8444);
nor U8504 (N_8504,N_8491,N_8440);
nor U8505 (N_8505,N_8443,N_8415);
or U8506 (N_8506,N_8405,N_8448);
nand U8507 (N_8507,N_8449,N_8463);
xnor U8508 (N_8508,N_8434,N_8432);
nor U8509 (N_8509,N_8471,N_8493);
xor U8510 (N_8510,N_8404,N_8413);
and U8511 (N_8511,N_8456,N_8467);
nand U8512 (N_8512,N_8464,N_8478);
xor U8513 (N_8513,N_8480,N_8441);
or U8514 (N_8514,N_8459,N_8427);
and U8515 (N_8515,N_8424,N_8474);
nand U8516 (N_8516,N_8458,N_8412);
or U8517 (N_8517,N_8472,N_8494);
and U8518 (N_8518,N_8421,N_8416);
and U8519 (N_8519,N_8436,N_8439);
or U8520 (N_8520,N_8431,N_8429);
xor U8521 (N_8521,N_8497,N_8406);
xnor U8522 (N_8522,N_8447,N_8408);
or U8523 (N_8523,N_8461,N_8473);
xnor U8524 (N_8524,N_8479,N_8453);
or U8525 (N_8525,N_8430,N_8410);
nor U8526 (N_8526,N_8435,N_8454);
and U8527 (N_8527,N_8411,N_8482);
nor U8528 (N_8528,N_8483,N_8451);
nand U8529 (N_8529,N_8452,N_8446);
and U8530 (N_8530,N_8420,N_8442);
and U8531 (N_8531,N_8469,N_8489);
or U8532 (N_8532,N_8428,N_8426);
nor U8533 (N_8533,N_8407,N_8486);
nor U8534 (N_8534,N_8476,N_8438);
nand U8535 (N_8535,N_8496,N_8462);
xnor U8536 (N_8536,N_8466,N_8419);
nor U8537 (N_8537,N_8495,N_8460);
and U8538 (N_8538,N_8418,N_8481);
xnor U8539 (N_8539,N_8401,N_8468);
nand U8540 (N_8540,N_8433,N_8475);
and U8541 (N_8541,N_8498,N_8417);
and U8542 (N_8542,N_8488,N_8423);
nand U8543 (N_8543,N_8400,N_8484);
nor U8544 (N_8544,N_8499,N_8422);
nand U8545 (N_8545,N_8470,N_8487);
or U8546 (N_8546,N_8403,N_8465);
nand U8547 (N_8547,N_8425,N_8477);
and U8548 (N_8548,N_8437,N_8445);
and U8549 (N_8549,N_8485,N_8402);
nand U8550 (N_8550,N_8430,N_8403);
xor U8551 (N_8551,N_8485,N_8419);
nor U8552 (N_8552,N_8495,N_8415);
xor U8553 (N_8553,N_8422,N_8412);
and U8554 (N_8554,N_8446,N_8488);
nor U8555 (N_8555,N_8425,N_8428);
xor U8556 (N_8556,N_8411,N_8498);
nand U8557 (N_8557,N_8486,N_8481);
or U8558 (N_8558,N_8445,N_8420);
nor U8559 (N_8559,N_8469,N_8464);
xnor U8560 (N_8560,N_8490,N_8435);
nand U8561 (N_8561,N_8431,N_8434);
xnor U8562 (N_8562,N_8438,N_8416);
nand U8563 (N_8563,N_8402,N_8427);
nor U8564 (N_8564,N_8492,N_8451);
nor U8565 (N_8565,N_8445,N_8414);
nor U8566 (N_8566,N_8422,N_8426);
or U8567 (N_8567,N_8490,N_8482);
nor U8568 (N_8568,N_8462,N_8463);
and U8569 (N_8569,N_8423,N_8483);
and U8570 (N_8570,N_8475,N_8497);
or U8571 (N_8571,N_8434,N_8459);
and U8572 (N_8572,N_8425,N_8414);
xnor U8573 (N_8573,N_8474,N_8411);
xnor U8574 (N_8574,N_8477,N_8427);
or U8575 (N_8575,N_8473,N_8402);
and U8576 (N_8576,N_8405,N_8444);
or U8577 (N_8577,N_8465,N_8407);
nor U8578 (N_8578,N_8401,N_8414);
nor U8579 (N_8579,N_8429,N_8493);
and U8580 (N_8580,N_8488,N_8414);
and U8581 (N_8581,N_8405,N_8421);
and U8582 (N_8582,N_8435,N_8475);
nand U8583 (N_8583,N_8451,N_8427);
nand U8584 (N_8584,N_8458,N_8479);
xor U8585 (N_8585,N_8407,N_8470);
xnor U8586 (N_8586,N_8444,N_8491);
and U8587 (N_8587,N_8436,N_8450);
and U8588 (N_8588,N_8415,N_8430);
xor U8589 (N_8589,N_8499,N_8415);
or U8590 (N_8590,N_8459,N_8452);
and U8591 (N_8591,N_8410,N_8441);
or U8592 (N_8592,N_8485,N_8405);
and U8593 (N_8593,N_8495,N_8458);
nor U8594 (N_8594,N_8418,N_8412);
or U8595 (N_8595,N_8403,N_8456);
or U8596 (N_8596,N_8485,N_8499);
xnor U8597 (N_8597,N_8443,N_8491);
or U8598 (N_8598,N_8455,N_8487);
xnor U8599 (N_8599,N_8436,N_8440);
or U8600 (N_8600,N_8591,N_8585);
or U8601 (N_8601,N_8566,N_8590);
nor U8602 (N_8602,N_8576,N_8500);
nand U8603 (N_8603,N_8545,N_8547);
nand U8604 (N_8604,N_8517,N_8515);
nor U8605 (N_8605,N_8529,N_8501);
and U8606 (N_8606,N_8553,N_8587);
and U8607 (N_8607,N_8595,N_8537);
and U8608 (N_8608,N_8575,N_8544);
nor U8609 (N_8609,N_8561,N_8514);
nor U8610 (N_8610,N_8534,N_8543);
nor U8611 (N_8611,N_8584,N_8552);
and U8612 (N_8612,N_8569,N_8535);
or U8613 (N_8613,N_8551,N_8546);
or U8614 (N_8614,N_8573,N_8507);
nand U8615 (N_8615,N_8586,N_8548);
or U8616 (N_8616,N_8568,N_8509);
or U8617 (N_8617,N_8571,N_8557);
nor U8618 (N_8618,N_8516,N_8554);
and U8619 (N_8619,N_8531,N_8583);
nor U8620 (N_8620,N_8511,N_8556);
nor U8621 (N_8621,N_8563,N_8570);
nor U8622 (N_8622,N_8592,N_8597);
or U8623 (N_8623,N_8588,N_8527);
and U8624 (N_8624,N_8521,N_8542);
or U8625 (N_8625,N_8503,N_8510);
nand U8626 (N_8626,N_8508,N_8505);
and U8627 (N_8627,N_8574,N_8578);
nor U8628 (N_8628,N_8565,N_8502);
or U8629 (N_8629,N_8530,N_8581);
nor U8630 (N_8630,N_8593,N_8532);
nor U8631 (N_8631,N_8522,N_8599);
xnor U8632 (N_8632,N_8533,N_8519);
nand U8633 (N_8633,N_8538,N_8512);
and U8634 (N_8634,N_8540,N_8518);
and U8635 (N_8635,N_8594,N_8596);
xor U8636 (N_8636,N_8560,N_8541);
xnor U8637 (N_8637,N_8528,N_8567);
xor U8638 (N_8638,N_8526,N_8564);
nand U8639 (N_8639,N_8555,N_8524);
xnor U8640 (N_8640,N_8558,N_8523);
nand U8641 (N_8641,N_8598,N_8562);
or U8642 (N_8642,N_8582,N_8579);
or U8643 (N_8643,N_8580,N_8520);
nand U8644 (N_8644,N_8559,N_8577);
or U8645 (N_8645,N_8550,N_8504);
xor U8646 (N_8646,N_8536,N_8539);
nand U8647 (N_8647,N_8549,N_8589);
nand U8648 (N_8648,N_8506,N_8513);
or U8649 (N_8649,N_8572,N_8525);
nand U8650 (N_8650,N_8573,N_8511);
nor U8651 (N_8651,N_8544,N_8550);
xnor U8652 (N_8652,N_8571,N_8594);
nor U8653 (N_8653,N_8548,N_8539);
nand U8654 (N_8654,N_8508,N_8528);
xor U8655 (N_8655,N_8538,N_8584);
and U8656 (N_8656,N_8590,N_8581);
xnor U8657 (N_8657,N_8538,N_8572);
nand U8658 (N_8658,N_8590,N_8586);
xnor U8659 (N_8659,N_8529,N_8561);
nand U8660 (N_8660,N_8583,N_8595);
nor U8661 (N_8661,N_8510,N_8577);
and U8662 (N_8662,N_8532,N_8543);
xor U8663 (N_8663,N_8565,N_8590);
xor U8664 (N_8664,N_8548,N_8567);
nand U8665 (N_8665,N_8513,N_8581);
nand U8666 (N_8666,N_8509,N_8593);
xor U8667 (N_8667,N_8546,N_8565);
or U8668 (N_8668,N_8506,N_8524);
and U8669 (N_8669,N_8508,N_8558);
nand U8670 (N_8670,N_8540,N_8571);
nand U8671 (N_8671,N_8582,N_8564);
nor U8672 (N_8672,N_8517,N_8565);
xor U8673 (N_8673,N_8576,N_8598);
xor U8674 (N_8674,N_8552,N_8542);
xor U8675 (N_8675,N_8584,N_8501);
nand U8676 (N_8676,N_8530,N_8570);
nor U8677 (N_8677,N_8594,N_8540);
nor U8678 (N_8678,N_8558,N_8528);
or U8679 (N_8679,N_8587,N_8582);
or U8680 (N_8680,N_8590,N_8540);
nor U8681 (N_8681,N_8580,N_8583);
nand U8682 (N_8682,N_8582,N_8528);
nand U8683 (N_8683,N_8549,N_8545);
and U8684 (N_8684,N_8560,N_8576);
nand U8685 (N_8685,N_8533,N_8571);
xnor U8686 (N_8686,N_8584,N_8591);
xnor U8687 (N_8687,N_8582,N_8599);
and U8688 (N_8688,N_8573,N_8537);
or U8689 (N_8689,N_8589,N_8582);
xnor U8690 (N_8690,N_8526,N_8537);
and U8691 (N_8691,N_8513,N_8537);
nand U8692 (N_8692,N_8500,N_8570);
xor U8693 (N_8693,N_8594,N_8525);
xnor U8694 (N_8694,N_8561,N_8530);
xnor U8695 (N_8695,N_8560,N_8543);
and U8696 (N_8696,N_8507,N_8598);
nor U8697 (N_8697,N_8578,N_8544);
xor U8698 (N_8698,N_8576,N_8567);
or U8699 (N_8699,N_8599,N_8502);
or U8700 (N_8700,N_8631,N_8623);
and U8701 (N_8701,N_8687,N_8607);
xor U8702 (N_8702,N_8652,N_8697);
nand U8703 (N_8703,N_8609,N_8693);
nand U8704 (N_8704,N_8620,N_8663);
or U8705 (N_8705,N_8622,N_8675);
xor U8706 (N_8706,N_8624,N_8658);
nor U8707 (N_8707,N_8629,N_8603);
xnor U8708 (N_8708,N_8659,N_8639);
nor U8709 (N_8709,N_8617,N_8679);
or U8710 (N_8710,N_8648,N_8626);
xor U8711 (N_8711,N_8656,N_8606);
xnor U8712 (N_8712,N_8612,N_8602);
or U8713 (N_8713,N_8673,N_8664);
nor U8714 (N_8714,N_8689,N_8614);
xor U8715 (N_8715,N_8666,N_8676);
nor U8716 (N_8716,N_8677,N_8699);
nand U8717 (N_8717,N_8650,N_8644);
and U8718 (N_8718,N_8691,N_8642);
xnor U8719 (N_8719,N_8695,N_8653);
and U8720 (N_8720,N_8627,N_8655);
or U8721 (N_8721,N_8665,N_8698);
nor U8722 (N_8722,N_8601,N_8635);
and U8723 (N_8723,N_8613,N_8660);
and U8724 (N_8724,N_8681,N_8683);
and U8725 (N_8725,N_8696,N_8645);
nor U8726 (N_8726,N_8657,N_8647);
or U8727 (N_8727,N_8662,N_8651);
nor U8728 (N_8728,N_8616,N_8661);
nand U8729 (N_8729,N_8628,N_8685);
nor U8730 (N_8730,N_8600,N_8605);
nand U8731 (N_8731,N_8680,N_8625);
nand U8732 (N_8732,N_8649,N_8688);
xnor U8733 (N_8733,N_8672,N_8674);
nor U8734 (N_8734,N_8610,N_8686);
nand U8735 (N_8735,N_8690,N_8621);
nand U8736 (N_8736,N_8643,N_8638);
and U8737 (N_8737,N_8671,N_8604);
nor U8738 (N_8738,N_8611,N_8667);
xnor U8739 (N_8739,N_8633,N_8668);
or U8740 (N_8740,N_8636,N_8670);
xor U8741 (N_8741,N_8654,N_8637);
nand U8742 (N_8742,N_8618,N_8608);
and U8743 (N_8743,N_8630,N_8619);
xnor U8744 (N_8744,N_8646,N_8641);
xnor U8745 (N_8745,N_8694,N_8692);
nand U8746 (N_8746,N_8682,N_8678);
and U8747 (N_8747,N_8684,N_8615);
nand U8748 (N_8748,N_8632,N_8640);
or U8749 (N_8749,N_8634,N_8669);
nand U8750 (N_8750,N_8689,N_8690);
nor U8751 (N_8751,N_8683,N_8671);
xor U8752 (N_8752,N_8616,N_8647);
and U8753 (N_8753,N_8694,N_8625);
or U8754 (N_8754,N_8618,N_8697);
nor U8755 (N_8755,N_8640,N_8623);
nor U8756 (N_8756,N_8641,N_8675);
and U8757 (N_8757,N_8603,N_8683);
xnor U8758 (N_8758,N_8600,N_8614);
and U8759 (N_8759,N_8657,N_8684);
nor U8760 (N_8760,N_8648,N_8638);
or U8761 (N_8761,N_8654,N_8685);
and U8762 (N_8762,N_8668,N_8670);
or U8763 (N_8763,N_8619,N_8607);
or U8764 (N_8764,N_8651,N_8683);
nor U8765 (N_8765,N_8629,N_8658);
and U8766 (N_8766,N_8613,N_8674);
or U8767 (N_8767,N_8609,N_8603);
nand U8768 (N_8768,N_8619,N_8635);
nor U8769 (N_8769,N_8677,N_8655);
nor U8770 (N_8770,N_8688,N_8693);
and U8771 (N_8771,N_8637,N_8662);
nor U8772 (N_8772,N_8634,N_8601);
or U8773 (N_8773,N_8609,N_8613);
and U8774 (N_8774,N_8603,N_8627);
nor U8775 (N_8775,N_8662,N_8695);
or U8776 (N_8776,N_8602,N_8679);
or U8777 (N_8777,N_8603,N_8656);
and U8778 (N_8778,N_8627,N_8607);
nand U8779 (N_8779,N_8683,N_8660);
nor U8780 (N_8780,N_8630,N_8656);
nor U8781 (N_8781,N_8657,N_8670);
or U8782 (N_8782,N_8650,N_8646);
or U8783 (N_8783,N_8603,N_8621);
nand U8784 (N_8784,N_8696,N_8663);
nand U8785 (N_8785,N_8637,N_8679);
xor U8786 (N_8786,N_8676,N_8634);
xor U8787 (N_8787,N_8672,N_8607);
xor U8788 (N_8788,N_8681,N_8644);
xor U8789 (N_8789,N_8667,N_8640);
nand U8790 (N_8790,N_8697,N_8662);
nor U8791 (N_8791,N_8691,N_8660);
nor U8792 (N_8792,N_8621,N_8657);
or U8793 (N_8793,N_8628,N_8629);
nor U8794 (N_8794,N_8659,N_8688);
and U8795 (N_8795,N_8660,N_8665);
and U8796 (N_8796,N_8612,N_8629);
or U8797 (N_8797,N_8667,N_8678);
or U8798 (N_8798,N_8669,N_8659);
nor U8799 (N_8799,N_8602,N_8625);
nor U8800 (N_8800,N_8756,N_8735);
nor U8801 (N_8801,N_8719,N_8760);
nand U8802 (N_8802,N_8741,N_8715);
xnor U8803 (N_8803,N_8733,N_8782);
and U8804 (N_8804,N_8749,N_8716);
and U8805 (N_8805,N_8779,N_8737);
nor U8806 (N_8806,N_8796,N_8799);
or U8807 (N_8807,N_8770,N_8758);
and U8808 (N_8808,N_8728,N_8711);
nor U8809 (N_8809,N_8710,N_8738);
nand U8810 (N_8810,N_8767,N_8776);
and U8811 (N_8811,N_8724,N_8722);
nor U8812 (N_8812,N_8708,N_8751);
xor U8813 (N_8813,N_8745,N_8721);
xor U8814 (N_8814,N_8766,N_8714);
nor U8815 (N_8815,N_8753,N_8713);
nand U8816 (N_8816,N_8784,N_8752);
or U8817 (N_8817,N_8706,N_8747);
and U8818 (N_8818,N_8717,N_8769);
nand U8819 (N_8819,N_8775,N_8754);
or U8820 (N_8820,N_8789,N_8720);
and U8821 (N_8821,N_8790,N_8763);
and U8822 (N_8822,N_8734,N_8778);
and U8823 (N_8823,N_8787,N_8765);
nor U8824 (N_8824,N_8742,N_8704);
nor U8825 (N_8825,N_8707,N_8774);
and U8826 (N_8826,N_8727,N_8750);
or U8827 (N_8827,N_8757,N_8772);
and U8828 (N_8828,N_8740,N_8773);
or U8829 (N_8829,N_8781,N_8761);
nand U8830 (N_8830,N_8709,N_8783);
or U8831 (N_8831,N_8712,N_8795);
nor U8832 (N_8832,N_8703,N_8777);
nor U8833 (N_8833,N_8771,N_8736);
nor U8834 (N_8834,N_8718,N_8744);
nand U8835 (N_8835,N_8791,N_8702);
xor U8836 (N_8836,N_8700,N_8729);
and U8837 (N_8837,N_8723,N_8743);
and U8838 (N_8838,N_8730,N_8788);
nand U8839 (N_8839,N_8726,N_8705);
nor U8840 (N_8840,N_8731,N_8793);
and U8841 (N_8841,N_8748,N_8762);
and U8842 (N_8842,N_8764,N_8785);
and U8843 (N_8843,N_8701,N_8797);
nand U8844 (N_8844,N_8780,N_8732);
or U8845 (N_8845,N_8798,N_8786);
nand U8846 (N_8846,N_8755,N_8792);
nand U8847 (N_8847,N_8768,N_8725);
xnor U8848 (N_8848,N_8794,N_8759);
nand U8849 (N_8849,N_8746,N_8739);
and U8850 (N_8850,N_8776,N_8793);
nand U8851 (N_8851,N_8773,N_8721);
nor U8852 (N_8852,N_8727,N_8770);
nor U8853 (N_8853,N_8720,N_8744);
or U8854 (N_8854,N_8724,N_8768);
or U8855 (N_8855,N_8742,N_8702);
xnor U8856 (N_8856,N_8775,N_8739);
xnor U8857 (N_8857,N_8751,N_8753);
or U8858 (N_8858,N_8763,N_8729);
nor U8859 (N_8859,N_8733,N_8750);
nor U8860 (N_8860,N_8761,N_8787);
nor U8861 (N_8861,N_8767,N_8739);
or U8862 (N_8862,N_8722,N_8778);
xor U8863 (N_8863,N_8734,N_8795);
and U8864 (N_8864,N_8705,N_8700);
nand U8865 (N_8865,N_8771,N_8770);
and U8866 (N_8866,N_8722,N_8750);
nor U8867 (N_8867,N_8748,N_8789);
xor U8868 (N_8868,N_8734,N_8776);
nor U8869 (N_8869,N_8702,N_8798);
or U8870 (N_8870,N_8727,N_8745);
nor U8871 (N_8871,N_8795,N_8718);
and U8872 (N_8872,N_8776,N_8705);
nand U8873 (N_8873,N_8766,N_8715);
nor U8874 (N_8874,N_8787,N_8727);
or U8875 (N_8875,N_8750,N_8798);
or U8876 (N_8876,N_8748,N_8720);
nand U8877 (N_8877,N_8702,N_8760);
xnor U8878 (N_8878,N_8704,N_8759);
nor U8879 (N_8879,N_8768,N_8700);
or U8880 (N_8880,N_8708,N_8739);
or U8881 (N_8881,N_8707,N_8795);
nor U8882 (N_8882,N_8742,N_8761);
nor U8883 (N_8883,N_8799,N_8758);
nor U8884 (N_8884,N_8745,N_8790);
nor U8885 (N_8885,N_8712,N_8730);
xor U8886 (N_8886,N_8708,N_8758);
and U8887 (N_8887,N_8751,N_8730);
or U8888 (N_8888,N_8758,N_8771);
xor U8889 (N_8889,N_8734,N_8735);
xnor U8890 (N_8890,N_8713,N_8747);
or U8891 (N_8891,N_8768,N_8758);
or U8892 (N_8892,N_8752,N_8771);
nand U8893 (N_8893,N_8787,N_8753);
and U8894 (N_8894,N_8740,N_8775);
xnor U8895 (N_8895,N_8732,N_8765);
xnor U8896 (N_8896,N_8701,N_8759);
xor U8897 (N_8897,N_8751,N_8721);
or U8898 (N_8898,N_8777,N_8786);
or U8899 (N_8899,N_8705,N_8727);
and U8900 (N_8900,N_8873,N_8845);
or U8901 (N_8901,N_8848,N_8894);
or U8902 (N_8902,N_8840,N_8854);
nand U8903 (N_8903,N_8898,N_8881);
and U8904 (N_8904,N_8816,N_8849);
nand U8905 (N_8905,N_8871,N_8855);
and U8906 (N_8906,N_8824,N_8812);
and U8907 (N_8907,N_8852,N_8828);
nor U8908 (N_8908,N_8893,N_8833);
or U8909 (N_8909,N_8832,N_8826);
and U8910 (N_8910,N_8823,N_8861);
nand U8911 (N_8911,N_8883,N_8880);
and U8912 (N_8912,N_8835,N_8866);
and U8913 (N_8913,N_8869,N_8856);
and U8914 (N_8914,N_8800,N_8841);
nand U8915 (N_8915,N_8885,N_8818);
nand U8916 (N_8916,N_8819,N_8810);
or U8917 (N_8917,N_8860,N_8872);
xnor U8918 (N_8918,N_8825,N_8837);
nand U8919 (N_8919,N_8878,N_8851);
xnor U8920 (N_8920,N_8865,N_8806);
nor U8921 (N_8921,N_8843,N_8867);
or U8922 (N_8922,N_8820,N_8827);
nand U8923 (N_8923,N_8846,N_8875);
or U8924 (N_8924,N_8815,N_8814);
nand U8925 (N_8925,N_8802,N_8884);
nor U8926 (N_8926,N_8879,N_8877);
and U8927 (N_8927,N_8887,N_8863);
and U8928 (N_8928,N_8892,N_8831);
or U8929 (N_8929,N_8817,N_8888);
nor U8930 (N_8930,N_8899,N_8813);
xor U8931 (N_8931,N_8842,N_8805);
or U8932 (N_8932,N_8821,N_8839);
nor U8933 (N_8933,N_8801,N_8895);
or U8934 (N_8934,N_8886,N_8809);
and U8935 (N_8935,N_8811,N_8874);
or U8936 (N_8936,N_8830,N_8829);
xor U8937 (N_8937,N_8870,N_8807);
and U8938 (N_8938,N_8889,N_8862);
nor U8939 (N_8939,N_8896,N_8803);
xor U8940 (N_8940,N_8847,N_8864);
xnor U8941 (N_8941,N_8857,N_8808);
or U8942 (N_8942,N_8858,N_8891);
nand U8943 (N_8943,N_8838,N_8853);
or U8944 (N_8944,N_8876,N_8836);
xor U8945 (N_8945,N_8850,N_8868);
xor U8946 (N_8946,N_8897,N_8834);
and U8947 (N_8947,N_8890,N_8844);
xnor U8948 (N_8948,N_8882,N_8822);
or U8949 (N_8949,N_8859,N_8804);
xor U8950 (N_8950,N_8819,N_8847);
and U8951 (N_8951,N_8877,N_8813);
nand U8952 (N_8952,N_8817,N_8809);
nand U8953 (N_8953,N_8894,N_8850);
or U8954 (N_8954,N_8804,N_8891);
and U8955 (N_8955,N_8879,N_8886);
nor U8956 (N_8956,N_8844,N_8851);
xnor U8957 (N_8957,N_8865,N_8866);
or U8958 (N_8958,N_8892,N_8882);
and U8959 (N_8959,N_8879,N_8885);
and U8960 (N_8960,N_8897,N_8874);
or U8961 (N_8961,N_8804,N_8877);
xnor U8962 (N_8962,N_8859,N_8883);
nand U8963 (N_8963,N_8860,N_8893);
and U8964 (N_8964,N_8869,N_8897);
nor U8965 (N_8965,N_8832,N_8818);
or U8966 (N_8966,N_8899,N_8838);
and U8967 (N_8967,N_8853,N_8806);
or U8968 (N_8968,N_8852,N_8858);
nand U8969 (N_8969,N_8878,N_8841);
or U8970 (N_8970,N_8857,N_8845);
nand U8971 (N_8971,N_8832,N_8810);
and U8972 (N_8972,N_8820,N_8837);
or U8973 (N_8973,N_8877,N_8831);
nor U8974 (N_8974,N_8893,N_8837);
or U8975 (N_8975,N_8856,N_8853);
or U8976 (N_8976,N_8862,N_8847);
and U8977 (N_8977,N_8884,N_8895);
xnor U8978 (N_8978,N_8890,N_8828);
xor U8979 (N_8979,N_8845,N_8828);
or U8980 (N_8980,N_8829,N_8886);
nand U8981 (N_8981,N_8882,N_8824);
nand U8982 (N_8982,N_8829,N_8807);
or U8983 (N_8983,N_8857,N_8877);
xor U8984 (N_8984,N_8829,N_8841);
and U8985 (N_8985,N_8802,N_8861);
or U8986 (N_8986,N_8868,N_8803);
or U8987 (N_8987,N_8820,N_8833);
and U8988 (N_8988,N_8882,N_8883);
xnor U8989 (N_8989,N_8864,N_8827);
and U8990 (N_8990,N_8811,N_8813);
or U8991 (N_8991,N_8830,N_8818);
and U8992 (N_8992,N_8807,N_8873);
or U8993 (N_8993,N_8812,N_8842);
and U8994 (N_8994,N_8811,N_8898);
nor U8995 (N_8995,N_8867,N_8859);
and U8996 (N_8996,N_8811,N_8879);
or U8997 (N_8997,N_8891,N_8854);
or U8998 (N_8998,N_8836,N_8844);
xor U8999 (N_8999,N_8809,N_8875);
nand U9000 (N_9000,N_8933,N_8990);
nor U9001 (N_9001,N_8976,N_8972);
nand U9002 (N_9002,N_8965,N_8907);
or U9003 (N_9003,N_8941,N_8920);
xor U9004 (N_9004,N_8902,N_8936);
or U9005 (N_9005,N_8993,N_8946);
xnor U9006 (N_9006,N_8904,N_8967);
or U9007 (N_9007,N_8999,N_8984);
or U9008 (N_9008,N_8908,N_8923);
and U9009 (N_9009,N_8981,N_8925);
xnor U9010 (N_9010,N_8914,N_8901);
or U9011 (N_9011,N_8996,N_8959);
and U9012 (N_9012,N_8906,N_8948);
xor U9013 (N_9013,N_8935,N_8950);
or U9014 (N_9014,N_8992,N_8956);
or U9015 (N_9015,N_8942,N_8932);
xnor U9016 (N_9016,N_8963,N_8998);
or U9017 (N_9017,N_8943,N_8947);
xor U9018 (N_9018,N_8939,N_8916);
and U9019 (N_9019,N_8960,N_8930);
nor U9020 (N_9020,N_8921,N_8980);
and U9021 (N_9021,N_8979,N_8903);
or U9022 (N_9022,N_8966,N_8919);
and U9023 (N_9023,N_8912,N_8911);
or U9024 (N_9024,N_8997,N_8927);
and U9025 (N_9025,N_8937,N_8961);
nor U9026 (N_9026,N_8982,N_8958);
xnor U9027 (N_9027,N_8971,N_8938);
and U9028 (N_9028,N_8985,N_8909);
nand U9029 (N_9029,N_8974,N_8949);
nand U9030 (N_9030,N_8968,N_8962);
and U9031 (N_9031,N_8964,N_8991);
or U9032 (N_9032,N_8955,N_8973);
nor U9033 (N_9033,N_8917,N_8957);
nor U9034 (N_9034,N_8995,N_8975);
nand U9035 (N_9035,N_8931,N_8986);
nor U9036 (N_9036,N_8918,N_8905);
xor U9037 (N_9037,N_8988,N_8987);
nand U9038 (N_9038,N_8940,N_8952);
nand U9039 (N_9039,N_8994,N_8945);
nand U9040 (N_9040,N_8951,N_8970);
nor U9041 (N_9041,N_8953,N_8954);
xor U9042 (N_9042,N_8924,N_8978);
and U9043 (N_9043,N_8928,N_8929);
or U9044 (N_9044,N_8915,N_8977);
and U9045 (N_9045,N_8944,N_8934);
xor U9046 (N_9046,N_8969,N_8900);
and U9047 (N_9047,N_8913,N_8922);
and U9048 (N_9048,N_8989,N_8983);
nor U9049 (N_9049,N_8926,N_8910);
nand U9050 (N_9050,N_8964,N_8930);
nand U9051 (N_9051,N_8928,N_8965);
or U9052 (N_9052,N_8918,N_8962);
xnor U9053 (N_9053,N_8919,N_8973);
and U9054 (N_9054,N_8919,N_8998);
nand U9055 (N_9055,N_8918,N_8999);
or U9056 (N_9056,N_8947,N_8986);
nand U9057 (N_9057,N_8939,N_8947);
nor U9058 (N_9058,N_8993,N_8904);
nor U9059 (N_9059,N_8916,N_8972);
or U9060 (N_9060,N_8942,N_8951);
and U9061 (N_9061,N_8926,N_8981);
or U9062 (N_9062,N_8925,N_8975);
xnor U9063 (N_9063,N_8943,N_8973);
xor U9064 (N_9064,N_8973,N_8977);
and U9065 (N_9065,N_8992,N_8929);
xnor U9066 (N_9066,N_8964,N_8974);
and U9067 (N_9067,N_8954,N_8935);
or U9068 (N_9068,N_8901,N_8977);
or U9069 (N_9069,N_8923,N_8948);
xnor U9070 (N_9070,N_8916,N_8957);
and U9071 (N_9071,N_8929,N_8922);
and U9072 (N_9072,N_8978,N_8927);
or U9073 (N_9073,N_8903,N_8992);
xnor U9074 (N_9074,N_8911,N_8929);
and U9075 (N_9075,N_8989,N_8922);
nor U9076 (N_9076,N_8998,N_8936);
and U9077 (N_9077,N_8947,N_8976);
nand U9078 (N_9078,N_8970,N_8905);
nor U9079 (N_9079,N_8999,N_8943);
nand U9080 (N_9080,N_8909,N_8908);
nand U9081 (N_9081,N_8911,N_8907);
nand U9082 (N_9082,N_8984,N_8905);
and U9083 (N_9083,N_8990,N_8961);
nor U9084 (N_9084,N_8972,N_8917);
nor U9085 (N_9085,N_8968,N_8988);
nand U9086 (N_9086,N_8907,N_8956);
nor U9087 (N_9087,N_8915,N_8900);
nand U9088 (N_9088,N_8932,N_8944);
and U9089 (N_9089,N_8961,N_8988);
and U9090 (N_9090,N_8943,N_8939);
or U9091 (N_9091,N_8905,N_8962);
xor U9092 (N_9092,N_8914,N_8992);
nand U9093 (N_9093,N_8971,N_8967);
xor U9094 (N_9094,N_8993,N_8925);
nand U9095 (N_9095,N_8987,N_8938);
nand U9096 (N_9096,N_8986,N_8995);
or U9097 (N_9097,N_8922,N_8918);
nand U9098 (N_9098,N_8915,N_8903);
and U9099 (N_9099,N_8931,N_8905);
or U9100 (N_9100,N_9031,N_9045);
or U9101 (N_9101,N_9032,N_9099);
xnor U9102 (N_9102,N_9040,N_9090);
xnor U9103 (N_9103,N_9005,N_9097);
or U9104 (N_9104,N_9025,N_9024);
nor U9105 (N_9105,N_9049,N_9014);
xnor U9106 (N_9106,N_9079,N_9036);
nor U9107 (N_9107,N_9053,N_9064);
or U9108 (N_9108,N_9018,N_9093);
nor U9109 (N_9109,N_9012,N_9086);
nand U9110 (N_9110,N_9088,N_9047);
or U9111 (N_9111,N_9075,N_9046);
or U9112 (N_9112,N_9077,N_9095);
nor U9113 (N_9113,N_9019,N_9000);
xnor U9114 (N_9114,N_9066,N_9001);
or U9115 (N_9115,N_9041,N_9062);
or U9116 (N_9116,N_9092,N_9085);
xnor U9117 (N_9117,N_9030,N_9034);
nand U9118 (N_9118,N_9058,N_9042);
xor U9119 (N_9119,N_9098,N_9052);
or U9120 (N_9120,N_9094,N_9009);
nand U9121 (N_9121,N_9087,N_9089);
and U9122 (N_9122,N_9013,N_9082);
or U9123 (N_9123,N_9057,N_9070);
nand U9124 (N_9124,N_9026,N_9011);
nand U9125 (N_9125,N_9023,N_9055);
and U9126 (N_9126,N_9033,N_9050);
and U9127 (N_9127,N_9027,N_9096);
or U9128 (N_9128,N_9074,N_9061);
and U9129 (N_9129,N_9037,N_9068);
and U9130 (N_9130,N_9039,N_9051);
or U9131 (N_9131,N_9016,N_9007);
and U9132 (N_9132,N_9038,N_9004);
and U9133 (N_9133,N_9017,N_9069);
or U9134 (N_9134,N_9044,N_9015);
xnor U9135 (N_9135,N_9003,N_9048);
and U9136 (N_9136,N_9028,N_9006);
nor U9137 (N_9137,N_9084,N_9054);
or U9138 (N_9138,N_9010,N_9056);
and U9139 (N_9139,N_9091,N_9060);
and U9140 (N_9140,N_9029,N_9071);
nand U9141 (N_9141,N_9043,N_9081);
xor U9142 (N_9142,N_9072,N_9083);
nor U9143 (N_9143,N_9078,N_9067);
and U9144 (N_9144,N_9022,N_9059);
nor U9145 (N_9145,N_9065,N_9076);
xnor U9146 (N_9146,N_9035,N_9021);
nand U9147 (N_9147,N_9008,N_9002);
nor U9148 (N_9148,N_9063,N_9080);
xor U9149 (N_9149,N_9020,N_9073);
and U9150 (N_9150,N_9087,N_9035);
xnor U9151 (N_9151,N_9052,N_9090);
and U9152 (N_9152,N_9011,N_9095);
and U9153 (N_9153,N_9048,N_9069);
and U9154 (N_9154,N_9013,N_9035);
nand U9155 (N_9155,N_9029,N_9027);
nor U9156 (N_9156,N_9027,N_9062);
or U9157 (N_9157,N_9094,N_9076);
nor U9158 (N_9158,N_9088,N_9051);
nand U9159 (N_9159,N_9090,N_9091);
or U9160 (N_9160,N_9067,N_9041);
nand U9161 (N_9161,N_9014,N_9057);
nand U9162 (N_9162,N_9075,N_9021);
and U9163 (N_9163,N_9023,N_9082);
nor U9164 (N_9164,N_9062,N_9018);
xor U9165 (N_9165,N_9091,N_9014);
and U9166 (N_9166,N_9074,N_9006);
and U9167 (N_9167,N_9099,N_9017);
xnor U9168 (N_9168,N_9018,N_9007);
xnor U9169 (N_9169,N_9062,N_9084);
or U9170 (N_9170,N_9049,N_9071);
or U9171 (N_9171,N_9058,N_9085);
nor U9172 (N_9172,N_9053,N_9016);
xnor U9173 (N_9173,N_9089,N_9051);
xnor U9174 (N_9174,N_9076,N_9028);
or U9175 (N_9175,N_9043,N_9053);
or U9176 (N_9176,N_9065,N_9016);
or U9177 (N_9177,N_9076,N_9081);
xor U9178 (N_9178,N_9084,N_9044);
nor U9179 (N_9179,N_9089,N_9069);
xor U9180 (N_9180,N_9065,N_9029);
and U9181 (N_9181,N_9025,N_9001);
xnor U9182 (N_9182,N_9024,N_9063);
nor U9183 (N_9183,N_9069,N_9057);
xnor U9184 (N_9184,N_9071,N_9060);
and U9185 (N_9185,N_9052,N_9048);
xor U9186 (N_9186,N_9016,N_9010);
nand U9187 (N_9187,N_9096,N_9059);
nor U9188 (N_9188,N_9024,N_9057);
or U9189 (N_9189,N_9017,N_9059);
nand U9190 (N_9190,N_9055,N_9015);
nor U9191 (N_9191,N_9031,N_9089);
or U9192 (N_9192,N_9010,N_9036);
or U9193 (N_9193,N_9056,N_9038);
and U9194 (N_9194,N_9094,N_9062);
or U9195 (N_9195,N_9005,N_9003);
nor U9196 (N_9196,N_9012,N_9082);
and U9197 (N_9197,N_9041,N_9071);
nand U9198 (N_9198,N_9092,N_9082);
nor U9199 (N_9199,N_9019,N_9095);
or U9200 (N_9200,N_9148,N_9138);
and U9201 (N_9201,N_9126,N_9131);
xnor U9202 (N_9202,N_9125,N_9112);
nor U9203 (N_9203,N_9183,N_9143);
or U9204 (N_9204,N_9171,N_9191);
xnor U9205 (N_9205,N_9108,N_9151);
and U9206 (N_9206,N_9167,N_9107);
and U9207 (N_9207,N_9113,N_9114);
nand U9208 (N_9208,N_9160,N_9110);
nor U9209 (N_9209,N_9116,N_9109);
nand U9210 (N_9210,N_9139,N_9169);
xor U9211 (N_9211,N_9128,N_9129);
xor U9212 (N_9212,N_9115,N_9154);
xnor U9213 (N_9213,N_9192,N_9137);
or U9214 (N_9214,N_9168,N_9177);
nand U9215 (N_9215,N_9117,N_9103);
and U9216 (N_9216,N_9144,N_9140);
xor U9217 (N_9217,N_9172,N_9174);
or U9218 (N_9218,N_9142,N_9179);
nand U9219 (N_9219,N_9185,N_9146);
nor U9220 (N_9220,N_9135,N_9181);
nor U9221 (N_9221,N_9180,N_9150);
nand U9222 (N_9222,N_9111,N_9159);
nand U9223 (N_9223,N_9106,N_9195);
nand U9224 (N_9224,N_9161,N_9188);
or U9225 (N_9225,N_9175,N_9120);
or U9226 (N_9226,N_9101,N_9127);
nand U9227 (N_9227,N_9102,N_9141);
nor U9228 (N_9228,N_9153,N_9193);
nor U9229 (N_9229,N_9122,N_9157);
nand U9230 (N_9230,N_9190,N_9100);
xnor U9231 (N_9231,N_9158,N_9194);
nor U9232 (N_9232,N_9134,N_9152);
nand U9233 (N_9233,N_9118,N_9132);
or U9234 (N_9234,N_9163,N_9189);
xor U9235 (N_9235,N_9178,N_9147);
nand U9236 (N_9236,N_9176,N_9187);
nor U9237 (N_9237,N_9173,N_9166);
or U9238 (N_9238,N_9149,N_9186);
or U9239 (N_9239,N_9133,N_9199);
nor U9240 (N_9240,N_9197,N_9156);
xor U9241 (N_9241,N_9124,N_9196);
nand U9242 (N_9242,N_9123,N_9170);
nor U9243 (N_9243,N_9136,N_9164);
xor U9244 (N_9244,N_9165,N_9155);
xnor U9245 (N_9245,N_9182,N_9119);
nand U9246 (N_9246,N_9130,N_9105);
xor U9247 (N_9247,N_9184,N_9145);
nor U9248 (N_9248,N_9162,N_9121);
or U9249 (N_9249,N_9104,N_9198);
xnor U9250 (N_9250,N_9166,N_9120);
and U9251 (N_9251,N_9165,N_9149);
xnor U9252 (N_9252,N_9140,N_9153);
xor U9253 (N_9253,N_9119,N_9123);
and U9254 (N_9254,N_9127,N_9123);
xnor U9255 (N_9255,N_9150,N_9139);
or U9256 (N_9256,N_9199,N_9127);
or U9257 (N_9257,N_9165,N_9182);
xnor U9258 (N_9258,N_9117,N_9136);
or U9259 (N_9259,N_9195,N_9145);
nor U9260 (N_9260,N_9115,N_9122);
nor U9261 (N_9261,N_9193,N_9154);
and U9262 (N_9262,N_9129,N_9167);
nor U9263 (N_9263,N_9117,N_9108);
nor U9264 (N_9264,N_9143,N_9193);
nor U9265 (N_9265,N_9195,N_9126);
nor U9266 (N_9266,N_9134,N_9174);
or U9267 (N_9267,N_9164,N_9118);
and U9268 (N_9268,N_9171,N_9192);
nand U9269 (N_9269,N_9156,N_9102);
and U9270 (N_9270,N_9140,N_9127);
and U9271 (N_9271,N_9118,N_9161);
or U9272 (N_9272,N_9146,N_9160);
nand U9273 (N_9273,N_9199,N_9130);
nor U9274 (N_9274,N_9157,N_9142);
nand U9275 (N_9275,N_9121,N_9158);
or U9276 (N_9276,N_9148,N_9125);
xnor U9277 (N_9277,N_9124,N_9190);
nor U9278 (N_9278,N_9155,N_9129);
or U9279 (N_9279,N_9119,N_9135);
nor U9280 (N_9280,N_9173,N_9149);
nand U9281 (N_9281,N_9197,N_9118);
or U9282 (N_9282,N_9128,N_9187);
or U9283 (N_9283,N_9170,N_9112);
nand U9284 (N_9284,N_9144,N_9134);
or U9285 (N_9285,N_9153,N_9114);
and U9286 (N_9286,N_9116,N_9154);
nand U9287 (N_9287,N_9140,N_9199);
nand U9288 (N_9288,N_9132,N_9128);
xor U9289 (N_9289,N_9139,N_9170);
and U9290 (N_9290,N_9119,N_9151);
xnor U9291 (N_9291,N_9129,N_9100);
nor U9292 (N_9292,N_9146,N_9104);
xor U9293 (N_9293,N_9111,N_9118);
nor U9294 (N_9294,N_9188,N_9195);
nor U9295 (N_9295,N_9115,N_9100);
or U9296 (N_9296,N_9132,N_9182);
and U9297 (N_9297,N_9149,N_9156);
xnor U9298 (N_9298,N_9136,N_9141);
or U9299 (N_9299,N_9172,N_9132);
nand U9300 (N_9300,N_9265,N_9223);
xnor U9301 (N_9301,N_9248,N_9275);
nor U9302 (N_9302,N_9243,N_9209);
and U9303 (N_9303,N_9210,N_9250);
nor U9304 (N_9304,N_9227,N_9281);
xor U9305 (N_9305,N_9235,N_9279);
nor U9306 (N_9306,N_9283,N_9284);
nand U9307 (N_9307,N_9202,N_9290);
nor U9308 (N_9308,N_9222,N_9291);
or U9309 (N_9309,N_9269,N_9207);
or U9310 (N_9310,N_9262,N_9219);
xnor U9311 (N_9311,N_9236,N_9232);
xor U9312 (N_9312,N_9220,N_9251);
or U9313 (N_9313,N_9212,N_9211);
nand U9314 (N_9314,N_9257,N_9256);
xnor U9315 (N_9315,N_9225,N_9252);
nor U9316 (N_9316,N_9263,N_9258);
nor U9317 (N_9317,N_9289,N_9267);
or U9318 (N_9318,N_9285,N_9214);
nand U9319 (N_9319,N_9260,N_9268);
nor U9320 (N_9320,N_9244,N_9273);
or U9321 (N_9321,N_9218,N_9204);
or U9322 (N_9322,N_9295,N_9217);
and U9323 (N_9323,N_9255,N_9297);
or U9324 (N_9324,N_9270,N_9292);
or U9325 (N_9325,N_9200,N_9205);
nor U9326 (N_9326,N_9278,N_9293);
or U9327 (N_9327,N_9282,N_9298);
and U9328 (N_9328,N_9233,N_9238);
or U9329 (N_9329,N_9261,N_9208);
nor U9330 (N_9330,N_9277,N_9229);
xnor U9331 (N_9331,N_9254,N_9213);
and U9332 (N_9332,N_9239,N_9215);
xor U9333 (N_9333,N_9224,N_9226);
or U9334 (N_9334,N_9280,N_9287);
or U9335 (N_9335,N_9266,N_9246);
or U9336 (N_9336,N_9242,N_9247);
nor U9337 (N_9337,N_9240,N_9294);
or U9338 (N_9338,N_9264,N_9231);
nand U9339 (N_9339,N_9253,N_9271);
xnor U9340 (N_9340,N_9228,N_9286);
xnor U9341 (N_9341,N_9216,N_9249);
and U9342 (N_9342,N_9234,N_9259);
nand U9343 (N_9343,N_9272,N_9201);
xor U9344 (N_9344,N_9206,N_9245);
xnor U9345 (N_9345,N_9221,N_9288);
nand U9346 (N_9346,N_9203,N_9296);
or U9347 (N_9347,N_9241,N_9237);
or U9348 (N_9348,N_9299,N_9274);
or U9349 (N_9349,N_9230,N_9276);
or U9350 (N_9350,N_9244,N_9201);
or U9351 (N_9351,N_9246,N_9220);
nand U9352 (N_9352,N_9279,N_9273);
nand U9353 (N_9353,N_9249,N_9206);
and U9354 (N_9354,N_9264,N_9234);
and U9355 (N_9355,N_9229,N_9265);
or U9356 (N_9356,N_9266,N_9233);
nor U9357 (N_9357,N_9286,N_9298);
nand U9358 (N_9358,N_9234,N_9273);
or U9359 (N_9359,N_9292,N_9248);
nand U9360 (N_9360,N_9236,N_9269);
and U9361 (N_9361,N_9248,N_9218);
or U9362 (N_9362,N_9254,N_9272);
xnor U9363 (N_9363,N_9253,N_9259);
nor U9364 (N_9364,N_9246,N_9237);
or U9365 (N_9365,N_9232,N_9260);
and U9366 (N_9366,N_9293,N_9267);
nand U9367 (N_9367,N_9206,N_9246);
xor U9368 (N_9368,N_9284,N_9230);
xnor U9369 (N_9369,N_9273,N_9274);
or U9370 (N_9370,N_9200,N_9287);
nand U9371 (N_9371,N_9277,N_9218);
or U9372 (N_9372,N_9226,N_9264);
nand U9373 (N_9373,N_9272,N_9258);
nand U9374 (N_9374,N_9252,N_9288);
nand U9375 (N_9375,N_9275,N_9217);
and U9376 (N_9376,N_9250,N_9253);
xnor U9377 (N_9377,N_9282,N_9297);
nand U9378 (N_9378,N_9290,N_9204);
xor U9379 (N_9379,N_9262,N_9272);
nand U9380 (N_9380,N_9266,N_9272);
xnor U9381 (N_9381,N_9230,N_9246);
or U9382 (N_9382,N_9207,N_9225);
nor U9383 (N_9383,N_9201,N_9232);
or U9384 (N_9384,N_9213,N_9265);
and U9385 (N_9385,N_9282,N_9214);
nand U9386 (N_9386,N_9220,N_9222);
nor U9387 (N_9387,N_9253,N_9266);
or U9388 (N_9388,N_9211,N_9243);
nor U9389 (N_9389,N_9239,N_9259);
xnor U9390 (N_9390,N_9228,N_9261);
xnor U9391 (N_9391,N_9226,N_9228);
nor U9392 (N_9392,N_9237,N_9275);
xnor U9393 (N_9393,N_9238,N_9247);
nor U9394 (N_9394,N_9233,N_9299);
nand U9395 (N_9395,N_9213,N_9203);
or U9396 (N_9396,N_9270,N_9230);
xnor U9397 (N_9397,N_9203,N_9236);
xor U9398 (N_9398,N_9260,N_9227);
or U9399 (N_9399,N_9219,N_9266);
xor U9400 (N_9400,N_9328,N_9372);
xor U9401 (N_9401,N_9301,N_9337);
xor U9402 (N_9402,N_9313,N_9343);
nand U9403 (N_9403,N_9310,N_9389);
and U9404 (N_9404,N_9362,N_9391);
xor U9405 (N_9405,N_9342,N_9374);
or U9406 (N_9406,N_9380,N_9358);
nor U9407 (N_9407,N_9361,N_9333);
nor U9408 (N_9408,N_9327,N_9302);
or U9409 (N_9409,N_9352,N_9365);
or U9410 (N_9410,N_9395,N_9335);
and U9411 (N_9411,N_9363,N_9306);
or U9412 (N_9412,N_9368,N_9318);
nor U9413 (N_9413,N_9378,N_9324);
xnor U9414 (N_9414,N_9314,N_9329);
or U9415 (N_9415,N_9323,N_9396);
nand U9416 (N_9416,N_9387,N_9311);
and U9417 (N_9417,N_9382,N_9367);
or U9418 (N_9418,N_9347,N_9394);
and U9419 (N_9419,N_9312,N_9336);
nor U9420 (N_9420,N_9340,N_9307);
or U9421 (N_9421,N_9345,N_9317);
nor U9422 (N_9422,N_9341,N_9353);
or U9423 (N_9423,N_9351,N_9392);
or U9424 (N_9424,N_9393,N_9308);
and U9425 (N_9425,N_9356,N_9379);
and U9426 (N_9426,N_9386,N_9300);
and U9427 (N_9427,N_9377,N_9364);
or U9428 (N_9428,N_9331,N_9399);
nand U9429 (N_9429,N_9388,N_9390);
xnor U9430 (N_9430,N_9360,N_9320);
nor U9431 (N_9431,N_9383,N_9381);
nor U9432 (N_9432,N_9366,N_9369);
or U9433 (N_9433,N_9321,N_9338);
xor U9434 (N_9434,N_9332,N_9397);
or U9435 (N_9435,N_9350,N_9304);
nor U9436 (N_9436,N_9315,N_9309);
nor U9437 (N_9437,N_9376,N_9370);
nor U9438 (N_9438,N_9357,N_9384);
xor U9439 (N_9439,N_9373,N_9359);
and U9440 (N_9440,N_9322,N_9348);
and U9441 (N_9441,N_9326,N_9371);
or U9442 (N_9442,N_9354,N_9325);
and U9443 (N_9443,N_9346,N_9339);
nor U9444 (N_9444,N_9319,N_9316);
nand U9445 (N_9445,N_9305,N_9398);
nand U9446 (N_9446,N_9385,N_9355);
nand U9447 (N_9447,N_9344,N_9330);
or U9448 (N_9448,N_9303,N_9375);
or U9449 (N_9449,N_9334,N_9349);
or U9450 (N_9450,N_9329,N_9313);
and U9451 (N_9451,N_9361,N_9344);
nand U9452 (N_9452,N_9346,N_9337);
xnor U9453 (N_9453,N_9384,N_9388);
and U9454 (N_9454,N_9382,N_9301);
and U9455 (N_9455,N_9350,N_9314);
nand U9456 (N_9456,N_9391,N_9370);
nor U9457 (N_9457,N_9374,N_9313);
or U9458 (N_9458,N_9368,N_9351);
nor U9459 (N_9459,N_9365,N_9328);
nor U9460 (N_9460,N_9396,N_9300);
or U9461 (N_9461,N_9377,N_9342);
or U9462 (N_9462,N_9325,N_9305);
nand U9463 (N_9463,N_9350,N_9305);
nand U9464 (N_9464,N_9397,N_9399);
xnor U9465 (N_9465,N_9378,N_9376);
nand U9466 (N_9466,N_9355,N_9345);
xor U9467 (N_9467,N_9322,N_9306);
or U9468 (N_9468,N_9310,N_9301);
or U9469 (N_9469,N_9304,N_9364);
nand U9470 (N_9470,N_9396,N_9349);
nor U9471 (N_9471,N_9379,N_9369);
nand U9472 (N_9472,N_9363,N_9384);
nor U9473 (N_9473,N_9342,N_9370);
xnor U9474 (N_9474,N_9326,N_9332);
or U9475 (N_9475,N_9379,N_9325);
xnor U9476 (N_9476,N_9388,N_9385);
xnor U9477 (N_9477,N_9305,N_9320);
nand U9478 (N_9478,N_9365,N_9315);
and U9479 (N_9479,N_9370,N_9397);
and U9480 (N_9480,N_9347,N_9342);
and U9481 (N_9481,N_9377,N_9399);
and U9482 (N_9482,N_9372,N_9344);
xnor U9483 (N_9483,N_9350,N_9347);
xnor U9484 (N_9484,N_9381,N_9309);
nor U9485 (N_9485,N_9303,N_9312);
xor U9486 (N_9486,N_9343,N_9300);
and U9487 (N_9487,N_9321,N_9363);
xor U9488 (N_9488,N_9345,N_9370);
or U9489 (N_9489,N_9335,N_9332);
and U9490 (N_9490,N_9380,N_9355);
and U9491 (N_9491,N_9339,N_9342);
xnor U9492 (N_9492,N_9346,N_9307);
nand U9493 (N_9493,N_9326,N_9380);
or U9494 (N_9494,N_9355,N_9396);
nand U9495 (N_9495,N_9307,N_9303);
nand U9496 (N_9496,N_9382,N_9361);
and U9497 (N_9497,N_9332,N_9347);
nor U9498 (N_9498,N_9398,N_9319);
nor U9499 (N_9499,N_9387,N_9379);
nor U9500 (N_9500,N_9403,N_9401);
nand U9501 (N_9501,N_9454,N_9430);
or U9502 (N_9502,N_9414,N_9494);
nor U9503 (N_9503,N_9442,N_9436);
and U9504 (N_9504,N_9460,N_9418);
xnor U9505 (N_9505,N_9416,N_9408);
and U9506 (N_9506,N_9409,N_9423);
xor U9507 (N_9507,N_9496,N_9448);
nand U9508 (N_9508,N_9417,N_9437);
nand U9509 (N_9509,N_9459,N_9455);
nor U9510 (N_9510,N_9480,N_9491);
and U9511 (N_9511,N_9485,N_9488);
or U9512 (N_9512,N_9434,N_9464);
or U9513 (N_9513,N_9478,N_9486);
or U9514 (N_9514,N_9477,N_9407);
xor U9515 (N_9515,N_9429,N_9481);
or U9516 (N_9516,N_9427,N_9497);
or U9517 (N_9517,N_9405,N_9440);
xnor U9518 (N_9518,N_9465,N_9461);
nor U9519 (N_9519,N_9411,N_9487);
and U9520 (N_9520,N_9449,N_9447);
and U9521 (N_9521,N_9475,N_9467);
nor U9522 (N_9522,N_9483,N_9473);
xor U9523 (N_9523,N_9492,N_9446);
or U9524 (N_9524,N_9443,N_9439);
nor U9525 (N_9525,N_9462,N_9428);
and U9526 (N_9526,N_9466,N_9404);
xor U9527 (N_9527,N_9471,N_9433);
nor U9528 (N_9528,N_9435,N_9472);
and U9529 (N_9529,N_9463,N_9490);
or U9530 (N_9530,N_9484,N_9402);
xor U9531 (N_9531,N_9426,N_9489);
and U9532 (N_9532,N_9498,N_9476);
and U9533 (N_9533,N_9450,N_9441);
xor U9534 (N_9534,N_9432,N_9419);
nand U9535 (N_9535,N_9420,N_9451);
nand U9536 (N_9536,N_9452,N_9456);
nand U9537 (N_9537,N_9431,N_9406);
and U9538 (N_9538,N_9438,N_9410);
or U9539 (N_9539,N_9474,N_9458);
xnor U9540 (N_9540,N_9415,N_9422);
and U9541 (N_9541,N_9445,N_9413);
nand U9542 (N_9542,N_9412,N_9499);
or U9543 (N_9543,N_9444,N_9493);
and U9544 (N_9544,N_9469,N_9479);
xnor U9545 (N_9545,N_9421,N_9468);
xnor U9546 (N_9546,N_9495,N_9457);
nor U9547 (N_9547,N_9424,N_9482);
and U9548 (N_9548,N_9425,N_9453);
or U9549 (N_9549,N_9470,N_9400);
nand U9550 (N_9550,N_9438,N_9444);
nand U9551 (N_9551,N_9490,N_9425);
or U9552 (N_9552,N_9421,N_9477);
nand U9553 (N_9553,N_9411,N_9456);
xor U9554 (N_9554,N_9498,N_9484);
nor U9555 (N_9555,N_9430,N_9462);
nand U9556 (N_9556,N_9465,N_9428);
and U9557 (N_9557,N_9421,N_9475);
or U9558 (N_9558,N_9463,N_9472);
nor U9559 (N_9559,N_9453,N_9467);
nor U9560 (N_9560,N_9405,N_9445);
xnor U9561 (N_9561,N_9431,N_9473);
nor U9562 (N_9562,N_9419,N_9445);
xor U9563 (N_9563,N_9445,N_9406);
or U9564 (N_9564,N_9401,N_9433);
nand U9565 (N_9565,N_9468,N_9450);
xor U9566 (N_9566,N_9483,N_9480);
and U9567 (N_9567,N_9404,N_9497);
xnor U9568 (N_9568,N_9447,N_9470);
and U9569 (N_9569,N_9446,N_9458);
or U9570 (N_9570,N_9473,N_9470);
nand U9571 (N_9571,N_9411,N_9446);
xor U9572 (N_9572,N_9477,N_9404);
nor U9573 (N_9573,N_9429,N_9400);
and U9574 (N_9574,N_9498,N_9440);
nor U9575 (N_9575,N_9407,N_9487);
xor U9576 (N_9576,N_9459,N_9475);
and U9577 (N_9577,N_9484,N_9444);
or U9578 (N_9578,N_9445,N_9484);
xnor U9579 (N_9579,N_9411,N_9430);
or U9580 (N_9580,N_9454,N_9419);
or U9581 (N_9581,N_9403,N_9453);
or U9582 (N_9582,N_9459,N_9418);
nand U9583 (N_9583,N_9449,N_9412);
and U9584 (N_9584,N_9430,N_9472);
xor U9585 (N_9585,N_9455,N_9412);
nor U9586 (N_9586,N_9410,N_9432);
and U9587 (N_9587,N_9416,N_9452);
xor U9588 (N_9588,N_9462,N_9455);
and U9589 (N_9589,N_9427,N_9490);
or U9590 (N_9590,N_9409,N_9474);
and U9591 (N_9591,N_9432,N_9493);
or U9592 (N_9592,N_9402,N_9411);
xnor U9593 (N_9593,N_9486,N_9414);
or U9594 (N_9594,N_9485,N_9460);
or U9595 (N_9595,N_9444,N_9481);
nor U9596 (N_9596,N_9452,N_9463);
nor U9597 (N_9597,N_9462,N_9447);
nor U9598 (N_9598,N_9419,N_9428);
and U9599 (N_9599,N_9489,N_9429);
xnor U9600 (N_9600,N_9533,N_9501);
nand U9601 (N_9601,N_9507,N_9544);
or U9602 (N_9602,N_9550,N_9591);
xnor U9603 (N_9603,N_9578,N_9529);
nand U9604 (N_9604,N_9521,N_9536);
or U9605 (N_9605,N_9569,N_9534);
nand U9606 (N_9606,N_9508,N_9598);
nand U9607 (N_9607,N_9543,N_9581);
or U9608 (N_9608,N_9509,N_9575);
nand U9609 (N_9609,N_9535,N_9545);
nand U9610 (N_9610,N_9519,N_9585);
or U9611 (N_9611,N_9551,N_9587);
xor U9612 (N_9612,N_9574,N_9559);
nor U9613 (N_9613,N_9566,N_9557);
and U9614 (N_9614,N_9546,N_9553);
and U9615 (N_9615,N_9531,N_9511);
xor U9616 (N_9616,N_9554,N_9512);
nand U9617 (N_9617,N_9570,N_9594);
xor U9618 (N_9618,N_9586,N_9523);
nor U9619 (N_9619,N_9580,N_9571);
or U9620 (N_9620,N_9518,N_9515);
nor U9621 (N_9621,N_9597,N_9549);
nor U9622 (N_9622,N_9592,N_9505);
or U9623 (N_9623,N_9541,N_9522);
and U9624 (N_9624,N_9567,N_9526);
and U9625 (N_9625,N_9540,N_9556);
and U9626 (N_9626,N_9506,N_9542);
and U9627 (N_9627,N_9514,N_9583);
xor U9628 (N_9628,N_9524,N_9568);
and U9629 (N_9629,N_9577,N_9547);
nand U9630 (N_9630,N_9510,N_9528);
xnor U9631 (N_9631,N_9596,N_9517);
or U9632 (N_9632,N_9503,N_9563);
or U9633 (N_9633,N_9589,N_9537);
nand U9634 (N_9634,N_9565,N_9572);
xor U9635 (N_9635,N_9538,N_9579);
nor U9636 (N_9636,N_9582,N_9576);
or U9637 (N_9637,N_9564,N_9560);
or U9638 (N_9638,N_9593,N_9527);
xnor U9639 (N_9639,N_9513,N_9555);
nand U9640 (N_9640,N_9590,N_9502);
or U9641 (N_9641,N_9599,N_9573);
nor U9642 (N_9642,N_9584,N_9532);
or U9643 (N_9643,N_9500,N_9562);
and U9644 (N_9644,N_9561,N_9530);
or U9645 (N_9645,N_9525,N_9548);
nand U9646 (N_9646,N_9539,N_9516);
xnor U9647 (N_9647,N_9504,N_9520);
nor U9648 (N_9648,N_9558,N_9588);
and U9649 (N_9649,N_9595,N_9552);
nand U9650 (N_9650,N_9540,N_9562);
xor U9651 (N_9651,N_9533,N_9587);
xnor U9652 (N_9652,N_9560,N_9504);
nor U9653 (N_9653,N_9567,N_9548);
or U9654 (N_9654,N_9567,N_9506);
and U9655 (N_9655,N_9513,N_9516);
or U9656 (N_9656,N_9514,N_9597);
nor U9657 (N_9657,N_9539,N_9595);
or U9658 (N_9658,N_9595,N_9585);
xor U9659 (N_9659,N_9584,N_9586);
and U9660 (N_9660,N_9551,N_9560);
xor U9661 (N_9661,N_9505,N_9511);
or U9662 (N_9662,N_9583,N_9542);
nor U9663 (N_9663,N_9563,N_9585);
or U9664 (N_9664,N_9558,N_9509);
or U9665 (N_9665,N_9585,N_9567);
or U9666 (N_9666,N_9554,N_9535);
nand U9667 (N_9667,N_9546,N_9535);
nor U9668 (N_9668,N_9529,N_9512);
xor U9669 (N_9669,N_9541,N_9579);
or U9670 (N_9670,N_9581,N_9517);
nor U9671 (N_9671,N_9589,N_9561);
xnor U9672 (N_9672,N_9553,N_9508);
nor U9673 (N_9673,N_9548,N_9588);
nor U9674 (N_9674,N_9540,N_9559);
nor U9675 (N_9675,N_9506,N_9527);
xor U9676 (N_9676,N_9590,N_9545);
or U9677 (N_9677,N_9594,N_9513);
nor U9678 (N_9678,N_9517,N_9502);
nand U9679 (N_9679,N_9535,N_9597);
nor U9680 (N_9680,N_9535,N_9569);
and U9681 (N_9681,N_9504,N_9595);
nand U9682 (N_9682,N_9593,N_9554);
and U9683 (N_9683,N_9520,N_9543);
nand U9684 (N_9684,N_9551,N_9554);
and U9685 (N_9685,N_9560,N_9597);
or U9686 (N_9686,N_9564,N_9509);
nor U9687 (N_9687,N_9591,N_9596);
xnor U9688 (N_9688,N_9591,N_9521);
and U9689 (N_9689,N_9506,N_9589);
nand U9690 (N_9690,N_9598,N_9592);
nand U9691 (N_9691,N_9509,N_9585);
nor U9692 (N_9692,N_9531,N_9592);
xor U9693 (N_9693,N_9547,N_9500);
or U9694 (N_9694,N_9564,N_9568);
nand U9695 (N_9695,N_9532,N_9543);
nor U9696 (N_9696,N_9510,N_9511);
nand U9697 (N_9697,N_9580,N_9566);
xnor U9698 (N_9698,N_9537,N_9506);
nor U9699 (N_9699,N_9543,N_9531);
nand U9700 (N_9700,N_9653,N_9656);
nand U9701 (N_9701,N_9634,N_9646);
and U9702 (N_9702,N_9639,N_9647);
and U9703 (N_9703,N_9660,N_9674);
nand U9704 (N_9704,N_9636,N_9612);
nand U9705 (N_9705,N_9682,N_9607);
or U9706 (N_9706,N_9611,N_9615);
nand U9707 (N_9707,N_9625,N_9618);
xor U9708 (N_9708,N_9680,N_9694);
xnor U9709 (N_9709,N_9635,N_9619);
or U9710 (N_9710,N_9604,N_9666);
nor U9711 (N_9711,N_9690,N_9672);
or U9712 (N_9712,N_9693,N_9630);
nand U9713 (N_9713,N_9628,N_9663);
or U9714 (N_9714,N_9600,N_9652);
nand U9715 (N_9715,N_9687,N_9629);
xnor U9716 (N_9716,N_9622,N_9621);
and U9717 (N_9717,N_9698,N_9685);
xnor U9718 (N_9718,N_9673,N_9627);
xor U9719 (N_9719,N_9648,N_9601);
nor U9720 (N_9720,N_9662,N_9679);
nor U9721 (N_9721,N_9632,N_9605);
and U9722 (N_9722,N_9633,N_9624);
xnor U9723 (N_9723,N_9691,N_9603);
or U9724 (N_9724,N_9642,N_9677);
and U9725 (N_9725,N_9670,N_9692);
xor U9726 (N_9726,N_9610,N_9637);
or U9727 (N_9727,N_9608,N_9631);
nand U9728 (N_9728,N_9683,N_9609);
nand U9729 (N_9729,N_9658,N_9684);
xnor U9730 (N_9730,N_9699,N_9678);
or U9731 (N_9731,N_9688,N_9614);
nand U9732 (N_9732,N_9657,N_9626);
and U9733 (N_9733,N_9649,N_9659);
xnor U9734 (N_9734,N_9606,N_9697);
nand U9735 (N_9735,N_9669,N_9668);
nor U9736 (N_9736,N_9623,N_9664);
nor U9737 (N_9737,N_9644,N_9645);
and U9738 (N_9738,N_9643,N_9661);
or U9739 (N_9739,N_9641,N_9686);
and U9740 (N_9740,N_9617,N_9638);
nand U9741 (N_9741,N_9616,N_9671);
nor U9742 (N_9742,N_9620,N_9689);
nor U9743 (N_9743,N_9675,N_9650);
nand U9744 (N_9744,N_9602,N_9613);
or U9745 (N_9745,N_9665,N_9651);
xnor U9746 (N_9746,N_9667,N_9681);
and U9747 (N_9747,N_9695,N_9654);
or U9748 (N_9748,N_9696,N_9655);
nor U9749 (N_9749,N_9676,N_9640);
and U9750 (N_9750,N_9637,N_9631);
or U9751 (N_9751,N_9600,N_9627);
nor U9752 (N_9752,N_9628,N_9662);
nor U9753 (N_9753,N_9639,N_9664);
nor U9754 (N_9754,N_9669,N_9600);
or U9755 (N_9755,N_9614,N_9639);
and U9756 (N_9756,N_9616,N_9658);
nand U9757 (N_9757,N_9677,N_9661);
or U9758 (N_9758,N_9613,N_9637);
or U9759 (N_9759,N_9615,N_9685);
and U9760 (N_9760,N_9642,N_9687);
and U9761 (N_9761,N_9698,N_9649);
nand U9762 (N_9762,N_9619,N_9607);
nor U9763 (N_9763,N_9668,N_9617);
and U9764 (N_9764,N_9685,N_9617);
xor U9765 (N_9765,N_9688,N_9627);
or U9766 (N_9766,N_9649,N_9678);
nand U9767 (N_9767,N_9691,N_9643);
nor U9768 (N_9768,N_9634,N_9641);
nand U9769 (N_9769,N_9606,N_9693);
and U9770 (N_9770,N_9660,N_9651);
or U9771 (N_9771,N_9624,N_9605);
nand U9772 (N_9772,N_9630,N_9683);
or U9773 (N_9773,N_9676,N_9697);
nand U9774 (N_9774,N_9603,N_9695);
nor U9775 (N_9775,N_9669,N_9683);
nand U9776 (N_9776,N_9691,N_9681);
xor U9777 (N_9777,N_9698,N_9628);
or U9778 (N_9778,N_9670,N_9612);
xnor U9779 (N_9779,N_9686,N_9683);
and U9780 (N_9780,N_9620,N_9644);
and U9781 (N_9781,N_9681,N_9647);
nor U9782 (N_9782,N_9625,N_9685);
and U9783 (N_9783,N_9627,N_9613);
nand U9784 (N_9784,N_9614,N_9690);
nor U9785 (N_9785,N_9697,N_9609);
xor U9786 (N_9786,N_9636,N_9606);
and U9787 (N_9787,N_9620,N_9627);
or U9788 (N_9788,N_9604,N_9645);
and U9789 (N_9789,N_9635,N_9600);
xnor U9790 (N_9790,N_9619,N_9689);
and U9791 (N_9791,N_9670,N_9604);
xnor U9792 (N_9792,N_9609,N_9649);
xor U9793 (N_9793,N_9673,N_9601);
xor U9794 (N_9794,N_9684,N_9646);
xor U9795 (N_9795,N_9692,N_9631);
nor U9796 (N_9796,N_9694,N_9614);
nor U9797 (N_9797,N_9624,N_9659);
or U9798 (N_9798,N_9622,N_9616);
or U9799 (N_9799,N_9676,N_9636);
nor U9800 (N_9800,N_9781,N_9727);
nor U9801 (N_9801,N_9728,N_9709);
and U9802 (N_9802,N_9759,N_9716);
and U9803 (N_9803,N_9708,N_9723);
xnor U9804 (N_9804,N_9717,N_9786);
or U9805 (N_9805,N_9740,N_9747);
xor U9806 (N_9806,N_9751,N_9736);
nand U9807 (N_9807,N_9731,N_9772);
and U9808 (N_9808,N_9720,N_9700);
xnor U9809 (N_9809,N_9719,N_9792);
and U9810 (N_9810,N_9732,N_9707);
and U9811 (N_9811,N_9788,N_9785);
and U9812 (N_9812,N_9758,N_9710);
xor U9813 (N_9813,N_9743,N_9755);
or U9814 (N_9814,N_9765,N_9715);
nand U9815 (N_9815,N_9799,N_9722);
nor U9816 (N_9816,N_9741,N_9771);
xor U9817 (N_9817,N_9783,N_9795);
nor U9818 (N_9818,N_9791,N_9711);
nand U9819 (N_9819,N_9763,N_9746);
or U9820 (N_9820,N_9729,N_9738);
and U9821 (N_9821,N_9737,N_9750);
nand U9822 (N_9822,N_9770,N_9757);
xnor U9823 (N_9823,N_9773,N_9744);
nand U9824 (N_9824,N_9724,N_9735);
nand U9825 (N_9825,N_9793,N_9718);
xnor U9826 (N_9826,N_9797,N_9730);
nand U9827 (N_9827,N_9752,N_9742);
nand U9828 (N_9828,N_9733,N_9714);
xor U9829 (N_9829,N_9767,N_9725);
nor U9830 (N_9830,N_9777,N_9721);
nand U9831 (N_9831,N_9774,N_9753);
and U9832 (N_9832,N_9794,N_9779);
or U9833 (N_9833,N_9701,N_9748);
nor U9834 (N_9834,N_9796,N_9798);
and U9835 (N_9835,N_9745,N_9734);
and U9836 (N_9836,N_9789,N_9787);
nand U9837 (N_9837,N_9754,N_9782);
nand U9838 (N_9838,N_9778,N_9739);
nand U9839 (N_9839,N_9705,N_9756);
xnor U9840 (N_9840,N_9780,N_9790);
nand U9841 (N_9841,N_9713,N_9760);
and U9842 (N_9842,N_9776,N_9704);
nor U9843 (N_9843,N_9784,N_9703);
nand U9844 (N_9844,N_9702,N_9762);
and U9845 (N_9845,N_9726,N_9712);
and U9846 (N_9846,N_9775,N_9764);
or U9847 (N_9847,N_9768,N_9766);
nand U9848 (N_9848,N_9749,N_9769);
nor U9849 (N_9849,N_9761,N_9706);
nand U9850 (N_9850,N_9766,N_9795);
xnor U9851 (N_9851,N_9744,N_9746);
nand U9852 (N_9852,N_9735,N_9752);
nor U9853 (N_9853,N_9706,N_9733);
nor U9854 (N_9854,N_9767,N_9745);
nor U9855 (N_9855,N_9788,N_9754);
xor U9856 (N_9856,N_9716,N_9764);
nor U9857 (N_9857,N_9719,N_9780);
nand U9858 (N_9858,N_9721,N_9700);
nand U9859 (N_9859,N_9749,N_9787);
nand U9860 (N_9860,N_9763,N_9755);
and U9861 (N_9861,N_9704,N_9740);
xnor U9862 (N_9862,N_9731,N_9785);
xor U9863 (N_9863,N_9730,N_9786);
nor U9864 (N_9864,N_9746,N_9765);
and U9865 (N_9865,N_9747,N_9798);
or U9866 (N_9866,N_9748,N_9772);
xor U9867 (N_9867,N_9787,N_9791);
or U9868 (N_9868,N_9719,N_9733);
or U9869 (N_9869,N_9780,N_9770);
and U9870 (N_9870,N_9717,N_9796);
nand U9871 (N_9871,N_9744,N_9735);
nand U9872 (N_9872,N_9717,N_9728);
xnor U9873 (N_9873,N_9753,N_9776);
nor U9874 (N_9874,N_9721,N_9722);
nand U9875 (N_9875,N_9777,N_9758);
nor U9876 (N_9876,N_9753,N_9710);
and U9877 (N_9877,N_9791,N_9703);
and U9878 (N_9878,N_9790,N_9794);
or U9879 (N_9879,N_9785,N_9777);
xor U9880 (N_9880,N_9783,N_9794);
nand U9881 (N_9881,N_9702,N_9774);
nor U9882 (N_9882,N_9714,N_9717);
nand U9883 (N_9883,N_9789,N_9762);
xor U9884 (N_9884,N_9742,N_9759);
nor U9885 (N_9885,N_9727,N_9782);
nand U9886 (N_9886,N_9737,N_9711);
nor U9887 (N_9887,N_9722,N_9753);
or U9888 (N_9888,N_9761,N_9745);
nor U9889 (N_9889,N_9711,N_9734);
xnor U9890 (N_9890,N_9781,N_9780);
or U9891 (N_9891,N_9754,N_9727);
nand U9892 (N_9892,N_9794,N_9745);
nor U9893 (N_9893,N_9793,N_9717);
nor U9894 (N_9894,N_9798,N_9782);
and U9895 (N_9895,N_9745,N_9738);
nand U9896 (N_9896,N_9799,N_9760);
nand U9897 (N_9897,N_9731,N_9712);
xnor U9898 (N_9898,N_9751,N_9739);
and U9899 (N_9899,N_9792,N_9784);
nor U9900 (N_9900,N_9809,N_9816);
or U9901 (N_9901,N_9832,N_9848);
nand U9902 (N_9902,N_9887,N_9895);
and U9903 (N_9903,N_9889,N_9833);
nor U9904 (N_9904,N_9899,N_9877);
or U9905 (N_9905,N_9853,N_9883);
xnor U9906 (N_9906,N_9852,N_9825);
and U9907 (N_9907,N_9885,N_9893);
or U9908 (N_9908,N_9827,N_9836);
nor U9909 (N_9909,N_9828,N_9842);
xor U9910 (N_9910,N_9850,N_9864);
xnor U9911 (N_9911,N_9865,N_9826);
nor U9912 (N_9912,N_9841,N_9886);
nand U9913 (N_9913,N_9837,N_9805);
xor U9914 (N_9914,N_9811,N_9878);
nand U9915 (N_9915,N_9803,N_9846);
xnor U9916 (N_9916,N_9856,N_9849);
nor U9917 (N_9917,N_9874,N_9822);
nor U9918 (N_9918,N_9892,N_9804);
nor U9919 (N_9919,N_9834,N_9843);
or U9920 (N_9920,N_9808,N_9830);
or U9921 (N_9921,N_9857,N_9800);
nor U9922 (N_9922,N_9835,N_9819);
xnor U9923 (N_9923,N_9847,N_9840);
nor U9924 (N_9924,N_9894,N_9838);
nor U9925 (N_9925,N_9817,N_9813);
nand U9926 (N_9926,N_9801,N_9862);
xor U9927 (N_9927,N_9875,N_9882);
xor U9928 (N_9928,N_9860,N_9814);
and U9929 (N_9929,N_9851,N_9897);
nor U9930 (N_9930,N_9858,N_9867);
nor U9931 (N_9931,N_9879,N_9880);
nor U9932 (N_9932,N_9871,N_9812);
nand U9933 (N_9933,N_9855,N_9820);
and U9934 (N_9934,N_9818,N_9815);
or U9935 (N_9935,N_9839,N_9845);
and U9936 (N_9936,N_9863,N_9888);
xnor U9937 (N_9937,N_9866,N_9861);
and U9938 (N_9938,N_9890,N_9898);
xor U9939 (N_9939,N_9831,N_9896);
and U9940 (N_9940,N_9810,N_9873);
or U9941 (N_9941,N_9854,N_9872);
and U9942 (N_9942,N_9876,N_9881);
xnor U9943 (N_9943,N_9829,N_9806);
or U9944 (N_9944,N_9859,N_9823);
xnor U9945 (N_9945,N_9802,N_9869);
and U9946 (N_9946,N_9884,N_9891);
xnor U9947 (N_9947,N_9824,N_9868);
and U9948 (N_9948,N_9807,N_9870);
or U9949 (N_9949,N_9821,N_9844);
nor U9950 (N_9950,N_9831,N_9854);
xor U9951 (N_9951,N_9859,N_9845);
nand U9952 (N_9952,N_9833,N_9852);
and U9953 (N_9953,N_9899,N_9826);
or U9954 (N_9954,N_9894,N_9802);
nand U9955 (N_9955,N_9893,N_9866);
nand U9956 (N_9956,N_9880,N_9872);
nor U9957 (N_9957,N_9835,N_9897);
nor U9958 (N_9958,N_9804,N_9882);
xor U9959 (N_9959,N_9887,N_9810);
nand U9960 (N_9960,N_9892,N_9805);
xor U9961 (N_9961,N_9807,N_9879);
xnor U9962 (N_9962,N_9878,N_9847);
nor U9963 (N_9963,N_9831,N_9884);
xor U9964 (N_9964,N_9821,N_9865);
nor U9965 (N_9965,N_9889,N_9844);
xor U9966 (N_9966,N_9873,N_9862);
or U9967 (N_9967,N_9850,N_9832);
nor U9968 (N_9968,N_9805,N_9808);
nor U9969 (N_9969,N_9874,N_9850);
nor U9970 (N_9970,N_9887,N_9862);
nand U9971 (N_9971,N_9836,N_9889);
or U9972 (N_9972,N_9830,N_9875);
nand U9973 (N_9973,N_9801,N_9886);
or U9974 (N_9974,N_9828,N_9836);
xor U9975 (N_9975,N_9844,N_9895);
xnor U9976 (N_9976,N_9855,N_9869);
nand U9977 (N_9977,N_9862,N_9826);
nand U9978 (N_9978,N_9873,N_9871);
xor U9979 (N_9979,N_9857,N_9804);
nand U9980 (N_9980,N_9889,N_9897);
xor U9981 (N_9981,N_9829,N_9832);
and U9982 (N_9982,N_9874,N_9846);
and U9983 (N_9983,N_9876,N_9863);
nand U9984 (N_9984,N_9819,N_9896);
nand U9985 (N_9985,N_9869,N_9895);
or U9986 (N_9986,N_9860,N_9818);
xor U9987 (N_9987,N_9805,N_9898);
or U9988 (N_9988,N_9878,N_9809);
and U9989 (N_9989,N_9837,N_9806);
or U9990 (N_9990,N_9880,N_9809);
nor U9991 (N_9991,N_9848,N_9890);
xnor U9992 (N_9992,N_9807,N_9839);
xnor U9993 (N_9993,N_9865,N_9888);
or U9994 (N_9994,N_9821,N_9840);
xnor U9995 (N_9995,N_9833,N_9813);
xnor U9996 (N_9996,N_9883,N_9831);
and U9997 (N_9997,N_9860,N_9844);
nand U9998 (N_9998,N_9893,N_9810);
xor U9999 (N_9999,N_9859,N_9890);
xor UO_0 (O_0,N_9969,N_9941);
xor UO_1 (O_1,N_9959,N_9949);
or UO_2 (O_2,N_9929,N_9993);
or UO_3 (O_3,N_9908,N_9913);
and UO_4 (O_4,N_9980,N_9922);
and UO_5 (O_5,N_9911,N_9910);
and UO_6 (O_6,N_9924,N_9972);
nor UO_7 (O_7,N_9914,N_9920);
xnor UO_8 (O_8,N_9971,N_9947);
and UO_9 (O_9,N_9940,N_9997);
and UO_10 (O_10,N_9944,N_9932);
and UO_11 (O_11,N_9902,N_9936);
nand UO_12 (O_12,N_9937,N_9990);
nand UO_13 (O_13,N_9954,N_9968);
and UO_14 (O_14,N_9953,N_9943);
xor UO_15 (O_15,N_9916,N_9927);
or UO_16 (O_16,N_9984,N_9967);
xnor UO_17 (O_17,N_9994,N_9991);
and UO_18 (O_18,N_9973,N_9939);
nor UO_19 (O_19,N_9963,N_9956);
xor UO_20 (O_20,N_9983,N_9962);
nor UO_21 (O_21,N_9900,N_9903);
or UO_22 (O_22,N_9930,N_9907);
or UO_23 (O_23,N_9964,N_9975);
and UO_24 (O_24,N_9942,N_9934);
or UO_25 (O_25,N_9912,N_9950);
nand UO_26 (O_26,N_9951,N_9901);
nor UO_27 (O_27,N_9952,N_9928);
nor UO_28 (O_28,N_9935,N_9988);
nand UO_29 (O_29,N_9982,N_9958);
nor UO_30 (O_30,N_9909,N_9926);
or UO_31 (O_31,N_9981,N_9985);
and UO_32 (O_32,N_9957,N_9974);
xnor UO_33 (O_33,N_9946,N_9965);
nand UO_34 (O_34,N_9918,N_9978);
and UO_35 (O_35,N_9986,N_9919);
or UO_36 (O_36,N_9989,N_9955);
xor UO_37 (O_37,N_9999,N_9961);
and UO_38 (O_38,N_9995,N_9917);
and UO_39 (O_39,N_9945,N_9998);
nor UO_40 (O_40,N_9925,N_9992);
nand UO_41 (O_41,N_9906,N_9904);
and UO_42 (O_42,N_9960,N_9938);
xnor UO_43 (O_43,N_9933,N_9966);
and UO_44 (O_44,N_9977,N_9948);
or UO_45 (O_45,N_9976,N_9931);
or UO_46 (O_46,N_9905,N_9915);
nand UO_47 (O_47,N_9996,N_9923);
or UO_48 (O_48,N_9979,N_9921);
nor UO_49 (O_49,N_9970,N_9987);
or UO_50 (O_50,N_9979,N_9902);
or UO_51 (O_51,N_9906,N_9957);
or UO_52 (O_52,N_9984,N_9941);
nor UO_53 (O_53,N_9974,N_9913);
nor UO_54 (O_54,N_9907,N_9929);
xnor UO_55 (O_55,N_9919,N_9904);
or UO_56 (O_56,N_9977,N_9958);
nand UO_57 (O_57,N_9901,N_9930);
and UO_58 (O_58,N_9922,N_9901);
or UO_59 (O_59,N_9994,N_9997);
nor UO_60 (O_60,N_9938,N_9948);
or UO_61 (O_61,N_9934,N_9993);
or UO_62 (O_62,N_9959,N_9900);
nor UO_63 (O_63,N_9922,N_9911);
xnor UO_64 (O_64,N_9940,N_9977);
nor UO_65 (O_65,N_9923,N_9907);
nand UO_66 (O_66,N_9906,N_9935);
nand UO_67 (O_67,N_9917,N_9991);
nand UO_68 (O_68,N_9984,N_9980);
and UO_69 (O_69,N_9965,N_9906);
or UO_70 (O_70,N_9996,N_9974);
and UO_71 (O_71,N_9988,N_9947);
nor UO_72 (O_72,N_9947,N_9931);
nand UO_73 (O_73,N_9900,N_9964);
and UO_74 (O_74,N_9989,N_9910);
and UO_75 (O_75,N_9956,N_9908);
nand UO_76 (O_76,N_9930,N_9968);
nor UO_77 (O_77,N_9972,N_9979);
nand UO_78 (O_78,N_9999,N_9919);
or UO_79 (O_79,N_9984,N_9954);
nor UO_80 (O_80,N_9941,N_9931);
nand UO_81 (O_81,N_9940,N_9948);
and UO_82 (O_82,N_9900,N_9913);
or UO_83 (O_83,N_9987,N_9960);
nor UO_84 (O_84,N_9918,N_9997);
nor UO_85 (O_85,N_9989,N_9916);
xnor UO_86 (O_86,N_9977,N_9913);
or UO_87 (O_87,N_9941,N_9968);
or UO_88 (O_88,N_9905,N_9956);
xnor UO_89 (O_89,N_9953,N_9936);
xnor UO_90 (O_90,N_9965,N_9901);
xor UO_91 (O_91,N_9989,N_9918);
nor UO_92 (O_92,N_9993,N_9921);
and UO_93 (O_93,N_9996,N_9901);
xnor UO_94 (O_94,N_9994,N_9995);
or UO_95 (O_95,N_9959,N_9954);
or UO_96 (O_96,N_9977,N_9939);
or UO_97 (O_97,N_9963,N_9988);
and UO_98 (O_98,N_9911,N_9918);
and UO_99 (O_99,N_9951,N_9936);
or UO_100 (O_100,N_9923,N_9998);
nand UO_101 (O_101,N_9961,N_9964);
nor UO_102 (O_102,N_9990,N_9914);
or UO_103 (O_103,N_9937,N_9997);
nand UO_104 (O_104,N_9992,N_9982);
nand UO_105 (O_105,N_9974,N_9972);
or UO_106 (O_106,N_9976,N_9934);
or UO_107 (O_107,N_9953,N_9980);
and UO_108 (O_108,N_9977,N_9931);
nor UO_109 (O_109,N_9947,N_9903);
and UO_110 (O_110,N_9918,N_9971);
nand UO_111 (O_111,N_9929,N_9955);
xor UO_112 (O_112,N_9999,N_9925);
and UO_113 (O_113,N_9931,N_9961);
xor UO_114 (O_114,N_9930,N_9949);
and UO_115 (O_115,N_9960,N_9975);
nand UO_116 (O_116,N_9995,N_9947);
xnor UO_117 (O_117,N_9996,N_9985);
or UO_118 (O_118,N_9935,N_9984);
nand UO_119 (O_119,N_9965,N_9990);
xnor UO_120 (O_120,N_9971,N_9911);
and UO_121 (O_121,N_9942,N_9980);
and UO_122 (O_122,N_9936,N_9965);
xnor UO_123 (O_123,N_9993,N_9990);
nand UO_124 (O_124,N_9964,N_9993);
or UO_125 (O_125,N_9926,N_9985);
and UO_126 (O_126,N_9916,N_9932);
nand UO_127 (O_127,N_9996,N_9947);
nor UO_128 (O_128,N_9939,N_9946);
nand UO_129 (O_129,N_9999,N_9943);
nand UO_130 (O_130,N_9947,N_9919);
nand UO_131 (O_131,N_9944,N_9988);
nand UO_132 (O_132,N_9958,N_9988);
nor UO_133 (O_133,N_9985,N_9915);
xnor UO_134 (O_134,N_9955,N_9903);
or UO_135 (O_135,N_9957,N_9958);
xor UO_136 (O_136,N_9968,N_9993);
or UO_137 (O_137,N_9957,N_9943);
and UO_138 (O_138,N_9904,N_9987);
nand UO_139 (O_139,N_9994,N_9990);
xnor UO_140 (O_140,N_9988,N_9999);
and UO_141 (O_141,N_9913,N_9961);
nand UO_142 (O_142,N_9957,N_9920);
xor UO_143 (O_143,N_9947,N_9967);
nand UO_144 (O_144,N_9991,N_9924);
and UO_145 (O_145,N_9990,N_9950);
xnor UO_146 (O_146,N_9949,N_9927);
or UO_147 (O_147,N_9963,N_9907);
nor UO_148 (O_148,N_9903,N_9926);
and UO_149 (O_149,N_9971,N_9955);
nand UO_150 (O_150,N_9942,N_9948);
or UO_151 (O_151,N_9929,N_9923);
and UO_152 (O_152,N_9977,N_9965);
nand UO_153 (O_153,N_9909,N_9922);
xnor UO_154 (O_154,N_9991,N_9995);
nor UO_155 (O_155,N_9956,N_9975);
and UO_156 (O_156,N_9958,N_9947);
xor UO_157 (O_157,N_9948,N_9964);
xor UO_158 (O_158,N_9996,N_9904);
nor UO_159 (O_159,N_9925,N_9991);
or UO_160 (O_160,N_9981,N_9900);
and UO_161 (O_161,N_9965,N_9980);
and UO_162 (O_162,N_9938,N_9945);
nand UO_163 (O_163,N_9953,N_9928);
xor UO_164 (O_164,N_9939,N_9936);
and UO_165 (O_165,N_9991,N_9935);
xnor UO_166 (O_166,N_9965,N_9987);
nand UO_167 (O_167,N_9958,N_9914);
and UO_168 (O_168,N_9998,N_9980);
nand UO_169 (O_169,N_9919,N_9984);
and UO_170 (O_170,N_9928,N_9923);
nand UO_171 (O_171,N_9967,N_9926);
and UO_172 (O_172,N_9987,N_9986);
or UO_173 (O_173,N_9909,N_9951);
and UO_174 (O_174,N_9967,N_9979);
or UO_175 (O_175,N_9957,N_9984);
and UO_176 (O_176,N_9905,N_9944);
and UO_177 (O_177,N_9987,N_9996);
nand UO_178 (O_178,N_9930,N_9925);
nand UO_179 (O_179,N_9937,N_9992);
nor UO_180 (O_180,N_9959,N_9938);
or UO_181 (O_181,N_9924,N_9963);
nand UO_182 (O_182,N_9940,N_9961);
and UO_183 (O_183,N_9964,N_9912);
nand UO_184 (O_184,N_9971,N_9929);
xor UO_185 (O_185,N_9905,N_9919);
nor UO_186 (O_186,N_9984,N_9943);
and UO_187 (O_187,N_9905,N_9990);
nand UO_188 (O_188,N_9972,N_9965);
or UO_189 (O_189,N_9916,N_9922);
xnor UO_190 (O_190,N_9944,N_9997);
nand UO_191 (O_191,N_9953,N_9961);
nor UO_192 (O_192,N_9997,N_9964);
nor UO_193 (O_193,N_9993,N_9935);
and UO_194 (O_194,N_9910,N_9941);
nor UO_195 (O_195,N_9993,N_9948);
nand UO_196 (O_196,N_9982,N_9930);
nand UO_197 (O_197,N_9982,N_9907);
or UO_198 (O_198,N_9982,N_9940);
nor UO_199 (O_199,N_9903,N_9941);
and UO_200 (O_200,N_9965,N_9925);
nor UO_201 (O_201,N_9960,N_9981);
and UO_202 (O_202,N_9924,N_9988);
or UO_203 (O_203,N_9950,N_9930);
and UO_204 (O_204,N_9913,N_9992);
nor UO_205 (O_205,N_9954,N_9992);
nand UO_206 (O_206,N_9922,N_9971);
and UO_207 (O_207,N_9900,N_9907);
nor UO_208 (O_208,N_9981,N_9968);
xor UO_209 (O_209,N_9962,N_9946);
or UO_210 (O_210,N_9942,N_9963);
nor UO_211 (O_211,N_9957,N_9968);
nor UO_212 (O_212,N_9908,N_9902);
and UO_213 (O_213,N_9974,N_9973);
nor UO_214 (O_214,N_9923,N_9987);
or UO_215 (O_215,N_9985,N_9918);
or UO_216 (O_216,N_9961,N_9959);
or UO_217 (O_217,N_9998,N_9908);
xnor UO_218 (O_218,N_9905,N_9903);
or UO_219 (O_219,N_9998,N_9946);
nor UO_220 (O_220,N_9900,N_9933);
nand UO_221 (O_221,N_9922,N_9986);
xnor UO_222 (O_222,N_9952,N_9959);
and UO_223 (O_223,N_9955,N_9962);
and UO_224 (O_224,N_9900,N_9911);
nor UO_225 (O_225,N_9944,N_9918);
or UO_226 (O_226,N_9937,N_9930);
and UO_227 (O_227,N_9918,N_9937);
and UO_228 (O_228,N_9955,N_9944);
nand UO_229 (O_229,N_9923,N_9916);
or UO_230 (O_230,N_9999,N_9903);
nand UO_231 (O_231,N_9960,N_9922);
nor UO_232 (O_232,N_9941,N_9990);
nand UO_233 (O_233,N_9961,N_9974);
or UO_234 (O_234,N_9967,N_9975);
or UO_235 (O_235,N_9913,N_9965);
or UO_236 (O_236,N_9942,N_9926);
and UO_237 (O_237,N_9989,N_9935);
nor UO_238 (O_238,N_9976,N_9952);
nand UO_239 (O_239,N_9931,N_9916);
and UO_240 (O_240,N_9991,N_9938);
nand UO_241 (O_241,N_9920,N_9941);
xnor UO_242 (O_242,N_9940,N_9960);
or UO_243 (O_243,N_9980,N_9960);
nand UO_244 (O_244,N_9990,N_9957);
and UO_245 (O_245,N_9931,N_9920);
xor UO_246 (O_246,N_9971,N_9952);
nand UO_247 (O_247,N_9954,N_9901);
nand UO_248 (O_248,N_9981,N_9938);
nor UO_249 (O_249,N_9953,N_9941);
and UO_250 (O_250,N_9947,N_9973);
nor UO_251 (O_251,N_9990,N_9949);
nand UO_252 (O_252,N_9919,N_9962);
or UO_253 (O_253,N_9964,N_9973);
xor UO_254 (O_254,N_9939,N_9985);
nand UO_255 (O_255,N_9976,N_9905);
and UO_256 (O_256,N_9917,N_9960);
or UO_257 (O_257,N_9974,N_9911);
or UO_258 (O_258,N_9932,N_9972);
nor UO_259 (O_259,N_9976,N_9922);
and UO_260 (O_260,N_9915,N_9995);
and UO_261 (O_261,N_9975,N_9963);
or UO_262 (O_262,N_9904,N_9947);
or UO_263 (O_263,N_9981,N_9948);
xor UO_264 (O_264,N_9936,N_9966);
and UO_265 (O_265,N_9932,N_9953);
or UO_266 (O_266,N_9950,N_9994);
and UO_267 (O_267,N_9989,N_9964);
or UO_268 (O_268,N_9904,N_9924);
or UO_269 (O_269,N_9962,N_9922);
nor UO_270 (O_270,N_9967,N_9991);
nor UO_271 (O_271,N_9993,N_9946);
or UO_272 (O_272,N_9938,N_9985);
nand UO_273 (O_273,N_9946,N_9997);
nand UO_274 (O_274,N_9933,N_9980);
xor UO_275 (O_275,N_9935,N_9902);
and UO_276 (O_276,N_9935,N_9981);
xor UO_277 (O_277,N_9966,N_9952);
xor UO_278 (O_278,N_9926,N_9955);
nor UO_279 (O_279,N_9912,N_9930);
and UO_280 (O_280,N_9949,N_9988);
and UO_281 (O_281,N_9999,N_9922);
and UO_282 (O_282,N_9903,N_9977);
and UO_283 (O_283,N_9900,N_9991);
xor UO_284 (O_284,N_9989,N_9909);
or UO_285 (O_285,N_9932,N_9934);
or UO_286 (O_286,N_9916,N_9918);
nand UO_287 (O_287,N_9972,N_9954);
xor UO_288 (O_288,N_9951,N_9982);
xnor UO_289 (O_289,N_9918,N_9938);
or UO_290 (O_290,N_9909,N_9908);
or UO_291 (O_291,N_9939,N_9996);
or UO_292 (O_292,N_9924,N_9938);
xor UO_293 (O_293,N_9971,N_9985);
and UO_294 (O_294,N_9905,N_9941);
nand UO_295 (O_295,N_9974,N_9921);
xnor UO_296 (O_296,N_9910,N_9939);
nor UO_297 (O_297,N_9903,N_9928);
nor UO_298 (O_298,N_9902,N_9978);
xor UO_299 (O_299,N_9942,N_9930);
or UO_300 (O_300,N_9977,N_9901);
and UO_301 (O_301,N_9922,N_9936);
xnor UO_302 (O_302,N_9946,N_9930);
nand UO_303 (O_303,N_9980,N_9971);
and UO_304 (O_304,N_9902,N_9941);
or UO_305 (O_305,N_9981,N_9990);
nor UO_306 (O_306,N_9973,N_9999);
xnor UO_307 (O_307,N_9982,N_9967);
nand UO_308 (O_308,N_9983,N_9948);
xnor UO_309 (O_309,N_9943,N_9947);
or UO_310 (O_310,N_9968,N_9923);
nor UO_311 (O_311,N_9962,N_9904);
nor UO_312 (O_312,N_9976,N_9948);
nand UO_313 (O_313,N_9937,N_9949);
nor UO_314 (O_314,N_9944,N_9974);
and UO_315 (O_315,N_9951,N_9935);
or UO_316 (O_316,N_9908,N_9904);
or UO_317 (O_317,N_9909,N_9991);
nand UO_318 (O_318,N_9927,N_9938);
or UO_319 (O_319,N_9914,N_9944);
or UO_320 (O_320,N_9903,N_9923);
xor UO_321 (O_321,N_9942,N_9979);
nor UO_322 (O_322,N_9928,N_9999);
xor UO_323 (O_323,N_9932,N_9912);
nand UO_324 (O_324,N_9947,N_9986);
xor UO_325 (O_325,N_9948,N_9932);
nor UO_326 (O_326,N_9989,N_9959);
or UO_327 (O_327,N_9953,N_9979);
xor UO_328 (O_328,N_9950,N_9957);
xnor UO_329 (O_329,N_9951,N_9975);
xor UO_330 (O_330,N_9911,N_9990);
nand UO_331 (O_331,N_9953,N_9935);
or UO_332 (O_332,N_9933,N_9918);
and UO_333 (O_333,N_9976,N_9987);
and UO_334 (O_334,N_9995,N_9945);
xor UO_335 (O_335,N_9902,N_9916);
nor UO_336 (O_336,N_9951,N_9957);
xnor UO_337 (O_337,N_9964,N_9903);
and UO_338 (O_338,N_9945,N_9944);
or UO_339 (O_339,N_9979,N_9946);
or UO_340 (O_340,N_9908,N_9969);
nand UO_341 (O_341,N_9987,N_9930);
nand UO_342 (O_342,N_9940,N_9981);
xnor UO_343 (O_343,N_9953,N_9983);
nor UO_344 (O_344,N_9988,N_9910);
nor UO_345 (O_345,N_9966,N_9961);
nand UO_346 (O_346,N_9980,N_9900);
and UO_347 (O_347,N_9920,N_9977);
nand UO_348 (O_348,N_9917,N_9918);
and UO_349 (O_349,N_9979,N_9927);
or UO_350 (O_350,N_9938,N_9913);
and UO_351 (O_351,N_9940,N_9906);
or UO_352 (O_352,N_9975,N_9942);
and UO_353 (O_353,N_9986,N_9983);
nor UO_354 (O_354,N_9992,N_9926);
xnor UO_355 (O_355,N_9932,N_9976);
or UO_356 (O_356,N_9937,N_9969);
xnor UO_357 (O_357,N_9977,N_9905);
or UO_358 (O_358,N_9917,N_9947);
xor UO_359 (O_359,N_9946,N_9977);
nor UO_360 (O_360,N_9911,N_9982);
nor UO_361 (O_361,N_9940,N_9921);
and UO_362 (O_362,N_9947,N_9937);
or UO_363 (O_363,N_9944,N_9950);
nor UO_364 (O_364,N_9991,N_9905);
or UO_365 (O_365,N_9981,N_9989);
and UO_366 (O_366,N_9957,N_9911);
nand UO_367 (O_367,N_9933,N_9964);
or UO_368 (O_368,N_9994,N_9961);
nor UO_369 (O_369,N_9988,N_9928);
or UO_370 (O_370,N_9907,N_9997);
nand UO_371 (O_371,N_9915,N_9903);
nor UO_372 (O_372,N_9931,N_9948);
nor UO_373 (O_373,N_9983,N_9965);
nand UO_374 (O_374,N_9973,N_9980);
nand UO_375 (O_375,N_9999,N_9985);
nand UO_376 (O_376,N_9970,N_9989);
nor UO_377 (O_377,N_9954,N_9905);
nand UO_378 (O_378,N_9913,N_9946);
nor UO_379 (O_379,N_9958,N_9928);
xnor UO_380 (O_380,N_9993,N_9900);
and UO_381 (O_381,N_9920,N_9980);
nor UO_382 (O_382,N_9986,N_9944);
nand UO_383 (O_383,N_9907,N_9936);
nand UO_384 (O_384,N_9938,N_9992);
nor UO_385 (O_385,N_9924,N_9949);
xnor UO_386 (O_386,N_9992,N_9986);
nand UO_387 (O_387,N_9983,N_9971);
or UO_388 (O_388,N_9910,N_9968);
nand UO_389 (O_389,N_9977,N_9912);
and UO_390 (O_390,N_9990,N_9982);
or UO_391 (O_391,N_9966,N_9915);
nor UO_392 (O_392,N_9969,N_9960);
nor UO_393 (O_393,N_9979,N_9947);
xnor UO_394 (O_394,N_9938,N_9926);
nand UO_395 (O_395,N_9907,N_9931);
xnor UO_396 (O_396,N_9910,N_9931);
nand UO_397 (O_397,N_9913,N_9969);
nand UO_398 (O_398,N_9953,N_9964);
and UO_399 (O_399,N_9904,N_9969);
xor UO_400 (O_400,N_9914,N_9946);
xor UO_401 (O_401,N_9984,N_9933);
nand UO_402 (O_402,N_9983,N_9939);
and UO_403 (O_403,N_9905,N_9911);
or UO_404 (O_404,N_9934,N_9988);
or UO_405 (O_405,N_9959,N_9975);
or UO_406 (O_406,N_9925,N_9960);
and UO_407 (O_407,N_9986,N_9972);
or UO_408 (O_408,N_9969,N_9914);
nor UO_409 (O_409,N_9922,N_9978);
nand UO_410 (O_410,N_9905,N_9963);
nor UO_411 (O_411,N_9942,N_9955);
nand UO_412 (O_412,N_9907,N_9986);
and UO_413 (O_413,N_9921,N_9957);
and UO_414 (O_414,N_9951,N_9993);
xor UO_415 (O_415,N_9991,N_9983);
and UO_416 (O_416,N_9907,N_9954);
and UO_417 (O_417,N_9920,N_9903);
xor UO_418 (O_418,N_9994,N_9982);
and UO_419 (O_419,N_9937,N_9929);
or UO_420 (O_420,N_9969,N_9995);
nor UO_421 (O_421,N_9948,N_9908);
xor UO_422 (O_422,N_9977,N_9947);
nand UO_423 (O_423,N_9958,N_9968);
nand UO_424 (O_424,N_9950,N_9988);
or UO_425 (O_425,N_9956,N_9973);
xor UO_426 (O_426,N_9948,N_9902);
xor UO_427 (O_427,N_9996,N_9906);
or UO_428 (O_428,N_9934,N_9989);
nand UO_429 (O_429,N_9934,N_9908);
xor UO_430 (O_430,N_9915,N_9982);
or UO_431 (O_431,N_9948,N_9914);
and UO_432 (O_432,N_9985,N_9975);
xor UO_433 (O_433,N_9903,N_9933);
xor UO_434 (O_434,N_9929,N_9976);
xor UO_435 (O_435,N_9955,N_9948);
nand UO_436 (O_436,N_9979,N_9971);
nand UO_437 (O_437,N_9902,N_9917);
and UO_438 (O_438,N_9933,N_9905);
or UO_439 (O_439,N_9971,N_9931);
or UO_440 (O_440,N_9996,N_9930);
and UO_441 (O_441,N_9941,N_9919);
xor UO_442 (O_442,N_9950,N_9967);
or UO_443 (O_443,N_9925,N_9953);
xnor UO_444 (O_444,N_9975,N_9946);
and UO_445 (O_445,N_9908,N_9915);
xnor UO_446 (O_446,N_9925,N_9997);
nand UO_447 (O_447,N_9952,N_9900);
nor UO_448 (O_448,N_9941,N_9926);
nor UO_449 (O_449,N_9945,N_9987);
xnor UO_450 (O_450,N_9944,N_9943);
and UO_451 (O_451,N_9972,N_9957);
or UO_452 (O_452,N_9989,N_9907);
or UO_453 (O_453,N_9993,N_9982);
nor UO_454 (O_454,N_9934,N_9955);
xnor UO_455 (O_455,N_9959,N_9913);
nand UO_456 (O_456,N_9922,N_9983);
or UO_457 (O_457,N_9937,N_9923);
and UO_458 (O_458,N_9955,N_9977);
xor UO_459 (O_459,N_9902,N_9912);
and UO_460 (O_460,N_9951,N_9988);
or UO_461 (O_461,N_9901,N_9952);
nor UO_462 (O_462,N_9991,N_9997);
and UO_463 (O_463,N_9968,N_9946);
or UO_464 (O_464,N_9958,N_9959);
or UO_465 (O_465,N_9991,N_9989);
and UO_466 (O_466,N_9998,N_9964);
xnor UO_467 (O_467,N_9904,N_9926);
and UO_468 (O_468,N_9982,N_9970);
nand UO_469 (O_469,N_9980,N_9905);
nand UO_470 (O_470,N_9900,N_9923);
or UO_471 (O_471,N_9950,N_9958);
or UO_472 (O_472,N_9931,N_9967);
nand UO_473 (O_473,N_9983,N_9935);
xor UO_474 (O_474,N_9957,N_9989);
nor UO_475 (O_475,N_9968,N_9913);
nand UO_476 (O_476,N_9944,N_9903);
and UO_477 (O_477,N_9939,N_9978);
xor UO_478 (O_478,N_9979,N_9915);
or UO_479 (O_479,N_9925,N_9905);
and UO_480 (O_480,N_9972,N_9911);
or UO_481 (O_481,N_9978,N_9998);
nand UO_482 (O_482,N_9941,N_9985);
nor UO_483 (O_483,N_9978,N_9983);
nor UO_484 (O_484,N_9970,N_9917);
xor UO_485 (O_485,N_9975,N_9939);
xnor UO_486 (O_486,N_9924,N_9994);
and UO_487 (O_487,N_9932,N_9911);
and UO_488 (O_488,N_9990,N_9966);
and UO_489 (O_489,N_9941,N_9940);
and UO_490 (O_490,N_9985,N_9973);
nor UO_491 (O_491,N_9933,N_9950);
nand UO_492 (O_492,N_9911,N_9933);
nor UO_493 (O_493,N_9928,N_9965);
nor UO_494 (O_494,N_9965,N_9916);
nor UO_495 (O_495,N_9975,N_9954);
and UO_496 (O_496,N_9970,N_9961);
and UO_497 (O_497,N_9973,N_9975);
and UO_498 (O_498,N_9973,N_9977);
xor UO_499 (O_499,N_9974,N_9912);
xnor UO_500 (O_500,N_9936,N_9910);
or UO_501 (O_501,N_9976,N_9980);
nand UO_502 (O_502,N_9998,N_9992);
nor UO_503 (O_503,N_9921,N_9958);
nand UO_504 (O_504,N_9957,N_9918);
nor UO_505 (O_505,N_9921,N_9919);
xor UO_506 (O_506,N_9983,N_9944);
and UO_507 (O_507,N_9948,N_9924);
or UO_508 (O_508,N_9967,N_9904);
nor UO_509 (O_509,N_9961,N_9977);
xnor UO_510 (O_510,N_9969,N_9912);
nand UO_511 (O_511,N_9924,N_9917);
xnor UO_512 (O_512,N_9979,N_9974);
xor UO_513 (O_513,N_9998,N_9949);
nor UO_514 (O_514,N_9995,N_9961);
or UO_515 (O_515,N_9926,N_9921);
nor UO_516 (O_516,N_9929,N_9934);
or UO_517 (O_517,N_9922,N_9968);
xnor UO_518 (O_518,N_9966,N_9995);
and UO_519 (O_519,N_9947,N_9987);
nand UO_520 (O_520,N_9971,N_9910);
xnor UO_521 (O_521,N_9973,N_9997);
and UO_522 (O_522,N_9958,N_9978);
xnor UO_523 (O_523,N_9916,N_9908);
or UO_524 (O_524,N_9927,N_9956);
nor UO_525 (O_525,N_9928,N_9917);
nand UO_526 (O_526,N_9904,N_9961);
nor UO_527 (O_527,N_9920,N_9968);
nand UO_528 (O_528,N_9958,N_9935);
nor UO_529 (O_529,N_9916,N_9966);
nor UO_530 (O_530,N_9999,N_9941);
xor UO_531 (O_531,N_9930,N_9999);
or UO_532 (O_532,N_9914,N_9924);
nand UO_533 (O_533,N_9947,N_9946);
nor UO_534 (O_534,N_9905,N_9996);
nor UO_535 (O_535,N_9946,N_9980);
xnor UO_536 (O_536,N_9967,N_9968);
or UO_537 (O_537,N_9991,N_9941);
or UO_538 (O_538,N_9980,N_9916);
and UO_539 (O_539,N_9913,N_9998);
or UO_540 (O_540,N_9907,N_9925);
xor UO_541 (O_541,N_9993,N_9962);
nor UO_542 (O_542,N_9983,N_9992);
xnor UO_543 (O_543,N_9955,N_9993);
or UO_544 (O_544,N_9998,N_9936);
nor UO_545 (O_545,N_9923,N_9965);
or UO_546 (O_546,N_9945,N_9946);
nor UO_547 (O_547,N_9983,N_9961);
nand UO_548 (O_548,N_9924,N_9969);
nand UO_549 (O_549,N_9988,N_9921);
and UO_550 (O_550,N_9946,N_9984);
or UO_551 (O_551,N_9994,N_9974);
xor UO_552 (O_552,N_9912,N_9953);
or UO_553 (O_553,N_9916,N_9912);
and UO_554 (O_554,N_9925,N_9917);
nand UO_555 (O_555,N_9944,N_9917);
xor UO_556 (O_556,N_9990,N_9908);
nor UO_557 (O_557,N_9917,N_9992);
or UO_558 (O_558,N_9980,N_9993);
xnor UO_559 (O_559,N_9904,N_9970);
xor UO_560 (O_560,N_9941,N_9988);
nor UO_561 (O_561,N_9982,N_9935);
nand UO_562 (O_562,N_9939,N_9901);
and UO_563 (O_563,N_9984,N_9995);
or UO_564 (O_564,N_9918,N_9996);
nand UO_565 (O_565,N_9953,N_9970);
xnor UO_566 (O_566,N_9913,N_9905);
or UO_567 (O_567,N_9917,N_9932);
xnor UO_568 (O_568,N_9946,N_9908);
and UO_569 (O_569,N_9982,N_9977);
or UO_570 (O_570,N_9940,N_9931);
and UO_571 (O_571,N_9967,N_9955);
xnor UO_572 (O_572,N_9945,N_9904);
or UO_573 (O_573,N_9937,N_9934);
or UO_574 (O_574,N_9938,N_9996);
nor UO_575 (O_575,N_9907,N_9933);
or UO_576 (O_576,N_9970,N_9903);
nand UO_577 (O_577,N_9958,N_9986);
nand UO_578 (O_578,N_9979,N_9911);
nand UO_579 (O_579,N_9900,N_9931);
nand UO_580 (O_580,N_9909,N_9954);
nor UO_581 (O_581,N_9960,N_9924);
nor UO_582 (O_582,N_9979,N_9905);
or UO_583 (O_583,N_9973,N_9937);
or UO_584 (O_584,N_9944,N_9942);
xor UO_585 (O_585,N_9997,N_9948);
or UO_586 (O_586,N_9998,N_9906);
xnor UO_587 (O_587,N_9961,N_9901);
xnor UO_588 (O_588,N_9932,N_9960);
or UO_589 (O_589,N_9921,N_9916);
nor UO_590 (O_590,N_9975,N_9974);
and UO_591 (O_591,N_9968,N_9933);
xor UO_592 (O_592,N_9933,N_9967);
nand UO_593 (O_593,N_9990,N_9918);
xor UO_594 (O_594,N_9925,N_9933);
nor UO_595 (O_595,N_9951,N_9980);
xor UO_596 (O_596,N_9902,N_9974);
or UO_597 (O_597,N_9945,N_9971);
nand UO_598 (O_598,N_9920,N_9916);
xnor UO_599 (O_599,N_9955,N_9905);
xor UO_600 (O_600,N_9996,N_9941);
nor UO_601 (O_601,N_9902,N_9931);
nand UO_602 (O_602,N_9986,N_9964);
nand UO_603 (O_603,N_9951,N_9983);
nor UO_604 (O_604,N_9991,N_9919);
or UO_605 (O_605,N_9913,N_9942);
and UO_606 (O_606,N_9935,N_9972);
nand UO_607 (O_607,N_9991,N_9945);
nand UO_608 (O_608,N_9939,N_9955);
and UO_609 (O_609,N_9934,N_9923);
nor UO_610 (O_610,N_9930,N_9972);
nor UO_611 (O_611,N_9941,N_9976);
nor UO_612 (O_612,N_9959,N_9976);
nor UO_613 (O_613,N_9922,N_9934);
nand UO_614 (O_614,N_9982,N_9974);
xnor UO_615 (O_615,N_9977,N_9917);
and UO_616 (O_616,N_9989,N_9986);
xnor UO_617 (O_617,N_9969,N_9963);
nand UO_618 (O_618,N_9951,N_9949);
and UO_619 (O_619,N_9946,N_9949);
nor UO_620 (O_620,N_9984,N_9955);
and UO_621 (O_621,N_9929,N_9962);
nor UO_622 (O_622,N_9921,N_9984);
nor UO_623 (O_623,N_9950,N_9947);
nor UO_624 (O_624,N_9914,N_9935);
nor UO_625 (O_625,N_9992,N_9935);
or UO_626 (O_626,N_9974,N_9950);
and UO_627 (O_627,N_9969,N_9976);
nand UO_628 (O_628,N_9954,N_9929);
nand UO_629 (O_629,N_9955,N_9904);
and UO_630 (O_630,N_9911,N_9942);
or UO_631 (O_631,N_9909,N_9906);
and UO_632 (O_632,N_9914,N_9983);
xnor UO_633 (O_633,N_9940,N_9962);
and UO_634 (O_634,N_9913,N_9903);
xor UO_635 (O_635,N_9930,N_9965);
and UO_636 (O_636,N_9915,N_9913);
nand UO_637 (O_637,N_9949,N_9936);
nor UO_638 (O_638,N_9968,N_9983);
nand UO_639 (O_639,N_9918,N_9967);
and UO_640 (O_640,N_9988,N_9969);
nor UO_641 (O_641,N_9902,N_9987);
or UO_642 (O_642,N_9907,N_9901);
and UO_643 (O_643,N_9991,N_9908);
and UO_644 (O_644,N_9936,N_9934);
or UO_645 (O_645,N_9958,N_9900);
xnor UO_646 (O_646,N_9972,N_9956);
or UO_647 (O_647,N_9996,N_9956);
and UO_648 (O_648,N_9939,N_9911);
nor UO_649 (O_649,N_9959,N_9951);
and UO_650 (O_650,N_9935,N_9939);
nor UO_651 (O_651,N_9934,N_9992);
or UO_652 (O_652,N_9984,N_9969);
xor UO_653 (O_653,N_9992,N_9994);
xnor UO_654 (O_654,N_9928,N_9969);
xnor UO_655 (O_655,N_9924,N_9990);
nand UO_656 (O_656,N_9956,N_9925);
nor UO_657 (O_657,N_9946,N_9981);
and UO_658 (O_658,N_9916,N_9907);
and UO_659 (O_659,N_9908,N_9941);
xnor UO_660 (O_660,N_9928,N_9963);
or UO_661 (O_661,N_9965,N_9971);
nor UO_662 (O_662,N_9958,N_9983);
xor UO_663 (O_663,N_9955,N_9961);
or UO_664 (O_664,N_9939,N_9932);
or UO_665 (O_665,N_9956,N_9904);
or UO_666 (O_666,N_9989,N_9963);
nor UO_667 (O_667,N_9924,N_9937);
nand UO_668 (O_668,N_9994,N_9955);
and UO_669 (O_669,N_9931,N_9960);
nor UO_670 (O_670,N_9988,N_9931);
nor UO_671 (O_671,N_9925,N_9970);
or UO_672 (O_672,N_9953,N_9972);
nand UO_673 (O_673,N_9963,N_9901);
or UO_674 (O_674,N_9916,N_9945);
or UO_675 (O_675,N_9901,N_9945);
and UO_676 (O_676,N_9936,N_9952);
nand UO_677 (O_677,N_9948,N_9933);
nor UO_678 (O_678,N_9915,N_9937);
nor UO_679 (O_679,N_9955,N_9975);
and UO_680 (O_680,N_9981,N_9927);
or UO_681 (O_681,N_9977,N_9916);
or UO_682 (O_682,N_9986,N_9991);
and UO_683 (O_683,N_9971,N_9904);
and UO_684 (O_684,N_9973,N_9991);
nand UO_685 (O_685,N_9935,N_9996);
nand UO_686 (O_686,N_9944,N_9976);
xnor UO_687 (O_687,N_9908,N_9971);
xnor UO_688 (O_688,N_9997,N_9965);
and UO_689 (O_689,N_9965,N_9988);
xnor UO_690 (O_690,N_9930,N_9908);
nor UO_691 (O_691,N_9945,N_9943);
nand UO_692 (O_692,N_9970,N_9922);
nor UO_693 (O_693,N_9999,N_9970);
nand UO_694 (O_694,N_9986,N_9998);
or UO_695 (O_695,N_9991,N_9946);
or UO_696 (O_696,N_9962,N_9933);
xnor UO_697 (O_697,N_9958,N_9931);
xnor UO_698 (O_698,N_9941,N_9946);
nand UO_699 (O_699,N_9904,N_9943);
or UO_700 (O_700,N_9967,N_9902);
and UO_701 (O_701,N_9994,N_9912);
xor UO_702 (O_702,N_9911,N_9948);
xnor UO_703 (O_703,N_9904,N_9978);
nor UO_704 (O_704,N_9957,N_9931);
nor UO_705 (O_705,N_9927,N_9959);
or UO_706 (O_706,N_9976,N_9910);
or UO_707 (O_707,N_9990,N_9933);
and UO_708 (O_708,N_9992,N_9999);
or UO_709 (O_709,N_9931,N_9946);
or UO_710 (O_710,N_9945,N_9950);
and UO_711 (O_711,N_9960,N_9999);
nor UO_712 (O_712,N_9924,N_9982);
nor UO_713 (O_713,N_9939,N_9945);
and UO_714 (O_714,N_9927,N_9908);
nand UO_715 (O_715,N_9915,N_9953);
or UO_716 (O_716,N_9905,N_9957);
xnor UO_717 (O_717,N_9903,N_9952);
nand UO_718 (O_718,N_9905,N_9992);
or UO_719 (O_719,N_9978,N_9923);
nand UO_720 (O_720,N_9944,N_9934);
nand UO_721 (O_721,N_9981,N_9995);
nand UO_722 (O_722,N_9908,N_9994);
nand UO_723 (O_723,N_9993,N_9938);
or UO_724 (O_724,N_9984,N_9944);
and UO_725 (O_725,N_9972,N_9958);
and UO_726 (O_726,N_9932,N_9989);
and UO_727 (O_727,N_9938,N_9950);
nand UO_728 (O_728,N_9997,N_9909);
nor UO_729 (O_729,N_9992,N_9981);
or UO_730 (O_730,N_9912,N_9915);
or UO_731 (O_731,N_9938,N_9908);
or UO_732 (O_732,N_9929,N_9939);
or UO_733 (O_733,N_9942,N_9907);
xor UO_734 (O_734,N_9989,N_9926);
and UO_735 (O_735,N_9948,N_9918);
and UO_736 (O_736,N_9993,N_9925);
or UO_737 (O_737,N_9915,N_9976);
or UO_738 (O_738,N_9955,N_9983);
and UO_739 (O_739,N_9976,N_9914);
and UO_740 (O_740,N_9956,N_9909);
xor UO_741 (O_741,N_9966,N_9964);
and UO_742 (O_742,N_9928,N_9979);
xor UO_743 (O_743,N_9921,N_9951);
or UO_744 (O_744,N_9988,N_9961);
xor UO_745 (O_745,N_9994,N_9967);
nor UO_746 (O_746,N_9936,N_9959);
nand UO_747 (O_747,N_9935,N_9934);
or UO_748 (O_748,N_9982,N_9987);
nor UO_749 (O_749,N_9985,N_9967);
xnor UO_750 (O_750,N_9962,N_9908);
nor UO_751 (O_751,N_9943,N_9935);
and UO_752 (O_752,N_9902,N_9993);
xnor UO_753 (O_753,N_9967,N_9963);
and UO_754 (O_754,N_9991,N_9907);
and UO_755 (O_755,N_9975,N_9984);
and UO_756 (O_756,N_9993,N_9984);
or UO_757 (O_757,N_9984,N_9923);
nor UO_758 (O_758,N_9993,N_9932);
nand UO_759 (O_759,N_9966,N_9984);
and UO_760 (O_760,N_9910,N_9960);
and UO_761 (O_761,N_9998,N_9952);
nand UO_762 (O_762,N_9972,N_9947);
or UO_763 (O_763,N_9935,N_9919);
or UO_764 (O_764,N_9968,N_9955);
nand UO_765 (O_765,N_9955,N_9943);
and UO_766 (O_766,N_9984,N_9904);
xor UO_767 (O_767,N_9919,N_9916);
and UO_768 (O_768,N_9955,N_9918);
and UO_769 (O_769,N_9981,N_9903);
and UO_770 (O_770,N_9963,N_9906);
nor UO_771 (O_771,N_9919,N_9922);
or UO_772 (O_772,N_9964,N_9984);
xor UO_773 (O_773,N_9991,N_9982);
and UO_774 (O_774,N_9993,N_9905);
nand UO_775 (O_775,N_9920,N_9961);
xnor UO_776 (O_776,N_9918,N_9936);
and UO_777 (O_777,N_9974,N_9949);
and UO_778 (O_778,N_9949,N_9901);
nor UO_779 (O_779,N_9965,N_9951);
nand UO_780 (O_780,N_9987,N_9983);
nor UO_781 (O_781,N_9915,N_9932);
and UO_782 (O_782,N_9909,N_9917);
nand UO_783 (O_783,N_9996,N_9971);
or UO_784 (O_784,N_9916,N_9962);
or UO_785 (O_785,N_9979,N_9962);
nand UO_786 (O_786,N_9993,N_9908);
xor UO_787 (O_787,N_9926,N_9966);
and UO_788 (O_788,N_9934,N_9921);
xnor UO_789 (O_789,N_9974,N_9980);
nor UO_790 (O_790,N_9972,N_9925);
nand UO_791 (O_791,N_9976,N_9992);
xor UO_792 (O_792,N_9996,N_9925);
nand UO_793 (O_793,N_9985,N_9916);
and UO_794 (O_794,N_9993,N_9974);
and UO_795 (O_795,N_9922,N_9981);
xnor UO_796 (O_796,N_9965,N_9966);
and UO_797 (O_797,N_9921,N_9969);
nor UO_798 (O_798,N_9947,N_9959);
or UO_799 (O_799,N_9991,N_9955);
nand UO_800 (O_800,N_9930,N_9995);
and UO_801 (O_801,N_9967,N_9958);
and UO_802 (O_802,N_9929,N_9995);
nand UO_803 (O_803,N_9928,N_9904);
nand UO_804 (O_804,N_9917,N_9942);
xnor UO_805 (O_805,N_9949,N_9981);
nor UO_806 (O_806,N_9987,N_9929);
nand UO_807 (O_807,N_9922,N_9992);
xnor UO_808 (O_808,N_9910,N_9933);
nor UO_809 (O_809,N_9963,N_9927);
xnor UO_810 (O_810,N_9992,N_9947);
or UO_811 (O_811,N_9916,N_9979);
nor UO_812 (O_812,N_9957,N_9998);
and UO_813 (O_813,N_9967,N_9944);
and UO_814 (O_814,N_9966,N_9923);
xnor UO_815 (O_815,N_9946,N_9920);
xor UO_816 (O_816,N_9924,N_9975);
nor UO_817 (O_817,N_9967,N_9941);
or UO_818 (O_818,N_9936,N_9994);
nor UO_819 (O_819,N_9928,N_9902);
xnor UO_820 (O_820,N_9939,N_9959);
and UO_821 (O_821,N_9929,N_9932);
or UO_822 (O_822,N_9959,N_9995);
nor UO_823 (O_823,N_9928,N_9943);
and UO_824 (O_824,N_9938,N_9941);
xor UO_825 (O_825,N_9934,N_9958);
nand UO_826 (O_826,N_9978,N_9924);
nor UO_827 (O_827,N_9970,N_9951);
nor UO_828 (O_828,N_9942,N_9905);
nor UO_829 (O_829,N_9991,N_9975);
xor UO_830 (O_830,N_9932,N_9983);
nand UO_831 (O_831,N_9966,N_9963);
nand UO_832 (O_832,N_9924,N_9916);
or UO_833 (O_833,N_9991,N_9963);
nand UO_834 (O_834,N_9946,N_9938);
or UO_835 (O_835,N_9923,N_9950);
or UO_836 (O_836,N_9925,N_9968);
and UO_837 (O_837,N_9964,N_9960);
nor UO_838 (O_838,N_9976,N_9972);
xor UO_839 (O_839,N_9985,N_9954);
nand UO_840 (O_840,N_9973,N_9990);
and UO_841 (O_841,N_9928,N_9994);
and UO_842 (O_842,N_9908,N_9907);
nand UO_843 (O_843,N_9943,N_9915);
xor UO_844 (O_844,N_9908,N_9979);
nand UO_845 (O_845,N_9979,N_9935);
xor UO_846 (O_846,N_9910,N_9962);
and UO_847 (O_847,N_9930,N_9926);
nor UO_848 (O_848,N_9963,N_9951);
nand UO_849 (O_849,N_9939,N_9968);
nor UO_850 (O_850,N_9945,N_9994);
nor UO_851 (O_851,N_9909,N_9910);
xor UO_852 (O_852,N_9925,N_9943);
or UO_853 (O_853,N_9972,N_9904);
nand UO_854 (O_854,N_9919,N_9903);
nor UO_855 (O_855,N_9918,N_9941);
nor UO_856 (O_856,N_9906,N_9900);
and UO_857 (O_857,N_9933,N_9961);
and UO_858 (O_858,N_9947,N_9909);
and UO_859 (O_859,N_9935,N_9904);
nor UO_860 (O_860,N_9930,N_9958);
or UO_861 (O_861,N_9913,N_9996);
nand UO_862 (O_862,N_9994,N_9947);
and UO_863 (O_863,N_9989,N_9987);
xor UO_864 (O_864,N_9934,N_9925);
xor UO_865 (O_865,N_9913,N_9976);
nand UO_866 (O_866,N_9902,N_9996);
xor UO_867 (O_867,N_9929,N_9982);
xnor UO_868 (O_868,N_9998,N_9944);
and UO_869 (O_869,N_9901,N_9982);
xor UO_870 (O_870,N_9909,N_9939);
nand UO_871 (O_871,N_9970,N_9960);
and UO_872 (O_872,N_9999,N_9931);
xnor UO_873 (O_873,N_9929,N_9915);
nor UO_874 (O_874,N_9964,N_9979);
or UO_875 (O_875,N_9917,N_9974);
or UO_876 (O_876,N_9943,N_9985);
or UO_877 (O_877,N_9986,N_9969);
xor UO_878 (O_878,N_9923,N_9959);
or UO_879 (O_879,N_9931,N_9970);
or UO_880 (O_880,N_9984,N_9931);
or UO_881 (O_881,N_9927,N_9930);
or UO_882 (O_882,N_9916,N_9967);
nand UO_883 (O_883,N_9957,N_9993);
or UO_884 (O_884,N_9933,N_9938);
or UO_885 (O_885,N_9935,N_9995);
nand UO_886 (O_886,N_9950,N_9934);
and UO_887 (O_887,N_9937,N_9936);
nand UO_888 (O_888,N_9938,N_9901);
or UO_889 (O_889,N_9939,N_9943);
nand UO_890 (O_890,N_9924,N_9954);
or UO_891 (O_891,N_9987,N_9977);
and UO_892 (O_892,N_9924,N_9983);
nand UO_893 (O_893,N_9975,N_9952);
xnor UO_894 (O_894,N_9911,N_9908);
nand UO_895 (O_895,N_9975,N_9905);
or UO_896 (O_896,N_9943,N_9982);
nand UO_897 (O_897,N_9962,N_9998);
nand UO_898 (O_898,N_9942,N_9974);
xor UO_899 (O_899,N_9981,N_9970);
and UO_900 (O_900,N_9967,N_9946);
nand UO_901 (O_901,N_9962,N_9982);
xnor UO_902 (O_902,N_9966,N_9906);
xor UO_903 (O_903,N_9912,N_9904);
and UO_904 (O_904,N_9907,N_9953);
nor UO_905 (O_905,N_9929,N_9927);
or UO_906 (O_906,N_9968,N_9952);
and UO_907 (O_907,N_9944,N_9963);
and UO_908 (O_908,N_9919,N_9951);
or UO_909 (O_909,N_9995,N_9952);
xor UO_910 (O_910,N_9923,N_9901);
or UO_911 (O_911,N_9935,N_9924);
nor UO_912 (O_912,N_9988,N_9987);
xnor UO_913 (O_913,N_9926,N_9905);
nand UO_914 (O_914,N_9941,N_9949);
or UO_915 (O_915,N_9914,N_9954);
or UO_916 (O_916,N_9979,N_9945);
nor UO_917 (O_917,N_9905,N_9938);
or UO_918 (O_918,N_9970,N_9962);
xnor UO_919 (O_919,N_9990,N_9970);
nor UO_920 (O_920,N_9999,N_9972);
and UO_921 (O_921,N_9981,N_9957);
nand UO_922 (O_922,N_9922,N_9930);
nand UO_923 (O_923,N_9903,N_9906);
xnor UO_924 (O_924,N_9912,N_9917);
and UO_925 (O_925,N_9918,N_9902);
and UO_926 (O_926,N_9989,N_9903);
nand UO_927 (O_927,N_9943,N_9938);
nand UO_928 (O_928,N_9949,N_9975);
and UO_929 (O_929,N_9998,N_9972);
or UO_930 (O_930,N_9982,N_9938);
xnor UO_931 (O_931,N_9986,N_9957);
nand UO_932 (O_932,N_9971,N_9925);
xnor UO_933 (O_933,N_9975,N_9986);
and UO_934 (O_934,N_9961,N_9932);
xor UO_935 (O_935,N_9960,N_9997);
nand UO_936 (O_936,N_9935,N_9956);
or UO_937 (O_937,N_9953,N_9974);
and UO_938 (O_938,N_9981,N_9974);
xnor UO_939 (O_939,N_9946,N_9976);
xnor UO_940 (O_940,N_9985,N_9979);
or UO_941 (O_941,N_9976,N_9958);
nor UO_942 (O_942,N_9994,N_9956);
nand UO_943 (O_943,N_9955,N_9935);
and UO_944 (O_944,N_9998,N_9910);
nor UO_945 (O_945,N_9976,N_9956);
xor UO_946 (O_946,N_9951,N_9912);
or UO_947 (O_947,N_9954,N_9951);
nand UO_948 (O_948,N_9940,N_9911);
nand UO_949 (O_949,N_9997,N_9953);
or UO_950 (O_950,N_9974,N_9920);
nor UO_951 (O_951,N_9916,N_9915);
nand UO_952 (O_952,N_9957,N_9926);
nor UO_953 (O_953,N_9996,N_9986);
xnor UO_954 (O_954,N_9967,N_9949);
nand UO_955 (O_955,N_9977,N_9921);
xor UO_956 (O_956,N_9938,N_9962);
xnor UO_957 (O_957,N_9902,N_9914);
nor UO_958 (O_958,N_9964,N_9978);
nand UO_959 (O_959,N_9933,N_9936);
nor UO_960 (O_960,N_9995,N_9982);
xnor UO_961 (O_961,N_9995,N_9970);
and UO_962 (O_962,N_9914,N_9997);
or UO_963 (O_963,N_9958,N_9999);
nor UO_964 (O_964,N_9974,N_9978);
or UO_965 (O_965,N_9909,N_9903);
nor UO_966 (O_966,N_9948,N_9917);
xnor UO_967 (O_967,N_9940,N_9989);
nand UO_968 (O_968,N_9940,N_9925);
and UO_969 (O_969,N_9910,N_9979);
or UO_970 (O_970,N_9916,N_9999);
nor UO_971 (O_971,N_9989,N_9983);
and UO_972 (O_972,N_9910,N_9926);
nor UO_973 (O_973,N_9941,N_9915);
nand UO_974 (O_974,N_9928,N_9936);
nor UO_975 (O_975,N_9934,N_9941);
or UO_976 (O_976,N_9981,N_9926);
xnor UO_977 (O_977,N_9912,N_9958);
or UO_978 (O_978,N_9951,N_9950);
or UO_979 (O_979,N_9956,N_9950);
nand UO_980 (O_980,N_9909,N_9957);
nand UO_981 (O_981,N_9948,N_9951);
xnor UO_982 (O_982,N_9940,N_9945);
and UO_983 (O_983,N_9911,N_9930);
nand UO_984 (O_984,N_9917,N_9914);
nor UO_985 (O_985,N_9980,N_9928);
nand UO_986 (O_986,N_9904,N_9921);
or UO_987 (O_987,N_9954,N_9945);
and UO_988 (O_988,N_9950,N_9913);
or UO_989 (O_989,N_9937,N_9951);
nor UO_990 (O_990,N_9962,N_9939);
nand UO_991 (O_991,N_9945,N_9949);
nand UO_992 (O_992,N_9970,N_9928);
nor UO_993 (O_993,N_9962,N_9973);
and UO_994 (O_994,N_9961,N_9948);
nor UO_995 (O_995,N_9928,N_9942);
nor UO_996 (O_996,N_9933,N_9957);
nand UO_997 (O_997,N_9917,N_9905);
xor UO_998 (O_998,N_9924,N_9992);
nand UO_999 (O_999,N_9921,N_9994);
or UO_1000 (O_1000,N_9997,N_9943);
nand UO_1001 (O_1001,N_9971,N_9927);
or UO_1002 (O_1002,N_9915,N_9940);
or UO_1003 (O_1003,N_9923,N_9979);
or UO_1004 (O_1004,N_9915,N_9975);
nor UO_1005 (O_1005,N_9966,N_9980);
nor UO_1006 (O_1006,N_9979,N_9919);
nor UO_1007 (O_1007,N_9969,N_9927);
xnor UO_1008 (O_1008,N_9901,N_9950);
and UO_1009 (O_1009,N_9970,N_9941);
nor UO_1010 (O_1010,N_9962,N_9971);
nand UO_1011 (O_1011,N_9982,N_9996);
nand UO_1012 (O_1012,N_9991,N_9953);
nor UO_1013 (O_1013,N_9964,N_9963);
or UO_1014 (O_1014,N_9901,N_9918);
and UO_1015 (O_1015,N_9966,N_9941);
or UO_1016 (O_1016,N_9958,N_9916);
nor UO_1017 (O_1017,N_9949,N_9908);
xor UO_1018 (O_1018,N_9983,N_9940);
or UO_1019 (O_1019,N_9919,N_9926);
and UO_1020 (O_1020,N_9945,N_9980);
xnor UO_1021 (O_1021,N_9921,N_9968);
xnor UO_1022 (O_1022,N_9922,N_9927);
and UO_1023 (O_1023,N_9987,N_9934);
nand UO_1024 (O_1024,N_9973,N_9953);
or UO_1025 (O_1025,N_9977,N_9985);
or UO_1026 (O_1026,N_9926,N_9978);
and UO_1027 (O_1027,N_9961,N_9907);
nand UO_1028 (O_1028,N_9918,N_9914);
nor UO_1029 (O_1029,N_9988,N_9943);
nand UO_1030 (O_1030,N_9990,N_9901);
nor UO_1031 (O_1031,N_9999,N_9906);
nand UO_1032 (O_1032,N_9949,N_9964);
or UO_1033 (O_1033,N_9981,N_9930);
nor UO_1034 (O_1034,N_9920,N_9956);
and UO_1035 (O_1035,N_9978,N_9971);
and UO_1036 (O_1036,N_9991,N_9961);
nand UO_1037 (O_1037,N_9965,N_9958);
or UO_1038 (O_1038,N_9982,N_9932);
nand UO_1039 (O_1039,N_9952,N_9990);
nor UO_1040 (O_1040,N_9929,N_9984);
xor UO_1041 (O_1041,N_9901,N_9983);
nand UO_1042 (O_1042,N_9942,N_9987);
or UO_1043 (O_1043,N_9952,N_9989);
nor UO_1044 (O_1044,N_9961,N_9985);
or UO_1045 (O_1045,N_9920,N_9938);
and UO_1046 (O_1046,N_9994,N_9954);
and UO_1047 (O_1047,N_9928,N_9973);
xnor UO_1048 (O_1048,N_9930,N_9939);
xnor UO_1049 (O_1049,N_9992,N_9961);
nor UO_1050 (O_1050,N_9974,N_9900);
xnor UO_1051 (O_1051,N_9956,N_9978);
or UO_1052 (O_1052,N_9912,N_9956);
or UO_1053 (O_1053,N_9901,N_9972);
nand UO_1054 (O_1054,N_9993,N_9979);
nand UO_1055 (O_1055,N_9945,N_9928);
nor UO_1056 (O_1056,N_9921,N_9912);
nand UO_1057 (O_1057,N_9995,N_9908);
xor UO_1058 (O_1058,N_9987,N_9952);
nand UO_1059 (O_1059,N_9967,N_9948);
or UO_1060 (O_1060,N_9967,N_9960);
or UO_1061 (O_1061,N_9906,N_9929);
xor UO_1062 (O_1062,N_9982,N_9949);
and UO_1063 (O_1063,N_9917,N_9939);
nand UO_1064 (O_1064,N_9901,N_9912);
xnor UO_1065 (O_1065,N_9965,N_9914);
and UO_1066 (O_1066,N_9954,N_9926);
or UO_1067 (O_1067,N_9975,N_9941);
nor UO_1068 (O_1068,N_9939,N_9976);
xnor UO_1069 (O_1069,N_9935,N_9945);
or UO_1070 (O_1070,N_9964,N_9913);
and UO_1071 (O_1071,N_9937,N_9971);
and UO_1072 (O_1072,N_9920,N_9943);
or UO_1073 (O_1073,N_9974,N_9935);
or UO_1074 (O_1074,N_9999,N_9962);
or UO_1075 (O_1075,N_9938,N_9902);
or UO_1076 (O_1076,N_9948,N_9937);
nand UO_1077 (O_1077,N_9935,N_9975);
xnor UO_1078 (O_1078,N_9964,N_9944);
nand UO_1079 (O_1079,N_9959,N_9910);
and UO_1080 (O_1080,N_9975,N_9990);
and UO_1081 (O_1081,N_9973,N_9969);
nor UO_1082 (O_1082,N_9911,N_9928);
nand UO_1083 (O_1083,N_9918,N_9994);
or UO_1084 (O_1084,N_9958,N_9942);
nor UO_1085 (O_1085,N_9970,N_9980);
nand UO_1086 (O_1086,N_9906,N_9955);
and UO_1087 (O_1087,N_9974,N_9963);
nor UO_1088 (O_1088,N_9958,N_9902);
or UO_1089 (O_1089,N_9919,N_9942);
and UO_1090 (O_1090,N_9919,N_9973);
or UO_1091 (O_1091,N_9940,N_9914);
nand UO_1092 (O_1092,N_9974,N_9984);
nand UO_1093 (O_1093,N_9985,N_9934);
nor UO_1094 (O_1094,N_9914,N_9967);
and UO_1095 (O_1095,N_9984,N_9912);
xor UO_1096 (O_1096,N_9926,N_9982);
and UO_1097 (O_1097,N_9969,N_9964);
nor UO_1098 (O_1098,N_9970,N_9934);
nand UO_1099 (O_1099,N_9988,N_9975);
nor UO_1100 (O_1100,N_9995,N_9957);
or UO_1101 (O_1101,N_9936,N_9990);
and UO_1102 (O_1102,N_9982,N_9979);
and UO_1103 (O_1103,N_9953,N_9921);
nor UO_1104 (O_1104,N_9997,N_9931);
or UO_1105 (O_1105,N_9957,N_9928);
and UO_1106 (O_1106,N_9906,N_9983);
or UO_1107 (O_1107,N_9975,N_9922);
or UO_1108 (O_1108,N_9977,N_9900);
or UO_1109 (O_1109,N_9957,N_9922);
and UO_1110 (O_1110,N_9907,N_9911);
or UO_1111 (O_1111,N_9987,N_9957);
nor UO_1112 (O_1112,N_9934,N_9902);
nand UO_1113 (O_1113,N_9971,N_9954);
and UO_1114 (O_1114,N_9997,N_9974);
and UO_1115 (O_1115,N_9938,N_9925);
nor UO_1116 (O_1116,N_9949,N_9971);
xor UO_1117 (O_1117,N_9935,N_9947);
or UO_1118 (O_1118,N_9980,N_9992);
nor UO_1119 (O_1119,N_9913,N_9919);
and UO_1120 (O_1120,N_9914,N_9951);
nand UO_1121 (O_1121,N_9925,N_9959);
nand UO_1122 (O_1122,N_9993,N_9978);
nand UO_1123 (O_1123,N_9917,N_9906);
nor UO_1124 (O_1124,N_9978,N_9911);
and UO_1125 (O_1125,N_9928,N_9995);
nor UO_1126 (O_1126,N_9948,N_9904);
and UO_1127 (O_1127,N_9907,N_9985);
or UO_1128 (O_1128,N_9903,N_9993);
or UO_1129 (O_1129,N_9980,N_9968);
and UO_1130 (O_1130,N_9936,N_9964);
xnor UO_1131 (O_1131,N_9988,N_9973);
nor UO_1132 (O_1132,N_9993,N_9952);
xnor UO_1133 (O_1133,N_9953,N_9926);
or UO_1134 (O_1134,N_9960,N_9958);
or UO_1135 (O_1135,N_9904,N_9925);
nand UO_1136 (O_1136,N_9941,N_9911);
nand UO_1137 (O_1137,N_9920,N_9901);
nand UO_1138 (O_1138,N_9907,N_9948);
or UO_1139 (O_1139,N_9982,N_9908);
or UO_1140 (O_1140,N_9922,N_9974);
nor UO_1141 (O_1141,N_9988,N_9912);
nor UO_1142 (O_1142,N_9941,N_9927);
and UO_1143 (O_1143,N_9952,N_9951);
xor UO_1144 (O_1144,N_9954,N_9956);
or UO_1145 (O_1145,N_9908,N_9965);
xnor UO_1146 (O_1146,N_9999,N_9981);
nand UO_1147 (O_1147,N_9943,N_9946);
or UO_1148 (O_1148,N_9993,N_9942);
and UO_1149 (O_1149,N_9924,N_9931);
or UO_1150 (O_1150,N_9965,N_9975);
nor UO_1151 (O_1151,N_9939,N_9965);
nor UO_1152 (O_1152,N_9963,N_9926);
and UO_1153 (O_1153,N_9917,N_9975);
and UO_1154 (O_1154,N_9920,N_9922);
xnor UO_1155 (O_1155,N_9910,N_9945);
xnor UO_1156 (O_1156,N_9970,N_9997);
xnor UO_1157 (O_1157,N_9951,N_9928);
and UO_1158 (O_1158,N_9957,N_9954);
xor UO_1159 (O_1159,N_9947,N_9976);
or UO_1160 (O_1160,N_9956,N_9989);
xnor UO_1161 (O_1161,N_9981,N_9951);
nand UO_1162 (O_1162,N_9967,N_9957);
and UO_1163 (O_1163,N_9987,N_9995);
and UO_1164 (O_1164,N_9969,N_9958);
nor UO_1165 (O_1165,N_9967,N_9953);
or UO_1166 (O_1166,N_9972,N_9970);
and UO_1167 (O_1167,N_9937,N_9920);
nand UO_1168 (O_1168,N_9978,N_9938);
nand UO_1169 (O_1169,N_9974,N_9916);
xor UO_1170 (O_1170,N_9985,N_9978);
and UO_1171 (O_1171,N_9915,N_9962);
or UO_1172 (O_1172,N_9966,N_9911);
xor UO_1173 (O_1173,N_9999,N_9938);
and UO_1174 (O_1174,N_9990,N_9960);
and UO_1175 (O_1175,N_9938,N_9942);
and UO_1176 (O_1176,N_9902,N_9937);
nand UO_1177 (O_1177,N_9905,N_9920);
or UO_1178 (O_1178,N_9953,N_9942);
nor UO_1179 (O_1179,N_9957,N_9961);
or UO_1180 (O_1180,N_9991,N_9904);
and UO_1181 (O_1181,N_9991,N_9980);
or UO_1182 (O_1182,N_9942,N_9936);
or UO_1183 (O_1183,N_9961,N_9939);
nor UO_1184 (O_1184,N_9957,N_9952);
xor UO_1185 (O_1185,N_9986,N_9916);
nand UO_1186 (O_1186,N_9960,N_9972);
or UO_1187 (O_1187,N_9976,N_9919);
or UO_1188 (O_1188,N_9981,N_9929);
xor UO_1189 (O_1189,N_9996,N_9998);
and UO_1190 (O_1190,N_9945,N_9983);
nor UO_1191 (O_1191,N_9966,N_9992);
and UO_1192 (O_1192,N_9959,N_9922);
and UO_1193 (O_1193,N_9991,N_9976);
nand UO_1194 (O_1194,N_9971,N_9917);
and UO_1195 (O_1195,N_9966,N_9925);
nor UO_1196 (O_1196,N_9956,N_9916);
nand UO_1197 (O_1197,N_9983,N_9916);
nand UO_1198 (O_1198,N_9986,N_9980);
nand UO_1199 (O_1199,N_9950,N_9985);
and UO_1200 (O_1200,N_9946,N_9960);
nor UO_1201 (O_1201,N_9945,N_9961);
and UO_1202 (O_1202,N_9950,N_9983);
nand UO_1203 (O_1203,N_9949,N_9903);
nand UO_1204 (O_1204,N_9971,N_9946);
nor UO_1205 (O_1205,N_9919,N_9906);
nor UO_1206 (O_1206,N_9976,N_9928);
nand UO_1207 (O_1207,N_9924,N_9953);
and UO_1208 (O_1208,N_9954,N_9911);
and UO_1209 (O_1209,N_9999,N_9963);
nor UO_1210 (O_1210,N_9923,N_9952);
xnor UO_1211 (O_1211,N_9913,N_9982);
and UO_1212 (O_1212,N_9926,N_9914);
nor UO_1213 (O_1213,N_9942,N_9946);
nand UO_1214 (O_1214,N_9937,N_9917);
nand UO_1215 (O_1215,N_9903,N_9983);
nand UO_1216 (O_1216,N_9939,N_9949);
nand UO_1217 (O_1217,N_9945,N_9972);
nor UO_1218 (O_1218,N_9923,N_9927);
or UO_1219 (O_1219,N_9988,N_9932);
xor UO_1220 (O_1220,N_9999,N_9990);
and UO_1221 (O_1221,N_9923,N_9920);
or UO_1222 (O_1222,N_9962,N_9936);
and UO_1223 (O_1223,N_9984,N_9951);
and UO_1224 (O_1224,N_9937,N_9907);
or UO_1225 (O_1225,N_9958,N_9943);
xnor UO_1226 (O_1226,N_9954,N_9949);
and UO_1227 (O_1227,N_9957,N_9942);
nor UO_1228 (O_1228,N_9921,N_9932);
and UO_1229 (O_1229,N_9954,N_9933);
nand UO_1230 (O_1230,N_9959,N_9965);
and UO_1231 (O_1231,N_9965,N_9981);
nor UO_1232 (O_1232,N_9947,N_9900);
xnor UO_1233 (O_1233,N_9932,N_9918);
nor UO_1234 (O_1234,N_9987,N_9973);
xor UO_1235 (O_1235,N_9920,N_9967);
xnor UO_1236 (O_1236,N_9978,N_9960);
xnor UO_1237 (O_1237,N_9950,N_9973);
and UO_1238 (O_1238,N_9955,N_9932);
nor UO_1239 (O_1239,N_9974,N_9925);
nand UO_1240 (O_1240,N_9998,N_9916);
nor UO_1241 (O_1241,N_9916,N_9933);
or UO_1242 (O_1242,N_9932,N_9937);
xor UO_1243 (O_1243,N_9954,N_9915);
xor UO_1244 (O_1244,N_9972,N_9926);
nor UO_1245 (O_1245,N_9964,N_9951);
or UO_1246 (O_1246,N_9921,N_9922);
xor UO_1247 (O_1247,N_9973,N_9907);
nor UO_1248 (O_1248,N_9928,N_9959);
nor UO_1249 (O_1249,N_9933,N_9901);
nor UO_1250 (O_1250,N_9908,N_9966);
or UO_1251 (O_1251,N_9914,N_9964);
or UO_1252 (O_1252,N_9942,N_9971);
xor UO_1253 (O_1253,N_9900,N_9929);
nor UO_1254 (O_1254,N_9939,N_9940);
and UO_1255 (O_1255,N_9929,N_9936);
or UO_1256 (O_1256,N_9972,N_9980);
nand UO_1257 (O_1257,N_9952,N_9985);
and UO_1258 (O_1258,N_9977,N_9907);
xor UO_1259 (O_1259,N_9939,N_9970);
nand UO_1260 (O_1260,N_9978,N_9973);
xnor UO_1261 (O_1261,N_9952,N_9948);
and UO_1262 (O_1262,N_9974,N_9940);
nor UO_1263 (O_1263,N_9914,N_9962);
nor UO_1264 (O_1264,N_9934,N_9996);
nand UO_1265 (O_1265,N_9953,N_9994);
or UO_1266 (O_1266,N_9909,N_9914);
and UO_1267 (O_1267,N_9925,N_9923);
and UO_1268 (O_1268,N_9932,N_9967);
or UO_1269 (O_1269,N_9942,N_9923);
or UO_1270 (O_1270,N_9978,N_9949);
nand UO_1271 (O_1271,N_9953,N_9945);
nor UO_1272 (O_1272,N_9963,N_9945);
xnor UO_1273 (O_1273,N_9951,N_9961);
xnor UO_1274 (O_1274,N_9987,N_9964);
or UO_1275 (O_1275,N_9973,N_9900);
nand UO_1276 (O_1276,N_9903,N_9982);
or UO_1277 (O_1277,N_9940,N_9976);
and UO_1278 (O_1278,N_9928,N_9924);
and UO_1279 (O_1279,N_9921,N_9978);
nand UO_1280 (O_1280,N_9932,N_9959);
nand UO_1281 (O_1281,N_9915,N_9964);
and UO_1282 (O_1282,N_9955,N_9969);
nor UO_1283 (O_1283,N_9962,N_9959);
nor UO_1284 (O_1284,N_9990,N_9909);
xor UO_1285 (O_1285,N_9981,N_9984);
and UO_1286 (O_1286,N_9950,N_9932);
xor UO_1287 (O_1287,N_9946,N_9964);
xnor UO_1288 (O_1288,N_9971,N_9956);
nor UO_1289 (O_1289,N_9958,N_9946);
xnor UO_1290 (O_1290,N_9980,N_9982);
and UO_1291 (O_1291,N_9967,N_9987);
xor UO_1292 (O_1292,N_9906,N_9938);
nand UO_1293 (O_1293,N_9930,N_9914);
or UO_1294 (O_1294,N_9903,N_9930);
and UO_1295 (O_1295,N_9947,N_9920);
or UO_1296 (O_1296,N_9953,N_9990);
nand UO_1297 (O_1297,N_9906,N_9953);
and UO_1298 (O_1298,N_9987,N_9920);
xor UO_1299 (O_1299,N_9972,N_9916);
or UO_1300 (O_1300,N_9983,N_9993);
xor UO_1301 (O_1301,N_9928,N_9966);
or UO_1302 (O_1302,N_9931,N_9953);
and UO_1303 (O_1303,N_9968,N_9909);
xor UO_1304 (O_1304,N_9939,N_9922);
nand UO_1305 (O_1305,N_9946,N_9969);
or UO_1306 (O_1306,N_9957,N_9956);
nor UO_1307 (O_1307,N_9910,N_9930);
and UO_1308 (O_1308,N_9999,N_9940);
xnor UO_1309 (O_1309,N_9946,N_9992);
nand UO_1310 (O_1310,N_9929,N_9983);
and UO_1311 (O_1311,N_9927,N_9978);
and UO_1312 (O_1312,N_9940,N_9985);
and UO_1313 (O_1313,N_9938,N_9956);
or UO_1314 (O_1314,N_9957,N_9927);
and UO_1315 (O_1315,N_9900,N_9976);
or UO_1316 (O_1316,N_9955,N_9966);
and UO_1317 (O_1317,N_9937,N_9919);
xor UO_1318 (O_1318,N_9922,N_9931);
xor UO_1319 (O_1319,N_9954,N_9953);
xor UO_1320 (O_1320,N_9967,N_9956);
nor UO_1321 (O_1321,N_9937,N_9986);
nand UO_1322 (O_1322,N_9922,N_9979);
and UO_1323 (O_1323,N_9953,N_9960);
xor UO_1324 (O_1324,N_9996,N_9942);
nand UO_1325 (O_1325,N_9985,N_9922);
or UO_1326 (O_1326,N_9929,N_9911);
or UO_1327 (O_1327,N_9914,N_9949);
nor UO_1328 (O_1328,N_9993,N_9933);
and UO_1329 (O_1329,N_9980,N_9923);
or UO_1330 (O_1330,N_9931,N_9908);
xor UO_1331 (O_1331,N_9916,N_9959);
nand UO_1332 (O_1332,N_9998,N_9905);
nand UO_1333 (O_1333,N_9956,N_9917);
and UO_1334 (O_1334,N_9902,N_9972);
nor UO_1335 (O_1335,N_9987,N_9906);
and UO_1336 (O_1336,N_9918,N_9952);
xor UO_1337 (O_1337,N_9903,N_9973);
nor UO_1338 (O_1338,N_9915,N_9973);
nor UO_1339 (O_1339,N_9980,N_9902);
nor UO_1340 (O_1340,N_9959,N_9917);
nor UO_1341 (O_1341,N_9942,N_9941);
nand UO_1342 (O_1342,N_9944,N_9936);
or UO_1343 (O_1343,N_9916,N_9948);
nor UO_1344 (O_1344,N_9908,N_9935);
nor UO_1345 (O_1345,N_9907,N_9909);
nand UO_1346 (O_1346,N_9941,N_9995);
xnor UO_1347 (O_1347,N_9940,N_9965);
and UO_1348 (O_1348,N_9951,N_9943);
or UO_1349 (O_1349,N_9980,N_9930);
or UO_1350 (O_1350,N_9963,N_9916);
or UO_1351 (O_1351,N_9928,N_9932);
xnor UO_1352 (O_1352,N_9911,N_9917);
xor UO_1353 (O_1353,N_9973,N_9945);
or UO_1354 (O_1354,N_9948,N_9960);
and UO_1355 (O_1355,N_9938,N_9919);
xor UO_1356 (O_1356,N_9937,N_9943);
xnor UO_1357 (O_1357,N_9928,N_9971);
xnor UO_1358 (O_1358,N_9903,N_9904);
and UO_1359 (O_1359,N_9944,N_9929);
nor UO_1360 (O_1360,N_9964,N_9976);
and UO_1361 (O_1361,N_9970,N_9949);
xor UO_1362 (O_1362,N_9906,N_9926);
xnor UO_1363 (O_1363,N_9975,N_9938);
nand UO_1364 (O_1364,N_9978,N_9957);
or UO_1365 (O_1365,N_9965,N_9900);
or UO_1366 (O_1366,N_9991,N_9968);
nor UO_1367 (O_1367,N_9915,N_9990);
nor UO_1368 (O_1368,N_9991,N_9922);
xnor UO_1369 (O_1369,N_9981,N_9934);
nor UO_1370 (O_1370,N_9927,N_9921);
and UO_1371 (O_1371,N_9994,N_9940);
nor UO_1372 (O_1372,N_9901,N_9984);
and UO_1373 (O_1373,N_9947,N_9915);
and UO_1374 (O_1374,N_9992,N_9928);
xnor UO_1375 (O_1375,N_9960,N_9939);
xor UO_1376 (O_1376,N_9927,N_9964);
or UO_1377 (O_1377,N_9968,N_9919);
nor UO_1378 (O_1378,N_9942,N_9965);
or UO_1379 (O_1379,N_9990,N_9923);
nor UO_1380 (O_1380,N_9952,N_9944);
nand UO_1381 (O_1381,N_9995,N_9933);
or UO_1382 (O_1382,N_9945,N_9903);
or UO_1383 (O_1383,N_9986,N_9935);
xnor UO_1384 (O_1384,N_9959,N_9930);
or UO_1385 (O_1385,N_9907,N_9957);
nand UO_1386 (O_1386,N_9997,N_9915);
nor UO_1387 (O_1387,N_9992,N_9975);
nor UO_1388 (O_1388,N_9907,N_9935);
nand UO_1389 (O_1389,N_9972,N_9984);
xnor UO_1390 (O_1390,N_9933,N_9958);
nand UO_1391 (O_1391,N_9904,N_9901);
or UO_1392 (O_1392,N_9976,N_9994);
nand UO_1393 (O_1393,N_9980,N_9995);
and UO_1394 (O_1394,N_9994,N_9944);
and UO_1395 (O_1395,N_9972,N_9978);
nor UO_1396 (O_1396,N_9973,N_9949);
xnor UO_1397 (O_1397,N_9966,N_9935);
and UO_1398 (O_1398,N_9966,N_9903);
nand UO_1399 (O_1399,N_9900,N_9917);
nand UO_1400 (O_1400,N_9985,N_9909);
or UO_1401 (O_1401,N_9970,N_9909);
nor UO_1402 (O_1402,N_9987,N_9924);
and UO_1403 (O_1403,N_9938,N_9986);
nand UO_1404 (O_1404,N_9907,N_9967);
nor UO_1405 (O_1405,N_9958,N_9997);
nor UO_1406 (O_1406,N_9925,N_9951);
nor UO_1407 (O_1407,N_9945,N_9941);
nor UO_1408 (O_1408,N_9951,N_9958);
nand UO_1409 (O_1409,N_9910,N_9957);
or UO_1410 (O_1410,N_9982,N_9966);
nor UO_1411 (O_1411,N_9912,N_9941);
nand UO_1412 (O_1412,N_9974,N_9928);
xor UO_1413 (O_1413,N_9933,N_9949);
xor UO_1414 (O_1414,N_9920,N_9982);
and UO_1415 (O_1415,N_9909,N_9993);
nor UO_1416 (O_1416,N_9987,N_9954);
nand UO_1417 (O_1417,N_9959,N_9984);
nand UO_1418 (O_1418,N_9904,N_9913);
xor UO_1419 (O_1419,N_9969,N_9985);
or UO_1420 (O_1420,N_9984,N_9936);
and UO_1421 (O_1421,N_9901,N_9936);
or UO_1422 (O_1422,N_9948,N_9903);
xnor UO_1423 (O_1423,N_9916,N_9942);
nand UO_1424 (O_1424,N_9984,N_9917);
nor UO_1425 (O_1425,N_9934,N_9953);
nor UO_1426 (O_1426,N_9961,N_9910);
nand UO_1427 (O_1427,N_9990,N_9920);
xnor UO_1428 (O_1428,N_9954,N_9912);
nor UO_1429 (O_1429,N_9934,N_9926);
nand UO_1430 (O_1430,N_9967,N_9959);
or UO_1431 (O_1431,N_9904,N_9965);
nand UO_1432 (O_1432,N_9993,N_9972);
nand UO_1433 (O_1433,N_9987,N_9993);
and UO_1434 (O_1434,N_9931,N_9986);
nor UO_1435 (O_1435,N_9918,N_9946);
xor UO_1436 (O_1436,N_9993,N_9973);
and UO_1437 (O_1437,N_9945,N_9900);
nor UO_1438 (O_1438,N_9976,N_9965);
xor UO_1439 (O_1439,N_9988,N_9908);
xor UO_1440 (O_1440,N_9961,N_9903);
or UO_1441 (O_1441,N_9907,N_9921);
xnor UO_1442 (O_1442,N_9957,N_9930);
nand UO_1443 (O_1443,N_9907,N_9969);
nor UO_1444 (O_1444,N_9986,N_9904);
nor UO_1445 (O_1445,N_9966,N_9918);
nor UO_1446 (O_1446,N_9978,N_9915);
or UO_1447 (O_1447,N_9966,N_9905);
or UO_1448 (O_1448,N_9914,N_9945);
and UO_1449 (O_1449,N_9981,N_9939);
nor UO_1450 (O_1450,N_9945,N_9920);
or UO_1451 (O_1451,N_9950,N_9925);
and UO_1452 (O_1452,N_9966,N_9919);
and UO_1453 (O_1453,N_9957,N_9900);
and UO_1454 (O_1454,N_9998,N_9912);
xor UO_1455 (O_1455,N_9952,N_9999);
or UO_1456 (O_1456,N_9937,N_9939);
nor UO_1457 (O_1457,N_9923,N_9960);
xor UO_1458 (O_1458,N_9959,N_9968);
nand UO_1459 (O_1459,N_9971,N_9994);
xnor UO_1460 (O_1460,N_9957,N_9936);
and UO_1461 (O_1461,N_9926,N_9979);
nand UO_1462 (O_1462,N_9916,N_9969);
nand UO_1463 (O_1463,N_9918,N_9929);
nor UO_1464 (O_1464,N_9903,N_9917);
xor UO_1465 (O_1465,N_9962,N_9925);
nor UO_1466 (O_1466,N_9940,N_9949);
nand UO_1467 (O_1467,N_9916,N_9993);
xnor UO_1468 (O_1468,N_9969,N_9903);
nand UO_1469 (O_1469,N_9976,N_9975);
nand UO_1470 (O_1470,N_9969,N_9956);
nand UO_1471 (O_1471,N_9905,N_9940);
and UO_1472 (O_1472,N_9978,N_9969);
nand UO_1473 (O_1473,N_9997,N_9930);
or UO_1474 (O_1474,N_9987,N_9941);
nor UO_1475 (O_1475,N_9918,N_9913);
and UO_1476 (O_1476,N_9922,N_9996);
or UO_1477 (O_1477,N_9900,N_9932);
or UO_1478 (O_1478,N_9929,N_9935);
and UO_1479 (O_1479,N_9945,N_9966);
or UO_1480 (O_1480,N_9959,N_9985);
xnor UO_1481 (O_1481,N_9934,N_9912);
nand UO_1482 (O_1482,N_9954,N_9993);
or UO_1483 (O_1483,N_9952,N_9938);
or UO_1484 (O_1484,N_9997,N_9933);
nand UO_1485 (O_1485,N_9968,N_9978);
xnor UO_1486 (O_1486,N_9915,N_9935);
and UO_1487 (O_1487,N_9955,N_9946);
and UO_1488 (O_1488,N_9945,N_9952);
xnor UO_1489 (O_1489,N_9927,N_9902);
and UO_1490 (O_1490,N_9937,N_9925);
or UO_1491 (O_1491,N_9938,N_9916);
xor UO_1492 (O_1492,N_9993,N_9947);
nand UO_1493 (O_1493,N_9910,N_9975);
xnor UO_1494 (O_1494,N_9964,N_9928);
nor UO_1495 (O_1495,N_9981,N_9983);
and UO_1496 (O_1496,N_9996,N_9936);
and UO_1497 (O_1497,N_9994,N_9942);
nand UO_1498 (O_1498,N_9902,N_9983);
nand UO_1499 (O_1499,N_9985,N_9964);
endmodule