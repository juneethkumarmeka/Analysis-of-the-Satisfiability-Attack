module basic_500_3000_500_30_levels_1xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_432,In_450);
xnor U1 (N_1,In_71,In_438);
or U2 (N_2,In_240,In_238);
nand U3 (N_3,In_108,In_17);
nand U4 (N_4,In_217,In_123);
nor U5 (N_5,In_357,In_124);
nor U6 (N_6,In_88,In_247);
and U7 (N_7,In_193,In_322);
or U8 (N_8,In_480,In_11);
nand U9 (N_9,In_142,In_202);
nor U10 (N_10,In_246,In_407);
and U11 (N_11,In_220,In_268);
nand U12 (N_12,In_93,In_199);
xnor U13 (N_13,In_448,In_59);
or U14 (N_14,In_434,In_209);
or U15 (N_15,In_308,In_212);
nand U16 (N_16,In_368,In_398);
nor U17 (N_17,In_230,In_82);
and U18 (N_18,In_478,In_295);
and U19 (N_19,In_376,In_215);
and U20 (N_20,In_239,In_43);
nor U21 (N_21,In_281,In_97);
xor U22 (N_22,In_63,In_185);
and U23 (N_23,In_152,In_305);
nand U24 (N_24,In_80,In_416);
and U25 (N_25,In_360,In_331);
and U26 (N_26,In_203,In_481);
or U27 (N_27,In_380,In_207);
and U28 (N_28,In_126,In_61);
nor U29 (N_29,In_29,In_19);
nand U30 (N_30,In_6,In_26);
or U31 (N_31,In_428,In_286);
nand U32 (N_32,In_187,In_447);
or U33 (N_33,In_266,In_275);
or U34 (N_34,In_355,In_329);
and U35 (N_35,In_2,In_184);
nor U36 (N_36,In_235,In_326);
and U37 (N_37,In_39,In_323);
nand U38 (N_38,In_221,In_405);
nor U39 (N_39,In_421,In_433);
nand U40 (N_40,In_435,In_468);
and U41 (N_41,In_89,In_206);
nand U42 (N_42,In_412,In_77);
and U43 (N_43,In_149,In_38);
nand U44 (N_44,In_437,In_12);
or U45 (N_45,In_301,In_191);
or U46 (N_46,In_482,In_312);
and U47 (N_47,In_351,In_13);
nand U48 (N_48,In_464,In_289);
or U49 (N_49,In_34,In_99);
nor U50 (N_50,In_440,In_200);
or U51 (N_51,In_245,In_455);
nor U52 (N_52,In_271,In_466);
and U53 (N_53,In_287,In_411);
and U54 (N_54,In_392,In_177);
or U55 (N_55,In_188,In_75);
or U56 (N_56,In_48,In_53);
nand U57 (N_57,In_95,In_430);
nor U58 (N_58,In_313,In_137);
and U59 (N_59,In_138,In_297);
nor U60 (N_60,In_121,In_84);
and U61 (N_61,In_255,In_315);
nor U62 (N_62,In_366,In_128);
xor U63 (N_63,In_181,In_79);
nand U64 (N_64,In_379,In_141);
nor U65 (N_65,In_408,In_106);
nand U66 (N_66,In_476,In_417);
nand U67 (N_67,In_498,In_348);
nor U68 (N_68,In_208,In_98);
nor U69 (N_69,In_36,In_40);
and U70 (N_70,In_165,In_429);
or U71 (N_71,In_248,In_33);
and U72 (N_72,In_324,In_342);
nand U73 (N_73,In_216,In_131);
nand U74 (N_74,In_422,In_51);
and U75 (N_75,In_499,In_50);
nor U76 (N_76,In_330,In_495);
or U77 (N_77,In_47,In_413);
nor U78 (N_78,In_284,In_58);
and U79 (N_79,In_104,In_136);
or U80 (N_80,In_171,In_332);
and U81 (N_81,In_192,In_439);
and U82 (N_82,In_160,In_65);
and U83 (N_83,In_122,In_484);
nor U84 (N_84,In_118,In_86);
and U85 (N_85,In_78,In_69);
and U86 (N_86,In_443,In_353);
nor U87 (N_87,In_496,In_190);
nor U88 (N_88,In_120,In_402);
nand U89 (N_89,In_117,In_234);
or U90 (N_90,In_306,In_356);
and U91 (N_91,In_163,In_249);
nor U92 (N_92,In_114,In_479);
and U93 (N_93,In_335,In_22);
and U94 (N_94,In_135,In_172);
nand U95 (N_95,In_487,In_244);
or U96 (N_96,In_57,In_401);
nor U97 (N_97,In_218,In_290);
or U98 (N_98,In_399,In_283);
or U99 (N_99,In_213,In_180);
xnor U100 (N_100,In_389,In_317);
nand U101 (N_101,In_375,In_258);
and U102 (N_102,In_186,In_169);
nor U103 (N_103,In_253,In_85);
or U104 (N_104,In_219,In_293);
nor U105 (N_105,In_103,N_38);
nor U106 (N_106,N_54,N_16);
or U107 (N_107,N_30,N_45);
and U108 (N_108,In_129,N_21);
or U109 (N_109,In_223,In_201);
or U110 (N_110,In_102,In_362);
nand U111 (N_111,In_475,In_497);
nor U112 (N_112,N_2,In_204);
nor U113 (N_113,In_489,In_56);
or U114 (N_114,In_377,In_394);
and U115 (N_115,In_345,In_96);
and U116 (N_116,In_307,N_97);
nand U117 (N_117,In_211,N_41);
nand U118 (N_118,In_66,In_373);
or U119 (N_119,N_42,In_274);
nand U120 (N_120,In_445,In_383);
or U121 (N_121,In_146,In_463);
and U122 (N_122,In_473,In_278);
nand U123 (N_123,N_20,In_277);
nor U124 (N_124,In_35,In_397);
and U125 (N_125,In_304,In_251);
nor U126 (N_126,N_12,N_60);
and U127 (N_127,In_371,In_349);
nor U128 (N_128,In_64,In_272);
or U129 (N_129,N_85,In_343);
or U130 (N_130,In_175,N_24);
or U131 (N_131,In_189,In_45);
nor U132 (N_132,In_400,In_147);
nand U133 (N_133,N_49,N_33);
nand U134 (N_134,In_228,In_302);
nor U135 (N_135,In_153,In_196);
nand U136 (N_136,In_456,In_431);
nand U137 (N_137,In_467,In_242);
nand U138 (N_138,In_83,N_84);
nor U139 (N_139,In_325,In_471);
xnor U140 (N_140,In_16,In_382);
and U141 (N_141,In_352,In_25);
nand U142 (N_142,In_309,N_28);
and U143 (N_143,In_337,In_132);
nor U144 (N_144,In_420,In_350);
xor U145 (N_145,In_173,In_474);
nand U146 (N_146,In_404,N_26);
or U147 (N_147,N_29,N_37);
or U148 (N_148,In_250,In_395);
and U149 (N_149,N_25,In_494);
and U150 (N_150,In_110,In_260);
and U151 (N_151,In_321,In_465);
or U152 (N_152,N_76,In_130);
nand U153 (N_153,N_17,In_340);
nor U154 (N_154,N_82,In_460);
and U155 (N_155,In_363,In_391);
nand U156 (N_156,N_55,In_488);
nor U157 (N_157,In_280,In_195);
or U158 (N_158,In_205,In_101);
nand U159 (N_159,In_170,In_354);
nand U160 (N_160,N_32,N_67);
and U161 (N_161,In_446,In_361);
nand U162 (N_162,In_358,In_457);
nor U163 (N_163,N_78,N_75);
or U164 (N_164,In_424,In_470);
nand U165 (N_165,In_210,In_113);
nand U166 (N_166,N_83,In_336);
and U167 (N_167,In_90,In_94);
nor U168 (N_168,N_19,N_43);
or U169 (N_169,N_69,In_270);
or U170 (N_170,In_257,In_359);
nand U171 (N_171,In_396,N_93);
nor U172 (N_172,In_176,N_66);
nor U173 (N_173,N_81,In_491);
nand U174 (N_174,In_303,N_91);
nand U175 (N_175,N_88,In_107);
nor U176 (N_176,N_3,In_267);
nand U177 (N_177,In_333,In_462);
and U178 (N_178,N_0,In_459);
nand U179 (N_179,In_311,N_86);
nor U180 (N_180,In_384,In_310);
or U181 (N_181,In_154,In_32);
or U182 (N_182,In_21,In_365);
and U183 (N_183,In_37,In_139);
nor U184 (N_184,N_52,In_105);
xnor U185 (N_185,In_162,N_11);
and U186 (N_186,N_8,In_227);
nor U187 (N_187,In_320,In_406);
or U188 (N_188,In_20,In_452);
nor U189 (N_189,N_6,N_80);
nor U190 (N_190,In_436,In_369);
and U191 (N_191,In_116,In_338);
nand U192 (N_192,In_92,In_299);
or U193 (N_193,In_18,In_224);
nand U194 (N_194,In_276,In_150);
nand U195 (N_195,N_98,N_58);
and U196 (N_196,In_0,In_291);
and U197 (N_197,In_418,In_388);
or U198 (N_198,In_461,In_72);
or U199 (N_199,In_490,N_89);
nand U200 (N_200,In_485,In_341);
and U201 (N_201,In_74,N_138);
nor U202 (N_202,N_174,In_55);
and U203 (N_203,In_441,In_231);
or U204 (N_204,N_118,In_100);
or U205 (N_205,N_191,N_105);
and U206 (N_206,In_23,N_199);
and U207 (N_207,N_154,In_263);
and U208 (N_208,N_157,In_9);
nand U209 (N_209,N_101,N_170);
nor U210 (N_210,In_419,N_46);
and U211 (N_211,In_168,N_1);
nor U212 (N_212,In_5,N_65);
nor U213 (N_213,N_150,In_285);
nor U214 (N_214,N_5,In_469);
nand U215 (N_215,In_31,N_186);
nand U216 (N_216,In_27,N_74);
or U217 (N_217,In_314,N_48);
and U218 (N_218,In_269,In_296);
nand U219 (N_219,In_237,N_167);
nor U220 (N_220,In_133,N_178);
nand U221 (N_221,In_194,N_165);
nor U222 (N_222,In_279,In_44);
nor U223 (N_223,N_134,N_166);
or U224 (N_224,In_115,N_179);
and U225 (N_225,N_168,N_47);
and U226 (N_226,N_147,N_155);
nand U227 (N_227,N_145,In_339);
and U228 (N_228,N_185,N_63);
or U229 (N_229,N_127,In_449);
or U230 (N_230,In_226,N_161);
nand U231 (N_231,In_387,N_187);
and U232 (N_232,In_492,In_367);
or U233 (N_233,In_159,In_241);
nor U234 (N_234,In_182,In_214);
nor U235 (N_235,In_1,N_177);
and U236 (N_236,N_64,N_44);
nor U237 (N_237,N_96,N_120);
nor U238 (N_238,N_102,In_261);
nor U239 (N_239,In_233,In_483);
and U240 (N_240,In_347,In_109);
nor U241 (N_241,N_111,N_194);
and U242 (N_242,In_453,N_59);
or U243 (N_243,In_151,N_13);
and U244 (N_244,N_142,N_193);
nand U245 (N_245,N_110,N_151);
xnor U246 (N_246,N_50,N_136);
nor U247 (N_247,N_183,In_386);
nor U248 (N_248,In_444,N_56);
and U249 (N_249,N_131,N_173);
and U250 (N_250,N_95,In_328);
xor U251 (N_251,In_197,In_143);
or U252 (N_252,In_486,N_112);
nor U253 (N_253,In_236,In_334);
nand U254 (N_254,In_166,N_72);
nor U255 (N_255,N_40,In_222);
nor U256 (N_256,In_183,N_163);
nand U257 (N_257,N_125,N_22);
nor U258 (N_258,In_427,In_54);
nor U259 (N_259,N_18,N_143);
or U260 (N_260,In_125,In_344);
and U261 (N_261,N_34,In_157);
nand U262 (N_262,N_73,N_190);
nand U263 (N_263,In_316,N_158);
nor U264 (N_264,In_174,In_119);
or U265 (N_265,In_167,In_393);
nand U266 (N_266,In_477,N_23);
and U267 (N_267,In_127,N_172);
and U268 (N_268,In_46,N_176);
nor U269 (N_269,In_425,N_100);
nand U270 (N_270,In_145,N_113);
or U271 (N_271,N_135,In_164);
nand U272 (N_272,In_52,In_91);
or U273 (N_273,In_8,N_87);
or U274 (N_274,N_126,N_68);
nor U275 (N_275,N_140,N_7);
nor U276 (N_276,In_294,N_106);
nor U277 (N_277,In_265,N_71);
and U278 (N_278,In_179,N_192);
nor U279 (N_279,N_162,In_252);
or U280 (N_280,N_109,In_229);
nor U281 (N_281,N_160,N_115);
and U282 (N_282,N_156,In_178);
nand U283 (N_283,In_24,N_119);
and U284 (N_284,In_81,N_27);
nor U285 (N_285,In_87,N_195);
nand U286 (N_286,N_122,In_300);
or U287 (N_287,N_139,N_129);
nand U288 (N_288,In_254,In_60);
nand U289 (N_289,N_117,In_298);
nand U290 (N_290,In_390,N_10);
nand U291 (N_291,N_99,In_140);
and U292 (N_292,In_414,N_92);
and U293 (N_293,N_36,In_15);
and U294 (N_294,In_225,In_472);
nor U295 (N_295,In_410,In_70);
nor U296 (N_296,N_164,In_385);
or U297 (N_297,N_79,N_104);
and U298 (N_298,In_426,In_161);
nor U299 (N_299,N_133,In_259);
nor U300 (N_300,N_159,N_277);
and U301 (N_301,N_205,N_144);
nand U302 (N_302,N_223,N_279);
nor U303 (N_303,In_372,In_292);
and U304 (N_304,N_225,In_73);
and U305 (N_305,N_130,N_128);
nor U306 (N_306,In_7,N_149);
nor U307 (N_307,In_148,N_242);
nor U308 (N_308,In_144,N_61);
and U309 (N_309,N_270,N_53);
or U310 (N_310,N_189,In_273);
nor U311 (N_311,N_227,N_240);
nand U312 (N_312,N_247,N_70);
nand U313 (N_313,N_35,N_235);
or U314 (N_314,N_267,In_112);
nor U315 (N_315,N_188,N_15);
nand U316 (N_316,N_271,N_77);
and U317 (N_317,N_236,N_299);
nor U318 (N_318,N_218,N_39);
nor U319 (N_319,N_215,N_261);
or U320 (N_320,N_248,In_3);
or U321 (N_321,N_273,In_156);
nor U322 (N_322,N_243,N_239);
xor U323 (N_323,In_370,N_224);
nor U324 (N_324,N_294,In_327);
and U325 (N_325,In_198,N_296);
and U326 (N_326,N_124,In_14);
and U327 (N_327,N_275,N_266);
nand U328 (N_328,In_111,In_67);
and U329 (N_329,N_229,N_292);
nand U330 (N_330,N_290,N_175);
nand U331 (N_331,N_249,N_57);
nand U332 (N_332,N_291,N_278);
nor U333 (N_333,N_121,N_226);
nand U334 (N_334,N_214,N_254);
nand U335 (N_335,N_232,N_123);
xor U336 (N_336,N_288,N_116);
nor U337 (N_337,N_209,In_28);
nor U338 (N_338,In_454,N_201);
or U339 (N_339,N_216,N_200);
and U340 (N_340,In_264,N_257);
and U341 (N_341,In_134,N_219);
nand U342 (N_342,In_68,In_364);
and U343 (N_343,In_76,N_231);
or U344 (N_344,N_103,In_423);
nor U345 (N_345,N_244,N_146);
nand U346 (N_346,N_210,N_169);
or U347 (N_347,N_241,N_253);
nand U348 (N_348,In_458,In_493);
nand U349 (N_349,N_259,In_30);
nand U350 (N_350,N_31,In_318);
and U351 (N_351,In_158,N_237);
and U352 (N_352,N_107,N_283);
or U353 (N_353,N_228,In_378);
and U354 (N_354,N_286,N_260);
and U355 (N_355,In_403,N_282);
nor U356 (N_356,N_181,In_319);
nand U357 (N_357,N_297,N_251);
or U358 (N_358,In_256,In_442);
nor U359 (N_359,N_246,N_184);
and U360 (N_360,N_250,N_207);
nor U361 (N_361,N_287,In_243);
and U362 (N_362,N_137,N_298);
and U363 (N_363,N_153,N_256);
nor U364 (N_364,In_262,N_62);
nand U365 (N_365,N_203,N_171);
nor U366 (N_366,In_155,N_198);
nor U367 (N_367,N_255,N_202);
and U368 (N_368,N_148,N_9);
nor U369 (N_369,In_282,N_141);
and U370 (N_370,N_182,N_114);
or U371 (N_371,N_284,N_152);
and U372 (N_372,N_230,N_211);
and U373 (N_373,In_232,N_274);
or U374 (N_374,N_217,N_213);
and U375 (N_375,N_289,N_238);
and U376 (N_376,N_220,In_415);
nand U377 (N_377,N_245,In_4);
nor U378 (N_378,In_41,N_180);
nor U379 (N_379,N_233,N_51);
nor U380 (N_380,N_14,N_262);
or U381 (N_381,In_62,N_221);
and U382 (N_382,In_10,N_258);
or U383 (N_383,N_4,In_374);
and U384 (N_384,In_49,In_288);
nand U385 (N_385,N_295,N_212);
nor U386 (N_386,N_252,In_451);
and U387 (N_387,In_409,N_272);
and U388 (N_388,In_42,N_234);
nor U389 (N_389,N_208,N_90);
and U390 (N_390,N_197,N_280);
nor U391 (N_391,In_346,N_132);
nor U392 (N_392,N_263,N_276);
nand U393 (N_393,N_264,N_281);
nand U394 (N_394,N_285,In_381);
or U395 (N_395,N_265,N_222);
nand U396 (N_396,N_268,N_293);
or U397 (N_397,N_206,N_269);
nand U398 (N_398,N_196,N_204);
nor U399 (N_399,N_108,N_94);
and U400 (N_400,N_361,N_355);
nor U401 (N_401,N_330,N_368);
nor U402 (N_402,N_393,N_315);
nand U403 (N_403,N_327,N_376);
nor U404 (N_404,N_391,N_387);
nand U405 (N_405,N_335,N_338);
and U406 (N_406,N_350,N_307);
and U407 (N_407,N_331,N_333);
and U408 (N_408,N_319,N_348);
or U409 (N_409,N_347,N_369);
and U410 (N_410,N_300,N_358);
and U411 (N_411,N_377,N_353);
and U412 (N_412,N_362,N_375);
or U413 (N_413,N_308,N_356);
nand U414 (N_414,N_344,N_334);
and U415 (N_415,N_381,N_352);
nor U416 (N_416,N_366,N_396);
or U417 (N_417,N_397,N_303);
and U418 (N_418,N_367,N_378);
nand U419 (N_419,N_314,N_371);
or U420 (N_420,N_317,N_394);
nand U421 (N_421,N_386,N_341);
and U422 (N_422,N_329,N_398);
nand U423 (N_423,N_340,N_304);
nand U424 (N_424,N_302,N_354);
nor U425 (N_425,N_324,N_389);
or U426 (N_426,N_399,N_383);
and U427 (N_427,N_360,N_310);
nand U428 (N_428,N_346,N_385);
nand U429 (N_429,N_342,N_332);
nor U430 (N_430,N_313,N_326);
or U431 (N_431,N_343,N_328);
and U432 (N_432,N_312,N_301);
nor U433 (N_433,N_384,N_306);
nor U434 (N_434,N_316,N_309);
nor U435 (N_435,N_390,N_351);
nor U436 (N_436,N_323,N_382);
nor U437 (N_437,N_374,N_380);
nor U438 (N_438,N_322,N_373);
nand U439 (N_439,N_349,N_392);
and U440 (N_440,N_395,N_318);
nand U441 (N_441,N_325,N_372);
and U442 (N_442,N_388,N_336);
nor U443 (N_443,N_311,N_345);
or U444 (N_444,N_305,N_357);
and U445 (N_445,N_379,N_365);
or U446 (N_446,N_363,N_364);
and U447 (N_447,N_321,N_337);
nor U448 (N_448,N_320,N_339);
and U449 (N_449,N_370,N_359);
and U450 (N_450,N_316,N_391);
or U451 (N_451,N_362,N_326);
nand U452 (N_452,N_324,N_399);
nand U453 (N_453,N_378,N_362);
or U454 (N_454,N_361,N_390);
nor U455 (N_455,N_382,N_367);
or U456 (N_456,N_348,N_379);
nand U457 (N_457,N_378,N_361);
and U458 (N_458,N_388,N_384);
and U459 (N_459,N_343,N_305);
nor U460 (N_460,N_369,N_386);
or U461 (N_461,N_360,N_300);
or U462 (N_462,N_318,N_330);
and U463 (N_463,N_302,N_367);
and U464 (N_464,N_318,N_300);
nor U465 (N_465,N_343,N_349);
nor U466 (N_466,N_337,N_306);
and U467 (N_467,N_377,N_378);
or U468 (N_468,N_355,N_376);
and U469 (N_469,N_314,N_341);
nor U470 (N_470,N_353,N_320);
nand U471 (N_471,N_378,N_324);
or U472 (N_472,N_316,N_353);
nor U473 (N_473,N_317,N_323);
and U474 (N_474,N_305,N_370);
or U475 (N_475,N_396,N_304);
or U476 (N_476,N_385,N_307);
nor U477 (N_477,N_357,N_314);
and U478 (N_478,N_333,N_332);
nand U479 (N_479,N_342,N_370);
nand U480 (N_480,N_395,N_368);
nor U481 (N_481,N_303,N_313);
nor U482 (N_482,N_323,N_378);
nor U483 (N_483,N_334,N_397);
nand U484 (N_484,N_312,N_359);
and U485 (N_485,N_389,N_325);
and U486 (N_486,N_396,N_307);
nor U487 (N_487,N_363,N_396);
and U488 (N_488,N_371,N_331);
nand U489 (N_489,N_326,N_311);
or U490 (N_490,N_350,N_377);
nand U491 (N_491,N_390,N_396);
and U492 (N_492,N_386,N_397);
nor U493 (N_493,N_377,N_368);
and U494 (N_494,N_314,N_377);
nand U495 (N_495,N_333,N_352);
or U496 (N_496,N_345,N_347);
and U497 (N_497,N_356,N_313);
and U498 (N_498,N_311,N_391);
and U499 (N_499,N_374,N_341);
or U500 (N_500,N_406,N_400);
and U501 (N_501,N_472,N_448);
nand U502 (N_502,N_441,N_496);
or U503 (N_503,N_451,N_428);
nor U504 (N_504,N_409,N_421);
or U505 (N_505,N_447,N_414);
and U506 (N_506,N_465,N_498);
and U507 (N_507,N_488,N_453);
nor U508 (N_508,N_499,N_477);
and U509 (N_509,N_471,N_426);
nor U510 (N_510,N_446,N_422);
xnor U511 (N_511,N_455,N_450);
or U512 (N_512,N_443,N_424);
or U513 (N_513,N_405,N_423);
nand U514 (N_514,N_412,N_467);
nand U515 (N_515,N_431,N_401);
nor U516 (N_516,N_460,N_403);
nand U517 (N_517,N_438,N_466);
and U518 (N_518,N_482,N_486);
nor U519 (N_519,N_495,N_417);
or U520 (N_520,N_429,N_410);
or U521 (N_521,N_485,N_458);
nand U522 (N_522,N_407,N_419);
or U523 (N_523,N_478,N_449);
or U524 (N_524,N_456,N_420);
or U525 (N_525,N_445,N_469);
nor U526 (N_526,N_484,N_416);
nand U527 (N_527,N_491,N_497);
nor U528 (N_528,N_468,N_463);
and U529 (N_529,N_411,N_436);
and U530 (N_530,N_452,N_494);
nor U531 (N_531,N_457,N_427);
or U532 (N_532,N_425,N_439);
nor U533 (N_533,N_408,N_435);
nand U534 (N_534,N_462,N_402);
and U535 (N_535,N_430,N_413);
and U536 (N_536,N_444,N_461);
nand U537 (N_537,N_483,N_470);
nor U538 (N_538,N_415,N_490);
and U539 (N_539,N_454,N_459);
or U540 (N_540,N_474,N_404);
or U541 (N_541,N_475,N_481);
and U542 (N_542,N_476,N_464);
nor U543 (N_543,N_492,N_434);
nor U544 (N_544,N_489,N_440);
or U545 (N_545,N_418,N_442);
or U546 (N_546,N_493,N_480);
nand U547 (N_547,N_433,N_473);
xor U548 (N_548,N_479,N_432);
nand U549 (N_549,N_487,N_437);
nor U550 (N_550,N_402,N_482);
nand U551 (N_551,N_439,N_434);
or U552 (N_552,N_471,N_450);
nand U553 (N_553,N_437,N_464);
nor U554 (N_554,N_463,N_427);
nand U555 (N_555,N_457,N_473);
and U556 (N_556,N_467,N_425);
nand U557 (N_557,N_439,N_453);
nor U558 (N_558,N_464,N_450);
nor U559 (N_559,N_404,N_416);
and U560 (N_560,N_411,N_422);
or U561 (N_561,N_464,N_405);
nor U562 (N_562,N_409,N_494);
and U563 (N_563,N_454,N_443);
nor U564 (N_564,N_462,N_424);
nand U565 (N_565,N_423,N_486);
nand U566 (N_566,N_476,N_466);
nand U567 (N_567,N_434,N_404);
nor U568 (N_568,N_402,N_409);
nor U569 (N_569,N_447,N_496);
nor U570 (N_570,N_447,N_469);
or U571 (N_571,N_487,N_471);
nand U572 (N_572,N_427,N_493);
and U573 (N_573,N_465,N_455);
or U574 (N_574,N_490,N_496);
nand U575 (N_575,N_402,N_436);
nand U576 (N_576,N_415,N_462);
nor U577 (N_577,N_477,N_426);
nand U578 (N_578,N_478,N_410);
nor U579 (N_579,N_462,N_420);
nor U580 (N_580,N_444,N_488);
nor U581 (N_581,N_483,N_449);
nand U582 (N_582,N_485,N_421);
nor U583 (N_583,N_457,N_496);
nand U584 (N_584,N_448,N_499);
nor U585 (N_585,N_452,N_418);
nand U586 (N_586,N_453,N_467);
nor U587 (N_587,N_439,N_407);
nand U588 (N_588,N_410,N_443);
or U589 (N_589,N_415,N_444);
or U590 (N_590,N_408,N_404);
nand U591 (N_591,N_495,N_407);
nor U592 (N_592,N_431,N_429);
and U593 (N_593,N_437,N_468);
or U594 (N_594,N_409,N_445);
nand U595 (N_595,N_472,N_427);
nand U596 (N_596,N_446,N_402);
nor U597 (N_597,N_417,N_446);
and U598 (N_598,N_425,N_499);
and U599 (N_599,N_455,N_424);
nand U600 (N_600,N_540,N_536);
and U601 (N_601,N_514,N_597);
or U602 (N_602,N_551,N_595);
nor U603 (N_603,N_549,N_557);
or U604 (N_604,N_518,N_571);
nand U605 (N_605,N_504,N_568);
or U606 (N_606,N_545,N_510);
nor U607 (N_607,N_554,N_593);
nor U608 (N_608,N_592,N_563);
nor U609 (N_609,N_525,N_587);
and U610 (N_610,N_576,N_535);
nor U611 (N_611,N_555,N_558);
or U612 (N_612,N_511,N_581);
or U613 (N_613,N_594,N_574);
nand U614 (N_614,N_596,N_584);
or U615 (N_615,N_552,N_515);
and U616 (N_616,N_529,N_516);
and U617 (N_617,N_556,N_570);
nor U618 (N_618,N_585,N_531);
nand U619 (N_619,N_569,N_520);
nor U620 (N_620,N_527,N_533);
and U621 (N_621,N_524,N_562);
nand U622 (N_622,N_505,N_537);
and U623 (N_623,N_579,N_548);
and U624 (N_624,N_591,N_538);
nor U625 (N_625,N_580,N_598);
and U626 (N_626,N_502,N_541);
nand U627 (N_627,N_507,N_561);
nand U628 (N_628,N_526,N_542);
or U629 (N_629,N_532,N_590);
nand U630 (N_630,N_589,N_577);
nor U631 (N_631,N_513,N_572);
nor U632 (N_632,N_501,N_582);
nor U633 (N_633,N_539,N_547);
and U634 (N_634,N_544,N_528);
nor U635 (N_635,N_586,N_530);
and U636 (N_636,N_522,N_566);
and U637 (N_637,N_560,N_575);
or U638 (N_638,N_573,N_534);
nor U639 (N_639,N_599,N_519);
and U640 (N_640,N_578,N_559);
nor U641 (N_641,N_523,N_508);
nand U642 (N_642,N_588,N_512);
or U643 (N_643,N_565,N_506);
or U644 (N_644,N_543,N_564);
nand U645 (N_645,N_509,N_517);
or U646 (N_646,N_550,N_583);
xor U647 (N_647,N_553,N_521);
or U648 (N_648,N_500,N_503);
nand U649 (N_649,N_546,N_567);
nand U650 (N_650,N_511,N_597);
or U651 (N_651,N_547,N_588);
nor U652 (N_652,N_516,N_505);
nand U653 (N_653,N_578,N_500);
and U654 (N_654,N_595,N_564);
or U655 (N_655,N_549,N_596);
and U656 (N_656,N_529,N_530);
nand U657 (N_657,N_554,N_503);
or U658 (N_658,N_553,N_534);
or U659 (N_659,N_562,N_534);
and U660 (N_660,N_508,N_522);
or U661 (N_661,N_515,N_593);
nand U662 (N_662,N_520,N_539);
nor U663 (N_663,N_535,N_549);
or U664 (N_664,N_525,N_590);
nand U665 (N_665,N_525,N_556);
and U666 (N_666,N_510,N_596);
nand U667 (N_667,N_537,N_554);
and U668 (N_668,N_504,N_546);
and U669 (N_669,N_502,N_544);
nand U670 (N_670,N_504,N_525);
or U671 (N_671,N_502,N_560);
nor U672 (N_672,N_580,N_503);
nor U673 (N_673,N_542,N_524);
nor U674 (N_674,N_576,N_575);
nand U675 (N_675,N_507,N_503);
nand U676 (N_676,N_573,N_530);
nor U677 (N_677,N_569,N_598);
and U678 (N_678,N_533,N_520);
or U679 (N_679,N_536,N_556);
nand U680 (N_680,N_521,N_554);
and U681 (N_681,N_571,N_591);
nand U682 (N_682,N_552,N_554);
nand U683 (N_683,N_538,N_544);
or U684 (N_684,N_554,N_519);
and U685 (N_685,N_588,N_529);
nor U686 (N_686,N_513,N_574);
or U687 (N_687,N_599,N_556);
or U688 (N_688,N_534,N_518);
and U689 (N_689,N_549,N_593);
and U690 (N_690,N_598,N_582);
or U691 (N_691,N_588,N_556);
and U692 (N_692,N_596,N_520);
and U693 (N_693,N_509,N_503);
nand U694 (N_694,N_585,N_560);
nor U695 (N_695,N_532,N_513);
nor U696 (N_696,N_522,N_528);
nand U697 (N_697,N_564,N_560);
or U698 (N_698,N_539,N_556);
nor U699 (N_699,N_581,N_558);
nor U700 (N_700,N_698,N_695);
nand U701 (N_701,N_622,N_629);
nor U702 (N_702,N_608,N_601);
and U703 (N_703,N_681,N_636);
nand U704 (N_704,N_615,N_686);
or U705 (N_705,N_672,N_600);
nand U706 (N_706,N_628,N_697);
nand U707 (N_707,N_641,N_635);
nor U708 (N_708,N_637,N_633);
nand U709 (N_709,N_671,N_604);
and U710 (N_710,N_658,N_677);
or U711 (N_711,N_620,N_607);
or U712 (N_712,N_662,N_609);
and U713 (N_713,N_696,N_653);
nor U714 (N_714,N_640,N_626);
or U715 (N_715,N_652,N_647);
nand U716 (N_716,N_643,N_668);
nor U717 (N_717,N_699,N_621);
nor U718 (N_718,N_669,N_654);
nand U719 (N_719,N_648,N_638);
nand U720 (N_720,N_678,N_670);
and U721 (N_721,N_676,N_694);
nor U722 (N_722,N_673,N_674);
nand U723 (N_723,N_691,N_664);
or U724 (N_724,N_625,N_657);
nand U725 (N_725,N_689,N_612);
or U726 (N_726,N_630,N_644);
or U727 (N_727,N_682,N_690);
nor U728 (N_728,N_679,N_659);
nor U729 (N_729,N_649,N_650);
or U730 (N_730,N_605,N_606);
nand U731 (N_731,N_675,N_634);
and U732 (N_732,N_680,N_666);
nand U733 (N_733,N_663,N_684);
nand U734 (N_734,N_687,N_645);
and U735 (N_735,N_646,N_692);
nor U736 (N_736,N_614,N_603);
or U737 (N_737,N_632,N_618);
nand U738 (N_738,N_610,N_665);
and U739 (N_739,N_619,N_623);
nand U740 (N_740,N_656,N_602);
nand U741 (N_741,N_613,N_683);
nand U742 (N_742,N_616,N_661);
and U743 (N_743,N_642,N_660);
or U744 (N_744,N_611,N_624);
nor U745 (N_745,N_627,N_651);
or U746 (N_746,N_685,N_693);
nor U747 (N_747,N_631,N_688);
nor U748 (N_748,N_617,N_667);
nor U749 (N_749,N_639,N_655);
nor U750 (N_750,N_667,N_673);
nand U751 (N_751,N_642,N_606);
nor U752 (N_752,N_616,N_614);
and U753 (N_753,N_618,N_639);
or U754 (N_754,N_650,N_602);
and U755 (N_755,N_671,N_697);
or U756 (N_756,N_626,N_610);
or U757 (N_757,N_696,N_669);
or U758 (N_758,N_644,N_632);
or U759 (N_759,N_643,N_621);
and U760 (N_760,N_620,N_657);
and U761 (N_761,N_666,N_630);
nor U762 (N_762,N_677,N_670);
and U763 (N_763,N_616,N_683);
nor U764 (N_764,N_603,N_671);
and U765 (N_765,N_622,N_611);
nand U766 (N_766,N_663,N_616);
and U767 (N_767,N_679,N_610);
nor U768 (N_768,N_609,N_696);
nor U769 (N_769,N_698,N_670);
nor U770 (N_770,N_695,N_622);
and U771 (N_771,N_663,N_674);
or U772 (N_772,N_674,N_688);
nand U773 (N_773,N_693,N_650);
nor U774 (N_774,N_687,N_617);
nor U775 (N_775,N_626,N_670);
nand U776 (N_776,N_675,N_690);
nand U777 (N_777,N_625,N_600);
nor U778 (N_778,N_675,N_605);
nor U779 (N_779,N_612,N_678);
nor U780 (N_780,N_630,N_614);
or U781 (N_781,N_622,N_677);
nand U782 (N_782,N_615,N_662);
or U783 (N_783,N_658,N_687);
nand U784 (N_784,N_685,N_663);
nor U785 (N_785,N_618,N_645);
and U786 (N_786,N_642,N_616);
and U787 (N_787,N_649,N_679);
and U788 (N_788,N_623,N_690);
nand U789 (N_789,N_665,N_633);
or U790 (N_790,N_606,N_658);
nand U791 (N_791,N_655,N_647);
nor U792 (N_792,N_607,N_637);
nor U793 (N_793,N_694,N_645);
nand U794 (N_794,N_603,N_660);
or U795 (N_795,N_657,N_632);
nand U796 (N_796,N_669,N_680);
nand U797 (N_797,N_676,N_670);
and U798 (N_798,N_603,N_632);
nor U799 (N_799,N_699,N_616);
or U800 (N_800,N_790,N_777);
or U801 (N_801,N_764,N_755);
and U802 (N_802,N_713,N_719);
or U803 (N_803,N_789,N_754);
nand U804 (N_804,N_772,N_778);
or U805 (N_805,N_722,N_741);
nor U806 (N_806,N_727,N_781);
or U807 (N_807,N_715,N_773);
and U808 (N_808,N_792,N_729);
nor U809 (N_809,N_737,N_703);
xor U810 (N_810,N_770,N_783);
or U811 (N_811,N_736,N_760);
nor U812 (N_812,N_780,N_785);
xnor U813 (N_813,N_743,N_776);
and U814 (N_814,N_716,N_718);
and U815 (N_815,N_730,N_701);
nand U816 (N_816,N_732,N_717);
xor U817 (N_817,N_751,N_775);
nand U818 (N_818,N_712,N_750);
or U819 (N_819,N_706,N_767);
nand U820 (N_820,N_723,N_787);
nor U821 (N_821,N_740,N_725);
nor U822 (N_822,N_700,N_711);
nand U823 (N_823,N_797,N_748);
and U824 (N_824,N_794,N_774);
nor U825 (N_825,N_708,N_707);
nand U826 (N_826,N_762,N_739);
nor U827 (N_827,N_724,N_752);
and U828 (N_828,N_731,N_746);
xnor U829 (N_829,N_786,N_768);
and U830 (N_830,N_734,N_702);
and U831 (N_831,N_766,N_798);
or U832 (N_832,N_742,N_784);
and U833 (N_833,N_721,N_759);
nand U834 (N_834,N_795,N_735);
nand U835 (N_835,N_757,N_744);
nor U836 (N_836,N_793,N_709);
and U837 (N_837,N_761,N_782);
nor U838 (N_838,N_765,N_745);
nor U839 (N_839,N_799,N_728);
or U840 (N_840,N_753,N_720);
and U841 (N_841,N_733,N_710);
nand U842 (N_842,N_749,N_771);
nor U843 (N_843,N_714,N_788);
and U844 (N_844,N_763,N_758);
nand U845 (N_845,N_791,N_705);
or U846 (N_846,N_726,N_779);
nand U847 (N_847,N_769,N_747);
and U848 (N_848,N_756,N_738);
or U849 (N_849,N_796,N_704);
and U850 (N_850,N_733,N_744);
nor U851 (N_851,N_727,N_719);
or U852 (N_852,N_775,N_765);
nand U853 (N_853,N_785,N_776);
or U854 (N_854,N_715,N_744);
and U855 (N_855,N_745,N_721);
and U856 (N_856,N_782,N_796);
nor U857 (N_857,N_718,N_710);
nand U858 (N_858,N_740,N_743);
and U859 (N_859,N_748,N_708);
nand U860 (N_860,N_779,N_768);
nor U861 (N_861,N_781,N_742);
and U862 (N_862,N_738,N_713);
nand U863 (N_863,N_735,N_770);
nand U864 (N_864,N_731,N_797);
or U865 (N_865,N_733,N_711);
and U866 (N_866,N_737,N_776);
nand U867 (N_867,N_708,N_772);
or U868 (N_868,N_754,N_793);
nor U869 (N_869,N_710,N_706);
nor U870 (N_870,N_799,N_727);
and U871 (N_871,N_741,N_751);
or U872 (N_872,N_747,N_754);
nor U873 (N_873,N_767,N_715);
nor U874 (N_874,N_787,N_789);
nand U875 (N_875,N_761,N_733);
and U876 (N_876,N_712,N_708);
nand U877 (N_877,N_704,N_728);
or U878 (N_878,N_731,N_790);
nor U879 (N_879,N_759,N_766);
nor U880 (N_880,N_770,N_778);
nor U881 (N_881,N_714,N_768);
nand U882 (N_882,N_717,N_759);
and U883 (N_883,N_733,N_734);
nand U884 (N_884,N_725,N_788);
nand U885 (N_885,N_758,N_734);
or U886 (N_886,N_777,N_747);
nand U887 (N_887,N_778,N_752);
nand U888 (N_888,N_753,N_755);
nor U889 (N_889,N_711,N_756);
nand U890 (N_890,N_726,N_757);
nor U891 (N_891,N_792,N_730);
and U892 (N_892,N_785,N_747);
nand U893 (N_893,N_706,N_782);
nor U894 (N_894,N_738,N_751);
nor U895 (N_895,N_769,N_792);
and U896 (N_896,N_782,N_718);
nor U897 (N_897,N_779,N_788);
nand U898 (N_898,N_796,N_724);
nand U899 (N_899,N_774,N_701);
nand U900 (N_900,N_856,N_828);
and U901 (N_901,N_846,N_858);
nor U902 (N_902,N_859,N_876);
and U903 (N_903,N_874,N_888);
nand U904 (N_904,N_841,N_838);
nor U905 (N_905,N_818,N_843);
and U906 (N_906,N_823,N_892);
nor U907 (N_907,N_883,N_875);
or U908 (N_908,N_839,N_881);
nand U909 (N_909,N_821,N_861);
and U910 (N_910,N_851,N_826);
or U911 (N_911,N_804,N_837);
or U912 (N_912,N_868,N_865);
nand U913 (N_913,N_840,N_852);
nor U914 (N_914,N_848,N_869);
nor U915 (N_915,N_806,N_815);
nor U916 (N_916,N_860,N_817);
and U917 (N_917,N_877,N_895);
and U918 (N_918,N_849,N_800);
and U919 (N_919,N_827,N_824);
nor U920 (N_920,N_814,N_889);
and U921 (N_921,N_842,N_884);
nand U922 (N_922,N_811,N_822);
nand U923 (N_923,N_887,N_819);
or U924 (N_924,N_820,N_897);
and U925 (N_925,N_857,N_885);
nor U926 (N_926,N_805,N_802);
nor U927 (N_927,N_855,N_829);
nand U928 (N_928,N_813,N_890);
or U929 (N_929,N_844,N_886);
nor U930 (N_930,N_834,N_873);
nor U931 (N_931,N_833,N_879);
nand U932 (N_932,N_810,N_866);
nor U933 (N_933,N_836,N_899);
or U934 (N_934,N_825,N_893);
nor U935 (N_935,N_832,N_847);
nor U936 (N_936,N_809,N_898);
nand U937 (N_937,N_850,N_867);
nand U938 (N_938,N_853,N_830);
nor U939 (N_939,N_891,N_862);
nand U940 (N_940,N_882,N_812);
nor U941 (N_941,N_894,N_801);
nand U942 (N_942,N_807,N_872);
nor U943 (N_943,N_863,N_845);
nor U944 (N_944,N_870,N_896);
and U945 (N_945,N_871,N_835);
nand U946 (N_946,N_854,N_803);
or U947 (N_947,N_816,N_808);
nand U948 (N_948,N_880,N_864);
and U949 (N_949,N_878,N_831);
and U950 (N_950,N_878,N_857);
or U951 (N_951,N_802,N_843);
nand U952 (N_952,N_883,N_887);
nand U953 (N_953,N_809,N_883);
or U954 (N_954,N_859,N_817);
or U955 (N_955,N_858,N_803);
nand U956 (N_956,N_839,N_899);
and U957 (N_957,N_816,N_898);
nand U958 (N_958,N_833,N_851);
and U959 (N_959,N_810,N_804);
and U960 (N_960,N_834,N_821);
and U961 (N_961,N_896,N_877);
nor U962 (N_962,N_850,N_859);
or U963 (N_963,N_878,N_856);
and U964 (N_964,N_884,N_878);
nand U965 (N_965,N_886,N_834);
nand U966 (N_966,N_804,N_889);
nor U967 (N_967,N_840,N_838);
nor U968 (N_968,N_845,N_864);
and U969 (N_969,N_896,N_892);
nand U970 (N_970,N_809,N_887);
or U971 (N_971,N_898,N_868);
or U972 (N_972,N_818,N_839);
nand U973 (N_973,N_869,N_873);
and U974 (N_974,N_838,N_817);
nor U975 (N_975,N_871,N_889);
nor U976 (N_976,N_885,N_809);
and U977 (N_977,N_869,N_860);
or U978 (N_978,N_813,N_852);
nor U979 (N_979,N_899,N_833);
or U980 (N_980,N_800,N_801);
nand U981 (N_981,N_820,N_845);
and U982 (N_982,N_896,N_829);
nand U983 (N_983,N_806,N_830);
or U984 (N_984,N_805,N_896);
nand U985 (N_985,N_821,N_894);
nor U986 (N_986,N_821,N_853);
nor U987 (N_987,N_818,N_869);
nor U988 (N_988,N_880,N_829);
or U989 (N_989,N_867,N_868);
nor U990 (N_990,N_881,N_850);
or U991 (N_991,N_886,N_837);
or U992 (N_992,N_844,N_898);
and U993 (N_993,N_825,N_802);
or U994 (N_994,N_820,N_819);
or U995 (N_995,N_836,N_845);
or U996 (N_996,N_893,N_865);
nor U997 (N_997,N_831,N_803);
xnor U998 (N_998,N_815,N_800);
or U999 (N_999,N_807,N_878);
and U1000 (N_1000,N_905,N_953);
or U1001 (N_1001,N_957,N_987);
and U1002 (N_1002,N_969,N_981);
or U1003 (N_1003,N_960,N_919);
or U1004 (N_1004,N_955,N_918);
or U1005 (N_1005,N_984,N_932);
nor U1006 (N_1006,N_937,N_997);
and U1007 (N_1007,N_959,N_989);
and U1008 (N_1008,N_965,N_961);
nand U1009 (N_1009,N_970,N_943);
nand U1010 (N_1010,N_972,N_927);
nand U1011 (N_1011,N_942,N_928);
nand U1012 (N_1012,N_964,N_940);
and U1013 (N_1013,N_944,N_949);
nand U1014 (N_1014,N_921,N_910);
nor U1015 (N_1015,N_936,N_903);
and U1016 (N_1016,N_966,N_945);
nor U1017 (N_1017,N_985,N_926);
nand U1018 (N_1018,N_999,N_929);
nand U1019 (N_1019,N_952,N_994);
nor U1020 (N_1020,N_973,N_907);
nand U1021 (N_1021,N_902,N_930);
and U1022 (N_1022,N_998,N_982);
nor U1023 (N_1023,N_980,N_967);
and U1024 (N_1024,N_978,N_925);
or U1025 (N_1025,N_924,N_993);
and U1026 (N_1026,N_920,N_904);
nor U1027 (N_1027,N_947,N_968);
or U1028 (N_1028,N_977,N_914);
and U1029 (N_1029,N_963,N_974);
and U1030 (N_1030,N_938,N_933);
nand U1031 (N_1031,N_922,N_906);
nor U1032 (N_1032,N_916,N_946);
or U1033 (N_1033,N_975,N_931);
or U1034 (N_1034,N_992,N_941);
nor U1035 (N_1035,N_956,N_909);
nor U1036 (N_1036,N_901,N_990);
or U1037 (N_1037,N_958,N_995);
or U1038 (N_1038,N_913,N_951);
nand U1039 (N_1039,N_986,N_976);
and U1040 (N_1040,N_911,N_900);
or U1041 (N_1041,N_939,N_948);
nand U1042 (N_1042,N_954,N_988);
or U1043 (N_1043,N_983,N_917);
nand U1044 (N_1044,N_908,N_934);
nand U1045 (N_1045,N_915,N_962);
and U1046 (N_1046,N_923,N_935);
and U1047 (N_1047,N_971,N_979);
or U1048 (N_1048,N_912,N_991);
and U1049 (N_1049,N_996,N_950);
nor U1050 (N_1050,N_935,N_971);
nor U1051 (N_1051,N_925,N_984);
or U1052 (N_1052,N_945,N_941);
nor U1053 (N_1053,N_984,N_940);
or U1054 (N_1054,N_991,N_960);
nand U1055 (N_1055,N_997,N_984);
nand U1056 (N_1056,N_992,N_924);
nand U1057 (N_1057,N_946,N_972);
nand U1058 (N_1058,N_913,N_972);
nor U1059 (N_1059,N_971,N_945);
nor U1060 (N_1060,N_939,N_966);
nand U1061 (N_1061,N_942,N_919);
and U1062 (N_1062,N_952,N_941);
nand U1063 (N_1063,N_936,N_918);
nand U1064 (N_1064,N_969,N_947);
and U1065 (N_1065,N_949,N_960);
or U1066 (N_1066,N_963,N_908);
or U1067 (N_1067,N_980,N_948);
or U1068 (N_1068,N_982,N_977);
nand U1069 (N_1069,N_958,N_967);
nand U1070 (N_1070,N_944,N_932);
nor U1071 (N_1071,N_970,N_930);
nand U1072 (N_1072,N_976,N_971);
or U1073 (N_1073,N_979,N_943);
nand U1074 (N_1074,N_943,N_983);
or U1075 (N_1075,N_916,N_938);
nand U1076 (N_1076,N_974,N_917);
or U1077 (N_1077,N_920,N_934);
or U1078 (N_1078,N_958,N_982);
nor U1079 (N_1079,N_991,N_938);
and U1080 (N_1080,N_959,N_992);
nor U1081 (N_1081,N_945,N_964);
nor U1082 (N_1082,N_909,N_901);
or U1083 (N_1083,N_932,N_926);
xnor U1084 (N_1084,N_921,N_941);
nand U1085 (N_1085,N_947,N_907);
or U1086 (N_1086,N_956,N_974);
nand U1087 (N_1087,N_984,N_930);
nor U1088 (N_1088,N_980,N_936);
or U1089 (N_1089,N_947,N_900);
nand U1090 (N_1090,N_954,N_994);
and U1091 (N_1091,N_900,N_982);
or U1092 (N_1092,N_971,N_922);
or U1093 (N_1093,N_978,N_977);
or U1094 (N_1094,N_993,N_994);
and U1095 (N_1095,N_944,N_965);
nor U1096 (N_1096,N_996,N_924);
nor U1097 (N_1097,N_904,N_946);
and U1098 (N_1098,N_991,N_956);
nor U1099 (N_1099,N_901,N_957);
and U1100 (N_1100,N_1053,N_1023);
or U1101 (N_1101,N_1008,N_1098);
and U1102 (N_1102,N_1041,N_1052);
and U1103 (N_1103,N_1014,N_1019);
or U1104 (N_1104,N_1021,N_1058);
nor U1105 (N_1105,N_1044,N_1092);
and U1106 (N_1106,N_1097,N_1026);
or U1107 (N_1107,N_1007,N_1096);
nor U1108 (N_1108,N_1011,N_1065);
nand U1109 (N_1109,N_1069,N_1063);
nor U1110 (N_1110,N_1033,N_1031);
nor U1111 (N_1111,N_1006,N_1038);
or U1112 (N_1112,N_1076,N_1068);
nand U1113 (N_1113,N_1036,N_1070);
nor U1114 (N_1114,N_1040,N_1054);
nand U1115 (N_1115,N_1000,N_1018);
nor U1116 (N_1116,N_1039,N_1066);
or U1117 (N_1117,N_1029,N_1043);
and U1118 (N_1118,N_1013,N_1024);
nor U1119 (N_1119,N_1091,N_1046);
or U1120 (N_1120,N_1035,N_1034);
or U1121 (N_1121,N_1042,N_1009);
nor U1122 (N_1122,N_1073,N_1020);
nand U1123 (N_1123,N_1055,N_1060);
nor U1124 (N_1124,N_1010,N_1090);
or U1125 (N_1125,N_1088,N_1004);
or U1126 (N_1126,N_1080,N_1089);
or U1127 (N_1127,N_1049,N_1027);
nor U1128 (N_1128,N_1059,N_1071);
or U1129 (N_1129,N_1017,N_1099);
or U1130 (N_1130,N_1048,N_1061);
nand U1131 (N_1131,N_1082,N_1062);
nor U1132 (N_1132,N_1074,N_1056);
and U1133 (N_1133,N_1083,N_1085);
nand U1134 (N_1134,N_1057,N_1022);
nand U1135 (N_1135,N_1002,N_1064);
and U1136 (N_1136,N_1086,N_1015);
nand U1137 (N_1137,N_1025,N_1030);
nor U1138 (N_1138,N_1078,N_1016);
or U1139 (N_1139,N_1047,N_1093);
or U1140 (N_1140,N_1079,N_1072);
or U1141 (N_1141,N_1028,N_1001);
or U1142 (N_1142,N_1095,N_1012);
nor U1143 (N_1143,N_1081,N_1094);
and U1144 (N_1144,N_1003,N_1084);
nand U1145 (N_1145,N_1087,N_1075);
nand U1146 (N_1146,N_1050,N_1077);
nand U1147 (N_1147,N_1037,N_1045);
nand U1148 (N_1148,N_1067,N_1032);
or U1149 (N_1149,N_1051,N_1005);
or U1150 (N_1150,N_1065,N_1042);
nand U1151 (N_1151,N_1004,N_1038);
and U1152 (N_1152,N_1078,N_1001);
nor U1153 (N_1153,N_1023,N_1033);
and U1154 (N_1154,N_1066,N_1084);
or U1155 (N_1155,N_1045,N_1033);
or U1156 (N_1156,N_1077,N_1084);
or U1157 (N_1157,N_1017,N_1096);
or U1158 (N_1158,N_1014,N_1064);
nand U1159 (N_1159,N_1069,N_1027);
or U1160 (N_1160,N_1064,N_1041);
nor U1161 (N_1161,N_1043,N_1085);
or U1162 (N_1162,N_1093,N_1036);
nor U1163 (N_1163,N_1076,N_1030);
and U1164 (N_1164,N_1086,N_1008);
or U1165 (N_1165,N_1075,N_1038);
nand U1166 (N_1166,N_1016,N_1087);
xor U1167 (N_1167,N_1068,N_1013);
and U1168 (N_1168,N_1022,N_1092);
nor U1169 (N_1169,N_1077,N_1052);
and U1170 (N_1170,N_1004,N_1082);
nand U1171 (N_1171,N_1063,N_1027);
or U1172 (N_1172,N_1024,N_1072);
nor U1173 (N_1173,N_1086,N_1081);
and U1174 (N_1174,N_1072,N_1019);
nand U1175 (N_1175,N_1051,N_1088);
or U1176 (N_1176,N_1065,N_1020);
xor U1177 (N_1177,N_1056,N_1013);
nand U1178 (N_1178,N_1052,N_1071);
or U1179 (N_1179,N_1081,N_1061);
nand U1180 (N_1180,N_1061,N_1020);
nand U1181 (N_1181,N_1086,N_1014);
and U1182 (N_1182,N_1002,N_1039);
nand U1183 (N_1183,N_1088,N_1017);
nor U1184 (N_1184,N_1038,N_1077);
nand U1185 (N_1185,N_1079,N_1077);
or U1186 (N_1186,N_1096,N_1043);
nand U1187 (N_1187,N_1080,N_1091);
or U1188 (N_1188,N_1061,N_1011);
and U1189 (N_1189,N_1047,N_1064);
and U1190 (N_1190,N_1069,N_1061);
nand U1191 (N_1191,N_1059,N_1055);
and U1192 (N_1192,N_1015,N_1008);
and U1193 (N_1193,N_1022,N_1003);
nor U1194 (N_1194,N_1062,N_1034);
and U1195 (N_1195,N_1069,N_1072);
or U1196 (N_1196,N_1020,N_1003);
or U1197 (N_1197,N_1022,N_1049);
and U1198 (N_1198,N_1008,N_1030);
nor U1199 (N_1199,N_1082,N_1076);
or U1200 (N_1200,N_1162,N_1179);
and U1201 (N_1201,N_1139,N_1163);
or U1202 (N_1202,N_1114,N_1193);
or U1203 (N_1203,N_1156,N_1192);
and U1204 (N_1204,N_1127,N_1113);
nand U1205 (N_1205,N_1183,N_1104);
nor U1206 (N_1206,N_1166,N_1184);
and U1207 (N_1207,N_1137,N_1194);
nand U1208 (N_1208,N_1141,N_1172);
or U1209 (N_1209,N_1105,N_1198);
and U1210 (N_1210,N_1157,N_1161);
or U1211 (N_1211,N_1129,N_1171);
nand U1212 (N_1212,N_1190,N_1107);
nor U1213 (N_1213,N_1119,N_1153);
or U1214 (N_1214,N_1146,N_1109);
nand U1215 (N_1215,N_1145,N_1134);
and U1216 (N_1216,N_1135,N_1103);
nand U1217 (N_1217,N_1154,N_1191);
nor U1218 (N_1218,N_1177,N_1188);
nand U1219 (N_1219,N_1116,N_1195);
and U1220 (N_1220,N_1197,N_1131);
and U1221 (N_1221,N_1102,N_1110);
nor U1222 (N_1222,N_1196,N_1144);
or U1223 (N_1223,N_1128,N_1180);
nand U1224 (N_1224,N_1187,N_1118);
or U1225 (N_1225,N_1165,N_1174);
and U1226 (N_1226,N_1169,N_1126);
or U1227 (N_1227,N_1159,N_1121);
and U1228 (N_1228,N_1112,N_1108);
nor U1229 (N_1229,N_1160,N_1130);
nand U1230 (N_1230,N_1182,N_1125);
nand U1231 (N_1231,N_1147,N_1133);
nor U1232 (N_1232,N_1155,N_1173);
nand U1233 (N_1233,N_1100,N_1122);
and U1234 (N_1234,N_1117,N_1168);
or U1235 (N_1235,N_1106,N_1167);
nor U1236 (N_1236,N_1149,N_1111);
nor U1237 (N_1237,N_1185,N_1158);
nor U1238 (N_1238,N_1143,N_1138);
and U1239 (N_1239,N_1186,N_1124);
nor U1240 (N_1240,N_1170,N_1136);
nand U1241 (N_1241,N_1164,N_1189);
xnor U1242 (N_1242,N_1101,N_1142);
or U1243 (N_1243,N_1140,N_1150);
nor U1244 (N_1244,N_1123,N_1120);
and U1245 (N_1245,N_1178,N_1148);
or U1246 (N_1246,N_1199,N_1175);
nor U1247 (N_1247,N_1115,N_1151);
or U1248 (N_1248,N_1152,N_1132);
and U1249 (N_1249,N_1176,N_1181);
and U1250 (N_1250,N_1165,N_1157);
or U1251 (N_1251,N_1115,N_1180);
nor U1252 (N_1252,N_1168,N_1105);
nor U1253 (N_1253,N_1129,N_1147);
or U1254 (N_1254,N_1191,N_1146);
nand U1255 (N_1255,N_1112,N_1153);
nand U1256 (N_1256,N_1173,N_1144);
or U1257 (N_1257,N_1110,N_1135);
nor U1258 (N_1258,N_1193,N_1159);
and U1259 (N_1259,N_1100,N_1173);
or U1260 (N_1260,N_1199,N_1165);
or U1261 (N_1261,N_1195,N_1137);
nand U1262 (N_1262,N_1144,N_1146);
nand U1263 (N_1263,N_1139,N_1189);
or U1264 (N_1264,N_1177,N_1183);
nand U1265 (N_1265,N_1194,N_1174);
nand U1266 (N_1266,N_1179,N_1148);
or U1267 (N_1267,N_1179,N_1147);
and U1268 (N_1268,N_1105,N_1199);
nand U1269 (N_1269,N_1155,N_1197);
or U1270 (N_1270,N_1137,N_1180);
nand U1271 (N_1271,N_1129,N_1164);
and U1272 (N_1272,N_1140,N_1131);
nand U1273 (N_1273,N_1110,N_1104);
nand U1274 (N_1274,N_1189,N_1133);
and U1275 (N_1275,N_1183,N_1188);
nand U1276 (N_1276,N_1182,N_1126);
nor U1277 (N_1277,N_1140,N_1129);
or U1278 (N_1278,N_1142,N_1135);
and U1279 (N_1279,N_1117,N_1185);
nand U1280 (N_1280,N_1159,N_1100);
or U1281 (N_1281,N_1148,N_1130);
or U1282 (N_1282,N_1181,N_1133);
nor U1283 (N_1283,N_1114,N_1106);
and U1284 (N_1284,N_1197,N_1106);
nor U1285 (N_1285,N_1186,N_1169);
nand U1286 (N_1286,N_1107,N_1110);
nor U1287 (N_1287,N_1174,N_1135);
and U1288 (N_1288,N_1129,N_1174);
or U1289 (N_1289,N_1150,N_1184);
nor U1290 (N_1290,N_1189,N_1169);
or U1291 (N_1291,N_1128,N_1153);
and U1292 (N_1292,N_1191,N_1139);
nor U1293 (N_1293,N_1101,N_1111);
or U1294 (N_1294,N_1191,N_1107);
nand U1295 (N_1295,N_1168,N_1198);
nor U1296 (N_1296,N_1104,N_1132);
and U1297 (N_1297,N_1175,N_1151);
or U1298 (N_1298,N_1137,N_1159);
nand U1299 (N_1299,N_1171,N_1159);
nand U1300 (N_1300,N_1232,N_1205);
or U1301 (N_1301,N_1202,N_1284);
and U1302 (N_1302,N_1228,N_1208);
nor U1303 (N_1303,N_1215,N_1262);
and U1304 (N_1304,N_1261,N_1244);
and U1305 (N_1305,N_1206,N_1214);
nand U1306 (N_1306,N_1240,N_1235);
and U1307 (N_1307,N_1213,N_1264);
and U1308 (N_1308,N_1278,N_1289);
or U1309 (N_1309,N_1210,N_1286);
nor U1310 (N_1310,N_1282,N_1217);
and U1311 (N_1311,N_1231,N_1230);
nand U1312 (N_1312,N_1241,N_1292);
nand U1313 (N_1313,N_1255,N_1259);
nand U1314 (N_1314,N_1263,N_1276);
nor U1315 (N_1315,N_1257,N_1252);
nor U1316 (N_1316,N_1221,N_1265);
nand U1317 (N_1317,N_1258,N_1236);
nor U1318 (N_1318,N_1219,N_1267);
nand U1319 (N_1319,N_1256,N_1296);
nor U1320 (N_1320,N_1290,N_1297);
nand U1321 (N_1321,N_1253,N_1218);
nand U1322 (N_1322,N_1266,N_1272);
or U1323 (N_1323,N_1222,N_1268);
nand U1324 (N_1324,N_1203,N_1239);
nand U1325 (N_1325,N_1250,N_1287);
and U1326 (N_1326,N_1248,N_1293);
and U1327 (N_1327,N_1288,N_1298);
or U1328 (N_1328,N_1299,N_1280);
nand U1329 (N_1329,N_1247,N_1283);
or U1330 (N_1330,N_1226,N_1201);
or U1331 (N_1331,N_1204,N_1224);
or U1332 (N_1332,N_1220,N_1260);
and U1333 (N_1333,N_1251,N_1216);
nor U1334 (N_1334,N_1243,N_1285);
and U1335 (N_1335,N_1270,N_1245);
and U1336 (N_1336,N_1212,N_1200);
and U1337 (N_1337,N_1225,N_1238);
nand U1338 (N_1338,N_1277,N_1254);
nor U1339 (N_1339,N_1234,N_1207);
or U1340 (N_1340,N_1294,N_1279);
nor U1341 (N_1341,N_1275,N_1242);
nand U1342 (N_1342,N_1291,N_1211);
nand U1343 (N_1343,N_1271,N_1274);
and U1344 (N_1344,N_1227,N_1229);
nand U1345 (N_1345,N_1273,N_1246);
or U1346 (N_1346,N_1281,N_1233);
nor U1347 (N_1347,N_1223,N_1209);
nand U1348 (N_1348,N_1237,N_1295);
or U1349 (N_1349,N_1269,N_1249);
or U1350 (N_1350,N_1257,N_1215);
and U1351 (N_1351,N_1273,N_1272);
and U1352 (N_1352,N_1265,N_1204);
and U1353 (N_1353,N_1265,N_1218);
nand U1354 (N_1354,N_1234,N_1208);
nor U1355 (N_1355,N_1268,N_1233);
and U1356 (N_1356,N_1201,N_1258);
nor U1357 (N_1357,N_1217,N_1298);
or U1358 (N_1358,N_1249,N_1245);
or U1359 (N_1359,N_1258,N_1245);
nand U1360 (N_1360,N_1203,N_1288);
and U1361 (N_1361,N_1262,N_1268);
nand U1362 (N_1362,N_1218,N_1283);
nand U1363 (N_1363,N_1260,N_1206);
and U1364 (N_1364,N_1254,N_1268);
nand U1365 (N_1365,N_1239,N_1263);
nand U1366 (N_1366,N_1212,N_1298);
nand U1367 (N_1367,N_1283,N_1269);
or U1368 (N_1368,N_1221,N_1279);
or U1369 (N_1369,N_1230,N_1257);
and U1370 (N_1370,N_1262,N_1246);
nor U1371 (N_1371,N_1268,N_1240);
nor U1372 (N_1372,N_1272,N_1278);
nor U1373 (N_1373,N_1249,N_1243);
and U1374 (N_1374,N_1211,N_1224);
or U1375 (N_1375,N_1299,N_1292);
or U1376 (N_1376,N_1275,N_1239);
or U1377 (N_1377,N_1232,N_1299);
and U1378 (N_1378,N_1217,N_1281);
and U1379 (N_1379,N_1261,N_1248);
nand U1380 (N_1380,N_1241,N_1243);
and U1381 (N_1381,N_1294,N_1242);
or U1382 (N_1382,N_1223,N_1298);
nand U1383 (N_1383,N_1237,N_1219);
nor U1384 (N_1384,N_1207,N_1201);
nand U1385 (N_1385,N_1266,N_1279);
nor U1386 (N_1386,N_1252,N_1217);
nand U1387 (N_1387,N_1238,N_1271);
nor U1388 (N_1388,N_1219,N_1265);
nand U1389 (N_1389,N_1217,N_1272);
and U1390 (N_1390,N_1293,N_1277);
and U1391 (N_1391,N_1284,N_1252);
nand U1392 (N_1392,N_1229,N_1244);
and U1393 (N_1393,N_1234,N_1267);
and U1394 (N_1394,N_1222,N_1285);
nand U1395 (N_1395,N_1274,N_1210);
nand U1396 (N_1396,N_1253,N_1278);
or U1397 (N_1397,N_1205,N_1284);
nor U1398 (N_1398,N_1211,N_1250);
and U1399 (N_1399,N_1241,N_1267);
or U1400 (N_1400,N_1330,N_1372);
nor U1401 (N_1401,N_1310,N_1307);
and U1402 (N_1402,N_1398,N_1303);
or U1403 (N_1403,N_1313,N_1354);
and U1404 (N_1404,N_1367,N_1332);
xor U1405 (N_1405,N_1317,N_1327);
or U1406 (N_1406,N_1338,N_1381);
or U1407 (N_1407,N_1341,N_1324);
nand U1408 (N_1408,N_1333,N_1320);
nor U1409 (N_1409,N_1318,N_1393);
nand U1410 (N_1410,N_1355,N_1383);
nor U1411 (N_1411,N_1391,N_1350);
or U1412 (N_1412,N_1343,N_1358);
and U1413 (N_1413,N_1308,N_1379);
nand U1414 (N_1414,N_1380,N_1377);
or U1415 (N_1415,N_1346,N_1392);
or U1416 (N_1416,N_1315,N_1305);
and U1417 (N_1417,N_1375,N_1331);
or U1418 (N_1418,N_1335,N_1314);
nand U1419 (N_1419,N_1362,N_1389);
and U1420 (N_1420,N_1394,N_1360);
nor U1421 (N_1421,N_1349,N_1388);
and U1422 (N_1422,N_1347,N_1322);
nand U1423 (N_1423,N_1373,N_1337);
and U1424 (N_1424,N_1374,N_1306);
nor U1425 (N_1425,N_1316,N_1370);
nand U1426 (N_1426,N_1353,N_1364);
nand U1427 (N_1427,N_1323,N_1351);
nand U1428 (N_1428,N_1352,N_1369);
and U1429 (N_1429,N_1386,N_1342);
and U1430 (N_1430,N_1395,N_1396);
or U1431 (N_1431,N_1361,N_1325);
nor U1432 (N_1432,N_1357,N_1384);
nand U1433 (N_1433,N_1376,N_1312);
and U1434 (N_1434,N_1339,N_1397);
or U1435 (N_1435,N_1321,N_1326);
and U1436 (N_1436,N_1300,N_1368);
or U1437 (N_1437,N_1334,N_1359);
nor U1438 (N_1438,N_1301,N_1382);
and U1439 (N_1439,N_1345,N_1399);
nor U1440 (N_1440,N_1365,N_1344);
nand U1441 (N_1441,N_1366,N_1328);
and U1442 (N_1442,N_1311,N_1302);
nor U1443 (N_1443,N_1385,N_1309);
and U1444 (N_1444,N_1371,N_1319);
nand U1445 (N_1445,N_1304,N_1348);
or U1446 (N_1446,N_1378,N_1336);
nor U1447 (N_1447,N_1363,N_1329);
or U1448 (N_1448,N_1390,N_1387);
and U1449 (N_1449,N_1340,N_1356);
nand U1450 (N_1450,N_1317,N_1389);
nor U1451 (N_1451,N_1320,N_1343);
nand U1452 (N_1452,N_1313,N_1369);
and U1453 (N_1453,N_1381,N_1392);
nor U1454 (N_1454,N_1392,N_1343);
xor U1455 (N_1455,N_1358,N_1328);
nand U1456 (N_1456,N_1307,N_1358);
and U1457 (N_1457,N_1327,N_1393);
nor U1458 (N_1458,N_1338,N_1365);
nor U1459 (N_1459,N_1368,N_1316);
nor U1460 (N_1460,N_1307,N_1390);
nor U1461 (N_1461,N_1355,N_1373);
xnor U1462 (N_1462,N_1340,N_1308);
and U1463 (N_1463,N_1329,N_1382);
nand U1464 (N_1464,N_1379,N_1302);
nand U1465 (N_1465,N_1305,N_1365);
nand U1466 (N_1466,N_1363,N_1349);
nand U1467 (N_1467,N_1362,N_1340);
nand U1468 (N_1468,N_1358,N_1398);
nor U1469 (N_1469,N_1300,N_1378);
nand U1470 (N_1470,N_1325,N_1337);
nand U1471 (N_1471,N_1303,N_1366);
and U1472 (N_1472,N_1341,N_1322);
or U1473 (N_1473,N_1369,N_1373);
and U1474 (N_1474,N_1345,N_1370);
nand U1475 (N_1475,N_1324,N_1370);
nor U1476 (N_1476,N_1368,N_1376);
nand U1477 (N_1477,N_1308,N_1319);
and U1478 (N_1478,N_1384,N_1347);
nor U1479 (N_1479,N_1321,N_1301);
nor U1480 (N_1480,N_1325,N_1350);
and U1481 (N_1481,N_1378,N_1366);
nand U1482 (N_1482,N_1318,N_1346);
or U1483 (N_1483,N_1390,N_1333);
nor U1484 (N_1484,N_1336,N_1350);
and U1485 (N_1485,N_1392,N_1342);
and U1486 (N_1486,N_1355,N_1374);
nor U1487 (N_1487,N_1387,N_1354);
nand U1488 (N_1488,N_1348,N_1309);
nor U1489 (N_1489,N_1342,N_1303);
and U1490 (N_1490,N_1376,N_1332);
and U1491 (N_1491,N_1338,N_1316);
nand U1492 (N_1492,N_1369,N_1364);
or U1493 (N_1493,N_1379,N_1397);
nand U1494 (N_1494,N_1321,N_1325);
xnor U1495 (N_1495,N_1346,N_1379);
nor U1496 (N_1496,N_1321,N_1342);
and U1497 (N_1497,N_1372,N_1317);
and U1498 (N_1498,N_1384,N_1313);
nor U1499 (N_1499,N_1350,N_1321);
or U1500 (N_1500,N_1445,N_1453);
or U1501 (N_1501,N_1438,N_1428);
or U1502 (N_1502,N_1471,N_1414);
and U1503 (N_1503,N_1429,N_1402);
and U1504 (N_1504,N_1493,N_1469);
nor U1505 (N_1505,N_1432,N_1486);
nand U1506 (N_1506,N_1431,N_1491);
nor U1507 (N_1507,N_1456,N_1461);
nor U1508 (N_1508,N_1465,N_1479);
or U1509 (N_1509,N_1457,N_1415);
nand U1510 (N_1510,N_1455,N_1446);
or U1511 (N_1511,N_1498,N_1416);
or U1512 (N_1512,N_1443,N_1483);
or U1513 (N_1513,N_1475,N_1449);
or U1514 (N_1514,N_1441,N_1458);
nor U1515 (N_1515,N_1489,N_1401);
or U1516 (N_1516,N_1448,N_1407);
or U1517 (N_1517,N_1464,N_1462);
or U1518 (N_1518,N_1425,N_1434);
and U1519 (N_1519,N_1452,N_1480);
nand U1520 (N_1520,N_1436,N_1419);
and U1521 (N_1521,N_1466,N_1460);
and U1522 (N_1522,N_1422,N_1442);
nor U1523 (N_1523,N_1410,N_1421);
nor U1524 (N_1524,N_1450,N_1485);
nand U1525 (N_1525,N_1435,N_1412);
nand U1526 (N_1526,N_1440,N_1492);
nand U1527 (N_1527,N_1463,N_1437);
or U1528 (N_1528,N_1404,N_1454);
and U1529 (N_1529,N_1496,N_1484);
nand U1530 (N_1530,N_1474,N_1439);
or U1531 (N_1531,N_1424,N_1418);
or U1532 (N_1532,N_1487,N_1403);
nand U1533 (N_1533,N_1490,N_1444);
nand U1534 (N_1534,N_1476,N_1451);
or U1535 (N_1535,N_1481,N_1477);
and U1536 (N_1536,N_1499,N_1400);
or U1537 (N_1537,N_1417,N_1406);
nor U1538 (N_1538,N_1420,N_1405);
nor U1539 (N_1539,N_1447,N_1467);
or U1540 (N_1540,N_1426,N_1433);
and U1541 (N_1541,N_1472,N_1495);
and U1542 (N_1542,N_1459,N_1488);
nor U1543 (N_1543,N_1411,N_1482);
or U1544 (N_1544,N_1473,N_1408);
or U1545 (N_1545,N_1478,N_1423);
nand U1546 (N_1546,N_1430,N_1409);
nor U1547 (N_1547,N_1494,N_1470);
nor U1548 (N_1548,N_1497,N_1468);
nand U1549 (N_1549,N_1427,N_1413);
nor U1550 (N_1550,N_1495,N_1402);
or U1551 (N_1551,N_1475,N_1461);
or U1552 (N_1552,N_1408,N_1416);
nand U1553 (N_1553,N_1478,N_1416);
nand U1554 (N_1554,N_1420,N_1492);
nand U1555 (N_1555,N_1461,N_1458);
and U1556 (N_1556,N_1473,N_1469);
nor U1557 (N_1557,N_1463,N_1400);
nand U1558 (N_1558,N_1405,N_1425);
or U1559 (N_1559,N_1444,N_1445);
nor U1560 (N_1560,N_1414,N_1402);
nand U1561 (N_1561,N_1473,N_1498);
xnor U1562 (N_1562,N_1427,N_1441);
nand U1563 (N_1563,N_1466,N_1417);
and U1564 (N_1564,N_1428,N_1477);
or U1565 (N_1565,N_1498,N_1436);
and U1566 (N_1566,N_1496,N_1478);
nor U1567 (N_1567,N_1445,N_1474);
nand U1568 (N_1568,N_1496,N_1434);
nand U1569 (N_1569,N_1442,N_1463);
nand U1570 (N_1570,N_1418,N_1474);
or U1571 (N_1571,N_1493,N_1435);
nand U1572 (N_1572,N_1458,N_1480);
or U1573 (N_1573,N_1410,N_1411);
nor U1574 (N_1574,N_1442,N_1408);
or U1575 (N_1575,N_1441,N_1415);
or U1576 (N_1576,N_1450,N_1496);
and U1577 (N_1577,N_1468,N_1499);
nor U1578 (N_1578,N_1448,N_1456);
nand U1579 (N_1579,N_1474,N_1423);
or U1580 (N_1580,N_1459,N_1490);
nor U1581 (N_1581,N_1442,N_1424);
nand U1582 (N_1582,N_1423,N_1468);
nand U1583 (N_1583,N_1412,N_1482);
and U1584 (N_1584,N_1499,N_1414);
or U1585 (N_1585,N_1465,N_1470);
nor U1586 (N_1586,N_1493,N_1498);
nor U1587 (N_1587,N_1406,N_1450);
nand U1588 (N_1588,N_1475,N_1404);
or U1589 (N_1589,N_1462,N_1410);
nand U1590 (N_1590,N_1402,N_1451);
nor U1591 (N_1591,N_1435,N_1490);
and U1592 (N_1592,N_1422,N_1428);
nor U1593 (N_1593,N_1457,N_1435);
nand U1594 (N_1594,N_1430,N_1414);
and U1595 (N_1595,N_1468,N_1470);
and U1596 (N_1596,N_1465,N_1467);
and U1597 (N_1597,N_1495,N_1440);
nor U1598 (N_1598,N_1446,N_1467);
nor U1599 (N_1599,N_1409,N_1410);
nand U1600 (N_1600,N_1596,N_1553);
and U1601 (N_1601,N_1544,N_1563);
nand U1602 (N_1602,N_1552,N_1571);
and U1603 (N_1603,N_1501,N_1586);
or U1604 (N_1604,N_1525,N_1582);
nor U1605 (N_1605,N_1531,N_1595);
and U1606 (N_1606,N_1562,N_1580);
or U1607 (N_1607,N_1532,N_1581);
nand U1608 (N_1608,N_1516,N_1518);
nand U1609 (N_1609,N_1576,N_1597);
and U1610 (N_1610,N_1585,N_1570);
nand U1611 (N_1611,N_1590,N_1507);
and U1612 (N_1612,N_1529,N_1589);
and U1613 (N_1613,N_1538,N_1502);
or U1614 (N_1614,N_1547,N_1545);
nand U1615 (N_1615,N_1541,N_1565);
and U1616 (N_1616,N_1530,N_1568);
and U1617 (N_1617,N_1535,N_1519);
or U1618 (N_1618,N_1591,N_1567);
nand U1619 (N_1619,N_1524,N_1555);
and U1620 (N_1620,N_1592,N_1569);
nand U1621 (N_1621,N_1599,N_1546);
nor U1622 (N_1622,N_1526,N_1549);
or U1623 (N_1623,N_1574,N_1523);
and U1624 (N_1624,N_1500,N_1514);
and U1625 (N_1625,N_1583,N_1548);
and U1626 (N_1626,N_1578,N_1537);
nor U1627 (N_1627,N_1543,N_1527);
and U1628 (N_1628,N_1575,N_1551);
and U1629 (N_1629,N_1593,N_1566);
nor U1630 (N_1630,N_1521,N_1533);
and U1631 (N_1631,N_1528,N_1588);
nand U1632 (N_1632,N_1564,N_1540);
nor U1633 (N_1633,N_1513,N_1573);
or U1634 (N_1634,N_1510,N_1506);
and U1635 (N_1635,N_1515,N_1557);
or U1636 (N_1636,N_1554,N_1572);
nand U1637 (N_1637,N_1594,N_1508);
or U1638 (N_1638,N_1504,N_1560);
nor U1639 (N_1639,N_1512,N_1522);
nand U1640 (N_1640,N_1536,N_1505);
or U1641 (N_1641,N_1561,N_1534);
nand U1642 (N_1642,N_1511,N_1556);
and U1643 (N_1643,N_1584,N_1539);
nand U1644 (N_1644,N_1550,N_1517);
or U1645 (N_1645,N_1520,N_1587);
and U1646 (N_1646,N_1558,N_1577);
nor U1647 (N_1647,N_1598,N_1509);
nand U1648 (N_1648,N_1542,N_1559);
and U1649 (N_1649,N_1503,N_1579);
and U1650 (N_1650,N_1501,N_1567);
nand U1651 (N_1651,N_1538,N_1593);
nand U1652 (N_1652,N_1589,N_1558);
nor U1653 (N_1653,N_1527,N_1560);
nand U1654 (N_1654,N_1533,N_1588);
nand U1655 (N_1655,N_1544,N_1522);
or U1656 (N_1656,N_1578,N_1543);
or U1657 (N_1657,N_1554,N_1507);
nor U1658 (N_1658,N_1514,N_1545);
or U1659 (N_1659,N_1539,N_1570);
nand U1660 (N_1660,N_1580,N_1514);
nand U1661 (N_1661,N_1516,N_1571);
nor U1662 (N_1662,N_1542,N_1507);
and U1663 (N_1663,N_1577,N_1559);
nand U1664 (N_1664,N_1557,N_1540);
nand U1665 (N_1665,N_1567,N_1518);
or U1666 (N_1666,N_1540,N_1533);
nor U1667 (N_1667,N_1547,N_1506);
or U1668 (N_1668,N_1578,N_1557);
or U1669 (N_1669,N_1575,N_1506);
or U1670 (N_1670,N_1501,N_1545);
and U1671 (N_1671,N_1526,N_1536);
or U1672 (N_1672,N_1531,N_1504);
nand U1673 (N_1673,N_1572,N_1547);
or U1674 (N_1674,N_1522,N_1500);
or U1675 (N_1675,N_1570,N_1579);
nand U1676 (N_1676,N_1556,N_1553);
and U1677 (N_1677,N_1500,N_1541);
nand U1678 (N_1678,N_1559,N_1504);
nand U1679 (N_1679,N_1546,N_1531);
nand U1680 (N_1680,N_1507,N_1525);
or U1681 (N_1681,N_1511,N_1582);
nor U1682 (N_1682,N_1556,N_1544);
nor U1683 (N_1683,N_1508,N_1557);
nand U1684 (N_1684,N_1578,N_1596);
nor U1685 (N_1685,N_1567,N_1595);
nor U1686 (N_1686,N_1576,N_1594);
nand U1687 (N_1687,N_1509,N_1566);
nand U1688 (N_1688,N_1594,N_1517);
or U1689 (N_1689,N_1585,N_1587);
and U1690 (N_1690,N_1505,N_1524);
nor U1691 (N_1691,N_1522,N_1513);
and U1692 (N_1692,N_1579,N_1587);
nand U1693 (N_1693,N_1518,N_1569);
or U1694 (N_1694,N_1528,N_1524);
nand U1695 (N_1695,N_1582,N_1521);
or U1696 (N_1696,N_1521,N_1569);
nor U1697 (N_1697,N_1541,N_1572);
and U1698 (N_1698,N_1558,N_1587);
nor U1699 (N_1699,N_1542,N_1533);
and U1700 (N_1700,N_1657,N_1665);
and U1701 (N_1701,N_1610,N_1603);
nand U1702 (N_1702,N_1695,N_1606);
nand U1703 (N_1703,N_1636,N_1649);
nor U1704 (N_1704,N_1645,N_1687);
or U1705 (N_1705,N_1647,N_1685);
or U1706 (N_1706,N_1644,N_1617);
and U1707 (N_1707,N_1611,N_1607);
xor U1708 (N_1708,N_1686,N_1650);
or U1709 (N_1709,N_1620,N_1662);
nand U1710 (N_1710,N_1683,N_1638);
or U1711 (N_1711,N_1697,N_1688);
nand U1712 (N_1712,N_1681,N_1653);
nor U1713 (N_1713,N_1671,N_1609);
and U1714 (N_1714,N_1663,N_1625);
or U1715 (N_1715,N_1693,N_1612);
or U1716 (N_1716,N_1623,N_1690);
and U1717 (N_1717,N_1602,N_1624);
nor U1718 (N_1718,N_1694,N_1627);
and U1719 (N_1719,N_1605,N_1670);
xor U1720 (N_1720,N_1646,N_1656);
or U1721 (N_1721,N_1613,N_1640);
and U1722 (N_1722,N_1633,N_1639);
nand U1723 (N_1723,N_1684,N_1641);
or U1724 (N_1724,N_1618,N_1619);
nand U1725 (N_1725,N_1635,N_1667);
and U1726 (N_1726,N_1673,N_1668);
and U1727 (N_1727,N_1608,N_1601);
or U1728 (N_1728,N_1634,N_1672);
or U1729 (N_1729,N_1626,N_1637);
nand U1730 (N_1730,N_1622,N_1628);
nor U1731 (N_1731,N_1691,N_1615);
and U1732 (N_1732,N_1614,N_1664);
and U1733 (N_1733,N_1696,N_1675);
nand U1734 (N_1734,N_1682,N_1629);
nand U1735 (N_1735,N_1674,N_1600);
and U1736 (N_1736,N_1648,N_1651);
nor U1737 (N_1737,N_1679,N_1692);
nor U1738 (N_1738,N_1616,N_1655);
and U1739 (N_1739,N_1631,N_1642);
nand U1740 (N_1740,N_1699,N_1643);
and U1741 (N_1741,N_1654,N_1669);
and U1742 (N_1742,N_1680,N_1621);
nor U1743 (N_1743,N_1678,N_1661);
and U1744 (N_1744,N_1666,N_1676);
nand U1745 (N_1745,N_1658,N_1604);
or U1746 (N_1746,N_1689,N_1632);
or U1747 (N_1747,N_1698,N_1677);
nand U1748 (N_1748,N_1660,N_1630);
nand U1749 (N_1749,N_1652,N_1659);
nand U1750 (N_1750,N_1660,N_1696);
nor U1751 (N_1751,N_1660,N_1680);
nand U1752 (N_1752,N_1600,N_1654);
and U1753 (N_1753,N_1666,N_1609);
nor U1754 (N_1754,N_1676,N_1619);
and U1755 (N_1755,N_1642,N_1635);
nand U1756 (N_1756,N_1646,N_1626);
nand U1757 (N_1757,N_1635,N_1611);
or U1758 (N_1758,N_1699,N_1658);
nor U1759 (N_1759,N_1697,N_1603);
nor U1760 (N_1760,N_1682,N_1600);
and U1761 (N_1761,N_1632,N_1678);
nor U1762 (N_1762,N_1698,N_1653);
nor U1763 (N_1763,N_1680,N_1692);
nor U1764 (N_1764,N_1635,N_1619);
nand U1765 (N_1765,N_1603,N_1636);
or U1766 (N_1766,N_1688,N_1637);
nor U1767 (N_1767,N_1642,N_1658);
nor U1768 (N_1768,N_1658,N_1635);
nor U1769 (N_1769,N_1664,N_1654);
nor U1770 (N_1770,N_1610,N_1627);
nand U1771 (N_1771,N_1649,N_1677);
or U1772 (N_1772,N_1673,N_1642);
nand U1773 (N_1773,N_1620,N_1671);
nand U1774 (N_1774,N_1632,N_1629);
and U1775 (N_1775,N_1676,N_1629);
nand U1776 (N_1776,N_1694,N_1685);
or U1777 (N_1777,N_1621,N_1637);
nor U1778 (N_1778,N_1665,N_1607);
nand U1779 (N_1779,N_1663,N_1623);
nor U1780 (N_1780,N_1653,N_1619);
or U1781 (N_1781,N_1683,N_1670);
nor U1782 (N_1782,N_1668,N_1651);
nand U1783 (N_1783,N_1602,N_1626);
nor U1784 (N_1784,N_1649,N_1668);
nand U1785 (N_1785,N_1682,N_1693);
and U1786 (N_1786,N_1665,N_1606);
and U1787 (N_1787,N_1645,N_1651);
nand U1788 (N_1788,N_1670,N_1629);
nand U1789 (N_1789,N_1625,N_1607);
or U1790 (N_1790,N_1687,N_1693);
nor U1791 (N_1791,N_1687,N_1628);
and U1792 (N_1792,N_1694,N_1608);
nor U1793 (N_1793,N_1675,N_1698);
or U1794 (N_1794,N_1624,N_1695);
and U1795 (N_1795,N_1643,N_1646);
nand U1796 (N_1796,N_1653,N_1622);
and U1797 (N_1797,N_1693,N_1657);
nor U1798 (N_1798,N_1651,N_1698);
nand U1799 (N_1799,N_1683,N_1665);
or U1800 (N_1800,N_1728,N_1762);
or U1801 (N_1801,N_1710,N_1752);
nor U1802 (N_1802,N_1791,N_1787);
or U1803 (N_1803,N_1753,N_1749);
nor U1804 (N_1804,N_1764,N_1788);
or U1805 (N_1805,N_1724,N_1735);
nand U1806 (N_1806,N_1755,N_1777);
nand U1807 (N_1807,N_1763,N_1797);
or U1808 (N_1808,N_1712,N_1718);
nand U1809 (N_1809,N_1727,N_1746);
nor U1810 (N_1810,N_1775,N_1737);
nand U1811 (N_1811,N_1780,N_1731);
nand U1812 (N_1812,N_1756,N_1717);
nand U1813 (N_1813,N_1748,N_1771);
nand U1814 (N_1814,N_1734,N_1706);
or U1815 (N_1815,N_1740,N_1751);
nand U1816 (N_1816,N_1736,N_1704);
or U1817 (N_1817,N_1725,N_1790);
nand U1818 (N_1818,N_1719,N_1792);
nand U1819 (N_1819,N_1742,N_1744);
and U1820 (N_1820,N_1723,N_1721);
nor U1821 (N_1821,N_1781,N_1714);
and U1822 (N_1822,N_1758,N_1711);
nor U1823 (N_1823,N_1769,N_1702);
and U1824 (N_1824,N_1754,N_1761);
nor U1825 (N_1825,N_1703,N_1715);
and U1826 (N_1826,N_1733,N_1778);
xor U1827 (N_1827,N_1794,N_1765);
nor U1828 (N_1828,N_1779,N_1705);
nand U1829 (N_1829,N_1750,N_1716);
nor U1830 (N_1830,N_1783,N_1770);
nor U1831 (N_1831,N_1768,N_1726);
or U1832 (N_1832,N_1707,N_1709);
nand U1833 (N_1833,N_1789,N_1730);
and U1834 (N_1834,N_1798,N_1759);
and U1835 (N_1835,N_1776,N_1700);
and U1836 (N_1836,N_1738,N_1773);
nand U1837 (N_1837,N_1766,N_1729);
and U1838 (N_1838,N_1722,N_1774);
and U1839 (N_1839,N_1757,N_1795);
nand U1840 (N_1840,N_1701,N_1785);
nor U1841 (N_1841,N_1741,N_1782);
nor U1842 (N_1842,N_1720,N_1747);
nand U1843 (N_1843,N_1732,N_1784);
and U1844 (N_1844,N_1745,N_1760);
nand U1845 (N_1845,N_1743,N_1713);
nand U1846 (N_1846,N_1796,N_1708);
or U1847 (N_1847,N_1786,N_1793);
and U1848 (N_1848,N_1799,N_1739);
and U1849 (N_1849,N_1772,N_1767);
nor U1850 (N_1850,N_1795,N_1754);
or U1851 (N_1851,N_1775,N_1757);
and U1852 (N_1852,N_1781,N_1713);
or U1853 (N_1853,N_1762,N_1722);
nor U1854 (N_1854,N_1719,N_1744);
and U1855 (N_1855,N_1721,N_1771);
nor U1856 (N_1856,N_1731,N_1712);
and U1857 (N_1857,N_1792,N_1734);
nand U1858 (N_1858,N_1750,N_1721);
or U1859 (N_1859,N_1729,N_1797);
or U1860 (N_1860,N_1775,N_1739);
or U1861 (N_1861,N_1724,N_1752);
nor U1862 (N_1862,N_1732,N_1700);
and U1863 (N_1863,N_1744,N_1788);
nand U1864 (N_1864,N_1771,N_1779);
and U1865 (N_1865,N_1778,N_1732);
and U1866 (N_1866,N_1793,N_1785);
nor U1867 (N_1867,N_1766,N_1786);
nor U1868 (N_1868,N_1757,N_1781);
nor U1869 (N_1869,N_1702,N_1796);
and U1870 (N_1870,N_1794,N_1795);
and U1871 (N_1871,N_1703,N_1706);
and U1872 (N_1872,N_1745,N_1732);
nor U1873 (N_1873,N_1780,N_1747);
nand U1874 (N_1874,N_1779,N_1707);
and U1875 (N_1875,N_1763,N_1709);
or U1876 (N_1876,N_1743,N_1710);
or U1877 (N_1877,N_1701,N_1764);
nor U1878 (N_1878,N_1745,N_1722);
nor U1879 (N_1879,N_1734,N_1750);
nand U1880 (N_1880,N_1783,N_1710);
nor U1881 (N_1881,N_1718,N_1722);
and U1882 (N_1882,N_1795,N_1788);
nor U1883 (N_1883,N_1750,N_1789);
and U1884 (N_1884,N_1752,N_1708);
nor U1885 (N_1885,N_1709,N_1761);
or U1886 (N_1886,N_1796,N_1762);
nor U1887 (N_1887,N_1757,N_1778);
nor U1888 (N_1888,N_1733,N_1706);
and U1889 (N_1889,N_1729,N_1709);
or U1890 (N_1890,N_1775,N_1771);
nand U1891 (N_1891,N_1718,N_1705);
nand U1892 (N_1892,N_1742,N_1767);
nand U1893 (N_1893,N_1711,N_1736);
nor U1894 (N_1894,N_1790,N_1799);
and U1895 (N_1895,N_1743,N_1738);
or U1896 (N_1896,N_1759,N_1777);
nor U1897 (N_1897,N_1742,N_1751);
nand U1898 (N_1898,N_1784,N_1701);
nor U1899 (N_1899,N_1718,N_1744);
and U1900 (N_1900,N_1896,N_1802);
and U1901 (N_1901,N_1884,N_1815);
nand U1902 (N_1902,N_1804,N_1876);
nand U1903 (N_1903,N_1806,N_1808);
or U1904 (N_1904,N_1854,N_1810);
and U1905 (N_1905,N_1897,N_1841);
or U1906 (N_1906,N_1843,N_1838);
or U1907 (N_1907,N_1893,N_1831);
nor U1908 (N_1908,N_1875,N_1823);
nand U1909 (N_1909,N_1847,N_1842);
and U1910 (N_1910,N_1826,N_1874);
or U1911 (N_1911,N_1818,N_1898);
and U1912 (N_1912,N_1828,N_1836);
and U1913 (N_1913,N_1853,N_1824);
nor U1914 (N_1914,N_1861,N_1873);
xor U1915 (N_1915,N_1800,N_1850);
nor U1916 (N_1916,N_1811,N_1890);
nand U1917 (N_1917,N_1885,N_1868);
nand U1918 (N_1918,N_1886,N_1872);
and U1919 (N_1919,N_1805,N_1870);
or U1920 (N_1920,N_1863,N_1877);
nand U1921 (N_1921,N_1892,N_1899);
and U1922 (N_1922,N_1867,N_1801);
nor U1923 (N_1923,N_1840,N_1888);
and U1924 (N_1924,N_1871,N_1803);
nand U1925 (N_1925,N_1862,N_1835);
nor U1926 (N_1926,N_1887,N_1839);
or U1927 (N_1927,N_1866,N_1851);
or U1928 (N_1928,N_1878,N_1837);
nor U1929 (N_1929,N_1889,N_1879);
or U1930 (N_1930,N_1844,N_1807);
and U1931 (N_1931,N_1852,N_1881);
nor U1932 (N_1932,N_1829,N_1819);
and U1933 (N_1933,N_1834,N_1858);
and U1934 (N_1934,N_1812,N_1895);
nor U1935 (N_1935,N_1827,N_1833);
nor U1936 (N_1936,N_1865,N_1816);
nand U1937 (N_1937,N_1857,N_1830);
or U1938 (N_1938,N_1894,N_1860);
nor U1939 (N_1939,N_1880,N_1849);
and U1940 (N_1940,N_1817,N_1809);
nor U1941 (N_1941,N_1813,N_1814);
and U1942 (N_1942,N_1882,N_1825);
nor U1943 (N_1943,N_1820,N_1864);
nor U1944 (N_1944,N_1869,N_1832);
or U1945 (N_1945,N_1848,N_1855);
nor U1946 (N_1946,N_1821,N_1891);
nand U1947 (N_1947,N_1856,N_1883);
and U1948 (N_1948,N_1822,N_1846);
nand U1949 (N_1949,N_1845,N_1859);
nand U1950 (N_1950,N_1841,N_1842);
nand U1951 (N_1951,N_1812,N_1869);
and U1952 (N_1952,N_1849,N_1800);
or U1953 (N_1953,N_1823,N_1877);
or U1954 (N_1954,N_1853,N_1815);
and U1955 (N_1955,N_1824,N_1848);
or U1956 (N_1956,N_1814,N_1857);
nor U1957 (N_1957,N_1804,N_1843);
nand U1958 (N_1958,N_1835,N_1849);
nand U1959 (N_1959,N_1854,N_1887);
nand U1960 (N_1960,N_1862,N_1802);
nor U1961 (N_1961,N_1899,N_1850);
nor U1962 (N_1962,N_1880,N_1897);
and U1963 (N_1963,N_1888,N_1811);
and U1964 (N_1964,N_1807,N_1891);
and U1965 (N_1965,N_1837,N_1811);
or U1966 (N_1966,N_1850,N_1837);
nor U1967 (N_1967,N_1830,N_1865);
and U1968 (N_1968,N_1867,N_1800);
or U1969 (N_1969,N_1896,N_1817);
and U1970 (N_1970,N_1844,N_1858);
nand U1971 (N_1971,N_1870,N_1874);
nand U1972 (N_1972,N_1879,N_1804);
or U1973 (N_1973,N_1886,N_1821);
or U1974 (N_1974,N_1816,N_1820);
nand U1975 (N_1975,N_1893,N_1833);
nand U1976 (N_1976,N_1853,N_1828);
or U1977 (N_1977,N_1891,N_1887);
nor U1978 (N_1978,N_1882,N_1852);
or U1979 (N_1979,N_1833,N_1849);
nor U1980 (N_1980,N_1842,N_1845);
or U1981 (N_1981,N_1852,N_1893);
or U1982 (N_1982,N_1863,N_1823);
or U1983 (N_1983,N_1880,N_1823);
and U1984 (N_1984,N_1843,N_1858);
nand U1985 (N_1985,N_1888,N_1895);
nor U1986 (N_1986,N_1893,N_1860);
and U1987 (N_1987,N_1839,N_1801);
nand U1988 (N_1988,N_1843,N_1865);
nor U1989 (N_1989,N_1845,N_1899);
and U1990 (N_1990,N_1838,N_1852);
nor U1991 (N_1991,N_1832,N_1811);
and U1992 (N_1992,N_1863,N_1843);
nor U1993 (N_1993,N_1831,N_1833);
nand U1994 (N_1994,N_1832,N_1864);
nor U1995 (N_1995,N_1877,N_1853);
or U1996 (N_1996,N_1820,N_1843);
or U1997 (N_1997,N_1803,N_1870);
nand U1998 (N_1998,N_1832,N_1862);
and U1999 (N_1999,N_1847,N_1802);
or U2000 (N_2000,N_1975,N_1976);
nor U2001 (N_2001,N_1929,N_1954);
or U2002 (N_2002,N_1965,N_1978);
and U2003 (N_2003,N_1916,N_1909);
nor U2004 (N_2004,N_1987,N_1932);
nand U2005 (N_2005,N_1947,N_1927);
or U2006 (N_2006,N_1912,N_1900);
nor U2007 (N_2007,N_1918,N_1949);
nand U2008 (N_2008,N_1911,N_1951);
nand U2009 (N_2009,N_1950,N_1917);
nand U2010 (N_2010,N_1944,N_1923);
or U2011 (N_2011,N_1968,N_1983);
nand U2012 (N_2012,N_1902,N_1963);
nor U2013 (N_2013,N_1933,N_1919);
and U2014 (N_2014,N_1939,N_1980);
or U2015 (N_2015,N_1967,N_1989);
and U2016 (N_2016,N_1931,N_1942);
and U2017 (N_2017,N_1990,N_1937);
or U2018 (N_2018,N_1910,N_1940);
or U2019 (N_2019,N_1999,N_1984);
or U2020 (N_2020,N_1908,N_1958);
or U2021 (N_2021,N_1998,N_1921);
nor U2022 (N_2022,N_1982,N_1973);
nand U2023 (N_2023,N_1903,N_1991);
and U2024 (N_2024,N_1934,N_1981);
nand U2025 (N_2025,N_1995,N_1959);
or U2026 (N_2026,N_1926,N_1948);
nand U2027 (N_2027,N_1985,N_1936);
nand U2028 (N_2028,N_1966,N_1946);
or U2029 (N_2029,N_1920,N_1935);
and U2030 (N_2030,N_1977,N_1955);
or U2031 (N_2031,N_1924,N_1906);
and U2032 (N_2032,N_1964,N_1996);
or U2033 (N_2033,N_1904,N_1960);
and U2034 (N_2034,N_1938,N_1992);
nand U2035 (N_2035,N_1928,N_1979);
nor U2036 (N_2036,N_1997,N_1974);
nor U2037 (N_2037,N_1969,N_1972);
or U2038 (N_2038,N_1993,N_1953);
and U2039 (N_2039,N_1971,N_1914);
nor U2040 (N_2040,N_1915,N_1905);
or U2041 (N_2041,N_1988,N_1930);
nand U2042 (N_2042,N_1957,N_1970);
and U2043 (N_2043,N_1922,N_1907);
and U2044 (N_2044,N_1941,N_1986);
or U2045 (N_2045,N_1961,N_1901);
and U2046 (N_2046,N_1956,N_1913);
nand U2047 (N_2047,N_1925,N_1945);
and U2048 (N_2048,N_1952,N_1994);
and U2049 (N_2049,N_1943,N_1962);
nand U2050 (N_2050,N_1901,N_1942);
nor U2051 (N_2051,N_1929,N_1952);
nor U2052 (N_2052,N_1942,N_1927);
and U2053 (N_2053,N_1962,N_1947);
nand U2054 (N_2054,N_1965,N_1921);
nor U2055 (N_2055,N_1934,N_1950);
and U2056 (N_2056,N_1908,N_1947);
and U2057 (N_2057,N_1985,N_1935);
nand U2058 (N_2058,N_1921,N_1909);
or U2059 (N_2059,N_1960,N_1966);
nor U2060 (N_2060,N_1921,N_1912);
and U2061 (N_2061,N_1924,N_1980);
nor U2062 (N_2062,N_1928,N_1931);
or U2063 (N_2063,N_1999,N_1908);
nor U2064 (N_2064,N_1961,N_1960);
nor U2065 (N_2065,N_1976,N_1972);
nand U2066 (N_2066,N_1956,N_1929);
and U2067 (N_2067,N_1981,N_1917);
nand U2068 (N_2068,N_1926,N_1933);
or U2069 (N_2069,N_1916,N_1913);
and U2070 (N_2070,N_1916,N_1956);
and U2071 (N_2071,N_1901,N_1928);
nor U2072 (N_2072,N_1996,N_1954);
or U2073 (N_2073,N_1978,N_1921);
or U2074 (N_2074,N_1994,N_1958);
or U2075 (N_2075,N_1910,N_1943);
nor U2076 (N_2076,N_1983,N_1927);
nand U2077 (N_2077,N_1960,N_1972);
nor U2078 (N_2078,N_1948,N_1916);
or U2079 (N_2079,N_1916,N_1900);
nor U2080 (N_2080,N_1996,N_1948);
and U2081 (N_2081,N_1950,N_1923);
and U2082 (N_2082,N_1984,N_1962);
or U2083 (N_2083,N_1977,N_1979);
nand U2084 (N_2084,N_1938,N_1903);
nor U2085 (N_2085,N_1968,N_1922);
nor U2086 (N_2086,N_1915,N_1948);
or U2087 (N_2087,N_1910,N_1923);
or U2088 (N_2088,N_1955,N_1913);
xor U2089 (N_2089,N_1918,N_1902);
nor U2090 (N_2090,N_1997,N_1925);
nand U2091 (N_2091,N_1917,N_1913);
or U2092 (N_2092,N_1920,N_1930);
xor U2093 (N_2093,N_1973,N_1903);
nor U2094 (N_2094,N_1981,N_1919);
and U2095 (N_2095,N_1950,N_1963);
nor U2096 (N_2096,N_1942,N_1967);
nor U2097 (N_2097,N_1916,N_1911);
or U2098 (N_2098,N_1973,N_1905);
nand U2099 (N_2099,N_1957,N_1950);
nor U2100 (N_2100,N_2089,N_2069);
nand U2101 (N_2101,N_2033,N_2027);
nor U2102 (N_2102,N_2060,N_2042);
nand U2103 (N_2103,N_2016,N_2023);
and U2104 (N_2104,N_2072,N_2007);
nand U2105 (N_2105,N_2077,N_2034);
or U2106 (N_2106,N_2006,N_2012);
nor U2107 (N_2107,N_2078,N_2085);
nor U2108 (N_2108,N_2049,N_2010);
nand U2109 (N_2109,N_2079,N_2032);
nand U2110 (N_2110,N_2075,N_2059);
and U2111 (N_2111,N_2050,N_2044);
and U2112 (N_2112,N_2009,N_2003);
nor U2113 (N_2113,N_2028,N_2091);
and U2114 (N_2114,N_2064,N_2074);
nand U2115 (N_2115,N_2039,N_2002);
nand U2116 (N_2116,N_2022,N_2057);
and U2117 (N_2117,N_2013,N_2030);
and U2118 (N_2118,N_2004,N_2025);
nand U2119 (N_2119,N_2058,N_2036);
or U2120 (N_2120,N_2056,N_2073);
or U2121 (N_2121,N_2063,N_2037);
nand U2122 (N_2122,N_2005,N_2043);
nand U2123 (N_2123,N_2094,N_2082);
or U2124 (N_2124,N_2061,N_2019);
nand U2125 (N_2125,N_2029,N_2031);
nor U2126 (N_2126,N_2015,N_2052);
or U2127 (N_2127,N_2098,N_2035);
or U2128 (N_2128,N_2095,N_2097);
and U2129 (N_2129,N_2099,N_2070);
or U2130 (N_2130,N_2020,N_2011);
nand U2131 (N_2131,N_2071,N_2076);
or U2132 (N_2132,N_2038,N_2018);
or U2133 (N_2133,N_2080,N_2088);
nor U2134 (N_2134,N_2024,N_2026);
nand U2135 (N_2135,N_2086,N_2041);
nand U2136 (N_2136,N_2001,N_2096);
nor U2137 (N_2137,N_2055,N_2067);
nor U2138 (N_2138,N_2046,N_2017);
and U2139 (N_2139,N_2051,N_2092);
and U2140 (N_2140,N_2084,N_2083);
nand U2141 (N_2141,N_2040,N_2021);
nor U2142 (N_2142,N_2068,N_2048);
nor U2143 (N_2143,N_2090,N_2093);
nand U2144 (N_2144,N_2054,N_2045);
or U2145 (N_2145,N_2087,N_2081);
nand U2146 (N_2146,N_2062,N_2065);
and U2147 (N_2147,N_2000,N_2014);
and U2148 (N_2148,N_2008,N_2053);
nand U2149 (N_2149,N_2047,N_2066);
or U2150 (N_2150,N_2015,N_2051);
nor U2151 (N_2151,N_2060,N_2083);
or U2152 (N_2152,N_2070,N_2015);
or U2153 (N_2153,N_2075,N_2025);
or U2154 (N_2154,N_2046,N_2033);
nand U2155 (N_2155,N_2071,N_2043);
nor U2156 (N_2156,N_2056,N_2018);
nand U2157 (N_2157,N_2013,N_2012);
nand U2158 (N_2158,N_2068,N_2069);
nand U2159 (N_2159,N_2086,N_2066);
nand U2160 (N_2160,N_2035,N_2003);
nand U2161 (N_2161,N_2084,N_2071);
nand U2162 (N_2162,N_2085,N_2001);
nor U2163 (N_2163,N_2067,N_2049);
nor U2164 (N_2164,N_2009,N_2010);
or U2165 (N_2165,N_2068,N_2025);
and U2166 (N_2166,N_2011,N_2053);
nor U2167 (N_2167,N_2003,N_2097);
nand U2168 (N_2168,N_2000,N_2088);
nor U2169 (N_2169,N_2003,N_2039);
nand U2170 (N_2170,N_2022,N_2091);
nand U2171 (N_2171,N_2064,N_2091);
and U2172 (N_2172,N_2039,N_2085);
or U2173 (N_2173,N_2026,N_2065);
nand U2174 (N_2174,N_2046,N_2095);
nand U2175 (N_2175,N_2040,N_2003);
nor U2176 (N_2176,N_2071,N_2042);
or U2177 (N_2177,N_2076,N_2093);
nor U2178 (N_2178,N_2094,N_2073);
and U2179 (N_2179,N_2049,N_2094);
nor U2180 (N_2180,N_2062,N_2056);
or U2181 (N_2181,N_2099,N_2054);
nor U2182 (N_2182,N_2056,N_2069);
nor U2183 (N_2183,N_2015,N_2046);
nor U2184 (N_2184,N_2057,N_2070);
nor U2185 (N_2185,N_2021,N_2004);
or U2186 (N_2186,N_2023,N_2035);
nor U2187 (N_2187,N_2067,N_2089);
nand U2188 (N_2188,N_2084,N_2070);
nand U2189 (N_2189,N_2053,N_2056);
nand U2190 (N_2190,N_2075,N_2061);
and U2191 (N_2191,N_2081,N_2021);
and U2192 (N_2192,N_2096,N_2053);
and U2193 (N_2193,N_2071,N_2026);
xnor U2194 (N_2194,N_2017,N_2009);
xor U2195 (N_2195,N_2012,N_2054);
or U2196 (N_2196,N_2019,N_2001);
nand U2197 (N_2197,N_2017,N_2032);
nand U2198 (N_2198,N_2002,N_2005);
nor U2199 (N_2199,N_2053,N_2065);
nand U2200 (N_2200,N_2109,N_2151);
and U2201 (N_2201,N_2197,N_2168);
nand U2202 (N_2202,N_2100,N_2160);
or U2203 (N_2203,N_2195,N_2154);
nor U2204 (N_2204,N_2117,N_2174);
nor U2205 (N_2205,N_2133,N_2176);
nand U2206 (N_2206,N_2136,N_2166);
or U2207 (N_2207,N_2182,N_2131);
or U2208 (N_2208,N_2145,N_2191);
nand U2209 (N_2209,N_2164,N_2186);
nand U2210 (N_2210,N_2193,N_2121);
and U2211 (N_2211,N_2125,N_2127);
and U2212 (N_2212,N_2188,N_2138);
nor U2213 (N_2213,N_2135,N_2144);
and U2214 (N_2214,N_2115,N_2167);
or U2215 (N_2215,N_2140,N_2155);
and U2216 (N_2216,N_2190,N_2134);
and U2217 (N_2217,N_2104,N_2194);
nor U2218 (N_2218,N_2184,N_2106);
xnor U2219 (N_2219,N_2108,N_2139);
nand U2220 (N_2220,N_2119,N_2185);
or U2221 (N_2221,N_2142,N_2170);
or U2222 (N_2222,N_2177,N_2178);
or U2223 (N_2223,N_2180,N_2105);
or U2224 (N_2224,N_2149,N_2156);
and U2225 (N_2225,N_2124,N_2152);
nor U2226 (N_2226,N_2126,N_2111);
nor U2227 (N_2227,N_2162,N_2116);
nand U2228 (N_2228,N_2132,N_2196);
and U2229 (N_2229,N_2147,N_2113);
nor U2230 (N_2230,N_2128,N_2129);
nand U2231 (N_2231,N_2173,N_2102);
nor U2232 (N_2232,N_2181,N_2199);
and U2233 (N_2233,N_2183,N_2143);
nand U2234 (N_2234,N_2171,N_2112);
nor U2235 (N_2235,N_2123,N_2158);
and U2236 (N_2236,N_2175,N_2157);
nor U2237 (N_2237,N_2198,N_2148);
nor U2238 (N_2238,N_2179,N_2118);
nand U2239 (N_2239,N_2172,N_2122);
and U2240 (N_2240,N_2150,N_2107);
nor U2241 (N_2241,N_2141,N_2110);
nand U2242 (N_2242,N_2163,N_2114);
or U2243 (N_2243,N_2153,N_2101);
nor U2244 (N_2244,N_2165,N_2130);
nor U2245 (N_2245,N_2192,N_2103);
and U2246 (N_2246,N_2137,N_2120);
and U2247 (N_2247,N_2146,N_2187);
and U2248 (N_2248,N_2161,N_2159);
or U2249 (N_2249,N_2169,N_2189);
and U2250 (N_2250,N_2187,N_2159);
and U2251 (N_2251,N_2181,N_2106);
nor U2252 (N_2252,N_2116,N_2138);
or U2253 (N_2253,N_2131,N_2149);
nor U2254 (N_2254,N_2117,N_2160);
or U2255 (N_2255,N_2172,N_2153);
nand U2256 (N_2256,N_2170,N_2174);
nor U2257 (N_2257,N_2130,N_2105);
nand U2258 (N_2258,N_2188,N_2136);
or U2259 (N_2259,N_2149,N_2128);
or U2260 (N_2260,N_2132,N_2148);
nand U2261 (N_2261,N_2161,N_2143);
or U2262 (N_2262,N_2197,N_2127);
nor U2263 (N_2263,N_2145,N_2129);
or U2264 (N_2264,N_2154,N_2156);
nor U2265 (N_2265,N_2162,N_2165);
nand U2266 (N_2266,N_2162,N_2199);
and U2267 (N_2267,N_2196,N_2197);
xnor U2268 (N_2268,N_2176,N_2193);
nand U2269 (N_2269,N_2152,N_2111);
nor U2270 (N_2270,N_2173,N_2136);
nor U2271 (N_2271,N_2180,N_2106);
nand U2272 (N_2272,N_2125,N_2187);
nor U2273 (N_2273,N_2132,N_2195);
nand U2274 (N_2274,N_2157,N_2176);
and U2275 (N_2275,N_2154,N_2187);
and U2276 (N_2276,N_2160,N_2170);
and U2277 (N_2277,N_2142,N_2194);
or U2278 (N_2278,N_2109,N_2113);
or U2279 (N_2279,N_2155,N_2112);
and U2280 (N_2280,N_2163,N_2154);
or U2281 (N_2281,N_2127,N_2155);
nor U2282 (N_2282,N_2162,N_2107);
or U2283 (N_2283,N_2148,N_2118);
and U2284 (N_2284,N_2108,N_2135);
nand U2285 (N_2285,N_2191,N_2152);
or U2286 (N_2286,N_2194,N_2137);
or U2287 (N_2287,N_2113,N_2178);
or U2288 (N_2288,N_2118,N_2109);
and U2289 (N_2289,N_2122,N_2102);
nand U2290 (N_2290,N_2157,N_2111);
nand U2291 (N_2291,N_2163,N_2128);
nor U2292 (N_2292,N_2156,N_2195);
nand U2293 (N_2293,N_2113,N_2138);
or U2294 (N_2294,N_2199,N_2118);
and U2295 (N_2295,N_2188,N_2191);
or U2296 (N_2296,N_2178,N_2116);
and U2297 (N_2297,N_2115,N_2171);
nor U2298 (N_2298,N_2113,N_2128);
nor U2299 (N_2299,N_2147,N_2159);
nor U2300 (N_2300,N_2270,N_2287);
nand U2301 (N_2301,N_2250,N_2204);
and U2302 (N_2302,N_2289,N_2246);
nand U2303 (N_2303,N_2249,N_2245);
or U2304 (N_2304,N_2278,N_2206);
nor U2305 (N_2305,N_2213,N_2228);
or U2306 (N_2306,N_2294,N_2219);
and U2307 (N_2307,N_2276,N_2247);
nand U2308 (N_2308,N_2293,N_2282);
nand U2309 (N_2309,N_2243,N_2272);
nand U2310 (N_2310,N_2281,N_2223);
or U2311 (N_2311,N_2200,N_2214);
nand U2312 (N_2312,N_2296,N_2216);
or U2313 (N_2313,N_2222,N_2238);
and U2314 (N_2314,N_2234,N_2207);
nor U2315 (N_2315,N_2298,N_2210);
or U2316 (N_2316,N_2221,N_2224);
or U2317 (N_2317,N_2226,N_2274);
and U2318 (N_2318,N_2218,N_2215);
or U2319 (N_2319,N_2261,N_2286);
or U2320 (N_2320,N_2241,N_2255);
nor U2321 (N_2321,N_2288,N_2225);
nor U2322 (N_2322,N_2217,N_2230);
xnor U2323 (N_2323,N_2208,N_2205);
nand U2324 (N_2324,N_2201,N_2229);
nor U2325 (N_2325,N_2236,N_2269);
xor U2326 (N_2326,N_2257,N_2231);
nor U2327 (N_2327,N_2254,N_2283);
nand U2328 (N_2328,N_2299,N_2290);
nand U2329 (N_2329,N_2291,N_2237);
or U2330 (N_2330,N_2256,N_2233);
and U2331 (N_2331,N_2292,N_2267);
or U2332 (N_2332,N_2297,N_2244);
nand U2333 (N_2333,N_2259,N_2248);
or U2334 (N_2334,N_2262,N_2284);
nand U2335 (N_2335,N_2279,N_2251);
nor U2336 (N_2336,N_2266,N_2209);
nor U2337 (N_2337,N_2227,N_2263);
nor U2338 (N_2338,N_2268,N_2275);
and U2339 (N_2339,N_2211,N_2212);
nor U2340 (N_2340,N_2260,N_2280);
nor U2341 (N_2341,N_2240,N_2220);
nor U2342 (N_2342,N_2239,N_2271);
or U2343 (N_2343,N_2252,N_2232);
nand U2344 (N_2344,N_2258,N_2285);
nand U2345 (N_2345,N_2264,N_2235);
nor U2346 (N_2346,N_2265,N_2295);
or U2347 (N_2347,N_2253,N_2203);
nor U2348 (N_2348,N_2242,N_2273);
nand U2349 (N_2349,N_2202,N_2277);
nand U2350 (N_2350,N_2285,N_2207);
nor U2351 (N_2351,N_2220,N_2215);
and U2352 (N_2352,N_2200,N_2264);
nand U2353 (N_2353,N_2231,N_2225);
or U2354 (N_2354,N_2270,N_2292);
or U2355 (N_2355,N_2248,N_2265);
and U2356 (N_2356,N_2246,N_2290);
nor U2357 (N_2357,N_2216,N_2243);
nand U2358 (N_2358,N_2241,N_2257);
nand U2359 (N_2359,N_2265,N_2280);
nand U2360 (N_2360,N_2271,N_2284);
and U2361 (N_2361,N_2282,N_2262);
xor U2362 (N_2362,N_2201,N_2248);
nand U2363 (N_2363,N_2293,N_2260);
and U2364 (N_2364,N_2276,N_2241);
nand U2365 (N_2365,N_2226,N_2218);
nor U2366 (N_2366,N_2206,N_2269);
or U2367 (N_2367,N_2270,N_2200);
or U2368 (N_2368,N_2234,N_2266);
nor U2369 (N_2369,N_2246,N_2230);
and U2370 (N_2370,N_2228,N_2254);
nand U2371 (N_2371,N_2260,N_2269);
and U2372 (N_2372,N_2237,N_2200);
nor U2373 (N_2373,N_2256,N_2240);
and U2374 (N_2374,N_2244,N_2266);
nand U2375 (N_2375,N_2215,N_2273);
nand U2376 (N_2376,N_2250,N_2296);
nor U2377 (N_2377,N_2290,N_2259);
or U2378 (N_2378,N_2273,N_2290);
nor U2379 (N_2379,N_2237,N_2238);
and U2380 (N_2380,N_2249,N_2227);
or U2381 (N_2381,N_2257,N_2283);
or U2382 (N_2382,N_2239,N_2235);
nor U2383 (N_2383,N_2206,N_2256);
nor U2384 (N_2384,N_2225,N_2282);
or U2385 (N_2385,N_2239,N_2205);
nand U2386 (N_2386,N_2276,N_2204);
xnor U2387 (N_2387,N_2258,N_2230);
nand U2388 (N_2388,N_2219,N_2243);
and U2389 (N_2389,N_2248,N_2217);
nor U2390 (N_2390,N_2223,N_2205);
or U2391 (N_2391,N_2214,N_2209);
nand U2392 (N_2392,N_2262,N_2203);
nand U2393 (N_2393,N_2231,N_2290);
or U2394 (N_2394,N_2274,N_2289);
nand U2395 (N_2395,N_2247,N_2236);
nor U2396 (N_2396,N_2224,N_2212);
nor U2397 (N_2397,N_2270,N_2254);
nor U2398 (N_2398,N_2257,N_2239);
and U2399 (N_2399,N_2282,N_2202);
or U2400 (N_2400,N_2376,N_2304);
nor U2401 (N_2401,N_2339,N_2360);
or U2402 (N_2402,N_2393,N_2323);
nand U2403 (N_2403,N_2301,N_2356);
and U2404 (N_2404,N_2395,N_2315);
nand U2405 (N_2405,N_2374,N_2385);
or U2406 (N_2406,N_2392,N_2319);
and U2407 (N_2407,N_2316,N_2357);
nor U2408 (N_2408,N_2305,N_2353);
or U2409 (N_2409,N_2350,N_2358);
nand U2410 (N_2410,N_2372,N_2344);
nor U2411 (N_2411,N_2382,N_2387);
nor U2412 (N_2412,N_2333,N_2329);
nor U2413 (N_2413,N_2306,N_2310);
nand U2414 (N_2414,N_2379,N_2377);
nand U2415 (N_2415,N_2375,N_2390);
nor U2416 (N_2416,N_2332,N_2326);
and U2417 (N_2417,N_2321,N_2336);
or U2418 (N_2418,N_2368,N_2364);
and U2419 (N_2419,N_2383,N_2359);
nand U2420 (N_2420,N_2361,N_2328);
nand U2421 (N_2421,N_2346,N_2363);
or U2422 (N_2422,N_2380,N_2327);
or U2423 (N_2423,N_2345,N_2320);
nand U2424 (N_2424,N_2352,N_2355);
nand U2425 (N_2425,N_2334,N_2307);
or U2426 (N_2426,N_2348,N_2351);
or U2427 (N_2427,N_2386,N_2391);
and U2428 (N_2428,N_2384,N_2300);
nand U2429 (N_2429,N_2343,N_2325);
nand U2430 (N_2430,N_2318,N_2366);
xnor U2431 (N_2431,N_2396,N_2331);
nand U2432 (N_2432,N_2308,N_2309);
or U2433 (N_2433,N_2330,N_2378);
nor U2434 (N_2434,N_2373,N_2317);
or U2435 (N_2435,N_2312,N_2371);
or U2436 (N_2436,N_2399,N_2313);
nand U2437 (N_2437,N_2389,N_2367);
and U2438 (N_2438,N_2311,N_2388);
nand U2439 (N_2439,N_2397,N_2381);
nand U2440 (N_2440,N_2342,N_2303);
and U2441 (N_2441,N_2349,N_2341);
and U2442 (N_2442,N_2340,N_2338);
nor U2443 (N_2443,N_2362,N_2347);
nand U2444 (N_2444,N_2335,N_2370);
and U2445 (N_2445,N_2398,N_2337);
or U2446 (N_2446,N_2354,N_2314);
and U2447 (N_2447,N_2394,N_2365);
or U2448 (N_2448,N_2322,N_2302);
nand U2449 (N_2449,N_2369,N_2324);
and U2450 (N_2450,N_2371,N_2384);
nand U2451 (N_2451,N_2353,N_2352);
nand U2452 (N_2452,N_2303,N_2335);
nand U2453 (N_2453,N_2359,N_2339);
or U2454 (N_2454,N_2331,N_2312);
nor U2455 (N_2455,N_2366,N_2337);
nand U2456 (N_2456,N_2302,N_2313);
nand U2457 (N_2457,N_2357,N_2325);
nand U2458 (N_2458,N_2383,N_2338);
and U2459 (N_2459,N_2342,N_2331);
nor U2460 (N_2460,N_2359,N_2375);
nand U2461 (N_2461,N_2367,N_2368);
or U2462 (N_2462,N_2348,N_2345);
nand U2463 (N_2463,N_2333,N_2379);
or U2464 (N_2464,N_2369,N_2381);
and U2465 (N_2465,N_2302,N_2380);
nor U2466 (N_2466,N_2368,N_2331);
or U2467 (N_2467,N_2322,N_2395);
or U2468 (N_2468,N_2395,N_2336);
or U2469 (N_2469,N_2348,N_2383);
and U2470 (N_2470,N_2346,N_2315);
and U2471 (N_2471,N_2385,N_2338);
and U2472 (N_2472,N_2397,N_2398);
nor U2473 (N_2473,N_2358,N_2399);
nand U2474 (N_2474,N_2342,N_2314);
and U2475 (N_2475,N_2311,N_2304);
and U2476 (N_2476,N_2364,N_2337);
nand U2477 (N_2477,N_2381,N_2307);
or U2478 (N_2478,N_2319,N_2350);
nor U2479 (N_2479,N_2357,N_2349);
and U2480 (N_2480,N_2312,N_2382);
nand U2481 (N_2481,N_2331,N_2340);
and U2482 (N_2482,N_2394,N_2327);
nand U2483 (N_2483,N_2363,N_2306);
nand U2484 (N_2484,N_2312,N_2316);
nor U2485 (N_2485,N_2388,N_2363);
nand U2486 (N_2486,N_2354,N_2367);
nor U2487 (N_2487,N_2354,N_2396);
nor U2488 (N_2488,N_2345,N_2393);
or U2489 (N_2489,N_2341,N_2392);
nand U2490 (N_2490,N_2387,N_2328);
nand U2491 (N_2491,N_2355,N_2377);
nand U2492 (N_2492,N_2306,N_2372);
and U2493 (N_2493,N_2380,N_2394);
or U2494 (N_2494,N_2354,N_2381);
nand U2495 (N_2495,N_2312,N_2321);
nor U2496 (N_2496,N_2362,N_2365);
or U2497 (N_2497,N_2349,N_2383);
or U2498 (N_2498,N_2392,N_2393);
and U2499 (N_2499,N_2371,N_2394);
nand U2500 (N_2500,N_2434,N_2456);
or U2501 (N_2501,N_2499,N_2483);
nand U2502 (N_2502,N_2481,N_2457);
nand U2503 (N_2503,N_2479,N_2448);
and U2504 (N_2504,N_2437,N_2424);
nor U2505 (N_2505,N_2484,N_2433);
nand U2506 (N_2506,N_2444,N_2445);
nand U2507 (N_2507,N_2401,N_2428);
nand U2508 (N_2508,N_2440,N_2490);
nor U2509 (N_2509,N_2454,N_2426);
and U2510 (N_2510,N_2447,N_2460);
and U2511 (N_2511,N_2459,N_2488);
nor U2512 (N_2512,N_2436,N_2404);
nand U2513 (N_2513,N_2475,N_2491);
nand U2514 (N_2514,N_2414,N_2458);
or U2515 (N_2515,N_2449,N_2411);
or U2516 (N_2516,N_2415,N_2430);
nand U2517 (N_2517,N_2425,N_2439);
and U2518 (N_2518,N_2492,N_2467);
or U2519 (N_2519,N_2464,N_2487);
or U2520 (N_2520,N_2423,N_2416);
or U2521 (N_2521,N_2453,N_2461);
nor U2522 (N_2522,N_2442,N_2493);
and U2523 (N_2523,N_2455,N_2400);
nand U2524 (N_2524,N_2462,N_2407);
or U2525 (N_2525,N_2443,N_2452);
and U2526 (N_2526,N_2473,N_2427);
nand U2527 (N_2527,N_2413,N_2405);
nor U2528 (N_2528,N_2470,N_2496);
nor U2529 (N_2529,N_2419,N_2476);
or U2530 (N_2530,N_2408,N_2450);
and U2531 (N_2531,N_2446,N_2463);
nor U2532 (N_2532,N_2410,N_2417);
and U2533 (N_2533,N_2497,N_2465);
nand U2534 (N_2534,N_2418,N_2466);
and U2535 (N_2535,N_2474,N_2486);
nand U2536 (N_2536,N_2409,N_2422);
nand U2537 (N_2537,N_2480,N_2435);
or U2538 (N_2538,N_2468,N_2498);
nand U2539 (N_2539,N_2403,N_2441);
nand U2540 (N_2540,N_2451,N_2438);
nor U2541 (N_2541,N_2489,N_2494);
or U2542 (N_2542,N_2431,N_2495);
nand U2543 (N_2543,N_2402,N_2469);
or U2544 (N_2544,N_2406,N_2420);
and U2545 (N_2545,N_2412,N_2485);
or U2546 (N_2546,N_2421,N_2477);
nand U2547 (N_2547,N_2432,N_2478);
nand U2548 (N_2548,N_2482,N_2472);
and U2549 (N_2549,N_2471,N_2429);
nor U2550 (N_2550,N_2405,N_2464);
and U2551 (N_2551,N_2449,N_2405);
nor U2552 (N_2552,N_2436,N_2483);
and U2553 (N_2553,N_2407,N_2419);
and U2554 (N_2554,N_2434,N_2475);
or U2555 (N_2555,N_2431,N_2407);
nand U2556 (N_2556,N_2438,N_2414);
nand U2557 (N_2557,N_2420,N_2475);
nor U2558 (N_2558,N_2449,N_2452);
or U2559 (N_2559,N_2418,N_2409);
nand U2560 (N_2560,N_2430,N_2422);
nand U2561 (N_2561,N_2420,N_2491);
and U2562 (N_2562,N_2491,N_2430);
or U2563 (N_2563,N_2413,N_2419);
or U2564 (N_2564,N_2480,N_2424);
nand U2565 (N_2565,N_2455,N_2495);
or U2566 (N_2566,N_2434,N_2416);
nand U2567 (N_2567,N_2453,N_2416);
nor U2568 (N_2568,N_2434,N_2446);
nand U2569 (N_2569,N_2489,N_2493);
nor U2570 (N_2570,N_2488,N_2472);
nand U2571 (N_2571,N_2489,N_2452);
nor U2572 (N_2572,N_2495,N_2458);
or U2573 (N_2573,N_2402,N_2434);
and U2574 (N_2574,N_2417,N_2426);
nor U2575 (N_2575,N_2414,N_2436);
nor U2576 (N_2576,N_2469,N_2484);
nand U2577 (N_2577,N_2428,N_2443);
nor U2578 (N_2578,N_2492,N_2493);
or U2579 (N_2579,N_2415,N_2492);
or U2580 (N_2580,N_2422,N_2487);
or U2581 (N_2581,N_2479,N_2449);
nor U2582 (N_2582,N_2483,N_2482);
nor U2583 (N_2583,N_2478,N_2457);
and U2584 (N_2584,N_2407,N_2487);
or U2585 (N_2585,N_2402,N_2447);
nor U2586 (N_2586,N_2435,N_2456);
nand U2587 (N_2587,N_2431,N_2415);
nand U2588 (N_2588,N_2488,N_2464);
nand U2589 (N_2589,N_2497,N_2426);
and U2590 (N_2590,N_2492,N_2442);
or U2591 (N_2591,N_2442,N_2432);
nor U2592 (N_2592,N_2412,N_2423);
or U2593 (N_2593,N_2474,N_2440);
and U2594 (N_2594,N_2448,N_2459);
and U2595 (N_2595,N_2470,N_2443);
nor U2596 (N_2596,N_2405,N_2459);
or U2597 (N_2597,N_2467,N_2453);
and U2598 (N_2598,N_2478,N_2485);
nand U2599 (N_2599,N_2457,N_2476);
and U2600 (N_2600,N_2527,N_2512);
and U2601 (N_2601,N_2506,N_2564);
nand U2602 (N_2602,N_2500,N_2559);
nand U2603 (N_2603,N_2502,N_2549);
nor U2604 (N_2604,N_2561,N_2528);
nand U2605 (N_2605,N_2551,N_2568);
nor U2606 (N_2606,N_2596,N_2597);
xor U2607 (N_2607,N_2553,N_2524);
and U2608 (N_2608,N_2554,N_2516);
and U2609 (N_2609,N_2592,N_2537);
or U2610 (N_2610,N_2504,N_2569);
nand U2611 (N_2611,N_2513,N_2519);
nor U2612 (N_2612,N_2534,N_2589);
and U2613 (N_2613,N_2582,N_2580);
nor U2614 (N_2614,N_2578,N_2546);
or U2615 (N_2615,N_2571,N_2508);
or U2616 (N_2616,N_2574,N_2501);
and U2617 (N_2617,N_2594,N_2584);
and U2618 (N_2618,N_2567,N_2581);
nand U2619 (N_2619,N_2510,N_2529);
or U2620 (N_2620,N_2585,N_2509);
nand U2621 (N_2621,N_2530,N_2507);
nand U2622 (N_2622,N_2517,N_2586);
nand U2623 (N_2623,N_2550,N_2598);
nor U2624 (N_2624,N_2560,N_2520);
or U2625 (N_2625,N_2541,N_2525);
and U2626 (N_2626,N_2576,N_2565);
or U2627 (N_2627,N_2536,N_2543);
nand U2628 (N_2628,N_2538,N_2505);
nand U2629 (N_2629,N_2523,N_2531);
nor U2630 (N_2630,N_2542,N_2590);
or U2631 (N_2631,N_2563,N_2547);
nor U2632 (N_2632,N_2599,N_2515);
and U2633 (N_2633,N_2514,N_2532);
nor U2634 (N_2634,N_2583,N_2539);
nor U2635 (N_2635,N_2573,N_2503);
nor U2636 (N_2636,N_2556,N_2518);
and U2637 (N_2637,N_2558,N_2579);
nor U2638 (N_2638,N_2557,N_2572);
nand U2639 (N_2639,N_2522,N_2545);
nor U2640 (N_2640,N_2575,N_2552);
nand U2641 (N_2641,N_2526,N_2593);
and U2642 (N_2642,N_2570,N_2562);
and U2643 (N_2643,N_2591,N_2533);
and U2644 (N_2644,N_2544,N_2535);
and U2645 (N_2645,N_2540,N_2577);
nor U2646 (N_2646,N_2566,N_2588);
or U2647 (N_2647,N_2511,N_2595);
nand U2648 (N_2648,N_2587,N_2555);
nand U2649 (N_2649,N_2521,N_2548);
and U2650 (N_2650,N_2540,N_2543);
and U2651 (N_2651,N_2527,N_2508);
nand U2652 (N_2652,N_2538,N_2522);
and U2653 (N_2653,N_2594,N_2551);
or U2654 (N_2654,N_2548,N_2584);
nor U2655 (N_2655,N_2551,N_2556);
nand U2656 (N_2656,N_2580,N_2567);
and U2657 (N_2657,N_2531,N_2576);
and U2658 (N_2658,N_2583,N_2587);
xnor U2659 (N_2659,N_2556,N_2541);
nor U2660 (N_2660,N_2523,N_2524);
and U2661 (N_2661,N_2571,N_2549);
nand U2662 (N_2662,N_2586,N_2569);
nor U2663 (N_2663,N_2553,N_2510);
nor U2664 (N_2664,N_2597,N_2521);
nand U2665 (N_2665,N_2599,N_2565);
nor U2666 (N_2666,N_2555,N_2595);
nor U2667 (N_2667,N_2561,N_2544);
nor U2668 (N_2668,N_2533,N_2518);
nand U2669 (N_2669,N_2559,N_2560);
and U2670 (N_2670,N_2559,N_2565);
nand U2671 (N_2671,N_2568,N_2513);
nand U2672 (N_2672,N_2558,N_2547);
or U2673 (N_2673,N_2580,N_2554);
and U2674 (N_2674,N_2582,N_2515);
and U2675 (N_2675,N_2522,N_2595);
nor U2676 (N_2676,N_2550,N_2585);
or U2677 (N_2677,N_2539,N_2518);
nor U2678 (N_2678,N_2567,N_2564);
and U2679 (N_2679,N_2548,N_2504);
or U2680 (N_2680,N_2507,N_2527);
and U2681 (N_2681,N_2562,N_2500);
nor U2682 (N_2682,N_2513,N_2582);
nor U2683 (N_2683,N_2567,N_2513);
nand U2684 (N_2684,N_2559,N_2593);
and U2685 (N_2685,N_2578,N_2593);
and U2686 (N_2686,N_2563,N_2574);
nand U2687 (N_2687,N_2571,N_2502);
nor U2688 (N_2688,N_2523,N_2552);
or U2689 (N_2689,N_2554,N_2523);
nand U2690 (N_2690,N_2539,N_2593);
nor U2691 (N_2691,N_2545,N_2542);
and U2692 (N_2692,N_2512,N_2509);
nor U2693 (N_2693,N_2548,N_2589);
or U2694 (N_2694,N_2532,N_2537);
nand U2695 (N_2695,N_2587,N_2505);
nor U2696 (N_2696,N_2585,N_2590);
nand U2697 (N_2697,N_2571,N_2538);
nand U2698 (N_2698,N_2566,N_2598);
and U2699 (N_2699,N_2500,N_2560);
nand U2700 (N_2700,N_2654,N_2682);
nand U2701 (N_2701,N_2648,N_2666);
nand U2702 (N_2702,N_2687,N_2698);
or U2703 (N_2703,N_2607,N_2623);
nand U2704 (N_2704,N_2678,N_2652);
nand U2705 (N_2705,N_2632,N_2617);
nor U2706 (N_2706,N_2657,N_2670);
nand U2707 (N_2707,N_2693,N_2661);
nand U2708 (N_2708,N_2667,N_2645);
and U2709 (N_2709,N_2639,N_2642);
nand U2710 (N_2710,N_2611,N_2691);
or U2711 (N_2711,N_2643,N_2695);
and U2712 (N_2712,N_2614,N_2647);
nor U2713 (N_2713,N_2694,N_2689);
nand U2714 (N_2714,N_2640,N_2636);
nand U2715 (N_2715,N_2658,N_2609);
nor U2716 (N_2716,N_2627,N_2608);
nand U2717 (N_2717,N_2618,N_2692);
nor U2718 (N_2718,N_2697,N_2602);
nand U2719 (N_2719,N_2651,N_2635);
or U2720 (N_2720,N_2662,N_2624);
or U2721 (N_2721,N_2673,N_2656);
and U2722 (N_2722,N_2610,N_2625);
nor U2723 (N_2723,N_2603,N_2660);
or U2724 (N_2724,N_2674,N_2630);
nand U2725 (N_2725,N_2615,N_2684);
nor U2726 (N_2726,N_2628,N_2650);
nand U2727 (N_2727,N_2629,N_2622);
and U2728 (N_2728,N_2637,N_2631);
nor U2729 (N_2729,N_2601,N_2675);
nand U2730 (N_2730,N_2620,N_2696);
nand U2731 (N_2731,N_2616,N_2664);
or U2732 (N_2732,N_2619,N_2672);
and U2733 (N_2733,N_2612,N_2613);
and U2734 (N_2734,N_2604,N_2683);
xor U2735 (N_2735,N_2600,N_2688);
xor U2736 (N_2736,N_2685,N_2641);
and U2737 (N_2737,N_2680,N_2638);
and U2738 (N_2738,N_2668,N_2679);
nor U2739 (N_2739,N_2659,N_2665);
and U2740 (N_2740,N_2644,N_2677);
nand U2741 (N_2741,N_2646,N_2626);
nor U2742 (N_2742,N_2621,N_2655);
or U2743 (N_2743,N_2634,N_2681);
nand U2744 (N_2744,N_2649,N_2690);
or U2745 (N_2745,N_2671,N_2606);
and U2746 (N_2746,N_2663,N_2669);
or U2747 (N_2747,N_2699,N_2633);
or U2748 (N_2748,N_2653,N_2676);
nand U2749 (N_2749,N_2605,N_2686);
nand U2750 (N_2750,N_2699,N_2669);
nand U2751 (N_2751,N_2622,N_2654);
nor U2752 (N_2752,N_2631,N_2647);
or U2753 (N_2753,N_2656,N_2639);
nand U2754 (N_2754,N_2637,N_2620);
nand U2755 (N_2755,N_2681,N_2607);
or U2756 (N_2756,N_2622,N_2684);
nand U2757 (N_2757,N_2657,N_2698);
nand U2758 (N_2758,N_2623,N_2660);
nand U2759 (N_2759,N_2677,N_2613);
and U2760 (N_2760,N_2644,N_2659);
or U2761 (N_2761,N_2649,N_2672);
and U2762 (N_2762,N_2674,N_2671);
nand U2763 (N_2763,N_2648,N_2626);
nor U2764 (N_2764,N_2683,N_2622);
nor U2765 (N_2765,N_2678,N_2624);
nor U2766 (N_2766,N_2622,N_2606);
nand U2767 (N_2767,N_2629,N_2618);
nand U2768 (N_2768,N_2642,N_2666);
nor U2769 (N_2769,N_2615,N_2600);
and U2770 (N_2770,N_2641,N_2617);
nor U2771 (N_2771,N_2630,N_2656);
nand U2772 (N_2772,N_2642,N_2623);
nor U2773 (N_2773,N_2602,N_2689);
or U2774 (N_2774,N_2610,N_2636);
or U2775 (N_2775,N_2656,N_2668);
nor U2776 (N_2776,N_2677,N_2686);
nand U2777 (N_2777,N_2656,N_2615);
and U2778 (N_2778,N_2688,N_2670);
nand U2779 (N_2779,N_2626,N_2633);
nand U2780 (N_2780,N_2624,N_2671);
nor U2781 (N_2781,N_2642,N_2655);
or U2782 (N_2782,N_2673,N_2616);
and U2783 (N_2783,N_2674,N_2677);
and U2784 (N_2784,N_2651,N_2665);
and U2785 (N_2785,N_2629,N_2699);
and U2786 (N_2786,N_2693,N_2683);
or U2787 (N_2787,N_2604,N_2606);
and U2788 (N_2788,N_2640,N_2675);
and U2789 (N_2789,N_2675,N_2670);
nand U2790 (N_2790,N_2668,N_2698);
or U2791 (N_2791,N_2603,N_2664);
or U2792 (N_2792,N_2673,N_2697);
nand U2793 (N_2793,N_2695,N_2690);
and U2794 (N_2794,N_2673,N_2611);
or U2795 (N_2795,N_2613,N_2673);
nor U2796 (N_2796,N_2626,N_2649);
nand U2797 (N_2797,N_2620,N_2683);
or U2798 (N_2798,N_2644,N_2650);
or U2799 (N_2799,N_2638,N_2655);
nor U2800 (N_2800,N_2793,N_2752);
and U2801 (N_2801,N_2797,N_2743);
nor U2802 (N_2802,N_2778,N_2726);
nor U2803 (N_2803,N_2741,N_2774);
and U2804 (N_2804,N_2708,N_2776);
nand U2805 (N_2805,N_2719,N_2715);
nand U2806 (N_2806,N_2710,N_2749);
nor U2807 (N_2807,N_2730,N_2733);
nor U2808 (N_2808,N_2707,N_2788);
nand U2809 (N_2809,N_2772,N_2702);
or U2810 (N_2810,N_2756,N_2761);
nand U2811 (N_2811,N_2735,N_2742);
nor U2812 (N_2812,N_2728,N_2732);
nor U2813 (N_2813,N_2706,N_2718);
nand U2814 (N_2814,N_2757,N_2763);
or U2815 (N_2815,N_2747,N_2760);
nand U2816 (N_2816,N_2783,N_2789);
or U2817 (N_2817,N_2736,N_2767);
or U2818 (N_2818,N_2745,N_2751);
nand U2819 (N_2819,N_2777,N_2794);
and U2820 (N_2820,N_2795,N_2725);
or U2821 (N_2821,N_2711,N_2770);
and U2822 (N_2822,N_2705,N_2786);
and U2823 (N_2823,N_2787,N_2720);
nor U2824 (N_2824,N_2768,N_2721);
nor U2825 (N_2825,N_2799,N_2779);
nand U2826 (N_2826,N_2701,N_2773);
nand U2827 (N_2827,N_2754,N_2714);
nor U2828 (N_2828,N_2782,N_2722);
nor U2829 (N_2829,N_2729,N_2798);
nor U2830 (N_2830,N_2791,N_2759);
nand U2831 (N_2831,N_2723,N_2764);
nand U2832 (N_2832,N_2734,N_2731);
or U2833 (N_2833,N_2785,N_2771);
nand U2834 (N_2834,N_2712,N_2703);
nand U2835 (N_2835,N_2704,N_2713);
nand U2836 (N_2836,N_2746,N_2758);
nand U2837 (N_2837,N_2790,N_2700);
nand U2838 (N_2838,N_2781,N_2744);
or U2839 (N_2839,N_2762,N_2755);
nor U2840 (N_2840,N_2769,N_2753);
and U2841 (N_2841,N_2737,N_2766);
nor U2842 (N_2842,N_2724,N_2709);
or U2843 (N_2843,N_2717,N_2796);
and U2844 (N_2844,N_2716,N_2738);
or U2845 (N_2845,N_2740,N_2775);
nor U2846 (N_2846,N_2780,N_2784);
or U2847 (N_2847,N_2765,N_2748);
and U2848 (N_2848,N_2739,N_2727);
nor U2849 (N_2849,N_2792,N_2750);
nor U2850 (N_2850,N_2739,N_2784);
xnor U2851 (N_2851,N_2785,N_2746);
or U2852 (N_2852,N_2738,N_2759);
nand U2853 (N_2853,N_2718,N_2747);
or U2854 (N_2854,N_2737,N_2745);
or U2855 (N_2855,N_2769,N_2750);
or U2856 (N_2856,N_2741,N_2746);
nand U2857 (N_2857,N_2763,N_2775);
nor U2858 (N_2858,N_2703,N_2791);
nand U2859 (N_2859,N_2793,N_2745);
nand U2860 (N_2860,N_2772,N_2746);
nor U2861 (N_2861,N_2700,N_2708);
and U2862 (N_2862,N_2714,N_2706);
or U2863 (N_2863,N_2733,N_2755);
nor U2864 (N_2864,N_2797,N_2705);
nand U2865 (N_2865,N_2792,N_2783);
or U2866 (N_2866,N_2717,N_2775);
or U2867 (N_2867,N_2777,N_2786);
or U2868 (N_2868,N_2718,N_2703);
and U2869 (N_2869,N_2745,N_2775);
nand U2870 (N_2870,N_2798,N_2740);
or U2871 (N_2871,N_2788,N_2708);
nand U2872 (N_2872,N_2781,N_2743);
and U2873 (N_2873,N_2717,N_2720);
or U2874 (N_2874,N_2789,N_2721);
xor U2875 (N_2875,N_2768,N_2782);
nor U2876 (N_2876,N_2725,N_2700);
nor U2877 (N_2877,N_2714,N_2799);
and U2878 (N_2878,N_2709,N_2748);
and U2879 (N_2879,N_2783,N_2758);
or U2880 (N_2880,N_2799,N_2793);
or U2881 (N_2881,N_2719,N_2767);
nand U2882 (N_2882,N_2701,N_2726);
or U2883 (N_2883,N_2770,N_2737);
and U2884 (N_2884,N_2738,N_2776);
or U2885 (N_2885,N_2759,N_2796);
nand U2886 (N_2886,N_2720,N_2723);
or U2887 (N_2887,N_2718,N_2752);
and U2888 (N_2888,N_2756,N_2709);
nand U2889 (N_2889,N_2717,N_2779);
or U2890 (N_2890,N_2791,N_2735);
and U2891 (N_2891,N_2786,N_2729);
and U2892 (N_2892,N_2752,N_2712);
or U2893 (N_2893,N_2734,N_2713);
or U2894 (N_2894,N_2781,N_2786);
and U2895 (N_2895,N_2770,N_2757);
or U2896 (N_2896,N_2732,N_2755);
or U2897 (N_2897,N_2782,N_2728);
or U2898 (N_2898,N_2754,N_2763);
or U2899 (N_2899,N_2755,N_2731);
and U2900 (N_2900,N_2892,N_2816);
nand U2901 (N_2901,N_2831,N_2832);
nand U2902 (N_2902,N_2894,N_2882);
or U2903 (N_2903,N_2873,N_2859);
nor U2904 (N_2904,N_2839,N_2880);
and U2905 (N_2905,N_2808,N_2818);
or U2906 (N_2906,N_2837,N_2847);
and U2907 (N_2907,N_2820,N_2819);
nand U2908 (N_2908,N_2891,N_2851);
nor U2909 (N_2909,N_2821,N_2840);
or U2910 (N_2910,N_2805,N_2849);
nor U2911 (N_2911,N_2872,N_2812);
nand U2912 (N_2912,N_2807,N_2815);
or U2913 (N_2913,N_2874,N_2867);
or U2914 (N_2914,N_2826,N_2877);
nor U2915 (N_2915,N_2884,N_2813);
nand U2916 (N_2916,N_2887,N_2801);
nand U2917 (N_2917,N_2865,N_2822);
nor U2918 (N_2918,N_2848,N_2855);
or U2919 (N_2919,N_2829,N_2869);
nand U2920 (N_2920,N_2883,N_2856);
or U2921 (N_2921,N_2852,N_2889);
nand U2922 (N_2922,N_2863,N_2836);
or U2923 (N_2923,N_2841,N_2828);
nor U2924 (N_2924,N_2834,N_2838);
and U2925 (N_2925,N_2800,N_2854);
nand U2926 (N_2926,N_2817,N_2864);
and U2927 (N_2927,N_2876,N_2897);
and U2928 (N_2928,N_2844,N_2850);
nand U2929 (N_2929,N_2846,N_2888);
or U2930 (N_2930,N_2862,N_2833);
nor U2931 (N_2931,N_2806,N_2825);
nand U2932 (N_2932,N_2893,N_2830);
nor U2933 (N_2933,N_2881,N_2811);
or U2934 (N_2934,N_2875,N_2853);
nand U2935 (N_2935,N_2827,N_2809);
nand U2936 (N_2936,N_2823,N_2890);
or U2937 (N_2937,N_2858,N_2871);
nand U2938 (N_2938,N_2899,N_2860);
nor U2939 (N_2939,N_2861,N_2885);
or U2940 (N_2940,N_2898,N_2866);
or U2941 (N_2941,N_2879,N_2810);
and U2942 (N_2942,N_2896,N_2814);
and U2943 (N_2943,N_2868,N_2895);
nor U2944 (N_2944,N_2878,N_2843);
nor U2945 (N_2945,N_2804,N_2824);
nand U2946 (N_2946,N_2842,N_2835);
and U2947 (N_2947,N_2802,N_2886);
and U2948 (N_2948,N_2857,N_2803);
nor U2949 (N_2949,N_2845,N_2870);
or U2950 (N_2950,N_2886,N_2806);
nor U2951 (N_2951,N_2846,N_2886);
or U2952 (N_2952,N_2814,N_2810);
or U2953 (N_2953,N_2837,N_2870);
and U2954 (N_2954,N_2825,N_2841);
nand U2955 (N_2955,N_2885,N_2873);
or U2956 (N_2956,N_2801,N_2895);
nand U2957 (N_2957,N_2873,N_2850);
or U2958 (N_2958,N_2835,N_2858);
nand U2959 (N_2959,N_2862,N_2873);
and U2960 (N_2960,N_2895,N_2835);
and U2961 (N_2961,N_2864,N_2837);
and U2962 (N_2962,N_2854,N_2820);
and U2963 (N_2963,N_2849,N_2847);
nor U2964 (N_2964,N_2832,N_2804);
nor U2965 (N_2965,N_2866,N_2807);
nand U2966 (N_2966,N_2827,N_2896);
nor U2967 (N_2967,N_2800,N_2823);
nand U2968 (N_2968,N_2850,N_2872);
or U2969 (N_2969,N_2811,N_2894);
nor U2970 (N_2970,N_2896,N_2860);
nor U2971 (N_2971,N_2823,N_2888);
nor U2972 (N_2972,N_2862,N_2867);
or U2973 (N_2973,N_2813,N_2815);
or U2974 (N_2974,N_2850,N_2852);
and U2975 (N_2975,N_2867,N_2871);
or U2976 (N_2976,N_2811,N_2897);
nor U2977 (N_2977,N_2802,N_2851);
or U2978 (N_2978,N_2875,N_2829);
nand U2979 (N_2979,N_2879,N_2833);
nor U2980 (N_2980,N_2879,N_2897);
nor U2981 (N_2981,N_2837,N_2874);
xor U2982 (N_2982,N_2838,N_2864);
or U2983 (N_2983,N_2809,N_2826);
nand U2984 (N_2984,N_2817,N_2872);
nand U2985 (N_2985,N_2895,N_2855);
nand U2986 (N_2986,N_2862,N_2876);
xnor U2987 (N_2987,N_2850,N_2858);
and U2988 (N_2988,N_2876,N_2853);
or U2989 (N_2989,N_2883,N_2848);
or U2990 (N_2990,N_2813,N_2863);
or U2991 (N_2991,N_2883,N_2867);
and U2992 (N_2992,N_2840,N_2834);
or U2993 (N_2993,N_2829,N_2817);
nor U2994 (N_2994,N_2888,N_2838);
or U2995 (N_2995,N_2867,N_2878);
nand U2996 (N_2996,N_2876,N_2867);
or U2997 (N_2997,N_2899,N_2877);
nand U2998 (N_2998,N_2896,N_2813);
or U2999 (N_2999,N_2839,N_2829);
xor UO_0 (O_0,N_2908,N_2902);
nor UO_1 (O_1,N_2905,N_2964);
or UO_2 (O_2,N_2984,N_2990);
nor UO_3 (O_3,N_2942,N_2943);
or UO_4 (O_4,N_2903,N_2963);
or UO_5 (O_5,N_2931,N_2989);
and UO_6 (O_6,N_2945,N_2976);
and UO_7 (O_7,N_2944,N_2995);
or UO_8 (O_8,N_2971,N_2993);
nor UO_9 (O_9,N_2994,N_2983);
nor UO_10 (O_10,N_2914,N_2978);
and UO_11 (O_11,N_2939,N_2965);
or UO_12 (O_12,N_2958,N_2987);
and UO_13 (O_13,N_2952,N_2909);
nor UO_14 (O_14,N_2949,N_2985);
nand UO_15 (O_15,N_2925,N_2938);
nor UO_16 (O_16,N_2954,N_2979);
nand UO_17 (O_17,N_2906,N_2972);
nor UO_18 (O_18,N_2946,N_2910);
nor UO_19 (O_19,N_2973,N_2920);
nand UO_20 (O_20,N_2966,N_2999);
nand UO_21 (O_21,N_2975,N_2998);
or UO_22 (O_22,N_2967,N_2934);
nand UO_23 (O_23,N_2923,N_2961);
nand UO_24 (O_24,N_2922,N_2913);
nor UO_25 (O_25,N_2981,N_2941);
xnor UO_26 (O_26,N_2997,N_2916);
and UO_27 (O_27,N_2900,N_2960);
nand UO_28 (O_28,N_2927,N_2912);
and UO_29 (O_29,N_2926,N_2936);
and UO_30 (O_30,N_2951,N_2940);
or UO_31 (O_31,N_2955,N_2924);
nand UO_32 (O_32,N_2911,N_2935);
nand UO_33 (O_33,N_2947,N_2930);
and UO_34 (O_34,N_2921,N_2980);
nand UO_35 (O_35,N_2950,N_2928);
nor UO_36 (O_36,N_2933,N_2974);
nand UO_37 (O_37,N_2957,N_2996);
nor UO_38 (O_38,N_2915,N_2988);
nor UO_39 (O_39,N_2982,N_2956);
and UO_40 (O_40,N_2953,N_2904);
nor UO_41 (O_41,N_2901,N_2919);
nand UO_42 (O_42,N_2932,N_2918);
and UO_43 (O_43,N_2969,N_2991);
or UO_44 (O_44,N_2937,N_2959);
nand UO_45 (O_45,N_2962,N_2929);
nand UO_46 (O_46,N_2986,N_2977);
nand UO_47 (O_47,N_2968,N_2970);
and UO_48 (O_48,N_2917,N_2992);
nand UO_49 (O_49,N_2948,N_2907);
and UO_50 (O_50,N_2995,N_2998);
nor UO_51 (O_51,N_2900,N_2969);
or UO_52 (O_52,N_2965,N_2900);
nor UO_53 (O_53,N_2974,N_2928);
nand UO_54 (O_54,N_2931,N_2905);
or UO_55 (O_55,N_2928,N_2972);
nor UO_56 (O_56,N_2981,N_2966);
and UO_57 (O_57,N_2989,N_2982);
nor UO_58 (O_58,N_2916,N_2915);
or UO_59 (O_59,N_2944,N_2943);
and UO_60 (O_60,N_2952,N_2935);
nor UO_61 (O_61,N_2996,N_2982);
nor UO_62 (O_62,N_2918,N_2913);
and UO_63 (O_63,N_2973,N_2915);
nor UO_64 (O_64,N_2935,N_2905);
nand UO_65 (O_65,N_2981,N_2984);
nor UO_66 (O_66,N_2976,N_2963);
nand UO_67 (O_67,N_2962,N_2948);
nor UO_68 (O_68,N_2997,N_2967);
nor UO_69 (O_69,N_2983,N_2946);
nand UO_70 (O_70,N_2975,N_2919);
or UO_71 (O_71,N_2984,N_2907);
and UO_72 (O_72,N_2992,N_2957);
nand UO_73 (O_73,N_2925,N_2931);
nand UO_74 (O_74,N_2928,N_2907);
or UO_75 (O_75,N_2991,N_2965);
and UO_76 (O_76,N_2917,N_2951);
and UO_77 (O_77,N_2989,N_2925);
or UO_78 (O_78,N_2922,N_2932);
or UO_79 (O_79,N_2940,N_2999);
nor UO_80 (O_80,N_2974,N_2941);
xor UO_81 (O_81,N_2961,N_2940);
or UO_82 (O_82,N_2942,N_2981);
nand UO_83 (O_83,N_2911,N_2970);
or UO_84 (O_84,N_2923,N_2909);
or UO_85 (O_85,N_2955,N_2988);
nor UO_86 (O_86,N_2920,N_2957);
nand UO_87 (O_87,N_2972,N_2913);
nand UO_88 (O_88,N_2974,N_2980);
or UO_89 (O_89,N_2989,N_2904);
or UO_90 (O_90,N_2943,N_2962);
nand UO_91 (O_91,N_2996,N_2983);
nor UO_92 (O_92,N_2996,N_2988);
nand UO_93 (O_93,N_2931,N_2949);
or UO_94 (O_94,N_2954,N_2974);
nand UO_95 (O_95,N_2959,N_2995);
nor UO_96 (O_96,N_2938,N_2927);
nor UO_97 (O_97,N_2999,N_2955);
or UO_98 (O_98,N_2969,N_2920);
nor UO_99 (O_99,N_2955,N_2990);
nand UO_100 (O_100,N_2970,N_2944);
or UO_101 (O_101,N_2997,N_2904);
nor UO_102 (O_102,N_2908,N_2925);
nor UO_103 (O_103,N_2904,N_2937);
or UO_104 (O_104,N_2920,N_2994);
and UO_105 (O_105,N_2961,N_2920);
or UO_106 (O_106,N_2959,N_2981);
or UO_107 (O_107,N_2944,N_2954);
or UO_108 (O_108,N_2959,N_2965);
nor UO_109 (O_109,N_2913,N_2925);
nand UO_110 (O_110,N_2966,N_2954);
and UO_111 (O_111,N_2959,N_2904);
or UO_112 (O_112,N_2965,N_2969);
or UO_113 (O_113,N_2922,N_2949);
nor UO_114 (O_114,N_2961,N_2933);
or UO_115 (O_115,N_2932,N_2906);
nand UO_116 (O_116,N_2980,N_2986);
nor UO_117 (O_117,N_2940,N_2930);
nor UO_118 (O_118,N_2992,N_2935);
and UO_119 (O_119,N_2960,N_2927);
nor UO_120 (O_120,N_2997,N_2924);
and UO_121 (O_121,N_2919,N_2932);
nand UO_122 (O_122,N_2999,N_2989);
nor UO_123 (O_123,N_2970,N_2926);
or UO_124 (O_124,N_2924,N_2952);
nor UO_125 (O_125,N_2997,N_2927);
nor UO_126 (O_126,N_2970,N_2918);
nand UO_127 (O_127,N_2911,N_2920);
nand UO_128 (O_128,N_2932,N_2946);
or UO_129 (O_129,N_2903,N_2911);
nor UO_130 (O_130,N_2924,N_2932);
nand UO_131 (O_131,N_2971,N_2982);
and UO_132 (O_132,N_2972,N_2994);
and UO_133 (O_133,N_2989,N_2976);
nor UO_134 (O_134,N_2912,N_2996);
nand UO_135 (O_135,N_2911,N_2905);
nor UO_136 (O_136,N_2917,N_2949);
nand UO_137 (O_137,N_2985,N_2991);
and UO_138 (O_138,N_2955,N_2984);
and UO_139 (O_139,N_2914,N_2933);
and UO_140 (O_140,N_2931,N_2933);
nor UO_141 (O_141,N_2934,N_2937);
and UO_142 (O_142,N_2961,N_2934);
nor UO_143 (O_143,N_2991,N_2937);
or UO_144 (O_144,N_2935,N_2900);
nor UO_145 (O_145,N_2933,N_2919);
nor UO_146 (O_146,N_2914,N_2902);
and UO_147 (O_147,N_2976,N_2969);
or UO_148 (O_148,N_2953,N_2925);
nor UO_149 (O_149,N_2914,N_2999);
nand UO_150 (O_150,N_2952,N_2933);
nor UO_151 (O_151,N_2933,N_2999);
and UO_152 (O_152,N_2932,N_2991);
xor UO_153 (O_153,N_2946,N_2995);
nor UO_154 (O_154,N_2983,N_2932);
and UO_155 (O_155,N_2905,N_2959);
nand UO_156 (O_156,N_2941,N_2979);
and UO_157 (O_157,N_2973,N_2956);
nor UO_158 (O_158,N_2966,N_2903);
or UO_159 (O_159,N_2942,N_2911);
nand UO_160 (O_160,N_2963,N_2937);
and UO_161 (O_161,N_2989,N_2997);
and UO_162 (O_162,N_2990,N_2940);
nor UO_163 (O_163,N_2951,N_2985);
nor UO_164 (O_164,N_2904,N_2995);
nor UO_165 (O_165,N_2938,N_2961);
or UO_166 (O_166,N_2971,N_2936);
and UO_167 (O_167,N_2961,N_2951);
nor UO_168 (O_168,N_2988,N_2971);
nor UO_169 (O_169,N_2955,N_2920);
and UO_170 (O_170,N_2921,N_2968);
nor UO_171 (O_171,N_2958,N_2911);
nor UO_172 (O_172,N_2908,N_2906);
nor UO_173 (O_173,N_2901,N_2968);
and UO_174 (O_174,N_2999,N_2990);
nor UO_175 (O_175,N_2944,N_2934);
or UO_176 (O_176,N_2952,N_2981);
and UO_177 (O_177,N_2917,N_2976);
and UO_178 (O_178,N_2985,N_2953);
nor UO_179 (O_179,N_2975,N_2973);
or UO_180 (O_180,N_2978,N_2944);
or UO_181 (O_181,N_2945,N_2911);
and UO_182 (O_182,N_2919,N_2929);
nor UO_183 (O_183,N_2988,N_2967);
or UO_184 (O_184,N_2901,N_2911);
or UO_185 (O_185,N_2916,N_2952);
nor UO_186 (O_186,N_2924,N_2971);
or UO_187 (O_187,N_2953,N_2971);
nand UO_188 (O_188,N_2959,N_2935);
or UO_189 (O_189,N_2988,N_2953);
and UO_190 (O_190,N_2993,N_2934);
nor UO_191 (O_191,N_2972,N_2963);
xor UO_192 (O_192,N_2913,N_2943);
nor UO_193 (O_193,N_2976,N_2985);
nand UO_194 (O_194,N_2942,N_2936);
nand UO_195 (O_195,N_2941,N_2945);
or UO_196 (O_196,N_2911,N_2977);
and UO_197 (O_197,N_2972,N_2902);
or UO_198 (O_198,N_2969,N_2997);
and UO_199 (O_199,N_2928,N_2993);
nor UO_200 (O_200,N_2984,N_2961);
nor UO_201 (O_201,N_2915,N_2942);
or UO_202 (O_202,N_2979,N_2902);
nand UO_203 (O_203,N_2996,N_2961);
or UO_204 (O_204,N_2988,N_2907);
nor UO_205 (O_205,N_2991,N_2971);
nand UO_206 (O_206,N_2960,N_2999);
or UO_207 (O_207,N_2928,N_2992);
nand UO_208 (O_208,N_2940,N_2959);
nor UO_209 (O_209,N_2993,N_2965);
and UO_210 (O_210,N_2943,N_2979);
nor UO_211 (O_211,N_2953,N_2926);
and UO_212 (O_212,N_2925,N_2962);
nor UO_213 (O_213,N_2913,N_2966);
and UO_214 (O_214,N_2975,N_2920);
nand UO_215 (O_215,N_2907,N_2911);
nor UO_216 (O_216,N_2976,N_2998);
nor UO_217 (O_217,N_2916,N_2901);
and UO_218 (O_218,N_2991,N_2931);
or UO_219 (O_219,N_2980,N_2945);
nor UO_220 (O_220,N_2982,N_2901);
nand UO_221 (O_221,N_2987,N_2934);
nand UO_222 (O_222,N_2948,N_2922);
nor UO_223 (O_223,N_2987,N_2984);
or UO_224 (O_224,N_2960,N_2946);
and UO_225 (O_225,N_2953,N_2932);
nand UO_226 (O_226,N_2994,N_2924);
or UO_227 (O_227,N_2917,N_2922);
nor UO_228 (O_228,N_2960,N_2975);
nand UO_229 (O_229,N_2937,N_2994);
nand UO_230 (O_230,N_2908,N_2904);
and UO_231 (O_231,N_2923,N_2994);
and UO_232 (O_232,N_2905,N_2948);
and UO_233 (O_233,N_2977,N_2912);
or UO_234 (O_234,N_2916,N_2904);
nand UO_235 (O_235,N_2934,N_2999);
and UO_236 (O_236,N_2971,N_2949);
nand UO_237 (O_237,N_2962,N_2923);
nand UO_238 (O_238,N_2905,N_2924);
nor UO_239 (O_239,N_2999,N_2924);
and UO_240 (O_240,N_2925,N_2923);
or UO_241 (O_241,N_2919,N_2985);
nor UO_242 (O_242,N_2996,N_2987);
or UO_243 (O_243,N_2981,N_2924);
xnor UO_244 (O_244,N_2958,N_2997);
and UO_245 (O_245,N_2930,N_2917);
and UO_246 (O_246,N_2951,N_2991);
nand UO_247 (O_247,N_2929,N_2926);
nor UO_248 (O_248,N_2906,N_2921);
nand UO_249 (O_249,N_2939,N_2994);
nor UO_250 (O_250,N_2905,N_2926);
nand UO_251 (O_251,N_2929,N_2995);
nor UO_252 (O_252,N_2931,N_2979);
and UO_253 (O_253,N_2925,N_2993);
and UO_254 (O_254,N_2993,N_2997);
nor UO_255 (O_255,N_2954,N_2968);
nand UO_256 (O_256,N_2950,N_2962);
nand UO_257 (O_257,N_2990,N_2909);
or UO_258 (O_258,N_2928,N_2906);
nor UO_259 (O_259,N_2909,N_2920);
or UO_260 (O_260,N_2954,N_2975);
nand UO_261 (O_261,N_2977,N_2961);
and UO_262 (O_262,N_2964,N_2997);
and UO_263 (O_263,N_2995,N_2917);
nor UO_264 (O_264,N_2913,N_2921);
nor UO_265 (O_265,N_2992,N_2943);
and UO_266 (O_266,N_2923,N_2944);
nand UO_267 (O_267,N_2982,N_2949);
and UO_268 (O_268,N_2903,N_2940);
or UO_269 (O_269,N_2904,N_2913);
nand UO_270 (O_270,N_2976,N_2911);
and UO_271 (O_271,N_2904,N_2944);
and UO_272 (O_272,N_2994,N_2948);
nor UO_273 (O_273,N_2939,N_2919);
or UO_274 (O_274,N_2960,N_2950);
nor UO_275 (O_275,N_2973,N_2930);
nor UO_276 (O_276,N_2931,N_2938);
and UO_277 (O_277,N_2935,N_2903);
or UO_278 (O_278,N_2953,N_2978);
nand UO_279 (O_279,N_2983,N_2944);
or UO_280 (O_280,N_2929,N_2939);
nand UO_281 (O_281,N_2907,N_2906);
nor UO_282 (O_282,N_2904,N_2960);
nand UO_283 (O_283,N_2948,N_2959);
nand UO_284 (O_284,N_2935,N_2977);
and UO_285 (O_285,N_2951,N_2987);
or UO_286 (O_286,N_2907,N_2920);
or UO_287 (O_287,N_2947,N_2906);
nand UO_288 (O_288,N_2917,N_2936);
and UO_289 (O_289,N_2979,N_2990);
or UO_290 (O_290,N_2943,N_2981);
and UO_291 (O_291,N_2943,N_2959);
or UO_292 (O_292,N_2953,N_2962);
or UO_293 (O_293,N_2993,N_2982);
or UO_294 (O_294,N_2934,N_2928);
nor UO_295 (O_295,N_2994,N_2916);
nand UO_296 (O_296,N_2948,N_2915);
and UO_297 (O_297,N_2981,N_2988);
and UO_298 (O_298,N_2900,N_2921);
and UO_299 (O_299,N_2961,N_2909);
nand UO_300 (O_300,N_2901,N_2934);
and UO_301 (O_301,N_2977,N_2950);
or UO_302 (O_302,N_2974,N_2917);
or UO_303 (O_303,N_2913,N_2998);
or UO_304 (O_304,N_2924,N_2980);
or UO_305 (O_305,N_2968,N_2992);
nor UO_306 (O_306,N_2956,N_2924);
nand UO_307 (O_307,N_2974,N_2949);
and UO_308 (O_308,N_2985,N_2911);
and UO_309 (O_309,N_2996,N_2969);
and UO_310 (O_310,N_2933,N_2994);
nand UO_311 (O_311,N_2968,N_2965);
nor UO_312 (O_312,N_2966,N_2996);
nor UO_313 (O_313,N_2986,N_2994);
nor UO_314 (O_314,N_2900,N_2949);
xor UO_315 (O_315,N_2999,N_2993);
nand UO_316 (O_316,N_2953,N_2996);
and UO_317 (O_317,N_2906,N_2978);
nand UO_318 (O_318,N_2967,N_2912);
xor UO_319 (O_319,N_2952,N_2960);
or UO_320 (O_320,N_2952,N_2915);
nand UO_321 (O_321,N_2903,N_2930);
nand UO_322 (O_322,N_2935,N_2919);
and UO_323 (O_323,N_2997,N_2945);
and UO_324 (O_324,N_2961,N_2987);
nor UO_325 (O_325,N_2902,N_2982);
and UO_326 (O_326,N_2965,N_2997);
nand UO_327 (O_327,N_2916,N_2978);
and UO_328 (O_328,N_2956,N_2905);
nand UO_329 (O_329,N_2925,N_2972);
nand UO_330 (O_330,N_2951,N_2910);
nand UO_331 (O_331,N_2982,N_2938);
and UO_332 (O_332,N_2975,N_2963);
and UO_333 (O_333,N_2999,N_2982);
nor UO_334 (O_334,N_2926,N_2935);
nand UO_335 (O_335,N_2942,N_2956);
nand UO_336 (O_336,N_2957,N_2926);
and UO_337 (O_337,N_2933,N_2993);
and UO_338 (O_338,N_2927,N_2972);
and UO_339 (O_339,N_2909,N_2949);
or UO_340 (O_340,N_2932,N_2956);
nand UO_341 (O_341,N_2997,N_2962);
nor UO_342 (O_342,N_2950,N_2927);
and UO_343 (O_343,N_2967,N_2926);
or UO_344 (O_344,N_2923,N_2903);
or UO_345 (O_345,N_2917,N_2980);
xor UO_346 (O_346,N_2909,N_2951);
or UO_347 (O_347,N_2925,N_2917);
nand UO_348 (O_348,N_2993,N_2969);
nand UO_349 (O_349,N_2924,N_2930);
nand UO_350 (O_350,N_2960,N_2986);
nor UO_351 (O_351,N_2902,N_2904);
or UO_352 (O_352,N_2936,N_2910);
or UO_353 (O_353,N_2943,N_2941);
nand UO_354 (O_354,N_2929,N_2941);
nor UO_355 (O_355,N_2979,N_2978);
or UO_356 (O_356,N_2940,N_2955);
nor UO_357 (O_357,N_2986,N_2911);
nor UO_358 (O_358,N_2938,N_2901);
nor UO_359 (O_359,N_2973,N_2903);
nor UO_360 (O_360,N_2982,N_2917);
nand UO_361 (O_361,N_2925,N_2994);
and UO_362 (O_362,N_2960,N_2984);
and UO_363 (O_363,N_2943,N_2924);
and UO_364 (O_364,N_2951,N_2964);
and UO_365 (O_365,N_2960,N_2979);
nor UO_366 (O_366,N_2940,N_2965);
or UO_367 (O_367,N_2961,N_2954);
and UO_368 (O_368,N_2936,N_2920);
and UO_369 (O_369,N_2988,N_2980);
nand UO_370 (O_370,N_2977,N_2963);
and UO_371 (O_371,N_2929,N_2983);
or UO_372 (O_372,N_2985,N_2926);
or UO_373 (O_373,N_2934,N_2977);
nor UO_374 (O_374,N_2995,N_2903);
or UO_375 (O_375,N_2937,N_2961);
nor UO_376 (O_376,N_2971,N_2954);
and UO_377 (O_377,N_2929,N_2932);
nand UO_378 (O_378,N_2992,N_2937);
nor UO_379 (O_379,N_2975,N_2964);
nand UO_380 (O_380,N_2961,N_2990);
or UO_381 (O_381,N_2995,N_2987);
or UO_382 (O_382,N_2908,N_2982);
or UO_383 (O_383,N_2922,N_2963);
nand UO_384 (O_384,N_2910,N_2918);
nand UO_385 (O_385,N_2933,N_2934);
or UO_386 (O_386,N_2910,N_2915);
nor UO_387 (O_387,N_2963,N_2984);
and UO_388 (O_388,N_2933,N_2922);
and UO_389 (O_389,N_2970,N_2981);
or UO_390 (O_390,N_2957,N_2950);
nor UO_391 (O_391,N_2932,N_2990);
and UO_392 (O_392,N_2960,N_2976);
and UO_393 (O_393,N_2905,N_2977);
or UO_394 (O_394,N_2988,N_2940);
and UO_395 (O_395,N_2936,N_2998);
nand UO_396 (O_396,N_2989,N_2986);
or UO_397 (O_397,N_2993,N_2970);
and UO_398 (O_398,N_2939,N_2963);
or UO_399 (O_399,N_2936,N_2986);
nand UO_400 (O_400,N_2909,N_2947);
nor UO_401 (O_401,N_2940,N_2915);
and UO_402 (O_402,N_2933,N_2970);
nor UO_403 (O_403,N_2999,N_2931);
nand UO_404 (O_404,N_2949,N_2943);
and UO_405 (O_405,N_2933,N_2966);
and UO_406 (O_406,N_2902,N_2901);
or UO_407 (O_407,N_2986,N_2914);
nand UO_408 (O_408,N_2931,N_2959);
and UO_409 (O_409,N_2995,N_2916);
and UO_410 (O_410,N_2992,N_2902);
nor UO_411 (O_411,N_2954,N_2905);
nand UO_412 (O_412,N_2946,N_2993);
and UO_413 (O_413,N_2923,N_2992);
nor UO_414 (O_414,N_2929,N_2996);
or UO_415 (O_415,N_2990,N_2935);
nor UO_416 (O_416,N_2952,N_2921);
nand UO_417 (O_417,N_2996,N_2964);
and UO_418 (O_418,N_2954,N_2941);
and UO_419 (O_419,N_2972,N_2905);
nor UO_420 (O_420,N_2969,N_2949);
nor UO_421 (O_421,N_2997,N_2931);
or UO_422 (O_422,N_2963,N_2908);
or UO_423 (O_423,N_2926,N_2960);
nor UO_424 (O_424,N_2953,N_2990);
nor UO_425 (O_425,N_2935,N_2923);
and UO_426 (O_426,N_2957,N_2970);
or UO_427 (O_427,N_2994,N_2944);
or UO_428 (O_428,N_2948,N_2990);
or UO_429 (O_429,N_2907,N_2938);
xor UO_430 (O_430,N_2903,N_2993);
or UO_431 (O_431,N_2930,N_2985);
nand UO_432 (O_432,N_2916,N_2972);
and UO_433 (O_433,N_2979,N_2928);
and UO_434 (O_434,N_2973,N_2957);
or UO_435 (O_435,N_2993,N_2951);
and UO_436 (O_436,N_2969,N_2923);
or UO_437 (O_437,N_2970,N_2996);
or UO_438 (O_438,N_2958,N_2917);
and UO_439 (O_439,N_2991,N_2925);
or UO_440 (O_440,N_2988,N_2993);
or UO_441 (O_441,N_2990,N_2920);
or UO_442 (O_442,N_2930,N_2983);
nand UO_443 (O_443,N_2994,N_2997);
and UO_444 (O_444,N_2909,N_2940);
nand UO_445 (O_445,N_2963,N_2973);
nand UO_446 (O_446,N_2962,N_2973);
nand UO_447 (O_447,N_2949,N_2991);
nor UO_448 (O_448,N_2982,N_2960);
or UO_449 (O_449,N_2902,N_2945);
nand UO_450 (O_450,N_2967,N_2917);
nand UO_451 (O_451,N_2916,N_2980);
and UO_452 (O_452,N_2908,N_2970);
nand UO_453 (O_453,N_2925,N_2939);
or UO_454 (O_454,N_2972,N_2990);
nand UO_455 (O_455,N_2901,N_2905);
and UO_456 (O_456,N_2947,N_2936);
nor UO_457 (O_457,N_2909,N_2904);
or UO_458 (O_458,N_2907,N_2952);
and UO_459 (O_459,N_2935,N_2981);
or UO_460 (O_460,N_2959,N_2987);
and UO_461 (O_461,N_2903,N_2915);
nand UO_462 (O_462,N_2932,N_2969);
and UO_463 (O_463,N_2907,N_2926);
nand UO_464 (O_464,N_2936,N_2981);
nand UO_465 (O_465,N_2912,N_2937);
nor UO_466 (O_466,N_2984,N_2904);
or UO_467 (O_467,N_2985,N_2980);
nand UO_468 (O_468,N_2945,N_2933);
nor UO_469 (O_469,N_2986,N_2927);
and UO_470 (O_470,N_2978,N_2940);
nand UO_471 (O_471,N_2934,N_2919);
and UO_472 (O_472,N_2927,N_2917);
and UO_473 (O_473,N_2988,N_2973);
nand UO_474 (O_474,N_2902,N_2903);
or UO_475 (O_475,N_2977,N_2933);
nand UO_476 (O_476,N_2952,N_2955);
nor UO_477 (O_477,N_2987,N_2937);
or UO_478 (O_478,N_2991,N_2930);
nor UO_479 (O_479,N_2903,N_2901);
or UO_480 (O_480,N_2993,N_2974);
nor UO_481 (O_481,N_2904,N_2917);
and UO_482 (O_482,N_2983,N_2925);
nor UO_483 (O_483,N_2977,N_2959);
and UO_484 (O_484,N_2967,N_2986);
nand UO_485 (O_485,N_2980,N_2970);
and UO_486 (O_486,N_2973,N_2944);
nand UO_487 (O_487,N_2900,N_2950);
or UO_488 (O_488,N_2958,N_2944);
and UO_489 (O_489,N_2955,N_2915);
nor UO_490 (O_490,N_2994,N_2901);
xor UO_491 (O_491,N_2991,N_2970);
and UO_492 (O_492,N_2958,N_2913);
nor UO_493 (O_493,N_2939,N_2935);
or UO_494 (O_494,N_2918,N_2978);
or UO_495 (O_495,N_2939,N_2915);
nand UO_496 (O_496,N_2958,N_2959);
nor UO_497 (O_497,N_2917,N_2973);
and UO_498 (O_498,N_2958,N_2916);
nor UO_499 (O_499,N_2962,N_2959);
endmodule